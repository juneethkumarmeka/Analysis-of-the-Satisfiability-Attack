module basic_2500_25000_3000_4_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18801,N_18802,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18939,N_18940,N_18941,N_18942,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18965,N_18966,N_18967,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19119,N_19120,N_19121,N_19122,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19600,N_19601,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19838,N_19839,N_19840,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20074,N_20075,N_20076,N_20077,N_20078,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20662,N_20663,N_20664,N_20665,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20944,N_20945,N_20946,N_20948,N_20950,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21070,N_21071,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21279,N_21280,N_21282,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21417,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21576,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21754,N_21755,N_21756,N_21757,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21818,N_21819,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22045,N_22046,N_22047,N_22048,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22250,N_22251,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22552,N_22553,N_22554,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22574,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23249,N_23250,N_23251,N_23252,N_23253,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23357,N_23358,N_23359,N_23360,N_23362,N_23364,N_23365,N_23366,N_23367,N_23368,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23390,N_23391,N_23392,N_23393,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23571,N_23572,N_23573,N_23574,N_23575,N_23577,N_23578,N_23579,N_23580,N_23581,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23706,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24118,N_24120,N_24121,N_24122,N_24123,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24209,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24300,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24319,N_24320,N_24321,N_24322,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24472,N_24473,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24576,N_24577,N_24578,N_24579,N_24581,N_24582,N_24583,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24642,N_24643,N_24644,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24776,N_24777,N_24778,N_24779,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1631,In_303);
nand U1 (N_1,In_2223,In_1471);
nand U2 (N_2,In_725,In_1397);
nand U3 (N_3,In_2441,In_2058);
nor U4 (N_4,In_567,In_450);
nand U5 (N_5,In_1080,In_40);
nand U6 (N_6,In_1548,In_1799);
and U7 (N_7,In_2099,In_1567);
and U8 (N_8,In_448,In_261);
nor U9 (N_9,In_1501,In_2287);
and U10 (N_10,In_1193,In_601);
nand U11 (N_11,In_131,In_1026);
or U12 (N_12,In_263,In_1381);
nand U13 (N_13,In_2045,In_489);
or U14 (N_14,In_1691,In_629);
nand U15 (N_15,In_1335,In_1771);
and U16 (N_16,In_476,In_292);
and U17 (N_17,In_1334,In_1173);
nand U18 (N_18,In_198,In_1769);
nand U19 (N_19,In_279,In_1185);
nand U20 (N_20,In_511,In_1070);
and U21 (N_21,In_1086,In_434);
and U22 (N_22,In_2197,In_777);
and U23 (N_23,In_523,In_955);
or U24 (N_24,In_1667,In_453);
or U25 (N_25,In_2331,In_2440);
and U26 (N_26,In_861,In_2327);
or U27 (N_27,In_1260,In_789);
and U28 (N_28,In_2211,In_902);
and U29 (N_29,In_1916,In_1433);
nand U30 (N_30,In_965,In_1187);
nand U31 (N_31,In_319,In_176);
and U32 (N_32,In_2401,In_560);
nor U33 (N_33,In_9,In_2356);
and U34 (N_34,In_2003,In_1459);
nor U35 (N_35,In_1581,In_1475);
nor U36 (N_36,In_1216,In_1431);
nor U37 (N_37,In_1784,In_149);
nand U38 (N_38,In_77,In_1764);
nor U39 (N_39,In_1956,In_467);
nor U40 (N_40,In_158,In_1557);
and U41 (N_41,In_934,In_1103);
nor U42 (N_42,In_1361,In_178);
and U43 (N_43,In_2173,In_1255);
nor U44 (N_44,In_1698,In_1790);
nor U45 (N_45,In_45,In_689);
nor U46 (N_46,In_1109,In_1474);
nor U47 (N_47,In_962,In_16);
or U48 (N_48,In_1296,In_2130);
xnor U49 (N_49,In_1283,In_2227);
and U50 (N_50,In_1354,In_2494);
nand U51 (N_51,In_2113,In_2009);
and U52 (N_52,In_1546,In_1344);
or U53 (N_53,In_2177,In_2449);
and U54 (N_54,In_623,In_889);
and U55 (N_55,In_868,In_1214);
and U56 (N_56,In_1179,In_1785);
or U57 (N_57,In_1676,In_1521);
or U58 (N_58,In_415,In_2493);
and U59 (N_59,In_2210,In_713);
or U60 (N_60,In_99,In_1419);
and U61 (N_61,In_21,In_990);
nand U62 (N_62,In_1097,In_1838);
nor U63 (N_63,In_549,In_1774);
nand U64 (N_64,In_1262,In_2396);
and U65 (N_65,In_690,In_2395);
and U66 (N_66,In_508,In_852);
xor U67 (N_67,In_2106,In_203);
and U68 (N_68,In_1966,In_1904);
nor U69 (N_69,In_614,In_483);
nor U70 (N_70,In_1378,In_1299);
and U71 (N_71,In_546,In_738);
nor U72 (N_72,In_520,In_799);
and U73 (N_73,In_1908,In_225);
nor U74 (N_74,In_2178,In_1719);
nor U75 (N_75,In_2139,In_2434);
nor U76 (N_76,In_1509,In_2151);
nor U77 (N_77,In_1887,In_1245);
or U78 (N_78,In_269,In_264);
and U79 (N_79,In_1540,In_648);
nor U80 (N_80,In_1266,In_1543);
nand U81 (N_81,In_1484,In_2275);
nand U82 (N_82,In_1519,In_1999);
nand U83 (N_83,In_181,In_222);
nor U84 (N_84,In_1244,In_218);
nand U85 (N_85,In_1695,In_907);
and U86 (N_86,In_1039,In_1977);
nor U87 (N_87,In_968,In_1886);
nor U88 (N_88,In_2219,In_1280);
and U89 (N_89,In_82,In_1294);
and U90 (N_90,In_1043,In_374);
and U91 (N_91,In_1563,In_2246);
or U92 (N_92,In_573,In_2377);
and U93 (N_93,In_204,In_446);
and U94 (N_94,In_233,In_1541);
and U95 (N_95,In_2324,In_2161);
nor U96 (N_96,In_1578,In_1851);
nand U97 (N_97,In_228,In_2482);
or U98 (N_98,In_1879,In_111);
and U99 (N_99,In_819,In_1278);
and U100 (N_100,In_2014,In_437);
or U101 (N_101,In_1135,In_1826);
or U102 (N_102,In_1493,In_991);
or U103 (N_103,In_1289,In_932);
or U104 (N_104,In_1709,In_668);
nor U105 (N_105,In_1095,In_2008);
and U106 (N_106,In_1951,In_212);
or U107 (N_107,In_1456,In_897);
and U108 (N_108,In_1846,In_1057);
and U109 (N_109,In_719,In_786);
nand U110 (N_110,In_2148,In_997);
nor U111 (N_111,In_57,In_1352);
or U112 (N_112,In_698,In_1812);
nand U113 (N_113,In_2262,In_2047);
nand U114 (N_114,In_357,In_186);
nand U115 (N_115,In_1842,In_1045);
nor U116 (N_116,In_1365,In_1576);
and U117 (N_117,In_1938,In_1082);
nand U118 (N_118,In_1840,In_1226);
or U119 (N_119,In_2230,In_2436);
nand U120 (N_120,In_818,In_2424);
nand U121 (N_121,In_2084,In_704);
or U122 (N_122,In_1268,In_973);
nand U123 (N_123,In_436,In_1735);
and U124 (N_124,In_433,In_2306);
or U125 (N_125,In_1110,In_324);
or U126 (N_126,In_1834,In_253);
and U127 (N_127,In_68,In_1229);
and U128 (N_128,In_1473,In_827);
and U129 (N_129,In_496,In_885);
nor U130 (N_130,In_2183,In_1559);
nand U131 (N_131,In_46,In_1894);
or U132 (N_132,In_2267,In_1787);
and U133 (N_133,In_1041,In_1011);
or U134 (N_134,In_1297,In_1892);
nor U135 (N_135,In_2248,In_503);
or U136 (N_136,In_71,In_1169);
nand U137 (N_137,In_1801,In_958);
nand U138 (N_138,In_1428,In_2114);
and U139 (N_139,In_556,In_53);
nand U140 (N_140,In_1034,In_1412);
or U141 (N_141,In_947,In_2066);
or U142 (N_142,In_217,In_2477);
or U143 (N_143,In_1596,In_321);
or U144 (N_144,In_238,In_382);
and U145 (N_145,In_2476,In_1944);
and U146 (N_146,In_553,In_1706);
and U147 (N_147,In_1393,In_380);
and U148 (N_148,In_1724,In_1154);
xnor U149 (N_149,In_1228,In_1816);
xor U150 (N_150,In_557,In_2038);
and U151 (N_151,In_1194,In_2000);
and U152 (N_152,In_1092,In_1233);
or U153 (N_153,In_1783,In_26);
nor U154 (N_154,In_900,In_837);
and U155 (N_155,In_2149,In_1128);
nor U156 (N_156,In_569,In_1516);
and U157 (N_157,In_908,In_2204);
and U158 (N_158,In_1176,In_2015);
and U159 (N_159,In_379,In_442);
xor U160 (N_160,In_2442,In_2315);
nor U161 (N_161,In_2174,In_384);
or U162 (N_162,In_2072,In_262);
nor U163 (N_163,In_1482,In_1742);
or U164 (N_164,In_2200,In_440);
nand U165 (N_165,In_2206,In_665);
nor U166 (N_166,In_1775,In_1220);
nand U167 (N_167,In_235,In_518);
or U168 (N_168,In_543,In_140);
or U169 (N_169,In_419,In_1403);
nand U170 (N_170,In_65,In_456);
nor U171 (N_171,In_2495,In_2354);
nor U172 (N_172,In_529,In_697);
nand U173 (N_173,In_764,In_540);
nor U174 (N_174,In_1534,In_147);
and U175 (N_175,In_1860,In_1111);
nand U176 (N_176,In_676,In_1313);
nor U177 (N_177,In_477,In_1167);
and U178 (N_178,In_1942,In_1981);
nand U179 (N_179,In_2329,In_585);
nor U180 (N_180,In_1374,In_609);
or U181 (N_181,In_1978,In_1457);
nor U182 (N_182,In_322,In_1995);
nor U183 (N_183,In_527,In_780);
nor U184 (N_184,In_1394,In_2128);
nand U185 (N_185,In_1224,In_245);
or U186 (N_186,In_2484,In_485);
nand U187 (N_187,In_1672,In_2092);
nand U188 (N_188,In_320,In_353);
nand U189 (N_189,In_1902,In_922);
or U190 (N_190,In_452,In_405);
and U191 (N_191,In_693,In_1003);
nand U192 (N_192,In_63,In_715);
and U193 (N_193,In_27,In_2368);
nor U194 (N_194,In_1300,In_414);
and U195 (N_195,In_917,In_2328);
or U196 (N_196,In_125,In_1654);
nor U197 (N_197,In_1808,In_1796);
or U198 (N_198,In_1642,In_839);
nand U199 (N_199,In_1186,In_1531);
nand U200 (N_200,In_1539,In_1325);
nor U201 (N_201,In_1630,In_363);
or U202 (N_202,In_2403,In_950);
nand U203 (N_203,In_1196,In_1212);
or U204 (N_204,In_2202,In_132);
nor U205 (N_205,In_2428,In_1051);
nand U206 (N_206,In_621,In_1637);
nor U207 (N_207,In_1148,In_1592);
nor U208 (N_208,In_1614,In_1588);
nor U209 (N_209,In_1303,In_1207);
and U210 (N_210,In_1157,In_492);
or U211 (N_211,In_413,In_175);
xor U212 (N_212,In_1740,In_1001);
and U213 (N_213,In_1249,In_1213);
nand U214 (N_214,In_2480,In_1726);
and U215 (N_215,In_784,In_2089);
or U216 (N_216,In_162,In_255);
or U217 (N_217,In_1275,In_202);
nand U218 (N_218,In_2029,In_2060);
nor U219 (N_219,In_2242,In_1217);
and U220 (N_220,In_924,In_1006);
nor U221 (N_221,In_1991,In_1858);
or U222 (N_222,In_887,In_936);
nand U223 (N_223,In_1124,In_367);
nor U224 (N_224,In_1651,In_74);
nand U225 (N_225,In_1119,In_570);
nor U226 (N_226,In_1499,In_333);
nand U227 (N_227,In_1989,In_873);
or U228 (N_228,In_2192,In_2125);
nand U229 (N_229,In_2413,In_2144);
and U230 (N_230,In_574,In_1583);
nor U231 (N_231,In_1091,In_291);
nor U232 (N_232,In_361,In_1505);
or U233 (N_233,In_960,In_1708);
nor U234 (N_234,In_551,In_1147);
and U235 (N_235,In_1702,In_2407);
or U236 (N_236,In_2470,In_1568);
and U237 (N_237,In_2111,In_1738);
or U238 (N_238,In_2102,In_2031);
nand U239 (N_239,In_2004,In_1199);
or U240 (N_240,In_1373,In_572);
or U241 (N_241,In_1237,In_1286);
nand U242 (N_242,In_2411,In_1472);
and U243 (N_243,In_2450,In_1321);
nor U244 (N_244,In_2108,In_660);
nand U245 (N_245,In_1416,In_770);
nor U246 (N_246,In_2237,In_2138);
nor U247 (N_247,In_2367,In_2313);
or U248 (N_248,In_154,In_2259);
nor U249 (N_249,In_334,In_1030);
nor U250 (N_250,In_1205,In_1360);
nor U251 (N_251,In_661,In_1112);
nand U252 (N_252,In_2446,In_1862);
nand U253 (N_253,In_1919,In_1754);
nand U254 (N_254,In_912,In_2425);
nand U255 (N_255,In_435,In_2293);
and U256 (N_256,In_344,In_1849);
nor U257 (N_257,In_519,In_387);
nor U258 (N_258,In_644,In_242);
or U259 (N_259,In_1158,In_1607);
nand U260 (N_260,In_1971,In_1551);
nor U261 (N_261,In_2002,In_1564);
nand U262 (N_262,In_1670,In_426);
nand U263 (N_263,In_1432,In_351);
nor U264 (N_264,In_4,In_270);
nor U265 (N_265,In_2245,In_248);
nor U266 (N_266,In_2453,In_684);
and U267 (N_267,In_308,In_317);
and U268 (N_268,In_1720,In_156);
nor U269 (N_269,In_1375,In_1830);
nor U270 (N_270,In_2117,In_2310);
nand U271 (N_271,In_365,In_612);
and U272 (N_272,In_25,In_1747);
nand U273 (N_273,In_1443,In_1079);
nor U274 (N_274,In_875,In_1678);
nor U275 (N_275,In_13,In_381);
or U276 (N_276,In_735,In_1671);
and U277 (N_277,In_402,In_832);
nor U278 (N_278,In_2188,In_2466);
nor U279 (N_279,In_964,In_1797);
and U280 (N_280,In_666,In_2147);
and U281 (N_281,In_58,In_1018);
and U282 (N_282,In_1714,In_2299);
or U283 (N_283,In_1666,In_1496);
or U284 (N_284,In_535,In_136);
or U285 (N_285,In_488,In_224);
and U286 (N_286,In_591,In_60);
or U287 (N_287,In_844,In_304);
or U288 (N_288,In_2392,In_1831);
nor U289 (N_289,In_946,In_1021);
nand U290 (N_290,In_672,In_107);
nand U291 (N_291,In_1138,In_1231);
or U292 (N_292,In_1175,In_1312);
nand U293 (N_293,In_695,In_2362);
nor U294 (N_294,In_701,In_298);
or U295 (N_295,In_1760,In_576);
nand U296 (N_296,In_1986,In_2349);
or U297 (N_297,In_169,In_2340);
nand U298 (N_298,In_2110,In_1096);
nor U299 (N_299,In_2120,In_1064);
nor U300 (N_300,In_2062,In_1259);
nand U301 (N_301,In_2376,In_1889);
or U302 (N_302,In_2228,In_241);
or U303 (N_303,In_191,In_935);
and U304 (N_304,In_368,In_2043);
nand U305 (N_305,In_2143,In_1813);
nand U306 (N_306,In_876,In_742);
nand U307 (N_307,In_1017,In_933);
nor U308 (N_308,In_1750,In_555);
nor U309 (N_309,In_345,In_2285);
nand U310 (N_310,In_438,In_1263);
nor U311 (N_311,In_1319,In_385);
or U312 (N_312,In_1730,In_1985);
nor U313 (N_313,In_208,In_1968);
and U314 (N_314,In_1716,In_685);
nand U315 (N_315,In_56,In_1298);
nor U316 (N_316,In_1005,In_1322);
and U317 (N_317,In_1446,In_1640);
and U318 (N_318,In_1932,In_256);
nand U319 (N_319,In_957,In_2071);
and U320 (N_320,In_1617,In_2104);
nand U321 (N_321,In_1125,In_2185);
nand U322 (N_322,In_487,In_1055);
nor U323 (N_323,In_920,In_1227);
or U324 (N_324,In_1538,In_901);
and U325 (N_325,In_811,In_1087);
nor U326 (N_326,In_812,In_1940);
and U327 (N_327,In_2257,In_2079);
nand U328 (N_328,In_31,In_1483);
or U329 (N_329,In_372,In_775);
nor U330 (N_330,In_2271,In_458);
nor U331 (N_331,In_1625,In_1022);
nand U332 (N_332,In_1903,In_772);
nand U333 (N_333,In_1060,In_1414);
and U334 (N_334,In_377,In_1643);
or U335 (N_335,In_2443,In_1946);
or U336 (N_336,In_2418,In_1779);
and U337 (N_337,In_788,In_637);
or U338 (N_338,In_1172,In_1409);
nor U339 (N_339,In_2412,In_2105);
and U340 (N_340,In_653,In_8);
and U341 (N_341,In_753,In_785);
and U342 (N_342,In_544,In_2055);
and U343 (N_343,In_1565,In_2260);
nor U344 (N_344,In_2321,In_2168);
nor U345 (N_345,In_878,In_100);
nand U346 (N_346,In_2420,In_2046);
nor U347 (N_347,In_2498,In_1770);
and U348 (N_348,In_664,In_2053);
and U349 (N_349,In_1608,In_2006);
nor U350 (N_350,In_445,In_674);
nand U351 (N_351,In_2157,In_195);
or U352 (N_352,In_79,In_1434);
nand U353 (N_353,In_1960,In_1897);
nor U354 (N_354,In_2318,In_1009);
or U355 (N_355,In_1837,In_1350);
and U356 (N_356,In_2253,In_761);
or U357 (N_357,In_2135,In_307);
nand U358 (N_358,In_1983,In_1177);
nor U359 (N_359,In_2346,In_454);
and U360 (N_360,In_825,In_1390);
or U361 (N_361,In_2387,In_170);
nand U362 (N_362,In_1878,In_1604);
nand U363 (N_363,In_575,In_1180);
and U364 (N_364,In_998,In_851);
nand U365 (N_365,In_823,In_2247);
or U366 (N_366,In_856,In_840);
or U367 (N_367,In_2437,In_2405);
and U368 (N_368,In_914,In_1852);
nor U369 (N_369,In_1000,In_1494);
or U370 (N_370,In_441,In_123);
and U371 (N_371,In_1054,In_2445);
nor U372 (N_372,In_1339,In_1282);
xor U373 (N_373,In_2308,In_148);
or U374 (N_374,In_1572,In_2369);
and U375 (N_375,In_1683,In_2037);
nor U376 (N_376,In_1669,In_1445);
nand U377 (N_377,In_1497,In_2464);
nand U378 (N_378,In_2086,In_160);
nand U379 (N_379,In_2217,In_550);
nor U380 (N_380,In_841,In_257);
nor U381 (N_381,In_1803,In_1257);
nand U382 (N_382,In_422,In_1533);
or U383 (N_383,In_266,In_707);
nand U384 (N_384,In_478,In_881);
nand U385 (N_385,In_1848,In_1100);
nor U386 (N_386,In_710,In_971);
and U387 (N_387,In_1662,In_632);
nor U388 (N_388,In_1418,In_466);
or U389 (N_389,In_15,In_213);
or U390 (N_390,In_499,In_1441);
nor U391 (N_391,In_1184,In_539);
nor U392 (N_392,In_1982,In_711);
nand U393 (N_393,In_2175,In_2077);
nand U394 (N_394,In_43,In_2316);
nand U395 (N_395,In_815,In_792);
or U396 (N_396,In_2064,In_1717);
and U397 (N_397,In_533,In_1686);
or U398 (N_398,In_1917,In_1198);
nand U399 (N_399,In_490,In_854);
nor U400 (N_400,In_2345,In_2456);
nor U401 (N_401,In_1363,In_81);
nand U402 (N_402,In_2468,In_11);
nand U403 (N_403,In_2007,In_699);
or U404 (N_404,In_2121,In_1700);
or U405 (N_405,In_12,In_462);
nor U406 (N_406,In_2309,In_1950);
nor U407 (N_407,In_2292,In_1859);
and U408 (N_408,In_1636,In_1072);
and U409 (N_409,In_2301,In_1014);
nor U410 (N_410,In_1411,In_619);
and U411 (N_411,In_2073,In_1274);
nor U412 (N_412,In_748,In_278);
or U413 (N_413,In_6,In_2300);
or U414 (N_414,In_1537,In_51);
nor U415 (N_415,In_1680,In_2052);
and U416 (N_416,In_2365,In_2155);
nor U417 (N_417,In_1346,In_2061);
nand U418 (N_418,In_2444,In_1211);
nor U419 (N_419,In_95,In_1906);
or U420 (N_420,In_1815,In_646);
and U421 (N_421,In_765,In_1468);
or U422 (N_422,In_2291,In_1032);
and U423 (N_423,In_2430,In_153);
nand U424 (N_424,In_1866,In_1115);
and U425 (N_425,In_444,In_196);
nor U426 (N_426,In_271,In_1911);
nor U427 (N_427,In_2010,In_1907);
nor U428 (N_428,In_247,In_758);
nor U429 (N_429,In_729,In_1491);
or U430 (N_430,In_297,In_1454);
nand U431 (N_431,In_999,In_117);
nand U432 (N_432,In_1663,In_1800);
nand U433 (N_433,In_1593,In_211);
or U434 (N_434,In_2485,In_1687);
nor U435 (N_435,In_1697,In_1798);
and U436 (N_436,In_2457,In_1063);
nor U437 (N_437,In_622,In_1256);
and U438 (N_438,In_1290,In_299);
nand U439 (N_439,In_1447,In_2330);
and U440 (N_440,In_1398,In_55);
or U441 (N_441,In_952,In_1914);
or U442 (N_442,In_2112,In_326);
and U443 (N_443,In_2098,In_1477);
nor U444 (N_444,In_1439,In_1379);
or U445 (N_445,In_842,In_1622);
or U446 (N_446,In_756,In_78);
and U447 (N_447,In_1078,In_328);
and U448 (N_448,In_87,In_2091);
nand U449 (N_449,In_386,In_1107);
or U450 (N_450,In_1139,In_530);
xnor U451 (N_451,In_1577,In_250);
nor U452 (N_452,In_904,In_717);
or U453 (N_453,In_2279,In_1131);
xnor U454 (N_454,In_1618,In_774);
nor U455 (N_455,In_1466,In_1033);
nor U456 (N_456,In_2491,In_2471);
nand U457 (N_457,In_2481,In_517);
and U458 (N_458,In_2193,In_524);
and U459 (N_459,In_2421,In_391);
nor U460 (N_460,In_2252,In_1969);
or U461 (N_461,In_987,In_1470);
nand U462 (N_462,In_229,In_1552);
and U463 (N_463,In_1182,In_930);
nor U464 (N_464,In_1421,In_1273);
or U465 (N_465,In_1550,In_669);
and U466 (N_466,In_358,In_1802);
nand U467 (N_467,In_44,In_2284);
nor U468 (N_468,In_1395,In_2207);
or U469 (N_469,In_1710,In_1143);
or U470 (N_470,In_1238,In_128);
nor U471 (N_471,In_1122,In_598);
and U472 (N_472,In_1646,In_73);
nand U473 (N_473,In_1913,In_2129);
or U474 (N_474,In_1804,In_400);
nor U475 (N_475,In_610,In_2017);
nand U476 (N_476,In_2496,In_1674);
nand U477 (N_477,In_24,In_2410);
nor U478 (N_478,In_2265,In_2069);
and U479 (N_479,In_1929,In_2243);
nand U480 (N_480,In_165,In_2090);
and U481 (N_481,In_1504,In_1461);
or U482 (N_482,In_1314,In_2272);
or U483 (N_483,In_583,In_431);
and U484 (N_484,In_70,In_1423);
and U485 (N_485,In_631,In_1874);
or U486 (N_486,In_2294,In_2153);
nor U487 (N_487,In_2458,In_2063);
nor U488 (N_488,In_867,In_953);
nand U489 (N_489,In_460,In_1073);
and U490 (N_490,In_145,In_349);
nor U491 (N_491,In_663,In_2281);
nand U492 (N_492,In_749,In_1518);
or U493 (N_493,In_1959,In_36);
nor U494 (N_494,In_337,In_85);
and U495 (N_495,In_677,In_853);
or U496 (N_496,In_769,In_1495);
and U497 (N_497,In_986,In_421);
and U498 (N_498,In_923,In_1141);
or U499 (N_499,In_1606,In_2163);
nand U500 (N_500,In_2134,In_2371);
nor U501 (N_501,In_804,In_268);
or U502 (N_502,In_1150,In_1727);
or U503 (N_503,In_1655,In_1376);
and U504 (N_504,In_1701,In_1258);
and U505 (N_505,In_398,In_1025);
nand U506 (N_506,In_1992,In_432);
or U507 (N_507,In_1881,In_1164);
or U508 (N_508,In_2370,In_2295);
and U509 (N_509,In_1965,In_721);
and U510 (N_510,In_192,In_2338);
nor U511 (N_511,In_1529,In_64);
or U512 (N_512,In_1668,In_1463);
nand U513 (N_513,In_2431,In_2042);
and U514 (N_514,In_1309,In_548);
and U515 (N_515,In_2320,In_159);
or U516 (N_516,In_1053,In_2082);
or U517 (N_517,In_2028,In_504);
or U518 (N_518,In_1225,In_656);
and U519 (N_519,In_884,In_243);
nand U520 (N_520,In_1042,In_396);
or U521 (N_521,In_1062,In_103);
and U522 (N_522,In_172,In_2335);
and U523 (N_523,In_747,In_532);
or U524 (N_524,In_1190,In_1828);
or U525 (N_525,In_2158,In_1440);
or U526 (N_526,In_1219,In_667);
or U527 (N_527,In_586,In_926);
or U528 (N_528,In_940,In_88);
nor U529 (N_529,In_1382,In_782);
or U530 (N_530,In_223,In_634);
nand U531 (N_531,In_1704,In_135);
nor U532 (N_532,In_1340,In_29);
or U533 (N_533,In_1085,In_2085);
nor U534 (N_534,In_1284,In_272);
or U535 (N_535,In_2166,In_2162);
or U536 (N_536,In_1641,In_210);
nand U537 (N_537,In_1739,In_1031);
and U538 (N_538,In_17,In_2036);
nand U539 (N_539,In_311,In_1023);
nand U540 (N_540,In_1613,In_1571);
nor U541 (N_541,In_1331,In_1647);
or U542 (N_542,In_2499,In_2039);
nand U543 (N_543,In_403,In_507);
or U544 (N_544,In_2176,In_2132);
or U545 (N_545,In_113,In_1380);
or U546 (N_546,In_2234,In_2027);
nand U547 (N_547,In_2189,In_2273);
and U548 (N_548,In_984,In_509);
or U549 (N_549,In_1920,In_1629);
and U550 (N_550,In_118,In_2263);
nand U551 (N_551,In_1424,In_356);
or U552 (N_552,In_820,In_2032);
or U553 (N_553,In_671,In_536);
nand U554 (N_554,In_1012,In_69);
nand U555 (N_555,In_393,In_1357);
or U556 (N_556,In_2429,In_428);
nand U557 (N_557,In_497,In_1696);
and U558 (N_558,In_903,In_910);
or U559 (N_559,In_945,In_143);
and U560 (N_560,In_52,In_2026);
and U561 (N_561,In_723,In_209);
nand U562 (N_562,In_1272,In_1963);
nor U563 (N_563,In_833,In_2323);
or U564 (N_564,In_1925,In_394);
nand U565 (N_565,In_1635,In_2359);
or U566 (N_566,In_590,In_2363);
or U567 (N_567,In_805,In_993);
and U568 (N_568,In_1694,In_471);
nor U569 (N_569,In_801,In_1949);
or U570 (N_570,In_906,In_1612);
nand U571 (N_571,In_1067,In_472);
and U572 (N_572,In_1876,In_331);
and U573 (N_573,In_1234,In_407);
nand U574 (N_574,In_2332,In_1984);
nor U575 (N_575,In_2297,In_139);
or U576 (N_576,In_1961,In_726);
and U577 (N_577,In_97,In_1728);
and U578 (N_578,In_1855,In_768);
or U579 (N_579,In_1809,In_1203);
nand U580 (N_580,In_1628,In_1508);
or U581 (N_581,In_1104,In_2404);
nand U582 (N_582,In_2304,In_2081);
nand U583 (N_583,In_1029,In_893);
or U584 (N_584,In_2278,In_2416);
nor U585 (N_585,In_2013,In_1383);
nor U586 (N_586,In_397,In_565);
nor U587 (N_587,In_708,In_1435);
and U588 (N_588,In_762,In_1870);
nor U589 (N_589,In_1899,In_2286);
and U590 (N_590,In_751,In_2075);
nor U591 (N_591,In_1208,In_647);
and U592 (N_592,In_2402,In_872);
nand U593 (N_593,In_2463,In_1332);
nand U594 (N_594,In_846,In_2447);
nor U595 (N_595,In_1677,In_1480);
and U596 (N_596,In_745,In_869);
nor U597 (N_597,In_1755,In_1453);
nand U598 (N_598,In_2136,In_2422);
or U599 (N_599,In_1088,In_1718);
and U600 (N_600,In_1161,In_1118);
and U601 (N_601,In_1648,In_1699);
nor U602 (N_602,In_890,In_352);
nor U603 (N_603,In_1239,In_401);
and U604 (N_604,In_1108,In_2214);
or U605 (N_605,In_2373,In_2465);
nor U606 (N_606,In_1598,In_1478);
nand U607 (N_607,In_977,In_227);
nand U608 (N_608,In_891,In_231);
and U609 (N_609,In_994,In_187);
nor U610 (N_610,In_286,In_2094);
nor U611 (N_611,In_120,In_182);
and U612 (N_612,In_2238,In_966);
or U613 (N_613,In_339,In_1449);
nor U614 (N_614,In_681,In_96);
and U615 (N_615,In_1292,In_2400);
or U616 (N_616,In_1140,In_1362);
nor U617 (N_617,In_164,In_254);
nor U618 (N_618,In_2030,In_643);
and U619 (N_619,In_92,In_2325);
or U620 (N_620,In_1895,In_937);
nor U621 (N_621,In_1980,In_1707);
nor U622 (N_622,In_939,In_1780);
and U623 (N_623,In_2474,In_2357);
and U624 (N_624,In_455,In_19);
nor U625 (N_625,In_2488,In_578);
or U626 (N_626,In_1074,In_949);
nand U627 (N_627,In_151,In_327);
and U628 (N_628,In_2251,In_1355);
and U629 (N_629,In_680,In_581);
nand U630 (N_630,In_67,In_137);
nand U631 (N_631,In_1392,In_1910);
nand U632 (N_632,In_563,In_1988);
nand U633 (N_633,In_2317,In_2380);
nand U634 (N_634,In_1044,In_709);
or U635 (N_635,In_2068,In_658);
or U636 (N_636,In_2483,In_838);
nor U637 (N_637,In_1287,In_1582);
nand U638 (N_638,In_411,In_892);
nand U639 (N_639,In_338,In_1500);
and U640 (N_640,In_537,In_2388);
nand U641 (N_641,In_564,In_1271);
or U642 (N_642,In_1868,In_1048);
and U643 (N_643,In_2433,In_599);
nor U644 (N_644,In_1767,In_1737);
or U645 (N_645,In_412,In_425);
or U646 (N_646,In_2415,In_1430);
or U647 (N_647,In_1144,In_896);
nor U648 (N_648,In_1372,In_898);
and U649 (N_649,In_1936,In_1133);
nand U650 (N_650,In_1781,In_2366);
or U651 (N_651,In_1345,In_1885);
and U652 (N_652,In_2384,In_1330);
and U653 (N_653,In_1389,In_670);
nor U654 (N_654,In_944,In_2351);
or U655 (N_655,In_959,In_1240);
or U656 (N_656,In_929,In_972);
and U657 (N_657,In_2288,In_615);
nand U658 (N_658,In_1276,In_1488);
nor U659 (N_659,In_2093,In_1869);
nor U660 (N_660,In_1427,In_1594);
and U661 (N_661,In_457,In_1083);
and U662 (N_662,In_595,In_1438);
and U663 (N_663,In_350,In_1713);
or U664 (N_664,In_114,In_2201);
and U665 (N_665,In_2435,In_985);
or U666 (N_666,In_2167,In_1326);
nor U667 (N_667,In_1391,In_1444);
and U668 (N_668,In_1269,In_2393);
nor U669 (N_669,In_2419,In_1285);
nor U670 (N_670,In_1997,In_461);
or U671 (N_671,In_173,In_2012);
nor U672 (N_672,In_1821,In_20);
or U673 (N_673,In_577,In_757);
or U674 (N_674,In_1099,In_1587);
or U675 (N_675,In_655,In_309);
and U676 (N_676,In_1254,In_275);
nand U677 (N_677,In_163,In_1310);
and U678 (N_678,In_2460,In_1805);
and U679 (N_679,In_915,In_482);
nand U680 (N_680,In_2191,In_1134);
or U681 (N_681,In_1328,In_850);
nor U682 (N_682,In_2195,In_2205);
nor U683 (N_683,In_251,In_2140);
xnor U684 (N_684,In_1232,In_2360);
and U685 (N_685,In_625,In_2254);
nor U686 (N_686,In_1777,In_325);
and U687 (N_687,In_1998,In_2239);
nor U688 (N_688,In_102,In_1132);
and U689 (N_689,In_1820,In_650);
and U690 (N_690,In_2255,In_1120);
nor U691 (N_691,In_2146,In_1673);
nand U692 (N_692,In_318,In_127);
or U693 (N_693,In_1952,In_1329);
and U694 (N_694,In_1306,In_475);
or U695 (N_695,In_1554,In_371);
and U696 (N_696,In_1010,In_755);
xnor U697 (N_697,In_486,In_1915);
nor U698 (N_698,In_39,In_1723);
or U699 (N_699,In_879,In_1145);
or U700 (N_700,In_10,In_1008);
and U701 (N_701,In_2221,In_983);
and U702 (N_702,In_1602,In_1945);
or U703 (N_703,In_720,In_1151);
nor U704 (N_704,In_1358,In_863);
nor U705 (N_705,In_2137,In_1342);
and U706 (N_706,In_1832,In_722);
nor U707 (N_707,In_888,In_829);
or U708 (N_708,In_406,In_2005);
or U709 (N_709,In_1758,In_179);
nor U710 (N_710,In_313,In_1349);
nand U711 (N_711,In_1974,In_604);
or U712 (N_712,In_1442,In_305);
or U713 (N_713,In_568,In_733);
nor U714 (N_714,In_1890,In_30);
or U715 (N_715,In_1941,In_817);
and U716 (N_716,In_1658,In_1528);
or U717 (N_717,In_1307,In_718);
nor U718 (N_718,In_1202,In_2180);
nor U719 (N_719,In_1705,In_1102);
and U720 (N_720,In_547,In_1101);
and U721 (N_721,In_849,In_18);
and U722 (N_722,In_617,In_542);
nor U723 (N_723,In_1996,In_2215);
and U724 (N_724,In_280,In_1437);
or U725 (N_725,In_2383,In_2187);
or U726 (N_726,In_1388,In_1749);
and U727 (N_727,In_793,In_1734);
nor U728 (N_728,In_2198,In_2312);
nand U729 (N_729,In_541,In_956);
and U730 (N_730,In_1279,In_2124);
nor U731 (N_731,In_284,In_86);
nor U732 (N_732,In_963,In_252);
nand U733 (N_733,In_2472,In_1729);
nor U734 (N_734,In_1489,In_2172);
and U735 (N_735,In_1341,In_2427);
and U736 (N_736,In_806,In_1241);
or U737 (N_737,In_37,In_552);
and U738 (N_738,In_1356,In_1338);
and U739 (N_739,In_1377,In_2080);
or U740 (N_740,In_1002,In_822);
nor U741 (N_741,In_2269,In_290);
nor U742 (N_742,In_588,In_686);
or U743 (N_743,In_1649,In_2226);
and U744 (N_744,In_2492,In_141);
or U745 (N_745,In_1311,In_94);
or U746 (N_746,In_1609,In_1733);
nand U747 (N_747,In_1270,In_2385);
and U748 (N_748,In_285,In_1506);
or U749 (N_749,In_1512,In_146);
nand U750 (N_750,In_2341,In_174);
nand U751 (N_751,In_559,In_142);
and U752 (N_752,In_494,In_1865);
and U753 (N_753,In_1603,In_1317);
and U754 (N_754,In_809,In_1530);
and U755 (N_755,In_2133,In_104);
nor U756 (N_756,In_2070,In_161);
and U757 (N_757,In_2067,In_388);
xnor U758 (N_758,In_1450,In_787);
nor U759 (N_759,In_627,In_183);
or U760 (N_760,In_1975,In_1793);
or U761 (N_761,In_1569,In_2044);
or U762 (N_762,In_230,In_1465);
and U763 (N_763,In_115,In_2109);
or U764 (N_764,In_1833,In_1933);
or U765 (N_765,In_2344,In_1027);
or U766 (N_766,In_1261,In_2);
nor U767 (N_767,In_607,In_1656);
nor U768 (N_768,In_2049,In_2001);
nand U769 (N_769,In_1215,In_2229);
nor U770 (N_770,In_692,In_1861);
and U771 (N_771,In_1152,In_1050);
nor U772 (N_772,In_961,In_1544);
and U773 (N_773,In_1399,In_1458);
and U774 (N_774,In_1084,In_899);
nor U775 (N_775,In_516,In_293);
nor U776 (N_776,In_1819,In_534);
nor U777 (N_777,In_2322,In_2115);
or U778 (N_778,In_600,In_925);
nor U779 (N_779,In_2241,In_193);
nor U780 (N_780,In_1515,In_1685);
nand U781 (N_781,In_831,In_724);
or U782 (N_782,In_1049,In_1586);
or U783 (N_783,In_427,In_1850);
and U784 (N_784,In_808,In_728);
or U785 (N_785,In_355,In_1451);
nor U786 (N_786,In_1056,In_2194);
nand U787 (N_787,In_566,In_2479);
nand U788 (N_788,In_866,In_1841);
and U789 (N_789,In_2342,In_592);
or U790 (N_790,In_1924,In_2451);
and U791 (N_791,In_2289,In_696);
or U792 (N_792,In_54,In_240);
nand U793 (N_793,In_199,In_459);
nor U794 (N_794,In_249,In_1327);
and U795 (N_795,In_1763,In_2347);
and U796 (N_796,In_2196,In_2350);
or U797 (N_797,In_2448,In_1632);
and U798 (N_798,In_468,In_2222);
and U799 (N_799,In_651,In_122);
or U800 (N_800,In_731,In_1318);
nor U801 (N_801,In_1759,In_1660);
xnor U802 (N_802,In_525,In_1736);
nor U803 (N_803,In_214,In_1600);
nor U804 (N_804,In_613,In_206);
nand U805 (N_805,In_855,In_2182);
or U806 (N_806,In_2164,In_702);
nand U807 (N_807,In_1081,In_1368);
nand U808 (N_808,In_232,In_1829);
and U809 (N_809,In_754,In_2209);
and U810 (N_810,In_1425,In_980);
and U811 (N_811,In_66,In_981);
and U812 (N_812,In_1511,In_1221);
and U813 (N_813,In_2298,In_1302);
nor U814 (N_814,In_1137,In_1794);
and U815 (N_815,In_2467,In_943);
or U816 (N_816,In_1864,In_1591);
nor U817 (N_817,In_1408,In_1746);
nor U818 (N_818,In_1448,In_616);
and U819 (N_819,In_2409,In_783);
or U820 (N_820,In_1007,In_369);
nand U821 (N_821,In_948,In_1953);
or U822 (N_822,In_1856,In_447);
nor U823 (N_823,In_1575,In_347);
or U824 (N_824,In_1404,In_635);
nand U825 (N_825,In_265,In_2212);
and U826 (N_826,In_32,In_909);
nor U827 (N_827,In_1429,In_1013);
nor U828 (N_828,In_2033,In_1958);
or U829 (N_829,In_180,In_810);
and U830 (N_830,In_2156,In_1513);
or U831 (N_831,In_493,In_1127);
and U832 (N_832,In_329,In_2224);
and U833 (N_833,In_982,In_1822);
and U834 (N_834,In_2141,In_38);
and U835 (N_835,In_1201,In_636);
or U836 (N_836,In_1204,In_1693);
and U837 (N_837,In_642,In_2282);
and U838 (N_838,In_1934,In_979);
nand U839 (N_839,In_340,In_1597);
and U840 (N_840,In_860,In_1492);
and U841 (N_841,In_91,In_1210);
nand U842 (N_842,In_1170,In_1935);
nor U843 (N_843,In_1065,In_185);
and U844 (N_844,In_877,In_1028);
nor U845 (N_845,In_2216,In_1410);
nor U846 (N_846,In_2336,In_1153);
nand U847 (N_847,In_2054,In_1943);
or U848 (N_848,In_1930,In_1987);
and U849 (N_849,In_1047,In_1405);
nor U850 (N_850,In_1316,In_797);
nand U851 (N_851,In_1744,In_207);
nand U852 (N_852,In_390,In_1400);
nand U853 (N_853,In_260,In_639);
nand U854 (N_854,In_2199,In_376);
and U855 (N_855,In_221,In_2048);
and U856 (N_856,In_1366,In_359);
or U857 (N_857,In_1171,In_1301);
xor U858 (N_858,In_1748,In_538);
nor U859 (N_859,In_1873,In_2249);
or U860 (N_860,In_2326,In_2181);
or U861 (N_861,In_1016,In_3);
or U862 (N_862,In_2432,In_750);
and U863 (N_863,In_1615,In_1364);
or U864 (N_864,In_1420,In_1973);
or U865 (N_865,In_2119,In_2021);
or U866 (N_866,In_35,In_886);
or U867 (N_867,In_417,In_911);
nand U868 (N_868,In_597,In_2399);
nand U869 (N_869,In_2088,In_714);
nor U870 (N_870,In_1789,In_1896);
and U871 (N_871,In_894,In_124);
or U872 (N_872,In_760,In_1384);
and U873 (N_873,In_1288,In_1200);
and U874 (N_874,In_845,In_1703);
nand U875 (N_875,In_1192,In_2050);
or U876 (N_876,In_675,In_28);
or U877 (N_877,In_1645,In_1498);
nor U878 (N_878,In_2203,In_1562);
nand U879 (N_879,In_473,In_1954);
nor U880 (N_880,In_521,In_116);
nand U881 (N_881,In_362,In_194);
nor U882 (N_882,In_2179,In_989);
nand U883 (N_883,In_967,In_14);
nor U884 (N_884,In_1415,In_424);
and U885 (N_885,In_1639,In_1681);
nand U886 (N_886,In_1807,In_1333);
and U887 (N_887,In_1979,In_1555);
or U888 (N_888,In_2307,In_580);
and U889 (N_889,In_705,In_2264);
nor U890 (N_890,In_512,In_1788);
nand U891 (N_891,In_267,In_1634);
nand U892 (N_892,In_274,In_1659);
nand U893 (N_893,In_589,In_129);
and U894 (N_894,In_287,In_2097);
and U895 (N_895,In_1888,In_1126);
nor U896 (N_896,In_342,In_283);
nand U897 (N_897,In_2218,In_34);
nand U898 (N_898,In_294,In_2381);
nand U899 (N_899,In_1467,In_1967);
nor U900 (N_900,In_2100,In_2225);
or U901 (N_901,In_1955,In_155);
or U902 (N_902,In_430,In_2096);
nor U903 (N_903,In_1776,In_144);
or U904 (N_904,In_1166,In_618);
and U905 (N_905,In_928,In_1347);
and U906 (N_906,In_1653,In_1165);
nor U907 (N_907,In_2382,In_119);
and U908 (N_908,In_836,In_716);
nand U909 (N_909,In_871,In_1741);
nor U910 (N_910,In_1485,In_1665);
or U911 (N_911,In_226,In_528);
nor U912 (N_912,In_2378,In_157);
nand U913 (N_913,In_1690,In_1772);
nand U914 (N_914,In_420,In_1181);
nand U915 (N_915,In_2283,In_1481);
and U916 (N_916,In_1348,In_703);
and U917 (N_917,In_1035,In_1743);
or U918 (N_918,In_1523,In_2462);
or U919 (N_919,In_1019,In_740);
nand U920 (N_920,In_816,In_1197);
nor U921 (N_921,In_1545,In_741);
or U922 (N_922,In_150,In_1939);
nand U923 (N_923,In_767,In_2489);
nor U924 (N_924,In_399,In_469);
and U925 (N_925,In_659,In_883);
nand U926 (N_926,In_2302,In_1560);
nor U927 (N_927,In_1845,In_691);
xor U928 (N_928,In_1136,In_491);
nor U929 (N_929,In_449,In_1066);
and U930 (N_930,In_1370,In_410);
and U931 (N_931,In_1359,In_2150);
nor U932 (N_932,In_1058,In_649);
or U933 (N_933,In_2353,In_2040);
and U934 (N_934,In_1059,In_220);
nor U935 (N_935,In_795,In_1757);
or U936 (N_936,In_188,In_1123);
nand U937 (N_937,In_1195,In_2116);
or U938 (N_938,In_2469,In_1526);
and U939 (N_939,In_638,In_366);
and U940 (N_940,In_1305,In_330);
nor U941 (N_941,In_1517,In_1657);
nand U942 (N_942,In_443,In_913);
and U943 (N_943,In_582,In_1579);
nor U944 (N_944,In_2256,In_2408);
and U945 (N_945,In_1209,In_281);
nand U946 (N_946,In_824,In_992);
nor U947 (N_947,In_1682,In_273);
and U948 (N_948,In_2473,In_1993);
and U949 (N_949,In_439,In_2426);
and U950 (N_950,In_931,In_974);
nor U951 (N_951,In_2490,In_1661);
nand U952 (N_952,In_662,In_1778);
nor U953 (N_953,In_2319,In_1462);
or U954 (N_954,In_1753,In_1623);
nand U955 (N_955,In_1711,In_1223);
nor U956 (N_956,In_969,In_1937);
nand U957 (N_957,In_1121,In_168);
and U958 (N_958,In_593,In_1206);
nor U959 (N_959,In_2364,In_2171);
and U960 (N_960,In_640,In_1163);
nand U961 (N_961,In_288,In_2059);
or U962 (N_962,In_2389,In_184);
and U963 (N_963,In_101,In_41);
and U964 (N_964,In_1323,In_2074);
and U965 (N_965,In_1964,In_1542);
nor U966 (N_966,In_501,In_2145);
or U967 (N_967,In_90,In_33);
or U968 (N_968,In_1715,In_1839);
nand U969 (N_969,In_1684,In_1105);
and U970 (N_970,In_1912,In_236);
nor U971 (N_971,In_2452,In_348);
nand U972 (N_972,In_197,In_2277);
nand U973 (N_973,In_109,In_106);
nor U974 (N_974,In_423,In_1731);
or U975 (N_975,In_2303,In_1814);
or U976 (N_976,In_1004,In_1304);
nor U977 (N_977,In_2083,In_554);
nor U978 (N_978,In_1957,In_2334);
or U979 (N_979,In_1460,In_237);
and U980 (N_980,In_2280,In_1610);
nand U981 (N_981,In_1624,In_2414);
nor U982 (N_982,In_976,In_791);
or U983 (N_983,In_739,In_1590);
and U984 (N_984,In_1324,In_0);
nor U985 (N_985,In_1487,In_1644);
nor U986 (N_986,In_2296,In_2235);
or U987 (N_987,In_641,In_2095);
or U988 (N_988,In_289,In_1825);
nand U989 (N_989,In_2186,In_1926);
nand U990 (N_990,In_1069,In_130);
nand U991 (N_991,In_2348,In_1795);
and U992 (N_992,In_418,In_2379);
nand U993 (N_993,In_2486,In_2455);
nand U994 (N_994,In_1351,In_2220);
nor U995 (N_995,In_1527,In_50);
and U996 (N_996,In_1765,In_2078);
nor U997 (N_997,In_2261,In_2142);
or U998 (N_998,In_1129,In_880);
nor U999 (N_999,In_657,In_1371);
and U1000 (N_1000,In_1156,In_1510);
and U1001 (N_1001,In_620,In_1168);
or U1002 (N_1002,In_1584,In_2152);
and U1003 (N_1003,In_1502,In_216);
nand U1004 (N_1004,In_1162,In_1061);
or U1005 (N_1005,In_630,In_1626);
nand U1006 (N_1006,In_2118,In_1020);
or U1007 (N_1007,In_1619,In_1247);
nand U1008 (N_1008,In_2034,In_2159);
or U1009 (N_1009,In_688,In_771);
and U1010 (N_1010,In_1417,In_1792);
or U1011 (N_1011,In_1159,In_2170);
or U1012 (N_1012,In_978,In_1752);
and U1013 (N_1013,In_370,In_1455);
or U1014 (N_1014,In_1535,In_679);
nand U1015 (N_1015,In_470,In_451);
nor U1016 (N_1016,In_138,In_2035);
or U1017 (N_1017,In_1146,In_759);
and U1018 (N_1018,In_905,In_558);
nor U1019 (N_1019,In_495,In_1407);
and U1020 (N_1020,In_1871,In_1077);
and U1021 (N_1021,In_874,In_1267);
nor U1022 (N_1022,In_1621,In_2236);
or U1023 (N_1023,In_2391,In_752);
or U1024 (N_1024,In_954,In_2423);
or U1025 (N_1025,In_2011,In_5);
nor U1026 (N_1026,In_1464,In_364);
nand U1027 (N_1027,In_828,In_1452);
nor U1028 (N_1028,In_1675,In_1337);
and U1029 (N_1029,In_807,In_1627);
nand U1030 (N_1030,In_465,In_847);
nand U1031 (N_1031,In_98,In_1252);
or U1032 (N_1032,In_1406,In_1847);
nor U1033 (N_1033,In_2065,In_995);
or U1034 (N_1034,In_1343,In_526);
or U1035 (N_1035,In_2244,In_1863);
nor U1036 (N_1036,In_2190,In_1923);
or U1037 (N_1037,In_1265,In_859);
nor U1038 (N_1038,In_1823,In_171);
and U1039 (N_1039,In_2024,In_938);
or U1040 (N_1040,In_1692,In_1558);
and U1041 (N_1041,In_1525,In_857);
or U1042 (N_1042,In_778,In_481);
nand U1043 (N_1043,In_1253,In_49);
and U1044 (N_1044,In_1222,In_1507);
or U1045 (N_1045,In_1573,In_1522);
xnor U1046 (N_1046,In_2016,In_1422);
and U1047 (N_1047,In_1514,In_712);
and U1048 (N_1048,In_919,In_1503);
or U1049 (N_1049,In_1264,In_61);
nor U1050 (N_1050,In_2107,In_2497);
and U1051 (N_1051,In_803,In_1191);
nand U1052 (N_1052,In_295,In_1490);
and U1053 (N_1053,In_678,In_1549);
nor U1054 (N_1054,In_1570,In_895);
or U1055 (N_1055,In_1725,In_282);
nand U1056 (N_1056,In_1402,In_802);
nor U1057 (N_1057,In_1246,In_343);
and U1058 (N_1058,In_596,In_796);
or U1059 (N_1059,In_927,In_744);
and U1060 (N_1060,In_975,In_258);
and U1061 (N_1061,In_1293,In_2123);
or U1062 (N_1062,In_730,In_1117);
nor U1063 (N_1063,In_316,In_1867);
nand U1064 (N_1064,In_1745,In_1556);
nor U1065 (N_1065,In_2025,In_244);
nand U1066 (N_1066,In_1396,In_766);
nor U1067 (N_1067,In_276,In_882);
and U1068 (N_1068,In_2461,In_310);
nand U1069 (N_1069,In_734,In_2018);
or U1070 (N_1070,In_743,In_2305);
and U1071 (N_1071,In_1599,In_2386);
nand U1072 (N_1072,In_341,In_166);
nand U1073 (N_1073,In_1601,In_498);
nand U1074 (N_1074,In_1574,In_1611);
nor U1075 (N_1075,In_1251,In_1761);
and U1076 (N_1076,In_2361,In_112);
nand U1077 (N_1077,In_1036,In_1106);
nor U1078 (N_1078,In_1880,In_1901);
nand U1079 (N_1079,In_1972,In_1843);
and U1080 (N_1080,In_300,In_673);
and U1081 (N_1081,In_1068,In_2459);
nor U1082 (N_1082,In_346,In_2022);
xnor U1083 (N_1083,In_416,In_1075);
nand U1084 (N_1084,In_1155,In_1854);
and U1085 (N_1085,In_312,In_1291);
and U1086 (N_1086,In_1835,In_2337);
or U1087 (N_1087,In_1605,In_474);
xnor U1088 (N_1088,In_126,In_1962);
nor U1089 (N_1089,In_246,In_727);
and U1090 (N_1090,In_200,In_1336);
and U1091 (N_1091,In_1090,In_813);
nand U1092 (N_1092,In_2439,In_1773);
nand U1093 (N_1093,In_315,In_219);
and U1094 (N_1094,In_1386,In_513);
nand U1095 (N_1095,In_395,In_1469);
and U1096 (N_1096,In_1928,In_332);
or U1097 (N_1097,In_354,In_259);
and U1098 (N_1098,In_835,In_918);
or U1099 (N_1099,In_514,In_502);
xnor U1100 (N_1100,In_1038,In_652);
nand U1101 (N_1101,In_1921,In_479);
xor U1102 (N_1102,In_737,In_89);
and U1103 (N_1103,In_916,In_1218);
nor U1104 (N_1104,In_1883,In_409);
and U1105 (N_1105,In_505,In_1189);
and U1106 (N_1106,In_2406,In_134);
and U1107 (N_1107,In_2311,In_2390);
and U1108 (N_1108,In_2051,In_1436);
or U1109 (N_1109,In_1638,In_2231);
nor U1110 (N_1110,In_1040,In_190);
nor U1111 (N_1111,In_335,In_1827);
or U1112 (N_1112,In_826,In_1948);
and U1113 (N_1113,In_239,In_1142);
xnor U1114 (N_1114,In_531,In_105);
or U1115 (N_1115,In_1836,In_2268);
nor U1116 (N_1116,In_1712,In_108);
nor U1117 (N_1117,In_2394,In_1884);
and U1118 (N_1118,In_389,In_205);
nand U1119 (N_1119,In_1616,In_1990);
nor U1120 (N_1120,In_645,In_858);
nand U1121 (N_1121,In_1235,In_314);
nor U1122 (N_1122,In_378,In_1242);
nor U1123 (N_1123,In_1385,In_2122);
and U1124 (N_1124,In_746,In_215);
nor U1125 (N_1125,In_996,In_1098);
nand U1126 (N_1126,In_1689,In_1905);
or U1127 (N_1127,In_2314,In_865);
nor U1128 (N_1128,In_1188,In_2475);
and U1129 (N_1129,In_1918,In_683);
or U1130 (N_1130,In_1116,In_2372);
and U1131 (N_1131,In_1791,In_773);
or U1132 (N_1132,In_1320,In_602);
nand U1133 (N_1133,In_1532,In_624);
and U1134 (N_1134,In_83,In_1633);
nor U1135 (N_1135,In_633,In_814);
or U1136 (N_1136,In_7,In_1688);
or U1137 (N_1137,In_1093,In_848);
or U1138 (N_1138,In_201,In_62);
and U1139 (N_1139,In_1113,In_1178);
nor U1140 (N_1140,In_22,In_1553);
and U1141 (N_1141,In_694,In_2233);
nand U1142 (N_1142,In_1768,In_603);
or U1143 (N_1143,In_167,In_628);
nand U1144 (N_1144,In_133,In_429);
or U1145 (N_1145,In_2397,In_2240);
nor U1146 (N_1146,In_189,In_47);
nor U1147 (N_1147,In_2258,In_1250);
and U1148 (N_1148,In_1353,In_522);
nand U1149 (N_1149,In_2352,In_1762);
nand U1150 (N_1150,In_1585,In_2131);
and U1151 (N_1151,In_1536,In_373);
nor U1152 (N_1152,In_561,In_80);
and U1153 (N_1153,In_484,In_1806);
nor U1154 (N_1154,In_1308,In_2041);
nor U1155 (N_1155,In_383,In_152);
or U1156 (N_1156,In_2087,In_1580);
and U1157 (N_1157,In_2019,In_584);
and U1158 (N_1158,In_2250,In_2023);
xnor U1159 (N_1159,In_1931,In_1922);
nand U1160 (N_1160,In_2454,In_1947);
nand U1161 (N_1161,In_1909,In_2169);
nor U1162 (N_1162,In_1520,In_84);
or U1163 (N_1163,In_1369,In_1811);
nand U1164 (N_1164,In_515,In_830);
or U1165 (N_1165,In_121,In_800);
or U1166 (N_1166,In_654,In_2343);
or U1167 (N_1167,In_2375,In_1872);
or U1168 (N_1168,In_2057,In_1566);
and U1169 (N_1169,In_545,In_942);
and U1170 (N_1170,In_1174,In_1248);
nand U1171 (N_1171,In_1230,In_1089);
or U1172 (N_1172,In_1524,In_941);
nand U1173 (N_1173,In_1732,In_1824);
and U1174 (N_1174,In_23,In_1766);
nand U1175 (N_1175,In_408,In_1882);
or U1176 (N_1176,In_2208,In_1620);
or U1177 (N_1177,In_1877,In_1547);
nor U1178 (N_1178,In_1160,In_72);
and U1179 (N_1179,In_500,In_862);
nand U1180 (N_1180,In_2274,In_2266);
or U1181 (N_1181,In_2154,In_2213);
and U1182 (N_1182,In_779,In_2374);
or U1183 (N_1183,In_1076,In_1751);
nor U1184 (N_1184,In_763,In_1898);
nand U1185 (N_1185,In_870,In_336);
nand U1186 (N_1186,In_579,In_1722);
or U1187 (N_1187,In_864,In_2076);
or U1188 (N_1188,In_301,In_392);
nor U1189 (N_1189,In_1857,In_2276);
and U1190 (N_1190,In_296,In_1114);
nand U1191 (N_1191,In_2290,In_776);
nand U1192 (N_1192,In_1130,In_2339);
or U1193 (N_1193,In_1,In_1927);
or U1194 (N_1194,In_1052,In_794);
and U1195 (N_1195,In_1650,In_75);
and U1196 (N_1196,In_790,In_1476);
and U1197 (N_1197,In_1295,In_606);
nor U1198 (N_1198,In_2232,In_1664);
nor U1199 (N_1199,In_736,In_277);
nand U1200 (N_1200,In_1786,In_2417);
and U1201 (N_1201,In_988,In_234);
and U1202 (N_1202,In_177,In_302);
and U1203 (N_1203,In_360,In_687);
nand U1204 (N_1204,In_2333,In_1891);
nor U1205 (N_1205,In_1236,In_587);
or U1206 (N_1206,In_2126,In_834);
nor U1207 (N_1207,In_1015,In_951);
and U1208 (N_1208,In_1994,In_76);
nand U1209 (N_1209,In_1046,In_1900);
nor U1210 (N_1210,In_1486,In_2101);
nor U1211 (N_1211,In_594,In_562);
or U1212 (N_1212,In_682,In_1401);
nand U1213 (N_1213,In_970,In_464);
xnor U1214 (N_1214,In_1893,In_1367);
nor U1215 (N_1215,In_821,In_463);
nand U1216 (N_1216,In_1243,In_1024);
nand U1217 (N_1217,In_2478,In_1426);
or U1218 (N_1218,In_306,In_2355);
nor U1219 (N_1219,In_1183,In_611);
or U1220 (N_1220,In_1595,In_2160);
or U1221 (N_1221,In_1875,In_110);
nor U1222 (N_1222,In_1281,In_375);
xor U1223 (N_1223,In_608,In_93);
nor U1224 (N_1224,In_1589,In_1652);
and U1225 (N_1225,In_1149,In_781);
nand U1226 (N_1226,In_1094,In_1818);
or U1227 (N_1227,In_1277,In_48);
and U1228 (N_1228,In_1976,In_700);
nand U1229 (N_1229,In_2056,In_1970);
and U1230 (N_1230,In_2184,In_2270);
or U1231 (N_1231,In_732,In_1721);
nand U1232 (N_1232,In_1413,In_626);
nor U1233 (N_1233,In_42,In_2438);
nor U1234 (N_1234,In_59,In_921);
and U1235 (N_1235,In_798,In_2487);
or U1236 (N_1236,In_506,In_1844);
and U1237 (N_1237,In_605,In_1387);
nor U1238 (N_1238,In_2020,In_1817);
or U1239 (N_1239,In_2127,In_1756);
or U1240 (N_1240,In_571,In_480);
nand U1241 (N_1241,In_1853,In_843);
nor U1242 (N_1242,In_323,In_2103);
nand U1243 (N_1243,In_404,In_1315);
and U1244 (N_1244,In_2398,In_706);
nor U1245 (N_1245,In_2358,In_1037);
and U1246 (N_1246,In_510,In_2165);
or U1247 (N_1247,In_1561,In_1479);
nor U1248 (N_1248,In_1071,In_1782);
and U1249 (N_1249,In_1679,In_1810);
and U1250 (N_1250,In_175,In_1477);
nand U1251 (N_1251,In_2236,In_736);
nor U1252 (N_1252,In_294,In_1369);
nor U1253 (N_1253,In_419,In_931);
xor U1254 (N_1254,In_1582,In_1760);
nor U1255 (N_1255,In_2149,In_1668);
nor U1256 (N_1256,In_2109,In_799);
nand U1257 (N_1257,In_2408,In_2268);
or U1258 (N_1258,In_1218,In_554);
and U1259 (N_1259,In_799,In_557);
and U1260 (N_1260,In_1370,In_119);
or U1261 (N_1261,In_162,In_1622);
nand U1262 (N_1262,In_1718,In_600);
nand U1263 (N_1263,In_939,In_30);
or U1264 (N_1264,In_1389,In_1632);
nor U1265 (N_1265,In_1937,In_2333);
or U1266 (N_1266,In_791,In_876);
or U1267 (N_1267,In_2441,In_211);
nand U1268 (N_1268,In_768,In_2269);
or U1269 (N_1269,In_92,In_271);
or U1270 (N_1270,In_464,In_1118);
or U1271 (N_1271,In_1708,In_1056);
nor U1272 (N_1272,In_918,In_1371);
nand U1273 (N_1273,In_830,In_1890);
and U1274 (N_1274,In_2464,In_1613);
nand U1275 (N_1275,In_2184,In_2014);
and U1276 (N_1276,In_119,In_905);
nand U1277 (N_1277,In_1002,In_720);
or U1278 (N_1278,In_278,In_1728);
or U1279 (N_1279,In_1603,In_1167);
nor U1280 (N_1280,In_416,In_1860);
nand U1281 (N_1281,In_113,In_2469);
nand U1282 (N_1282,In_2183,In_959);
and U1283 (N_1283,In_245,In_1323);
nor U1284 (N_1284,In_2241,In_631);
and U1285 (N_1285,In_1726,In_174);
and U1286 (N_1286,In_1731,In_1423);
nand U1287 (N_1287,In_257,In_1793);
and U1288 (N_1288,In_2248,In_1012);
and U1289 (N_1289,In_218,In_1845);
nor U1290 (N_1290,In_1728,In_820);
nand U1291 (N_1291,In_763,In_2343);
and U1292 (N_1292,In_876,In_1065);
and U1293 (N_1293,In_807,In_1915);
nor U1294 (N_1294,In_95,In_1941);
nor U1295 (N_1295,In_666,In_2124);
nor U1296 (N_1296,In_1651,In_1239);
nand U1297 (N_1297,In_803,In_922);
or U1298 (N_1298,In_574,In_1295);
nor U1299 (N_1299,In_1021,In_422);
and U1300 (N_1300,In_748,In_377);
or U1301 (N_1301,In_614,In_1195);
or U1302 (N_1302,In_2494,In_1284);
xnor U1303 (N_1303,In_117,In_2001);
nor U1304 (N_1304,In_445,In_1376);
or U1305 (N_1305,In_2326,In_1436);
and U1306 (N_1306,In_1169,In_1548);
nand U1307 (N_1307,In_1506,In_1603);
and U1308 (N_1308,In_2454,In_587);
nor U1309 (N_1309,In_1968,In_2337);
nand U1310 (N_1310,In_711,In_1742);
and U1311 (N_1311,In_1763,In_1323);
or U1312 (N_1312,In_36,In_1901);
and U1313 (N_1313,In_1584,In_657);
and U1314 (N_1314,In_540,In_2021);
and U1315 (N_1315,In_1237,In_422);
nand U1316 (N_1316,In_1111,In_371);
and U1317 (N_1317,In_140,In_394);
and U1318 (N_1318,In_2176,In_1896);
or U1319 (N_1319,In_2067,In_2300);
nand U1320 (N_1320,In_651,In_1694);
and U1321 (N_1321,In_2071,In_1267);
or U1322 (N_1322,In_1307,In_1814);
and U1323 (N_1323,In_88,In_227);
or U1324 (N_1324,In_1489,In_1605);
or U1325 (N_1325,In_922,In_41);
or U1326 (N_1326,In_2302,In_1801);
nand U1327 (N_1327,In_1794,In_331);
nand U1328 (N_1328,In_292,In_2477);
or U1329 (N_1329,In_94,In_1943);
nor U1330 (N_1330,In_946,In_2484);
or U1331 (N_1331,In_1357,In_2159);
nand U1332 (N_1332,In_1701,In_1483);
or U1333 (N_1333,In_1872,In_1251);
and U1334 (N_1334,In_2318,In_2141);
and U1335 (N_1335,In_196,In_2397);
nand U1336 (N_1336,In_2406,In_1680);
nand U1337 (N_1337,In_1488,In_1315);
nand U1338 (N_1338,In_1544,In_1784);
xnor U1339 (N_1339,In_1019,In_2443);
nand U1340 (N_1340,In_1456,In_121);
or U1341 (N_1341,In_2268,In_182);
or U1342 (N_1342,In_618,In_1802);
and U1343 (N_1343,In_1789,In_739);
nor U1344 (N_1344,In_1260,In_467);
nor U1345 (N_1345,In_1458,In_1359);
nand U1346 (N_1346,In_268,In_978);
or U1347 (N_1347,In_1669,In_2056);
nor U1348 (N_1348,In_806,In_1496);
and U1349 (N_1349,In_1585,In_1154);
or U1350 (N_1350,In_1492,In_2008);
nand U1351 (N_1351,In_32,In_2288);
nor U1352 (N_1352,In_208,In_1075);
or U1353 (N_1353,In_1424,In_2010);
nand U1354 (N_1354,In_2195,In_2382);
nand U1355 (N_1355,In_1983,In_1237);
nor U1356 (N_1356,In_526,In_2202);
or U1357 (N_1357,In_1740,In_597);
and U1358 (N_1358,In_2497,In_910);
nand U1359 (N_1359,In_2,In_1188);
nor U1360 (N_1360,In_1872,In_1027);
and U1361 (N_1361,In_1509,In_1374);
and U1362 (N_1362,In_1490,In_2293);
nand U1363 (N_1363,In_2317,In_2276);
or U1364 (N_1364,In_2131,In_527);
nor U1365 (N_1365,In_2292,In_1210);
or U1366 (N_1366,In_1799,In_1063);
and U1367 (N_1367,In_2163,In_1206);
nor U1368 (N_1368,In_811,In_492);
nor U1369 (N_1369,In_705,In_2178);
and U1370 (N_1370,In_2146,In_1140);
or U1371 (N_1371,In_2294,In_2143);
or U1372 (N_1372,In_2072,In_2365);
or U1373 (N_1373,In_633,In_473);
or U1374 (N_1374,In_733,In_411);
nand U1375 (N_1375,In_1582,In_1118);
and U1376 (N_1376,In_40,In_566);
and U1377 (N_1377,In_2282,In_1298);
nor U1378 (N_1378,In_426,In_443);
and U1379 (N_1379,In_1621,In_2361);
nor U1380 (N_1380,In_1580,In_590);
or U1381 (N_1381,In_76,In_985);
nor U1382 (N_1382,In_93,In_267);
nor U1383 (N_1383,In_2153,In_468);
nand U1384 (N_1384,In_396,In_337);
nor U1385 (N_1385,In_1993,In_1827);
nor U1386 (N_1386,In_877,In_800);
nor U1387 (N_1387,In_2486,In_991);
and U1388 (N_1388,In_1573,In_840);
nand U1389 (N_1389,In_256,In_1024);
or U1390 (N_1390,In_1075,In_519);
or U1391 (N_1391,In_2282,In_633);
nand U1392 (N_1392,In_271,In_605);
nor U1393 (N_1393,In_1160,In_2312);
and U1394 (N_1394,In_1950,In_2417);
and U1395 (N_1395,In_322,In_335);
or U1396 (N_1396,In_1526,In_1484);
or U1397 (N_1397,In_1372,In_262);
or U1398 (N_1398,In_1650,In_1739);
or U1399 (N_1399,In_1502,In_1250);
nor U1400 (N_1400,In_1715,In_2110);
xor U1401 (N_1401,In_1254,In_946);
and U1402 (N_1402,In_2058,In_1673);
nor U1403 (N_1403,In_372,In_1838);
or U1404 (N_1404,In_724,In_2271);
or U1405 (N_1405,In_1451,In_77);
and U1406 (N_1406,In_556,In_519);
and U1407 (N_1407,In_1279,In_870);
nand U1408 (N_1408,In_1030,In_175);
and U1409 (N_1409,In_441,In_876);
nand U1410 (N_1410,In_1956,In_1466);
and U1411 (N_1411,In_1302,In_1814);
nand U1412 (N_1412,In_1589,In_579);
nand U1413 (N_1413,In_2332,In_1115);
nand U1414 (N_1414,In_2493,In_213);
and U1415 (N_1415,In_572,In_2193);
nor U1416 (N_1416,In_1505,In_2067);
or U1417 (N_1417,In_1063,In_2336);
nand U1418 (N_1418,In_758,In_160);
nor U1419 (N_1419,In_478,In_842);
nand U1420 (N_1420,In_1729,In_761);
and U1421 (N_1421,In_1280,In_2413);
and U1422 (N_1422,In_2374,In_1145);
and U1423 (N_1423,In_1679,In_1087);
nor U1424 (N_1424,In_2390,In_1022);
or U1425 (N_1425,In_2295,In_1395);
nor U1426 (N_1426,In_1393,In_2378);
and U1427 (N_1427,In_336,In_729);
and U1428 (N_1428,In_1624,In_414);
and U1429 (N_1429,In_1802,In_1294);
and U1430 (N_1430,In_1346,In_1500);
or U1431 (N_1431,In_1732,In_28);
nand U1432 (N_1432,In_1303,In_2434);
nand U1433 (N_1433,In_1498,In_1646);
nand U1434 (N_1434,In_572,In_2328);
nand U1435 (N_1435,In_581,In_788);
and U1436 (N_1436,In_2456,In_912);
nor U1437 (N_1437,In_150,In_1929);
nor U1438 (N_1438,In_2184,In_2254);
nand U1439 (N_1439,In_605,In_854);
or U1440 (N_1440,In_2258,In_529);
nand U1441 (N_1441,In_1735,In_809);
and U1442 (N_1442,In_378,In_1382);
nand U1443 (N_1443,In_1134,In_889);
nand U1444 (N_1444,In_1888,In_1063);
nand U1445 (N_1445,In_515,In_135);
or U1446 (N_1446,In_1964,In_1908);
nand U1447 (N_1447,In_2394,In_1154);
and U1448 (N_1448,In_569,In_874);
and U1449 (N_1449,In_1519,In_2408);
and U1450 (N_1450,In_1997,In_440);
and U1451 (N_1451,In_1382,In_79);
nor U1452 (N_1452,In_2146,In_45);
nand U1453 (N_1453,In_2161,In_538);
nand U1454 (N_1454,In_2238,In_281);
or U1455 (N_1455,In_2287,In_2465);
or U1456 (N_1456,In_1074,In_125);
nor U1457 (N_1457,In_767,In_2077);
or U1458 (N_1458,In_11,In_262);
and U1459 (N_1459,In_1435,In_187);
nand U1460 (N_1460,In_2318,In_248);
nor U1461 (N_1461,In_489,In_1461);
nand U1462 (N_1462,In_2149,In_1038);
xnor U1463 (N_1463,In_667,In_807);
or U1464 (N_1464,In_712,In_2409);
nand U1465 (N_1465,In_2267,In_338);
or U1466 (N_1466,In_1158,In_2221);
or U1467 (N_1467,In_118,In_2428);
nand U1468 (N_1468,In_1691,In_1745);
and U1469 (N_1469,In_267,In_2221);
or U1470 (N_1470,In_385,In_86);
nand U1471 (N_1471,In_645,In_1471);
xnor U1472 (N_1472,In_958,In_85);
or U1473 (N_1473,In_227,In_477);
and U1474 (N_1474,In_1365,In_1389);
nor U1475 (N_1475,In_265,In_2344);
or U1476 (N_1476,In_2117,In_2389);
or U1477 (N_1477,In_1041,In_536);
nor U1478 (N_1478,In_33,In_608);
nand U1479 (N_1479,In_1123,In_537);
and U1480 (N_1480,In_1000,In_939);
nor U1481 (N_1481,In_157,In_101);
and U1482 (N_1482,In_714,In_1998);
nand U1483 (N_1483,In_728,In_294);
or U1484 (N_1484,In_2477,In_1271);
or U1485 (N_1485,In_1615,In_1491);
and U1486 (N_1486,In_2149,In_1741);
or U1487 (N_1487,In_1521,In_662);
nand U1488 (N_1488,In_2389,In_504);
nor U1489 (N_1489,In_2342,In_2233);
or U1490 (N_1490,In_2255,In_2183);
and U1491 (N_1491,In_1338,In_236);
nand U1492 (N_1492,In_983,In_1621);
and U1493 (N_1493,In_2043,In_2133);
and U1494 (N_1494,In_1142,In_802);
nand U1495 (N_1495,In_759,In_1790);
and U1496 (N_1496,In_2102,In_2133);
nor U1497 (N_1497,In_541,In_1604);
or U1498 (N_1498,In_1674,In_1529);
and U1499 (N_1499,In_1513,In_1626);
or U1500 (N_1500,In_955,In_830);
nand U1501 (N_1501,In_1367,In_1114);
or U1502 (N_1502,In_1494,In_868);
nand U1503 (N_1503,In_33,In_1911);
and U1504 (N_1504,In_920,In_1867);
and U1505 (N_1505,In_672,In_847);
or U1506 (N_1506,In_674,In_1);
nand U1507 (N_1507,In_1556,In_1101);
and U1508 (N_1508,In_269,In_706);
or U1509 (N_1509,In_1255,In_125);
or U1510 (N_1510,In_382,In_2172);
nor U1511 (N_1511,In_1903,In_1684);
and U1512 (N_1512,In_1016,In_588);
and U1513 (N_1513,In_2376,In_2195);
nor U1514 (N_1514,In_793,In_510);
or U1515 (N_1515,In_1571,In_651);
or U1516 (N_1516,In_1706,In_182);
and U1517 (N_1517,In_2475,In_1882);
nand U1518 (N_1518,In_1396,In_2018);
or U1519 (N_1519,In_2459,In_652);
and U1520 (N_1520,In_2369,In_614);
or U1521 (N_1521,In_1203,In_2224);
nor U1522 (N_1522,In_2159,In_501);
nand U1523 (N_1523,In_517,In_1064);
and U1524 (N_1524,In_752,In_1045);
or U1525 (N_1525,In_1065,In_832);
or U1526 (N_1526,In_510,In_1804);
and U1527 (N_1527,In_1891,In_2118);
nor U1528 (N_1528,In_404,In_112);
or U1529 (N_1529,In_458,In_1125);
or U1530 (N_1530,In_31,In_1699);
nand U1531 (N_1531,In_1302,In_556);
or U1532 (N_1532,In_801,In_1591);
nand U1533 (N_1533,In_971,In_1868);
nor U1534 (N_1534,In_785,In_1864);
nand U1535 (N_1535,In_461,In_465);
and U1536 (N_1536,In_1095,In_1210);
nand U1537 (N_1537,In_319,In_1812);
or U1538 (N_1538,In_1031,In_1816);
or U1539 (N_1539,In_1764,In_1893);
nor U1540 (N_1540,In_1406,In_423);
nand U1541 (N_1541,In_2473,In_1060);
or U1542 (N_1542,In_2072,In_276);
nand U1543 (N_1543,In_1143,In_1561);
or U1544 (N_1544,In_1928,In_183);
nand U1545 (N_1545,In_776,In_262);
nand U1546 (N_1546,In_1681,In_200);
nor U1547 (N_1547,In_85,In_1743);
nor U1548 (N_1548,In_1001,In_1830);
or U1549 (N_1549,In_504,In_868);
nor U1550 (N_1550,In_2444,In_259);
nand U1551 (N_1551,In_1264,In_1389);
or U1552 (N_1552,In_2018,In_1891);
nand U1553 (N_1553,In_1300,In_2353);
or U1554 (N_1554,In_402,In_2091);
or U1555 (N_1555,In_2436,In_161);
nor U1556 (N_1556,In_1822,In_2372);
nor U1557 (N_1557,In_1819,In_1627);
or U1558 (N_1558,In_1968,In_1516);
nor U1559 (N_1559,In_598,In_1786);
nor U1560 (N_1560,In_1972,In_585);
nor U1561 (N_1561,In_2497,In_1605);
and U1562 (N_1562,In_2453,In_1138);
and U1563 (N_1563,In_301,In_138);
nand U1564 (N_1564,In_1517,In_1635);
and U1565 (N_1565,In_220,In_1154);
or U1566 (N_1566,In_1804,In_647);
nand U1567 (N_1567,In_2256,In_862);
nor U1568 (N_1568,In_374,In_2465);
or U1569 (N_1569,In_1077,In_250);
nand U1570 (N_1570,In_1554,In_1896);
nand U1571 (N_1571,In_2292,In_1368);
nor U1572 (N_1572,In_1165,In_725);
nor U1573 (N_1573,In_1383,In_52);
or U1574 (N_1574,In_1227,In_1895);
nor U1575 (N_1575,In_1132,In_553);
nor U1576 (N_1576,In_1970,In_349);
nand U1577 (N_1577,In_1989,In_660);
or U1578 (N_1578,In_502,In_879);
nand U1579 (N_1579,In_584,In_983);
nand U1580 (N_1580,In_754,In_621);
or U1581 (N_1581,In_483,In_2081);
and U1582 (N_1582,In_2419,In_570);
and U1583 (N_1583,In_618,In_1312);
or U1584 (N_1584,In_744,In_2331);
and U1585 (N_1585,In_1184,In_816);
or U1586 (N_1586,In_2299,In_253);
and U1587 (N_1587,In_1392,In_2290);
or U1588 (N_1588,In_7,In_527);
nor U1589 (N_1589,In_1008,In_229);
and U1590 (N_1590,In_2434,In_2343);
nand U1591 (N_1591,In_47,In_926);
nor U1592 (N_1592,In_2118,In_407);
and U1593 (N_1593,In_1967,In_138);
nand U1594 (N_1594,In_698,In_426);
nand U1595 (N_1595,In_403,In_704);
and U1596 (N_1596,In_436,In_1385);
or U1597 (N_1597,In_2177,In_757);
xor U1598 (N_1598,In_204,In_830);
nor U1599 (N_1599,In_1904,In_106);
nor U1600 (N_1600,In_275,In_55);
nand U1601 (N_1601,In_1842,In_1179);
nand U1602 (N_1602,In_1624,In_1496);
or U1603 (N_1603,In_2001,In_162);
nand U1604 (N_1604,In_621,In_2353);
or U1605 (N_1605,In_1233,In_1706);
and U1606 (N_1606,In_82,In_26);
and U1607 (N_1607,In_2307,In_103);
nor U1608 (N_1608,In_2434,In_1909);
nor U1609 (N_1609,In_2192,In_1586);
or U1610 (N_1610,In_2182,In_170);
nor U1611 (N_1611,In_672,In_349);
or U1612 (N_1612,In_946,In_2001);
and U1613 (N_1613,In_946,In_543);
and U1614 (N_1614,In_214,In_1459);
or U1615 (N_1615,In_2300,In_1491);
or U1616 (N_1616,In_697,In_1011);
nand U1617 (N_1617,In_435,In_1787);
and U1618 (N_1618,In_156,In_237);
nor U1619 (N_1619,In_1173,In_2202);
and U1620 (N_1620,In_990,In_1075);
and U1621 (N_1621,In_82,In_1652);
and U1622 (N_1622,In_877,In_1198);
nand U1623 (N_1623,In_1065,In_2138);
or U1624 (N_1624,In_1136,In_609);
or U1625 (N_1625,In_611,In_1203);
nor U1626 (N_1626,In_2160,In_538);
and U1627 (N_1627,In_2240,In_1940);
nand U1628 (N_1628,In_932,In_1482);
nor U1629 (N_1629,In_695,In_567);
nor U1630 (N_1630,In_586,In_1492);
and U1631 (N_1631,In_1910,In_1615);
and U1632 (N_1632,In_1630,In_2040);
nand U1633 (N_1633,In_2399,In_203);
nor U1634 (N_1634,In_2369,In_192);
and U1635 (N_1635,In_2211,In_1746);
or U1636 (N_1636,In_451,In_2158);
or U1637 (N_1637,In_2450,In_451);
and U1638 (N_1638,In_415,In_621);
nand U1639 (N_1639,In_854,In_899);
and U1640 (N_1640,In_99,In_1469);
and U1641 (N_1641,In_988,In_2401);
nand U1642 (N_1642,In_10,In_72);
or U1643 (N_1643,In_1812,In_1014);
nor U1644 (N_1644,In_1596,In_1104);
or U1645 (N_1645,In_332,In_1890);
nor U1646 (N_1646,In_2185,In_2365);
nand U1647 (N_1647,In_519,In_2287);
nor U1648 (N_1648,In_919,In_872);
nand U1649 (N_1649,In_1622,In_746);
nand U1650 (N_1650,In_276,In_745);
and U1651 (N_1651,In_1243,In_655);
or U1652 (N_1652,In_1869,In_796);
nand U1653 (N_1653,In_2230,In_2327);
nand U1654 (N_1654,In_1653,In_1890);
nor U1655 (N_1655,In_2397,In_304);
nor U1656 (N_1656,In_249,In_1004);
and U1657 (N_1657,In_1255,In_2244);
nor U1658 (N_1658,In_2440,In_361);
or U1659 (N_1659,In_2454,In_1669);
nor U1660 (N_1660,In_1664,In_1840);
or U1661 (N_1661,In_1051,In_247);
nand U1662 (N_1662,In_2223,In_340);
and U1663 (N_1663,In_1087,In_497);
nor U1664 (N_1664,In_2366,In_1618);
nor U1665 (N_1665,In_1706,In_1842);
nor U1666 (N_1666,In_897,In_1939);
nand U1667 (N_1667,In_936,In_2366);
and U1668 (N_1668,In_307,In_1445);
nand U1669 (N_1669,In_1585,In_1683);
and U1670 (N_1670,In_110,In_2175);
and U1671 (N_1671,In_2333,In_2457);
nand U1672 (N_1672,In_1602,In_1369);
and U1673 (N_1673,In_1598,In_2044);
nor U1674 (N_1674,In_866,In_124);
and U1675 (N_1675,In_498,In_9);
nor U1676 (N_1676,In_1,In_1311);
nor U1677 (N_1677,In_2106,In_1396);
nand U1678 (N_1678,In_1682,In_1797);
nand U1679 (N_1679,In_2402,In_95);
or U1680 (N_1680,In_1711,In_867);
or U1681 (N_1681,In_2361,In_1388);
and U1682 (N_1682,In_724,In_119);
or U1683 (N_1683,In_57,In_2209);
and U1684 (N_1684,In_184,In_156);
xor U1685 (N_1685,In_1110,In_1848);
or U1686 (N_1686,In_2310,In_1864);
nand U1687 (N_1687,In_1946,In_2053);
and U1688 (N_1688,In_1340,In_159);
nor U1689 (N_1689,In_835,In_409);
or U1690 (N_1690,In_71,In_365);
nand U1691 (N_1691,In_1325,In_915);
or U1692 (N_1692,In_1791,In_2346);
nand U1693 (N_1693,In_1731,In_1912);
nor U1694 (N_1694,In_18,In_50);
nor U1695 (N_1695,In_1718,In_2050);
or U1696 (N_1696,In_1513,In_1938);
and U1697 (N_1697,In_1022,In_1951);
nand U1698 (N_1698,In_1293,In_2299);
nor U1699 (N_1699,In_2482,In_1580);
and U1700 (N_1700,In_1332,In_785);
nand U1701 (N_1701,In_216,In_1492);
or U1702 (N_1702,In_931,In_629);
nor U1703 (N_1703,In_1500,In_238);
nand U1704 (N_1704,In_1584,In_996);
or U1705 (N_1705,In_700,In_1097);
and U1706 (N_1706,In_2320,In_392);
or U1707 (N_1707,In_368,In_764);
nand U1708 (N_1708,In_1384,In_363);
or U1709 (N_1709,In_1430,In_1746);
nor U1710 (N_1710,In_30,In_162);
nand U1711 (N_1711,In_652,In_1034);
xor U1712 (N_1712,In_2279,In_2061);
nor U1713 (N_1713,In_40,In_74);
nor U1714 (N_1714,In_255,In_1406);
nor U1715 (N_1715,In_1198,In_851);
nor U1716 (N_1716,In_1553,In_2076);
nor U1717 (N_1717,In_2023,In_871);
and U1718 (N_1718,In_465,In_568);
nor U1719 (N_1719,In_2422,In_2382);
or U1720 (N_1720,In_1665,In_1039);
nor U1721 (N_1721,In_1754,In_252);
or U1722 (N_1722,In_24,In_204);
or U1723 (N_1723,In_2278,In_613);
nand U1724 (N_1724,In_1228,In_1877);
nand U1725 (N_1725,In_342,In_1645);
nand U1726 (N_1726,In_841,In_1677);
nor U1727 (N_1727,In_1845,In_2443);
nand U1728 (N_1728,In_2324,In_461);
and U1729 (N_1729,In_2176,In_116);
nand U1730 (N_1730,In_105,In_2395);
or U1731 (N_1731,In_801,In_1593);
nor U1732 (N_1732,In_1358,In_2441);
and U1733 (N_1733,In_1876,In_196);
nand U1734 (N_1734,In_495,In_1758);
and U1735 (N_1735,In_474,In_86);
and U1736 (N_1736,In_2267,In_2075);
nor U1737 (N_1737,In_1079,In_49);
or U1738 (N_1738,In_379,In_155);
nand U1739 (N_1739,In_887,In_2208);
or U1740 (N_1740,In_2161,In_96);
and U1741 (N_1741,In_385,In_912);
and U1742 (N_1742,In_483,In_302);
and U1743 (N_1743,In_1841,In_54);
nand U1744 (N_1744,In_174,In_1248);
and U1745 (N_1745,In_1325,In_150);
and U1746 (N_1746,In_1942,In_1964);
or U1747 (N_1747,In_475,In_389);
or U1748 (N_1748,In_1554,In_2035);
or U1749 (N_1749,In_825,In_1476);
nand U1750 (N_1750,In_1611,In_1263);
nand U1751 (N_1751,In_615,In_21);
or U1752 (N_1752,In_2091,In_155);
or U1753 (N_1753,In_1708,In_1024);
nand U1754 (N_1754,In_1846,In_1000);
or U1755 (N_1755,In_954,In_1413);
nand U1756 (N_1756,In_1474,In_923);
and U1757 (N_1757,In_2131,In_2111);
nor U1758 (N_1758,In_78,In_1761);
and U1759 (N_1759,In_2249,In_1581);
or U1760 (N_1760,In_2095,In_2469);
nand U1761 (N_1761,In_2392,In_2012);
nand U1762 (N_1762,In_1029,In_1618);
and U1763 (N_1763,In_639,In_1500);
nor U1764 (N_1764,In_2000,In_2056);
nor U1765 (N_1765,In_2246,In_2054);
or U1766 (N_1766,In_1649,In_2429);
and U1767 (N_1767,In_199,In_1698);
and U1768 (N_1768,In_2491,In_1895);
nor U1769 (N_1769,In_1679,In_126);
or U1770 (N_1770,In_424,In_2330);
nor U1771 (N_1771,In_112,In_730);
xnor U1772 (N_1772,In_1498,In_701);
or U1773 (N_1773,In_2256,In_1787);
nand U1774 (N_1774,In_2369,In_892);
and U1775 (N_1775,In_808,In_1168);
nand U1776 (N_1776,In_327,In_709);
nor U1777 (N_1777,In_1815,In_1417);
or U1778 (N_1778,In_1022,In_434);
and U1779 (N_1779,In_2499,In_2058);
nand U1780 (N_1780,In_1439,In_533);
or U1781 (N_1781,In_2197,In_1603);
nand U1782 (N_1782,In_1456,In_1618);
nand U1783 (N_1783,In_2043,In_1527);
and U1784 (N_1784,In_919,In_2219);
nor U1785 (N_1785,In_1076,In_578);
nor U1786 (N_1786,In_669,In_791);
nor U1787 (N_1787,In_746,In_1556);
nand U1788 (N_1788,In_1472,In_1566);
nand U1789 (N_1789,In_255,In_1047);
nor U1790 (N_1790,In_787,In_1093);
nand U1791 (N_1791,In_631,In_1875);
or U1792 (N_1792,In_362,In_154);
nor U1793 (N_1793,In_808,In_137);
nand U1794 (N_1794,In_1629,In_611);
or U1795 (N_1795,In_1657,In_2169);
nor U1796 (N_1796,In_2109,In_1268);
nor U1797 (N_1797,In_861,In_1813);
or U1798 (N_1798,In_2335,In_931);
and U1799 (N_1799,In_1650,In_431);
and U1800 (N_1800,In_205,In_1392);
and U1801 (N_1801,In_684,In_1863);
nand U1802 (N_1802,In_2310,In_1321);
and U1803 (N_1803,In_1200,In_1679);
xor U1804 (N_1804,In_283,In_743);
nand U1805 (N_1805,In_1299,In_2064);
nor U1806 (N_1806,In_1994,In_2371);
and U1807 (N_1807,In_2185,In_1038);
nand U1808 (N_1808,In_1022,In_559);
nand U1809 (N_1809,In_146,In_1484);
nand U1810 (N_1810,In_2447,In_303);
nand U1811 (N_1811,In_21,In_518);
and U1812 (N_1812,In_2130,In_1726);
nand U1813 (N_1813,In_1385,In_1721);
or U1814 (N_1814,In_197,In_2252);
and U1815 (N_1815,In_1092,In_941);
or U1816 (N_1816,In_1428,In_1113);
or U1817 (N_1817,In_309,In_237);
nor U1818 (N_1818,In_1129,In_674);
nor U1819 (N_1819,In_1505,In_316);
or U1820 (N_1820,In_1344,In_2138);
or U1821 (N_1821,In_1363,In_1320);
and U1822 (N_1822,In_919,In_1755);
xnor U1823 (N_1823,In_2260,In_1309);
or U1824 (N_1824,In_1706,In_2077);
or U1825 (N_1825,In_1044,In_2251);
and U1826 (N_1826,In_2462,In_1298);
or U1827 (N_1827,In_1340,In_1707);
and U1828 (N_1828,In_189,In_527);
nor U1829 (N_1829,In_709,In_2003);
and U1830 (N_1830,In_1068,In_2015);
and U1831 (N_1831,In_1999,In_1513);
and U1832 (N_1832,In_1391,In_1903);
nand U1833 (N_1833,In_1392,In_2123);
or U1834 (N_1834,In_664,In_2220);
xnor U1835 (N_1835,In_968,In_2443);
nand U1836 (N_1836,In_1041,In_1228);
nor U1837 (N_1837,In_2423,In_1204);
or U1838 (N_1838,In_242,In_596);
or U1839 (N_1839,In_700,In_809);
nand U1840 (N_1840,In_1494,In_2334);
or U1841 (N_1841,In_1182,In_1025);
nor U1842 (N_1842,In_677,In_644);
nand U1843 (N_1843,In_1508,In_2338);
nor U1844 (N_1844,In_1839,In_542);
nand U1845 (N_1845,In_352,In_1368);
nor U1846 (N_1846,In_56,In_267);
nor U1847 (N_1847,In_1340,In_57);
nor U1848 (N_1848,In_1540,In_1529);
or U1849 (N_1849,In_546,In_589);
and U1850 (N_1850,In_2484,In_1680);
and U1851 (N_1851,In_1547,In_1978);
nand U1852 (N_1852,In_1867,In_230);
nor U1853 (N_1853,In_399,In_2198);
and U1854 (N_1854,In_1111,In_879);
nand U1855 (N_1855,In_2478,In_1719);
and U1856 (N_1856,In_2460,In_175);
or U1857 (N_1857,In_2250,In_231);
or U1858 (N_1858,In_841,In_231);
nand U1859 (N_1859,In_2147,In_458);
and U1860 (N_1860,In_1221,In_644);
and U1861 (N_1861,In_2221,In_1919);
and U1862 (N_1862,In_126,In_776);
nor U1863 (N_1863,In_1509,In_596);
or U1864 (N_1864,In_2387,In_699);
nand U1865 (N_1865,In_174,In_1188);
or U1866 (N_1866,In_820,In_2480);
and U1867 (N_1867,In_2150,In_99);
and U1868 (N_1868,In_477,In_1212);
and U1869 (N_1869,In_402,In_2418);
nand U1870 (N_1870,In_1906,In_949);
nand U1871 (N_1871,In_1134,In_2082);
and U1872 (N_1872,In_1068,In_1854);
or U1873 (N_1873,In_1160,In_344);
or U1874 (N_1874,In_17,In_1350);
nand U1875 (N_1875,In_662,In_2206);
and U1876 (N_1876,In_839,In_1230);
and U1877 (N_1877,In_124,In_2329);
nand U1878 (N_1878,In_800,In_1936);
or U1879 (N_1879,In_1579,In_646);
or U1880 (N_1880,In_467,In_2058);
and U1881 (N_1881,In_627,In_2328);
and U1882 (N_1882,In_508,In_2461);
nor U1883 (N_1883,In_242,In_1760);
or U1884 (N_1884,In_1866,In_2390);
or U1885 (N_1885,In_1170,In_2199);
nand U1886 (N_1886,In_2323,In_1575);
nand U1887 (N_1887,In_229,In_456);
and U1888 (N_1888,In_1687,In_1402);
or U1889 (N_1889,In_1088,In_105);
or U1890 (N_1890,In_2003,In_1123);
nor U1891 (N_1891,In_2130,In_167);
nand U1892 (N_1892,In_256,In_578);
nor U1893 (N_1893,In_100,In_1749);
nor U1894 (N_1894,In_2221,In_1079);
and U1895 (N_1895,In_1547,In_845);
nand U1896 (N_1896,In_2309,In_2193);
nor U1897 (N_1897,In_2404,In_1915);
nor U1898 (N_1898,In_1636,In_1204);
or U1899 (N_1899,In_1838,In_908);
and U1900 (N_1900,In_40,In_2376);
nor U1901 (N_1901,In_990,In_2272);
nor U1902 (N_1902,In_680,In_1958);
nand U1903 (N_1903,In_1171,In_542);
and U1904 (N_1904,In_450,In_1236);
or U1905 (N_1905,In_704,In_1021);
nor U1906 (N_1906,In_318,In_1606);
or U1907 (N_1907,In_1933,In_286);
and U1908 (N_1908,In_33,In_585);
and U1909 (N_1909,In_1956,In_341);
nand U1910 (N_1910,In_1371,In_1420);
nor U1911 (N_1911,In_1278,In_1064);
nor U1912 (N_1912,In_571,In_809);
and U1913 (N_1913,In_162,In_897);
nor U1914 (N_1914,In_1034,In_278);
and U1915 (N_1915,In_125,In_724);
nor U1916 (N_1916,In_1899,In_386);
and U1917 (N_1917,In_525,In_1957);
nor U1918 (N_1918,In_1906,In_2165);
or U1919 (N_1919,In_200,In_2173);
nor U1920 (N_1920,In_1843,In_2398);
nand U1921 (N_1921,In_876,In_1394);
and U1922 (N_1922,In_549,In_2460);
or U1923 (N_1923,In_809,In_532);
or U1924 (N_1924,In_382,In_741);
nor U1925 (N_1925,In_80,In_1615);
and U1926 (N_1926,In_2239,In_416);
nand U1927 (N_1927,In_452,In_1883);
nor U1928 (N_1928,In_187,In_1384);
or U1929 (N_1929,In_2129,In_699);
and U1930 (N_1930,In_2160,In_321);
nor U1931 (N_1931,In_1518,In_765);
or U1932 (N_1932,In_2373,In_119);
and U1933 (N_1933,In_1564,In_2240);
nor U1934 (N_1934,In_2306,In_307);
and U1935 (N_1935,In_957,In_929);
or U1936 (N_1936,In_587,In_2441);
and U1937 (N_1937,In_1622,In_1047);
and U1938 (N_1938,In_2007,In_278);
nor U1939 (N_1939,In_1119,In_354);
or U1940 (N_1940,In_357,In_237);
and U1941 (N_1941,In_468,In_245);
and U1942 (N_1942,In_1105,In_432);
or U1943 (N_1943,In_290,In_854);
nor U1944 (N_1944,In_1124,In_872);
and U1945 (N_1945,In_1947,In_1374);
nor U1946 (N_1946,In_1310,In_1115);
nand U1947 (N_1947,In_1661,In_969);
and U1948 (N_1948,In_119,In_1836);
nor U1949 (N_1949,In_1337,In_2349);
and U1950 (N_1950,In_2271,In_1681);
nor U1951 (N_1951,In_512,In_108);
nand U1952 (N_1952,In_720,In_438);
and U1953 (N_1953,In_2083,In_1194);
or U1954 (N_1954,In_2391,In_1861);
or U1955 (N_1955,In_1924,In_2052);
nor U1956 (N_1956,In_1561,In_21);
and U1957 (N_1957,In_2491,In_1374);
or U1958 (N_1958,In_202,In_104);
nor U1959 (N_1959,In_2289,In_43);
or U1960 (N_1960,In_1190,In_2081);
nand U1961 (N_1961,In_1608,In_344);
nand U1962 (N_1962,In_1838,In_590);
nor U1963 (N_1963,In_7,In_1743);
nor U1964 (N_1964,In_98,In_1712);
nand U1965 (N_1965,In_684,In_2427);
nor U1966 (N_1966,In_1264,In_2495);
nand U1967 (N_1967,In_149,In_1825);
nand U1968 (N_1968,In_746,In_167);
nand U1969 (N_1969,In_2128,In_1);
nor U1970 (N_1970,In_1800,In_1793);
nand U1971 (N_1971,In_602,In_1436);
nor U1972 (N_1972,In_570,In_719);
or U1973 (N_1973,In_1588,In_635);
nand U1974 (N_1974,In_759,In_2015);
and U1975 (N_1975,In_2386,In_2235);
nand U1976 (N_1976,In_1404,In_944);
nand U1977 (N_1977,In_159,In_418);
or U1978 (N_1978,In_1669,In_2442);
and U1979 (N_1979,In_1220,In_2278);
nor U1980 (N_1980,In_1630,In_908);
nor U1981 (N_1981,In_22,In_563);
or U1982 (N_1982,In_1775,In_1512);
and U1983 (N_1983,In_212,In_1255);
nor U1984 (N_1984,In_1807,In_1357);
and U1985 (N_1985,In_585,In_1223);
or U1986 (N_1986,In_897,In_1772);
nand U1987 (N_1987,In_1972,In_1265);
and U1988 (N_1988,In_2136,In_382);
and U1989 (N_1989,In_1810,In_1404);
nor U1990 (N_1990,In_2294,In_493);
or U1991 (N_1991,In_840,In_2222);
and U1992 (N_1992,In_712,In_1180);
or U1993 (N_1993,In_1793,In_2492);
nor U1994 (N_1994,In_2061,In_1395);
or U1995 (N_1995,In_1074,In_389);
and U1996 (N_1996,In_545,In_2071);
nor U1997 (N_1997,In_2254,In_1105);
nor U1998 (N_1998,In_647,In_1958);
or U1999 (N_1999,In_249,In_555);
nor U2000 (N_2000,In_2038,In_1670);
or U2001 (N_2001,In_1921,In_31);
nor U2002 (N_2002,In_93,In_1817);
and U2003 (N_2003,In_1649,In_999);
and U2004 (N_2004,In_40,In_1170);
nand U2005 (N_2005,In_1528,In_1937);
nor U2006 (N_2006,In_646,In_1388);
nand U2007 (N_2007,In_116,In_697);
nand U2008 (N_2008,In_1212,In_1122);
nand U2009 (N_2009,In_363,In_2175);
or U2010 (N_2010,In_1848,In_1780);
nand U2011 (N_2011,In_1312,In_1177);
or U2012 (N_2012,In_1424,In_562);
and U2013 (N_2013,In_442,In_211);
nor U2014 (N_2014,In_1626,In_1761);
or U2015 (N_2015,In_951,In_2283);
or U2016 (N_2016,In_953,In_2271);
or U2017 (N_2017,In_1688,In_2373);
nor U2018 (N_2018,In_1960,In_2460);
nor U2019 (N_2019,In_1903,In_444);
or U2020 (N_2020,In_982,In_455);
or U2021 (N_2021,In_2247,In_92);
or U2022 (N_2022,In_2384,In_124);
and U2023 (N_2023,In_2396,In_1480);
and U2024 (N_2024,In_423,In_394);
or U2025 (N_2025,In_1204,In_1271);
and U2026 (N_2026,In_1112,In_1706);
nor U2027 (N_2027,In_2125,In_1745);
nor U2028 (N_2028,In_974,In_1216);
and U2029 (N_2029,In_1308,In_1087);
nor U2030 (N_2030,In_486,In_1405);
and U2031 (N_2031,In_1217,In_1324);
and U2032 (N_2032,In_2124,In_1686);
nor U2033 (N_2033,In_2042,In_1941);
and U2034 (N_2034,In_1060,In_661);
and U2035 (N_2035,In_1684,In_2493);
nor U2036 (N_2036,In_1620,In_767);
nand U2037 (N_2037,In_1056,In_808);
nand U2038 (N_2038,In_377,In_2144);
and U2039 (N_2039,In_2315,In_817);
nand U2040 (N_2040,In_7,In_1003);
nor U2041 (N_2041,In_1479,In_1740);
nor U2042 (N_2042,In_1658,In_1069);
nand U2043 (N_2043,In_973,In_2211);
or U2044 (N_2044,In_1973,In_803);
nand U2045 (N_2045,In_1906,In_1903);
nor U2046 (N_2046,In_1001,In_2481);
nor U2047 (N_2047,In_925,In_781);
and U2048 (N_2048,In_733,In_96);
nor U2049 (N_2049,In_1300,In_1346);
nand U2050 (N_2050,In_1421,In_768);
or U2051 (N_2051,In_446,In_2454);
and U2052 (N_2052,In_999,In_593);
and U2053 (N_2053,In_329,In_1176);
and U2054 (N_2054,In_1685,In_1464);
nand U2055 (N_2055,In_54,In_1640);
xor U2056 (N_2056,In_332,In_1759);
or U2057 (N_2057,In_753,In_2094);
and U2058 (N_2058,In_931,In_880);
and U2059 (N_2059,In_2294,In_2199);
nor U2060 (N_2060,In_1943,In_366);
nand U2061 (N_2061,In_1084,In_1659);
nand U2062 (N_2062,In_1920,In_2205);
or U2063 (N_2063,In_1284,In_1381);
nor U2064 (N_2064,In_2181,In_1932);
nand U2065 (N_2065,In_2074,In_206);
nand U2066 (N_2066,In_1145,In_624);
nor U2067 (N_2067,In_885,In_1636);
and U2068 (N_2068,In_1088,In_572);
nor U2069 (N_2069,In_1396,In_618);
nand U2070 (N_2070,In_1016,In_707);
nand U2071 (N_2071,In_1119,In_2168);
and U2072 (N_2072,In_1399,In_1465);
nand U2073 (N_2073,In_1743,In_618);
and U2074 (N_2074,In_293,In_78);
or U2075 (N_2075,In_1529,In_888);
xor U2076 (N_2076,In_1150,In_722);
and U2077 (N_2077,In_410,In_1806);
nor U2078 (N_2078,In_1282,In_1685);
or U2079 (N_2079,In_1455,In_579);
and U2080 (N_2080,In_1615,In_1465);
and U2081 (N_2081,In_684,In_908);
or U2082 (N_2082,In_690,In_633);
and U2083 (N_2083,In_1205,In_2174);
and U2084 (N_2084,In_2137,In_772);
nor U2085 (N_2085,In_1496,In_2192);
and U2086 (N_2086,In_1941,In_1343);
nor U2087 (N_2087,In_2288,In_1296);
nor U2088 (N_2088,In_1646,In_1851);
nor U2089 (N_2089,In_200,In_970);
or U2090 (N_2090,In_98,In_779);
nand U2091 (N_2091,In_111,In_1633);
nor U2092 (N_2092,In_285,In_895);
nand U2093 (N_2093,In_1157,In_277);
nand U2094 (N_2094,In_499,In_165);
or U2095 (N_2095,In_1047,In_658);
and U2096 (N_2096,In_656,In_2294);
nand U2097 (N_2097,In_1728,In_1994);
or U2098 (N_2098,In_47,In_1820);
nand U2099 (N_2099,In_1631,In_2079);
nand U2100 (N_2100,In_844,In_1940);
and U2101 (N_2101,In_97,In_2207);
or U2102 (N_2102,In_2045,In_1519);
or U2103 (N_2103,In_708,In_1432);
nand U2104 (N_2104,In_515,In_1516);
nor U2105 (N_2105,In_1492,In_668);
or U2106 (N_2106,In_2225,In_888);
nor U2107 (N_2107,In_2267,In_2233);
and U2108 (N_2108,In_600,In_680);
or U2109 (N_2109,In_176,In_1895);
and U2110 (N_2110,In_1710,In_128);
nand U2111 (N_2111,In_1622,In_1608);
or U2112 (N_2112,In_97,In_564);
and U2113 (N_2113,In_1366,In_283);
nand U2114 (N_2114,In_934,In_2401);
nor U2115 (N_2115,In_195,In_2175);
and U2116 (N_2116,In_1399,In_994);
and U2117 (N_2117,In_663,In_1432);
and U2118 (N_2118,In_1581,In_2228);
nand U2119 (N_2119,In_181,In_1300);
or U2120 (N_2120,In_2413,In_2405);
nand U2121 (N_2121,In_1151,In_92);
and U2122 (N_2122,In_276,In_561);
and U2123 (N_2123,In_1932,In_2124);
and U2124 (N_2124,In_1786,In_790);
nand U2125 (N_2125,In_2451,In_191);
and U2126 (N_2126,In_256,In_909);
or U2127 (N_2127,In_2037,In_1529);
or U2128 (N_2128,In_645,In_2123);
and U2129 (N_2129,In_893,In_1651);
or U2130 (N_2130,In_2000,In_2421);
or U2131 (N_2131,In_1325,In_202);
and U2132 (N_2132,In_1939,In_594);
and U2133 (N_2133,In_1608,In_965);
nor U2134 (N_2134,In_851,In_1320);
nand U2135 (N_2135,In_1139,In_2266);
xor U2136 (N_2136,In_1770,In_1538);
or U2137 (N_2137,In_1253,In_1161);
nor U2138 (N_2138,In_607,In_1270);
nand U2139 (N_2139,In_963,In_2294);
and U2140 (N_2140,In_1935,In_2360);
or U2141 (N_2141,In_1128,In_284);
nor U2142 (N_2142,In_2213,In_614);
nor U2143 (N_2143,In_553,In_717);
nor U2144 (N_2144,In_1681,In_210);
nor U2145 (N_2145,In_973,In_2422);
or U2146 (N_2146,In_524,In_920);
nor U2147 (N_2147,In_1687,In_1056);
and U2148 (N_2148,In_364,In_2386);
nand U2149 (N_2149,In_690,In_2021);
nor U2150 (N_2150,In_898,In_1763);
nand U2151 (N_2151,In_1817,In_317);
nand U2152 (N_2152,In_592,In_1357);
nand U2153 (N_2153,In_2098,In_533);
nand U2154 (N_2154,In_1888,In_1758);
and U2155 (N_2155,In_572,In_1857);
and U2156 (N_2156,In_1349,In_108);
or U2157 (N_2157,In_187,In_2347);
nand U2158 (N_2158,In_856,In_293);
or U2159 (N_2159,In_1196,In_625);
nor U2160 (N_2160,In_133,In_145);
nor U2161 (N_2161,In_151,In_1226);
nand U2162 (N_2162,In_1229,In_910);
or U2163 (N_2163,In_608,In_987);
nand U2164 (N_2164,In_1357,In_413);
or U2165 (N_2165,In_1690,In_2353);
nand U2166 (N_2166,In_708,In_287);
nand U2167 (N_2167,In_1036,In_2088);
nand U2168 (N_2168,In_1895,In_1732);
and U2169 (N_2169,In_595,In_2391);
and U2170 (N_2170,In_1688,In_1974);
and U2171 (N_2171,In_1278,In_1618);
or U2172 (N_2172,In_361,In_2068);
or U2173 (N_2173,In_1187,In_1191);
nor U2174 (N_2174,In_2070,In_1335);
and U2175 (N_2175,In_2088,In_146);
or U2176 (N_2176,In_1900,In_1702);
nand U2177 (N_2177,In_2159,In_1770);
or U2178 (N_2178,In_1997,In_385);
nor U2179 (N_2179,In_2309,In_319);
nand U2180 (N_2180,In_1463,In_197);
xor U2181 (N_2181,In_1269,In_1723);
or U2182 (N_2182,In_1413,In_638);
nor U2183 (N_2183,In_2468,In_271);
nand U2184 (N_2184,In_107,In_144);
nor U2185 (N_2185,In_853,In_1503);
nand U2186 (N_2186,In_1492,In_1938);
nand U2187 (N_2187,In_1533,In_1694);
and U2188 (N_2188,In_1077,In_1880);
and U2189 (N_2189,In_450,In_1038);
or U2190 (N_2190,In_615,In_1739);
nor U2191 (N_2191,In_884,In_544);
or U2192 (N_2192,In_1635,In_1963);
nor U2193 (N_2193,In_1134,In_1039);
nand U2194 (N_2194,In_2071,In_1614);
nand U2195 (N_2195,In_731,In_1065);
and U2196 (N_2196,In_878,In_2184);
or U2197 (N_2197,In_2473,In_63);
or U2198 (N_2198,In_2340,In_592);
nand U2199 (N_2199,In_502,In_654);
nor U2200 (N_2200,In_1456,In_2235);
nand U2201 (N_2201,In_1571,In_884);
and U2202 (N_2202,In_381,In_1308);
nand U2203 (N_2203,In_1474,In_1336);
nand U2204 (N_2204,In_2020,In_366);
and U2205 (N_2205,In_441,In_2044);
and U2206 (N_2206,In_587,In_2137);
nand U2207 (N_2207,In_2314,In_478);
nand U2208 (N_2208,In_1464,In_1086);
nor U2209 (N_2209,In_1619,In_550);
nand U2210 (N_2210,In_2347,In_2133);
nand U2211 (N_2211,In_225,In_1394);
or U2212 (N_2212,In_588,In_1376);
and U2213 (N_2213,In_2373,In_1535);
and U2214 (N_2214,In_1359,In_2212);
nand U2215 (N_2215,In_671,In_2428);
xnor U2216 (N_2216,In_2339,In_2358);
or U2217 (N_2217,In_2404,In_2424);
nand U2218 (N_2218,In_1986,In_1466);
nand U2219 (N_2219,In_1060,In_276);
or U2220 (N_2220,In_880,In_1423);
nor U2221 (N_2221,In_1719,In_324);
nand U2222 (N_2222,In_2127,In_680);
nor U2223 (N_2223,In_77,In_42);
nor U2224 (N_2224,In_1592,In_1452);
nand U2225 (N_2225,In_179,In_2113);
nand U2226 (N_2226,In_2335,In_1736);
and U2227 (N_2227,In_1768,In_416);
nor U2228 (N_2228,In_1062,In_2033);
nand U2229 (N_2229,In_1187,In_1613);
and U2230 (N_2230,In_2393,In_386);
nor U2231 (N_2231,In_1235,In_1084);
or U2232 (N_2232,In_1684,In_2323);
and U2233 (N_2233,In_1367,In_1002);
nand U2234 (N_2234,In_1859,In_867);
or U2235 (N_2235,In_147,In_1073);
nand U2236 (N_2236,In_2094,In_1973);
nor U2237 (N_2237,In_1135,In_1692);
and U2238 (N_2238,In_1573,In_2202);
nand U2239 (N_2239,In_1883,In_1880);
nand U2240 (N_2240,In_1240,In_2175);
nand U2241 (N_2241,In_1861,In_1011);
nor U2242 (N_2242,In_2228,In_1617);
nor U2243 (N_2243,In_1704,In_1511);
or U2244 (N_2244,In_238,In_1189);
nand U2245 (N_2245,In_578,In_1818);
or U2246 (N_2246,In_48,In_119);
or U2247 (N_2247,In_759,In_1014);
xnor U2248 (N_2248,In_2342,In_2304);
nand U2249 (N_2249,In_2053,In_1191);
or U2250 (N_2250,In_174,In_1010);
and U2251 (N_2251,In_1821,In_2415);
and U2252 (N_2252,In_2358,In_2223);
nand U2253 (N_2253,In_262,In_1282);
nand U2254 (N_2254,In_645,In_1329);
or U2255 (N_2255,In_1071,In_877);
nor U2256 (N_2256,In_2460,In_2322);
or U2257 (N_2257,In_557,In_1694);
nand U2258 (N_2258,In_626,In_2086);
nand U2259 (N_2259,In_2415,In_2027);
nand U2260 (N_2260,In_506,In_584);
and U2261 (N_2261,In_2172,In_994);
nor U2262 (N_2262,In_1444,In_2290);
nor U2263 (N_2263,In_886,In_1065);
or U2264 (N_2264,In_928,In_255);
nor U2265 (N_2265,In_1570,In_1014);
nand U2266 (N_2266,In_2014,In_1334);
or U2267 (N_2267,In_1195,In_223);
or U2268 (N_2268,In_1036,In_2085);
nand U2269 (N_2269,In_1987,In_1027);
or U2270 (N_2270,In_1374,In_2413);
nand U2271 (N_2271,In_1992,In_656);
and U2272 (N_2272,In_1855,In_821);
or U2273 (N_2273,In_582,In_2100);
nor U2274 (N_2274,In_724,In_689);
nand U2275 (N_2275,In_1460,In_2002);
or U2276 (N_2276,In_948,In_206);
xnor U2277 (N_2277,In_849,In_1950);
nand U2278 (N_2278,In_2042,In_335);
nand U2279 (N_2279,In_2372,In_150);
or U2280 (N_2280,In_568,In_67);
nor U2281 (N_2281,In_1065,In_48);
nor U2282 (N_2282,In_949,In_290);
and U2283 (N_2283,In_950,In_1691);
nor U2284 (N_2284,In_1244,In_248);
nand U2285 (N_2285,In_172,In_2133);
and U2286 (N_2286,In_2464,In_1976);
nand U2287 (N_2287,In_518,In_2320);
nor U2288 (N_2288,In_269,In_1459);
or U2289 (N_2289,In_22,In_1677);
and U2290 (N_2290,In_1222,In_595);
nor U2291 (N_2291,In_1060,In_1229);
and U2292 (N_2292,In_2491,In_1704);
nand U2293 (N_2293,In_2381,In_1025);
nand U2294 (N_2294,In_698,In_666);
and U2295 (N_2295,In_2075,In_1200);
or U2296 (N_2296,In_194,In_1232);
and U2297 (N_2297,In_734,In_2280);
nand U2298 (N_2298,In_1003,In_494);
or U2299 (N_2299,In_219,In_1382);
or U2300 (N_2300,In_1652,In_530);
or U2301 (N_2301,In_1009,In_1650);
xnor U2302 (N_2302,In_1949,In_381);
and U2303 (N_2303,In_1233,In_1566);
and U2304 (N_2304,In_1298,In_1536);
and U2305 (N_2305,In_1970,In_1758);
and U2306 (N_2306,In_1122,In_1544);
and U2307 (N_2307,In_1006,In_1850);
nor U2308 (N_2308,In_2006,In_1178);
and U2309 (N_2309,In_449,In_804);
and U2310 (N_2310,In_691,In_313);
nor U2311 (N_2311,In_1452,In_200);
and U2312 (N_2312,In_1989,In_353);
nor U2313 (N_2313,In_289,In_1324);
or U2314 (N_2314,In_1045,In_228);
or U2315 (N_2315,In_591,In_2142);
and U2316 (N_2316,In_831,In_1593);
and U2317 (N_2317,In_192,In_1517);
nand U2318 (N_2318,In_968,In_1766);
nor U2319 (N_2319,In_2015,In_2202);
and U2320 (N_2320,In_50,In_1459);
nor U2321 (N_2321,In_644,In_1160);
nand U2322 (N_2322,In_1551,In_1303);
and U2323 (N_2323,In_2096,In_503);
or U2324 (N_2324,In_603,In_1780);
and U2325 (N_2325,In_2223,In_1744);
or U2326 (N_2326,In_988,In_2407);
nor U2327 (N_2327,In_1954,In_894);
or U2328 (N_2328,In_1171,In_2199);
and U2329 (N_2329,In_566,In_672);
nor U2330 (N_2330,In_2420,In_1566);
or U2331 (N_2331,In_1520,In_1865);
nor U2332 (N_2332,In_1925,In_1467);
or U2333 (N_2333,In_1938,In_221);
and U2334 (N_2334,In_2336,In_519);
or U2335 (N_2335,In_1349,In_1466);
or U2336 (N_2336,In_1507,In_133);
and U2337 (N_2337,In_455,In_211);
nand U2338 (N_2338,In_1393,In_1159);
nand U2339 (N_2339,In_109,In_1920);
or U2340 (N_2340,In_1256,In_2030);
and U2341 (N_2341,In_607,In_252);
nand U2342 (N_2342,In_29,In_1027);
nor U2343 (N_2343,In_628,In_2120);
and U2344 (N_2344,In_2417,In_2313);
and U2345 (N_2345,In_1041,In_669);
nor U2346 (N_2346,In_1079,In_2160);
nand U2347 (N_2347,In_1789,In_1847);
nor U2348 (N_2348,In_1582,In_1591);
nand U2349 (N_2349,In_1866,In_1887);
nor U2350 (N_2350,In_2058,In_1305);
nor U2351 (N_2351,In_2035,In_1080);
nand U2352 (N_2352,In_2071,In_29);
and U2353 (N_2353,In_13,In_1241);
nor U2354 (N_2354,In_2027,In_96);
and U2355 (N_2355,In_1704,In_1449);
or U2356 (N_2356,In_526,In_1146);
or U2357 (N_2357,In_1224,In_430);
nor U2358 (N_2358,In_1682,In_1865);
and U2359 (N_2359,In_1306,In_1534);
nand U2360 (N_2360,In_2451,In_1464);
and U2361 (N_2361,In_1803,In_1625);
and U2362 (N_2362,In_157,In_2188);
and U2363 (N_2363,In_2026,In_121);
nor U2364 (N_2364,In_1612,In_1180);
or U2365 (N_2365,In_185,In_380);
nand U2366 (N_2366,In_201,In_1985);
or U2367 (N_2367,In_2076,In_2450);
nor U2368 (N_2368,In_2096,In_108);
nand U2369 (N_2369,In_2488,In_493);
and U2370 (N_2370,In_1463,In_619);
nor U2371 (N_2371,In_2282,In_1824);
nand U2372 (N_2372,In_1605,In_1964);
nand U2373 (N_2373,In_645,In_2474);
nor U2374 (N_2374,In_841,In_719);
and U2375 (N_2375,In_2433,In_501);
and U2376 (N_2376,In_1885,In_323);
nand U2377 (N_2377,In_1093,In_308);
nand U2378 (N_2378,In_842,In_1930);
nor U2379 (N_2379,In_1278,In_2261);
nor U2380 (N_2380,In_1204,In_1035);
and U2381 (N_2381,In_1566,In_87);
or U2382 (N_2382,In_1088,In_2162);
and U2383 (N_2383,In_1746,In_2346);
or U2384 (N_2384,In_1457,In_1094);
nor U2385 (N_2385,In_1920,In_1355);
nand U2386 (N_2386,In_2366,In_623);
xor U2387 (N_2387,In_1367,In_1864);
or U2388 (N_2388,In_484,In_332);
nor U2389 (N_2389,In_929,In_844);
and U2390 (N_2390,In_1734,In_292);
and U2391 (N_2391,In_327,In_1094);
nor U2392 (N_2392,In_140,In_585);
and U2393 (N_2393,In_1163,In_1999);
or U2394 (N_2394,In_936,In_860);
or U2395 (N_2395,In_1725,In_587);
nor U2396 (N_2396,In_382,In_1098);
nand U2397 (N_2397,In_2147,In_123);
nor U2398 (N_2398,In_1344,In_75);
nand U2399 (N_2399,In_2471,In_1830);
and U2400 (N_2400,In_1573,In_675);
or U2401 (N_2401,In_1592,In_1383);
nand U2402 (N_2402,In_345,In_171);
nand U2403 (N_2403,In_1411,In_1727);
or U2404 (N_2404,In_143,In_1667);
nor U2405 (N_2405,In_1111,In_687);
and U2406 (N_2406,In_1344,In_783);
nor U2407 (N_2407,In_188,In_786);
or U2408 (N_2408,In_1618,In_1059);
nor U2409 (N_2409,In_2191,In_278);
and U2410 (N_2410,In_925,In_2147);
or U2411 (N_2411,In_2124,In_1726);
nor U2412 (N_2412,In_1125,In_1464);
nor U2413 (N_2413,In_1019,In_1119);
or U2414 (N_2414,In_641,In_1895);
nor U2415 (N_2415,In_176,In_1573);
nor U2416 (N_2416,In_524,In_1901);
or U2417 (N_2417,In_1935,In_785);
nand U2418 (N_2418,In_2230,In_2262);
and U2419 (N_2419,In_1985,In_2230);
and U2420 (N_2420,In_1227,In_258);
nor U2421 (N_2421,In_2270,In_1072);
nand U2422 (N_2422,In_1994,In_1694);
and U2423 (N_2423,In_2106,In_1328);
or U2424 (N_2424,In_1291,In_1673);
and U2425 (N_2425,In_1318,In_2002);
nand U2426 (N_2426,In_1076,In_1449);
or U2427 (N_2427,In_431,In_1402);
and U2428 (N_2428,In_454,In_86);
nor U2429 (N_2429,In_2490,In_1501);
nand U2430 (N_2430,In_1641,In_2337);
and U2431 (N_2431,In_804,In_1416);
and U2432 (N_2432,In_387,In_2299);
or U2433 (N_2433,In_224,In_2235);
or U2434 (N_2434,In_1734,In_2080);
nor U2435 (N_2435,In_1368,In_1468);
and U2436 (N_2436,In_158,In_1484);
or U2437 (N_2437,In_361,In_1799);
or U2438 (N_2438,In_1210,In_97);
nor U2439 (N_2439,In_1,In_1296);
and U2440 (N_2440,In_1611,In_1389);
and U2441 (N_2441,In_2377,In_969);
nor U2442 (N_2442,In_2006,In_1243);
nand U2443 (N_2443,In_278,In_860);
or U2444 (N_2444,In_1129,In_855);
nand U2445 (N_2445,In_805,In_1647);
and U2446 (N_2446,In_507,In_639);
or U2447 (N_2447,In_422,In_1712);
or U2448 (N_2448,In_982,In_1129);
nor U2449 (N_2449,In_532,In_1141);
and U2450 (N_2450,In_1894,In_956);
or U2451 (N_2451,In_388,In_957);
or U2452 (N_2452,In_1104,In_891);
nand U2453 (N_2453,In_1814,In_2499);
and U2454 (N_2454,In_759,In_575);
or U2455 (N_2455,In_2011,In_948);
or U2456 (N_2456,In_73,In_1065);
and U2457 (N_2457,In_1030,In_2112);
nand U2458 (N_2458,In_932,In_154);
nand U2459 (N_2459,In_1352,In_1614);
nand U2460 (N_2460,In_772,In_28);
nand U2461 (N_2461,In_374,In_193);
and U2462 (N_2462,In_2089,In_1821);
and U2463 (N_2463,In_1526,In_1429);
and U2464 (N_2464,In_1867,In_190);
nand U2465 (N_2465,In_2390,In_2394);
nor U2466 (N_2466,In_839,In_2166);
or U2467 (N_2467,In_634,In_2347);
and U2468 (N_2468,In_609,In_2085);
and U2469 (N_2469,In_171,In_166);
nor U2470 (N_2470,In_1306,In_852);
and U2471 (N_2471,In_63,In_1646);
nor U2472 (N_2472,In_1563,In_1206);
nand U2473 (N_2473,In_181,In_2250);
and U2474 (N_2474,In_2317,In_2293);
and U2475 (N_2475,In_2269,In_1887);
nand U2476 (N_2476,In_254,In_393);
and U2477 (N_2477,In_2456,In_394);
or U2478 (N_2478,In_2056,In_1607);
or U2479 (N_2479,In_37,In_591);
and U2480 (N_2480,In_803,In_423);
or U2481 (N_2481,In_782,In_249);
nor U2482 (N_2482,In_1649,In_1498);
or U2483 (N_2483,In_1738,In_975);
or U2484 (N_2484,In_196,In_1802);
nor U2485 (N_2485,In_321,In_1407);
nand U2486 (N_2486,In_1975,In_541);
or U2487 (N_2487,In_2490,In_67);
and U2488 (N_2488,In_2039,In_538);
nand U2489 (N_2489,In_1560,In_1368);
nand U2490 (N_2490,In_916,In_1609);
or U2491 (N_2491,In_712,In_1276);
nand U2492 (N_2492,In_734,In_906);
or U2493 (N_2493,In_932,In_2423);
and U2494 (N_2494,In_2479,In_2193);
nand U2495 (N_2495,In_1518,In_1513);
nor U2496 (N_2496,In_2335,In_94);
nor U2497 (N_2497,In_172,In_2143);
nor U2498 (N_2498,In_1287,In_1115);
nor U2499 (N_2499,In_1754,In_1780);
nor U2500 (N_2500,In_1914,In_434);
and U2501 (N_2501,In_879,In_1006);
nand U2502 (N_2502,In_66,In_298);
nor U2503 (N_2503,In_1247,In_2136);
nor U2504 (N_2504,In_912,In_1029);
nand U2505 (N_2505,In_1300,In_1988);
or U2506 (N_2506,In_1997,In_799);
and U2507 (N_2507,In_1987,In_2156);
or U2508 (N_2508,In_2361,In_1657);
and U2509 (N_2509,In_2153,In_597);
and U2510 (N_2510,In_2349,In_2228);
and U2511 (N_2511,In_459,In_1672);
or U2512 (N_2512,In_2474,In_1505);
and U2513 (N_2513,In_1130,In_1103);
or U2514 (N_2514,In_1549,In_1683);
nor U2515 (N_2515,In_849,In_625);
and U2516 (N_2516,In_705,In_1777);
nand U2517 (N_2517,In_1391,In_620);
and U2518 (N_2518,In_745,In_2411);
or U2519 (N_2519,In_2378,In_907);
nand U2520 (N_2520,In_1994,In_1792);
nor U2521 (N_2521,In_1112,In_1905);
nand U2522 (N_2522,In_997,In_854);
nor U2523 (N_2523,In_1663,In_16);
and U2524 (N_2524,In_773,In_521);
and U2525 (N_2525,In_2285,In_1470);
nor U2526 (N_2526,In_1161,In_1180);
nor U2527 (N_2527,In_2321,In_2042);
nand U2528 (N_2528,In_348,In_969);
or U2529 (N_2529,In_1787,In_2433);
and U2530 (N_2530,In_1013,In_1929);
nand U2531 (N_2531,In_1608,In_1620);
or U2532 (N_2532,In_1115,In_333);
xor U2533 (N_2533,In_153,In_2288);
or U2534 (N_2534,In_2114,In_1332);
and U2535 (N_2535,In_15,In_1782);
or U2536 (N_2536,In_2395,In_342);
or U2537 (N_2537,In_79,In_1741);
nand U2538 (N_2538,In_151,In_305);
nand U2539 (N_2539,In_1217,In_1861);
and U2540 (N_2540,In_175,In_2318);
nor U2541 (N_2541,In_882,In_542);
or U2542 (N_2542,In_1765,In_1292);
nor U2543 (N_2543,In_555,In_1509);
and U2544 (N_2544,In_1732,In_160);
or U2545 (N_2545,In_1667,In_388);
and U2546 (N_2546,In_1408,In_522);
nand U2547 (N_2547,In_18,In_1229);
nor U2548 (N_2548,In_957,In_1580);
and U2549 (N_2549,In_874,In_1492);
and U2550 (N_2550,In_1302,In_1255);
and U2551 (N_2551,In_2189,In_1794);
nor U2552 (N_2552,In_1345,In_2001);
and U2553 (N_2553,In_234,In_1299);
or U2554 (N_2554,In_1450,In_387);
nand U2555 (N_2555,In_2424,In_1841);
or U2556 (N_2556,In_1477,In_2461);
and U2557 (N_2557,In_1216,In_622);
nor U2558 (N_2558,In_1835,In_2191);
or U2559 (N_2559,In_826,In_775);
nand U2560 (N_2560,In_1967,In_1612);
nor U2561 (N_2561,In_624,In_2015);
or U2562 (N_2562,In_364,In_2178);
and U2563 (N_2563,In_2319,In_944);
or U2564 (N_2564,In_1723,In_2085);
or U2565 (N_2565,In_1114,In_812);
or U2566 (N_2566,In_587,In_559);
nor U2567 (N_2567,In_2076,In_865);
and U2568 (N_2568,In_628,In_1675);
or U2569 (N_2569,In_638,In_2120);
or U2570 (N_2570,In_596,In_619);
nand U2571 (N_2571,In_1151,In_259);
and U2572 (N_2572,In_1493,In_1699);
or U2573 (N_2573,In_1974,In_1734);
nor U2574 (N_2574,In_1482,In_1557);
nand U2575 (N_2575,In_1973,In_768);
and U2576 (N_2576,In_1321,In_1475);
nand U2577 (N_2577,In_2146,In_2339);
nor U2578 (N_2578,In_1766,In_1939);
nand U2579 (N_2579,In_242,In_1261);
or U2580 (N_2580,In_2294,In_734);
nor U2581 (N_2581,In_1654,In_1134);
and U2582 (N_2582,In_124,In_520);
and U2583 (N_2583,In_444,In_2333);
and U2584 (N_2584,In_1394,In_1620);
and U2585 (N_2585,In_1108,In_913);
nand U2586 (N_2586,In_41,In_1837);
nand U2587 (N_2587,In_2033,In_1760);
nor U2588 (N_2588,In_1266,In_1056);
nor U2589 (N_2589,In_1669,In_1119);
and U2590 (N_2590,In_461,In_119);
and U2591 (N_2591,In_310,In_2477);
nand U2592 (N_2592,In_1459,In_753);
nand U2593 (N_2593,In_1005,In_302);
or U2594 (N_2594,In_1460,In_964);
or U2595 (N_2595,In_1484,In_1745);
and U2596 (N_2596,In_1543,In_837);
nor U2597 (N_2597,In_1302,In_379);
nand U2598 (N_2598,In_357,In_657);
and U2599 (N_2599,In_2450,In_2018);
or U2600 (N_2600,In_1091,In_2282);
and U2601 (N_2601,In_1454,In_1311);
nand U2602 (N_2602,In_1035,In_1008);
and U2603 (N_2603,In_688,In_1002);
or U2604 (N_2604,In_743,In_1419);
nand U2605 (N_2605,In_2077,In_1479);
nand U2606 (N_2606,In_904,In_932);
and U2607 (N_2607,In_1585,In_722);
or U2608 (N_2608,In_2105,In_16);
nor U2609 (N_2609,In_879,In_1899);
nand U2610 (N_2610,In_1460,In_960);
nand U2611 (N_2611,In_1949,In_1768);
or U2612 (N_2612,In_1997,In_624);
and U2613 (N_2613,In_1156,In_1827);
nor U2614 (N_2614,In_923,In_2486);
and U2615 (N_2615,In_169,In_2160);
nand U2616 (N_2616,In_2364,In_1603);
nor U2617 (N_2617,In_1049,In_1999);
xnor U2618 (N_2618,In_347,In_263);
and U2619 (N_2619,In_2391,In_659);
and U2620 (N_2620,In_1425,In_1725);
nor U2621 (N_2621,In_304,In_370);
or U2622 (N_2622,In_943,In_2158);
or U2623 (N_2623,In_165,In_827);
nor U2624 (N_2624,In_1514,In_1202);
or U2625 (N_2625,In_2342,In_896);
or U2626 (N_2626,In_2025,In_1553);
or U2627 (N_2627,In_118,In_691);
nor U2628 (N_2628,In_493,In_579);
and U2629 (N_2629,In_1222,In_320);
and U2630 (N_2630,In_2086,In_320);
and U2631 (N_2631,In_2452,In_981);
nand U2632 (N_2632,In_1762,In_1185);
nor U2633 (N_2633,In_256,In_80);
nand U2634 (N_2634,In_457,In_843);
and U2635 (N_2635,In_214,In_1181);
nor U2636 (N_2636,In_556,In_1049);
nor U2637 (N_2637,In_1195,In_1488);
and U2638 (N_2638,In_1342,In_2134);
or U2639 (N_2639,In_2452,In_1109);
nor U2640 (N_2640,In_1752,In_2473);
nand U2641 (N_2641,In_1605,In_609);
and U2642 (N_2642,In_2333,In_897);
and U2643 (N_2643,In_1384,In_707);
nand U2644 (N_2644,In_2178,In_291);
nand U2645 (N_2645,In_1623,In_1418);
nor U2646 (N_2646,In_161,In_1079);
nand U2647 (N_2647,In_2279,In_1228);
nor U2648 (N_2648,In_510,In_610);
nor U2649 (N_2649,In_1907,In_1819);
and U2650 (N_2650,In_404,In_991);
nor U2651 (N_2651,In_887,In_1023);
and U2652 (N_2652,In_2318,In_2060);
or U2653 (N_2653,In_2032,In_399);
and U2654 (N_2654,In_1461,In_1844);
and U2655 (N_2655,In_542,In_1958);
nor U2656 (N_2656,In_1522,In_2409);
nor U2657 (N_2657,In_822,In_2285);
or U2658 (N_2658,In_172,In_1749);
nand U2659 (N_2659,In_1609,In_2284);
and U2660 (N_2660,In_1964,In_610);
and U2661 (N_2661,In_1685,In_593);
or U2662 (N_2662,In_2048,In_1776);
or U2663 (N_2663,In_1330,In_1282);
nand U2664 (N_2664,In_1282,In_60);
nand U2665 (N_2665,In_2041,In_215);
or U2666 (N_2666,In_2099,In_724);
and U2667 (N_2667,In_438,In_1988);
or U2668 (N_2668,In_1618,In_1404);
and U2669 (N_2669,In_290,In_1222);
nand U2670 (N_2670,In_737,In_1653);
or U2671 (N_2671,In_226,In_2194);
and U2672 (N_2672,In_1563,In_2286);
nor U2673 (N_2673,In_984,In_1989);
nand U2674 (N_2674,In_1834,In_990);
or U2675 (N_2675,In_474,In_2223);
nand U2676 (N_2676,In_1929,In_1351);
nor U2677 (N_2677,In_610,In_829);
nand U2678 (N_2678,In_22,In_1135);
and U2679 (N_2679,In_1772,In_1327);
nor U2680 (N_2680,In_2317,In_814);
and U2681 (N_2681,In_1488,In_2243);
and U2682 (N_2682,In_2450,In_817);
or U2683 (N_2683,In_2408,In_1271);
nand U2684 (N_2684,In_670,In_848);
and U2685 (N_2685,In_1423,In_256);
nand U2686 (N_2686,In_775,In_323);
nand U2687 (N_2687,In_2108,In_399);
or U2688 (N_2688,In_2054,In_792);
or U2689 (N_2689,In_1526,In_2132);
nand U2690 (N_2690,In_1065,In_1407);
or U2691 (N_2691,In_1033,In_2475);
nor U2692 (N_2692,In_826,In_1596);
nand U2693 (N_2693,In_1148,In_1335);
and U2694 (N_2694,In_2231,In_1265);
nor U2695 (N_2695,In_2481,In_217);
nand U2696 (N_2696,In_1563,In_2324);
nor U2697 (N_2697,In_1515,In_1033);
and U2698 (N_2698,In_945,In_2221);
or U2699 (N_2699,In_718,In_2360);
or U2700 (N_2700,In_1706,In_1522);
nand U2701 (N_2701,In_517,In_234);
or U2702 (N_2702,In_449,In_680);
nand U2703 (N_2703,In_2382,In_2328);
or U2704 (N_2704,In_1487,In_75);
nor U2705 (N_2705,In_144,In_89);
nand U2706 (N_2706,In_2373,In_2198);
nor U2707 (N_2707,In_1222,In_457);
nand U2708 (N_2708,In_896,In_649);
nor U2709 (N_2709,In_1701,In_2395);
nand U2710 (N_2710,In_1717,In_322);
and U2711 (N_2711,In_2310,In_187);
or U2712 (N_2712,In_444,In_2012);
nor U2713 (N_2713,In_1305,In_1947);
and U2714 (N_2714,In_1557,In_331);
and U2715 (N_2715,In_596,In_1832);
nand U2716 (N_2716,In_199,In_27);
or U2717 (N_2717,In_1928,In_2313);
or U2718 (N_2718,In_2350,In_2335);
nand U2719 (N_2719,In_103,In_1742);
or U2720 (N_2720,In_215,In_951);
or U2721 (N_2721,In_473,In_448);
nand U2722 (N_2722,In_2242,In_199);
nand U2723 (N_2723,In_2121,In_256);
or U2724 (N_2724,In_1050,In_1412);
or U2725 (N_2725,In_1480,In_1334);
or U2726 (N_2726,In_1393,In_866);
nor U2727 (N_2727,In_2106,In_110);
or U2728 (N_2728,In_985,In_56);
xor U2729 (N_2729,In_1172,In_1684);
nand U2730 (N_2730,In_968,In_902);
nand U2731 (N_2731,In_2292,In_2329);
and U2732 (N_2732,In_2038,In_2008);
and U2733 (N_2733,In_1223,In_2165);
or U2734 (N_2734,In_2279,In_1387);
nand U2735 (N_2735,In_479,In_963);
nor U2736 (N_2736,In_1061,In_1345);
nor U2737 (N_2737,In_1195,In_2069);
and U2738 (N_2738,In_1034,In_1904);
or U2739 (N_2739,In_1816,In_1742);
nand U2740 (N_2740,In_680,In_576);
and U2741 (N_2741,In_184,In_1306);
nor U2742 (N_2742,In_2066,In_2335);
nor U2743 (N_2743,In_969,In_760);
nand U2744 (N_2744,In_1581,In_626);
and U2745 (N_2745,In_1870,In_1097);
or U2746 (N_2746,In_743,In_436);
and U2747 (N_2747,In_978,In_1826);
nor U2748 (N_2748,In_320,In_2327);
nor U2749 (N_2749,In_2382,In_112);
nor U2750 (N_2750,In_2241,In_1794);
and U2751 (N_2751,In_858,In_802);
nand U2752 (N_2752,In_1187,In_1669);
or U2753 (N_2753,In_311,In_2251);
nor U2754 (N_2754,In_879,In_1396);
nand U2755 (N_2755,In_1413,In_1953);
and U2756 (N_2756,In_893,In_2455);
nor U2757 (N_2757,In_157,In_1992);
nand U2758 (N_2758,In_662,In_180);
and U2759 (N_2759,In_1383,In_621);
nand U2760 (N_2760,In_1531,In_1216);
or U2761 (N_2761,In_1454,In_955);
or U2762 (N_2762,In_140,In_882);
and U2763 (N_2763,In_2090,In_2005);
and U2764 (N_2764,In_39,In_1829);
and U2765 (N_2765,In_1525,In_593);
nand U2766 (N_2766,In_1849,In_377);
and U2767 (N_2767,In_2291,In_1422);
or U2768 (N_2768,In_189,In_1634);
nand U2769 (N_2769,In_2303,In_1015);
or U2770 (N_2770,In_506,In_2430);
and U2771 (N_2771,In_1248,In_1621);
or U2772 (N_2772,In_1513,In_651);
nor U2773 (N_2773,In_1491,In_2091);
or U2774 (N_2774,In_1670,In_1781);
and U2775 (N_2775,In_2095,In_1686);
or U2776 (N_2776,In_148,In_2156);
and U2777 (N_2777,In_1062,In_550);
nand U2778 (N_2778,In_2294,In_1011);
and U2779 (N_2779,In_2461,In_545);
nor U2780 (N_2780,In_812,In_1616);
nand U2781 (N_2781,In_2083,In_1142);
and U2782 (N_2782,In_2425,In_864);
nand U2783 (N_2783,In_2150,In_1857);
and U2784 (N_2784,In_1824,In_28);
or U2785 (N_2785,In_208,In_924);
nor U2786 (N_2786,In_25,In_1100);
nor U2787 (N_2787,In_800,In_1130);
and U2788 (N_2788,In_584,In_14);
or U2789 (N_2789,In_1716,In_2073);
nand U2790 (N_2790,In_538,In_1858);
or U2791 (N_2791,In_1069,In_1748);
and U2792 (N_2792,In_2264,In_586);
nand U2793 (N_2793,In_549,In_772);
nand U2794 (N_2794,In_126,In_2228);
or U2795 (N_2795,In_1660,In_2317);
nand U2796 (N_2796,In_1144,In_2091);
or U2797 (N_2797,In_1302,In_1048);
nand U2798 (N_2798,In_2488,In_2184);
or U2799 (N_2799,In_61,In_1094);
nor U2800 (N_2800,In_248,In_17);
or U2801 (N_2801,In_2118,In_872);
nor U2802 (N_2802,In_2346,In_585);
nor U2803 (N_2803,In_913,In_1645);
or U2804 (N_2804,In_33,In_176);
nand U2805 (N_2805,In_197,In_1080);
and U2806 (N_2806,In_1594,In_364);
nor U2807 (N_2807,In_2029,In_809);
or U2808 (N_2808,In_413,In_44);
nor U2809 (N_2809,In_1500,In_1402);
and U2810 (N_2810,In_1464,In_1300);
and U2811 (N_2811,In_2085,In_291);
and U2812 (N_2812,In_489,In_2237);
nand U2813 (N_2813,In_473,In_466);
or U2814 (N_2814,In_2294,In_2174);
and U2815 (N_2815,In_494,In_1819);
nor U2816 (N_2816,In_1560,In_799);
or U2817 (N_2817,In_214,In_175);
and U2818 (N_2818,In_879,In_890);
nor U2819 (N_2819,In_1588,In_345);
and U2820 (N_2820,In_223,In_1421);
and U2821 (N_2821,In_1523,In_2029);
nand U2822 (N_2822,In_1774,In_2162);
or U2823 (N_2823,In_1145,In_2356);
or U2824 (N_2824,In_2082,In_1510);
and U2825 (N_2825,In_1779,In_2187);
nor U2826 (N_2826,In_1688,In_461);
nand U2827 (N_2827,In_1798,In_1027);
and U2828 (N_2828,In_114,In_190);
nand U2829 (N_2829,In_449,In_462);
nand U2830 (N_2830,In_2130,In_645);
or U2831 (N_2831,In_503,In_66);
or U2832 (N_2832,In_2028,In_1522);
nor U2833 (N_2833,In_1646,In_1375);
and U2834 (N_2834,In_1655,In_22);
nor U2835 (N_2835,In_928,In_1105);
nand U2836 (N_2836,In_1209,In_1846);
nand U2837 (N_2837,In_1107,In_1740);
nor U2838 (N_2838,In_841,In_2300);
and U2839 (N_2839,In_2467,In_1495);
xnor U2840 (N_2840,In_1519,In_1631);
nand U2841 (N_2841,In_1249,In_392);
or U2842 (N_2842,In_1518,In_394);
nor U2843 (N_2843,In_1764,In_1570);
and U2844 (N_2844,In_1007,In_2127);
nor U2845 (N_2845,In_1278,In_2326);
nand U2846 (N_2846,In_1869,In_1694);
nor U2847 (N_2847,In_1800,In_218);
nand U2848 (N_2848,In_2060,In_1404);
or U2849 (N_2849,In_161,In_1591);
and U2850 (N_2850,In_2288,In_80);
or U2851 (N_2851,In_392,In_534);
or U2852 (N_2852,In_1383,In_529);
or U2853 (N_2853,In_2474,In_1032);
nor U2854 (N_2854,In_1810,In_876);
nand U2855 (N_2855,In_88,In_351);
or U2856 (N_2856,In_878,In_1707);
nor U2857 (N_2857,In_339,In_1546);
and U2858 (N_2858,In_2317,In_2102);
or U2859 (N_2859,In_810,In_494);
and U2860 (N_2860,In_1261,In_1716);
nand U2861 (N_2861,In_960,In_186);
and U2862 (N_2862,In_428,In_1893);
nor U2863 (N_2863,In_578,In_1656);
nand U2864 (N_2864,In_1083,In_694);
or U2865 (N_2865,In_689,In_2000);
or U2866 (N_2866,In_1792,In_1460);
and U2867 (N_2867,In_1873,In_1835);
nor U2868 (N_2868,In_905,In_962);
and U2869 (N_2869,In_1982,In_1788);
or U2870 (N_2870,In_1176,In_1168);
nor U2871 (N_2871,In_1701,In_374);
and U2872 (N_2872,In_1511,In_2260);
nor U2873 (N_2873,In_816,In_1489);
or U2874 (N_2874,In_2022,In_2315);
and U2875 (N_2875,In_670,In_442);
nor U2876 (N_2876,In_1416,In_430);
or U2877 (N_2877,In_931,In_1814);
nor U2878 (N_2878,In_1297,In_237);
or U2879 (N_2879,In_2268,In_1903);
nor U2880 (N_2880,In_447,In_1091);
and U2881 (N_2881,In_449,In_1345);
or U2882 (N_2882,In_2373,In_2236);
and U2883 (N_2883,In_2285,In_1582);
nor U2884 (N_2884,In_2273,In_623);
xnor U2885 (N_2885,In_639,In_199);
and U2886 (N_2886,In_2254,In_2412);
and U2887 (N_2887,In_1851,In_350);
nand U2888 (N_2888,In_903,In_1476);
nor U2889 (N_2889,In_633,In_1058);
and U2890 (N_2890,In_285,In_115);
xor U2891 (N_2891,In_1076,In_942);
nand U2892 (N_2892,In_2391,In_822);
and U2893 (N_2893,In_53,In_1283);
or U2894 (N_2894,In_1238,In_1362);
and U2895 (N_2895,In_812,In_484);
nand U2896 (N_2896,In_2390,In_752);
nor U2897 (N_2897,In_2238,In_519);
nand U2898 (N_2898,In_498,In_1554);
nand U2899 (N_2899,In_2012,In_368);
nor U2900 (N_2900,In_1186,In_2452);
nor U2901 (N_2901,In_2327,In_641);
nor U2902 (N_2902,In_1161,In_1668);
nand U2903 (N_2903,In_2179,In_929);
and U2904 (N_2904,In_1710,In_1543);
nand U2905 (N_2905,In_2093,In_1974);
and U2906 (N_2906,In_1929,In_882);
and U2907 (N_2907,In_779,In_454);
and U2908 (N_2908,In_608,In_239);
nand U2909 (N_2909,In_2150,In_1470);
nor U2910 (N_2910,In_105,In_1915);
or U2911 (N_2911,In_1186,In_809);
nor U2912 (N_2912,In_1093,In_1799);
nand U2913 (N_2913,In_1419,In_1609);
and U2914 (N_2914,In_2216,In_1978);
nand U2915 (N_2915,In_1582,In_725);
nand U2916 (N_2916,In_840,In_810);
and U2917 (N_2917,In_2075,In_867);
nor U2918 (N_2918,In_1606,In_1546);
or U2919 (N_2919,In_1954,In_796);
nor U2920 (N_2920,In_1927,In_2006);
nand U2921 (N_2921,In_489,In_1646);
and U2922 (N_2922,In_1468,In_240);
or U2923 (N_2923,In_1636,In_516);
nor U2924 (N_2924,In_109,In_686);
nand U2925 (N_2925,In_1253,In_820);
nand U2926 (N_2926,In_407,In_1158);
and U2927 (N_2927,In_1641,In_830);
or U2928 (N_2928,In_370,In_755);
nor U2929 (N_2929,In_194,In_2087);
and U2930 (N_2930,In_2224,In_1416);
and U2931 (N_2931,In_126,In_380);
nand U2932 (N_2932,In_2394,In_541);
or U2933 (N_2933,In_876,In_517);
nor U2934 (N_2934,In_697,In_199);
nand U2935 (N_2935,In_2143,In_972);
and U2936 (N_2936,In_580,In_1490);
xnor U2937 (N_2937,In_1364,In_741);
nand U2938 (N_2938,In_1018,In_980);
or U2939 (N_2939,In_154,In_645);
and U2940 (N_2940,In_576,In_1759);
or U2941 (N_2941,In_258,In_1089);
nor U2942 (N_2942,In_47,In_239);
nand U2943 (N_2943,In_1749,In_482);
and U2944 (N_2944,In_1465,In_1020);
nor U2945 (N_2945,In_115,In_1327);
and U2946 (N_2946,In_1846,In_1245);
nand U2947 (N_2947,In_1271,In_2430);
and U2948 (N_2948,In_748,In_320);
or U2949 (N_2949,In_924,In_1202);
or U2950 (N_2950,In_909,In_435);
nor U2951 (N_2951,In_1855,In_243);
nor U2952 (N_2952,In_155,In_2033);
nor U2953 (N_2953,In_1562,In_953);
or U2954 (N_2954,In_200,In_764);
nand U2955 (N_2955,In_1015,In_1182);
nor U2956 (N_2956,In_1609,In_2160);
nor U2957 (N_2957,In_731,In_1615);
and U2958 (N_2958,In_1426,In_1863);
or U2959 (N_2959,In_904,In_648);
nor U2960 (N_2960,In_474,In_1637);
nand U2961 (N_2961,In_302,In_1368);
nor U2962 (N_2962,In_2188,In_2046);
nand U2963 (N_2963,In_2155,In_1640);
or U2964 (N_2964,In_410,In_2223);
and U2965 (N_2965,In_1481,In_424);
or U2966 (N_2966,In_151,In_1646);
nor U2967 (N_2967,In_2417,In_359);
and U2968 (N_2968,In_2132,In_2340);
nor U2969 (N_2969,In_274,In_2145);
and U2970 (N_2970,In_62,In_286);
or U2971 (N_2971,In_779,In_989);
or U2972 (N_2972,In_1575,In_1898);
and U2973 (N_2973,In_1414,In_1967);
or U2974 (N_2974,In_1991,In_737);
nand U2975 (N_2975,In_761,In_2321);
and U2976 (N_2976,In_1928,In_2412);
nand U2977 (N_2977,In_928,In_1083);
nor U2978 (N_2978,In_167,In_2242);
nand U2979 (N_2979,In_1967,In_2175);
and U2980 (N_2980,In_1853,In_1067);
or U2981 (N_2981,In_601,In_1014);
nor U2982 (N_2982,In_1199,In_272);
and U2983 (N_2983,In_174,In_989);
and U2984 (N_2984,In_1268,In_1907);
nand U2985 (N_2985,In_194,In_2399);
and U2986 (N_2986,In_713,In_2047);
and U2987 (N_2987,In_2374,In_1482);
or U2988 (N_2988,In_2285,In_1958);
and U2989 (N_2989,In_1427,In_1328);
or U2990 (N_2990,In_2322,In_922);
nor U2991 (N_2991,In_424,In_1362);
nand U2992 (N_2992,In_10,In_2423);
nor U2993 (N_2993,In_1153,In_684);
nor U2994 (N_2994,In_2155,In_731);
or U2995 (N_2995,In_2075,In_431);
nand U2996 (N_2996,In_639,In_1699);
and U2997 (N_2997,In_1319,In_1977);
and U2998 (N_2998,In_1412,In_752);
and U2999 (N_2999,In_296,In_330);
nand U3000 (N_3000,In_1474,In_1176);
nor U3001 (N_3001,In_1022,In_1468);
or U3002 (N_3002,In_2152,In_2308);
nand U3003 (N_3003,In_1074,In_267);
nand U3004 (N_3004,In_2053,In_337);
or U3005 (N_3005,In_2074,In_2160);
or U3006 (N_3006,In_1469,In_1836);
and U3007 (N_3007,In_1883,In_838);
nand U3008 (N_3008,In_2105,In_1624);
and U3009 (N_3009,In_2009,In_24);
and U3010 (N_3010,In_168,In_48);
nor U3011 (N_3011,In_2371,In_110);
and U3012 (N_3012,In_1354,In_1665);
nor U3013 (N_3013,In_1296,In_2206);
nor U3014 (N_3014,In_636,In_953);
or U3015 (N_3015,In_2469,In_1651);
and U3016 (N_3016,In_1735,In_400);
nor U3017 (N_3017,In_562,In_1628);
nor U3018 (N_3018,In_1428,In_1049);
and U3019 (N_3019,In_176,In_1140);
nand U3020 (N_3020,In_84,In_1586);
or U3021 (N_3021,In_83,In_1897);
and U3022 (N_3022,In_1244,In_2478);
and U3023 (N_3023,In_2149,In_1676);
nor U3024 (N_3024,In_994,In_198);
nand U3025 (N_3025,In_709,In_91);
or U3026 (N_3026,In_1783,In_6);
nor U3027 (N_3027,In_1534,In_437);
and U3028 (N_3028,In_1456,In_2000);
and U3029 (N_3029,In_1444,In_979);
or U3030 (N_3030,In_423,In_2444);
or U3031 (N_3031,In_1142,In_1209);
nor U3032 (N_3032,In_159,In_2336);
xnor U3033 (N_3033,In_1192,In_1314);
nor U3034 (N_3034,In_1966,In_159);
or U3035 (N_3035,In_933,In_1327);
and U3036 (N_3036,In_224,In_904);
and U3037 (N_3037,In_2213,In_1355);
nor U3038 (N_3038,In_1450,In_310);
nor U3039 (N_3039,In_1098,In_1738);
xor U3040 (N_3040,In_339,In_389);
nor U3041 (N_3041,In_763,In_69);
nor U3042 (N_3042,In_401,In_1095);
nor U3043 (N_3043,In_2385,In_1591);
or U3044 (N_3044,In_277,In_57);
nand U3045 (N_3045,In_1473,In_151);
nand U3046 (N_3046,In_465,In_198);
nand U3047 (N_3047,In_2431,In_1934);
nor U3048 (N_3048,In_281,In_874);
or U3049 (N_3049,In_1146,In_987);
nand U3050 (N_3050,In_1355,In_1653);
or U3051 (N_3051,In_1267,In_1111);
nand U3052 (N_3052,In_816,In_1767);
nor U3053 (N_3053,In_2124,In_974);
nor U3054 (N_3054,In_1982,In_843);
nand U3055 (N_3055,In_1463,In_702);
and U3056 (N_3056,In_277,In_1083);
nor U3057 (N_3057,In_251,In_579);
or U3058 (N_3058,In_1084,In_2046);
and U3059 (N_3059,In_1812,In_536);
or U3060 (N_3060,In_2160,In_1193);
or U3061 (N_3061,In_1249,In_1498);
nor U3062 (N_3062,In_68,In_1236);
nand U3063 (N_3063,In_1377,In_320);
nand U3064 (N_3064,In_1164,In_1418);
nand U3065 (N_3065,In_695,In_262);
nand U3066 (N_3066,In_1872,In_281);
or U3067 (N_3067,In_430,In_1020);
xnor U3068 (N_3068,In_2068,In_421);
nand U3069 (N_3069,In_984,In_1029);
nand U3070 (N_3070,In_1123,In_1106);
nor U3071 (N_3071,In_1225,In_142);
and U3072 (N_3072,In_1162,In_1997);
nand U3073 (N_3073,In_411,In_1827);
or U3074 (N_3074,In_1575,In_1886);
nand U3075 (N_3075,In_1259,In_635);
nor U3076 (N_3076,In_2388,In_2070);
nor U3077 (N_3077,In_2304,In_1730);
nor U3078 (N_3078,In_570,In_1394);
and U3079 (N_3079,In_2441,In_2130);
nand U3080 (N_3080,In_306,In_836);
nand U3081 (N_3081,In_1014,In_1418);
or U3082 (N_3082,In_1525,In_804);
and U3083 (N_3083,In_775,In_868);
or U3084 (N_3084,In_831,In_189);
nand U3085 (N_3085,In_926,In_483);
nand U3086 (N_3086,In_2203,In_1811);
nor U3087 (N_3087,In_1565,In_1412);
nor U3088 (N_3088,In_1580,In_456);
and U3089 (N_3089,In_1560,In_1757);
or U3090 (N_3090,In_1584,In_1521);
nand U3091 (N_3091,In_849,In_403);
nand U3092 (N_3092,In_1429,In_1142);
and U3093 (N_3093,In_1807,In_415);
or U3094 (N_3094,In_2322,In_1228);
nor U3095 (N_3095,In_1515,In_964);
nor U3096 (N_3096,In_201,In_2311);
nand U3097 (N_3097,In_1493,In_240);
and U3098 (N_3098,In_1301,In_280);
nor U3099 (N_3099,In_1705,In_106);
nand U3100 (N_3100,In_290,In_944);
or U3101 (N_3101,In_1117,In_1860);
or U3102 (N_3102,In_128,In_1634);
nor U3103 (N_3103,In_360,In_2021);
nor U3104 (N_3104,In_1046,In_156);
nand U3105 (N_3105,In_1076,In_97);
or U3106 (N_3106,In_2389,In_1666);
or U3107 (N_3107,In_532,In_1502);
nor U3108 (N_3108,In_1441,In_1719);
xor U3109 (N_3109,In_1237,In_864);
or U3110 (N_3110,In_1213,In_76);
nor U3111 (N_3111,In_2391,In_2228);
and U3112 (N_3112,In_2223,In_2496);
nand U3113 (N_3113,In_372,In_553);
nor U3114 (N_3114,In_1374,In_1970);
nor U3115 (N_3115,In_2037,In_1870);
and U3116 (N_3116,In_1677,In_157);
or U3117 (N_3117,In_2495,In_315);
and U3118 (N_3118,In_1641,In_1509);
nor U3119 (N_3119,In_334,In_407);
nor U3120 (N_3120,In_865,In_852);
or U3121 (N_3121,In_549,In_787);
nor U3122 (N_3122,In_2368,In_1420);
nand U3123 (N_3123,In_585,In_286);
and U3124 (N_3124,In_1306,In_1257);
and U3125 (N_3125,In_201,In_1703);
and U3126 (N_3126,In_1174,In_794);
and U3127 (N_3127,In_257,In_2047);
and U3128 (N_3128,In_993,In_2200);
and U3129 (N_3129,In_2320,In_442);
nand U3130 (N_3130,In_1263,In_1880);
and U3131 (N_3131,In_378,In_338);
and U3132 (N_3132,In_1826,In_1150);
nor U3133 (N_3133,In_2026,In_2202);
nor U3134 (N_3134,In_362,In_1657);
nand U3135 (N_3135,In_2149,In_1887);
xor U3136 (N_3136,In_1436,In_2386);
and U3137 (N_3137,In_1519,In_2107);
nand U3138 (N_3138,In_1172,In_1389);
nor U3139 (N_3139,In_1994,In_2490);
nand U3140 (N_3140,In_385,In_963);
or U3141 (N_3141,In_1879,In_1779);
nor U3142 (N_3142,In_48,In_948);
nor U3143 (N_3143,In_1869,In_2355);
or U3144 (N_3144,In_28,In_219);
and U3145 (N_3145,In_722,In_933);
or U3146 (N_3146,In_2174,In_2213);
and U3147 (N_3147,In_1085,In_811);
nand U3148 (N_3148,In_1121,In_1114);
nand U3149 (N_3149,In_672,In_893);
or U3150 (N_3150,In_2324,In_949);
nor U3151 (N_3151,In_185,In_2065);
or U3152 (N_3152,In_271,In_898);
nand U3153 (N_3153,In_622,In_1056);
nand U3154 (N_3154,In_2008,In_895);
or U3155 (N_3155,In_171,In_1696);
and U3156 (N_3156,In_1354,In_186);
or U3157 (N_3157,In_1757,In_622);
nand U3158 (N_3158,In_547,In_278);
nand U3159 (N_3159,In_2006,In_1873);
nand U3160 (N_3160,In_1852,In_902);
xnor U3161 (N_3161,In_643,In_980);
nand U3162 (N_3162,In_161,In_887);
and U3163 (N_3163,In_866,In_311);
and U3164 (N_3164,In_2296,In_365);
nor U3165 (N_3165,In_644,In_904);
and U3166 (N_3166,In_1620,In_1549);
nand U3167 (N_3167,In_480,In_1497);
or U3168 (N_3168,In_1070,In_800);
nor U3169 (N_3169,In_2462,In_2235);
nor U3170 (N_3170,In_594,In_1804);
or U3171 (N_3171,In_76,In_1515);
and U3172 (N_3172,In_271,In_1145);
nor U3173 (N_3173,In_1484,In_1074);
nor U3174 (N_3174,In_1156,In_1711);
nand U3175 (N_3175,In_1634,In_1646);
and U3176 (N_3176,In_97,In_924);
or U3177 (N_3177,In_2407,In_2485);
or U3178 (N_3178,In_36,In_763);
nor U3179 (N_3179,In_2285,In_727);
nand U3180 (N_3180,In_408,In_1732);
nor U3181 (N_3181,In_2035,In_1001);
or U3182 (N_3182,In_1588,In_570);
nand U3183 (N_3183,In_537,In_2325);
nand U3184 (N_3184,In_912,In_1009);
or U3185 (N_3185,In_1899,In_1530);
and U3186 (N_3186,In_651,In_691);
and U3187 (N_3187,In_2193,In_579);
nor U3188 (N_3188,In_488,In_1460);
nand U3189 (N_3189,In_306,In_1356);
nand U3190 (N_3190,In_197,In_72);
nand U3191 (N_3191,In_714,In_2211);
nand U3192 (N_3192,In_516,In_2154);
or U3193 (N_3193,In_2074,In_438);
or U3194 (N_3194,In_640,In_619);
or U3195 (N_3195,In_818,In_156);
nor U3196 (N_3196,In_472,In_494);
and U3197 (N_3197,In_2257,In_1473);
and U3198 (N_3198,In_1312,In_336);
or U3199 (N_3199,In_683,In_1013);
or U3200 (N_3200,In_1865,In_1402);
or U3201 (N_3201,In_1952,In_1584);
nand U3202 (N_3202,In_6,In_2077);
and U3203 (N_3203,In_2323,In_1257);
and U3204 (N_3204,In_1775,In_870);
or U3205 (N_3205,In_1130,In_1045);
nand U3206 (N_3206,In_134,In_1061);
nand U3207 (N_3207,In_1951,In_1117);
and U3208 (N_3208,In_298,In_829);
nand U3209 (N_3209,In_1658,In_1246);
or U3210 (N_3210,In_229,In_1197);
nand U3211 (N_3211,In_1742,In_1972);
and U3212 (N_3212,In_871,In_1042);
nor U3213 (N_3213,In_202,In_2097);
and U3214 (N_3214,In_1405,In_2104);
nor U3215 (N_3215,In_1208,In_2342);
or U3216 (N_3216,In_313,In_1700);
nor U3217 (N_3217,In_2194,In_2003);
or U3218 (N_3218,In_2278,In_1418);
nor U3219 (N_3219,In_2251,In_2094);
nand U3220 (N_3220,In_1370,In_12);
and U3221 (N_3221,In_1057,In_758);
nand U3222 (N_3222,In_622,In_2369);
and U3223 (N_3223,In_2117,In_1976);
nor U3224 (N_3224,In_2284,In_175);
and U3225 (N_3225,In_1861,In_50);
and U3226 (N_3226,In_2051,In_21);
nor U3227 (N_3227,In_1547,In_1588);
and U3228 (N_3228,In_1869,In_82);
nor U3229 (N_3229,In_1741,In_620);
xnor U3230 (N_3230,In_1356,In_476);
or U3231 (N_3231,In_964,In_635);
nand U3232 (N_3232,In_1332,In_1837);
nand U3233 (N_3233,In_1548,In_1487);
nor U3234 (N_3234,In_1366,In_1611);
nand U3235 (N_3235,In_1332,In_679);
nand U3236 (N_3236,In_1959,In_2006);
or U3237 (N_3237,In_540,In_1592);
or U3238 (N_3238,In_630,In_1029);
xnor U3239 (N_3239,In_203,In_888);
or U3240 (N_3240,In_496,In_102);
nand U3241 (N_3241,In_704,In_2220);
nand U3242 (N_3242,In_1993,In_1043);
nand U3243 (N_3243,In_445,In_1256);
nand U3244 (N_3244,In_1873,In_385);
or U3245 (N_3245,In_79,In_1131);
nand U3246 (N_3246,In_356,In_1777);
nor U3247 (N_3247,In_2245,In_128);
and U3248 (N_3248,In_1140,In_320);
nor U3249 (N_3249,In_2329,In_1805);
and U3250 (N_3250,In_1684,In_1209);
nand U3251 (N_3251,In_2155,In_799);
and U3252 (N_3252,In_2127,In_2213);
nor U3253 (N_3253,In_1772,In_1271);
and U3254 (N_3254,In_2155,In_609);
nor U3255 (N_3255,In_1473,In_1702);
or U3256 (N_3256,In_564,In_313);
or U3257 (N_3257,In_175,In_1765);
nor U3258 (N_3258,In_160,In_750);
and U3259 (N_3259,In_1767,In_2284);
or U3260 (N_3260,In_1789,In_879);
and U3261 (N_3261,In_1337,In_104);
nor U3262 (N_3262,In_636,In_367);
and U3263 (N_3263,In_1603,In_615);
nand U3264 (N_3264,In_930,In_467);
nand U3265 (N_3265,In_2028,In_51);
and U3266 (N_3266,In_1585,In_1161);
and U3267 (N_3267,In_1756,In_957);
nor U3268 (N_3268,In_1989,In_1792);
or U3269 (N_3269,In_2084,In_916);
and U3270 (N_3270,In_243,In_1147);
or U3271 (N_3271,In_1198,In_2234);
nor U3272 (N_3272,In_2379,In_350);
and U3273 (N_3273,In_618,In_1804);
nand U3274 (N_3274,In_2214,In_2498);
nor U3275 (N_3275,In_407,In_484);
nor U3276 (N_3276,In_1381,In_2438);
nor U3277 (N_3277,In_178,In_23);
nor U3278 (N_3278,In_1873,In_453);
nor U3279 (N_3279,In_1880,In_1881);
nor U3280 (N_3280,In_710,In_781);
nor U3281 (N_3281,In_2045,In_2347);
or U3282 (N_3282,In_160,In_294);
or U3283 (N_3283,In_2458,In_1381);
or U3284 (N_3284,In_2319,In_962);
nor U3285 (N_3285,In_1040,In_1562);
nor U3286 (N_3286,In_1158,In_368);
nor U3287 (N_3287,In_1486,In_11);
nor U3288 (N_3288,In_1168,In_519);
nor U3289 (N_3289,In_1577,In_1752);
nand U3290 (N_3290,In_2303,In_1610);
nor U3291 (N_3291,In_2458,In_804);
or U3292 (N_3292,In_1269,In_1611);
or U3293 (N_3293,In_1636,In_469);
nor U3294 (N_3294,In_831,In_294);
or U3295 (N_3295,In_179,In_471);
xor U3296 (N_3296,In_163,In_1361);
or U3297 (N_3297,In_1523,In_764);
and U3298 (N_3298,In_1235,In_687);
nor U3299 (N_3299,In_1180,In_1422);
nand U3300 (N_3300,In_53,In_823);
xor U3301 (N_3301,In_1803,In_1848);
or U3302 (N_3302,In_451,In_1407);
and U3303 (N_3303,In_1099,In_381);
nor U3304 (N_3304,In_1120,In_1752);
or U3305 (N_3305,In_1296,In_498);
and U3306 (N_3306,In_2492,In_145);
nor U3307 (N_3307,In_2355,In_476);
nand U3308 (N_3308,In_973,In_396);
or U3309 (N_3309,In_1256,In_436);
nand U3310 (N_3310,In_372,In_1328);
nor U3311 (N_3311,In_1598,In_1977);
or U3312 (N_3312,In_1024,In_1345);
or U3313 (N_3313,In_2079,In_2496);
and U3314 (N_3314,In_281,In_1102);
or U3315 (N_3315,In_889,In_1813);
or U3316 (N_3316,In_2061,In_1527);
and U3317 (N_3317,In_1905,In_2060);
or U3318 (N_3318,In_225,In_1684);
xnor U3319 (N_3319,In_822,In_1359);
or U3320 (N_3320,In_2443,In_1078);
nand U3321 (N_3321,In_753,In_312);
or U3322 (N_3322,In_1392,In_1073);
nand U3323 (N_3323,In_1893,In_1259);
nor U3324 (N_3324,In_729,In_260);
nand U3325 (N_3325,In_415,In_871);
and U3326 (N_3326,In_1499,In_2021);
and U3327 (N_3327,In_1926,In_852);
nand U3328 (N_3328,In_755,In_1831);
nand U3329 (N_3329,In_1355,In_971);
nand U3330 (N_3330,In_1941,In_2346);
nand U3331 (N_3331,In_457,In_1551);
and U3332 (N_3332,In_160,In_1525);
or U3333 (N_3333,In_2448,In_1828);
or U3334 (N_3334,In_350,In_2321);
nand U3335 (N_3335,In_2104,In_1990);
and U3336 (N_3336,In_1184,In_253);
or U3337 (N_3337,In_2236,In_1332);
nand U3338 (N_3338,In_726,In_1550);
nand U3339 (N_3339,In_2122,In_1816);
nor U3340 (N_3340,In_2351,In_1210);
and U3341 (N_3341,In_1705,In_1930);
and U3342 (N_3342,In_660,In_1979);
nand U3343 (N_3343,In_14,In_4);
nor U3344 (N_3344,In_1701,In_1572);
and U3345 (N_3345,In_318,In_1762);
and U3346 (N_3346,In_2151,In_2343);
or U3347 (N_3347,In_31,In_1180);
nor U3348 (N_3348,In_1351,In_1914);
nor U3349 (N_3349,In_2201,In_1474);
or U3350 (N_3350,In_1060,In_598);
nor U3351 (N_3351,In_1579,In_1090);
nand U3352 (N_3352,In_95,In_2386);
and U3353 (N_3353,In_1521,In_1277);
or U3354 (N_3354,In_1322,In_2238);
and U3355 (N_3355,In_525,In_993);
or U3356 (N_3356,In_115,In_1599);
and U3357 (N_3357,In_2362,In_429);
or U3358 (N_3358,In_1018,In_1985);
nand U3359 (N_3359,In_968,In_1046);
nor U3360 (N_3360,In_555,In_3);
nand U3361 (N_3361,In_2475,In_1426);
nor U3362 (N_3362,In_963,In_1516);
and U3363 (N_3363,In_536,In_21);
nor U3364 (N_3364,In_1813,In_2282);
or U3365 (N_3365,In_1104,In_1715);
nand U3366 (N_3366,In_2,In_1675);
and U3367 (N_3367,In_1095,In_1723);
nand U3368 (N_3368,In_1947,In_757);
nand U3369 (N_3369,In_847,In_616);
nand U3370 (N_3370,In_331,In_2373);
nor U3371 (N_3371,In_2038,In_666);
nor U3372 (N_3372,In_552,In_967);
nand U3373 (N_3373,In_820,In_2445);
and U3374 (N_3374,In_1638,In_124);
nand U3375 (N_3375,In_1088,In_1771);
or U3376 (N_3376,In_408,In_2233);
or U3377 (N_3377,In_599,In_2443);
nor U3378 (N_3378,In_1821,In_1125);
and U3379 (N_3379,In_718,In_16);
nor U3380 (N_3380,In_479,In_60);
and U3381 (N_3381,In_2463,In_31);
or U3382 (N_3382,In_1428,In_597);
and U3383 (N_3383,In_640,In_1120);
and U3384 (N_3384,In_1444,In_745);
nand U3385 (N_3385,In_323,In_2259);
and U3386 (N_3386,In_2375,In_1774);
or U3387 (N_3387,In_350,In_130);
and U3388 (N_3388,In_2343,In_2040);
or U3389 (N_3389,In_2498,In_1611);
or U3390 (N_3390,In_13,In_18);
or U3391 (N_3391,In_189,In_1543);
and U3392 (N_3392,In_913,In_1124);
nor U3393 (N_3393,In_667,In_1718);
nand U3394 (N_3394,In_1849,In_1639);
nand U3395 (N_3395,In_2242,In_119);
nand U3396 (N_3396,In_2011,In_2194);
and U3397 (N_3397,In_238,In_363);
and U3398 (N_3398,In_175,In_2226);
and U3399 (N_3399,In_1837,In_1314);
and U3400 (N_3400,In_2187,In_280);
nand U3401 (N_3401,In_796,In_1286);
and U3402 (N_3402,In_2223,In_1700);
or U3403 (N_3403,In_1498,In_347);
and U3404 (N_3404,In_475,In_1707);
and U3405 (N_3405,In_841,In_2334);
nand U3406 (N_3406,In_998,In_920);
nand U3407 (N_3407,In_926,In_152);
nand U3408 (N_3408,In_294,In_2085);
nand U3409 (N_3409,In_1179,In_1369);
or U3410 (N_3410,In_2178,In_911);
nor U3411 (N_3411,In_1084,In_688);
nor U3412 (N_3412,In_270,In_846);
and U3413 (N_3413,In_1874,In_860);
nand U3414 (N_3414,In_1339,In_2384);
nand U3415 (N_3415,In_1234,In_1262);
or U3416 (N_3416,In_177,In_2094);
nor U3417 (N_3417,In_2096,In_1550);
nor U3418 (N_3418,In_346,In_2242);
nor U3419 (N_3419,In_2486,In_2201);
nand U3420 (N_3420,In_2093,In_1222);
nand U3421 (N_3421,In_1545,In_262);
nor U3422 (N_3422,In_955,In_1605);
and U3423 (N_3423,In_1288,In_495);
or U3424 (N_3424,In_1606,In_1519);
or U3425 (N_3425,In_1475,In_241);
nand U3426 (N_3426,In_492,In_608);
or U3427 (N_3427,In_1465,In_2172);
or U3428 (N_3428,In_1700,In_1462);
nand U3429 (N_3429,In_1034,In_783);
nor U3430 (N_3430,In_117,In_1020);
or U3431 (N_3431,In_2207,In_574);
nand U3432 (N_3432,In_1931,In_879);
or U3433 (N_3433,In_1181,In_282);
xnor U3434 (N_3434,In_1521,In_140);
nor U3435 (N_3435,In_821,In_1953);
and U3436 (N_3436,In_411,In_1106);
nor U3437 (N_3437,In_1520,In_1911);
nor U3438 (N_3438,In_743,In_2037);
nand U3439 (N_3439,In_2345,In_2173);
or U3440 (N_3440,In_2146,In_2098);
and U3441 (N_3441,In_1314,In_426);
and U3442 (N_3442,In_1904,In_1759);
nand U3443 (N_3443,In_2343,In_2045);
nand U3444 (N_3444,In_2272,In_318);
and U3445 (N_3445,In_477,In_1821);
and U3446 (N_3446,In_1071,In_164);
nand U3447 (N_3447,In_37,In_942);
or U3448 (N_3448,In_295,In_2389);
or U3449 (N_3449,In_827,In_2088);
nor U3450 (N_3450,In_2464,In_1222);
and U3451 (N_3451,In_2124,In_1653);
or U3452 (N_3452,In_992,In_2392);
nor U3453 (N_3453,In_1506,In_1003);
and U3454 (N_3454,In_1639,In_2031);
and U3455 (N_3455,In_1896,In_2060);
and U3456 (N_3456,In_948,In_2297);
or U3457 (N_3457,In_1893,In_1216);
nor U3458 (N_3458,In_894,In_1873);
nor U3459 (N_3459,In_1010,In_1119);
nand U3460 (N_3460,In_1460,In_1795);
nand U3461 (N_3461,In_421,In_346);
nand U3462 (N_3462,In_2492,In_254);
or U3463 (N_3463,In_91,In_293);
and U3464 (N_3464,In_66,In_2315);
and U3465 (N_3465,In_2349,In_1991);
and U3466 (N_3466,In_2041,In_1385);
or U3467 (N_3467,In_444,In_732);
or U3468 (N_3468,In_2463,In_1150);
and U3469 (N_3469,In_1588,In_344);
and U3470 (N_3470,In_282,In_2242);
nand U3471 (N_3471,In_2054,In_956);
or U3472 (N_3472,In_1516,In_1355);
nand U3473 (N_3473,In_2486,In_1503);
nand U3474 (N_3474,In_2493,In_10);
nand U3475 (N_3475,In_319,In_2379);
nand U3476 (N_3476,In_378,In_787);
or U3477 (N_3477,In_550,In_1716);
nand U3478 (N_3478,In_2131,In_733);
and U3479 (N_3479,In_2274,In_119);
xor U3480 (N_3480,In_1531,In_205);
nor U3481 (N_3481,In_2005,In_1994);
and U3482 (N_3482,In_1430,In_2113);
nand U3483 (N_3483,In_2076,In_1430);
nand U3484 (N_3484,In_2451,In_2456);
or U3485 (N_3485,In_925,In_1096);
or U3486 (N_3486,In_1844,In_388);
nand U3487 (N_3487,In_1035,In_1609);
or U3488 (N_3488,In_1033,In_484);
nand U3489 (N_3489,In_1028,In_2190);
and U3490 (N_3490,In_2409,In_79);
nand U3491 (N_3491,In_2488,In_579);
and U3492 (N_3492,In_2042,In_2084);
and U3493 (N_3493,In_1380,In_226);
nor U3494 (N_3494,In_1271,In_549);
or U3495 (N_3495,In_1272,In_2259);
or U3496 (N_3496,In_2178,In_1689);
nor U3497 (N_3497,In_2019,In_2380);
nand U3498 (N_3498,In_1596,In_578);
nor U3499 (N_3499,In_7,In_481);
and U3500 (N_3500,In_808,In_2377);
or U3501 (N_3501,In_764,In_467);
nand U3502 (N_3502,In_434,In_158);
and U3503 (N_3503,In_970,In_1630);
nor U3504 (N_3504,In_422,In_2185);
nor U3505 (N_3505,In_1037,In_1729);
nor U3506 (N_3506,In_2378,In_292);
nor U3507 (N_3507,In_1172,In_2231);
or U3508 (N_3508,In_1643,In_1248);
nand U3509 (N_3509,In_2183,In_612);
or U3510 (N_3510,In_1546,In_1548);
nor U3511 (N_3511,In_2212,In_2252);
nor U3512 (N_3512,In_185,In_482);
or U3513 (N_3513,In_768,In_960);
nand U3514 (N_3514,In_523,In_1923);
and U3515 (N_3515,In_2224,In_507);
or U3516 (N_3516,In_1107,In_583);
nor U3517 (N_3517,In_830,In_323);
nor U3518 (N_3518,In_450,In_2363);
and U3519 (N_3519,In_1312,In_1138);
nand U3520 (N_3520,In_1407,In_1968);
or U3521 (N_3521,In_497,In_573);
or U3522 (N_3522,In_2498,In_1936);
nand U3523 (N_3523,In_112,In_878);
and U3524 (N_3524,In_508,In_670);
and U3525 (N_3525,In_2241,In_1933);
nor U3526 (N_3526,In_669,In_1206);
or U3527 (N_3527,In_1265,In_1965);
nand U3528 (N_3528,In_1113,In_1248);
xor U3529 (N_3529,In_637,In_2040);
nand U3530 (N_3530,In_1504,In_1652);
or U3531 (N_3531,In_2487,In_270);
nand U3532 (N_3532,In_1814,In_696);
nor U3533 (N_3533,In_829,In_1697);
and U3534 (N_3534,In_2219,In_1505);
xnor U3535 (N_3535,In_420,In_1399);
or U3536 (N_3536,In_1263,In_122);
nor U3537 (N_3537,In_1586,In_1363);
or U3538 (N_3538,In_2178,In_915);
nand U3539 (N_3539,In_2306,In_1351);
nor U3540 (N_3540,In_1348,In_1173);
nor U3541 (N_3541,In_271,In_521);
nand U3542 (N_3542,In_1996,In_1904);
nand U3543 (N_3543,In_478,In_2254);
or U3544 (N_3544,In_839,In_163);
nor U3545 (N_3545,In_779,In_2417);
nand U3546 (N_3546,In_1899,In_761);
nor U3547 (N_3547,In_563,In_2270);
or U3548 (N_3548,In_1751,In_1774);
nor U3549 (N_3549,In_186,In_566);
nor U3550 (N_3550,In_2393,In_1427);
and U3551 (N_3551,In_1411,In_508);
nor U3552 (N_3552,In_2390,In_1959);
or U3553 (N_3553,In_1977,In_1156);
nand U3554 (N_3554,In_1159,In_2017);
nor U3555 (N_3555,In_860,In_2409);
nand U3556 (N_3556,In_1885,In_377);
or U3557 (N_3557,In_525,In_1680);
xor U3558 (N_3558,In_1717,In_1543);
nand U3559 (N_3559,In_655,In_1523);
or U3560 (N_3560,In_1373,In_290);
nand U3561 (N_3561,In_1628,In_1117);
nand U3562 (N_3562,In_2224,In_1800);
nor U3563 (N_3563,In_982,In_978);
nand U3564 (N_3564,In_1126,In_1014);
or U3565 (N_3565,In_1920,In_1389);
nand U3566 (N_3566,In_29,In_1046);
or U3567 (N_3567,In_35,In_522);
and U3568 (N_3568,In_233,In_2320);
nor U3569 (N_3569,In_425,In_339);
nand U3570 (N_3570,In_1209,In_478);
nor U3571 (N_3571,In_2127,In_130);
nor U3572 (N_3572,In_162,In_2241);
and U3573 (N_3573,In_2290,In_609);
nand U3574 (N_3574,In_2436,In_2102);
and U3575 (N_3575,In_1346,In_1874);
or U3576 (N_3576,In_1651,In_1424);
nand U3577 (N_3577,In_243,In_367);
or U3578 (N_3578,In_1216,In_1732);
or U3579 (N_3579,In_397,In_371);
and U3580 (N_3580,In_1255,In_563);
and U3581 (N_3581,In_168,In_1709);
and U3582 (N_3582,In_481,In_103);
nor U3583 (N_3583,In_1805,In_612);
nor U3584 (N_3584,In_1629,In_1621);
and U3585 (N_3585,In_1857,In_2033);
and U3586 (N_3586,In_511,In_687);
nor U3587 (N_3587,In_1421,In_1174);
and U3588 (N_3588,In_1001,In_2151);
or U3589 (N_3589,In_832,In_929);
and U3590 (N_3590,In_2167,In_1993);
and U3591 (N_3591,In_1998,In_2031);
nand U3592 (N_3592,In_357,In_781);
nor U3593 (N_3593,In_871,In_1385);
and U3594 (N_3594,In_1331,In_967);
and U3595 (N_3595,In_1134,In_56);
nor U3596 (N_3596,In_166,In_32);
nand U3597 (N_3597,In_1651,In_1855);
nor U3598 (N_3598,In_1815,In_1771);
and U3599 (N_3599,In_1071,In_2052);
xor U3600 (N_3600,In_1752,In_1925);
or U3601 (N_3601,In_243,In_995);
and U3602 (N_3602,In_1058,In_2156);
nor U3603 (N_3603,In_2281,In_1276);
or U3604 (N_3604,In_709,In_1218);
nor U3605 (N_3605,In_1685,In_1397);
nor U3606 (N_3606,In_513,In_1391);
nand U3607 (N_3607,In_827,In_1821);
or U3608 (N_3608,In_2349,In_886);
nand U3609 (N_3609,In_1685,In_7);
nor U3610 (N_3610,In_1509,In_1290);
nand U3611 (N_3611,In_1270,In_945);
and U3612 (N_3612,In_1951,In_1507);
and U3613 (N_3613,In_1766,In_1441);
nand U3614 (N_3614,In_2080,In_1778);
nor U3615 (N_3615,In_1155,In_863);
and U3616 (N_3616,In_1965,In_2160);
nor U3617 (N_3617,In_404,In_321);
nor U3618 (N_3618,In_607,In_2364);
nor U3619 (N_3619,In_561,In_312);
nor U3620 (N_3620,In_931,In_1588);
or U3621 (N_3621,In_630,In_2160);
nor U3622 (N_3622,In_931,In_2346);
and U3623 (N_3623,In_2295,In_153);
and U3624 (N_3624,In_327,In_1588);
nor U3625 (N_3625,In_461,In_515);
nor U3626 (N_3626,In_2410,In_1797);
and U3627 (N_3627,In_1639,In_126);
and U3628 (N_3628,In_2431,In_1912);
nand U3629 (N_3629,In_1734,In_1775);
and U3630 (N_3630,In_416,In_822);
or U3631 (N_3631,In_2366,In_1536);
nor U3632 (N_3632,In_490,In_2337);
nor U3633 (N_3633,In_2174,In_2204);
and U3634 (N_3634,In_716,In_397);
or U3635 (N_3635,In_1926,In_866);
and U3636 (N_3636,In_1554,In_2155);
and U3637 (N_3637,In_342,In_1635);
nand U3638 (N_3638,In_1251,In_2371);
nor U3639 (N_3639,In_565,In_1824);
nand U3640 (N_3640,In_69,In_1737);
nand U3641 (N_3641,In_1030,In_1453);
or U3642 (N_3642,In_115,In_995);
nand U3643 (N_3643,In_903,In_1379);
or U3644 (N_3644,In_61,In_501);
or U3645 (N_3645,In_1422,In_693);
nor U3646 (N_3646,In_2255,In_193);
and U3647 (N_3647,In_1002,In_2097);
nand U3648 (N_3648,In_662,In_1530);
nand U3649 (N_3649,In_1321,In_2129);
nand U3650 (N_3650,In_2349,In_1696);
and U3651 (N_3651,In_2162,In_2209);
nor U3652 (N_3652,In_601,In_2492);
or U3653 (N_3653,In_1249,In_1883);
and U3654 (N_3654,In_1189,In_675);
nor U3655 (N_3655,In_53,In_1501);
nand U3656 (N_3656,In_2053,In_705);
and U3657 (N_3657,In_1565,In_1361);
or U3658 (N_3658,In_200,In_629);
and U3659 (N_3659,In_1028,In_857);
and U3660 (N_3660,In_827,In_1284);
nor U3661 (N_3661,In_271,In_579);
nand U3662 (N_3662,In_350,In_742);
nor U3663 (N_3663,In_350,In_1068);
and U3664 (N_3664,In_1000,In_704);
xnor U3665 (N_3665,In_2333,In_1519);
nand U3666 (N_3666,In_587,In_27);
nand U3667 (N_3667,In_2005,In_1538);
and U3668 (N_3668,In_605,In_2160);
nand U3669 (N_3669,In_1431,In_1548);
or U3670 (N_3670,In_223,In_55);
and U3671 (N_3671,In_687,In_2458);
nor U3672 (N_3672,In_1159,In_2372);
nand U3673 (N_3673,In_1951,In_2355);
and U3674 (N_3674,In_2427,In_34);
or U3675 (N_3675,In_1795,In_721);
nor U3676 (N_3676,In_1495,In_1668);
nand U3677 (N_3677,In_1251,In_1414);
nor U3678 (N_3678,In_2054,In_1259);
and U3679 (N_3679,In_1953,In_127);
and U3680 (N_3680,In_59,In_1564);
nor U3681 (N_3681,In_269,In_2435);
and U3682 (N_3682,In_2019,In_1560);
nand U3683 (N_3683,In_26,In_368);
or U3684 (N_3684,In_1726,In_1297);
or U3685 (N_3685,In_1647,In_976);
nand U3686 (N_3686,In_1034,In_525);
or U3687 (N_3687,In_307,In_2420);
and U3688 (N_3688,In_111,In_1147);
nand U3689 (N_3689,In_1991,In_2051);
nand U3690 (N_3690,In_1740,In_726);
and U3691 (N_3691,In_2000,In_867);
and U3692 (N_3692,In_756,In_291);
nor U3693 (N_3693,In_524,In_2394);
or U3694 (N_3694,In_63,In_1812);
and U3695 (N_3695,In_2312,In_650);
nor U3696 (N_3696,In_46,In_127);
and U3697 (N_3697,In_4,In_817);
or U3698 (N_3698,In_974,In_1430);
and U3699 (N_3699,In_1474,In_960);
nand U3700 (N_3700,In_1538,In_1418);
nand U3701 (N_3701,In_891,In_647);
nand U3702 (N_3702,In_152,In_2136);
and U3703 (N_3703,In_2204,In_2117);
nand U3704 (N_3704,In_2131,In_1315);
or U3705 (N_3705,In_2261,In_1713);
and U3706 (N_3706,In_1845,In_209);
nand U3707 (N_3707,In_371,In_2472);
or U3708 (N_3708,In_2227,In_1497);
and U3709 (N_3709,In_1755,In_1436);
nand U3710 (N_3710,In_475,In_1775);
nor U3711 (N_3711,In_611,In_2479);
or U3712 (N_3712,In_685,In_597);
or U3713 (N_3713,In_1446,In_2152);
and U3714 (N_3714,In_984,In_2291);
nand U3715 (N_3715,In_1653,In_1650);
and U3716 (N_3716,In_933,In_190);
nand U3717 (N_3717,In_1704,In_1777);
or U3718 (N_3718,In_16,In_1706);
nand U3719 (N_3719,In_290,In_367);
or U3720 (N_3720,In_1020,In_345);
nand U3721 (N_3721,In_2329,In_2354);
or U3722 (N_3722,In_433,In_149);
nor U3723 (N_3723,In_1190,In_105);
nand U3724 (N_3724,In_1903,In_880);
or U3725 (N_3725,In_650,In_378);
and U3726 (N_3726,In_1882,In_2319);
and U3727 (N_3727,In_1071,In_2130);
and U3728 (N_3728,In_7,In_2454);
nand U3729 (N_3729,In_1634,In_158);
nor U3730 (N_3730,In_2498,In_477);
nor U3731 (N_3731,In_2222,In_772);
nand U3732 (N_3732,In_2196,In_1788);
nor U3733 (N_3733,In_1840,In_653);
nand U3734 (N_3734,In_1952,In_995);
and U3735 (N_3735,In_75,In_1599);
or U3736 (N_3736,In_86,In_369);
and U3737 (N_3737,In_953,In_2386);
and U3738 (N_3738,In_1544,In_2335);
or U3739 (N_3739,In_2202,In_799);
nand U3740 (N_3740,In_1327,In_2037);
and U3741 (N_3741,In_1214,In_855);
or U3742 (N_3742,In_2344,In_741);
and U3743 (N_3743,In_1571,In_2056);
nor U3744 (N_3744,In_2133,In_1266);
and U3745 (N_3745,In_1335,In_2237);
nand U3746 (N_3746,In_270,In_1804);
and U3747 (N_3747,In_236,In_1371);
nor U3748 (N_3748,In_419,In_1159);
nor U3749 (N_3749,In_1676,In_189);
nand U3750 (N_3750,In_825,In_1159);
and U3751 (N_3751,In_1494,In_2350);
nand U3752 (N_3752,In_455,In_832);
nand U3753 (N_3753,In_574,In_1600);
or U3754 (N_3754,In_1503,In_1139);
nor U3755 (N_3755,In_1649,In_1862);
nand U3756 (N_3756,In_435,In_1632);
or U3757 (N_3757,In_1577,In_1640);
nor U3758 (N_3758,In_7,In_1196);
nor U3759 (N_3759,In_1458,In_2316);
and U3760 (N_3760,In_1087,In_1080);
nor U3761 (N_3761,In_2495,In_2042);
or U3762 (N_3762,In_2105,In_48);
nand U3763 (N_3763,In_122,In_760);
nand U3764 (N_3764,In_1673,In_698);
and U3765 (N_3765,In_1924,In_1142);
and U3766 (N_3766,In_1491,In_1831);
and U3767 (N_3767,In_2225,In_970);
and U3768 (N_3768,In_624,In_788);
nor U3769 (N_3769,In_93,In_1672);
or U3770 (N_3770,In_83,In_205);
or U3771 (N_3771,In_1410,In_2221);
or U3772 (N_3772,In_721,In_2263);
nand U3773 (N_3773,In_2125,In_2170);
nand U3774 (N_3774,In_1619,In_208);
or U3775 (N_3775,In_938,In_562);
and U3776 (N_3776,In_1490,In_352);
and U3777 (N_3777,In_1696,In_956);
or U3778 (N_3778,In_2110,In_1557);
or U3779 (N_3779,In_1507,In_1633);
nand U3780 (N_3780,In_2129,In_1035);
nor U3781 (N_3781,In_1761,In_630);
nand U3782 (N_3782,In_574,In_68);
nor U3783 (N_3783,In_58,In_1394);
and U3784 (N_3784,In_1019,In_1120);
nor U3785 (N_3785,In_466,In_1416);
and U3786 (N_3786,In_1274,In_1247);
and U3787 (N_3787,In_1188,In_1769);
and U3788 (N_3788,In_440,In_879);
nand U3789 (N_3789,In_227,In_2166);
or U3790 (N_3790,In_319,In_903);
nand U3791 (N_3791,In_1584,In_368);
nand U3792 (N_3792,In_1653,In_2199);
nor U3793 (N_3793,In_945,In_2316);
and U3794 (N_3794,In_1676,In_441);
and U3795 (N_3795,In_1115,In_1686);
or U3796 (N_3796,In_904,In_1713);
and U3797 (N_3797,In_19,In_2361);
nor U3798 (N_3798,In_2177,In_2330);
nor U3799 (N_3799,In_407,In_2347);
nand U3800 (N_3800,In_1936,In_2245);
or U3801 (N_3801,In_2276,In_1083);
nor U3802 (N_3802,In_1771,In_235);
nor U3803 (N_3803,In_166,In_1881);
or U3804 (N_3804,In_676,In_541);
nand U3805 (N_3805,In_758,In_124);
nand U3806 (N_3806,In_1671,In_563);
or U3807 (N_3807,In_900,In_1810);
and U3808 (N_3808,In_1224,In_974);
nand U3809 (N_3809,In_1407,In_370);
or U3810 (N_3810,In_1933,In_108);
nand U3811 (N_3811,In_301,In_1010);
and U3812 (N_3812,In_1735,In_1196);
or U3813 (N_3813,In_1147,In_1399);
and U3814 (N_3814,In_1778,In_222);
nand U3815 (N_3815,In_1027,In_780);
nand U3816 (N_3816,In_245,In_517);
or U3817 (N_3817,In_11,In_2188);
and U3818 (N_3818,In_2185,In_1350);
nand U3819 (N_3819,In_102,In_80);
nand U3820 (N_3820,In_445,In_23);
or U3821 (N_3821,In_2437,In_500);
nand U3822 (N_3822,In_1217,In_679);
nor U3823 (N_3823,In_2023,In_1553);
nor U3824 (N_3824,In_1162,In_2282);
and U3825 (N_3825,In_44,In_457);
nand U3826 (N_3826,In_543,In_2352);
nor U3827 (N_3827,In_374,In_1297);
and U3828 (N_3828,In_922,In_1976);
nand U3829 (N_3829,In_2496,In_1130);
nand U3830 (N_3830,In_1279,In_1462);
and U3831 (N_3831,In_2375,In_1156);
or U3832 (N_3832,In_1839,In_2494);
nand U3833 (N_3833,In_1636,In_881);
nand U3834 (N_3834,In_1893,In_1293);
or U3835 (N_3835,In_1683,In_40);
or U3836 (N_3836,In_2371,In_1451);
nand U3837 (N_3837,In_2306,In_290);
nor U3838 (N_3838,In_332,In_193);
or U3839 (N_3839,In_1646,In_1262);
or U3840 (N_3840,In_822,In_1147);
and U3841 (N_3841,In_1848,In_46);
and U3842 (N_3842,In_1293,In_1390);
nand U3843 (N_3843,In_1187,In_2342);
or U3844 (N_3844,In_2257,In_911);
and U3845 (N_3845,In_2000,In_1411);
nand U3846 (N_3846,In_2431,In_1449);
and U3847 (N_3847,In_895,In_1218);
and U3848 (N_3848,In_2364,In_939);
and U3849 (N_3849,In_604,In_307);
and U3850 (N_3850,In_1314,In_2408);
nand U3851 (N_3851,In_592,In_703);
nor U3852 (N_3852,In_1916,In_1808);
nor U3853 (N_3853,In_716,In_2056);
and U3854 (N_3854,In_2073,In_144);
nor U3855 (N_3855,In_1897,In_1953);
nor U3856 (N_3856,In_1759,In_1374);
nand U3857 (N_3857,In_183,In_1203);
nand U3858 (N_3858,In_831,In_2393);
nor U3859 (N_3859,In_1352,In_31);
nor U3860 (N_3860,In_1903,In_1763);
nand U3861 (N_3861,In_785,In_950);
nor U3862 (N_3862,In_2447,In_770);
nand U3863 (N_3863,In_796,In_1150);
or U3864 (N_3864,In_1640,In_432);
or U3865 (N_3865,In_524,In_120);
nand U3866 (N_3866,In_241,In_1171);
nand U3867 (N_3867,In_953,In_1698);
or U3868 (N_3868,In_2283,In_1523);
and U3869 (N_3869,In_1410,In_2017);
nor U3870 (N_3870,In_1506,In_551);
and U3871 (N_3871,In_76,In_89);
nor U3872 (N_3872,In_386,In_715);
and U3873 (N_3873,In_1924,In_533);
and U3874 (N_3874,In_2268,In_2020);
or U3875 (N_3875,In_1696,In_1601);
and U3876 (N_3876,In_840,In_2069);
nor U3877 (N_3877,In_77,In_147);
nor U3878 (N_3878,In_798,In_719);
nor U3879 (N_3879,In_1835,In_665);
nand U3880 (N_3880,In_1732,In_1841);
nand U3881 (N_3881,In_1860,In_37);
or U3882 (N_3882,In_953,In_315);
nand U3883 (N_3883,In_949,In_854);
nor U3884 (N_3884,In_570,In_1334);
nor U3885 (N_3885,In_748,In_456);
or U3886 (N_3886,In_1818,In_1388);
nand U3887 (N_3887,In_696,In_1011);
nand U3888 (N_3888,In_532,In_794);
nor U3889 (N_3889,In_2195,In_2263);
and U3890 (N_3890,In_346,In_599);
nand U3891 (N_3891,In_2037,In_874);
and U3892 (N_3892,In_568,In_702);
nand U3893 (N_3893,In_39,In_2269);
nand U3894 (N_3894,In_1564,In_456);
nor U3895 (N_3895,In_281,In_947);
nand U3896 (N_3896,In_829,In_1266);
nand U3897 (N_3897,In_911,In_2021);
nor U3898 (N_3898,In_2442,In_121);
nor U3899 (N_3899,In_2352,In_148);
and U3900 (N_3900,In_1290,In_1714);
nand U3901 (N_3901,In_1446,In_533);
and U3902 (N_3902,In_465,In_924);
or U3903 (N_3903,In_1590,In_146);
nor U3904 (N_3904,In_1992,In_617);
or U3905 (N_3905,In_160,In_1075);
or U3906 (N_3906,In_1878,In_10);
or U3907 (N_3907,In_269,In_1786);
or U3908 (N_3908,In_2331,In_58);
nand U3909 (N_3909,In_1807,In_2305);
and U3910 (N_3910,In_1035,In_185);
nor U3911 (N_3911,In_666,In_82);
nor U3912 (N_3912,In_763,In_1973);
or U3913 (N_3913,In_2019,In_1072);
nand U3914 (N_3914,In_651,In_1128);
nand U3915 (N_3915,In_1020,In_340);
nor U3916 (N_3916,In_1180,In_41);
or U3917 (N_3917,In_1318,In_1460);
and U3918 (N_3918,In_389,In_1555);
and U3919 (N_3919,In_2004,In_200);
and U3920 (N_3920,In_2397,In_1362);
nor U3921 (N_3921,In_1735,In_1151);
nand U3922 (N_3922,In_2258,In_1721);
and U3923 (N_3923,In_1988,In_189);
nand U3924 (N_3924,In_2411,In_732);
xor U3925 (N_3925,In_1163,In_1148);
nand U3926 (N_3926,In_399,In_1526);
or U3927 (N_3927,In_2264,In_549);
nor U3928 (N_3928,In_1115,In_2254);
and U3929 (N_3929,In_577,In_1458);
and U3930 (N_3930,In_1457,In_431);
nor U3931 (N_3931,In_932,In_1465);
nand U3932 (N_3932,In_2435,In_2206);
or U3933 (N_3933,In_1193,In_241);
nor U3934 (N_3934,In_850,In_967);
or U3935 (N_3935,In_2308,In_500);
nor U3936 (N_3936,In_1630,In_1935);
or U3937 (N_3937,In_2078,In_1167);
nand U3938 (N_3938,In_925,In_2313);
and U3939 (N_3939,In_520,In_825);
nor U3940 (N_3940,In_187,In_2034);
and U3941 (N_3941,In_1517,In_698);
or U3942 (N_3942,In_2026,In_440);
or U3943 (N_3943,In_610,In_913);
nor U3944 (N_3944,In_775,In_780);
nor U3945 (N_3945,In_1186,In_1871);
nand U3946 (N_3946,In_1960,In_2303);
nor U3947 (N_3947,In_1256,In_736);
or U3948 (N_3948,In_1976,In_1578);
and U3949 (N_3949,In_183,In_1053);
and U3950 (N_3950,In_706,In_2022);
xnor U3951 (N_3951,In_967,In_1976);
nor U3952 (N_3952,In_1164,In_1830);
nor U3953 (N_3953,In_1211,In_1932);
or U3954 (N_3954,In_953,In_1749);
and U3955 (N_3955,In_2050,In_2071);
nor U3956 (N_3956,In_1103,In_1059);
and U3957 (N_3957,In_244,In_1628);
or U3958 (N_3958,In_1185,In_944);
nor U3959 (N_3959,In_1994,In_457);
nor U3960 (N_3960,In_1989,In_506);
nor U3961 (N_3961,In_1916,In_249);
or U3962 (N_3962,In_59,In_676);
nor U3963 (N_3963,In_2049,In_681);
nor U3964 (N_3964,In_2151,In_1915);
nand U3965 (N_3965,In_660,In_1648);
nor U3966 (N_3966,In_544,In_2414);
or U3967 (N_3967,In_1734,In_979);
nand U3968 (N_3968,In_2421,In_60);
nand U3969 (N_3969,In_481,In_1883);
nor U3970 (N_3970,In_253,In_322);
nand U3971 (N_3971,In_1999,In_2230);
or U3972 (N_3972,In_1274,In_1906);
and U3973 (N_3973,In_2340,In_84);
nor U3974 (N_3974,In_934,In_2167);
nand U3975 (N_3975,In_2496,In_667);
or U3976 (N_3976,In_1925,In_1466);
nor U3977 (N_3977,In_409,In_1333);
or U3978 (N_3978,In_2182,In_2078);
or U3979 (N_3979,In_1048,In_1293);
nand U3980 (N_3980,In_820,In_1086);
nor U3981 (N_3981,In_1540,In_169);
nor U3982 (N_3982,In_1058,In_2235);
nor U3983 (N_3983,In_2037,In_612);
nor U3984 (N_3984,In_10,In_140);
nand U3985 (N_3985,In_573,In_1048);
nor U3986 (N_3986,In_1065,In_21);
or U3987 (N_3987,In_2173,In_134);
and U3988 (N_3988,In_995,In_1342);
nor U3989 (N_3989,In_2246,In_1318);
or U3990 (N_3990,In_1640,In_973);
nand U3991 (N_3991,In_1442,In_1556);
and U3992 (N_3992,In_477,In_1784);
nand U3993 (N_3993,In_2340,In_2492);
nand U3994 (N_3994,In_1565,In_1390);
nand U3995 (N_3995,In_2275,In_828);
nand U3996 (N_3996,In_1429,In_812);
nor U3997 (N_3997,In_1416,In_1354);
or U3998 (N_3998,In_281,In_1439);
nor U3999 (N_3999,In_1914,In_301);
nand U4000 (N_4000,In_701,In_1242);
nand U4001 (N_4001,In_1384,In_1322);
nand U4002 (N_4002,In_484,In_83);
or U4003 (N_4003,In_2329,In_148);
and U4004 (N_4004,In_774,In_2269);
or U4005 (N_4005,In_667,In_2241);
nand U4006 (N_4006,In_1174,In_1319);
nor U4007 (N_4007,In_573,In_35);
and U4008 (N_4008,In_2116,In_1664);
nor U4009 (N_4009,In_2316,In_1062);
or U4010 (N_4010,In_1318,In_376);
nand U4011 (N_4011,In_1081,In_1211);
nor U4012 (N_4012,In_171,In_1222);
nor U4013 (N_4013,In_1777,In_1805);
nand U4014 (N_4014,In_494,In_484);
nand U4015 (N_4015,In_898,In_39);
nand U4016 (N_4016,In_101,In_1571);
or U4017 (N_4017,In_795,In_2227);
nand U4018 (N_4018,In_1902,In_329);
and U4019 (N_4019,In_820,In_1867);
and U4020 (N_4020,In_897,In_366);
and U4021 (N_4021,In_2349,In_52);
and U4022 (N_4022,In_1618,In_561);
nor U4023 (N_4023,In_1565,In_2292);
nor U4024 (N_4024,In_2217,In_1234);
and U4025 (N_4025,In_304,In_1998);
nand U4026 (N_4026,In_1019,In_885);
nor U4027 (N_4027,In_822,In_2310);
or U4028 (N_4028,In_1537,In_1194);
and U4029 (N_4029,In_1293,In_1915);
and U4030 (N_4030,In_1035,In_2146);
and U4031 (N_4031,In_2214,In_2129);
nand U4032 (N_4032,In_1595,In_1765);
nand U4033 (N_4033,In_31,In_1722);
nor U4034 (N_4034,In_2347,In_2025);
nor U4035 (N_4035,In_1169,In_280);
nor U4036 (N_4036,In_1638,In_580);
and U4037 (N_4037,In_1344,In_1699);
and U4038 (N_4038,In_99,In_502);
or U4039 (N_4039,In_2400,In_1651);
or U4040 (N_4040,In_1849,In_2478);
and U4041 (N_4041,In_2023,In_1256);
nor U4042 (N_4042,In_797,In_1333);
and U4043 (N_4043,In_1832,In_1224);
or U4044 (N_4044,In_2042,In_984);
or U4045 (N_4045,In_1992,In_2221);
nor U4046 (N_4046,In_2235,In_2228);
nand U4047 (N_4047,In_2092,In_988);
and U4048 (N_4048,In_2288,In_1612);
and U4049 (N_4049,In_1339,In_244);
nor U4050 (N_4050,In_1808,In_1098);
or U4051 (N_4051,In_1689,In_484);
and U4052 (N_4052,In_2412,In_1773);
or U4053 (N_4053,In_1553,In_244);
or U4054 (N_4054,In_2248,In_27);
or U4055 (N_4055,In_1606,In_999);
or U4056 (N_4056,In_424,In_1363);
nand U4057 (N_4057,In_1930,In_2304);
nand U4058 (N_4058,In_640,In_1248);
nand U4059 (N_4059,In_1380,In_1863);
and U4060 (N_4060,In_2464,In_554);
or U4061 (N_4061,In_639,In_1394);
nor U4062 (N_4062,In_1004,In_121);
nand U4063 (N_4063,In_1735,In_207);
nor U4064 (N_4064,In_255,In_521);
nand U4065 (N_4065,In_172,In_1830);
nand U4066 (N_4066,In_1126,In_2321);
and U4067 (N_4067,In_353,In_2400);
nor U4068 (N_4068,In_2064,In_2243);
or U4069 (N_4069,In_2049,In_1060);
nand U4070 (N_4070,In_1170,In_801);
nand U4071 (N_4071,In_999,In_430);
nor U4072 (N_4072,In_1731,In_507);
or U4073 (N_4073,In_1523,In_39);
nand U4074 (N_4074,In_1096,In_324);
nand U4075 (N_4075,In_229,In_663);
nor U4076 (N_4076,In_2299,In_2243);
or U4077 (N_4077,In_655,In_875);
and U4078 (N_4078,In_2399,In_1100);
and U4079 (N_4079,In_99,In_2209);
nor U4080 (N_4080,In_2233,In_1655);
nor U4081 (N_4081,In_890,In_558);
nand U4082 (N_4082,In_342,In_1166);
and U4083 (N_4083,In_672,In_1950);
or U4084 (N_4084,In_1733,In_1805);
and U4085 (N_4085,In_1525,In_2278);
and U4086 (N_4086,In_1204,In_1706);
and U4087 (N_4087,In_424,In_1125);
or U4088 (N_4088,In_31,In_1005);
or U4089 (N_4089,In_1611,In_2033);
nor U4090 (N_4090,In_1276,In_10);
or U4091 (N_4091,In_109,In_767);
nand U4092 (N_4092,In_559,In_860);
or U4093 (N_4093,In_1650,In_2167);
nor U4094 (N_4094,In_304,In_2259);
xor U4095 (N_4095,In_2105,In_1225);
nand U4096 (N_4096,In_499,In_669);
or U4097 (N_4097,In_1571,In_2310);
or U4098 (N_4098,In_996,In_1775);
xnor U4099 (N_4099,In_2133,In_798);
nor U4100 (N_4100,In_1989,In_993);
nand U4101 (N_4101,In_1860,In_2254);
or U4102 (N_4102,In_170,In_660);
nand U4103 (N_4103,In_2129,In_1992);
xnor U4104 (N_4104,In_1567,In_1174);
nand U4105 (N_4105,In_246,In_1122);
nand U4106 (N_4106,In_1636,In_2301);
or U4107 (N_4107,In_75,In_2151);
or U4108 (N_4108,In_2089,In_703);
and U4109 (N_4109,In_847,In_1955);
or U4110 (N_4110,In_293,In_2131);
nand U4111 (N_4111,In_2062,In_1774);
or U4112 (N_4112,In_1307,In_508);
or U4113 (N_4113,In_1045,In_1312);
or U4114 (N_4114,In_896,In_1935);
and U4115 (N_4115,In_1445,In_717);
nand U4116 (N_4116,In_1780,In_1575);
and U4117 (N_4117,In_1924,In_120);
and U4118 (N_4118,In_1473,In_2424);
or U4119 (N_4119,In_27,In_606);
nand U4120 (N_4120,In_2126,In_1052);
nor U4121 (N_4121,In_706,In_952);
and U4122 (N_4122,In_2296,In_1954);
and U4123 (N_4123,In_454,In_787);
or U4124 (N_4124,In_709,In_152);
and U4125 (N_4125,In_2173,In_1319);
xor U4126 (N_4126,In_1015,In_607);
or U4127 (N_4127,In_2433,In_2312);
or U4128 (N_4128,In_588,In_2046);
or U4129 (N_4129,In_761,In_1167);
nand U4130 (N_4130,In_2203,In_330);
nand U4131 (N_4131,In_2262,In_1197);
nand U4132 (N_4132,In_1347,In_313);
nand U4133 (N_4133,In_637,In_2030);
nand U4134 (N_4134,In_685,In_2448);
or U4135 (N_4135,In_880,In_1752);
and U4136 (N_4136,In_1234,In_1762);
nand U4137 (N_4137,In_1766,In_2310);
or U4138 (N_4138,In_1229,In_2003);
xnor U4139 (N_4139,In_961,In_1314);
or U4140 (N_4140,In_1374,In_2104);
or U4141 (N_4141,In_925,In_1550);
nand U4142 (N_4142,In_274,In_110);
or U4143 (N_4143,In_309,In_1455);
nand U4144 (N_4144,In_2215,In_1485);
nand U4145 (N_4145,In_1841,In_711);
and U4146 (N_4146,In_1031,In_2089);
or U4147 (N_4147,In_1389,In_2343);
nand U4148 (N_4148,In_1025,In_89);
nor U4149 (N_4149,In_1727,In_1931);
or U4150 (N_4150,In_157,In_386);
xor U4151 (N_4151,In_1806,In_487);
and U4152 (N_4152,In_471,In_2407);
nor U4153 (N_4153,In_1250,In_912);
or U4154 (N_4154,In_571,In_1873);
nor U4155 (N_4155,In_1189,In_1888);
or U4156 (N_4156,In_1956,In_542);
or U4157 (N_4157,In_1414,In_144);
and U4158 (N_4158,In_232,In_780);
nor U4159 (N_4159,In_2233,In_2015);
or U4160 (N_4160,In_2414,In_470);
nor U4161 (N_4161,In_1050,In_1139);
or U4162 (N_4162,In_2409,In_1222);
and U4163 (N_4163,In_1512,In_731);
nor U4164 (N_4164,In_1264,In_1170);
nor U4165 (N_4165,In_2129,In_1232);
nand U4166 (N_4166,In_244,In_2269);
xnor U4167 (N_4167,In_1104,In_1154);
and U4168 (N_4168,In_2118,In_276);
or U4169 (N_4169,In_2368,In_2052);
nor U4170 (N_4170,In_16,In_2182);
nor U4171 (N_4171,In_1955,In_142);
or U4172 (N_4172,In_1421,In_2033);
nor U4173 (N_4173,In_1753,In_1607);
or U4174 (N_4174,In_2388,In_576);
nand U4175 (N_4175,In_2433,In_1941);
and U4176 (N_4176,In_1209,In_266);
and U4177 (N_4177,In_1675,In_531);
nor U4178 (N_4178,In_1563,In_508);
nor U4179 (N_4179,In_2028,In_1328);
and U4180 (N_4180,In_346,In_392);
nand U4181 (N_4181,In_644,In_140);
nand U4182 (N_4182,In_2097,In_1704);
nor U4183 (N_4183,In_1817,In_11);
or U4184 (N_4184,In_915,In_1426);
and U4185 (N_4185,In_722,In_331);
or U4186 (N_4186,In_1057,In_147);
or U4187 (N_4187,In_957,In_1509);
or U4188 (N_4188,In_1283,In_1412);
and U4189 (N_4189,In_373,In_815);
or U4190 (N_4190,In_417,In_56);
nor U4191 (N_4191,In_2166,In_1795);
nor U4192 (N_4192,In_207,In_265);
or U4193 (N_4193,In_598,In_348);
nor U4194 (N_4194,In_2186,In_588);
nand U4195 (N_4195,In_1143,In_1102);
and U4196 (N_4196,In_1542,In_1509);
nor U4197 (N_4197,In_2215,In_1048);
and U4198 (N_4198,In_2290,In_588);
and U4199 (N_4199,In_1610,In_2138);
xor U4200 (N_4200,In_1439,In_1209);
or U4201 (N_4201,In_415,In_1418);
or U4202 (N_4202,In_1421,In_1028);
nand U4203 (N_4203,In_316,In_548);
nor U4204 (N_4204,In_789,In_446);
nor U4205 (N_4205,In_1828,In_910);
nand U4206 (N_4206,In_314,In_607);
or U4207 (N_4207,In_412,In_1649);
and U4208 (N_4208,In_1336,In_919);
and U4209 (N_4209,In_371,In_1063);
nor U4210 (N_4210,In_1740,In_428);
nor U4211 (N_4211,In_1160,In_2135);
nand U4212 (N_4212,In_508,In_1705);
or U4213 (N_4213,In_367,In_160);
or U4214 (N_4214,In_1136,In_367);
nor U4215 (N_4215,In_1059,In_1122);
nand U4216 (N_4216,In_2159,In_2229);
and U4217 (N_4217,In_897,In_712);
or U4218 (N_4218,In_2450,In_1203);
and U4219 (N_4219,In_1209,In_407);
nand U4220 (N_4220,In_983,In_2419);
nor U4221 (N_4221,In_2255,In_795);
nand U4222 (N_4222,In_1549,In_2023);
or U4223 (N_4223,In_1662,In_976);
and U4224 (N_4224,In_1566,In_1612);
and U4225 (N_4225,In_1542,In_1547);
nor U4226 (N_4226,In_2187,In_2165);
nand U4227 (N_4227,In_2230,In_634);
nor U4228 (N_4228,In_1633,In_1862);
and U4229 (N_4229,In_2118,In_506);
and U4230 (N_4230,In_2209,In_1911);
nor U4231 (N_4231,In_1566,In_438);
and U4232 (N_4232,In_1743,In_473);
nor U4233 (N_4233,In_1535,In_1473);
or U4234 (N_4234,In_2445,In_775);
nor U4235 (N_4235,In_732,In_413);
nand U4236 (N_4236,In_100,In_1937);
nor U4237 (N_4237,In_1988,In_2490);
nand U4238 (N_4238,In_985,In_2003);
and U4239 (N_4239,In_2276,In_2424);
or U4240 (N_4240,In_614,In_1158);
nand U4241 (N_4241,In_709,In_333);
nand U4242 (N_4242,In_723,In_1325);
nand U4243 (N_4243,In_1404,In_1995);
nor U4244 (N_4244,In_1474,In_72);
or U4245 (N_4245,In_1020,In_2234);
nand U4246 (N_4246,In_2090,In_2062);
nand U4247 (N_4247,In_563,In_1318);
nor U4248 (N_4248,In_2385,In_664);
or U4249 (N_4249,In_1497,In_1453);
and U4250 (N_4250,In_1602,In_41);
nand U4251 (N_4251,In_2333,In_545);
or U4252 (N_4252,In_270,In_708);
nor U4253 (N_4253,In_981,In_1973);
nand U4254 (N_4254,In_1542,In_1883);
or U4255 (N_4255,In_2417,In_1327);
or U4256 (N_4256,In_1827,In_723);
and U4257 (N_4257,In_2372,In_158);
nand U4258 (N_4258,In_1561,In_773);
nor U4259 (N_4259,In_1651,In_5);
and U4260 (N_4260,In_159,In_1283);
nand U4261 (N_4261,In_2335,In_251);
nand U4262 (N_4262,In_140,In_1190);
or U4263 (N_4263,In_1356,In_80);
and U4264 (N_4264,In_2473,In_368);
nor U4265 (N_4265,In_1760,In_986);
and U4266 (N_4266,In_49,In_1195);
or U4267 (N_4267,In_1679,In_2292);
and U4268 (N_4268,In_1102,In_671);
nor U4269 (N_4269,In_1795,In_2388);
nand U4270 (N_4270,In_380,In_363);
or U4271 (N_4271,In_1863,In_185);
and U4272 (N_4272,In_1923,In_1338);
nor U4273 (N_4273,In_910,In_536);
nor U4274 (N_4274,In_1413,In_455);
or U4275 (N_4275,In_550,In_2431);
or U4276 (N_4276,In_843,In_22);
and U4277 (N_4277,In_391,In_1536);
or U4278 (N_4278,In_851,In_1598);
and U4279 (N_4279,In_1958,In_1726);
xor U4280 (N_4280,In_155,In_950);
nor U4281 (N_4281,In_1609,In_1944);
xnor U4282 (N_4282,In_519,In_2269);
or U4283 (N_4283,In_1949,In_1415);
or U4284 (N_4284,In_1777,In_1555);
nand U4285 (N_4285,In_2151,In_1013);
nand U4286 (N_4286,In_635,In_2116);
and U4287 (N_4287,In_1565,In_1250);
nor U4288 (N_4288,In_1847,In_2214);
nor U4289 (N_4289,In_756,In_2433);
or U4290 (N_4290,In_1584,In_1739);
nand U4291 (N_4291,In_1881,In_2317);
and U4292 (N_4292,In_1002,In_1762);
or U4293 (N_4293,In_1775,In_1779);
or U4294 (N_4294,In_724,In_816);
or U4295 (N_4295,In_1991,In_1740);
or U4296 (N_4296,In_1780,In_1302);
or U4297 (N_4297,In_313,In_1457);
and U4298 (N_4298,In_1716,In_798);
or U4299 (N_4299,In_1671,In_1689);
or U4300 (N_4300,In_2142,In_666);
nand U4301 (N_4301,In_1937,In_703);
or U4302 (N_4302,In_1844,In_2012);
or U4303 (N_4303,In_2247,In_1251);
nand U4304 (N_4304,In_1131,In_616);
nand U4305 (N_4305,In_504,In_2056);
and U4306 (N_4306,In_1914,In_1920);
and U4307 (N_4307,In_2423,In_322);
nor U4308 (N_4308,In_2361,In_2129);
and U4309 (N_4309,In_2233,In_1115);
nor U4310 (N_4310,In_1959,In_2064);
or U4311 (N_4311,In_18,In_2014);
or U4312 (N_4312,In_834,In_621);
nand U4313 (N_4313,In_686,In_1807);
or U4314 (N_4314,In_1072,In_1103);
and U4315 (N_4315,In_455,In_1053);
and U4316 (N_4316,In_1929,In_1213);
nor U4317 (N_4317,In_987,In_790);
nor U4318 (N_4318,In_245,In_1491);
nand U4319 (N_4319,In_1513,In_8);
nand U4320 (N_4320,In_350,In_891);
nor U4321 (N_4321,In_2398,In_79);
or U4322 (N_4322,In_1044,In_2142);
nor U4323 (N_4323,In_945,In_1864);
and U4324 (N_4324,In_1034,In_1831);
or U4325 (N_4325,In_1346,In_1523);
or U4326 (N_4326,In_57,In_814);
or U4327 (N_4327,In_1253,In_1171);
or U4328 (N_4328,In_1556,In_2092);
and U4329 (N_4329,In_1932,In_463);
nor U4330 (N_4330,In_1300,In_1417);
or U4331 (N_4331,In_1202,In_1870);
xnor U4332 (N_4332,In_1739,In_1347);
and U4333 (N_4333,In_1433,In_981);
nand U4334 (N_4334,In_441,In_1173);
nand U4335 (N_4335,In_771,In_2085);
and U4336 (N_4336,In_350,In_2399);
and U4337 (N_4337,In_329,In_2278);
or U4338 (N_4338,In_162,In_1760);
nand U4339 (N_4339,In_709,In_1019);
nor U4340 (N_4340,In_1832,In_306);
or U4341 (N_4341,In_1668,In_1866);
nand U4342 (N_4342,In_742,In_579);
or U4343 (N_4343,In_2092,In_2447);
nand U4344 (N_4344,In_2139,In_231);
nor U4345 (N_4345,In_462,In_1466);
and U4346 (N_4346,In_2364,In_1002);
and U4347 (N_4347,In_552,In_756);
nor U4348 (N_4348,In_1755,In_1670);
nor U4349 (N_4349,In_1638,In_2336);
nor U4350 (N_4350,In_1568,In_2199);
and U4351 (N_4351,In_504,In_169);
nand U4352 (N_4352,In_1929,In_1328);
or U4353 (N_4353,In_384,In_568);
nand U4354 (N_4354,In_1752,In_1053);
or U4355 (N_4355,In_2214,In_1581);
and U4356 (N_4356,In_2114,In_1351);
and U4357 (N_4357,In_74,In_433);
and U4358 (N_4358,In_1286,In_1718);
or U4359 (N_4359,In_1243,In_2462);
nand U4360 (N_4360,In_1948,In_598);
nor U4361 (N_4361,In_118,In_42);
or U4362 (N_4362,In_2284,In_1519);
nor U4363 (N_4363,In_363,In_449);
nand U4364 (N_4364,In_241,In_1770);
nand U4365 (N_4365,In_1611,In_1690);
nor U4366 (N_4366,In_1171,In_1602);
nand U4367 (N_4367,In_198,In_203);
nor U4368 (N_4368,In_211,In_1310);
and U4369 (N_4369,In_1543,In_1513);
nand U4370 (N_4370,In_701,In_625);
or U4371 (N_4371,In_764,In_226);
nand U4372 (N_4372,In_692,In_277);
or U4373 (N_4373,In_1653,In_886);
or U4374 (N_4374,In_665,In_2198);
nand U4375 (N_4375,In_1973,In_1321);
or U4376 (N_4376,In_2201,In_298);
nand U4377 (N_4377,In_255,In_2338);
xnor U4378 (N_4378,In_1355,In_2420);
or U4379 (N_4379,In_1339,In_2007);
nand U4380 (N_4380,In_555,In_2256);
nor U4381 (N_4381,In_406,In_1595);
and U4382 (N_4382,In_617,In_572);
and U4383 (N_4383,In_4,In_1976);
or U4384 (N_4384,In_298,In_1247);
or U4385 (N_4385,In_2320,In_475);
or U4386 (N_4386,In_1357,In_570);
nor U4387 (N_4387,In_988,In_746);
nand U4388 (N_4388,In_1529,In_2196);
and U4389 (N_4389,In_2243,In_1692);
nand U4390 (N_4390,In_2085,In_60);
and U4391 (N_4391,In_239,In_454);
nor U4392 (N_4392,In_1948,In_1478);
nor U4393 (N_4393,In_1556,In_323);
and U4394 (N_4394,In_769,In_1640);
nand U4395 (N_4395,In_311,In_1877);
nand U4396 (N_4396,In_1524,In_813);
or U4397 (N_4397,In_2499,In_2249);
nand U4398 (N_4398,In_1467,In_1274);
nor U4399 (N_4399,In_150,In_1368);
and U4400 (N_4400,In_2401,In_642);
and U4401 (N_4401,In_95,In_1877);
nand U4402 (N_4402,In_1157,In_650);
nand U4403 (N_4403,In_329,In_2183);
nor U4404 (N_4404,In_1727,In_977);
or U4405 (N_4405,In_1614,In_700);
and U4406 (N_4406,In_490,In_1805);
nor U4407 (N_4407,In_1302,In_2300);
nand U4408 (N_4408,In_860,In_92);
nor U4409 (N_4409,In_1562,In_134);
or U4410 (N_4410,In_264,In_1201);
nor U4411 (N_4411,In_150,In_366);
or U4412 (N_4412,In_563,In_321);
or U4413 (N_4413,In_1503,In_188);
nand U4414 (N_4414,In_1554,In_1047);
nor U4415 (N_4415,In_1557,In_777);
and U4416 (N_4416,In_1132,In_1746);
nand U4417 (N_4417,In_2475,In_2352);
nor U4418 (N_4418,In_889,In_1836);
or U4419 (N_4419,In_876,In_1932);
and U4420 (N_4420,In_1582,In_263);
nand U4421 (N_4421,In_721,In_1601);
nor U4422 (N_4422,In_864,In_503);
and U4423 (N_4423,In_49,In_961);
or U4424 (N_4424,In_380,In_947);
xnor U4425 (N_4425,In_1661,In_818);
and U4426 (N_4426,In_2009,In_1593);
and U4427 (N_4427,In_1138,In_624);
nand U4428 (N_4428,In_2430,In_2128);
and U4429 (N_4429,In_702,In_1119);
and U4430 (N_4430,In_1226,In_1707);
or U4431 (N_4431,In_1022,In_1853);
nand U4432 (N_4432,In_1617,In_2005);
nand U4433 (N_4433,In_59,In_82);
nand U4434 (N_4434,In_2181,In_611);
or U4435 (N_4435,In_2430,In_1410);
or U4436 (N_4436,In_2364,In_2313);
nand U4437 (N_4437,In_948,In_1505);
or U4438 (N_4438,In_2451,In_1413);
nand U4439 (N_4439,In_2481,In_803);
or U4440 (N_4440,In_468,In_2024);
nand U4441 (N_4441,In_1659,In_1611);
and U4442 (N_4442,In_667,In_891);
and U4443 (N_4443,In_274,In_1502);
and U4444 (N_4444,In_442,In_1509);
nand U4445 (N_4445,In_1849,In_1211);
nand U4446 (N_4446,In_1960,In_187);
xnor U4447 (N_4447,In_1434,In_2198);
or U4448 (N_4448,In_1033,In_366);
nand U4449 (N_4449,In_880,In_432);
and U4450 (N_4450,In_488,In_757);
or U4451 (N_4451,In_269,In_1183);
or U4452 (N_4452,In_1421,In_213);
nand U4453 (N_4453,In_51,In_360);
or U4454 (N_4454,In_294,In_2102);
and U4455 (N_4455,In_429,In_982);
or U4456 (N_4456,In_419,In_380);
or U4457 (N_4457,In_1887,In_1506);
or U4458 (N_4458,In_2067,In_2358);
and U4459 (N_4459,In_1997,In_1480);
and U4460 (N_4460,In_2483,In_808);
and U4461 (N_4461,In_1307,In_1449);
and U4462 (N_4462,In_439,In_1837);
or U4463 (N_4463,In_2040,In_1576);
nand U4464 (N_4464,In_561,In_1804);
nor U4465 (N_4465,In_2405,In_1562);
and U4466 (N_4466,In_292,In_1326);
or U4467 (N_4467,In_1523,In_1314);
nor U4468 (N_4468,In_586,In_18);
and U4469 (N_4469,In_2161,In_2414);
and U4470 (N_4470,In_2367,In_596);
and U4471 (N_4471,In_5,In_1815);
and U4472 (N_4472,In_1967,In_790);
or U4473 (N_4473,In_922,In_132);
or U4474 (N_4474,In_1284,In_1657);
and U4475 (N_4475,In_293,In_455);
or U4476 (N_4476,In_1657,In_286);
nand U4477 (N_4477,In_1973,In_625);
nand U4478 (N_4478,In_1276,In_1466);
nand U4479 (N_4479,In_1953,In_1043);
and U4480 (N_4480,In_184,In_2);
and U4481 (N_4481,In_139,In_1979);
nor U4482 (N_4482,In_582,In_1459);
nor U4483 (N_4483,In_1350,In_992);
nand U4484 (N_4484,In_493,In_930);
nand U4485 (N_4485,In_1534,In_2412);
nand U4486 (N_4486,In_1257,In_1175);
nor U4487 (N_4487,In_1771,In_1289);
nor U4488 (N_4488,In_868,In_1801);
and U4489 (N_4489,In_2154,In_1604);
and U4490 (N_4490,In_1824,In_2327);
nor U4491 (N_4491,In_644,In_2399);
nor U4492 (N_4492,In_429,In_565);
and U4493 (N_4493,In_1587,In_2313);
or U4494 (N_4494,In_2240,In_1485);
and U4495 (N_4495,In_273,In_2338);
and U4496 (N_4496,In_1605,In_26);
or U4497 (N_4497,In_1911,In_2194);
and U4498 (N_4498,In_974,In_428);
nor U4499 (N_4499,In_1597,In_2451);
xor U4500 (N_4500,In_366,In_109);
nand U4501 (N_4501,In_286,In_1234);
nor U4502 (N_4502,In_2008,In_930);
or U4503 (N_4503,In_2336,In_795);
nand U4504 (N_4504,In_245,In_109);
nor U4505 (N_4505,In_326,In_249);
nand U4506 (N_4506,In_1744,In_1759);
nor U4507 (N_4507,In_2226,In_166);
nand U4508 (N_4508,In_434,In_577);
nand U4509 (N_4509,In_185,In_1626);
or U4510 (N_4510,In_2183,In_981);
nor U4511 (N_4511,In_726,In_175);
nand U4512 (N_4512,In_2190,In_577);
nor U4513 (N_4513,In_2250,In_768);
nand U4514 (N_4514,In_2310,In_336);
nand U4515 (N_4515,In_1112,In_1664);
nor U4516 (N_4516,In_1062,In_368);
and U4517 (N_4517,In_1595,In_1962);
or U4518 (N_4518,In_259,In_357);
and U4519 (N_4519,In_2499,In_1819);
or U4520 (N_4520,In_479,In_392);
nand U4521 (N_4521,In_829,In_473);
and U4522 (N_4522,In_1104,In_1308);
nor U4523 (N_4523,In_423,In_1421);
nand U4524 (N_4524,In_1136,In_349);
and U4525 (N_4525,In_868,In_66);
nor U4526 (N_4526,In_1190,In_1116);
and U4527 (N_4527,In_395,In_277);
or U4528 (N_4528,In_401,In_1069);
nor U4529 (N_4529,In_1771,In_486);
or U4530 (N_4530,In_1661,In_846);
and U4531 (N_4531,In_717,In_1346);
nand U4532 (N_4532,In_582,In_1428);
and U4533 (N_4533,In_1835,In_2404);
nand U4534 (N_4534,In_467,In_641);
nand U4535 (N_4535,In_561,In_273);
nand U4536 (N_4536,In_1413,In_969);
nor U4537 (N_4537,In_2300,In_102);
nor U4538 (N_4538,In_807,In_14);
nor U4539 (N_4539,In_24,In_576);
nor U4540 (N_4540,In_2286,In_1038);
nor U4541 (N_4541,In_95,In_817);
nor U4542 (N_4542,In_2457,In_792);
nand U4543 (N_4543,In_581,In_1051);
nor U4544 (N_4544,In_855,In_1161);
nand U4545 (N_4545,In_2019,In_1764);
nor U4546 (N_4546,In_1605,In_233);
and U4547 (N_4547,In_779,In_739);
nand U4548 (N_4548,In_1665,In_1803);
and U4549 (N_4549,In_1353,In_607);
or U4550 (N_4550,In_1219,In_1849);
nor U4551 (N_4551,In_2255,In_1457);
or U4552 (N_4552,In_1145,In_479);
nor U4553 (N_4553,In_591,In_1020);
nor U4554 (N_4554,In_1376,In_1094);
or U4555 (N_4555,In_460,In_349);
nand U4556 (N_4556,In_2330,In_498);
and U4557 (N_4557,In_1949,In_2299);
nor U4558 (N_4558,In_884,In_2447);
or U4559 (N_4559,In_2469,In_1913);
and U4560 (N_4560,In_1781,In_2110);
nand U4561 (N_4561,In_2224,In_1313);
or U4562 (N_4562,In_2052,In_567);
nor U4563 (N_4563,In_1048,In_1927);
nor U4564 (N_4564,In_635,In_52);
nor U4565 (N_4565,In_846,In_1070);
and U4566 (N_4566,In_903,In_123);
or U4567 (N_4567,In_815,In_1316);
nand U4568 (N_4568,In_129,In_790);
and U4569 (N_4569,In_2304,In_147);
nand U4570 (N_4570,In_509,In_662);
and U4571 (N_4571,In_2357,In_1032);
nor U4572 (N_4572,In_161,In_2387);
xor U4573 (N_4573,In_689,In_2487);
nor U4574 (N_4574,In_245,In_696);
nor U4575 (N_4575,In_1788,In_1300);
and U4576 (N_4576,In_118,In_1194);
xor U4577 (N_4577,In_2114,In_1490);
nand U4578 (N_4578,In_1553,In_926);
nand U4579 (N_4579,In_2256,In_905);
or U4580 (N_4580,In_429,In_1440);
nor U4581 (N_4581,In_1018,In_536);
nand U4582 (N_4582,In_705,In_175);
and U4583 (N_4583,In_504,In_2322);
and U4584 (N_4584,In_883,In_1904);
nor U4585 (N_4585,In_1677,In_1038);
nor U4586 (N_4586,In_1892,In_193);
nand U4587 (N_4587,In_923,In_2037);
nand U4588 (N_4588,In_838,In_536);
or U4589 (N_4589,In_634,In_2050);
nand U4590 (N_4590,In_1357,In_2346);
and U4591 (N_4591,In_1590,In_177);
and U4592 (N_4592,In_1746,In_1119);
and U4593 (N_4593,In_1776,In_382);
and U4594 (N_4594,In_320,In_1815);
and U4595 (N_4595,In_292,In_827);
or U4596 (N_4596,In_718,In_1733);
and U4597 (N_4597,In_1659,In_991);
and U4598 (N_4598,In_379,In_2239);
nor U4599 (N_4599,In_2004,In_1009);
or U4600 (N_4600,In_60,In_2375);
and U4601 (N_4601,In_1804,In_2439);
nor U4602 (N_4602,In_526,In_2428);
nor U4603 (N_4603,In_1035,In_2188);
nor U4604 (N_4604,In_1794,In_1635);
nor U4605 (N_4605,In_1008,In_1515);
and U4606 (N_4606,In_2352,In_445);
nor U4607 (N_4607,In_2183,In_1810);
and U4608 (N_4608,In_674,In_2155);
xor U4609 (N_4609,In_832,In_689);
or U4610 (N_4610,In_2374,In_1553);
nor U4611 (N_4611,In_1972,In_1680);
and U4612 (N_4612,In_1496,In_2024);
and U4613 (N_4613,In_497,In_107);
nand U4614 (N_4614,In_424,In_177);
and U4615 (N_4615,In_227,In_1527);
or U4616 (N_4616,In_1728,In_949);
and U4617 (N_4617,In_1725,In_2469);
xor U4618 (N_4618,In_1132,In_176);
nand U4619 (N_4619,In_1142,In_1326);
or U4620 (N_4620,In_2440,In_2266);
and U4621 (N_4621,In_2006,In_2449);
nor U4622 (N_4622,In_223,In_703);
nor U4623 (N_4623,In_1083,In_1122);
nor U4624 (N_4624,In_433,In_164);
nand U4625 (N_4625,In_2286,In_2411);
nor U4626 (N_4626,In_744,In_1103);
nand U4627 (N_4627,In_768,In_453);
or U4628 (N_4628,In_2347,In_382);
nand U4629 (N_4629,In_2188,In_1607);
or U4630 (N_4630,In_1186,In_1471);
or U4631 (N_4631,In_1256,In_1166);
and U4632 (N_4632,In_875,In_2495);
nand U4633 (N_4633,In_1742,In_1732);
nand U4634 (N_4634,In_515,In_218);
nand U4635 (N_4635,In_2331,In_2081);
or U4636 (N_4636,In_92,In_276);
and U4637 (N_4637,In_2415,In_1384);
nor U4638 (N_4638,In_1244,In_2007);
or U4639 (N_4639,In_479,In_1636);
or U4640 (N_4640,In_1783,In_605);
or U4641 (N_4641,In_522,In_258);
nor U4642 (N_4642,In_221,In_1329);
nand U4643 (N_4643,In_843,In_444);
and U4644 (N_4644,In_2347,In_1164);
nor U4645 (N_4645,In_83,In_680);
and U4646 (N_4646,In_1336,In_2050);
nor U4647 (N_4647,In_111,In_2129);
and U4648 (N_4648,In_2423,In_2096);
nor U4649 (N_4649,In_1935,In_1541);
nor U4650 (N_4650,In_2205,In_775);
and U4651 (N_4651,In_1913,In_1281);
or U4652 (N_4652,In_1469,In_1739);
or U4653 (N_4653,In_811,In_2086);
nand U4654 (N_4654,In_771,In_1414);
xor U4655 (N_4655,In_1279,In_108);
nor U4656 (N_4656,In_1847,In_1841);
and U4657 (N_4657,In_2314,In_569);
nand U4658 (N_4658,In_248,In_1965);
nand U4659 (N_4659,In_2120,In_2113);
and U4660 (N_4660,In_1196,In_368);
or U4661 (N_4661,In_998,In_1966);
or U4662 (N_4662,In_1009,In_380);
or U4663 (N_4663,In_1864,In_1402);
nor U4664 (N_4664,In_1828,In_1528);
and U4665 (N_4665,In_794,In_1568);
nand U4666 (N_4666,In_551,In_270);
nand U4667 (N_4667,In_432,In_1142);
nor U4668 (N_4668,In_362,In_1733);
or U4669 (N_4669,In_797,In_1314);
or U4670 (N_4670,In_1158,In_735);
nor U4671 (N_4671,In_876,In_737);
nor U4672 (N_4672,In_2092,In_683);
nand U4673 (N_4673,In_1772,In_2161);
nor U4674 (N_4674,In_1881,In_2287);
nand U4675 (N_4675,In_1726,In_159);
nor U4676 (N_4676,In_1261,In_2167);
nand U4677 (N_4677,In_1844,In_1823);
or U4678 (N_4678,In_565,In_2124);
nor U4679 (N_4679,In_207,In_378);
or U4680 (N_4680,In_294,In_1741);
or U4681 (N_4681,In_1202,In_1635);
nand U4682 (N_4682,In_347,In_1979);
nand U4683 (N_4683,In_2047,In_149);
and U4684 (N_4684,In_667,In_868);
nand U4685 (N_4685,In_964,In_1576);
or U4686 (N_4686,In_807,In_2130);
nand U4687 (N_4687,In_426,In_1901);
and U4688 (N_4688,In_1612,In_2402);
nor U4689 (N_4689,In_809,In_2202);
nor U4690 (N_4690,In_810,In_381);
and U4691 (N_4691,In_823,In_1469);
nand U4692 (N_4692,In_516,In_2207);
and U4693 (N_4693,In_1671,In_2371);
or U4694 (N_4694,In_2161,In_1423);
or U4695 (N_4695,In_909,In_1508);
and U4696 (N_4696,In_647,In_2282);
or U4697 (N_4697,In_702,In_1529);
nor U4698 (N_4698,In_2308,In_1530);
or U4699 (N_4699,In_1714,In_1873);
and U4700 (N_4700,In_1767,In_2432);
or U4701 (N_4701,In_1106,In_179);
or U4702 (N_4702,In_1167,In_28);
or U4703 (N_4703,In_2409,In_30);
and U4704 (N_4704,In_74,In_675);
or U4705 (N_4705,In_179,In_2186);
xnor U4706 (N_4706,In_909,In_1078);
and U4707 (N_4707,In_951,In_841);
or U4708 (N_4708,In_1606,In_1635);
nand U4709 (N_4709,In_2253,In_2381);
or U4710 (N_4710,In_2484,In_1862);
nand U4711 (N_4711,In_2440,In_1464);
nor U4712 (N_4712,In_1891,In_626);
nand U4713 (N_4713,In_1018,In_1058);
nor U4714 (N_4714,In_874,In_1822);
or U4715 (N_4715,In_1066,In_1850);
and U4716 (N_4716,In_2279,In_2034);
and U4717 (N_4717,In_1058,In_135);
nand U4718 (N_4718,In_350,In_1522);
or U4719 (N_4719,In_1116,In_513);
and U4720 (N_4720,In_1706,In_1935);
or U4721 (N_4721,In_1082,In_782);
nand U4722 (N_4722,In_346,In_1652);
or U4723 (N_4723,In_923,In_1105);
nor U4724 (N_4724,In_230,In_705);
and U4725 (N_4725,In_662,In_1421);
and U4726 (N_4726,In_336,In_241);
nand U4727 (N_4727,In_613,In_2059);
nand U4728 (N_4728,In_2230,In_2399);
and U4729 (N_4729,In_37,In_785);
nand U4730 (N_4730,In_1788,In_442);
or U4731 (N_4731,In_2081,In_1635);
or U4732 (N_4732,In_2320,In_2091);
nor U4733 (N_4733,In_945,In_986);
nor U4734 (N_4734,In_540,In_377);
or U4735 (N_4735,In_1409,In_120);
or U4736 (N_4736,In_1008,In_416);
or U4737 (N_4737,In_774,In_1697);
or U4738 (N_4738,In_1699,In_780);
or U4739 (N_4739,In_791,In_474);
nand U4740 (N_4740,In_114,In_2404);
and U4741 (N_4741,In_985,In_1396);
nor U4742 (N_4742,In_2012,In_298);
or U4743 (N_4743,In_298,In_1534);
nand U4744 (N_4744,In_1834,In_1552);
or U4745 (N_4745,In_2459,In_1361);
nand U4746 (N_4746,In_1149,In_508);
xnor U4747 (N_4747,In_820,In_1905);
or U4748 (N_4748,In_205,In_2100);
and U4749 (N_4749,In_2371,In_674);
or U4750 (N_4750,In_958,In_926);
and U4751 (N_4751,In_2466,In_1822);
and U4752 (N_4752,In_695,In_1841);
and U4753 (N_4753,In_578,In_651);
or U4754 (N_4754,In_1437,In_2152);
nor U4755 (N_4755,In_1633,In_1364);
or U4756 (N_4756,In_1028,In_263);
or U4757 (N_4757,In_1893,In_1872);
nand U4758 (N_4758,In_12,In_225);
nand U4759 (N_4759,In_2391,In_2307);
and U4760 (N_4760,In_2225,In_2038);
nor U4761 (N_4761,In_1947,In_372);
and U4762 (N_4762,In_1370,In_726);
or U4763 (N_4763,In_2169,In_536);
nand U4764 (N_4764,In_2248,In_835);
nand U4765 (N_4765,In_2076,In_778);
or U4766 (N_4766,In_2367,In_410);
or U4767 (N_4767,In_708,In_2453);
xor U4768 (N_4768,In_605,In_833);
and U4769 (N_4769,In_186,In_573);
and U4770 (N_4770,In_140,In_1941);
or U4771 (N_4771,In_463,In_1039);
nand U4772 (N_4772,In_798,In_362);
nand U4773 (N_4773,In_1543,In_1797);
and U4774 (N_4774,In_1194,In_1371);
nor U4775 (N_4775,In_529,In_1594);
nor U4776 (N_4776,In_1258,In_426);
nand U4777 (N_4777,In_1173,In_450);
or U4778 (N_4778,In_42,In_127);
or U4779 (N_4779,In_609,In_2350);
and U4780 (N_4780,In_2473,In_1654);
or U4781 (N_4781,In_2388,In_1705);
and U4782 (N_4782,In_1927,In_1650);
nand U4783 (N_4783,In_1151,In_1637);
nor U4784 (N_4784,In_522,In_1558);
nand U4785 (N_4785,In_1078,In_98);
nand U4786 (N_4786,In_2000,In_775);
nand U4787 (N_4787,In_1889,In_593);
nor U4788 (N_4788,In_339,In_1301);
or U4789 (N_4789,In_1983,In_2376);
nor U4790 (N_4790,In_541,In_820);
or U4791 (N_4791,In_445,In_1995);
nor U4792 (N_4792,In_2474,In_1247);
or U4793 (N_4793,In_2287,In_2262);
nor U4794 (N_4794,In_888,In_82);
nand U4795 (N_4795,In_1185,In_1678);
nand U4796 (N_4796,In_24,In_40);
nor U4797 (N_4797,In_857,In_768);
or U4798 (N_4798,In_1152,In_734);
nor U4799 (N_4799,In_785,In_1716);
or U4800 (N_4800,In_1989,In_2021);
and U4801 (N_4801,In_810,In_213);
or U4802 (N_4802,In_2030,In_427);
nor U4803 (N_4803,In_2489,In_2304);
or U4804 (N_4804,In_2001,In_170);
nand U4805 (N_4805,In_1011,In_1200);
nand U4806 (N_4806,In_1656,In_2444);
and U4807 (N_4807,In_856,In_751);
and U4808 (N_4808,In_1698,In_1650);
or U4809 (N_4809,In_2282,In_838);
and U4810 (N_4810,In_1057,In_1305);
and U4811 (N_4811,In_383,In_371);
or U4812 (N_4812,In_360,In_2034);
nor U4813 (N_4813,In_939,In_1081);
nor U4814 (N_4814,In_57,In_2233);
nand U4815 (N_4815,In_716,In_241);
nand U4816 (N_4816,In_2188,In_35);
xor U4817 (N_4817,In_1523,In_465);
and U4818 (N_4818,In_2480,In_1953);
or U4819 (N_4819,In_1684,In_2040);
xnor U4820 (N_4820,In_2175,In_877);
nand U4821 (N_4821,In_194,In_1100);
nand U4822 (N_4822,In_2106,In_2085);
and U4823 (N_4823,In_1900,In_782);
nor U4824 (N_4824,In_2090,In_2164);
nand U4825 (N_4825,In_850,In_92);
and U4826 (N_4826,In_1517,In_271);
or U4827 (N_4827,In_137,In_1337);
nor U4828 (N_4828,In_2247,In_1939);
xnor U4829 (N_4829,In_662,In_1439);
and U4830 (N_4830,In_2168,In_390);
or U4831 (N_4831,In_1148,In_1981);
and U4832 (N_4832,In_1078,In_424);
nor U4833 (N_4833,In_424,In_1036);
nor U4834 (N_4834,In_1542,In_1197);
nand U4835 (N_4835,In_1992,In_561);
nand U4836 (N_4836,In_430,In_1366);
nand U4837 (N_4837,In_199,In_1711);
nand U4838 (N_4838,In_265,In_1031);
or U4839 (N_4839,In_2327,In_429);
nor U4840 (N_4840,In_330,In_904);
nor U4841 (N_4841,In_629,In_532);
nand U4842 (N_4842,In_168,In_666);
or U4843 (N_4843,In_184,In_1641);
nand U4844 (N_4844,In_407,In_1849);
nand U4845 (N_4845,In_1165,In_1937);
or U4846 (N_4846,In_1213,In_1813);
nor U4847 (N_4847,In_438,In_2131);
or U4848 (N_4848,In_1895,In_1868);
nand U4849 (N_4849,In_189,In_86);
nand U4850 (N_4850,In_1330,In_755);
and U4851 (N_4851,In_467,In_938);
and U4852 (N_4852,In_1006,In_2045);
nand U4853 (N_4853,In_831,In_972);
nand U4854 (N_4854,In_2460,In_626);
nand U4855 (N_4855,In_1633,In_2244);
nand U4856 (N_4856,In_1016,In_104);
nor U4857 (N_4857,In_525,In_370);
and U4858 (N_4858,In_2236,In_1364);
nor U4859 (N_4859,In_1976,In_1970);
nand U4860 (N_4860,In_164,In_686);
nand U4861 (N_4861,In_208,In_904);
or U4862 (N_4862,In_1667,In_972);
nor U4863 (N_4863,In_91,In_642);
nand U4864 (N_4864,In_2224,In_1929);
or U4865 (N_4865,In_1640,In_2052);
nand U4866 (N_4866,In_1276,In_1876);
nand U4867 (N_4867,In_807,In_916);
nor U4868 (N_4868,In_550,In_1568);
nand U4869 (N_4869,In_2435,In_2278);
and U4870 (N_4870,In_1832,In_1804);
nand U4871 (N_4871,In_2244,In_982);
and U4872 (N_4872,In_962,In_80);
and U4873 (N_4873,In_1164,In_812);
or U4874 (N_4874,In_611,In_57);
xor U4875 (N_4875,In_120,In_2116);
nand U4876 (N_4876,In_1232,In_376);
and U4877 (N_4877,In_1493,In_934);
nand U4878 (N_4878,In_1851,In_1864);
nor U4879 (N_4879,In_2081,In_1159);
and U4880 (N_4880,In_1559,In_2237);
nand U4881 (N_4881,In_761,In_1209);
and U4882 (N_4882,In_81,In_732);
nor U4883 (N_4883,In_2060,In_205);
or U4884 (N_4884,In_1904,In_473);
nor U4885 (N_4885,In_1121,In_1601);
nand U4886 (N_4886,In_2056,In_1701);
nor U4887 (N_4887,In_925,In_135);
or U4888 (N_4888,In_454,In_1380);
nor U4889 (N_4889,In_1296,In_666);
or U4890 (N_4890,In_2482,In_222);
and U4891 (N_4891,In_880,In_507);
nand U4892 (N_4892,In_356,In_515);
and U4893 (N_4893,In_1531,In_614);
xor U4894 (N_4894,In_695,In_2257);
or U4895 (N_4895,In_1088,In_93);
nor U4896 (N_4896,In_2404,In_1591);
nand U4897 (N_4897,In_907,In_2460);
nand U4898 (N_4898,In_2466,In_132);
nand U4899 (N_4899,In_597,In_21);
and U4900 (N_4900,In_2498,In_493);
nor U4901 (N_4901,In_1795,In_1371);
nor U4902 (N_4902,In_28,In_2471);
or U4903 (N_4903,In_2368,In_1243);
nand U4904 (N_4904,In_2422,In_1083);
and U4905 (N_4905,In_1287,In_831);
or U4906 (N_4906,In_92,In_1055);
or U4907 (N_4907,In_1261,In_638);
nand U4908 (N_4908,In_2092,In_817);
xnor U4909 (N_4909,In_1396,In_2246);
nor U4910 (N_4910,In_892,In_1669);
and U4911 (N_4911,In_1327,In_1077);
nand U4912 (N_4912,In_1621,In_1900);
nor U4913 (N_4913,In_2245,In_1225);
nor U4914 (N_4914,In_2394,In_2175);
nor U4915 (N_4915,In_206,In_1732);
nand U4916 (N_4916,In_225,In_380);
nand U4917 (N_4917,In_2285,In_1136);
and U4918 (N_4918,In_926,In_1443);
and U4919 (N_4919,In_629,In_116);
or U4920 (N_4920,In_527,In_2418);
or U4921 (N_4921,In_15,In_1265);
xor U4922 (N_4922,In_2274,In_332);
and U4923 (N_4923,In_2101,In_2015);
and U4924 (N_4924,In_404,In_1814);
and U4925 (N_4925,In_1233,In_50);
nor U4926 (N_4926,In_1136,In_1173);
nand U4927 (N_4927,In_1697,In_207);
nand U4928 (N_4928,In_969,In_157);
or U4929 (N_4929,In_1977,In_481);
or U4930 (N_4930,In_840,In_382);
or U4931 (N_4931,In_1658,In_856);
nand U4932 (N_4932,In_469,In_781);
or U4933 (N_4933,In_87,In_1304);
or U4934 (N_4934,In_692,In_1557);
nand U4935 (N_4935,In_288,In_2361);
nor U4936 (N_4936,In_2190,In_1393);
nor U4937 (N_4937,In_1900,In_1415);
nor U4938 (N_4938,In_505,In_1872);
and U4939 (N_4939,In_334,In_1782);
nor U4940 (N_4940,In_2190,In_2068);
nor U4941 (N_4941,In_1325,In_260);
or U4942 (N_4942,In_789,In_1553);
nand U4943 (N_4943,In_742,In_1046);
nand U4944 (N_4944,In_1076,In_1423);
or U4945 (N_4945,In_1663,In_722);
nor U4946 (N_4946,In_803,In_1073);
or U4947 (N_4947,In_2032,In_644);
and U4948 (N_4948,In_254,In_1454);
or U4949 (N_4949,In_1898,In_1744);
nor U4950 (N_4950,In_743,In_2115);
nor U4951 (N_4951,In_2009,In_772);
or U4952 (N_4952,In_1860,In_2095);
and U4953 (N_4953,In_1306,In_2421);
or U4954 (N_4954,In_898,In_349);
and U4955 (N_4955,In_1826,In_1316);
nand U4956 (N_4956,In_690,In_2059);
nor U4957 (N_4957,In_404,In_1358);
nand U4958 (N_4958,In_386,In_1022);
or U4959 (N_4959,In_223,In_1975);
or U4960 (N_4960,In_1188,In_2329);
nor U4961 (N_4961,In_1349,In_1468);
nor U4962 (N_4962,In_2094,In_578);
and U4963 (N_4963,In_2177,In_448);
nand U4964 (N_4964,In_2232,In_1094);
nand U4965 (N_4965,In_1526,In_1);
and U4966 (N_4966,In_193,In_1890);
or U4967 (N_4967,In_1800,In_711);
nor U4968 (N_4968,In_765,In_2409);
and U4969 (N_4969,In_1100,In_1070);
nor U4970 (N_4970,In_781,In_2066);
or U4971 (N_4971,In_1734,In_423);
nand U4972 (N_4972,In_2247,In_1117);
nor U4973 (N_4973,In_2029,In_1850);
and U4974 (N_4974,In_1376,In_1795);
or U4975 (N_4975,In_1547,In_1945);
nor U4976 (N_4976,In_1598,In_1148);
nor U4977 (N_4977,In_1501,In_1832);
nor U4978 (N_4978,In_725,In_235);
or U4979 (N_4979,In_906,In_804);
and U4980 (N_4980,In_1852,In_702);
and U4981 (N_4981,In_1504,In_613);
nor U4982 (N_4982,In_525,In_2148);
or U4983 (N_4983,In_2371,In_1421);
and U4984 (N_4984,In_2166,In_1344);
and U4985 (N_4985,In_1716,In_1628);
nand U4986 (N_4986,In_1173,In_2090);
and U4987 (N_4987,In_847,In_1261);
or U4988 (N_4988,In_840,In_497);
and U4989 (N_4989,In_661,In_449);
or U4990 (N_4990,In_180,In_1945);
nor U4991 (N_4991,In_995,In_2409);
or U4992 (N_4992,In_2460,In_756);
nand U4993 (N_4993,In_2323,In_475);
nand U4994 (N_4994,In_2333,In_32);
nor U4995 (N_4995,In_950,In_173);
and U4996 (N_4996,In_1592,In_958);
or U4997 (N_4997,In_290,In_185);
and U4998 (N_4998,In_2004,In_1551);
and U4999 (N_4999,In_2024,In_2258);
and U5000 (N_5000,In_1235,In_1049);
and U5001 (N_5001,In_793,In_594);
or U5002 (N_5002,In_994,In_2264);
nor U5003 (N_5003,In_2387,In_1039);
nand U5004 (N_5004,In_2350,In_1598);
nor U5005 (N_5005,In_1921,In_1739);
nor U5006 (N_5006,In_490,In_2032);
and U5007 (N_5007,In_134,In_180);
nor U5008 (N_5008,In_2299,In_1092);
or U5009 (N_5009,In_1934,In_2250);
xnor U5010 (N_5010,In_605,In_1932);
or U5011 (N_5011,In_54,In_1123);
nor U5012 (N_5012,In_1738,In_909);
nand U5013 (N_5013,In_229,In_774);
or U5014 (N_5014,In_1016,In_743);
and U5015 (N_5015,In_1406,In_2404);
and U5016 (N_5016,In_2345,In_1247);
nor U5017 (N_5017,In_2322,In_167);
nor U5018 (N_5018,In_1318,In_653);
nor U5019 (N_5019,In_515,In_1139);
nor U5020 (N_5020,In_585,In_1936);
or U5021 (N_5021,In_1932,In_2145);
or U5022 (N_5022,In_666,In_2187);
nand U5023 (N_5023,In_2410,In_1898);
and U5024 (N_5024,In_571,In_1431);
nand U5025 (N_5025,In_162,In_1429);
and U5026 (N_5026,In_46,In_51);
xnor U5027 (N_5027,In_681,In_690);
nor U5028 (N_5028,In_1253,In_2387);
nor U5029 (N_5029,In_1915,In_1514);
nand U5030 (N_5030,In_1223,In_2238);
or U5031 (N_5031,In_206,In_1002);
nand U5032 (N_5032,In_652,In_741);
nand U5033 (N_5033,In_1033,In_1833);
and U5034 (N_5034,In_108,In_1631);
or U5035 (N_5035,In_1759,In_156);
nor U5036 (N_5036,In_1529,In_505);
and U5037 (N_5037,In_515,In_147);
and U5038 (N_5038,In_1525,In_2429);
and U5039 (N_5039,In_1942,In_1545);
or U5040 (N_5040,In_1841,In_136);
and U5041 (N_5041,In_1753,In_153);
or U5042 (N_5042,In_86,In_1125);
nor U5043 (N_5043,In_870,In_1337);
and U5044 (N_5044,In_886,In_1420);
nand U5045 (N_5045,In_1600,In_1921);
or U5046 (N_5046,In_1229,In_368);
or U5047 (N_5047,In_517,In_2465);
and U5048 (N_5048,In_1498,In_175);
and U5049 (N_5049,In_878,In_2307);
and U5050 (N_5050,In_1119,In_669);
or U5051 (N_5051,In_1681,In_1154);
and U5052 (N_5052,In_1132,In_2234);
nand U5053 (N_5053,In_1852,In_34);
or U5054 (N_5054,In_198,In_108);
nand U5055 (N_5055,In_565,In_699);
and U5056 (N_5056,In_1151,In_776);
nor U5057 (N_5057,In_1679,In_2140);
nand U5058 (N_5058,In_579,In_1660);
or U5059 (N_5059,In_2113,In_2006);
or U5060 (N_5060,In_2348,In_1537);
and U5061 (N_5061,In_79,In_2084);
nand U5062 (N_5062,In_1107,In_841);
nor U5063 (N_5063,In_1756,In_872);
nor U5064 (N_5064,In_175,In_799);
nor U5065 (N_5065,In_66,In_36);
nand U5066 (N_5066,In_785,In_1122);
and U5067 (N_5067,In_1153,In_1449);
and U5068 (N_5068,In_314,In_2458);
or U5069 (N_5069,In_356,In_2462);
and U5070 (N_5070,In_2166,In_500);
and U5071 (N_5071,In_1722,In_1517);
nand U5072 (N_5072,In_885,In_2093);
and U5073 (N_5073,In_1791,In_1107);
and U5074 (N_5074,In_666,In_2058);
xnor U5075 (N_5075,In_2025,In_1522);
or U5076 (N_5076,In_1168,In_2269);
nand U5077 (N_5077,In_767,In_2065);
nor U5078 (N_5078,In_116,In_794);
or U5079 (N_5079,In_2349,In_616);
nand U5080 (N_5080,In_2083,In_2044);
nor U5081 (N_5081,In_1076,In_570);
or U5082 (N_5082,In_576,In_2428);
nand U5083 (N_5083,In_836,In_986);
nor U5084 (N_5084,In_2431,In_658);
or U5085 (N_5085,In_1515,In_501);
nand U5086 (N_5086,In_2095,In_517);
or U5087 (N_5087,In_1116,In_1606);
nor U5088 (N_5088,In_685,In_101);
or U5089 (N_5089,In_939,In_2134);
or U5090 (N_5090,In_698,In_126);
and U5091 (N_5091,In_2438,In_407);
nand U5092 (N_5092,In_1169,In_1585);
and U5093 (N_5093,In_2396,In_1520);
xnor U5094 (N_5094,In_1475,In_2317);
or U5095 (N_5095,In_1628,In_1180);
or U5096 (N_5096,In_1517,In_1258);
and U5097 (N_5097,In_2174,In_1090);
or U5098 (N_5098,In_1220,In_1134);
nand U5099 (N_5099,In_208,In_1979);
nor U5100 (N_5100,In_493,In_1604);
and U5101 (N_5101,In_205,In_1746);
and U5102 (N_5102,In_2189,In_1988);
nand U5103 (N_5103,In_322,In_2210);
nand U5104 (N_5104,In_833,In_1029);
and U5105 (N_5105,In_1953,In_1053);
nand U5106 (N_5106,In_945,In_2163);
nor U5107 (N_5107,In_2497,In_1370);
and U5108 (N_5108,In_2121,In_786);
or U5109 (N_5109,In_1502,In_931);
nor U5110 (N_5110,In_2133,In_403);
and U5111 (N_5111,In_962,In_1361);
nor U5112 (N_5112,In_755,In_2143);
and U5113 (N_5113,In_1887,In_1382);
nand U5114 (N_5114,In_1148,In_1949);
nand U5115 (N_5115,In_275,In_92);
nor U5116 (N_5116,In_843,In_1091);
or U5117 (N_5117,In_636,In_1594);
or U5118 (N_5118,In_2250,In_644);
and U5119 (N_5119,In_530,In_1089);
nand U5120 (N_5120,In_1129,In_1533);
and U5121 (N_5121,In_914,In_2430);
and U5122 (N_5122,In_27,In_1556);
nand U5123 (N_5123,In_2313,In_440);
or U5124 (N_5124,In_1543,In_2096);
or U5125 (N_5125,In_1163,In_2229);
nor U5126 (N_5126,In_1617,In_1499);
nand U5127 (N_5127,In_925,In_316);
or U5128 (N_5128,In_246,In_324);
nand U5129 (N_5129,In_874,In_1900);
or U5130 (N_5130,In_511,In_1393);
nor U5131 (N_5131,In_1549,In_1592);
and U5132 (N_5132,In_626,In_1224);
or U5133 (N_5133,In_11,In_481);
nand U5134 (N_5134,In_1992,In_527);
nand U5135 (N_5135,In_731,In_436);
or U5136 (N_5136,In_767,In_879);
and U5137 (N_5137,In_123,In_325);
nor U5138 (N_5138,In_1649,In_1802);
nand U5139 (N_5139,In_472,In_909);
and U5140 (N_5140,In_374,In_1007);
nand U5141 (N_5141,In_2464,In_2471);
nand U5142 (N_5142,In_445,In_961);
nand U5143 (N_5143,In_1932,In_1518);
and U5144 (N_5144,In_1751,In_1509);
and U5145 (N_5145,In_1885,In_1613);
nor U5146 (N_5146,In_179,In_1953);
and U5147 (N_5147,In_1452,In_1829);
nand U5148 (N_5148,In_960,In_655);
nor U5149 (N_5149,In_921,In_616);
or U5150 (N_5150,In_821,In_1277);
nor U5151 (N_5151,In_1423,In_2370);
xnor U5152 (N_5152,In_656,In_1575);
and U5153 (N_5153,In_2101,In_1965);
nor U5154 (N_5154,In_274,In_655);
nand U5155 (N_5155,In_2004,In_1454);
and U5156 (N_5156,In_1332,In_167);
and U5157 (N_5157,In_903,In_650);
or U5158 (N_5158,In_1870,In_467);
nor U5159 (N_5159,In_2199,In_84);
nand U5160 (N_5160,In_2495,In_131);
and U5161 (N_5161,In_2013,In_1605);
and U5162 (N_5162,In_2263,In_1236);
nand U5163 (N_5163,In_2171,In_1020);
or U5164 (N_5164,In_2387,In_119);
nor U5165 (N_5165,In_2411,In_1470);
nand U5166 (N_5166,In_2143,In_201);
nand U5167 (N_5167,In_61,In_1178);
nand U5168 (N_5168,In_1182,In_1514);
or U5169 (N_5169,In_1791,In_681);
nor U5170 (N_5170,In_961,In_598);
and U5171 (N_5171,In_1719,In_143);
or U5172 (N_5172,In_1613,In_1661);
nor U5173 (N_5173,In_957,In_2210);
nand U5174 (N_5174,In_773,In_1379);
nand U5175 (N_5175,In_487,In_1634);
nor U5176 (N_5176,In_1981,In_2418);
and U5177 (N_5177,In_2057,In_2099);
nand U5178 (N_5178,In_1834,In_802);
nand U5179 (N_5179,In_1248,In_2249);
or U5180 (N_5180,In_1145,In_147);
or U5181 (N_5181,In_747,In_61);
nor U5182 (N_5182,In_1310,In_896);
or U5183 (N_5183,In_693,In_1446);
nand U5184 (N_5184,In_1612,In_1725);
nor U5185 (N_5185,In_2274,In_1774);
nand U5186 (N_5186,In_567,In_1419);
nor U5187 (N_5187,In_1885,In_1200);
and U5188 (N_5188,In_2248,In_853);
nand U5189 (N_5189,In_2278,In_1366);
nor U5190 (N_5190,In_1675,In_315);
or U5191 (N_5191,In_2422,In_1367);
and U5192 (N_5192,In_1983,In_2402);
or U5193 (N_5193,In_1955,In_1645);
or U5194 (N_5194,In_319,In_4);
or U5195 (N_5195,In_252,In_1887);
and U5196 (N_5196,In_466,In_1241);
nor U5197 (N_5197,In_287,In_1193);
or U5198 (N_5198,In_1042,In_129);
nor U5199 (N_5199,In_2068,In_1237);
and U5200 (N_5200,In_414,In_1991);
nor U5201 (N_5201,In_1087,In_1320);
and U5202 (N_5202,In_1758,In_1653);
or U5203 (N_5203,In_1823,In_473);
and U5204 (N_5204,In_1373,In_657);
nand U5205 (N_5205,In_1138,In_632);
and U5206 (N_5206,In_205,In_1591);
nand U5207 (N_5207,In_1819,In_1823);
nand U5208 (N_5208,In_1049,In_1025);
xnor U5209 (N_5209,In_618,In_156);
and U5210 (N_5210,In_1966,In_1355);
nand U5211 (N_5211,In_274,In_2457);
and U5212 (N_5212,In_1057,In_318);
nand U5213 (N_5213,In_1963,In_256);
nand U5214 (N_5214,In_1230,In_1132);
xor U5215 (N_5215,In_288,In_313);
or U5216 (N_5216,In_1074,In_1078);
and U5217 (N_5217,In_1628,In_942);
nor U5218 (N_5218,In_1185,In_2287);
or U5219 (N_5219,In_1170,In_1046);
and U5220 (N_5220,In_1078,In_2407);
or U5221 (N_5221,In_1013,In_2264);
and U5222 (N_5222,In_1898,In_1903);
nor U5223 (N_5223,In_667,In_2429);
nand U5224 (N_5224,In_903,In_2344);
or U5225 (N_5225,In_1074,In_1550);
nand U5226 (N_5226,In_798,In_894);
and U5227 (N_5227,In_1674,In_172);
nor U5228 (N_5228,In_955,In_1518);
and U5229 (N_5229,In_1920,In_1225);
or U5230 (N_5230,In_1899,In_141);
and U5231 (N_5231,In_888,In_2494);
nand U5232 (N_5232,In_2228,In_660);
and U5233 (N_5233,In_1719,In_1270);
nor U5234 (N_5234,In_989,In_2460);
nand U5235 (N_5235,In_1202,In_1759);
nand U5236 (N_5236,In_2383,In_2134);
and U5237 (N_5237,In_690,In_1951);
and U5238 (N_5238,In_1914,In_1367);
and U5239 (N_5239,In_171,In_517);
nand U5240 (N_5240,In_1749,In_2111);
nor U5241 (N_5241,In_1524,In_1972);
or U5242 (N_5242,In_1817,In_195);
nor U5243 (N_5243,In_2497,In_1327);
nor U5244 (N_5244,In_249,In_1698);
and U5245 (N_5245,In_35,In_1201);
or U5246 (N_5246,In_281,In_2015);
or U5247 (N_5247,In_1229,In_575);
and U5248 (N_5248,In_1791,In_269);
or U5249 (N_5249,In_1826,In_101);
nand U5250 (N_5250,In_899,In_1359);
nand U5251 (N_5251,In_672,In_1055);
and U5252 (N_5252,In_245,In_2193);
and U5253 (N_5253,In_348,In_1538);
and U5254 (N_5254,In_733,In_2237);
xnor U5255 (N_5255,In_1189,In_1014);
or U5256 (N_5256,In_1952,In_2027);
nor U5257 (N_5257,In_2176,In_1155);
and U5258 (N_5258,In_1035,In_2484);
nor U5259 (N_5259,In_1098,In_1205);
nand U5260 (N_5260,In_263,In_1452);
nor U5261 (N_5261,In_1739,In_1345);
and U5262 (N_5262,In_1367,In_587);
or U5263 (N_5263,In_1823,In_293);
or U5264 (N_5264,In_941,In_186);
or U5265 (N_5265,In_16,In_823);
or U5266 (N_5266,In_240,In_962);
nor U5267 (N_5267,In_795,In_2259);
or U5268 (N_5268,In_428,In_2375);
or U5269 (N_5269,In_2177,In_1679);
nand U5270 (N_5270,In_1483,In_227);
nor U5271 (N_5271,In_2260,In_1010);
nand U5272 (N_5272,In_722,In_1728);
nor U5273 (N_5273,In_488,In_2140);
nor U5274 (N_5274,In_765,In_699);
nor U5275 (N_5275,In_2124,In_660);
nor U5276 (N_5276,In_1982,In_871);
or U5277 (N_5277,In_2355,In_2472);
or U5278 (N_5278,In_1046,In_675);
and U5279 (N_5279,In_1977,In_2010);
nor U5280 (N_5280,In_1307,In_1491);
and U5281 (N_5281,In_1843,In_2012);
or U5282 (N_5282,In_2175,In_340);
or U5283 (N_5283,In_776,In_39);
and U5284 (N_5284,In_727,In_786);
or U5285 (N_5285,In_1705,In_883);
or U5286 (N_5286,In_1703,In_1444);
nor U5287 (N_5287,In_2290,In_2327);
nor U5288 (N_5288,In_1778,In_1437);
or U5289 (N_5289,In_455,In_406);
nand U5290 (N_5290,In_1992,In_3);
and U5291 (N_5291,In_1473,In_694);
nor U5292 (N_5292,In_38,In_153);
nor U5293 (N_5293,In_2362,In_2233);
or U5294 (N_5294,In_1919,In_1149);
nand U5295 (N_5295,In_2315,In_427);
nand U5296 (N_5296,In_2314,In_973);
nor U5297 (N_5297,In_951,In_1633);
nor U5298 (N_5298,In_1386,In_2455);
or U5299 (N_5299,In_2015,In_1535);
or U5300 (N_5300,In_122,In_807);
or U5301 (N_5301,In_2153,In_2386);
or U5302 (N_5302,In_1194,In_283);
nor U5303 (N_5303,In_2389,In_1219);
and U5304 (N_5304,In_1852,In_941);
nand U5305 (N_5305,In_103,In_1256);
and U5306 (N_5306,In_578,In_2342);
or U5307 (N_5307,In_850,In_2038);
and U5308 (N_5308,In_1001,In_1593);
nand U5309 (N_5309,In_2005,In_594);
nand U5310 (N_5310,In_1615,In_1245);
nor U5311 (N_5311,In_1075,In_2227);
xor U5312 (N_5312,In_1311,In_32);
nor U5313 (N_5313,In_109,In_1498);
nand U5314 (N_5314,In_660,In_617);
nor U5315 (N_5315,In_1606,In_852);
nor U5316 (N_5316,In_2211,In_2031);
and U5317 (N_5317,In_1087,In_108);
nor U5318 (N_5318,In_340,In_87);
nor U5319 (N_5319,In_772,In_1747);
nand U5320 (N_5320,In_329,In_171);
or U5321 (N_5321,In_1508,In_2022);
nand U5322 (N_5322,In_698,In_897);
nor U5323 (N_5323,In_1880,In_1878);
nand U5324 (N_5324,In_1177,In_1239);
nor U5325 (N_5325,In_1409,In_2449);
and U5326 (N_5326,In_25,In_919);
nand U5327 (N_5327,In_1852,In_1076);
nand U5328 (N_5328,In_240,In_1087);
and U5329 (N_5329,In_1635,In_2186);
or U5330 (N_5330,In_2142,In_1586);
nor U5331 (N_5331,In_727,In_1437);
nand U5332 (N_5332,In_1564,In_1933);
and U5333 (N_5333,In_1357,In_740);
nand U5334 (N_5334,In_2356,In_1645);
or U5335 (N_5335,In_2194,In_1519);
or U5336 (N_5336,In_1454,In_1966);
and U5337 (N_5337,In_2310,In_1230);
nand U5338 (N_5338,In_1681,In_1713);
nor U5339 (N_5339,In_2281,In_2405);
nand U5340 (N_5340,In_862,In_204);
or U5341 (N_5341,In_2243,In_1200);
nor U5342 (N_5342,In_904,In_1771);
nor U5343 (N_5343,In_1575,In_2389);
or U5344 (N_5344,In_151,In_345);
nand U5345 (N_5345,In_603,In_1738);
nand U5346 (N_5346,In_1939,In_1409);
xor U5347 (N_5347,In_1097,In_1320);
and U5348 (N_5348,In_1409,In_624);
nor U5349 (N_5349,In_1221,In_150);
and U5350 (N_5350,In_221,In_739);
or U5351 (N_5351,In_644,In_2340);
nand U5352 (N_5352,In_2020,In_799);
and U5353 (N_5353,In_2432,In_184);
and U5354 (N_5354,In_231,In_835);
or U5355 (N_5355,In_756,In_1047);
or U5356 (N_5356,In_1318,In_1819);
and U5357 (N_5357,In_1877,In_2023);
and U5358 (N_5358,In_732,In_1374);
nor U5359 (N_5359,In_2041,In_802);
nor U5360 (N_5360,In_1614,In_787);
and U5361 (N_5361,In_727,In_319);
or U5362 (N_5362,In_2076,In_790);
or U5363 (N_5363,In_1148,In_1871);
or U5364 (N_5364,In_1157,In_759);
nor U5365 (N_5365,In_2267,In_327);
or U5366 (N_5366,In_687,In_1230);
and U5367 (N_5367,In_2247,In_1304);
nand U5368 (N_5368,In_2403,In_2022);
nand U5369 (N_5369,In_923,In_647);
or U5370 (N_5370,In_2166,In_1167);
or U5371 (N_5371,In_1210,In_2008);
nor U5372 (N_5372,In_349,In_1260);
nor U5373 (N_5373,In_1453,In_1764);
nand U5374 (N_5374,In_274,In_1979);
and U5375 (N_5375,In_1888,In_597);
and U5376 (N_5376,In_794,In_304);
or U5377 (N_5377,In_478,In_1812);
nor U5378 (N_5378,In_2170,In_2085);
nand U5379 (N_5379,In_150,In_530);
nand U5380 (N_5380,In_717,In_71);
and U5381 (N_5381,In_1539,In_296);
nand U5382 (N_5382,In_994,In_1499);
nand U5383 (N_5383,In_1691,In_1697);
and U5384 (N_5384,In_1692,In_1875);
and U5385 (N_5385,In_1477,In_1222);
nand U5386 (N_5386,In_148,In_122);
nor U5387 (N_5387,In_1455,In_1494);
or U5388 (N_5388,In_1832,In_446);
nor U5389 (N_5389,In_1712,In_1709);
and U5390 (N_5390,In_57,In_2013);
and U5391 (N_5391,In_675,In_1493);
nor U5392 (N_5392,In_2432,In_1797);
nand U5393 (N_5393,In_2444,In_2320);
and U5394 (N_5394,In_2143,In_1556);
nand U5395 (N_5395,In_1506,In_524);
nor U5396 (N_5396,In_1021,In_850);
nand U5397 (N_5397,In_1626,In_1562);
nor U5398 (N_5398,In_1476,In_1750);
nor U5399 (N_5399,In_312,In_356);
or U5400 (N_5400,In_509,In_1488);
and U5401 (N_5401,In_874,In_1832);
nand U5402 (N_5402,In_1324,In_2094);
and U5403 (N_5403,In_1049,In_391);
and U5404 (N_5404,In_899,In_181);
and U5405 (N_5405,In_585,In_706);
or U5406 (N_5406,In_696,In_433);
nand U5407 (N_5407,In_2107,In_856);
nand U5408 (N_5408,In_483,In_1880);
and U5409 (N_5409,In_1442,In_2382);
nand U5410 (N_5410,In_1336,In_913);
nand U5411 (N_5411,In_1612,In_1165);
nand U5412 (N_5412,In_1816,In_1156);
nand U5413 (N_5413,In_972,In_445);
nand U5414 (N_5414,In_1428,In_1748);
and U5415 (N_5415,In_1291,In_1277);
and U5416 (N_5416,In_526,In_1066);
or U5417 (N_5417,In_304,In_2114);
nor U5418 (N_5418,In_1609,In_2308);
nor U5419 (N_5419,In_262,In_1267);
and U5420 (N_5420,In_893,In_1857);
and U5421 (N_5421,In_56,In_1919);
nand U5422 (N_5422,In_731,In_766);
nor U5423 (N_5423,In_798,In_967);
and U5424 (N_5424,In_503,In_2030);
nand U5425 (N_5425,In_478,In_431);
nand U5426 (N_5426,In_578,In_1037);
and U5427 (N_5427,In_2044,In_2326);
xor U5428 (N_5428,In_1994,In_1904);
nand U5429 (N_5429,In_1017,In_98);
or U5430 (N_5430,In_838,In_575);
nor U5431 (N_5431,In_1376,In_1046);
xnor U5432 (N_5432,In_1863,In_996);
nand U5433 (N_5433,In_140,In_1685);
or U5434 (N_5434,In_1980,In_270);
or U5435 (N_5435,In_1569,In_1851);
nor U5436 (N_5436,In_2207,In_1470);
nand U5437 (N_5437,In_1119,In_1980);
nand U5438 (N_5438,In_2348,In_695);
nand U5439 (N_5439,In_476,In_209);
nor U5440 (N_5440,In_324,In_1280);
nand U5441 (N_5441,In_2029,In_1696);
or U5442 (N_5442,In_1395,In_383);
or U5443 (N_5443,In_979,In_1487);
and U5444 (N_5444,In_404,In_487);
or U5445 (N_5445,In_621,In_2479);
or U5446 (N_5446,In_1688,In_2284);
and U5447 (N_5447,In_942,In_2309);
nand U5448 (N_5448,In_2472,In_1027);
and U5449 (N_5449,In_2418,In_807);
or U5450 (N_5450,In_1384,In_1918);
or U5451 (N_5451,In_601,In_785);
and U5452 (N_5452,In_1246,In_1039);
nor U5453 (N_5453,In_349,In_793);
and U5454 (N_5454,In_1381,In_2228);
or U5455 (N_5455,In_1333,In_1617);
nor U5456 (N_5456,In_762,In_2341);
and U5457 (N_5457,In_2009,In_694);
or U5458 (N_5458,In_1050,In_265);
nor U5459 (N_5459,In_1315,In_2045);
nand U5460 (N_5460,In_2252,In_463);
nand U5461 (N_5461,In_695,In_555);
and U5462 (N_5462,In_2253,In_229);
xor U5463 (N_5463,In_668,In_2299);
nor U5464 (N_5464,In_1220,In_826);
or U5465 (N_5465,In_609,In_1859);
and U5466 (N_5466,In_2081,In_1967);
nand U5467 (N_5467,In_961,In_943);
or U5468 (N_5468,In_1374,In_492);
nor U5469 (N_5469,In_150,In_1482);
nand U5470 (N_5470,In_1501,In_1279);
nor U5471 (N_5471,In_2486,In_1080);
nand U5472 (N_5472,In_275,In_1377);
or U5473 (N_5473,In_1631,In_2483);
and U5474 (N_5474,In_1901,In_1538);
xnor U5475 (N_5475,In_1693,In_761);
nor U5476 (N_5476,In_2155,In_1310);
or U5477 (N_5477,In_171,In_1875);
and U5478 (N_5478,In_819,In_587);
or U5479 (N_5479,In_1792,In_1363);
or U5480 (N_5480,In_122,In_1041);
or U5481 (N_5481,In_512,In_422);
or U5482 (N_5482,In_413,In_237);
or U5483 (N_5483,In_1980,In_1684);
nand U5484 (N_5484,In_189,In_638);
or U5485 (N_5485,In_858,In_1301);
nor U5486 (N_5486,In_298,In_2070);
nand U5487 (N_5487,In_1743,In_1865);
nand U5488 (N_5488,In_93,In_2311);
and U5489 (N_5489,In_176,In_1600);
or U5490 (N_5490,In_1392,In_206);
nand U5491 (N_5491,In_1532,In_962);
nand U5492 (N_5492,In_2009,In_384);
nor U5493 (N_5493,In_1142,In_1561);
nand U5494 (N_5494,In_235,In_746);
or U5495 (N_5495,In_1686,In_2212);
or U5496 (N_5496,In_2105,In_545);
and U5497 (N_5497,In_924,In_2441);
and U5498 (N_5498,In_1622,In_73);
nor U5499 (N_5499,In_81,In_704);
nand U5500 (N_5500,In_2099,In_2323);
nand U5501 (N_5501,In_2236,In_2031);
nor U5502 (N_5502,In_2059,In_1718);
or U5503 (N_5503,In_1949,In_1165);
nor U5504 (N_5504,In_508,In_1674);
and U5505 (N_5505,In_2419,In_1835);
and U5506 (N_5506,In_369,In_2223);
or U5507 (N_5507,In_317,In_1139);
nor U5508 (N_5508,In_2291,In_1512);
or U5509 (N_5509,In_1205,In_1928);
nand U5510 (N_5510,In_1949,In_2393);
or U5511 (N_5511,In_224,In_614);
and U5512 (N_5512,In_156,In_1257);
nand U5513 (N_5513,In_1926,In_1661);
or U5514 (N_5514,In_1518,In_1384);
and U5515 (N_5515,In_2460,In_1256);
nand U5516 (N_5516,In_698,In_19);
or U5517 (N_5517,In_1937,In_2055);
nor U5518 (N_5518,In_2029,In_965);
and U5519 (N_5519,In_2192,In_2254);
nor U5520 (N_5520,In_1435,In_1394);
nand U5521 (N_5521,In_398,In_2418);
nor U5522 (N_5522,In_2329,In_20);
or U5523 (N_5523,In_1810,In_537);
and U5524 (N_5524,In_655,In_974);
and U5525 (N_5525,In_910,In_1194);
or U5526 (N_5526,In_93,In_1823);
nor U5527 (N_5527,In_592,In_370);
nand U5528 (N_5528,In_1183,In_1137);
nand U5529 (N_5529,In_1640,In_1218);
nand U5530 (N_5530,In_2398,In_289);
nand U5531 (N_5531,In_955,In_1481);
nor U5532 (N_5532,In_2137,In_1616);
and U5533 (N_5533,In_2270,In_842);
and U5534 (N_5534,In_656,In_2146);
and U5535 (N_5535,In_153,In_1701);
nand U5536 (N_5536,In_693,In_822);
nor U5537 (N_5537,In_932,In_2129);
or U5538 (N_5538,In_534,In_2248);
and U5539 (N_5539,In_843,In_1693);
nor U5540 (N_5540,In_699,In_516);
or U5541 (N_5541,In_513,In_1742);
nand U5542 (N_5542,In_1687,In_871);
or U5543 (N_5543,In_1016,In_1909);
nand U5544 (N_5544,In_346,In_1489);
nand U5545 (N_5545,In_1813,In_971);
nor U5546 (N_5546,In_858,In_803);
nand U5547 (N_5547,In_1197,In_1003);
and U5548 (N_5548,In_1107,In_1392);
nor U5549 (N_5549,In_1894,In_627);
and U5550 (N_5550,In_545,In_655);
xor U5551 (N_5551,In_1234,In_2340);
or U5552 (N_5552,In_435,In_2079);
nor U5553 (N_5553,In_143,In_1601);
and U5554 (N_5554,In_1053,In_1700);
and U5555 (N_5555,In_1244,In_1011);
nand U5556 (N_5556,In_2117,In_2404);
or U5557 (N_5557,In_524,In_104);
nand U5558 (N_5558,In_1521,In_332);
nor U5559 (N_5559,In_2281,In_2454);
nor U5560 (N_5560,In_314,In_684);
or U5561 (N_5561,In_775,In_1079);
nor U5562 (N_5562,In_1504,In_975);
nand U5563 (N_5563,In_2494,In_694);
nor U5564 (N_5564,In_1523,In_715);
and U5565 (N_5565,In_835,In_534);
nor U5566 (N_5566,In_93,In_1309);
nand U5567 (N_5567,In_2166,In_1496);
and U5568 (N_5568,In_1970,In_309);
xor U5569 (N_5569,In_755,In_2386);
or U5570 (N_5570,In_954,In_640);
nor U5571 (N_5571,In_1244,In_1937);
nor U5572 (N_5572,In_2466,In_2436);
nand U5573 (N_5573,In_222,In_627);
and U5574 (N_5574,In_625,In_495);
and U5575 (N_5575,In_2255,In_1609);
or U5576 (N_5576,In_631,In_1991);
and U5577 (N_5577,In_2488,In_2424);
nor U5578 (N_5578,In_128,In_1947);
and U5579 (N_5579,In_1072,In_2347);
and U5580 (N_5580,In_643,In_152);
or U5581 (N_5581,In_914,In_2227);
or U5582 (N_5582,In_1425,In_2107);
or U5583 (N_5583,In_34,In_344);
nand U5584 (N_5584,In_2352,In_1149);
or U5585 (N_5585,In_510,In_386);
nor U5586 (N_5586,In_1408,In_170);
xnor U5587 (N_5587,In_1629,In_2356);
nor U5588 (N_5588,In_1118,In_2179);
or U5589 (N_5589,In_554,In_2002);
or U5590 (N_5590,In_1683,In_727);
nand U5591 (N_5591,In_742,In_642);
and U5592 (N_5592,In_1161,In_1830);
nor U5593 (N_5593,In_1865,In_1176);
nand U5594 (N_5594,In_2239,In_82);
nor U5595 (N_5595,In_1609,In_1207);
nor U5596 (N_5596,In_2095,In_2081);
and U5597 (N_5597,In_12,In_1040);
nor U5598 (N_5598,In_1038,In_2106);
nand U5599 (N_5599,In_1909,In_462);
and U5600 (N_5600,In_643,In_2231);
nand U5601 (N_5601,In_1853,In_1330);
nand U5602 (N_5602,In_631,In_2007);
or U5603 (N_5603,In_1574,In_1721);
nor U5604 (N_5604,In_1874,In_191);
or U5605 (N_5605,In_846,In_593);
or U5606 (N_5606,In_1255,In_2450);
xor U5607 (N_5607,In_717,In_579);
nand U5608 (N_5608,In_1605,In_1204);
nor U5609 (N_5609,In_169,In_267);
and U5610 (N_5610,In_1536,In_2494);
or U5611 (N_5611,In_1761,In_1464);
nand U5612 (N_5612,In_2011,In_1482);
nand U5613 (N_5613,In_165,In_1375);
or U5614 (N_5614,In_1453,In_1684);
nor U5615 (N_5615,In_1807,In_1823);
and U5616 (N_5616,In_583,In_238);
nand U5617 (N_5617,In_1198,In_1232);
or U5618 (N_5618,In_1862,In_2000);
nor U5619 (N_5619,In_883,In_1122);
nand U5620 (N_5620,In_595,In_2450);
and U5621 (N_5621,In_1163,In_815);
nor U5622 (N_5622,In_356,In_4);
nor U5623 (N_5623,In_366,In_2194);
or U5624 (N_5624,In_323,In_2126);
and U5625 (N_5625,In_1022,In_827);
nand U5626 (N_5626,In_2398,In_1184);
or U5627 (N_5627,In_879,In_275);
or U5628 (N_5628,In_560,In_908);
nand U5629 (N_5629,In_2122,In_1319);
nor U5630 (N_5630,In_2175,In_1277);
and U5631 (N_5631,In_1422,In_406);
nand U5632 (N_5632,In_708,In_132);
nor U5633 (N_5633,In_2179,In_982);
nor U5634 (N_5634,In_1785,In_2407);
nor U5635 (N_5635,In_860,In_1911);
and U5636 (N_5636,In_2147,In_1358);
nand U5637 (N_5637,In_1605,In_560);
or U5638 (N_5638,In_1785,In_2165);
nand U5639 (N_5639,In_1153,In_2268);
nand U5640 (N_5640,In_1311,In_1902);
nor U5641 (N_5641,In_413,In_1297);
xnor U5642 (N_5642,In_2370,In_15);
nor U5643 (N_5643,In_1410,In_1083);
or U5644 (N_5644,In_233,In_1526);
or U5645 (N_5645,In_1716,In_426);
nor U5646 (N_5646,In_922,In_1137);
and U5647 (N_5647,In_2089,In_1378);
nand U5648 (N_5648,In_2435,In_1880);
and U5649 (N_5649,In_1901,In_1529);
nand U5650 (N_5650,In_451,In_2040);
and U5651 (N_5651,In_1609,In_1005);
nor U5652 (N_5652,In_1130,In_1579);
nand U5653 (N_5653,In_921,In_1500);
nor U5654 (N_5654,In_691,In_1610);
and U5655 (N_5655,In_1021,In_1836);
nand U5656 (N_5656,In_465,In_411);
or U5657 (N_5657,In_137,In_838);
nor U5658 (N_5658,In_682,In_33);
xor U5659 (N_5659,In_1357,In_1811);
nand U5660 (N_5660,In_1222,In_226);
nor U5661 (N_5661,In_468,In_1244);
or U5662 (N_5662,In_224,In_2465);
or U5663 (N_5663,In_966,In_1827);
nand U5664 (N_5664,In_775,In_1436);
nand U5665 (N_5665,In_7,In_233);
nand U5666 (N_5666,In_840,In_386);
and U5667 (N_5667,In_498,In_15);
or U5668 (N_5668,In_343,In_418);
or U5669 (N_5669,In_1288,In_437);
or U5670 (N_5670,In_1180,In_215);
and U5671 (N_5671,In_2262,In_676);
and U5672 (N_5672,In_1420,In_1830);
nor U5673 (N_5673,In_2374,In_855);
nor U5674 (N_5674,In_1184,In_24);
and U5675 (N_5675,In_123,In_1648);
or U5676 (N_5676,In_2135,In_460);
nand U5677 (N_5677,In_453,In_1544);
and U5678 (N_5678,In_1453,In_1871);
or U5679 (N_5679,In_129,In_901);
nand U5680 (N_5680,In_951,In_691);
and U5681 (N_5681,In_243,In_1800);
or U5682 (N_5682,In_1987,In_328);
or U5683 (N_5683,In_2372,In_1585);
or U5684 (N_5684,In_1788,In_1522);
nor U5685 (N_5685,In_2133,In_284);
or U5686 (N_5686,In_1023,In_1931);
or U5687 (N_5687,In_494,In_445);
nand U5688 (N_5688,In_242,In_413);
nor U5689 (N_5689,In_822,In_2213);
or U5690 (N_5690,In_488,In_929);
nand U5691 (N_5691,In_1183,In_624);
and U5692 (N_5692,In_1582,In_661);
and U5693 (N_5693,In_2415,In_2315);
nor U5694 (N_5694,In_785,In_1593);
nor U5695 (N_5695,In_1974,In_653);
nand U5696 (N_5696,In_1140,In_544);
and U5697 (N_5697,In_1392,In_65);
and U5698 (N_5698,In_54,In_2192);
and U5699 (N_5699,In_950,In_1348);
nand U5700 (N_5700,In_1579,In_495);
or U5701 (N_5701,In_1546,In_131);
nand U5702 (N_5702,In_1253,In_2431);
nor U5703 (N_5703,In_198,In_502);
nor U5704 (N_5704,In_871,In_164);
or U5705 (N_5705,In_156,In_1629);
and U5706 (N_5706,In_2070,In_387);
nor U5707 (N_5707,In_736,In_1596);
nor U5708 (N_5708,In_316,In_284);
nor U5709 (N_5709,In_1132,In_579);
nand U5710 (N_5710,In_2083,In_2498);
or U5711 (N_5711,In_1017,In_840);
nor U5712 (N_5712,In_1879,In_2294);
or U5713 (N_5713,In_2011,In_1939);
nand U5714 (N_5714,In_431,In_953);
and U5715 (N_5715,In_1949,In_1830);
nor U5716 (N_5716,In_486,In_1420);
and U5717 (N_5717,In_756,In_2250);
or U5718 (N_5718,In_2355,In_47);
and U5719 (N_5719,In_1198,In_1710);
nor U5720 (N_5720,In_1353,In_793);
or U5721 (N_5721,In_928,In_2282);
nor U5722 (N_5722,In_2200,In_2066);
nand U5723 (N_5723,In_1175,In_832);
nor U5724 (N_5724,In_1331,In_650);
nor U5725 (N_5725,In_1372,In_513);
or U5726 (N_5726,In_243,In_1256);
and U5727 (N_5727,In_1549,In_374);
nand U5728 (N_5728,In_2329,In_57);
nand U5729 (N_5729,In_1452,In_506);
and U5730 (N_5730,In_905,In_271);
and U5731 (N_5731,In_129,In_259);
nor U5732 (N_5732,In_2219,In_2150);
or U5733 (N_5733,In_451,In_773);
or U5734 (N_5734,In_1567,In_491);
or U5735 (N_5735,In_121,In_933);
nand U5736 (N_5736,In_1069,In_1176);
xnor U5737 (N_5737,In_663,In_956);
nand U5738 (N_5738,In_1909,In_279);
or U5739 (N_5739,In_2364,In_2214);
nand U5740 (N_5740,In_1213,In_2010);
nor U5741 (N_5741,In_710,In_2405);
nor U5742 (N_5742,In_1536,In_826);
nor U5743 (N_5743,In_2305,In_2399);
and U5744 (N_5744,In_1643,In_195);
nand U5745 (N_5745,In_1646,In_2309);
nand U5746 (N_5746,In_1776,In_1593);
and U5747 (N_5747,In_2123,In_1816);
and U5748 (N_5748,In_1021,In_2449);
and U5749 (N_5749,In_1986,In_1994);
nand U5750 (N_5750,In_865,In_219);
and U5751 (N_5751,In_2383,In_122);
nor U5752 (N_5752,In_2106,In_653);
or U5753 (N_5753,In_1990,In_827);
or U5754 (N_5754,In_1507,In_1315);
or U5755 (N_5755,In_1021,In_1444);
and U5756 (N_5756,In_1052,In_2129);
nor U5757 (N_5757,In_735,In_1276);
nor U5758 (N_5758,In_1634,In_1694);
and U5759 (N_5759,In_1390,In_2232);
or U5760 (N_5760,In_2377,In_2367);
nor U5761 (N_5761,In_717,In_802);
and U5762 (N_5762,In_1843,In_700);
or U5763 (N_5763,In_1832,In_2048);
nand U5764 (N_5764,In_394,In_258);
xnor U5765 (N_5765,In_2346,In_528);
and U5766 (N_5766,In_93,In_586);
nor U5767 (N_5767,In_1011,In_215);
xnor U5768 (N_5768,In_1551,In_1750);
nor U5769 (N_5769,In_1197,In_1897);
nor U5770 (N_5770,In_1996,In_365);
or U5771 (N_5771,In_917,In_2074);
nand U5772 (N_5772,In_1217,In_265);
nand U5773 (N_5773,In_765,In_323);
xnor U5774 (N_5774,In_505,In_686);
or U5775 (N_5775,In_1219,In_1761);
nor U5776 (N_5776,In_555,In_591);
and U5777 (N_5777,In_627,In_1778);
and U5778 (N_5778,In_1881,In_1887);
and U5779 (N_5779,In_1791,In_1463);
or U5780 (N_5780,In_2488,In_2013);
and U5781 (N_5781,In_801,In_712);
and U5782 (N_5782,In_1602,In_1580);
or U5783 (N_5783,In_1120,In_1029);
or U5784 (N_5784,In_824,In_270);
or U5785 (N_5785,In_1893,In_1347);
and U5786 (N_5786,In_622,In_1886);
nor U5787 (N_5787,In_1288,In_32);
nor U5788 (N_5788,In_2196,In_271);
and U5789 (N_5789,In_1636,In_2234);
nand U5790 (N_5790,In_80,In_1510);
and U5791 (N_5791,In_1345,In_203);
or U5792 (N_5792,In_630,In_1921);
xor U5793 (N_5793,In_1639,In_121);
and U5794 (N_5794,In_2463,In_257);
nand U5795 (N_5795,In_1870,In_1513);
or U5796 (N_5796,In_1630,In_1184);
and U5797 (N_5797,In_1608,In_318);
and U5798 (N_5798,In_374,In_1768);
nand U5799 (N_5799,In_1270,In_619);
nor U5800 (N_5800,In_121,In_8);
nor U5801 (N_5801,In_16,In_1782);
and U5802 (N_5802,In_2320,In_1470);
or U5803 (N_5803,In_859,In_918);
nor U5804 (N_5804,In_509,In_423);
xor U5805 (N_5805,In_232,In_2);
or U5806 (N_5806,In_2364,In_1958);
and U5807 (N_5807,In_364,In_710);
and U5808 (N_5808,In_1732,In_709);
and U5809 (N_5809,In_1374,In_2156);
nor U5810 (N_5810,In_1254,In_290);
and U5811 (N_5811,In_157,In_192);
nand U5812 (N_5812,In_2105,In_2179);
xor U5813 (N_5813,In_2341,In_1282);
nand U5814 (N_5814,In_911,In_313);
nand U5815 (N_5815,In_2193,In_1700);
nand U5816 (N_5816,In_141,In_512);
nand U5817 (N_5817,In_1343,In_361);
nand U5818 (N_5818,In_363,In_592);
nor U5819 (N_5819,In_428,In_1837);
or U5820 (N_5820,In_1172,In_2141);
or U5821 (N_5821,In_1072,In_1614);
or U5822 (N_5822,In_2158,In_937);
and U5823 (N_5823,In_1682,In_1224);
or U5824 (N_5824,In_1786,In_1229);
or U5825 (N_5825,In_135,In_1251);
or U5826 (N_5826,In_96,In_1239);
or U5827 (N_5827,In_1272,In_54);
and U5828 (N_5828,In_1677,In_959);
or U5829 (N_5829,In_997,In_800);
nand U5830 (N_5830,In_1334,In_1624);
nor U5831 (N_5831,In_465,In_820);
nor U5832 (N_5832,In_1703,In_2452);
nor U5833 (N_5833,In_729,In_1059);
xor U5834 (N_5834,In_329,In_1288);
nor U5835 (N_5835,In_2365,In_55);
or U5836 (N_5836,In_2059,In_1490);
nand U5837 (N_5837,In_746,In_1936);
and U5838 (N_5838,In_1776,In_919);
and U5839 (N_5839,In_982,In_2457);
nor U5840 (N_5840,In_263,In_1858);
and U5841 (N_5841,In_400,In_1991);
and U5842 (N_5842,In_271,In_1895);
or U5843 (N_5843,In_166,In_1212);
nand U5844 (N_5844,In_1092,In_2249);
or U5845 (N_5845,In_1418,In_2304);
nand U5846 (N_5846,In_2137,In_1648);
and U5847 (N_5847,In_1558,In_1369);
nor U5848 (N_5848,In_1101,In_373);
nand U5849 (N_5849,In_974,In_1098);
or U5850 (N_5850,In_1886,In_1388);
or U5851 (N_5851,In_1973,In_297);
and U5852 (N_5852,In_1993,In_1600);
or U5853 (N_5853,In_409,In_1512);
nor U5854 (N_5854,In_379,In_483);
nand U5855 (N_5855,In_1335,In_1943);
or U5856 (N_5856,In_1654,In_1062);
nand U5857 (N_5857,In_9,In_2284);
or U5858 (N_5858,In_2192,In_1494);
nand U5859 (N_5859,In_1505,In_157);
or U5860 (N_5860,In_177,In_2006);
xor U5861 (N_5861,In_345,In_1904);
nand U5862 (N_5862,In_308,In_1547);
nand U5863 (N_5863,In_499,In_1453);
and U5864 (N_5864,In_49,In_1052);
and U5865 (N_5865,In_1348,In_2363);
and U5866 (N_5866,In_401,In_652);
nor U5867 (N_5867,In_133,In_774);
or U5868 (N_5868,In_1918,In_2071);
nand U5869 (N_5869,In_689,In_802);
nor U5870 (N_5870,In_472,In_4);
and U5871 (N_5871,In_1297,In_2309);
nand U5872 (N_5872,In_2019,In_2471);
or U5873 (N_5873,In_476,In_735);
nor U5874 (N_5874,In_667,In_2022);
or U5875 (N_5875,In_1333,In_1324);
and U5876 (N_5876,In_388,In_109);
and U5877 (N_5877,In_402,In_407);
or U5878 (N_5878,In_2197,In_2292);
and U5879 (N_5879,In_428,In_2073);
or U5880 (N_5880,In_816,In_285);
nor U5881 (N_5881,In_496,In_2459);
nor U5882 (N_5882,In_1586,In_784);
nand U5883 (N_5883,In_2292,In_995);
or U5884 (N_5884,In_146,In_2494);
nand U5885 (N_5885,In_1252,In_2446);
or U5886 (N_5886,In_306,In_284);
or U5887 (N_5887,In_1385,In_797);
or U5888 (N_5888,In_1349,In_689);
and U5889 (N_5889,In_2473,In_1315);
nand U5890 (N_5890,In_1047,In_1906);
nor U5891 (N_5891,In_495,In_277);
nand U5892 (N_5892,In_591,In_1903);
nor U5893 (N_5893,In_1008,In_2188);
nand U5894 (N_5894,In_833,In_1891);
xnor U5895 (N_5895,In_1672,In_1942);
or U5896 (N_5896,In_2337,In_1694);
or U5897 (N_5897,In_605,In_1643);
nor U5898 (N_5898,In_1965,In_2490);
nand U5899 (N_5899,In_2429,In_101);
nand U5900 (N_5900,In_1431,In_2249);
and U5901 (N_5901,In_961,In_2005);
and U5902 (N_5902,In_919,In_189);
and U5903 (N_5903,In_584,In_762);
and U5904 (N_5904,In_2423,In_595);
and U5905 (N_5905,In_1443,In_641);
nand U5906 (N_5906,In_360,In_281);
nor U5907 (N_5907,In_165,In_2294);
nor U5908 (N_5908,In_1457,In_1917);
nand U5909 (N_5909,In_1871,In_2226);
nor U5910 (N_5910,In_1173,In_603);
nor U5911 (N_5911,In_330,In_573);
xnor U5912 (N_5912,In_2297,In_583);
and U5913 (N_5913,In_2051,In_1921);
or U5914 (N_5914,In_1293,In_449);
or U5915 (N_5915,In_1521,In_1347);
and U5916 (N_5916,In_1669,In_2364);
and U5917 (N_5917,In_1234,In_125);
or U5918 (N_5918,In_873,In_1378);
or U5919 (N_5919,In_386,In_1755);
nand U5920 (N_5920,In_2275,In_770);
nand U5921 (N_5921,In_964,In_665);
nand U5922 (N_5922,In_1994,In_1342);
nor U5923 (N_5923,In_364,In_1978);
nor U5924 (N_5924,In_82,In_530);
or U5925 (N_5925,In_941,In_1921);
nand U5926 (N_5926,In_1021,In_731);
and U5927 (N_5927,In_1332,In_1742);
nor U5928 (N_5928,In_2444,In_1531);
nor U5929 (N_5929,In_2077,In_1438);
nor U5930 (N_5930,In_1474,In_1469);
or U5931 (N_5931,In_151,In_1255);
or U5932 (N_5932,In_1491,In_975);
or U5933 (N_5933,In_2015,In_1835);
or U5934 (N_5934,In_590,In_1832);
or U5935 (N_5935,In_1160,In_2068);
nor U5936 (N_5936,In_867,In_688);
and U5937 (N_5937,In_965,In_24);
and U5938 (N_5938,In_609,In_221);
and U5939 (N_5939,In_1137,In_1399);
and U5940 (N_5940,In_281,In_2258);
or U5941 (N_5941,In_784,In_1454);
and U5942 (N_5942,In_1524,In_1419);
nor U5943 (N_5943,In_2321,In_590);
nor U5944 (N_5944,In_2479,In_750);
xnor U5945 (N_5945,In_2310,In_2415);
nand U5946 (N_5946,In_971,In_296);
or U5947 (N_5947,In_1975,In_645);
or U5948 (N_5948,In_1796,In_2224);
nand U5949 (N_5949,In_27,In_840);
or U5950 (N_5950,In_851,In_2370);
nor U5951 (N_5951,In_1761,In_1954);
and U5952 (N_5952,In_50,In_1718);
or U5953 (N_5953,In_1059,In_874);
nand U5954 (N_5954,In_761,In_2027);
nor U5955 (N_5955,In_504,In_2212);
or U5956 (N_5956,In_1035,In_1548);
and U5957 (N_5957,In_2154,In_16);
or U5958 (N_5958,In_1209,In_2225);
nor U5959 (N_5959,In_924,In_2496);
nor U5960 (N_5960,In_1217,In_2092);
and U5961 (N_5961,In_2312,In_1626);
or U5962 (N_5962,In_1576,In_712);
and U5963 (N_5963,In_1788,In_1204);
nand U5964 (N_5964,In_1965,In_611);
nand U5965 (N_5965,In_798,In_1452);
nand U5966 (N_5966,In_1946,In_2076);
nand U5967 (N_5967,In_673,In_142);
and U5968 (N_5968,In_660,In_1129);
and U5969 (N_5969,In_285,In_2282);
nand U5970 (N_5970,In_1451,In_479);
nand U5971 (N_5971,In_1663,In_58);
or U5972 (N_5972,In_801,In_107);
and U5973 (N_5973,In_464,In_2171);
nand U5974 (N_5974,In_1132,In_627);
or U5975 (N_5975,In_1021,In_236);
or U5976 (N_5976,In_2096,In_270);
nor U5977 (N_5977,In_1121,In_1471);
or U5978 (N_5978,In_84,In_657);
or U5979 (N_5979,In_1205,In_1661);
and U5980 (N_5980,In_420,In_245);
and U5981 (N_5981,In_1852,In_2283);
and U5982 (N_5982,In_2078,In_2011);
nand U5983 (N_5983,In_2385,In_2097);
and U5984 (N_5984,In_1450,In_1347);
nor U5985 (N_5985,In_2215,In_614);
or U5986 (N_5986,In_219,In_1305);
nand U5987 (N_5987,In_2226,In_1377);
nand U5988 (N_5988,In_1635,In_802);
nor U5989 (N_5989,In_1708,In_243);
nand U5990 (N_5990,In_1209,In_568);
xnor U5991 (N_5991,In_1000,In_2294);
and U5992 (N_5992,In_51,In_2280);
or U5993 (N_5993,In_1468,In_1376);
or U5994 (N_5994,In_1041,In_752);
and U5995 (N_5995,In_2451,In_1443);
nor U5996 (N_5996,In_1491,In_2230);
nor U5997 (N_5997,In_1887,In_202);
and U5998 (N_5998,In_1883,In_2351);
nor U5999 (N_5999,In_982,In_1814);
nor U6000 (N_6000,In_89,In_910);
or U6001 (N_6001,In_1669,In_2);
nor U6002 (N_6002,In_160,In_1493);
or U6003 (N_6003,In_2138,In_2244);
nor U6004 (N_6004,In_325,In_2290);
nor U6005 (N_6005,In_2073,In_774);
or U6006 (N_6006,In_1261,In_1424);
nand U6007 (N_6007,In_2280,In_1082);
and U6008 (N_6008,In_2353,In_949);
nand U6009 (N_6009,In_1360,In_1694);
nand U6010 (N_6010,In_1059,In_2030);
or U6011 (N_6011,In_1876,In_2126);
and U6012 (N_6012,In_524,In_1183);
and U6013 (N_6013,In_1490,In_60);
nor U6014 (N_6014,In_1828,In_738);
nor U6015 (N_6015,In_1215,In_489);
nand U6016 (N_6016,In_1829,In_1480);
nor U6017 (N_6017,In_2185,In_1146);
and U6018 (N_6018,In_1141,In_2323);
or U6019 (N_6019,In_602,In_888);
nand U6020 (N_6020,In_232,In_727);
or U6021 (N_6021,In_162,In_1697);
and U6022 (N_6022,In_512,In_78);
and U6023 (N_6023,In_339,In_2166);
and U6024 (N_6024,In_1004,In_241);
and U6025 (N_6025,In_2397,In_302);
nand U6026 (N_6026,In_1317,In_1977);
or U6027 (N_6027,In_1336,In_2349);
or U6028 (N_6028,In_1528,In_1064);
or U6029 (N_6029,In_856,In_2374);
nand U6030 (N_6030,In_539,In_2421);
nor U6031 (N_6031,In_314,In_1057);
and U6032 (N_6032,In_1060,In_2383);
or U6033 (N_6033,In_389,In_1683);
nor U6034 (N_6034,In_955,In_2359);
nor U6035 (N_6035,In_369,In_1358);
or U6036 (N_6036,In_1513,In_377);
nor U6037 (N_6037,In_1742,In_1158);
or U6038 (N_6038,In_1531,In_2058);
and U6039 (N_6039,In_478,In_790);
and U6040 (N_6040,In_200,In_2387);
or U6041 (N_6041,In_1438,In_2189);
nor U6042 (N_6042,In_1731,In_137);
xnor U6043 (N_6043,In_1538,In_1642);
or U6044 (N_6044,In_969,In_1565);
nand U6045 (N_6045,In_261,In_804);
and U6046 (N_6046,In_2290,In_901);
and U6047 (N_6047,In_2470,In_1939);
and U6048 (N_6048,In_108,In_799);
nand U6049 (N_6049,In_1929,In_1283);
or U6050 (N_6050,In_1489,In_1895);
and U6051 (N_6051,In_611,In_1282);
or U6052 (N_6052,In_752,In_1246);
or U6053 (N_6053,In_2343,In_2491);
or U6054 (N_6054,In_2494,In_108);
and U6055 (N_6055,In_1968,In_380);
nor U6056 (N_6056,In_790,In_2258);
and U6057 (N_6057,In_2217,In_542);
nand U6058 (N_6058,In_438,In_72);
nand U6059 (N_6059,In_102,In_1089);
nor U6060 (N_6060,In_1989,In_934);
nand U6061 (N_6061,In_2492,In_2202);
or U6062 (N_6062,In_1036,In_1249);
nand U6063 (N_6063,In_2190,In_1175);
or U6064 (N_6064,In_368,In_1923);
or U6065 (N_6065,In_467,In_817);
nand U6066 (N_6066,In_1638,In_1877);
nor U6067 (N_6067,In_2266,In_1084);
or U6068 (N_6068,In_164,In_1968);
and U6069 (N_6069,In_1342,In_1436);
nand U6070 (N_6070,In_682,In_2001);
or U6071 (N_6071,In_931,In_574);
nor U6072 (N_6072,In_1902,In_1303);
nor U6073 (N_6073,In_1181,In_1044);
nor U6074 (N_6074,In_2148,In_930);
nor U6075 (N_6075,In_2174,In_57);
and U6076 (N_6076,In_1459,In_1602);
nand U6077 (N_6077,In_2354,In_2349);
or U6078 (N_6078,In_151,In_1278);
or U6079 (N_6079,In_1444,In_1063);
nand U6080 (N_6080,In_928,In_101);
nand U6081 (N_6081,In_524,In_1209);
nand U6082 (N_6082,In_1672,In_1290);
or U6083 (N_6083,In_1882,In_1668);
nor U6084 (N_6084,In_982,In_1755);
or U6085 (N_6085,In_2306,In_883);
and U6086 (N_6086,In_314,In_765);
and U6087 (N_6087,In_250,In_2321);
or U6088 (N_6088,In_1825,In_1679);
and U6089 (N_6089,In_202,In_477);
and U6090 (N_6090,In_767,In_435);
nor U6091 (N_6091,In_1689,In_827);
nand U6092 (N_6092,In_1201,In_2106);
xor U6093 (N_6093,In_2345,In_328);
and U6094 (N_6094,In_1309,In_2308);
or U6095 (N_6095,In_768,In_1197);
nand U6096 (N_6096,In_1521,In_2269);
nor U6097 (N_6097,In_1786,In_520);
or U6098 (N_6098,In_2490,In_180);
or U6099 (N_6099,In_2321,In_856);
nand U6100 (N_6100,In_1108,In_1548);
nand U6101 (N_6101,In_1659,In_1156);
and U6102 (N_6102,In_2147,In_1629);
nand U6103 (N_6103,In_95,In_1838);
and U6104 (N_6104,In_2098,In_1978);
and U6105 (N_6105,In_1122,In_819);
or U6106 (N_6106,In_115,In_1037);
nand U6107 (N_6107,In_1691,In_1404);
and U6108 (N_6108,In_540,In_1167);
nand U6109 (N_6109,In_757,In_1328);
nor U6110 (N_6110,In_137,In_97);
nor U6111 (N_6111,In_2300,In_1383);
or U6112 (N_6112,In_254,In_2235);
nand U6113 (N_6113,In_1799,In_241);
nor U6114 (N_6114,In_1807,In_1262);
nand U6115 (N_6115,In_1534,In_909);
and U6116 (N_6116,In_1552,In_1967);
or U6117 (N_6117,In_309,In_2013);
and U6118 (N_6118,In_2378,In_873);
or U6119 (N_6119,In_2164,In_1892);
nor U6120 (N_6120,In_2028,In_467);
nand U6121 (N_6121,In_872,In_1882);
nand U6122 (N_6122,In_38,In_739);
nand U6123 (N_6123,In_1800,In_1303);
nor U6124 (N_6124,In_2188,In_1312);
nand U6125 (N_6125,In_2270,In_1102);
or U6126 (N_6126,In_3,In_88);
or U6127 (N_6127,In_398,In_2298);
or U6128 (N_6128,In_429,In_1497);
or U6129 (N_6129,In_1509,In_2471);
and U6130 (N_6130,In_2094,In_1854);
and U6131 (N_6131,In_165,In_2049);
nor U6132 (N_6132,In_2311,In_382);
nand U6133 (N_6133,In_1897,In_213);
nand U6134 (N_6134,In_2248,In_310);
nor U6135 (N_6135,In_520,In_1363);
nor U6136 (N_6136,In_1666,In_150);
and U6137 (N_6137,In_2120,In_982);
or U6138 (N_6138,In_933,In_1317);
or U6139 (N_6139,In_203,In_1075);
or U6140 (N_6140,In_1032,In_277);
nand U6141 (N_6141,In_280,In_1737);
nor U6142 (N_6142,In_2459,In_1156);
or U6143 (N_6143,In_1784,In_426);
or U6144 (N_6144,In_2130,In_16);
or U6145 (N_6145,In_1622,In_254);
nor U6146 (N_6146,In_1148,In_1230);
nand U6147 (N_6147,In_2423,In_1437);
or U6148 (N_6148,In_2283,In_1096);
or U6149 (N_6149,In_1027,In_571);
nor U6150 (N_6150,In_2342,In_1035);
nand U6151 (N_6151,In_13,In_1814);
and U6152 (N_6152,In_1334,In_2155);
nor U6153 (N_6153,In_2250,In_1318);
nand U6154 (N_6154,In_1095,In_2048);
nand U6155 (N_6155,In_2012,In_332);
nand U6156 (N_6156,In_1123,In_1460);
or U6157 (N_6157,In_2126,In_2372);
nand U6158 (N_6158,In_2462,In_2090);
or U6159 (N_6159,In_2028,In_439);
nor U6160 (N_6160,In_1315,In_512);
or U6161 (N_6161,In_2161,In_995);
nor U6162 (N_6162,In_894,In_1744);
and U6163 (N_6163,In_137,In_56);
and U6164 (N_6164,In_2435,In_2197);
nand U6165 (N_6165,In_801,In_1160);
nand U6166 (N_6166,In_1102,In_2020);
nor U6167 (N_6167,In_175,In_1957);
nand U6168 (N_6168,In_1652,In_1926);
nand U6169 (N_6169,In_436,In_1835);
and U6170 (N_6170,In_951,In_381);
nor U6171 (N_6171,In_705,In_1741);
or U6172 (N_6172,In_2166,In_1548);
nand U6173 (N_6173,In_2440,In_319);
nor U6174 (N_6174,In_1936,In_553);
nand U6175 (N_6175,In_218,In_1650);
nor U6176 (N_6176,In_1498,In_2346);
and U6177 (N_6177,In_1696,In_572);
and U6178 (N_6178,In_913,In_306);
nand U6179 (N_6179,In_300,In_1664);
or U6180 (N_6180,In_1599,In_719);
or U6181 (N_6181,In_1058,In_1169);
or U6182 (N_6182,In_511,In_1009);
nor U6183 (N_6183,In_902,In_1276);
nor U6184 (N_6184,In_1580,In_1836);
and U6185 (N_6185,In_367,In_1173);
and U6186 (N_6186,In_690,In_2007);
nor U6187 (N_6187,In_890,In_1290);
or U6188 (N_6188,In_2482,In_2104);
nand U6189 (N_6189,In_716,In_148);
and U6190 (N_6190,In_2226,In_688);
nand U6191 (N_6191,In_753,In_1188);
nor U6192 (N_6192,In_779,In_443);
nor U6193 (N_6193,In_906,In_1467);
nand U6194 (N_6194,In_1014,In_1095);
nand U6195 (N_6195,In_1551,In_2212);
nor U6196 (N_6196,In_1791,In_1200);
and U6197 (N_6197,In_484,In_1931);
nor U6198 (N_6198,In_514,In_839);
nor U6199 (N_6199,In_1829,In_1956);
and U6200 (N_6200,In_1772,In_1314);
nand U6201 (N_6201,In_1127,In_1490);
or U6202 (N_6202,In_1886,In_626);
or U6203 (N_6203,In_977,In_1989);
nor U6204 (N_6204,In_467,In_514);
nor U6205 (N_6205,In_2262,In_2150);
nand U6206 (N_6206,In_678,In_1526);
nand U6207 (N_6207,In_2014,In_1132);
nand U6208 (N_6208,In_967,In_1852);
and U6209 (N_6209,In_1103,In_1315);
and U6210 (N_6210,In_398,In_108);
nand U6211 (N_6211,In_134,In_1916);
nand U6212 (N_6212,In_2420,In_196);
or U6213 (N_6213,In_2149,In_1510);
nor U6214 (N_6214,In_705,In_426);
nand U6215 (N_6215,In_491,In_1221);
nor U6216 (N_6216,In_458,In_1706);
and U6217 (N_6217,In_1332,In_2437);
or U6218 (N_6218,In_2348,In_628);
nand U6219 (N_6219,In_2093,In_2106);
and U6220 (N_6220,In_1981,In_97);
and U6221 (N_6221,In_1033,In_39);
and U6222 (N_6222,In_1402,In_1316);
or U6223 (N_6223,In_2029,In_337);
nand U6224 (N_6224,In_1662,In_1041);
and U6225 (N_6225,In_1568,In_393);
or U6226 (N_6226,In_361,In_2118);
and U6227 (N_6227,In_1882,In_1560);
nor U6228 (N_6228,In_1627,In_145);
nand U6229 (N_6229,In_735,In_1915);
nand U6230 (N_6230,In_1341,In_370);
nor U6231 (N_6231,In_1327,In_2261);
nor U6232 (N_6232,In_59,In_70);
nand U6233 (N_6233,In_1378,In_2312);
nand U6234 (N_6234,In_426,In_132);
nand U6235 (N_6235,In_2302,In_1229);
nand U6236 (N_6236,In_2260,In_2359);
nand U6237 (N_6237,In_2213,In_423);
or U6238 (N_6238,In_2317,In_2105);
nand U6239 (N_6239,In_477,In_1555);
or U6240 (N_6240,In_319,In_42);
and U6241 (N_6241,In_800,In_601);
and U6242 (N_6242,In_347,In_631);
nor U6243 (N_6243,In_857,In_1552);
nand U6244 (N_6244,In_1222,In_233);
and U6245 (N_6245,In_742,In_2203);
and U6246 (N_6246,In_2280,In_1216);
xor U6247 (N_6247,In_730,In_2362);
nand U6248 (N_6248,In_1820,In_1088);
or U6249 (N_6249,In_1543,In_933);
or U6250 (N_6250,N_4218,N_3323);
nor U6251 (N_6251,N_2834,N_3108);
nand U6252 (N_6252,N_2389,N_1007);
nand U6253 (N_6253,N_1396,N_4844);
and U6254 (N_6254,N_1931,N_2383);
and U6255 (N_6255,N_4053,N_3624);
nand U6256 (N_6256,N_3876,N_5920);
and U6257 (N_6257,N_5971,N_2301);
and U6258 (N_6258,N_172,N_5727);
and U6259 (N_6259,N_2798,N_5872);
or U6260 (N_6260,N_4695,N_2329);
nor U6261 (N_6261,N_5293,N_3884);
nand U6262 (N_6262,N_449,N_5808);
nand U6263 (N_6263,N_3611,N_1034);
nor U6264 (N_6264,N_1964,N_5559);
nand U6265 (N_6265,N_4385,N_2796);
nor U6266 (N_6266,N_2658,N_5793);
or U6267 (N_6267,N_2226,N_2030);
nor U6268 (N_6268,N_5299,N_5327);
or U6269 (N_6269,N_2517,N_3093);
and U6270 (N_6270,N_4880,N_1326);
and U6271 (N_6271,N_2097,N_5387);
nor U6272 (N_6272,N_5516,N_3982);
and U6273 (N_6273,N_2403,N_1039);
and U6274 (N_6274,N_782,N_4669);
or U6275 (N_6275,N_1624,N_1162);
or U6276 (N_6276,N_2734,N_3685);
nand U6277 (N_6277,N_6088,N_1539);
nand U6278 (N_6278,N_5563,N_3182);
or U6279 (N_6279,N_5826,N_2059);
or U6280 (N_6280,N_2373,N_5152);
nand U6281 (N_6281,N_2762,N_5851);
nand U6282 (N_6282,N_4168,N_5319);
and U6283 (N_6283,N_3723,N_6206);
nor U6284 (N_6284,N_3449,N_999);
nor U6285 (N_6285,N_9,N_4322);
xnor U6286 (N_6286,N_5594,N_5999);
nor U6287 (N_6287,N_307,N_6097);
and U6288 (N_6288,N_3321,N_6177);
nand U6289 (N_6289,N_2421,N_2345);
nor U6290 (N_6290,N_4914,N_3291);
nor U6291 (N_6291,N_6182,N_4330);
nor U6292 (N_6292,N_5548,N_1156);
xor U6293 (N_6293,N_4278,N_3904);
nor U6294 (N_6294,N_5554,N_5948);
nor U6295 (N_6295,N_2575,N_3314);
nor U6296 (N_6296,N_5976,N_5970);
nand U6297 (N_6297,N_867,N_1938);
or U6298 (N_6298,N_2100,N_2662);
nor U6299 (N_6299,N_3845,N_1542);
or U6300 (N_6300,N_5310,N_2148);
nand U6301 (N_6301,N_4962,N_3622);
nor U6302 (N_6302,N_5823,N_2811);
or U6303 (N_6303,N_5663,N_4850);
nor U6304 (N_6304,N_982,N_1402);
nand U6305 (N_6305,N_5553,N_5778);
nand U6306 (N_6306,N_1531,N_1325);
nor U6307 (N_6307,N_5517,N_5480);
and U6308 (N_6308,N_5814,N_3236);
or U6309 (N_6309,N_1709,N_3041);
and U6310 (N_6310,N_448,N_2844);
or U6311 (N_6311,N_1585,N_1018);
nand U6312 (N_6312,N_1522,N_4743);
and U6313 (N_6313,N_5816,N_5998);
nor U6314 (N_6314,N_3172,N_4380);
and U6315 (N_6315,N_2807,N_3947);
and U6316 (N_6316,N_3202,N_5586);
or U6317 (N_6317,N_6222,N_4956);
nor U6318 (N_6318,N_1313,N_5499);
nor U6319 (N_6319,N_743,N_1098);
or U6320 (N_6320,N_2230,N_27);
and U6321 (N_6321,N_5994,N_3950);
nand U6322 (N_6322,N_5323,N_2559);
nand U6323 (N_6323,N_4276,N_3647);
nand U6324 (N_6324,N_334,N_3765);
or U6325 (N_6325,N_3692,N_1715);
nand U6326 (N_6326,N_2615,N_4697);
and U6327 (N_6327,N_4555,N_4199);
and U6328 (N_6328,N_1817,N_3697);
or U6329 (N_6329,N_200,N_4547);
nor U6330 (N_6330,N_868,N_2194);
or U6331 (N_6331,N_2262,N_5267);
nor U6332 (N_6332,N_5446,N_3453);
or U6333 (N_6333,N_5643,N_14);
nor U6334 (N_6334,N_996,N_3122);
or U6335 (N_6335,N_5588,N_1637);
or U6336 (N_6336,N_5218,N_238);
and U6337 (N_6337,N_4833,N_3059);
nand U6338 (N_6338,N_4519,N_5185);
nor U6339 (N_6339,N_3082,N_2471);
nor U6340 (N_6340,N_4560,N_6046);
and U6341 (N_6341,N_3981,N_2268);
nand U6342 (N_6342,N_1633,N_375);
nand U6343 (N_6343,N_3926,N_1602);
nor U6344 (N_6344,N_2554,N_3288);
and U6345 (N_6345,N_468,N_5658);
nor U6346 (N_6346,N_1381,N_4858);
nor U6347 (N_6347,N_1775,N_265);
and U6348 (N_6348,N_544,N_2987);
nor U6349 (N_6349,N_2646,N_1353);
or U6350 (N_6350,N_3251,N_3356);
nand U6351 (N_6351,N_6116,N_6141);
or U6352 (N_6352,N_2155,N_658);
nand U6353 (N_6353,N_4421,N_4122);
nor U6354 (N_6354,N_3392,N_4101);
and U6355 (N_6355,N_695,N_3777);
or U6356 (N_6356,N_5785,N_3631);
nor U6357 (N_6357,N_6194,N_5278);
nor U6358 (N_6358,N_4965,N_3580);
nor U6359 (N_6359,N_2368,N_2069);
nor U6360 (N_6360,N_5191,N_3381);
nor U6361 (N_6361,N_1631,N_1195);
nand U6362 (N_6362,N_3022,N_2772);
and U6363 (N_6363,N_4653,N_1414);
nand U6364 (N_6364,N_342,N_1880);
and U6365 (N_6365,N_2152,N_2033);
nand U6366 (N_6366,N_5346,N_5059);
nor U6367 (N_6367,N_3407,N_2758);
nor U6368 (N_6368,N_2854,N_5037);
or U6369 (N_6369,N_225,N_5507);
or U6370 (N_6370,N_902,N_133);
and U6371 (N_6371,N_450,N_2723);
and U6372 (N_6372,N_5277,N_5635);
nor U6373 (N_6373,N_5639,N_5725);
or U6374 (N_6374,N_6060,N_4698);
nand U6375 (N_6375,N_675,N_3858);
and U6376 (N_6376,N_3881,N_3357);
and U6377 (N_6377,N_4347,N_4207);
nor U6378 (N_6378,N_5492,N_4500);
or U6379 (N_6379,N_1655,N_6054);
nor U6380 (N_6380,N_2044,N_1661);
or U6381 (N_6381,N_6139,N_894);
nand U6382 (N_6382,N_3762,N_2296);
nor U6383 (N_6383,N_2034,N_5271);
nand U6384 (N_6384,N_5128,N_1696);
nand U6385 (N_6385,N_1209,N_571);
nor U6386 (N_6386,N_5961,N_5836);
or U6387 (N_6387,N_2372,N_2073);
and U6388 (N_6388,N_2998,N_929);
and U6389 (N_6389,N_318,N_3015);
and U6390 (N_6390,N_5339,N_1223);
nand U6391 (N_6391,N_1406,N_4942);
nor U6392 (N_6392,N_232,N_5662);
nor U6393 (N_6393,N_5476,N_1985);
or U6394 (N_6394,N_4245,N_3044);
and U6395 (N_6395,N_4447,N_5767);
nor U6396 (N_6396,N_4982,N_3485);
and U6397 (N_6397,N_528,N_2452);
nor U6398 (N_6398,N_5382,N_6134);
or U6399 (N_6399,N_3042,N_6100);
nand U6400 (N_6400,N_3009,N_1060);
and U6401 (N_6401,N_5459,N_5703);
nor U6402 (N_6402,N_2691,N_4883);
or U6403 (N_6403,N_2271,N_5627);
and U6404 (N_6404,N_3364,N_1541);
or U6405 (N_6405,N_5822,N_1606);
or U6406 (N_6406,N_2178,N_1788);
and U6407 (N_6407,N_1095,N_2254);
nor U6408 (N_6408,N_2355,N_274);
or U6409 (N_6409,N_4353,N_4938);
or U6410 (N_6410,N_5952,N_3584);
nor U6411 (N_6411,N_3717,N_5743);
or U6412 (N_6412,N_1456,N_2320);
or U6413 (N_6413,N_2989,N_3161);
nor U6414 (N_6414,N_1348,N_1844);
nor U6415 (N_6415,N_2509,N_2241);
nor U6416 (N_6416,N_5804,N_4992);
nor U6417 (N_6417,N_543,N_3703);
or U6418 (N_6418,N_5463,N_4180);
or U6419 (N_6419,N_5728,N_3706);
or U6420 (N_6420,N_1021,N_5049);
nor U6421 (N_6421,N_1062,N_2123);
and U6422 (N_6422,N_5631,N_1306);
nor U6423 (N_6423,N_2134,N_4201);
nand U6424 (N_6424,N_331,N_5646);
or U6425 (N_6425,N_2225,N_2205);
and U6426 (N_6426,N_3800,N_4445);
and U6427 (N_6427,N_6219,N_1438);
or U6428 (N_6428,N_874,N_5033);
nor U6429 (N_6429,N_5081,N_3940);
nand U6430 (N_6430,N_3260,N_4510);
or U6431 (N_6431,N_953,N_4798);
nand U6432 (N_6432,N_42,N_3462);
nor U6433 (N_6433,N_2050,N_4782);
and U6434 (N_6434,N_3416,N_1304);
or U6435 (N_6435,N_147,N_4220);
or U6436 (N_6436,N_3132,N_4606);
nand U6437 (N_6437,N_179,N_1070);
nor U6438 (N_6438,N_3229,N_3514);
or U6439 (N_6439,N_1442,N_4910);
nand U6440 (N_6440,N_4487,N_5958);
nor U6441 (N_6441,N_5163,N_1989);
nor U6442 (N_6442,N_3919,N_3867);
and U6443 (N_6443,N_437,N_2188);
and U6444 (N_6444,N_1214,N_1427);
nor U6445 (N_6445,N_1285,N_5250);
or U6446 (N_6446,N_3851,N_305);
and U6447 (N_6447,N_4726,N_236);
and U6448 (N_6448,N_5711,N_5526);
or U6449 (N_6449,N_5556,N_4328);
and U6450 (N_6450,N_2548,N_5605);
nand U6451 (N_6451,N_5352,N_4932);
and U6452 (N_6452,N_1305,N_5599);
or U6453 (N_6453,N_5745,N_5504);
and U6454 (N_6454,N_2853,N_832);
and U6455 (N_6455,N_1084,N_5018);
and U6456 (N_6456,N_1261,N_253);
nor U6457 (N_6457,N_3801,N_688);
and U6458 (N_6458,N_3724,N_1568);
nor U6459 (N_6459,N_525,N_6136);
nand U6460 (N_6460,N_178,N_650);
nor U6461 (N_6461,N_3659,N_2640);
or U6462 (N_6462,N_2207,N_3595);
nand U6463 (N_6463,N_1771,N_921);
nand U6464 (N_6464,N_5869,N_1733);
and U6465 (N_6465,N_1872,N_1660);
nand U6466 (N_6466,N_401,N_3597);
and U6467 (N_6467,N_4008,N_1913);
nor U6468 (N_6468,N_3903,N_2163);
or U6469 (N_6469,N_488,N_3586);
xnor U6470 (N_6470,N_3277,N_2478);
xnor U6471 (N_6471,N_992,N_3225);
or U6472 (N_6472,N_2896,N_106);
nand U6473 (N_6473,N_5094,N_1051);
or U6474 (N_6474,N_4652,N_154);
nand U6475 (N_6475,N_128,N_5210);
nand U6476 (N_6476,N_1740,N_1806);
nand U6477 (N_6477,N_257,N_4279);
nor U6478 (N_6478,N_1623,N_5207);
nor U6479 (N_6479,N_4724,N_5540);
nor U6480 (N_6480,N_3520,N_5722);
or U6481 (N_6481,N_2359,N_2788);
and U6482 (N_6482,N_1867,N_3193);
nand U6483 (N_6483,N_6105,N_432);
and U6484 (N_6484,N_5256,N_4955);
or U6485 (N_6485,N_1178,N_2009);
nand U6486 (N_6486,N_2906,N_3694);
xor U6487 (N_6487,N_5455,N_2287);
nor U6488 (N_6488,N_1901,N_1134);
or U6489 (N_6489,N_1268,N_1682);
or U6490 (N_6490,N_5176,N_5305);
and U6491 (N_6491,N_308,N_4513);
nand U6492 (N_6492,N_1701,N_804);
nor U6493 (N_6493,N_201,N_2008);
or U6494 (N_6494,N_5544,N_4419);
or U6495 (N_6495,N_730,N_4195);
and U6496 (N_6496,N_3306,N_1450);
nor U6497 (N_6497,N_2130,N_3319);
nor U6498 (N_6498,N_2810,N_5717);
and U6499 (N_6499,N_2838,N_1433);
nand U6500 (N_6500,N_692,N_1575);
or U6501 (N_6501,N_430,N_4535);
and U6502 (N_6502,N_5086,N_4277);
nor U6503 (N_6503,N_3083,N_2196);
and U6504 (N_6504,N_5098,N_3821);
and U6505 (N_6505,N_881,N_242);
nand U6506 (N_6506,N_823,N_1934);
nor U6507 (N_6507,N_4649,N_3722);
or U6508 (N_6508,N_1215,N_3571);
nand U6509 (N_6509,N_948,N_4538);
and U6510 (N_6510,N_4639,N_6085);
nor U6511 (N_6511,N_4356,N_3949);
and U6512 (N_6512,N_674,N_5226);
nand U6513 (N_6513,N_4524,N_434);
nor U6514 (N_6514,N_2154,N_11);
nor U6515 (N_6515,N_2956,N_1453);
nand U6516 (N_6516,N_4552,N_4483);
nand U6517 (N_6517,N_358,N_2036);
and U6518 (N_6518,N_3938,N_4988);
or U6519 (N_6519,N_1672,N_3602);
nand U6520 (N_6520,N_2971,N_5854);
nand U6521 (N_6521,N_1663,N_6211);
or U6522 (N_6522,N_5263,N_3741);
nor U6523 (N_6523,N_2719,N_1289);
nor U6524 (N_6524,N_1122,N_2292);
and U6525 (N_6525,N_4661,N_3387);
nand U6526 (N_6526,N_535,N_3523);
nand U6527 (N_6527,N_3578,N_4216);
and U6528 (N_6528,N_2480,N_1286);
nand U6529 (N_6529,N_296,N_5852);
or U6530 (N_6530,N_4332,N_3328);
or U6531 (N_6531,N_1206,N_3822);
or U6532 (N_6532,N_4898,N_1811);
nand U6533 (N_6533,N_4464,N_5150);
or U6534 (N_6534,N_3458,N_585);
and U6535 (N_6535,N_4198,N_5577);
nor U6536 (N_6536,N_187,N_357);
or U6537 (N_6537,N_327,N_1890);
nor U6538 (N_6538,N_2157,N_2941);
nand U6539 (N_6539,N_1249,N_1630);
nor U6540 (N_6540,N_5671,N_2282);
nor U6541 (N_6541,N_1327,N_3660);
nand U6542 (N_6542,N_50,N_6074);
nand U6543 (N_6543,N_3493,N_2416);
and U6544 (N_6544,N_1093,N_5502);
nand U6545 (N_6545,N_5413,N_1503);
nor U6546 (N_6546,N_2905,N_5932);
or U6547 (N_6547,N_1421,N_5221);
nor U6548 (N_6548,N_5261,N_5887);
and U6549 (N_6549,N_104,N_1257);
or U6550 (N_6550,N_1293,N_1557);
nor U6551 (N_6551,N_4469,N_3826);
nand U6552 (N_6552,N_1997,N_4739);
nand U6553 (N_6553,N_6243,N_2922);
or U6554 (N_6554,N_3080,N_3231);
or U6555 (N_6555,N_5070,N_5759);
nand U6556 (N_6556,N_1654,N_6247);
nand U6557 (N_6557,N_3859,N_1431);
and U6558 (N_6558,N_4542,N_676);
nor U6559 (N_6559,N_4571,N_5147);
or U6560 (N_6560,N_2555,N_1573);
or U6561 (N_6561,N_3307,N_566);
nor U6562 (N_6562,N_4505,N_1762);
and U6563 (N_6563,N_1213,N_2032);
nor U6564 (N_6564,N_977,N_6173);
or U6565 (N_6565,N_2609,N_5290);
or U6566 (N_6566,N_4246,N_5223);
nor U6567 (N_6567,N_1896,N_1594);
and U6568 (N_6568,N_5716,N_5036);
or U6569 (N_6569,N_1618,N_2293);
and U6570 (N_6570,N_3284,N_5988);
and U6571 (N_6571,N_1296,N_3233);
and U6572 (N_6572,N_1782,N_5460);
nand U6573 (N_6573,N_4359,N_4770);
and U6574 (N_6574,N_3969,N_4736);
nor U6575 (N_6575,N_1727,N_943);
nor U6576 (N_6576,N_109,N_3921);
or U6577 (N_6577,N_5704,N_114);
nand U6578 (N_6578,N_4372,N_947);
and U6579 (N_6579,N_5164,N_2654);
nor U6580 (N_6580,N_1831,N_1509);
or U6581 (N_6581,N_3145,N_3341);
and U6582 (N_6582,N_2051,N_210);
and U6583 (N_6583,N_6032,N_828);
or U6584 (N_6584,N_6113,N_2305);
or U6585 (N_6585,N_3179,N_3585);
or U6586 (N_6586,N_1322,N_3376);
nor U6587 (N_6587,N_4074,N_498);
nor U6588 (N_6588,N_1780,N_2197);
xor U6589 (N_6589,N_5350,N_1040);
nand U6590 (N_6590,N_5888,N_5736);
nand U6591 (N_6591,N_5571,N_2346);
xnor U6592 (N_6592,N_2603,N_2012);
nand U6593 (N_6593,N_5394,N_5418);
or U6594 (N_6594,N_2622,N_417);
or U6595 (N_6595,N_5072,N_5535);
or U6596 (N_6596,N_1377,N_813);
nand U6597 (N_6597,N_839,N_2379);
xor U6598 (N_6598,N_4397,N_3442);
and U6599 (N_6599,N_6019,N_5927);
and U6600 (N_6600,N_5737,N_6089);
nand U6601 (N_6601,N_624,N_4105);
or U6602 (N_6602,N_5938,N_3345);
and U6603 (N_6603,N_486,N_4699);
and U6604 (N_6604,N_1128,N_1083);
xnor U6605 (N_6605,N_875,N_4536);
or U6606 (N_6606,N_514,N_4738);
nand U6607 (N_6607,N_5963,N_1031);
nor U6608 (N_6608,N_49,N_1358);
nor U6609 (N_6609,N_4455,N_3983);
and U6610 (N_6610,N_3004,N_297);
nor U6611 (N_6611,N_2335,N_4232);
nor U6612 (N_6612,N_5587,N_272);
and U6613 (N_6613,N_3922,N_1187);
nand U6614 (N_6614,N_2897,N_5216);
nor U6615 (N_6615,N_279,N_887);
nor U6616 (N_6616,N_1620,N_1076);
nand U6617 (N_6617,N_5537,N_3238);
nand U6618 (N_6618,N_3355,N_945);
nand U6619 (N_6619,N_726,N_3732);
or U6620 (N_6620,N_6022,N_4874);
or U6621 (N_6621,N_910,N_1800);
nand U6622 (N_6622,N_245,N_6104);
and U6623 (N_6623,N_3184,N_4553);
and U6624 (N_6624,N_5832,N_6012);
and U6625 (N_6625,N_5124,N_2146);
nand U6626 (N_6626,N_5075,N_4048);
nand U6627 (N_6627,N_5016,N_5032);
and U6628 (N_6628,N_4377,N_4757);
or U6629 (N_6629,N_1336,N_3255);
and U6630 (N_6630,N_2106,N_4530);
or U6631 (N_6631,N_2806,N_226);
nand U6632 (N_6632,N_6122,N_4435);
or U6633 (N_6633,N_4060,N_5817);
or U6634 (N_6634,N_472,N_1192);
nor U6635 (N_6635,N_2975,N_2718);
nand U6636 (N_6636,N_2092,N_686);
or U6637 (N_6637,N_555,N_5435);
nand U6638 (N_6638,N_4482,N_6198);
or U6639 (N_6639,N_1949,N_5043);
and U6640 (N_6640,N_946,N_2898);
nor U6641 (N_6641,N_84,N_1004);
nand U6642 (N_6642,N_1046,N_481);
and U6643 (N_6643,N_2516,N_5469);
nor U6644 (N_6644,N_3467,N_1491);
nor U6645 (N_6645,N_4009,N_4769);
nand U6646 (N_6646,N_2664,N_5108);
or U6647 (N_6647,N_4637,N_1383);
or U6648 (N_6648,N_2692,N_408);
or U6649 (N_6649,N_2821,N_1743);
nand U6650 (N_6650,N_164,N_4226);
and U6651 (N_6651,N_4342,N_4428);
or U6652 (N_6652,N_2782,N_4273);
nor U6653 (N_6653,N_4974,N_633);
or U6654 (N_6654,N_6207,N_4793);
nand U6655 (N_6655,N_812,N_2514);
nor U6656 (N_6656,N_4717,N_182);
xor U6657 (N_6657,N_1382,N_1691);
or U6658 (N_6658,N_5083,N_3740);
nor U6659 (N_6659,N_4759,N_1244);
nor U6660 (N_6660,N_3473,N_3437);
nor U6661 (N_6661,N_3001,N_5084);
and U6662 (N_6662,N_1842,N_4696);
and U6663 (N_6663,N_1881,N_4734);
or U6664 (N_6664,N_4977,N_5845);
nand U6665 (N_6665,N_6015,N_994);
nor U6666 (N_6666,N_678,N_1921);
or U6667 (N_6667,N_3099,N_4900);
and U6668 (N_6668,N_5104,N_2611);
or U6669 (N_6669,N_745,N_2162);
nand U6670 (N_6670,N_351,N_5294);
and U6671 (N_6671,N_203,N_5570);
or U6672 (N_6672,N_1042,N_1317);
and U6673 (N_6673,N_2563,N_3218);
or U6674 (N_6674,N_5565,N_3394);
nand U6675 (N_6675,N_2535,N_313);
and U6676 (N_6676,N_4233,N_2974);
and U6677 (N_6677,N_5316,N_1479);
nand U6678 (N_6678,N_1115,N_3113);
nand U6679 (N_6679,N_2023,N_1189);
or U6680 (N_6680,N_3930,N_340);
nand U6681 (N_6681,N_362,N_4083);
or U6682 (N_6682,N_3297,N_549);
and U6683 (N_6683,N_299,N_3071);
nor U6684 (N_6684,N_4102,N_1833);
nand U6685 (N_6685,N_1930,N_1254);
or U6686 (N_6686,N_4203,N_4237);
nand U6687 (N_6687,N_2647,N_666);
nand U6688 (N_6688,N_1555,N_5986);
nand U6689 (N_6689,N_1,N_3154);
or U6690 (N_6690,N_2445,N_3490);
and U6691 (N_6691,N_2417,N_6135);
nor U6692 (N_6692,N_625,N_5886);
xor U6693 (N_6693,N_3978,N_3727);
nand U6694 (N_6694,N_2295,N_4271);
nand U6695 (N_6695,N_1235,N_4680);
nand U6696 (N_6696,N_3016,N_1439);
and U6697 (N_6697,N_5088,N_2767);
nor U6698 (N_6698,N_1357,N_2936);
nand U6699 (N_6699,N_2915,N_5109);
nor U6700 (N_6700,N_4033,N_1403);
or U6701 (N_6701,N_6158,N_998);
nand U6702 (N_6702,N_4887,N_1461);
xor U6703 (N_6703,N_614,N_3305);
and U6704 (N_6704,N_909,N_6205);
and U6705 (N_6705,N_1173,N_87);
and U6706 (N_6706,N_5876,N_5205);
and U6707 (N_6707,N_970,N_3395);
nand U6708 (N_6708,N_1126,N_3543);
nor U6709 (N_6709,N_188,N_91);
nor U6710 (N_6710,N_1702,N_4248);
nand U6711 (N_6711,N_151,N_1832);
nand U6712 (N_6712,N_775,N_2735);
nand U6713 (N_6713,N_1599,N_1664);
nand U6714 (N_6714,N_3857,N_905);
nor U6715 (N_6715,N_4158,N_5390);
nor U6716 (N_6716,N_2642,N_3948);
or U6717 (N_6717,N_3100,N_1725);
or U6718 (N_6718,N_112,N_5698);
xnor U6719 (N_6719,N_4622,N_316);
nor U6720 (N_6720,N_2102,N_2601);
or U6721 (N_6721,N_2730,N_328);
nor U6722 (N_6722,N_3003,N_3530);
and U6723 (N_6723,N_1879,N_1246);
nand U6724 (N_6724,N_6244,N_3961);
and U6725 (N_6725,N_5053,N_1596);
nand U6726 (N_6726,N_3928,N_4566);
xnor U6727 (N_6727,N_696,N_5863);
nand U6728 (N_6728,N_427,N_556);
nor U6729 (N_6729,N_3695,N_1125);
and U6730 (N_6730,N_4103,N_1245);
nand U6731 (N_6731,N_2945,N_2376);
and U6732 (N_6732,N_1129,N_4864);
nor U6733 (N_6733,N_3564,N_345);
and U6734 (N_6734,N_4523,N_3953);
and U6735 (N_6735,N_931,N_840);
nand U6736 (N_6736,N_4412,N_1375);
nor U6737 (N_6737,N_2749,N_2840);
and U6738 (N_6738,N_1634,N_78);
nor U6739 (N_6739,N_2337,N_4877);
or U6740 (N_6740,N_2229,N_5091);
nor U6741 (N_6741,N_1429,N_3511);
nor U6742 (N_6742,N_2583,N_2619);
nor U6743 (N_6743,N_2006,N_2536);
and U6744 (N_6744,N_2704,N_3866);
and U6745 (N_6745,N_3337,N_1861);
or U6746 (N_6746,N_3373,N_2712);
and U6747 (N_6747,N_2088,N_4768);
nand U6748 (N_6748,N_2506,N_4749);
nor U6749 (N_6749,N_5980,N_2473);
or U6750 (N_6750,N_3552,N_3986);
and U6751 (N_6751,N_2540,N_5905);
and U6752 (N_6752,N_255,N_5771);
nor U6753 (N_6753,N_2700,N_4299);
nor U6754 (N_6754,N_2022,N_3272);
nor U6755 (N_6755,N_321,N_231);
nor U6756 (N_6756,N_3211,N_6169);
or U6757 (N_6757,N_3217,N_5297);
or U6758 (N_6758,N_776,N_2940);
nor U6759 (N_6759,N_5539,N_5031);
or U6760 (N_6760,N_3128,N_1790);
or U6761 (N_6761,N_606,N_3436);
or U6762 (N_6762,N_4410,N_6131);
and U6763 (N_6763,N_2994,N_1563);
and U6764 (N_6764,N_2025,N_4230);
or U6765 (N_6765,N_3827,N_1053);
and U6766 (N_6766,N_3555,N_1311);
nor U6767 (N_6767,N_615,N_1174);
nand U6768 (N_6768,N_2641,N_2191);
or U6769 (N_6769,N_1678,N_5828);
and U6770 (N_6770,N_5601,N_3457);
and U6771 (N_6771,N_4559,N_3572);
nand U6772 (N_6772,N_2387,N_3936);
nor U6773 (N_6773,N_3208,N_2751);
nor U6774 (N_6774,N_288,N_1742);
or U6775 (N_6775,N_303,N_35);
nor U6776 (N_6776,N_1294,N_3501);
nand U6777 (N_6777,N_361,N_4466);
nor U6778 (N_6778,N_1907,N_4805);
and U6779 (N_6779,N_5006,N_1443);
and U6780 (N_6780,N_5111,N_4859);
and U6781 (N_6781,N_2895,N_1615);
or U6782 (N_6782,N_2110,N_1873);
nand U6783 (N_6783,N_4133,N_5925);
or U6784 (N_6784,N_191,N_5821);
xnor U6785 (N_6785,N_5200,N_2482);
nand U6786 (N_6786,N_256,N_1205);
or U6787 (N_6787,N_4106,N_661);
nand U6788 (N_6788,N_3576,N_6175);
nor U6789 (N_6789,N_691,N_2978);
nand U6790 (N_6790,N_2572,N_1781);
and U6791 (N_6791,N_2781,N_1912);
and U6792 (N_6792,N_1412,N_4119);
nand U6793 (N_6793,N_2189,N_2489);
nand U6794 (N_6794,N_3808,N_17);
nand U6795 (N_6795,N_4702,N_3201);
or U6796 (N_6796,N_1066,N_3589);
or U6797 (N_6797,N_3508,N_5733);
nand U6798 (N_6798,N_4934,N_3744);
nand U6799 (N_6799,N_4865,N_215);
and U6800 (N_6800,N_4068,N_4826);
or U6801 (N_6801,N_1036,N_2809);
nand U6802 (N_6802,N_2632,N_347);
nand U6803 (N_6803,N_310,N_4704);
or U6804 (N_6804,N_281,N_1006);
nor U6805 (N_6805,N_6045,N_5738);
nor U6806 (N_6806,N_1809,N_944);
or U6807 (N_6807,N_2602,N_2068);
nor U6808 (N_6808,N_5426,N_5842);
nand U6809 (N_6809,N_986,N_5061);
or U6810 (N_6810,N_234,N_2374);
nand U6811 (N_6811,N_2424,N_3220);
or U6812 (N_6812,N_5583,N_5353);
nand U6813 (N_6813,N_3036,N_30);
nor U6814 (N_6814,N_1180,N_1892);
nand U6815 (N_6815,N_2494,N_2900);
nor U6816 (N_6816,N_3792,N_4894);
or U6817 (N_6817,N_588,N_3518);
nor U6818 (N_6818,N_1807,N_5213);
nand U6819 (N_6819,N_409,N_5937);
nand U6820 (N_6820,N_1511,N_1299);
nor U6821 (N_6821,N_3065,N_460);
nand U6822 (N_6822,N_2057,N_2316);
nor U6823 (N_6823,N_471,N_2881);
nand U6824 (N_6824,N_2046,N_1218);
and U6825 (N_6825,N_402,N_1320);
or U6826 (N_6826,N_1392,N_2860);
nor U6827 (N_6827,N_2760,N_2669);
and U6828 (N_6828,N_1825,N_3556);
nor U6829 (N_6829,N_3619,N_6001);
nand U6830 (N_6830,N_1864,N_230);
or U6831 (N_6831,N_1621,N_5198);
nor U6832 (N_6832,N_3750,N_4902);
and U6833 (N_6833,N_4929,N_895);
nor U6834 (N_6834,N_3682,N_2541);
nand U6835 (N_6835,N_1155,N_732);
nand U6836 (N_6836,N_6249,N_2174);
nor U6837 (N_6837,N_1272,N_3283);
and U6838 (N_6838,N_3696,N_2929);
or U6839 (N_6839,N_4417,N_5028);
and U6840 (N_6840,N_2832,N_1356);
and U6841 (N_6841,N_1333,N_810);
nor U6842 (N_6842,N_4374,N_239);
and U6843 (N_6843,N_1203,N_4791);
nand U6844 (N_6844,N_3868,N_1560);
nor U6845 (N_6845,N_4022,N_3945);
nor U6846 (N_6846,N_3326,N_1543);
nand U6847 (N_6847,N_3796,N_4247);
nand U6848 (N_6848,N_3609,N_3365);
nand U6849 (N_6849,N_3242,N_2120);
nand U6850 (N_6850,N_3087,N_2070);
nor U6851 (N_6851,N_3806,N_6049);
or U6852 (N_6852,N_34,N_1351);
nand U6853 (N_6853,N_5580,N_405);
or U6854 (N_6854,N_2284,N_893);
or U6855 (N_6855,N_3106,N_6014);
or U6856 (N_6856,N_1789,N_3850);
and U6857 (N_6857,N_1891,N_3925);
and U6858 (N_6858,N_2290,N_859);
or U6859 (N_6859,N_1865,N_3397);
or U6860 (N_6860,N_1965,N_3130);
nor U6861 (N_6861,N_6165,N_2436);
and U6862 (N_6862,N_618,N_4870);
nand U6863 (N_6863,N_4645,N_487);
and U6864 (N_6864,N_2122,N_3495);
or U6865 (N_6865,N_4191,N_3751);
and U6866 (N_6866,N_4855,N_273);
nand U6867 (N_6867,N_2682,N_2438);
nor U6868 (N_6868,N_3124,N_184);
nor U6869 (N_6869,N_5555,N_1410);
nand U6870 (N_6870,N_3270,N_2495);
and U6871 (N_6871,N_5419,N_1119);
nand U6872 (N_6872,N_5853,N_491);
nor U6873 (N_6873,N_1883,N_3683);
or U6874 (N_6874,N_797,N_5997);
nor U6875 (N_6875,N_6057,N_136);
and U6876 (N_6876,N_2397,N_356);
nand U6877 (N_6877,N_4046,N_800);
nand U6878 (N_6878,N_2361,N_1698);
nand U6879 (N_6879,N_4011,N_4042);
and U6880 (N_6880,N_6009,N_1855);
nor U6881 (N_6881,N_4183,N_4650);
and U6882 (N_6882,N_1255,N_3795);
and U6883 (N_6883,N_1980,N_1339);
nor U6884 (N_6884,N_3303,N_5969);
and U6885 (N_6885,N_2098,N_134);
and U6886 (N_6886,N_1700,N_287);
nor U6887 (N_6887,N_4707,N_721);
or U6888 (N_6888,N_5772,N_395);
and U6889 (N_6889,N_5442,N_2054);
or U6890 (N_6890,N_1387,N_3327);
nor U6891 (N_6891,N_5103,N_3869);
nand U6892 (N_6892,N_3588,N_5051);
and U6893 (N_6893,N_3880,N_1230);
nand U6894 (N_6894,N_906,N_1489);
nand U6895 (N_6895,N_4326,N_5951);
or U6896 (N_6896,N_1520,N_6098);
and U6897 (N_6897,N_5073,N_3883);
and U6898 (N_6898,N_3011,N_4722);
or U6899 (N_6899,N_3568,N_3803);
and U6900 (N_6900,N_397,N_1280);
nand U6901 (N_6901,N_596,N_4169);
or U6902 (N_6902,N_1735,N_5186);
nand U6903 (N_6903,N_926,N_4387);
nor U6904 (N_6904,N_3417,N_5292);
nor U6905 (N_6905,N_5069,N_152);
nand U6906 (N_6906,N_4358,N_5742);
or U6907 (N_6907,N_2441,N_3206);
nor U6908 (N_6908,N_783,N_3246);
or U6909 (N_6909,N_3066,N_3549);
nand U6910 (N_6910,N_3424,N_3749);
xnor U6911 (N_6911,N_1184,N_1454);
nor U6912 (N_6912,N_3415,N_4597);
nand U6913 (N_6913,N_3012,N_2385);
and U6914 (N_6914,N_5973,N_4178);
nand U6915 (N_6915,N_2366,N_3053);
and U6916 (N_6916,N_5159,N_4537);
nor U6917 (N_6917,N_2133,N_3931);
or U6918 (N_6918,N_1355,N_563);
or U6919 (N_6919,N_6156,N_2710);
nor U6920 (N_6920,N_2223,N_6225);
nor U6921 (N_6921,N_1028,N_1474);
or U6922 (N_6922,N_5253,N_5365);
nand U6923 (N_6923,N_4922,N_5640);
and U6924 (N_6924,N_668,N_3715);
or U6925 (N_6925,N_5945,N_2726);
or U6926 (N_6926,N_5357,N_251);
xnor U6927 (N_6927,N_6008,N_876);
nor U6928 (N_6928,N_866,N_4809);
nor U6929 (N_6929,N_4710,N_4893);
and U6930 (N_6930,N_4100,N_2294);
and U6931 (N_6931,N_5114,N_1995);
nand U6932 (N_6932,N_4755,N_2841);
nor U6933 (N_6933,N_4810,N_2515);
nor U6934 (N_6934,N_1619,N_559);
and U6935 (N_6935,N_5399,N_6061);
and U6936 (N_6936,N_4061,N_2737);
nand U6937 (N_6937,N_1199,N_4655);
nor U6938 (N_6938,N_3638,N_4713);
and U6939 (N_6939,N_3092,N_4351);
nor U6940 (N_6940,N_1274,N_2880);
or U6941 (N_6941,N_4150,N_3738);
or U6942 (N_6942,N_1547,N_904);
and U6943 (N_6943,N_4983,N_419);
and U6944 (N_6944,N_2577,N_1011);
or U6945 (N_6945,N_6148,N_725);
nand U6946 (N_6946,N_4824,N_2454);
nand U6947 (N_6947,N_2423,N_2890);
nand U6948 (N_6948,N_2866,N_214);
and U6949 (N_6949,N_264,N_3384);
nor U6950 (N_6950,N_5783,N_312);
and U6951 (N_6951,N_922,N_3658);
or U6952 (N_6952,N_1653,N_5622);
and U6953 (N_6953,N_4413,N_5899);
and U6954 (N_6954,N_1273,N_4352);
and U6955 (N_6955,N_282,N_1281);
nor U6956 (N_6956,N_539,N_2910);
or U6957 (N_6957,N_5187,N_4234);
nor U6958 (N_6958,N_3125,N_5762);
and U6959 (N_6959,N_2265,N_1221);
nand U6960 (N_6960,N_4803,N_6228);
and U6961 (N_6961,N_1805,N_3725);
nand U6962 (N_6962,N_1549,N_2285);
or U6963 (N_6963,N_3652,N_4853);
or U6964 (N_6964,N_2972,N_3854);
or U6965 (N_6965,N_2396,N_143);
nor U6966 (N_6966,N_5231,N_4525);
nand U6967 (N_6967,N_928,N_5782);
nand U6968 (N_6968,N_3052,N_2743);
nand U6969 (N_6969,N_741,N_5288);
nor U6970 (N_6970,N_137,N_560);
or U6971 (N_6971,N_3654,N_3714);
and U6972 (N_6972,N_2886,N_1588);
and U6973 (N_6973,N_1001,N_4039);
nand U6974 (N_6974,N_2638,N_1761);
nand U6975 (N_6975,N_458,N_2139);
and U6976 (N_6976,N_3816,N_3933);
nand U6977 (N_6977,N_2644,N_1676);
or U6978 (N_6978,N_4527,N_118);
nand U6979 (N_6979,N_1535,N_5282);
nor U6980 (N_6980,N_1407,N_5792);
nand U6981 (N_6981,N_1561,N_2339);
or U6982 (N_6982,N_1567,N_2943);
and U6983 (N_6983,N_1813,N_1829);
and U6984 (N_6984,N_3718,N_5598);
nor U6985 (N_6985,N_5510,N_3655);
nand U6986 (N_6986,N_598,N_3002);
or U6987 (N_6987,N_2942,N_2356);
nor U6988 (N_6988,N_4467,N_5438);
xnor U6989 (N_6989,N_3275,N_5653);
and U6990 (N_6990,N_5274,N_3174);
nand U6991 (N_6991,N_5251,N_5017);
nand U6992 (N_6992,N_2117,N_3705);
nand U6993 (N_6993,N_4862,N_5153);
or U6994 (N_6994,N_1570,N_354);
nand U6995 (N_6995,N_4670,N_1315);
or U6996 (N_6996,N_3030,N_1978);
nor U6997 (N_6997,N_4317,N_917);
nand U6998 (N_6998,N_3605,N_3472);
and U6999 (N_6999,N_2882,N_1845);
nand U7000 (N_7000,N_835,N_2328);
or U7001 (N_7001,N_4863,N_275);
and U7002 (N_7002,N_1976,N_3223);
or U7003 (N_7003,N_2542,N_4861);
and U7004 (N_7004,N_6071,N_2175);
and U7005 (N_7005,N_2324,N_6002);
nand U7006 (N_7006,N_2636,N_176);
nor U7007 (N_7007,N_5637,N_4745);
xnor U7008 (N_7008,N_5982,N_5224);
or U7009 (N_7009,N_1635,N_1094);
or U7010 (N_7010,N_2386,N_5308);
nor U7011 (N_7011,N_1768,N_1342);
and U7012 (N_7012,N_1595,N_939);
and U7013 (N_7013,N_5203,N_3599);
nand U7014 (N_7014,N_4378,N_5373);
xnor U7015 (N_7015,N_967,N_6190);
nor U7016 (N_7016,N_3451,N_4959);
and U7017 (N_7017,N_2916,N_5359);
or U7018 (N_7018,N_5893,N_717);
and U7019 (N_7019,N_2508,N_4275);
nor U7020 (N_7020,N_5401,N_6037);
and U7021 (N_7021,N_1073,N_4913);
and U7022 (N_7022,N_557,N_4092);
and U7023 (N_7023,N_484,N_5585);
and U7024 (N_7024,N_2079,N_1256);
nand U7025 (N_7025,N_2058,N_1719);
and U7026 (N_7026,N_3121,N_2976);
and U7027 (N_7027,N_6174,N_5959);
nor U7028 (N_7028,N_5765,N_5404);
nand U7029 (N_7029,N_452,N_4324);
or U7030 (N_7030,N_1411,N_3278);
nor U7031 (N_7031,N_5107,N_366);
nand U7032 (N_7032,N_1510,N_1008);
and U7033 (N_7033,N_4957,N_4308);
or U7034 (N_7034,N_6083,N_3222);
nor U7035 (N_7035,N_5393,N_3534);
and U7036 (N_7036,N_5238,N_4564);
and U7037 (N_7037,N_1064,N_4140);
nor U7038 (N_7038,N_4215,N_5328);
nand U7039 (N_7039,N_5538,N_19);
nor U7040 (N_7040,N_228,N_608);
nor U7041 (N_7041,N_3375,N_5788);
nand U7042 (N_7042,N_5774,N_5770);
or U7043 (N_7043,N_2333,N_3133);
nor U7044 (N_7044,N_3623,N_3175);
nor U7045 (N_7045,N_4114,N_4866);
nor U7046 (N_7046,N_385,N_3965);
nand U7047 (N_7047,N_3425,N_3642);
nand U7048 (N_7048,N_5235,N_646);
and U7049 (N_7049,N_3097,N_1217);
nor U7050 (N_7050,N_1764,N_5609);
nor U7051 (N_7051,N_4077,N_1164);
nor U7052 (N_7052,N_4557,N_1504);
nand U7053 (N_7053,N_2019,N_4037);
nand U7054 (N_7054,N_3870,N_1363);
nand U7055 (N_7055,N_3551,N_788);
and U7056 (N_7056,N_3422,N_3807);
and U7057 (N_7057,N_2357,N_2545);
or U7058 (N_7058,N_2317,N_2061);
or U7059 (N_7059,N_4442,N_2210);
nand U7060 (N_7060,N_2931,N_1132);
or U7061 (N_7061,N_4642,N_5062);
and U7062 (N_7062,N_79,N_6048);
or U7063 (N_7063,N_3892,N_485);
or U7064 (N_7064,N_4574,N_2158);
and U7065 (N_7065,N_769,N_2626);
nor U7066 (N_7066,N_1988,N_702);
and U7067 (N_7067,N_4509,N_5928);
nand U7068 (N_7068,N_5739,N_750);
nor U7069 (N_7069,N_2425,N_5402);
or U7070 (N_7070,N_2460,N_3606);
or U7071 (N_7071,N_5489,N_3039);
or U7072 (N_7072,N_197,N_897);
nor U7073 (N_7073,N_4392,N_4672);
or U7074 (N_7074,N_2875,N_2754);
or U7075 (N_7075,N_5657,N_779);
nor U7076 (N_7076,N_3582,N_3285);
and U7077 (N_7077,N_1730,N_3257);
and U7078 (N_7078,N_217,N_5260);
or U7079 (N_7079,N_5208,N_2592);
nor U7080 (N_7080,N_4395,N_3524);
or U7081 (N_7081,N_5183,N_3267);
nor U7082 (N_7082,N_2449,N_1252);
or U7083 (N_7083,N_1086,N_5364);
nand U7084 (N_7084,N_4605,N_5196);
and U7085 (N_7085,N_5090,N_5667);
and U7086 (N_7086,N_2839,N_5650);
or U7087 (N_7087,N_3413,N_443);
nand U7088 (N_7088,N_2114,N_959);
nand U7089 (N_7089,N_3758,N_873);
or U7090 (N_7090,N_5689,N_4753);
nor U7091 (N_7091,N_398,N_1253);
nor U7092 (N_7092,N_4282,N_4217);
nand U7093 (N_7093,N_4406,N_2703);
nand U7094 (N_7094,N_459,N_4369);
or U7095 (N_7095,N_1518,N_5519);
nand U7096 (N_7096,N_2049,N_2149);
nand U7097 (N_7097,N_1586,N_190);
and U7098 (N_7098,N_1167,N_3499);
and U7099 (N_7099,N_960,N_4837);
nand U7100 (N_7100,N_3610,N_2075);
nand U7101 (N_7101,N_1636,N_3970);
or U7102 (N_7102,N_1319,N_1665);
or U7103 (N_7103,N_261,N_5482);
or U7104 (N_7104,N_5813,N_148);
nand U7105 (N_7105,N_4329,N_2927);
nor U7106 (N_7106,N_2472,N_1533);
or U7107 (N_7107,N_2401,N_5907);
and U7108 (N_7108,N_4823,N_1359);
and U7109 (N_7109,N_2016,N_4210);
nor U7110 (N_7110,N_3455,N_1905);
and U7111 (N_7111,N_5978,N_5315);
nor U7112 (N_7112,N_3618,N_292);
xor U7113 (N_7113,N_2273,N_3814);
or U7114 (N_7114,N_2222,N_4080);
nand U7115 (N_7115,N_521,N_4946);
or U7116 (N_7116,N_2307,N_4958);
nand U7117 (N_7117,N_5380,N_1451);
nand U7118 (N_7118,N_5701,N_638);
nor U7119 (N_7119,N_4817,N_5136);
and U7120 (N_7120,N_1394,N_399);
and U7121 (N_7121,N_4067,N_2326);
and U7122 (N_7122,N_5349,N_1827);
nor U7123 (N_7123,N_1836,N_3077);
and U7124 (N_7124,N_4801,N_1026);
or U7125 (N_7125,N_173,N_3414);
nor U7126 (N_7126,N_1884,N_2904);
and U7127 (N_7127,N_2099,N_3434);
nor U7128 (N_7128,N_5157,N_116);
nand U7129 (N_7129,N_1024,N_4058);
or U7130 (N_7130,N_6155,N_3441);
nand U7131 (N_7131,N_1266,N_3063);
or U7132 (N_7132,N_5252,N_963);
and U7133 (N_7133,N_2186,N_4882);
and U7134 (N_7134,N_2408,N_4588);
nand U7135 (N_7135,N_1374,N_4975);
and U7136 (N_7136,N_5007,N_740);
or U7137 (N_7137,N_247,N_1020);
and U7138 (N_7138,N_2878,N_3802);
and U7139 (N_7139,N_4323,N_6145);
nand U7140 (N_7140,N_5443,N_315);
nor U7141 (N_7141,N_2392,N_37);
and U7142 (N_7142,N_5296,N_2771);
and U7143 (N_7143,N_4927,N_5784);
nand U7144 (N_7144,N_2496,N_2944);
or U7145 (N_7145,N_949,N_2055);
nand U7146 (N_7146,N_5078,N_2255);
nand U7147 (N_7147,N_3329,N_241);
and U7148 (N_7148,N_388,N_5115);
nor U7149 (N_7149,N_1922,N_5596);
and U7150 (N_7150,N_3200,N_1943);
nor U7151 (N_7151,N_1078,N_973);
and U7152 (N_7152,N_3320,N_3516);
or U7153 (N_7153,N_4659,N_853);
or U7154 (N_7154,N_3198,N_2733);
and U7155 (N_7155,N_738,N_3143);
nand U7156 (N_7156,N_3196,N_1612);
nand U7157 (N_7157,N_742,N_3600);
and U7158 (N_7158,N_5477,N_2192);
or U7159 (N_7159,N_4767,N_1644);
nor U7160 (N_7160,N_5245,N_193);
nor U7161 (N_7161,N_5211,N_2456);
and U7162 (N_7162,N_4868,N_4460);
nor U7163 (N_7163,N_673,N_5332);
nand U7164 (N_7164,N_2042,N_5188);
nand U7165 (N_7165,N_671,N_2304);
nor U7166 (N_7166,N_1778,N_1373);
xnor U7167 (N_7167,N_4788,N_1759);
or U7168 (N_7168,N_4013,N_5655);
nand U7169 (N_7169,N_5360,N_3344);
or U7170 (N_7170,N_1100,N_3681);
or U7171 (N_7171,N_6086,N_3676);
and U7172 (N_7172,N_473,N_3460);
xnor U7173 (N_7173,N_3935,N_4185);
nand U7174 (N_7174,N_4972,N_3068);
nand U7175 (N_7175,N_5589,N_2497);
nor U7176 (N_7176,N_2909,N_5919);
nor U7177 (N_7177,N_4700,N_6120);
nand U7178 (N_7178,N_2512,N_2671);
nand U7179 (N_7179,N_2907,N_5097);
nand U7180 (N_7180,N_833,N_3781);
and U7181 (N_7181,N_5105,N_1300);
or U7182 (N_7182,N_5922,N_5696);
nor U7183 (N_7183,N_2746,N_1786);
nor U7184 (N_7184,N_1430,N_4831);
nor U7185 (N_7185,N_153,N_1389);
nor U7186 (N_7186,N_805,N_3468);
nand U7187 (N_7187,N_3023,N_4001);
nor U7188 (N_7188,N_1957,N_1035);
nand U7189 (N_7189,N_5331,N_1502);
nand U7190 (N_7190,N_4373,N_352);
nand U7191 (N_7191,N_4948,N_522);
and U7192 (N_7192,N_2484,N_3464);
or U7193 (N_7193,N_412,N_5597);
or U7194 (N_7194,N_1501,N_5162);
and U7195 (N_7195,N_4814,N_6020);
and U7196 (N_7196,N_3972,N_1145);
nor U7197 (N_7197,N_3558,N_2920);
nand U7198 (N_7198,N_394,N_2003);
and U7199 (N_7199,N_6041,N_4355);
nand U7200 (N_7200,N_2872,N_105);
and U7201 (N_7201,N_1010,N_58);
and U7202 (N_7202,N_6199,N_1690);
nand U7203 (N_7203,N_4239,N_2519);
or U7204 (N_7204,N_4097,N_2091);
nand U7205 (N_7205,N_2725,N_3136);
nor U7206 (N_7206,N_3944,N_2581);
nor U7207 (N_7207,N_2001,N_5871);
or U7208 (N_7208,N_1210,N_647);
nor U7209 (N_7209,N_4581,N_1838);
nor U7210 (N_7210,N_6056,N_5500);
and U7211 (N_7211,N_857,N_807);
nor U7212 (N_7212,N_2047,N_728);
nor U7213 (N_7213,N_4257,N_2272);
and U7214 (N_7214,N_751,N_3628);
nand U7215 (N_7215,N_3988,N_377);
nor U7216 (N_7216,N_1056,N_2645);
and U7217 (N_7217,N_4828,N_20);
nor U7218 (N_7218,N_3117,N_2127);
and U7219 (N_7219,N_1118,N_2985);
or U7220 (N_7220,N_5889,N_4027);
or U7221 (N_7221,N_762,N_506);
and U7222 (N_7222,N_26,N_1136);
and U7223 (N_7223,N_3232,N_3447);
and U7224 (N_7224,N_4819,N_4335);
nor U7225 (N_7225,N_4607,N_6082);
nor U7226 (N_7226,N_685,N_4402);
nor U7227 (N_7227,N_5719,N_768);
nand U7228 (N_7228,N_3707,N_5410);
nand U7229 (N_7229,N_61,N_2588);
and U7230 (N_7230,N_3127,N_2694);
and U7231 (N_7231,N_4111,N_4325);
nor U7232 (N_7232,N_6132,N_2492);
and U7233 (N_7233,N_5141,N_5432);
and U7234 (N_7234,N_3339,N_456);
nor U7235 (N_7235,N_1785,N_4686);
and U7236 (N_7236,N_3343,N_864);
and U7237 (N_7237,N_4115,N_3666);
and U7238 (N_7238,N_3378,N_4714);
and U7239 (N_7239,N_5190,N_1005);
nor U7240 (N_7240,N_5232,N_1259);
nand U7241 (N_7241,N_1366,N_2835);
nor U7242 (N_7242,N_952,N_3653);
nor U7243 (N_7243,N_5674,N_2695);
or U7244 (N_7244,N_3398,N_18);
nand U7245 (N_7245,N_2871,N_609);
nor U7246 (N_7246,N_1999,N_189);
and U7247 (N_7247,N_693,N_1689);
or U7248 (N_7248,N_5547,N_5142);
or U7249 (N_7249,N_3757,N_3797);
or U7250 (N_7250,N_3293,N_1919);
and U7251 (N_7251,N_6011,N_4889);
and U7252 (N_7252,N_474,N_1238);
or U7253 (N_7253,N_4166,N_1335);
nor U7254 (N_7254,N_3563,N_5529);
nand U7255 (N_7255,N_3924,N_3664);
and U7256 (N_7256,N_4486,N_6159);
or U7257 (N_7257,N_5769,N_2698);
or U7258 (N_7258,N_3630,N_1370);
and U7259 (N_7259,N_5173,N_5827);
and U7260 (N_7260,N_3581,N_749);
nand U7261 (N_7261,N_2558,N_4970);
nand U7262 (N_7262,N_40,N_3669);
and U7263 (N_7263,N_4420,N_177);
or U7264 (N_7264,N_3633,N_2297);
nor U7265 (N_7265,N_5819,N_2409);
nand U7266 (N_7266,N_3138,N_4427);
nor U7267 (N_7267,N_3756,N_4296);
nor U7268 (N_7268,N_5551,N_1393);
or U7269 (N_7269,N_1858,N_5668);
and U7270 (N_7270,N_6053,N_1731);
and U7271 (N_7271,N_2775,N_2676);
nor U7272 (N_7272,N_2950,N_2048);
nand U7273 (N_7273,N_5110,N_2215);
nor U7274 (N_7274,N_3977,N_4093);
nor U7275 (N_7275,N_2997,N_2378);
nand U7276 (N_7276,N_1981,N_2752);
nor U7277 (N_7277,N_2992,N_5881);
nand U7278 (N_7278,N_1493,N_5595);
or U7279 (N_7279,N_3151,N_2791);
nor U7280 (N_7280,N_5045,N_980);
nor U7281 (N_7281,N_583,N_4146);
and U7282 (N_7282,N_1863,N_5883);
nand U7283 (N_7283,N_3163,N_1113);
and U7284 (N_7284,N_4712,N_2027);
nor U7285 (N_7285,N_4036,N_6185);
nand U7286 (N_7286,N_1579,N_6027);
nor U7287 (N_7287,N_290,N_1264);
and U7288 (N_7288,N_1895,N_2453);
and U7289 (N_7289,N_4516,N_1841);
and U7290 (N_7290,N_656,N_4225);
nand U7291 (N_7291,N_6004,N_5713);
nand U7292 (N_7292,N_2949,N_4394);
or U7293 (N_7293,N_5757,N_2993);
nor U7294 (N_7294,N_285,N_1193);
nand U7295 (N_7295,N_1478,N_1154);
or U7296 (N_7296,N_5524,N_5992);
nor U7297 (N_7297,N_3710,N_5634);
nor U7298 (N_7298,N_2237,N_1288);
or U7299 (N_7299,N_5348,N_2015);
nor U7300 (N_7300,N_1862,N_107);
nand U7301 (N_7301,N_102,N_2402);
and U7302 (N_7302,N_5672,N_664);
nand U7303 (N_7303,N_1548,N_773);
or U7304 (N_7304,N_4879,N_2278);
or U7305 (N_7305,N_1159,N_5720);
or U7306 (N_7306,N_3929,N_4973);
nand U7307 (N_7307,N_1545,N_6162);
nor U7308 (N_7308,N_5661,N_2521);
nand U7309 (N_7309,N_76,N_1757);
or U7310 (N_7310,N_747,N_855);
or U7311 (N_7311,N_4030,N_6147);
or U7312 (N_7312,N_4263,N_706);
nor U7313 (N_7313,N_4625,N_1309);
and U7314 (N_7314,N_2300,N_5001);
nor U7315 (N_7315,N_2085,N_527);
nor U7316 (N_7316,N_47,N_4501);
or U7317 (N_7317,N_4534,N_5337);
nor U7318 (N_7318,N_6017,N_5838);
nor U7319 (N_7319,N_350,N_4675);
or U7320 (N_7320,N_5312,N_4961);
and U7321 (N_7321,N_1507,N_1935);
and U7322 (N_7322,N_3889,N_1120);
xnor U7323 (N_7323,N_605,N_5939);
or U7324 (N_7324,N_5775,N_592);
or U7325 (N_7325,N_3190,N_3994);
nor U7326 (N_7326,N_3429,N_3028);
nor U7327 (N_7327,N_3021,N_2395);
nor U7328 (N_7328,N_1483,N_2721);
and U7329 (N_7329,N_1148,N_1603);
and U7330 (N_7330,N_4176,N_6119);
nand U7331 (N_7331,N_5690,N_2930);
xor U7332 (N_7332,N_4243,N_5514);
nand U7333 (N_7333,N_1071,N_5830);
nand U7334 (N_7334,N_1044,N_4361);
and U7335 (N_7335,N_2414,N_4568);
nand U7336 (N_7336,N_3895,N_5303);
nor U7337 (N_7337,N_5946,N_161);
or U7338 (N_7338,N_4118,N_572);
and U7339 (N_7339,N_2031,N_1695);
nand U7340 (N_7340,N_1908,N_1183);
or U7341 (N_7341,N_1669,N_2267);
nand U7342 (N_7342,N_2778,N_3391);
nand U7343 (N_7343,N_1171,N_3423);
nor U7344 (N_7344,N_4227,N_1998);
or U7345 (N_7345,N_5840,N_3007);
and U7346 (N_7346,N_5891,N_2795);
xnor U7347 (N_7347,N_4422,N_5254);
nand U7348 (N_7348,N_2000,N_6180);
and U7349 (N_7349,N_2179,N_5405);
or U7350 (N_7350,N_4881,N_4546);
nor U7351 (N_7351,N_4020,N_508);
nor U7352 (N_7352,N_378,N_3119);
or U7353 (N_7353,N_3917,N_4113);
nand U7354 (N_7354,N_5194,N_5491);
and U7355 (N_7355,N_4384,N_3996);
and U7356 (N_7356,N_1792,N_2498);
nand U7357 (N_7357,N_2661,N_2336);
nor U7358 (N_7358,N_2984,N_1444);
nand U7359 (N_7359,N_789,N_4691);
or U7360 (N_7360,N_639,N_1401);
and U7361 (N_7361,N_4404,N_2848);
and U7362 (N_7362,N_5398,N_5910);
or U7363 (N_7363,N_4454,N_1496);
and U7364 (N_7364,N_2925,N_3700);
nor U7365 (N_7365,N_4512,N_3309);
nand U7366 (N_7366,N_3215,N_2150);
and U7367 (N_7367,N_294,N_2867);
and U7368 (N_7368,N_343,N_2208);
nor U7369 (N_7369,N_382,N_5630);
nor U7370 (N_7370,N_4572,N_5509);
nor U7371 (N_7371,N_4109,N_3786);
or U7372 (N_7372,N_2635,N_1554);
and U7373 (N_7373,N_2634,N_4235);
and U7374 (N_7374,N_2742,N_46);
nand U7375 (N_7375,N_513,N_760);
and U7376 (N_7376,N_5148,N_3672);
nand U7377 (N_7377,N_2109,N_4815);
and U7378 (N_7378,N_796,N_1876);
nor U7379 (N_7379,N_4398,N_2204);
nor U7380 (N_7380,N_3210,N_386);
nand U7381 (N_7381,N_1258,N_2250);
and U7382 (N_7382,N_4760,N_6170);
or U7383 (N_7383,N_1639,N_6030);
nor U7384 (N_7384,N_4917,N_3636);
nor U7385 (N_7385,N_5013,N_4069);
nor U7386 (N_7386,N_344,N_5805);
or U7387 (N_7387,N_4382,N_1077);
and U7388 (N_7388,N_6016,N_978);
nor U7389 (N_7389,N_1497,N_4165);
and U7390 (N_7390,N_3096,N_1014);
nand U7391 (N_7391,N_6110,N_284);
and U7392 (N_7392,N_1346,N_2648);
nor U7393 (N_7393,N_6237,N_914);
nand U7394 (N_7394,N_6223,N_5755);
nand U7395 (N_7395,N_1515,N_1262);
and U7396 (N_7396,N_997,N_5799);
or U7397 (N_7397,N_554,N_300);
or U7398 (N_7398,N_4476,N_5706);
or U7399 (N_7399,N_2817,N_1728);
and U7400 (N_7400,N_1590,N_4678);
or U7401 (N_7401,N_1075,N_2768);
nor U7402 (N_7402,N_4966,N_2303);
nor U7403 (N_7403,N_5751,N_4055);
or U7404 (N_7404,N_4852,N_5705);
nor U7405 (N_7405,N_5143,N_3346);
nand U7406 (N_7406,N_5497,N_5495);
or U7407 (N_7407,N_4784,N_3603);
nand U7408 (N_7408,N_4633,N_2584);
or U7409 (N_7409,N_4391,N_5444);
and U7410 (N_7410,N_97,N_3332);
and U7411 (N_7411,N_2870,N_4306);
and U7412 (N_7412,N_5985,N_3824);
nor U7413 (N_7413,N_5850,N_4532);
and U7414 (N_7414,N_3874,N_3712);
nor U7415 (N_7415,N_3891,N_25);
nand U7416 (N_7416,N_2256,N_24);
and U7417 (N_7417,N_5068,N_565);
or U7418 (N_7418,N_4281,N_3169);
nor U7419 (N_7419,N_3348,N_4725);
nor U7420 (N_7420,N_5462,N_5229);
or U7421 (N_7421,N_4170,N_5560);
or U7422 (N_7422,N_5322,N_4269);
or U7423 (N_7423,N_3393,N_1424);
xnor U7424 (N_7424,N_4045,N_5848);
or U7425 (N_7425,N_1130,N_850);
and U7426 (N_7426,N_3191,N_2983);
nor U7427 (N_7427,N_763,N_1343);
nor U7428 (N_7428,N_900,N_2119);
nand U7429 (N_7429,N_5616,N_1047);
nor U7430 (N_7430,N_3024,N_4086);
or U7431 (N_7431,N_4303,N_492);
nand U7432 (N_7432,N_1267,N_1968);
nand U7433 (N_7433,N_6109,N_6018);
and U7434 (N_7434,N_3112,N_1544);
and U7435 (N_7435,N_3118,N_4911);
and U7436 (N_7436,N_2876,N_3366);
nand U7437 (N_7437,N_3768,N_4495);
or U7438 (N_7438,N_6166,N_3546);
or U7439 (N_7439,N_5931,N_657);
nor U7440 (N_7440,N_4430,N_2243);
nor U7441 (N_7441,N_1769,N_1693);
nand U7442 (N_7442,N_4733,N_2819);
or U7443 (N_7443,N_507,N_830);
and U7444 (N_7444,N_1889,N_4492);
nand U7445 (N_7445,N_1840,N_1516);
nor U7446 (N_7446,N_5600,N_5314);
or U7447 (N_7447,N_4907,N_4162);
or U7448 (N_7448,N_3412,N_403);
xnor U7449 (N_7449,N_3998,N_323);
nor U7450 (N_7450,N_3562,N_3794);
nor U7451 (N_7451,N_5820,N_135);
and U7452 (N_7452,N_3975,N_541);
and U7453 (N_7453,N_1153,N_2251);
and U7454 (N_7454,N_3031,N_3678);
nor U7455 (N_7455,N_4498,N_824);
or U7456 (N_7456,N_3813,N_5035);
or U7457 (N_7457,N_5354,N_1558);
or U7458 (N_7458,N_4981,N_2729);
nand U7459 (N_7459,N_4890,N_2390);
nand U7460 (N_7460,N_2080,N_5764);
nor U7461 (N_7461,N_2578,N_5484);
or U7462 (N_7462,N_1766,N_1739);
nor U7463 (N_7463,N_5855,N_2206);
nor U7464 (N_7464,N_1971,N_1425);
nand U7465 (N_7465,N_2078,N_373);
and U7466 (N_7466,N_4339,N_1991);
nand U7467 (N_7467,N_103,N_4737);
nor U7468 (N_7468,N_2688,N_5987);
nor U7469 (N_7469,N_4010,N_1226);
and U7470 (N_7470,N_3898,N_2298);
and U7471 (N_7471,N_131,N_3195);
nand U7472 (N_7472,N_2856,N_3848);
nand U7473 (N_7473,N_3230,N_771);
nand U7474 (N_7474,N_581,N_1656);
nand U7475 (N_7475,N_4998,N_699);
nor U7476 (N_7476,N_2348,N_5962);
nand U7477 (N_7477,N_765,N_3909);
or U7478 (N_7478,N_3787,N_1041);
nor U7479 (N_7479,N_3056,N_2511);
and U7480 (N_7480,N_4314,N_3025);
nand U7481 (N_7481,N_1176,N_12);
xnor U7482 (N_7482,N_4873,N_3995);
and U7483 (N_7483,N_5718,N_2448);
nor U7484 (N_7484,N_3532,N_701);
or U7485 (N_7485,N_429,N_1745);
and U7486 (N_7486,N_2861,N_462);
nand U7487 (N_7487,N_1459,N_1546);
nor U7488 (N_7488,N_1794,N_884);
nand U7489 (N_7489,N_1506,N_4899);
or U7490 (N_7490,N_1477,N_5417);
nor U7491 (N_7491,N_4582,N_3844);
nor U7492 (N_7492,N_2145,N_710);
or U7493 (N_7493,N_3205,N_23);
nand U7494 (N_7494,N_6038,N_4579);
or U7495 (N_7495,N_5273,N_4209);
nand U7496 (N_7496,N_4472,N_983);
nand U7497 (N_7497,N_5747,N_393);
and U7498 (N_7498,N_5137,N_3374);
nor U7499 (N_7499,N_655,N_4808);
nor U7500 (N_7500,N_2013,N_3492);
nand U7501 (N_7501,N_3055,N_1688);
or U7502 (N_7502,N_5714,N_3342);
nor U7503 (N_7503,N_4663,N_5488);
or U7504 (N_7504,N_950,N_3736);
nor U7505 (N_7505,N_4857,N_2792);
or U7506 (N_7506,N_2037,N_5584);
nor U7507 (N_7507,N_3570,N_2325);
nand U7508 (N_7508,N_4346,N_383);
and U7509 (N_7509,N_6213,N_2020);
nor U7510 (N_7510,N_727,N_1196);
and U7511 (N_7511,N_856,N_3906);
or U7512 (N_7512,N_4360,N_4613);
or U7513 (N_7513,N_5612,N_1947);
or U7514 (N_7514,N_766,N_99);
nand U7515 (N_7515,N_1225,N_3665);
nor U7516 (N_7516,N_3008,N_5374);
nor U7517 (N_7517,N_4063,N_863);
or U7518 (N_7518,N_2913,N_4685);
nand U7519 (N_7519,N_2391,N_2776);
xnor U7520 (N_7520,N_2693,N_908);
nor U7521 (N_7521,N_579,N_1828);
nand U7522 (N_7522,N_2968,N_4078);
nor U7523 (N_7523,N_4820,N_2490);
and U7524 (N_7524,N_3153,N_4860);
nand U7525 (N_7525,N_1449,N_3878);
nor U7526 (N_7526,N_988,N_259);
or U7527 (N_7527,N_752,N_1109);
nand U7528 (N_7528,N_1472,N_1111);
or U7529 (N_7529,N_4660,N_489);
and U7530 (N_7530,N_2526,N_5501);
nor U7531 (N_7531,N_4813,N_611);
nand U7532 (N_7532,N_1019,N_1052);
nor U7533 (N_7533,N_4088,N_5562);
nand U7534 (N_7534,N_2935,N_2198);
nor U7535 (N_7535,N_2330,N_5485);
or U7536 (N_7536,N_3842,N_1909);
nor U7537 (N_7537,N_2094,N_3461);
or U7538 (N_7538,N_3377,N_2350);
nor U7539 (N_7539,N_6099,N_2879);
nand U7540 (N_7540,N_4711,N_4792);
or U7541 (N_7541,N_1826,N_53);
nand U7542 (N_7542,N_4504,N_1680);
nor U7543 (N_7543,N_1107,N_2426);
nand U7544 (N_7544,N_1488,N_5177);
nand U7545 (N_7545,N_2002,N_3566);
nor U7546 (N_7546,N_6149,N_493);
or U7547 (N_7547,N_1347,N_5474);
nand U7548 (N_7548,N_4363,N_5134);
nand U7549 (N_7549,N_3318,N_3300);
nor U7550 (N_7550,N_3199,N_2660);
or U7551 (N_7551,N_5131,N_1437);
and U7552 (N_7552,N_3081,N_1308);
nand U7553 (N_7553,N_4285,N_5730);
nand U7554 (N_7554,N_3783,N_2990);
or U7555 (N_7555,N_662,N_3265);
nor U7556 (N_7556,N_5175,N_2582);
and U7557 (N_7557,N_5222,N_4340);
nand U7558 (N_7558,N_6245,N_4334);
nor U7559 (N_7559,N_4297,N_4953);
nor U7560 (N_7560,N_2863,N_3536);
or U7561 (N_7561,N_1200,N_5803);
nor U7562 (N_7562,N_1791,N_2007);
or U7563 (N_7563,N_3410,N_4266);
and U7564 (N_7564,N_4781,N_3240);
and U7565 (N_7565,N_4591,N_5543);
or U7566 (N_7566,N_73,N_4436);
or U7567 (N_7567,N_5974,N_2461);
or U7568 (N_7568,N_2728,N_3463);
nor U7569 (N_7569,N_811,N_1049);
or U7570 (N_7570,N_477,N_3648);
and U7571 (N_7571,N_335,N_1202);
nand U7572 (N_7572,N_5361,N_3168);
nand U7573 (N_7573,N_5810,N_144);
nor U7574 (N_7574,N_4744,N_4256);
nand U7575 (N_7575,N_2952,N_4987);
and U7576 (N_7576,N_1467,N_4517);
nor U7577 (N_7577,N_4840,N_5247);
or U7578 (N_7578,N_155,N_4727);
nand U7579 (N_7579,N_836,N_163);
nand U7580 (N_7580,N_4389,N_1233);
nand U7581 (N_7581,N_3406,N_4706);
nand U7582 (N_7582,N_1729,N_1135);
nand U7583 (N_7583,N_4040,N_2804);
or U7584 (N_7584,N_5868,N_4261);
nand U7585 (N_7585,N_113,N_4969);
or U7586 (N_7586,N_3592,N_5913);
or U7587 (N_7587,N_3840,N_4758);
nand U7588 (N_7588,N_5675,N_3189);
and U7589 (N_7589,N_1085,N_5351);
or U7590 (N_7590,N_1354,N_2140);
or U7591 (N_7591,N_2486,N_3481);
nor U7592 (N_7592,N_2082,N_425);
or U7593 (N_7593,N_4825,N_2607);
nor U7594 (N_7594,N_1962,N_4264);
and U7595 (N_7595,N_3671,N_1749);
nand U7596 (N_7596,N_2842,N_764);
xnor U7597 (N_7597,N_5030,N_2537);
xor U7598 (N_7598,N_1108,N_799);
nand U7599 (N_7599,N_5989,N_4240);
and U7600 (N_7600,N_1753,N_2777);
nand U7601 (N_7601,N_442,N_3427);
or U7602 (N_7602,N_4940,N_4662);
and U7603 (N_7603,N_1593,N_2261);
nor U7604 (N_7604,N_74,N_1958);
nand U7605 (N_7605,N_2717,N_2557);
nand U7606 (N_7606,N_5960,N_5268);
and U7607 (N_7607,N_5926,N_5593);
and U7608 (N_7608,N_1513,N_4802);
and U7609 (N_7609,N_218,N_4295);
xnor U7610 (N_7610,N_4085,N_6031);
and U7611 (N_7611,N_5957,N_2846);
or U7612 (N_7612,N_4014,N_5561);
or U7613 (N_7613,N_1152,N_2911);
and U7614 (N_7614,N_3966,N_634);
nand U7615 (N_7615,N_6241,N_736);
or U7616 (N_7616,N_5020,N_5636);
xnor U7617 (N_7617,N_480,N_3939);
or U7618 (N_7618,N_3701,N_4811);
xnor U7619 (N_7619,N_4715,N_4854);
or U7620 (N_7620,N_5283,N_1774);
and U7621 (N_7621,N_4742,N_2538);
and U7622 (N_7622,N_1452,N_1368);
nand U7623 (N_7623,N_4159,N_923);
and U7624 (N_7624,N_965,N_3693);
nand U7625 (N_7625,N_3886,N_2597);
or U7626 (N_7626,N_5466,N_1640);
xor U7627 (N_7627,N_1138,N_2216);
xor U7628 (N_7628,N_3788,N_3134);
and U7629 (N_7629,N_185,N_142);
nand U7630 (N_7630,N_5106,N_5552);
nor U7631 (N_7631,N_3517,N_1364);
nand U7632 (N_7632,N_4963,N_2708);
nand U7633 (N_7633,N_1627,N_2686);
and U7634 (N_7634,N_4152,N_5686);
and U7635 (N_7635,N_4787,N_5847);
or U7636 (N_7636,N_711,N_1096);
nand U7637 (N_7637,N_1779,N_5023);
and U7638 (N_7638,N_1236,N_4265);
nor U7639 (N_7639,N_4238,N_2803);
xnor U7640 (N_7640,N_3322,N_4433);
nor U7641 (N_7641,N_424,N_5692);
and U7642 (N_7642,N_1417,N_537);
and U7643 (N_7643,N_4920,N_519);
and U7644 (N_7644,N_3316,N_3677);
nand U7645 (N_7645,N_5034,N_2544);
xor U7646 (N_7646,N_2236,N_1142);
or U7647 (N_7647,N_1344,N_694);
nand U7648 (N_7648,N_85,N_1291);
or U7649 (N_7649,N_2812,N_2481);
or U7650 (N_7650,N_3431,N_5753);
or U7651 (N_7651,N_3446,N_69);
and U7652 (N_7652,N_4049,N_38);
nand U7653 (N_7653,N_1345,N_6040);
nand U7654 (N_7654,N_3324,N_72);
nand U7655 (N_7655,N_5744,N_4007);
nand U7656 (N_7656,N_4473,N_2561);
nor U7657 (N_7657,N_5955,N_5396);
nor U7658 (N_7658,N_3061,N_1679);
and U7659 (N_7659,N_3967,N_5687);
or U7660 (N_7660,N_3216,N_3338);
nand U7661 (N_7661,N_6196,N_5777);
and U7662 (N_7662,N_2435,N_919);
nand U7663 (N_7663,N_3679,N_1227);
nor U7664 (N_7664,N_1065,N_5522);
nand U7665 (N_7665,N_400,N_4206);
and U7666 (N_7666,N_5325,N_2353);
nand U7667 (N_7667,N_5864,N_1983);
nor U7668 (N_7668,N_4867,N_4971);
or U7669 (N_7669,N_757,N_469);
nor U7670 (N_7670,N_1116,N_441);
nand U7671 (N_7671,N_1521,N_1967);
and U7672 (N_7672,N_4312,N_2315);
nand U7673 (N_7673,N_4979,N_5929);
nor U7674 (N_7674,N_1878,N_795);
or U7675 (N_7675,N_1536,N_138);
or U7676 (N_7676,N_4475,N_4117);
nand U7677 (N_7677,N_3847,N_911);
and U7678 (N_7678,N_3496,N_1422);
nand U7679 (N_7679,N_4924,N_5918);
nand U7680 (N_7680,N_3667,N_2589);
nand U7681 (N_7681,N_4618,N_5866);
and U7682 (N_7682,N_2072,N_1399);
nand U7683 (N_7683,N_2769,N_2770);
nand U7684 (N_7684,N_3385,N_5236);
or U7685 (N_7685,N_801,N_2858);
or U7686 (N_7686,N_3129,N_2052);
or U7687 (N_7687,N_536,N_4728);
or U7688 (N_7688,N_216,N_3029);
nor U7689 (N_7689,N_2958,N_5532);
nand U7690 (N_7690,N_1182,N_5345);
xor U7691 (N_7691,N_324,N_3386);
or U7692 (N_7692,N_5029,N_5791);
nor U7693 (N_7693,N_4596,N_3560);
and U7694 (N_7694,N_2606,N_1671);
nand U7695 (N_7695,N_4134,N_2797);
or U7696 (N_7696,N_461,N_1460);
nand U7697 (N_7697,N_4250,N_3539);
and U7698 (N_7698,N_542,N_5472);
nand U7699 (N_7699,N_5906,N_3815);
or U7700 (N_7700,N_714,N_3612);
nor U7701 (N_7701,N_1532,N_2849);
or U7702 (N_7702,N_3262,N_4666);
or U7703 (N_7703,N_3379,N_5214);
and U7704 (N_7704,N_2302,N_465);
and U7705 (N_7705,N_758,N_607);
and U7706 (N_7706,N_2986,N_5602);
and U7707 (N_7707,N_2736,N_5126);
or U7708 (N_7708,N_1290,N_4531);
nand U7709 (N_7709,N_550,N_139);
nand U7710 (N_7710,N_3060,N_4409);
nor U7711 (N_7711,N_3148,N_1803);
or U7712 (N_7712,N_620,N_4041);
nand U7713 (N_7713,N_3760,N_1668);
or U7714 (N_7714,N_4912,N_670);
and U7715 (N_7715,N_734,N_629);
nand U7716 (N_7716,N_709,N_1367);
and U7717 (N_7717,N_5607,N_5806);
nor U7718 (N_7718,N_2965,N_5118);
nand U7719 (N_7719,N_2398,N_280);
nor U7720 (N_7720,N_1012,N_2181);
nor U7721 (N_7721,N_5306,N_2894);
or U7722 (N_7722,N_5139,N_4054);
and U7723 (N_7723,N_5179,N_1569);
and U7724 (N_7724,N_2165,N_915);
and U7725 (N_7725,N_2026,N_4526);
nor U7726 (N_7726,N_4990,N_2785);
nand U7727 (N_7727,N_1498,N_4254);
nand U7728 (N_7728,N_1487,N_1854);
and U7729 (N_7729,N_6220,N_1376);
nand U7730 (N_7730,N_211,N_3440);
or U7731 (N_7731,N_6197,N_6042);
xor U7732 (N_7732,N_3779,N_4631);
nand U7733 (N_7733,N_3006,N_5422);
or U7734 (N_7734,N_5041,N_2630);
or U7735 (N_7735,N_4365,N_1659);
or U7736 (N_7736,N_5837,N_5395);
nor U7737 (N_7737,N_4778,N_5977);
nand U7738 (N_7738,N_368,N_5389);
nor U7739 (N_7739,N_1445,N_652);
nand U7740 (N_7740,N_3974,N_2040);
nor U7741 (N_7741,N_533,N_4869);
and U7742 (N_7742,N_1385,N_4488);
nand U7743 (N_7743,N_3656,N_365);
and U7744 (N_7744,N_5123,N_4762);
or U7745 (N_7745,N_4231,N_1524);
and U7746 (N_7746,N_3308,N_2847);
nand U7747 (N_7747,N_1600,N_1843);
nand U7748 (N_7748,N_157,N_3088);
and U7749 (N_7749,N_4836,N_1316);
and U7750 (N_7750,N_4371,N_5338);
xnor U7751 (N_7751,N_490,N_6123);
or U7752 (N_7752,N_3014,N_4026);
nand U7753 (N_7753,N_6208,N_3353);
and U7754 (N_7754,N_1859,N_4478);
or U7755 (N_7755,N_39,N_2629);
nand U7756 (N_7756,N_4136,N_4213);
or U7757 (N_7757,N_4157,N_1219);
nor U7758 (N_7758,N_6059,N_659);
or U7759 (N_7759,N_77,N_5458);
or U7760 (N_7760,N_3596,N_707);
nand U7761 (N_7761,N_3968,N_1242);
nor U7762 (N_7762,N_2864,N_4403);
or U7763 (N_7763,N_5763,N_2429);
or U7764 (N_7764,N_158,N_6184);
nand U7765 (N_7765,N_2502,N_140);
or U7766 (N_7766,N_86,N_890);
or U7767 (N_7767,N_2818,N_2260);
and U7768 (N_7768,N_6200,N_3358);
or U7769 (N_7769,N_2885,N_5633);
or U7770 (N_7770,N_4104,N_5478);
and U7771 (N_7771,N_2469,N_6231);
or U7772 (N_7772,N_43,N_341);
nand U7773 (N_7773,N_5531,N_2252);
or U7774 (N_7774,N_2487,N_5779);
or U7775 (N_7775,N_6230,N_1269);
nand U7776 (N_7776,N_3302,N_5831);
and U7777 (N_7777,N_2529,N_538);
nor U7778 (N_7778,N_3640,N_1795);
xnor U7779 (N_7779,N_496,N_1888);
nor U7780 (N_7780,N_2783,N_6248);
nor U7781 (N_7781,N_3856,N_1652);
nand U7782 (N_7782,N_6064,N_2217);
nand U7783 (N_7783,N_4600,N_3152);
nand U7784 (N_7784,N_3401,N_2399);
nand U7785 (N_7785,N_2917,N_6115);
nand U7786 (N_7786,N_3131,N_5750);
or U7787 (N_7787,N_6195,N_3491);
nor U7788 (N_7788,N_4561,N_5740);
nand U7789 (N_7789,N_1170,N_3748);
nand U7790 (N_7790,N_786,N_5521);
nand U7791 (N_7791,N_5901,N_1517);
nand U7792 (N_7792,N_4292,N_5699);
nand U7793 (N_7793,N_3817,N_3528);
nor U7794 (N_7794,N_3639,N_233);
or U7795 (N_7795,N_2991,N_4044);
nand U7796 (N_7796,N_4923,N_6112);
or U7797 (N_7797,N_3989,N_2129);
and U7798 (N_7798,N_2926,N_4321);
nand U7799 (N_7799,N_5412,N_2005);
and U7800 (N_7800,N_3170,N_2066);
and U7801 (N_7801,N_3668,N_2604);
nand U7802 (N_7802,N_3943,N_3430);
and U7803 (N_7803,N_2442,N_124);
or U7804 (N_7804,N_6050,N_5336);
xor U7805 (N_7805,N_755,N_5055);
nand U7806 (N_7806,N_4541,N_932);
nand U7807 (N_7807,N_621,N_3746);
or U7808 (N_7808,N_3704,N_2678);
and U7809 (N_7809,N_1067,N_2567);
nor U7810 (N_7810,N_3298,N_5679);
or U7811 (N_7811,N_2264,N_4628);
nand U7812 (N_7812,N_192,N_5903);
and U7813 (N_7813,N_2289,N_2801);
and U7814 (N_7814,N_6024,N_2960);
nor U7815 (N_7815,N_1638,N_6242);
nand U7816 (N_7816,N_254,N_3352);
and U7817 (N_7817,N_841,N_4144);
or U7818 (N_7818,N_4694,N_4554);
and U7819 (N_7819,N_3923,N_3139);
nor U7820 (N_7820,N_2135,N_871);
nand U7821 (N_7821,N_475,N_731);
nor U7822 (N_7822,N_2043,N_1194);
and U7823 (N_7823,N_518,N_100);
or U7824 (N_7824,N_2877,N_4138);
nor U7825 (N_7825,N_2653,N_4800);
nand U7826 (N_7826,N_1099,N_2657);
or U7827 (N_7827,N_5420,N_4730);
nor U7828 (N_7828,N_132,N_4835);
or U7829 (N_7829,N_1945,N_4260);
and U7830 (N_7830,N_1441,N_1270);
and U7831 (N_7831,N_1721,N_1025);
nand U7832 (N_7832,N_2380,N_3101);
or U7833 (N_7833,N_1814,N_229);
or U7834 (N_7834,N_2888,N_3331);
nor U7835 (N_7835,N_883,N_1801);
nor U7836 (N_7836,N_5217,N_4821);
nor U7837 (N_7837,N_6076,N_1301);
or U7838 (N_7838,N_2428,N_1243);
nand U7839 (N_7839,N_3793,N_2836);
or U7840 (N_7840,N_4773,N_5941);
and U7841 (N_7841,N_1856,N_2668);
and U7842 (N_7842,N_6095,N_612);
or U7843 (N_7843,N_1068,N_3711);
nand U7844 (N_7844,N_5617,N_2137);
nor U7845 (N_7845,N_5079,N_3547);
nor U7846 (N_7846,N_4127,N_2450);
nor U7847 (N_7847,N_6029,N_3157);
or U7848 (N_7848,N_5039,N_2126);
nor U7849 (N_7849,N_5219,N_5825);
and U7850 (N_7850,N_3990,N_935);
nor U7851 (N_7851,N_2209,N_4777);
or U7852 (N_7852,N_3073,N_1911);
or U7853 (N_7853,N_3166,N_4214);
nor U7854 (N_7854,N_4636,N_2826);
nor U7855 (N_7855,N_4539,N_4432);
nand U7856 (N_7856,N_1160,N_2352);
nor U7857 (N_7857,N_1251,N_6226);
nor U7858 (N_7858,N_5786,N_3810);
nand U7859 (N_7859,N_4255,N_4906);
nor U7860 (N_7860,N_1784,N_5112);
nand U7861 (N_7861,N_3040,N_4370);
nor U7862 (N_7862,N_4775,N_4681);
and U7863 (N_7863,N_4145,N_4849);
nand U7864 (N_7864,N_5525,N_4494);
or U7865 (N_7865,N_936,N_2153);
nor U7866 (N_7866,N_3531,N_3778);
nand U7867 (N_7867,N_4577,N_5695);
and U7868 (N_7868,N_5908,N_1707);
and U7869 (N_7869,N_4094,N_5966);
or U7870 (N_7870,N_770,N_374);
nor U7871 (N_7871,N_3264,N_2869);
nand U7872 (N_7872,N_5651,N_1201);
nand U7873 (N_7873,N_3690,N_3317);
nor U7874 (N_7874,N_2696,N_3888);
nand U7875 (N_7875,N_5800,N_4130);
or U7876 (N_7876,N_4161,N_3747);
and U7877 (N_7877,N_3367,N_3646);
nand U7878 (N_7878,N_5582,N_5342);
or U7879 (N_7879,N_5170,N_5754);
or U7880 (N_7880,N_3072,N_1822);
nor U7881 (N_7881,N_5333,N_3150);
and U7882 (N_7882,N_1512,N_127);
or U7883 (N_7883,N_4341,N_635);
nand U7884 (N_7884,N_4050,N_2551);
and U7885 (N_7885,N_5656,N_6171);
nor U7886 (N_7886,N_5712,N_4931);
nor U7887 (N_7887,N_1318,N_22);
or U7888 (N_7888,N_3382,N_6006);
and U7889 (N_7889,N_2171,N_4832);
nor U7890 (N_7890,N_2928,N_4903);
nand U7891 (N_7891,N_2643,N_4318);
nor U7892 (N_7892,N_5074,N_2912);
or U7893 (N_7893,N_4984,N_4065);
nand U7894 (N_7894,N_4073,N_6224);
nand U7895 (N_7895,N_1490,N_2681);
or U7896 (N_7896,N_4790,N_5487);
nand U7897 (N_7897,N_5875,N_3235);
and U7898 (N_7898,N_3043,N_643);
nand U7899 (N_7899,N_5206,N_3142);
or U7900 (N_7900,N_5669,N_6069);
nor U7901 (N_7901,N_5227,N_4905);
and U7902 (N_7902,N_1388,N_6227);
nand U7903 (N_7903,N_3439,N_3362);
nor U7904 (N_7904,N_4829,N_1677);
nor U7905 (N_7905,N_3770,N_3527);
and U7906 (N_7906,N_4615,N_3224);
nor U7907 (N_7907,N_2651,N_219);
nand U7908 (N_7908,N_2412,N_1711);
or U7909 (N_7909,N_3537,N_207);
nor U7910 (N_7910,N_5683,N_5857);
and U7911 (N_7911,N_2231,N_3688);
or U7912 (N_7912,N_708,N_2510);
nand U7913 (N_7913,N_1628,N_4479);
nand U7914 (N_7914,N_5789,N_523);
nand U7915 (N_7915,N_781,N_2283);
or U7916 (N_7916,N_3745,N_1578);
nand U7917 (N_7917,N_5257,N_421);
and U7918 (N_7918,N_2219,N_2418);
or U7919 (N_7919,N_364,N_3708);
or U7920 (N_7920,N_3046,N_5610);
nor U7921 (N_7921,N_1104,N_4667);
nor U7922 (N_7922,N_5697,N_4189);
and U7923 (N_7923,N_3497,N_5077);
nand U7924 (N_7924,N_2865,N_1712);
and U7925 (N_7925,N_5280,N_4431);
and U7926 (N_7926,N_2633,N_589);
nor U7927 (N_7927,N_6092,N_4624);
and U7928 (N_7928,N_6052,N_5161);
and U7929 (N_7929,N_1283,N_1526);
nor U7930 (N_7930,N_991,N_1552);
nand U7931 (N_7931,N_2212,N_4244);
or U7932 (N_7932,N_5011,N_4716);
or U7933 (N_7933,N_6178,N_5807);
or U7934 (N_7934,N_5564,N_3181);
or U7935 (N_7935,N_2447,N_1332);
and U7936 (N_7936,N_4876,N_6106);
nor U7937 (N_7937,N_4884,N_6021);
or U7938 (N_7938,N_66,N_1204);
or U7939 (N_7939,N_5166,N_4897);
and U7940 (N_7940,N_4181,N_3899);
nand U7941 (N_7941,N_1752,N_2605);
and U7942 (N_7942,N_4090,N_5042);
nor U7943 (N_7943,N_5520,N_4772);
or U7944 (N_7944,N_1993,N_2884);
nor U7945 (N_7945,N_3183,N_2499);
and U7946 (N_7946,N_145,N_1747);
nand U7947 (N_7947,N_1079,N_5414);
and U7948 (N_7948,N_2650,N_3281);
nand U7949 (N_7949,N_4132,N_6066);
nand U7950 (N_7950,N_1986,N_700);
and U7951 (N_7951,N_510,N_5909);
and U7952 (N_7952,N_83,N_790);
or U7953 (N_7953,N_3754,N_110);
nor U7954 (N_7954,N_5392,N_5797);
or U7955 (N_7955,N_2764,N_4490);
nor U7956 (N_7956,N_961,N_4841);
or U7957 (N_7957,N_1147,N_957);
or U7958 (N_7958,N_4038,N_754);
or U7959 (N_7959,N_5995,N_644);
and U7960 (N_7960,N_5790,N_698);
nand U7961 (N_7961,N_3593,N_2765);
nor U7962 (N_7962,N_3626,N_6160);
nor U7963 (N_7963,N_5508,N_5220);
and U7964 (N_7964,N_166,N_5996);
nand U7965 (N_7965,N_311,N_3952);
nand U7966 (N_7966,N_418,N_3167);
nand U7967 (N_7967,N_5424,N_2868);
and U7968 (N_7968,N_5993,N_5317);
nand U7969 (N_7969,N_4935,N_2528);
nor U7970 (N_7970,N_842,N_5731);
and U7971 (N_7971,N_4752,N_204);
nor U7972 (N_7972,N_5071,N_2195);
or U7973 (N_7973,N_4764,N_391);
nor U7974 (N_7974,N_1900,N_5388);
nand U7975 (N_7975,N_6070,N_3776);
or U7976 (N_7976,N_3204,N_2747);
nor U7977 (N_7977,N_2112,N_3286);
or U7978 (N_7978,N_1059,N_5542);
nand U7979 (N_7979,N_5849,N_447);
or U7980 (N_7980,N_2982,N_5279);
nor U7981 (N_7981,N_2446,N_5879);
or U7982 (N_7982,N_2874,N_1446);
or U7983 (N_7983,N_4357,N_4414);
nand U7984 (N_7984,N_4129,N_3860);
and U7985 (N_7985,N_3987,N_3616);
and U7986 (N_7986,N_5096,N_4602);
and U7987 (N_7987,N_4108,N_4502);
and U7988 (N_7988,N_3635,N_4567);
and U7989 (N_7989,N_5882,N_2520);
and U7990 (N_7990,N_5169,N_3079);
nand U7991 (N_7991,N_5878,N_5642);
nor U7992 (N_7992,N_3456,N_33);
or U7993 (N_7993,N_2141,N_1172);
and U7994 (N_7994,N_753,N_642);
nand U7995 (N_7995,N_4503,N_4193);
nor U7996 (N_7996,N_6221,N_545);
nor U7997 (N_7997,N_5060,N_1528);
nand U7998 (N_7998,N_1386,N_3192);
or U7999 (N_7999,N_5212,N_3956);
and U8000 (N_8000,N_2837,N_1016);
nand U8001 (N_8001,N_3567,N_3964);
or U8002 (N_8002,N_2627,N_1260);
nor U8003 (N_8003,N_3825,N_3486);
nor U8004 (N_8004,N_574,N_4004);
and U8005 (N_8005,N_3160,N_1589);
nand U8006 (N_8006,N_4967,N_5470);
nor U8007 (N_8007,N_338,N_2115);
nor U8008 (N_8008,N_2759,N_4804);
or U8009 (N_8009,N_4287,N_1924);
nor U8010 (N_8010,N_6186,N_5165);
xor U8011 (N_8011,N_1037,N_1419);
nor U8012 (N_8012,N_5781,N_3784);
and U8013 (N_8013,N_3094,N_4641);
nand U8014 (N_8014,N_878,N_4087);
or U8015 (N_8015,N_5291,N_793);
nor U8016 (N_8016,N_1124,N_3550);
and U8017 (N_8017,N_3197,N_2053);
and U8018 (N_8018,N_476,N_4619);
nor U8019 (N_8019,N_2276,N_3872);
nand U8020 (N_8020,N_682,N_938);
or U8021 (N_8021,N_1169,N_5890);
and U8022 (N_8022,N_5099,N_1229);
nand U8023 (N_8023,N_5449,N_1043);
and U8024 (N_8024,N_4921,N_2954);
or U8025 (N_8025,N_416,N_3673);
or U8026 (N_8026,N_5439,N_4081);
and U8027 (N_8027,N_4515,N_1869);
or U8028 (N_8028,N_3459,N_1163);
or U8029 (N_8029,N_5896,N_483);
or U8030 (N_8030,N_3259,N_5575);
or U8031 (N_8031,N_4110,N_2891);
and U8032 (N_8032,N_974,N_3843);
and U8033 (N_8033,N_5330,N_4309);
nor U8034 (N_8034,N_2081,N_4904);
nor U8035 (N_8035,N_1973,N_2652);
or U8036 (N_8036,N_1944,N_2981);
nand U8037 (N_8037,N_4592,N_1220);
nand U8038 (N_8038,N_2096,N_6168);
nor U8039 (N_8039,N_2951,N_3000);
nand U8040 (N_8040,N_258,N_3469);
nand U8041 (N_8041,N_2955,N_2744);
and U8042 (N_8042,N_3411,N_4400);
or U8043 (N_8043,N_5347,N_3649);
nor U8044 (N_8044,N_5085,N_3535);
or U8045 (N_8045,N_1960,N_1418);
and U8046 (N_8046,N_4057,N_5243);
or U8047 (N_8047,N_3247,N_5371);
nand U8048 (N_8048,N_5048,N_4748);
nor U8049 (N_8049,N_3102,N_4423);
nand U8050 (N_8050,N_4028,N_1576);
nor U8051 (N_8051,N_5383,N_785);
nor U8052 (N_8052,N_6183,N_5149);
nor U8053 (N_8053,N_1793,N_4806);
and U8054 (N_8054,N_3686,N_2440);
nand U8055 (N_8055,N_3540,N_3110);
or U8056 (N_8056,N_390,N_4960);
or U8057 (N_8057,N_1713,N_4583);
or U8058 (N_8058,N_2327,N_4416);
or U8059 (N_8059,N_120,N_4930);
or U8060 (N_8060,N_5844,N_438);
nor U8061 (N_8061,N_2369,N_4795);
or U8062 (N_8062,N_1466,N_3837);
nor U8063 (N_8063,N_68,N_561);
nand U8064 (N_8064,N_6210,N_4017);
or U8065 (N_8065,N_3363,N_3513);
and U8066 (N_8066,N_5904,N_3620);
nor U8067 (N_8067,N_2977,N_367);
nor U8068 (N_8068,N_3370,N_5381);
nor U8069 (N_8069,N_4497,N_2406);
nor U8070 (N_8070,N_3830,N_3533);
nand U8071 (N_8071,N_2371,N_3634);
nor U8072 (N_8072,N_1468,N_3887);
and U8073 (N_8073,N_5664,N_663);
nand U8074 (N_8074,N_1090,N_901);
or U8075 (N_8075,N_3862,N_3962);
and U8076 (N_8076,N_746,N_3698);
or U8077 (N_8077,N_2546,N_372);
or U8078 (N_8078,N_4025,N_1629);
nor U8079 (N_8079,N_1482,N_4156);
nor U8080 (N_8080,N_5604,N_4190);
nor U8081 (N_8081,N_5567,N_1898);
nand U8082 (N_8082,N_2957,N_641);
and U8083 (N_8083,N_3017,N_5680);
nor U8084 (N_8084,N_5021,N_3050);
nor U8085 (N_8085,N_2899,N_4797);
nand U8086 (N_8086,N_3089,N_4623);
or U8087 (N_8087,N_4480,N_2761);
or U8088 (N_8088,N_2468,N_5760);
nor U8089 (N_8089,N_5366,N_4364);
nand U8090 (N_8090,N_5749,N_981);
or U8091 (N_8091,N_1846,N_3399);
nor U8092 (N_8092,N_2280,N_1681);
and U8093 (N_8093,N_5225,N_2543);
nor U8094 (N_8094,N_4262,N_3573);
or U8095 (N_8095,N_817,N_4995);
and U8096 (N_8096,N_3301,N_2488);
and U8097 (N_8097,N_724,N_5684);
nand U8098 (N_8098,N_2714,N_4002);
nor U8099 (N_8099,N_619,N_2816);
or U8100 (N_8100,N_3927,N_4205);
or U8101 (N_8101,N_5012,N_5241);
or U8102 (N_8102,N_1240,N_6216);
nor U8103 (N_8103,N_3146,N_1029);
nand U8104 (N_8104,N_5615,N_2246);
and U8105 (N_8105,N_1955,N_4529);
or U8106 (N_8106,N_1571,N_3159);
nand U8107 (N_8107,N_1776,N_2288);
nor U8108 (N_8108,N_1058,N_6039);
or U8109 (N_8109,N_1380,N_627);
and U8110 (N_8110,N_5311,N_5320);
and U8111 (N_8111,N_5264,N_6191);
and U8112 (N_8112,N_349,N_3164);
and U8113 (N_8113,N_6129,N_1932);
nor U8114 (N_8114,N_5921,N_5936);
nand U8115 (N_8115,N_3709,N_1929);
or U8116 (N_8116,N_6051,N_3526);
or U8117 (N_8117,N_3176,N_2321);
nand U8118 (N_8118,N_4446,N_3450);
or U8119 (N_8119,N_1330,N_1651);
nand U8120 (N_8120,N_593,N_4540);
nor U8121 (N_8121,N_6218,N_2684);
and U8122 (N_8122,N_1553,N_4147);
or U8123 (N_8123,N_3629,N_4208);
nor U8124 (N_8124,N_4173,N_3853);
and U8125 (N_8125,N_5592,N_5591);
nor U8126 (N_8126,N_3085,N_3621);
nor U8127 (N_8127,N_2919,N_5578);
or U8128 (N_8128,N_5802,N_3512);
and U8129 (N_8129,N_3404,N_1222);
or U8130 (N_8130,N_1216,N_3643);
nand U8131 (N_8131,N_4827,N_1208);
nor U8132 (N_8132,N_5019,N_5127);
and U8133 (N_8133,N_3637,N_3069);
nand U8134 (N_8134,N_848,N_2713);
or U8135 (N_8135,N_5014,N_6108);
or U8136 (N_8136,N_5015,N_3010);
nand U8137 (N_8137,N_4786,N_976);
nor U8138 (N_8138,N_2388,N_2200);
nand U8139 (N_8139,N_4120,N_3419);
nor U8140 (N_8140,N_2504,N_435);
and U8141 (N_8141,N_2789,N_4407);
nand U8142 (N_8142,N_715,N_2218);
nor U8143 (N_8143,N_5425,N_826);
nand U8144 (N_8144,N_886,N_1271);
nand U8145 (N_8145,N_942,N_5067);
nor U8146 (N_8146,N_479,N_5066);
and U8147 (N_8147,N_5286,N_4126);
or U8148 (N_8148,N_2213,N_1984);
and U8149 (N_8149,N_1667,N_6013);
nor U8150 (N_8150,N_5624,N_1987);
or U8151 (N_8151,N_5385,N_4219);
nand U8152 (N_8152,N_1853,N_2711);
nor U8153 (N_8153,N_1819,N_3261);
and U8154 (N_8154,N_5040,N_4071);
or U8155 (N_8155,N_4453,N_933);
nand U8156 (N_8156,N_1626,N_504);
nor U8157 (N_8157,N_4438,N_4916);
nand U8158 (N_8158,N_1165,N_4846);
nand U8159 (N_8159,N_3836,N_2513);
nand U8160 (N_8160,N_577,N_3502);
nand U8161 (N_8161,N_4599,N_6161);
and U8162 (N_8162,N_1110,N_720);
nand U8163 (N_8163,N_2620,N_5773);
nor U8164 (N_8164,N_4851,N_4401);
nor U8165 (N_8165,N_3615,N_1851);
and U8166 (N_8166,N_2065,N_3914);
nand U8167 (N_8167,N_5341,N_4284);
and U8168 (N_8168,N_2550,N_2610);
nor U8169 (N_8169,N_3105,N_3340);
nand U8170 (N_8170,N_5433,N_4612);
or U8171 (N_8171,N_4188,N_2697);
or U8172 (N_8172,N_36,N_3388);
nand U8173 (N_8173,N_1457,N_5270);
nor U8174 (N_8174,N_4167,N_6080);
and U8175 (N_8175,N_5403,N_3334);
nand U8176 (N_8176,N_4656,N_3219);
and U8177 (N_8177,N_4367,N_2574);
and U8178 (N_8178,N_2045,N_6003);
and U8179 (N_8179,N_5057,N_2937);
and U8180 (N_8180,N_940,N_3212);
or U8181 (N_8181,N_3488,N_1724);
and U8182 (N_8182,N_654,N_1390);
and U8183 (N_8183,N_1758,N_2156);
or U8184 (N_8184,N_1114,N_4253);
nand U8185 (N_8185,N_4796,N_5902);
and U8186 (N_8186,N_206,N_3687);
nor U8187 (N_8187,N_6081,N_1143);
or U8188 (N_8188,N_3911,N_3614);
nor U8189 (N_8189,N_4444,N_5146);
nor U8190 (N_8190,N_1951,N_5550);
nand U8191 (N_8191,N_2560,N_2732);
nand U8192 (N_8192,N_4763,N_4204);
nor U8193 (N_8193,N_98,N_3311);
or U8194 (N_8194,N_3433,N_3846);
nor U8195 (N_8195,N_5003,N_3834);
nand U8196 (N_8196,N_2549,N_5729);
and U8197 (N_8197,N_632,N_1121);
or U8198 (N_8198,N_816,N_1471);
nand U8199 (N_8199,N_2144,N_2170);
nand U8200 (N_8200,N_2939,N_1198);
nor U8201 (N_8201,N_1871,N_5);
or U8202 (N_8202,N_1530,N_2235);
nand U8203 (N_8203,N_4508,N_2464);
xnor U8204 (N_8204,N_1583,N_2980);
and U8205 (N_8205,N_5914,N_2400);
nor U8206 (N_8206,N_2566,N_5168);
nand U8207 (N_8207,N_5981,N_1485);
nor U8208 (N_8208,N_5248,N_3973);
nand U8209 (N_8209,N_575,N_4551);
or U8210 (N_8210,N_4735,N_6125);
nor U8211 (N_8211,N_2995,N_3389);
and U8212 (N_8212,N_5239,N_2463);
or U8213 (N_8213,N_5576,N_1648);
and U8214 (N_8214,N_3361,N_4399);
nand U8215 (N_8215,N_1015,N_2573);
xor U8216 (N_8216,N_1063,N_918);
nor U8217 (N_8217,N_3489,N_4908);
and U8218 (N_8218,N_849,N_501);
or U8219 (N_8219,N_825,N_6101);
and U8220 (N_8220,N_4316,N_3115);
or U8221 (N_8221,N_2342,N_4047);
or U8222 (N_8222,N_3035,N_2716);
nand U8223 (N_8223,N_2458,N_4470);
xor U8224 (N_8224,N_5285,N_2600);
nor U8225 (N_8225,N_5723,N_1918);
nand U8226 (N_8226,N_3542,N_2360);
nand U8227 (N_8227,N_5249,N_5255);
nand U8228 (N_8228,N_156,N_591);
nand U8229 (N_8229,N_4679,N_719);
or U8230 (N_8230,N_2672,N_202);
nor U8231 (N_8231,N_5930,N_777);
or U8232 (N_8232,N_5457,N_1329);
and U8233 (N_8233,N_5151,N_2525);
or U8234 (N_8234,N_1564,N_4032);
and U8235 (N_8235,N_934,N_5943);
or U8236 (N_8236,N_4780,N_5080);
and U8237 (N_8237,N_4943,N_1850);
nor U8238 (N_8238,N_3538,N_2707);
nand U8239 (N_8239,N_1447,N_649);
nand U8240 (N_8240,N_1917,N_4616);
xnor U8241 (N_8241,N_4584,N_803);
nor U8242 (N_8242,N_5746,N_117);
or U8243 (N_8243,N_5809,N_4468);
nor U8244 (N_8244,N_1732,N_6124);
nand U8245 (N_8245,N_5409,N_1767);
or U8246 (N_8246,N_4337,N_5362);
and U8247 (N_8247,N_454,N_5197);
or U8248 (N_8248,N_6047,N_433);
and U8249 (N_8249,N_1601,N_2322);
or U8250 (N_8250,N_2108,N_5427);
nand U8251 (N_8251,N_4474,N_1287);
nor U8252 (N_8252,N_3730,N_1737);
and U8253 (N_8253,N_756,N_3268);
nor U8254 (N_8254,N_3963,N_4545);
or U8255 (N_8255,N_4228,N_1550);
nand U8256 (N_8256,N_2715,N_1982);
and U8257 (N_8257,N_224,N_2470);
nand U8258 (N_8258,N_2793,N_2921);
or U8259 (N_8259,N_4300,N_8);
or U8260 (N_8260,N_3503,N_3505);
and U8261 (N_8261,N_2089,N_227);
nand U8262 (N_8262,N_3086,N_4131);
nor U8263 (N_8263,N_6153,N_2571);
nand U8264 (N_8264,N_268,N_597);
nand U8265 (N_8265,N_2655,N_3617);
nor U8266 (N_8266,N_6163,N_1092);
or U8267 (N_8267,N_1340,N_3084);
nor U8268 (N_8268,N_1675,N_2534);
or U8269 (N_8269,N_4338,N_626);
or U8270 (N_8270,N_5566,N_52);
nor U8271 (N_8271,N_4771,N_3955);
and U8272 (N_8272,N_51,N_4112);
or U8273 (N_8273,N_3785,N_4283);
nand U8274 (N_8274,N_5189,N_2833);
or U8275 (N_8275,N_3782,N_1614);
and U8276 (N_8276,N_3766,N_4016);
or U8277 (N_8277,N_2334,N_1902);
nand U8278 (N_8278,N_2410,N_3383);
and U8279 (N_8279,N_125,N_6202);
nor U8280 (N_8280,N_6167,N_2562);
and U8281 (N_8281,N_3835,N_2614);
and U8282 (N_8282,N_2367,N_3992);
nor U8283 (N_8283,N_1649,N_5058);
nor U8284 (N_8284,N_2238,N_2591);
or U8285 (N_8285,N_3484,N_4816);
nand U8286 (N_8286,N_837,N_1032);
or U8287 (N_8287,N_3350,N_235);
and U8288 (N_8288,N_4658,N_6238);
and U8289 (N_8289,N_1915,N_1625);
and U8290 (N_8290,N_1839,N_5415);
nand U8291 (N_8291,N_1925,N_2116);
nand U8292 (N_8292,N_4740,N_5101);
nor U8293 (N_8293,N_1847,N_4878);
nor U8294 (N_8294,N_3254,N_16);
and U8295 (N_8295,N_568,N_4031);
or U8296 (N_8296,N_4937,N_913);
and U8297 (N_8297,N_5558,N_3294);
or U8298 (N_8298,N_4021,N_861);
nor U8299 (N_8299,N_1106,N_5038);
nor U8300 (N_8300,N_5228,N_3875);
or U8301 (N_8301,N_3728,N_1961);
and U8302 (N_8302,N_5452,N_729);
or U8303 (N_8303,N_2104,N_6144);
or U8304 (N_8304,N_5473,N_6193);
nor U8305 (N_8305,N_2176,N_3480);
or U8306 (N_8306,N_847,N_5884);
nand U8307 (N_8307,N_617,N_1717);
and U8308 (N_8308,N_3187,N_2530);
or U8309 (N_8309,N_5874,N_5027);
nor U8310 (N_8310,N_1349,N_5859);
nand U8311 (N_8311,N_955,N_4302);
and U8312 (N_8312,N_5856,N_15);
and U8313 (N_8313,N_1942,N_2933);
nand U8314 (N_8314,N_1475,N_2232);
or U8315 (N_8315,N_2503,N_1647);
and U8316 (N_8316,N_4229,N_1307);
nor U8317 (N_8317,N_4892,N_2349);
and U8318 (N_8318,N_1022,N_4587);
nand U8319 (N_8319,N_1897,N_4751);
or U8320 (N_8320,N_4258,N_2420);
nor U8321 (N_8321,N_3984,N_3221);
nor U8322 (N_8322,N_3165,N_1738);
nor U8323 (N_8323,N_1812,N_5326);
or U8324 (N_8324,N_1952,N_4186);
nand U8325 (N_8325,N_2724,N_1525);
or U8326 (N_8326,N_3759,N_831);
and U8327 (N_8327,N_3109,N_2706);
or U8328 (N_8328,N_4075,N_3274);
nand U8329 (N_8329,N_4289,N_1484);
nor U8330 (N_8330,N_5702,N_2314);
nand U8331 (N_8331,N_4941,N_2259);
and U8332 (N_8332,N_3209,N_2118);
or U8333 (N_8333,N_376,N_3396);
and U8334 (N_8334,N_4533,N_1605);
nor U8335 (N_8335,N_3444,N_2953);
nor U8336 (N_8336,N_4683,N_2124);
nor U8337 (N_8337,N_5511,N_5180);
nand U8338 (N_8338,N_21,N_2039);
or U8339 (N_8339,N_888,N_2553);
or U8340 (N_8340,N_4425,N_5135);
nand U8341 (N_8341,N_4562,N_553);
and U8342 (N_8342,N_5304,N_123);
nor U8343 (N_8343,N_160,N_3613);
and U8344 (N_8344,N_2479,N_3590);
nand U8345 (N_8345,N_5082,N_6078);
nand U8346 (N_8346,N_3049,N_3482);
or U8347 (N_8347,N_5376,N_1937);
or U8348 (N_8348,N_2505,N_4441);
nor U8349 (N_8349,N_1276,N_1685);
or U8350 (N_8350,N_843,N_4242);
and U8351 (N_8351,N_1565,N_1207);
nor U8352 (N_8352,N_6130,N_2242);
nand U8353 (N_8353,N_520,N_872);
nor U8354 (N_8354,N_96,N_6126);
nor U8355 (N_8355,N_1050,N_4124);
and U8356 (N_8356,N_2722,N_1081);
or U8357 (N_8357,N_2903,N_1662);
or U8358 (N_8358,N_2277,N_497);
nand U8359 (N_8359,N_1448,N_3369);
nand U8360 (N_8360,N_168,N_186);
nor U8361 (N_8361,N_3276,N_4754);
and U8362 (N_8362,N_4506,N_1436);
nand U8363 (N_8363,N_346,N_4223);
nand U8364 (N_8364,N_3896,N_495);
nand U8365 (N_8365,N_5475,N_2586);
nor U8366 (N_8366,N_4944,N_984);
nand U8367 (N_8367,N_4779,N_3252);
nand U8368 (N_8368,N_526,N_1117);
and U8369 (N_8369,N_384,N_3897);
nor U8370 (N_8370,N_3755,N_56);
and U8371 (N_8371,N_1582,N_2076);
nand U8372 (N_8372,N_3111,N_4549);
or U8373 (N_8373,N_4543,N_1799);
nor U8374 (N_8374,N_2087,N_603);
or U8375 (N_8375,N_4200,N_4673);
nor U8376 (N_8376,N_4274,N_64);
nor U8377 (N_8377,N_57,N_5423);
and U8378 (N_8378,N_4576,N_2613);
and U8379 (N_8379,N_4481,N_3699);
and U8380 (N_8380,N_2617,N_320);
nor U8381 (N_8381,N_5721,N_5732);
or U8382 (N_8382,N_2187,N_6036);
and U8383 (N_8383,N_5693,N_3645);
and U8384 (N_8384,N_2961,N_5434);
or U8385 (N_8385,N_767,N_759);
or U8386 (N_8386,N_4286,N_4082);
and U8387 (N_8387,N_505,N_2382);
and U8388 (N_8388,N_968,N_5965);
or U8389 (N_8389,N_5160,N_1295);
nand U8390 (N_8390,N_5025,N_4635);
or U8391 (N_8391,N_3478,N_1168);
and U8392 (N_8392,N_3380,N_1140);
nor U8393 (N_8393,N_2014,N_4630);
and U8394 (N_8394,N_3739,N_2824);
and U8395 (N_8395,N_4499,N_5132);
nand U8396 (N_8396,N_4690,N_1302);
nand U8397 (N_8397,N_5122,N_4909);
or U8398 (N_8398,N_3644,N_4570);
nor U8399 (N_8399,N_3893,N_6172);
nor U8400 (N_8400,N_4241,N_2959);
nor U8401 (N_8401,N_5950,N_5242);
and U8402 (N_8402,N_2666,N_5513);
or U8403 (N_8403,N_622,N_6235);
nor U8404 (N_8404,N_4617,N_1821);
or U8405 (N_8405,N_3905,N_3287);
nor U8406 (N_8406,N_1350,N_3295);
nor U8407 (N_8407,N_1137,N_1823);
nand U8408 (N_8408,N_4731,N_6067);
or U8409 (N_8409,N_3173,N_993);
and U8410 (N_8410,N_4997,N_569);
nor U8411 (N_8411,N_4362,N_4756);
nand U8412 (N_8412,N_2873,N_1397);
or U8413 (N_8413,N_3178,N_3890);
or U8414 (N_8414,N_243,N_573);
nand U8415 (N_8415,N_199,N_317);
nor U8416 (N_8416,N_2527,N_240);
nor U8417 (N_8417,N_4703,N_1069);
nand U8418 (N_8418,N_2612,N_3310);
and U8419 (N_8419,N_4629,N_882);
xnor U8420 (N_8420,N_325,N_5358);
or U8421 (N_8421,N_174,N_2062);
or U8422 (N_8422,N_420,N_809);
nor U8423 (N_8423,N_1994,N_2161);
and U8424 (N_8424,N_3811,N_5356);
and U8425 (N_8425,N_2375,N_3670);
and U8426 (N_8426,N_4052,N_562);
or U8427 (N_8427,N_1030,N_1027);
and U8428 (N_8428,N_6062,N_3608);
nand U8429 (N_8429,N_3280,N_428);
nand U8430 (N_8430,N_838,N_2234);
nand U8431 (N_8431,N_2547,N_423);
nand U8432 (N_8432,N_1716,N_1736);
nand U8433 (N_8433,N_2608,N_111);
and U8434 (N_8434,N_4651,N_4456);
and U8435 (N_8435,N_4496,N_4307);
and U8436 (N_8436,N_3494,N_2193);
or U8437 (N_8437,N_5900,N_3098);
nor U8438 (N_8438,N_5894,N_1405);
nor U8439 (N_8439,N_3902,N_2670);
nor U8440 (N_8440,N_1928,N_4452);
or U8441 (N_8441,N_2029,N_6152);
nor U8442 (N_8442,N_930,N_1835);
or U8443 (N_8443,N_4249,N_2131);
and U8444 (N_8444,N_5569,N_858);
nor U8445 (N_8445,N_355,N_3812);
nor U8446 (N_8446,N_2790,N_446);
nor U8447 (N_8447,N_2738,N_2598);
and U8448 (N_8448,N_3713,N_697);
or U8449 (N_8449,N_3483,N_2095);
or U8450 (N_8450,N_3545,N_3831);
and U8451 (N_8451,N_5421,N_3349);
nor U8452 (N_8452,N_2240,N_792);
and U8453 (N_8453,N_2524,N_1804);
nor U8454 (N_8454,N_3761,N_5483);
nand U8455 (N_8455,N_3203,N_5275);
nand U8456 (N_8456,N_337,N_2483);
or U8457 (N_8457,N_951,N_3716);
nand U8458 (N_8458,N_2814,N_1810);
and U8459 (N_8459,N_1587,N_5266);
nor U8460 (N_8460,N_2121,N_1706);
nor U8461 (N_8461,N_3877,N_2467);
and U8462 (N_8462,N_3663,N_1770);
nand U8463 (N_8463,N_4153,N_1404);
or U8464 (N_8464,N_1920,N_1906);
and U8465 (N_8465,N_3336,N_1893);
or U8466 (N_8466,N_733,N_3504);
nor U8467 (N_8467,N_2973,N_4933);
nand U8468 (N_8468,N_3292,N_3587);
nor U8469 (N_8469,N_4288,N_1185);
and U8470 (N_8470,N_5000,N_6203);
or U8471 (N_8471,N_2569,N_1017);
and U8472 (N_8472,N_1996,N_1003);
nor U8473 (N_8473,N_3005,N_3849);
nand U8474 (N_8474,N_4671,N_5533);
nand U8475 (N_8475,N_5456,N_6151);
nand U8476 (N_8476,N_5195,N_2485);
nand U8477 (N_8477,N_4465,N_4294);
or U8478 (N_8478,N_2318,N_2183);
nand U8479 (N_8479,N_2415,N_2946);
or U8480 (N_8480,N_4489,N_2892);
or U8481 (N_8481,N_2405,N_94);
or U8482 (N_8482,N_5880,N_3510);
nand U8483 (N_8483,N_5321,N_548);
or U8484 (N_8484,N_4601,N_4766);
nor U8485 (N_8485,N_6188,N_2159);
and U8486 (N_8486,N_1948,N_3335);
and U8487 (N_8487,N_3062,N_1360);
nand U8488 (N_8488,N_4585,N_4116);
or U8489 (N_8489,N_3684,N_594);
or U8490 (N_8490,N_5776,N_5209);
or U8491 (N_8491,N_1977,N_1023);
nand U8492 (N_8492,N_5174,N_2332);
nor U8493 (N_8493,N_1103,N_5391);
or U8494 (N_8494,N_267,N_5677);
and U8495 (N_8495,N_5787,N_1033);
or U8496 (N_8496,N_6077,N_2996);
and U8497 (N_8497,N_3915,N_121);
or U8498 (N_8498,N_4521,N_4459);
or U8499 (N_8499,N_1699,N_4175);
and U8500 (N_8500,N_892,N_4875);
nor U8501 (N_8501,N_2727,N_5065);
nand U8502 (N_8502,N_1045,N_1748);
or U8503 (N_8503,N_1750,N_2459);
nand U8504 (N_8504,N_5244,N_628);
nand U8505 (N_8505,N_2431,N_2914);
and U8506 (N_8506,N_4319,N_4164);
or U8507 (N_8507,N_547,N_5734);
or U8508 (N_8508,N_6072,N_6240);
and U8509 (N_8509,N_920,N_2637);
nor U8510 (N_8510,N_6090,N_89);
nand U8511 (N_8511,N_339,N_6007);
or U8512 (N_8512,N_532,N_1899);
and U8513 (N_8513,N_4807,N_3243);
nor U8514 (N_8514,N_6146,N_2113);
or U8515 (N_8515,N_5440,N_6005);
nor U8516 (N_8516,N_899,N_4575);
nand U8517 (N_8517,N_5681,N_3402);
or U8518 (N_8518,N_5130,N_5867);
and U8519 (N_8519,N_578,N_4701);
and U8520 (N_8520,N_6000,N_3241);
nand U8521 (N_8521,N_3541,N_2347);
nand U8522 (N_8522,N_4072,N_3601);
or U8523 (N_8523,N_4812,N_5536);
nor U8524 (N_8524,N_3347,N_722);
nand U8525 (N_8525,N_3095,N_3565);
and U8526 (N_8526,N_4544,N_5818);
nand U8527 (N_8527,N_5815,N_5155);
or U8528 (N_8528,N_1149,N_5156);
and U8529 (N_8529,N_3155,N_1013);
nor U8530 (N_8530,N_2756,N_2358);
nor U8531 (N_8531,N_4609,N_4729);
nand U8532 (N_8532,N_5167,N_5182);
and U8533 (N_8533,N_4848,N_6094);
nor U8534 (N_8534,N_271,N_3045);
nand U8535 (N_8535,N_5895,N_2855);
nor U8536 (N_8536,N_3506,N_1646);
and U8537 (N_8537,N_2299,N_3249);
or U8538 (N_8538,N_213,N_1610);
and U8539 (N_8539,N_2709,N_5372);
and U8540 (N_8540,N_1061,N_41);
nor U8541 (N_8541,N_5295,N_2343);
nor U8542 (N_8542,N_5752,N_1278);
nor U8543 (N_8543,N_5833,N_704);
nor U8544 (N_8544,N_5933,N_2384);
and U8545 (N_8545,N_2827,N_1894);
nand U8546 (N_8546,N_426,N_65);
nand U8547 (N_8547,N_2128,N_2201);
nand U8548 (N_8548,N_1608,N_2443);
nand U8549 (N_8549,N_4461,N_4440);
nor U8550 (N_8550,N_4950,N_5004);
or U8551 (N_8551,N_829,N_2624);
nor U8552 (N_8552,N_5968,N_5623);
and U8553 (N_8553,N_276,N_29);
or U8554 (N_8554,N_3438,N_3841);
nor U8555 (N_8555,N_1607,N_1282);
and U8556 (N_8556,N_6035,N_3632);
nor U8557 (N_8557,N_4439,N_4550);
or U8558 (N_8558,N_599,N_5240);
nand U8559 (N_8559,N_4015,N_1464);
nor U8560 (N_8560,N_631,N_2172);
nor U8561 (N_8561,N_1362,N_5375);
nor U8562 (N_8562,N_6034,N_2565);
nor U8563 (N_8563,N_3032,N_2518);
xor U8564 (N_8564,N_5949,N_1161);
or U8565 (N_8565,N_4964,N_3186);
nor U8566 (N_8566,N_2202,N_502);
nor U8567 (N_8567,N_4301,N_2474);
and U8568 (N_8568,N_1462,N_170);
or U8569 (N_8569,N_4172,N_2220);
and U8570 (N_8570,N_2270,N_3999);
nor U8571 (N_8571,N_862,N_2618);
nand U8572 (N_8572,N_2887,N_4);
and U8573 (N_8573,N_5367,N_1783);
and U8574 (N_8574,N_4062,N_1186);
nor U8575 (N_8575,N_5116,N_3207);
nand U8576 (N_8576,N_1979,N_1166);
and U8577 (N_8577,N_5199,N_2064);
and U8578 (N_8578,N_3027,N_3577);
or U8579 (N_8579,N_4620,N_3726);
nor U8580 (N_8580,N_3245,N_6140);
or U8581 (N_8581,N_6111,N_531);
xnor U8582 (N_8582,N_2918,N_5541);
nand U8583 (N_8583,N_336,N_3515);
nand U8584 (N_8584,N_6117,N_5384);
nor U8585 (N_8585,N_2587,N_5649);
nand U8586 (N_8586,N_2656,N_5573);
nand U8587 (N_8587,N_5935,N_2245);
nor U8588 (N_8588,N_4684,N_380);
and U8589 (N_8589,N_4885,N_1870);
or U8590 (N_8590,N_927,N_5629);
nor U8591 (N_8591,N_5010,N_183);
and U8592 (N_8592,N_194,N_4886);
nor U8593 (N_8593,N_5632,N_540);
nor U8594 (N_8594,N_1190,N_2805);
and U8595 (N_8595,N_2705,N_2038);
and U8596 (N_8596,N_3575,N_1939);
nand U8597 (N_8597,N_3674,N_3525);
nand U8598 (N_8598,N_2932,N_4411);
or U8599 (N_8599,N_1903,N_2649);
and U8600 (N_8600,N_4949,N_266);
nor U8601 (N_8601,N_2779,N_1465);
nand U8602 (N_8602,N_54,N_67);
nand U8603 (N_8603,N_1572,N_1642);
or U8604 (N_8604,N_3789,N_5917);
and U8605 (N_8605,N_5518,N_3894);
and U8606 (N_8606,N_5230,N_1686);
and U8607 (N_8607,N_3771,N_3116);
nor U8608 (N_8608,N_4563,N_2774);
nand U8609 (N_8609,N_4573,N_5877);
or U8610 (N_8610,N_92,N_2748);
and U8611 (N_8611,N_1371,N_4993);
or U8612 (N_8612,N_6236,N_924);
and U8613 (N_8613,N_716,N_3798);
nand U8614 (N_8614,N_1416,N_2552);
and U8615 (N_8615,N_6102,N_896);
nor U8616 (N_8616,N_3158,N_1658);
and U8617 (N_8617,N_3521,N_5812);
nor U8618 (N_8618,N_3838,N_3013);
and U8619 (N_8619,N_298,N_1089);
nor U8620 (N_8620,N_814,N_5281);
or U8621 (N_8621,N_5940,N_3244);
nor U8622 (N_8622,N_1234,N_1714);
or U8623 (N_8623,N_169,N_2060);
nand U8624 (N_8624,N_1365,N_791);
and U8625 (N_8625,N_413,N_3445);
nand U8626 (N_8626,N_5307,N_1263);
or U8627 (N_8627,N_4149,N_2439);
nor U8628 (N_8628,N_159,N_713);
nand U8629 (N_8629,N_5324,N_5685);
and U8630 (N_8630,N_623,N_63);
nand U8631 (N_8631,N_1133,N_4794);
nand U8632 (N_8632,N_1882,N_737);
and U8633 (N_8633,N_6033,N_5092);
nor U8634 (N_8634,N_0,N_333);
nand U8635 (N_8635,N_1754,N_1481);
xor U8636 (N_8636,N_2168,N_4343);
or U8637 (N_8637,N_2214,N_5454);
nor U8638 (N_8638,N_1720,N_3408);
and U8639 (N_8639,N_5530,N_5368);
or U8640 (N_8640,N_3226,N_2556);
nand U8641 (N_8641,N_5611,N_4856);
nand U8642 (N_8642,N_5666,N_774);
or U8643 (N_8643,N_4638,N_444);
nor U8644 (N_8644,N_5379,N_3871);
nor U8645 (N_8645,N_3256,N_2680);
or U8646 (N_8646,N_2319,N_5009);
and U8647 (N_8647,N_2825,N_5467);
or U8648 (N_8648,N_1331,N_558);
and U8649 (N_8649,N_410,N_5363);
or U8650 (N_8650,N_2164,N_4986);
nor U8651 (N_8651,N_5024,N_5688);
and U8652 (N_8652,N_648,N_3359);
nor U8653 (N_8653,N_1726,N_1101);
and U8654 (N_8654,N_5557,N_1080);
and U8655 (N_8655,N_3315,N_4096);
nor U8656 (N_8656,N_2829,N_3742);
nand U8657 (N_8657,N_3420,N_744);
nor U8658 (N_8658,N_5284,N_1458);
and U8659 (N_8659,N_5766,N_4732);
and U8660 (N_8660,N_2659,N_512);
and U8661 (N_8661,N_4590,N_979);
and U8662 (N_8662,N_2667,N_5301);
nor U8663 (N_8663,N_4051,N_703);
nand U8664 (N_8664,N_3641,N_6023);
or U8665 (N_8665,N_3885,N_4179);
nand U8666 (N_8666,N_2599,N_2823);
nand U8667 (N_8667,N_4789,N_2590);
nand U8668 (N_8668,N_677,N_2522);
nand U8669 (N_8669,N_4451,N_277);
nand U8670 (N_8670,N_1914,N_3263);
and U8671 (N_8671,N_4251,N_4746);
or U8672 (N_8672,N_1181,N_546);
or U8673 (N_8673,N_319,N_171);
nor U8674 (N_8674,N_5619,N_2041);
nor U8675 (N_8675,N_1211,N_414);
xor U8676 (N_8676,N_819,N_198);
or U8677 (N_8677,N_3126,N_5005);
or U8678 (N_8678,N_870,N_221);
nand U8679 (N_8679,N_237,N_1250);
nor U8680 (N_8680,N_4643,N_1463);
nand U8681 (N_8681,N_1055,N_2184);
nor U8682 (N_8682,N_2501,N_269);
or U8683 (N_8683,N_1723,N_3680);
and U8684 (N_8684,N_1188,N_4313);
nor U8685 (N_8685,N_4485,N_4194);
or U8686 (N_8686,N_3559,N_1875);
and U8687 (N_8687,N_1815,N_3279);
and U8688 (N_8688,N_1534,N_3934);
nand U8689 (N_8689,N_360,N_3507);
or U8690 (N_8690,N_1000,N_2341);
nand U8691 (N_8691,N_4437,N_4719);
or U8692 (N_8692,N_5125,N_1687);
nand U8693 (N_8693,N_4376,N_2576);
nand U8694 (N_8694,N_2902,N_5798);
nor U8695 (N_8695,N_1848,N_4139);
and U8696 (N_8696,N_6127,N_4280);
or U8697 (N_8697,N_4305,N_1123);
or U8698 (N_8698,N_6075,N_150);
nor U8699 (N_8699,N_2539,N_587);
nand U8700 (N_8700,N_2011,N_2323);
nor U8701 (N_8701,N_3932,N_1378);
or U8702 (N_8702,N_580,N_4705);
or U8703 (N_8703,N_371,N_1372);
nand U8704 (N_8704,N_4901,N_5046);
nand U8705 (N_8705,N_55,N_6164);
nor U8706 (N_8706,N_4006,N_5546);
nand U8707 (N_8707,N_3661,N_5724);
nor U8708 (N_8708,N_3997,N_4980);
nor U8709 (N_8709,N_1072,N_5829);
nor U8710 (N_8710,N_3579,N_5780);
or U8711 (N_8711,N_6143,N_1808);
nand U8712 (N_8712,N_576,N_5991);
and U8713 (N_8713,N_2970,N_4121);
nand U8714 (N_8714,N_4320,N_3522);
nand U8715 (N_8715,N_3731,N_4845);
nor U8716 (N_8716,N_2107,N_1494);
nor U8717 (N_8717,N_4708,N_175);
nor U8718 (N_8718,N_5735,N_5618);
or U8719 (N_8719,N_586,N_306);
or U8720 (N_8720,N_1886,N_5369);
nor U8721 (N_8721,N_5758,N_1609);
nand U8722 (N_8722,N_551,N_1241);
nand U8723 (N_8723,N_798,N_1824);
nand U8724 (N_8724,N_3702,N_3048);
nor U8725 (N_8725,N_1470,N_4996);
or U8726 (N_8726,N_1887,N_4621);
and U8727 (N_8727,N_1617,N_3790);
and U8728 (N_8728,N_5318,N_3372);
and U8729 (N_8729,N_4449,N_1395);
nand U8730 (N_8730,N_969,N_2101);
or U8731 (N_8731,N_222,N_1432);
nor U8732 (N_8732,N_5990,N_5121);
nor U8733 (N_8733,N_2988,N_44);
nor U8734 (N_8734,N_1277,N_5652);
nand U8735 (N_8735,N_1673,N_3171);
and U8736 (N_8736,N_5964,N_2979);
or U8737 (N_8737,N_1956,N_3368);
nand U8738 (N_8738,N_5979,N_5811);
and U8739 (N_8739,N_4064,N_4709);
or U8740 (N_8740,N_3,N_1708);
and U8741 (N_8741,N_4310,N_3554);
xnor U8742 (N_8742,N_6073,N_3916);
and U8743 (N_8743,N_457,N_6121);
nand U8744 (N_8744,N_3180,N_3104);
nand U8745 (N_8745,N_263,N_5008);
nor U8746 (N_8746,N_1247,N_636);
nand U8747 (N_8747,N_1279,N_126);
or U8748 (N_8748,N_4776,N_439);
and U8749 (N_8749,N_1500,N_260);
or U8750 (N_8750,N_1703,N_1704);
or U8751 (N_8751,N_3805,N_5858);
or U8752 (N_8752,N_1379,N_2883);
or U8753 (N_8753,N_5498,N_2248);
nor U8754 (N_8754,N_2808,N_5641);
and U8755 (N_8755,N_6026,N_534);
nor U8756 (N_8756,N_739,N_5534);
nor U8757 (N_8757,N_5192,N_5089);
and U8758 (N_8758,N_6010,N_162);
or U8759 (N_8759,N_1866,N_3583);
nand U8760 (N_8760,N_5794,N_5768);
nand U8761 (N_8761,N_4331,N_302);
and U8762 (N_8762,N_3735,N_5451);
nor U8763 (N_8763,N_975,N_5448);
or U8764 (N_8764,N_2090,N_5259);
and U8765 (N_8765,N_891,N_5276);
or U8766 (N_8766,N_869,N_1798);
and U8767 (N_8767,N_4211,N_4160);
nand U8768 (N_8768,N_4677,N_4936);
nand U8769 (N_8769,N_5100,N_3296);
nor U8770 (N_8770,N_2354,N_1413);
nor U8771 (N_8771,N_5490,N_4143);
and U8772 (N_8772,N_3544,N_5408);
nand U8773 (N_8773,N_6179,N_5064);
and U8774 (N_8774,N_3557,N_1992);
or U8775 (N_8775,N_4682,N_5340);
or U8776 (N_8776,N_5741,N_4066);
and U8777 (N_8777,N_71,N_2857);
nand U8778 (N_8778,N_2862,N_3729);
nand U8779 (N_8779,N_780,N_5044);
nor U8780 (N_8780,N_2286,N_1158);
or U8781 (N_8781,N_1197,N_5956);
nand U8782 (N_8782,N_5370,N_3360);
and U8783 (N_8783,N_4994,N_683);
nor U8784 (N_8784,N_778,N_2623);
and U8785 (N_8785,N_3466,N_2685);
nand U8786 (N_8786,N_5861,N_2851);
or U8787 (N_8787,N_2185,N_1303);
and U8788 (N_8788,N_5549,N_2702);
or U8789 (N_8789,N_987,N_1224);
and U8790 (N_8790,N_4415,N_5313);
nor U8791 (N_8791,N_3839,N_1645);
nand U8792 (N_8792,N_2763,N_2631);
and U8793 (N_8793,N_1523,N_4315);
and U8794 (N_8794,N_1885,N_3901);
and U8795 (N_8795,N_2831,N_212);
or U8796 (N_8796,N_5378,N_2138);
and U8797 (N_8797,N_379,N_5258);
or U8798 (N_8798,N_6157,N_2422);
and U8799 (N_8799,N_5898,N_1860);
nor U8800 (N_8800,N_3980,N_5140);
nor U8801 (N_8801,N_4187,N_1852);
nand U8802 (N_8802,N_6079,N_5302);
or U8803 (N_8803,N_220,N_6133);
nand U8804 (N_8804,N_1746,N_2457);
or U8805 (N_8805,N_3400,N_389);
nor U8806 (N_8806,N_4945,N_5233);
and U8807 (N_8807,N_2247,N_5309);
nand U8808 (N_8808,N_2755,N_3951);
and U8809 (N_8809,N_5523,N_1415);
or U8810 (N_8810,N_3852,N_5865);
and U8811 (N_8811,N_4569,N_329);
and U8812 (N_8812,N_1088,N_5154);
nor U8813 (N_8813,N_2967,N_834);
nand U8814 (N_8814,N_815,N_772);
nor U8815 (N_8815,N_1796,N_3569);
or U8816 (N_8816,N_1127,N_463);
nand U8817 (N_8817,N_3734,N_3657);
nor U8818 (N_8818,N_2455,N_3769);
and U8819 (N_8819,N_3034,N_2674);
or U8820 (N_8820,N_4548,N_5181);
and U8821 (N_8821,N_196,N_1916);
and U8822 (N_8822,N_1321,N_5272);
nand U8823 (N_8823,N_5824,N_1338);
or U8824 (N_8824,N_4350,N_3074);
nand U8825 (N_8825,N_180,N_3752);
and U8826 (N_8826,N_3421,N_601);
nand U8827 (N_8827,N_2451,N_4646);
or U8828 (N_8828,N_2177,N_4947);
nor U8829 (N_8829,N_2687,N_5144);
nand U8830 (N_8830,N_3775,N_4558);
nand U8831 (N_8831,N_2111,N_2843);
nor U8832 (N_8832,N_5428,N_167);
nand U8833 (N_8833,N_2444,N_1538);
or U8834 (N_8834,N_6246,N_5691);
and U8835 (N_8835,N_3773,N_1969);
or U8836 (N_8836,N_1492,N_672);
nand U8837 (N_8837,N_3282,N_3753);
and U8838 (N_8838,N_5795,N_1666);
nand U8839 (N_8839,N_332,N_5234);
nand U8840 (N_8840,N_5608,N_4018);
and U8841 (N_8841,N_5445,N_4594);
nand U8842 (N_8842,N_748,N_5897);
nor U8843 (N_8843,N_3237,N_4822);
and U8844 (N_8844,N_3194,N_4648);
and U8845 (N_8845,N_3405,N_4272);
and U8846 (N_8846,N_6217,N_1910);
or U8847 (N_8847,N_2859,N_3720);
and U8848 (N_8848,N_6103,N_5579);
or U8849 (N_8849,N_2739,N_4830);
and U8850 (N_8850,N_962,N_4603);
and U8851 (N_8851,N_1581,N_3500);
nand U8852 (N_8852,N_3662,N_2024);
or U8853 (N_8853,N_6025,N_3228);
nand U8854 (N_8854,N_865,N_252);
nand U8855 (N_8855,N_2249,N_369);
nand U8856 (N_8856,N_3070,N_4614);
and U8857 (N_8857,N_5581,N_5468);
and U8858 (N_8858,N_972,N_6229);
nand U8859 (N_8859,N_6176,N_3809);
nor U8860 (N_8860,N_5298,N_6043);
or U8861 (N_8861,N_1435,N_2533);
or U8862 (N_8862,N_3403,N_4196);
nand U8863 (N_8863,N_5119,N_1670);
nand U8864 (N_8864,N_3107,N_1756);
nand U8865 (N_8865,N_6096,N_4091);
and U8866 (N_8866,N_4236,N_2180);
nor U8867 (N_8867,N_4895,N_3418);
nor U8868 (N_8868,N_81,N_2813);
nor U8869 (N_8869,N_1486,N_3651);
nor U8870 (N_8870,N_879,N_3855);
or U8871 (N_8871,N_5648,N_3908);
nand U8872 (N_8872,N_885,N_4418);
nand U8873 (N_8873,N_645,N_4354);
nand U8874 (N_8874,N_5453,N_2570);
or U8875 (N_8875,N_4693,N_5942);
nand U8876 (N_8876,N_249,N_808);
nand U8877 (N_8877,N_283,N_5479);
and U8878 (N_8878,N_4434,N_4268);
or U8879 (N_8879,N_4137,N_2211);
and U8880 (N_8880,N_690,N_5670);
or U8881 (N_8881,N_687,N_1591);
nor U8882 (N_8882,N_5528,N_1830);
and U8883 (N_8883,N_304,N_509);
and U8884 (N_8884,N_4721,N_4799);
or U8885 (N_8885,N_5620,N_3625);
nor U8886 (N_8886,N_1975,N_4511);
nand U8887 (N_8887,N_3188,N_181);
and U8888 (N_8888,N_3057,N_3312);
and U8889 (N_8889,N_1495,N_5715);
nor U8890 (N_8890,N_2432,N_93);
and U8891 (N_8891,N_5411,N_2773);
nor U8892 (N_8892,N_4348,N_2966);
nor U8893 (N_8893,N_3819,N_3443);
nor U8894 (N_8894,N_4462,N_4991);
and U8895 (N_8895,N_1580,N_1150);
and U8896 (N_8896,N_2182,N_4891);
or U8897 (N_8897,N_5287,N_3147);
nor U8898 (N_8898,N_3804,N_1950);
nand U8899 (N_8899,N_353,N_4267);
nor U8900 (N_8900,N_5682,N_6044);
nor U8901 (N_8901,N_2802,N_2780);
and U8902 (N_8902,N_4141,N_1734);
nor U8903 (N_8903,N_3650,N_3330);
nor U8904 (N_8904,N_1527,N_59);
or U8905 (N_8905,N_1622,N_4919);
nor U8906 (N_8906,N_3691,N_5056);
nor U8907 (N_8907,N_1926,N_3873);
nor U8908 (N_8908,N_4393,N_1352);
nand U8909 (N_8909,N_1529,N_6091);
or U8910 (N_8910,N_422,N_5022);
or U8911 (N_8911,N_205,N_3137);
nor U8912 (N_8912,N_3435,N_6187);
nor U8913 (N_8913,N_5133,N_500);
and U8914 (N_8914,N_5626,N_4290);
or U8915 (N_8915,N_1592,N_4783);
nand U8916 (N_8916,N_4270,N_1284);
nor U8917 (N_8917,N_6084,N_4029);
and U8918 (N_8918,N_141,N_4349);
and U8919 (N_8919,N_4098,N_4163);
nand U8920 (N_8920,N_4626,N_2639);
nor U8921 (N_8921,N_846,N_517);
nand U8922 (N_8922,N_4135,N_2962);
or U8923 (N_8923,N_5574,N_326);
or U8924 (N_8924,N_2253,N_90);
and U8925 (N_8925,N_4989,N_5846);
nand U8926 (N_8926,N_5873,N_3452);
and U8927 (N_8927,N_3882,N_5644);
and U8928 (N_8928,N_1514,N_2580);
nor U8929 (N_8929,N_3772,N_2364);
nand U8930 (N_8930,N_1874,N_4604);
or U8931 (N_8931,N_3477,N_5761);
nand U8932 (N_8932,N_4056,N_2309);
nand U8933 (N_8933,N_3253,N_637);
nand U8934 (N_8934,N_6201,N_5625);
and U8935 (N_8935,N_5178,N_2532);
nor U8936 (N_8936,N_4654,N_3120);
nand U8937 (N_8937,N_3976,N_499);
nor U8938 (N_8938,N_1232,N_4507);
nor U8939 (N_8939,N_4586,N_4125);
nor U8940 (N_8940,N_3140,N_3454);
or U8941 (N_8941,N_971,N_4925);
nand U8942 (N_8942,N_2404,N_2465);
nand U8943 (N_8943,N_4099,N_3054);
or U8944 (N_8944,N_289,N_3038);
nor U8945 (N_8945,N_630,N_5184);
nor U8946 (N_8946,N_3743,N_3266);
or U8947 (N_8947,N_3960,N_1834);
nor U8948 (N_8948,N_1177,N_3594);
nor U8949 (N_8949,N_4741,N_4664);
or U8950 (N_8950,N_4059,N_4429);
nor U8951 (N_8951,N_2221,N_407);
nand U8952 (N_8952,N_4598,N_2924);
and U8953 (N_8953,N_1904,N_5953);
nor U8954 (N_8954,N_5397,N_108);
or U8955 (N_8955,N_3354,N_4381);
nand U8956 (N_8956,N_4689,N_660);
and U8957 (N_8957,N_2594,N_2233);
nor U8958 (N_8958,N_2279,N_5621);
nand U8959 (N_8959,N_5344,N_4939);
nor U8960 (N_8960,N_718,N_3780);
nand U8961 (N_8961,N_5628,N_2766);
or U8962 (N_8962,N_6118,N_4627);
or U8963 (N_8963,N_2071,N_1074);
and U8964 (N_8964,N_5215,N_1191);
nand U8965 (N_8965,N_2004,N_115);
and U8966 (N_8966,N_3548,N_2224);
and U8967 (N_8967,N_4528,N_5843);
nand U8968 (N_8968,N_396,N_941);
or U8969 (N_8969,N_2018,N_5707);
nor U8970 (N_8970,N_515,N_3258);
nor U8971 (N_8971,N_903,N_2377);
and U8972 (N_8972,N_2227,N_1777);
nand U8973 (N_8973,N_1048,N_5172);
nor U8974 (N_8974,N_1179,N_852);
and U8975 (N_8975,N_1537,N_392);
nand U8976 (N_8976,N_1923,N_5002);
and U8977 (N_8977,N_1476,N_5954);
nand U8978 (N_8978,N_937,N_1175);
nand U8979 (N_8979,N_802,N_2799);
and U8980 (N_8980,N_995,N_4688);
or U8981 (N_8981,N_4522,N_2596);
and U8982 (N_8982,N_3058,N_4871);
nand U8983 (N_8983,N_5934,N_3561);
and U8984 (N_8984,N_4184,N_4842);
and U8985 (N_8985,N_1426,N_582);
xnor U8986 (N_8986,N_2313,N_31);
nor U8987 (N_8987,N_3051,N_4221);
nor U8988 (N_8988,N_2132,N_5660);
or U8989 (N_8989,N_1323,N_4128);
or U8990 (N_8990,N_5400,N_2093);
or U8991 (N_8991,N_4291,N_2067);
nand U8992 (N_8992,N_440,N_2203);
or U8993 (N_8993,N_1974,N_5289);
or U8994 (N_8994,N_2310,N_4408);
and U8995 (N_8995,N_3075,N_2745);
and U8996 (N_8996,N_916,N_2585);
or U8997 (N_8997,N_5505,N_5416);
and U8998 (N_8998,N_2701,N_4450);
nor U8999 (N_8999,N_3833,N_5700);
nand U9000 (N_9000,N_2199,N_1002);
nor U9001 (N_9001,N_2228,N_2784);
and U9002 (N_9002,N_2312,N_3763);
and U9003 (N_9003,N_1857,N_4304);
or U9004 (N_9004,N_5659,N_3078);
nor U9005 (N_9005,N_616,N_4834);
and U9006 (N_9006,N_5407,N_5654);
or U9007 (N_9007,N_4951,N_3832);
or U9008 (N_9008,N_516,N_5202);
nor U9009 (N_9009,N_4774,N_1765);
nor U9010 (N_9010,N_4107,N_5947);
and U9011 (N_9011,N_2427,N_2084);
or U9012 (N_9012,N_4197,N_149);
nor U9013 (N_9013,N_5237,N_2083);
or U9014 (N_9014,N_6150,N_2340);
nor U9015 (N_9015,N_4222,N_130);
and U9016 (N_9016,N_2344,N_2173);
nand U9017 (N_9017,N_2969,N_877);
and U9018 (N_9018,N_1131,N_3487);
and U9019 (N_9019,N_3037,N_1102);
and U9020 (N_9020,N_5464,N_5120);
nor U9021 (N_9021,N_1741,N_3149);
nand U9022 (N_9022,N_2381,N_665);
nor U9023 (N_9023,N_2500,N_4491);
nand U9024 (N_9024,N_278,N_5515);
and U9025 (N_9025,N_28,N_4095);
nand U9026 (N_9026,N_2677,N_2934);
nand U9027 (N_9027,N_2274,N_5343);
and U9028 (N_9028,N_3498,N_330);
or U9029 (N_9029,N_4676,N_3123);
nand U9030 (N_9030,N_4366,N_4896);
nor U9031 (N_9031,N_1933,N_4926);
nor U9032 (N_9032,N_1455,N_1744);
or U9033 (N_9033,N_1641,N_5545);
nand U9034 (N_9034,N_209,N_1239);
nand U9035 (N_9035,N_5447,N_822);
nor U9036 (N_9036,N_2433,N_404);
nor U9037 (N_9037,N_5087,N_667);
nand U9038 (N_9038,N_451,N_5441);
nand U9039 (N_9039,N_4034,N_1480);
nor U9040 (N_9040,N_723,N_2258);
and U9041 (N_9041,N_3144,N_2275);
and U9042 (N_9042,N_1566,N_4718);
and U9043 (N_9043,N_4640,N_4076);
nand U9044 (N_9044,N_3371,N_2820);
nor U9045 (N_9045,N_5026,N_2673);
nor U9046 (N_9046,N_3993,N_5335);
and U9047 (N_9047,N_3351,N_2999);
nor U9048 (N_9048,N_5193,N_4838);
nor U9049 (N_9049,N_381,N_2021);
or U9050 (N_9050,N_2103,N_1146);
and U9051 (N_9051,N_3448,N_6114);
nor U9052 (N_9052,N_4578,N_4610);
nand U9053 (N_9053,N_1773,N_3946);
nor U9054 (N_9054,N_3574,N_4872);
nand U9055 (N_9055,N_3907,N_3509);
nand U9056 (N_9056,N_2786,N_3135);
or U9057 (N_9057,N_2311,N_2690);
and U9058 (N_9058,N_889,N_5436);
nand U9059 (N_9059,N_5496,N_3234);
nand U9060 (N_9060,N_1970,N_854);
or U9061 (N_9061,N_5972,N_1369);
nand U9062 (N_9062,N_1391,N_3959);
or U9063 (N_9063,N_348,N_2568);
or U9064 (N_9064,N_4003,N_1551);
nand U9065 (N_9065,N_208,N_4148);
nand U9066 (N_9066,N_1057,N_3865);
nor U9067 (N_9067,N_5334,N_5204);
nor U9068 (N_9068,N_5590,N_6107);
or U9069 (N_9069,N_5437,N_604);
and U9070 (N_9070,N_1718,N_5246);
nor U9071 (N_9071,N_270,N_4843);
or U9072 (N_9072,N_4484,N_1643);
nand U9073 (N_9073,N_1105,N_2407);
and U9074 (N_9074,N_5924,N_3474);
nand U9075 (N_9075,N_880,N_5377);
or U9076 (N_9076,N_1361,N_4457);
and U9077 (N_9077,N_1697,N_5406);
nand U9078 (N_9078,N_2430,N_122);
nand U9079 (N_9079,N_860,N_1297);
nand U9080 (N_9080,N_1384,N_4765);
or U9081 (N_9081,N_4692,N_2166);
nand U9082 (N_9082,N_4084,N_293);
nand U9083 (N_9083,N_1760,N_1556);
nand U9084 (N_9084,N_2683,N_4985);
nand U9085 (N_9085,N_4202,N_2125);
nor U9086 (N_9086,N_2963,N_1941);
nand U9087 (N_9087,N_3675,N_4390);
nand U9088 (N_9088,N_552,N_1946);
and U9089 (N_9089,N_1755,N_590);
nor U9090 (N_9090,N_295,N_455);
nand U9091 (N_9091,N_119,N_684);
and U9092 (N_9092,N_2263,N_3304);
nor U9093 (N_9093,N_4293,N_1157);
nor U9094 (N_9094,N_1868,N_511);
nand U9095 (N_9095,N_6233,N_146);
or U9096 (N_9096,N_4070,N_1314);
nand U9097 (N_9097,N_2815,N_2830);
or U9098 (N_9098,N_4388,N_1966);
or U9099 (N_9099,N_4368,N_301);
nor U9100 (N_9100,N_2466,N_2105);
nand U9101 (N_9101,N_964,N_2507);
nor U9102 (N_9102,N_3828,N_2331);
nor U9103 (N_9103,N_1657,N_4918);
or U9104 (N_9104,N_3141,N_4396);
nand U9105 (N_9105,N_5138,N_821);
nor U9106 (N_9106,N_3733,N_5834);
nor U9107 (N_9107,N_4344,N_2889);
and U9108 (N_9108,N_5673,N_898);
or U9109 (N_9109,N_2850,N_3020);
nor U9110 (N_9110,N_129,N_2035);
nor U9111 (N_9111,N_60,N_5983);
nor U9112 (N_9112,N_5638,N_6065);
or U9113 (N_9113,N_4379,N_4595);
nand U9114 (N_9114,N_5145,N_2675);
or U9115 (N_9115,N_2616,N_4345);
nor U9116 (N_9116,N_1540,N_845);
nor U9117 (N_9117,N_5450,N_1954);
xor U9118 (N_9118,N_4005,N_3470);
nor U9119 (N_9119,N_1144,N_3432);
nor U9120 (N_9120,N_1613,N_4978);
or U9121 (N_9121,N_3791,N_467);
nand U9122 (N_9122,N_2476,N_2169);
or U9123 (N_9123,N_3476,N_2800);
nor U9124 (N_9124,N_6204,N_3067);
nand U9125 (N_9125,N_2741,N_925);
nor U9126 (N_9126,N_1616,N_2434);
or U9127 (N_9127,N_1816,N_5915);
xnor U9128 (N_9128,N_3047,N_3937);
and U9129 (N_9129,N_4458,N_2028);
and U9130 (N_9130,N_2160,N_3604);
nor U9131 (N_9131,N_5047,N_4405);
and U9132 (N_9132,N_3991,N_4928);
and U9133 (N_9133,N_5603,N_5870);
nor U9134 (N_9134,N_3325,N_4785);
or U9135 (N_9135,N_3627,N_3213);
nand U9136 (N_9136,N_2901,N_3721);
nor U9137 (N_9137,N_2475,N_1772);
and U9138 (N_9138,N_3689,N_2351);
xor U9139 (N_9139,N_4089,N_5113);
nor U9140 (N_9140,N_5117,N_1692);
nand U9141 (N_9141,N_2017,N_1434);
or U9142 (N_9142,N_363,N_1097);
nor U9143 (N_9143,N_4589,N_2628);
and U9144 (N_9144,N_286,N_3519);
and U9145 (N_9145,N_223,N_958);
nand U9146 (N_9146,N_2086,N_1650);
nand U9147 (N_9147,N_4839,N_2308);
nor U9148 (N_9148,N_2077,N_4674);
nand U9149 (N_9149,N_5052,N_5748);
and U9150 (N_9150,N_1275,N_453);
nand U9151 (N_9151,N_5568,N_3289);
and U9152 (N_9152,N_4023,N_4976);
or U9153 (N_9153,N_4448,N_1959);
nor U9154 (N_9154,N_600,N_5967);
or U9155 (N_9155,N_3942,N_3971);
nor U9156 (N_9156,N_820,N_3064);
nor U9157 (N_9157,N_4611,N_4952);
and U9158 (N_9158,N_6055,N_1151);
and U9159 (N_9159,N_761,N_1802);
and U9160 (N_9160,N_4761,N_48);
or U9161 (N_9161,N_3156,N_1953);
nand U9162 (N_9162,N_4426,N_1469);
nand U9163 (N_9163,N_3076,N_5269);
nor U9164 (N_9164,N_2750,N_4580);
or U9165 (N_9165,N_4818,N_482);
nand U9166 (N_9166,N_5527,N_5916);
nor U9167 (N_9167,N_5171,N_5911);
nand U9168 (N_9168,N_3764,N_5486);
nand U9169 (N_9169,N_5095,N_3774);
nand U9170 (N_9170,N_470,N_1408);
nor U9171 (N_9171,N_5158,N_1499);
nand U9172 (N_9172,N_2593,N_3426);
or U9173 (N_9173,N_2306,N_4298);
nor U9174 (N_9174,N_1849,N_2947);
xnor U9175 (N_9175,N_3941,N_5975);
nor U9176 (N_9176,N_4720,N_1705);
nand U9177 (N_9177,N_406,N_4336);
nand U9178 (N_9178,N_5300,N_2151);
nand U9179 (N_9179,N_3979,N_5063);
and U9180 (N_9180,N_985,N_990);
nand U9181 (N_9181,N_95,N_5471);
nand U9182 (N_9182,N_3114,N_5431);
and U9183 (N_9183,N_524,N_262);
and U9184 (N_9184,N_4968,N_1559);
nor U9185 (N_9185,N_6063,N_6212);
nand U9186 (N_9186,N_912,N_5676);
and U9187 (N_9187,N_4123,N_6192);
or U9188 (N_9188,N_1820,N_3823);
or U9189 (N_9189,N_6137,N_5093);
nand U9190 (N_9190,N_3162,N_2365);
nor U9191 (N_9191,N_478,N_4723);
or U9192 (N_9192,N_88,N_2056);
nand U9193 (N_9193,N_62,N_827);
and U9194 (N_9194,N_2266,N_3957);
and U9195 (N_9195,N_2147,N_1990);
nand U9196 (N_9196,N_4171,N_1584);
and U9197 (N_9197,N_3607,N_322);
and U9198 (N_9198,N_1409,N_3912);
nand U9199 (N_9199,N_2964,N_1310);
and U9200 (N_9200,N_70,N_2291);
nor U9201 (N_9201,N_5839,N_1597);
nand U9202 (N_9202,N_5512,N_680);
and U9203 (N_9203,N_4514,N_4915);
or U9204 (N_9204,N_3475,N_907);
or U9205 (N_9205,N_2462,N_75);
nor U9206 (N_9206,N_5862,N_4750);
nand U9207 (N_9207,N_2699,N_4424);
nor U9208 (N_9208,N_2938,N_564);
nand U9209 (N_9209,N_1632,N_1787);
and U9210 (N_9210,N_4518,N_2411);
and U9211 (N_9211,N_3861,N_5572);
nand U9212 (N_9212,N_2794,N_3767);
nor U9213 (N_9213,N_431,N_5429);
and U9214 (N_9214,N_1797,N_3954);
nor U9215 (N_9215,N_2074,N_4520);
nor U9216 (N_9216,N_2370,N_4192);
nor U9217 (N_9217,N_32,N_584);
nand U9218 (N_9218,N_1328,N_6215);
and U9219 (N_9219,N_5355,N_5606);
or U9220 (N_9220,N_1237,N_5885);
nor U9221 (N_9221,N_3985,N_2393);
nor U9222 (N_9222,N_10,N_5647);
or U9223 (N_9223,N_5984,N_5054);
nand U9224 (N_9224,N_3018,N_5801);
nand U9225 (N_9225,N_954,N_5461);
and U9226 (N_9226,N_7,N_5481);
nand U9227 (N_9227,N_6239,N_1112);
and U9228 (N_9228,N_3090,N_466);
nor U9229 (N_9229,N_3920,N_3239);
and U9230 (N_9230,N_1038,N_2363);
or U9231 (N_9231,N_1248,N_5430);
nand U9232 (N_9232,N_244,N_1763);
or U9233 (N_9233,N_1324,N_5709);
nor U9234 (N_9234,N_6232,N_3719);
nand U9235 (N_9235,N_1936,N_1428);
or U9236 (N_9236,N_2167,N_1837);
nor U9237 (N_9237,N_4311,N_1694);
nor U9238 (N_9238,N_4375,N_2190);
nor U9239 (N_9239,N_653,N_1508);
nor U9240 (N_9240,N_6138,N_4999);
and U9241 (N_9241,N_2269,N_3471);
or U9242 (N_9242,N_1298,N_3177);
and U9243 (N_9243,N_387,N_1420);
nand U9244 (N_9244,N_2822,N_2338);
nor U9245 (N_9245,N_1505,N_669);
and U9246 (N_9246,N_5129,N_2753);
and U9247 (N_9247,N_2625,N_613);
nor U9248 (N_9248,N_1400,N_248);
and U9249 (N_9249,N_4019,N_2663);
or U9250 (N_9250,N_3290,N_6058);
and U9251 (N_9251,N_1312,N_3273);
and U9252 (N_9252,N_4151,N_4327);
nor U9253 (N_9253,N_735,N_4954);
nand U9254 (N_9254,N_1231,N_250);
nor U9255 (N_9255,N_2923,N_1212);
or U9256 (N_9256,N_1009,N_4888);
nor U9257 (N_9257,N_6214,N_787);
xnor U9258 (N_9258,N_651,N_309);
nor U9259 (N_9259,N_3910,N_595);
nand U9260 (N_9260,N_1683,N_844);
and U9261 (N_9261,N_494,N_3799);
and U9262 (N_9262,N_3598,N_5841);
nor U9263 (N_9263,N_1423,N_5923);
or U9264 (N_9264,N_3019,N_4665);
nand U9265 (N_9265,N_5665,N_2257);
and U9266 (N_9266,N_2689,N_4565);
nor U9267 (N_9267,N_2595,N_5265);
nand U9268 (N_9268,N_5710,N_2679);
nor U9269 (N_9269,N_2665,N_2948);
nor U9270 (N_9270,N_4024,N_411);
nor U9271 (N_9271,N_6,N_6068);
and U9272 (N_9272,N_4687,N_3271);
and U9273 (N_9273,N_784,N_1265);
or U9274 (N_9274,N_1139,N_679);
nor U9275 (N_9275,N_2531,N_2281);
and U9276 (N_9276,N_3409,N_1091);
and U9277 (N_9277,N_4333,N_2394);
nor U9278 (N_9278,N_3185,N_2621);
nor U9279 (N_9279,N_3227,N_3333);
xnor U9280 (N_9280,N_2142,N_4634);
nor U9281 (N_9281,N_2143,N_3900);
and U9282 (N_9282,N_2491,N_1341);
or U9283 (N_9283,N_2731,N_3269);
and U9284 (N_9284,N_4668,N_1141);
nand U9285 (N_9285,N_2564,N_291);
nand U9286 (N_9286,N_1963,N_1927);
or U9287 (N_9287,N_4177,N_3103);
nor U9288 (N_9288,N_851,N_5694);
and U9289 (N_9289,N_4252,N_966);
or U9290 (N_9290,N_4463,N_1082);
nor U9291 (N_9291,N_80,N_5892);
nor U9292 (N_9292,N_3313,N_3250);
or U9293 (N_9293,N_5678,N_2852);
nor U9294 (N_9294,N_101,N_3918);
nor U9295 (N_9295,N_2908,N_5944);
nor U9296 (N_9296,N_4155,N_989);
or U9297 (N_9297,N_3390,N_4154);
or U9298 (N_9298,N_4443,N_4259);
and U9299 (N_9299,N_1940,N_1292);
nor U9300 (N_9300,N_1751,N_5860);
nand U9301 (N_9301,N_1473,N_4012);
and U9302 (N_9302,N_3864,N_2579);
nor U9303 (N_9303,N_1334,N_6128);
xor U9304 (N_9304,N_3465,N_370);
nor U9305 (N_9305,N_610,N_2523);
nand U9306 (N_9306,N_3913,N_3091);
nand U9307 (N_9307,N_5796,N_45);
or U9308 (N_9308,N_503,N_602);
nand U9309 (N_9309,N_5912,N_5726);
or U9310 (N_9310,N_1562,N_3863);
nor U9311 (N_9311,N_165,N_6142);
nor U9312 (N_9312,N_436,N_806);
and U9313 (N_9313,N_5262,N_705);
nor U9314 (N_9314,N_4142,N_4657);
or U9315 (N_9315,N_2239,N_6028);
nand U9316 (N_9316,N_6093,N_5493);
nor U9317 (N_9317,N_5613,N_6181);
nor U9318 (N_9318,N_818,N_4383);
nor U9319 (N_9319,N_3737,N_2828);
nand U9320 (N_9320,N_6087,N_4647);
or U9321 (N_9321,N_1710,N_464);
or U9322 (N_9322,N_3299,N_5050);
nor U9323 (N_9323,N_13,N_82);
or U9324 (N_9324,N_1337,N_6234);
or U9325 (N_9325,N_4608,N_2413);
and U9326 (N_9326,N_2,N_5494);
or U9327 (N_9327,N_956,N_570);
nand U9328 (N_9328,N_640,N_712);
nand U9329 (N_9329,N_359,N_3248);
or U9330 (N_9330,N_2787,N_530);
nand U9331 (N_9331,N_2063,N_5503);
or U9332 (N_9332,N_1440,N_5708);
and U9333 (N_9333,N_1519,N_3879);
nor U9334 (N_9334,N_246,N_5386);
nand U9335 (N_9335,N_4182,N_1877);
or U9336 (N_9336,N_5645,N_2757);
or U9337 (N_9337,N_5076,N_1577);
and U9338 (N_9338,N_4212,N_2362);
or U9339 (N_9339,N_4471,N_2845);
or U9340 (N_9340,N_3958,N_4477);
or U9341 (N_9341,N_4079,N_2010);
nand U9342 (N_9342,N_2477,N_2437);
and U9343 (N_9343,N_3479,N_3829);
nor U9344 (N_9344,N_4035,N_1722);
nor U9345 (N_9345,N_1604,N_4000);
nor U9346 (N_9346,N_794,N_1972);
nor U9347 (N_9347,N_6154,N_3818);
and U9348 (N_9348,N_1398,N_1598);
nor U9349 (N_9349,N_3553,N_3033);
and U9350 (N_9350,N_3820,N_5506);
and U9351 (N_9351,N_6209,N_2740);
nand U9352 (N_9352,N_4747,N_5465);
or U9353 (N_9353,N_4174,N_529);
and U9354 (N_9354,N_314,N_3214);
xnor U9355 (N_9355,N_4644,N_415);
xnor U9356 (N_9356,N_4386,N_4593);
nor U9357 (N_9357,N_195,N_2893);
and U9358 (N_9358,N_1574,N_2244);
nor U9359 (N_9359,N_1054,N_1087);
and U9360 (N_9360,N_3428,N_3591);
nand U9361 (N_9361,N_2720,N_567);
nor U9362 (N_9362,N_4224,N_5102);
nor U9363 (N_9363,N_2493,N_681);
and U9364 (N_9364,N_1228,N_5329);
xnor U9365 (N_9365,N_5201,N_5756);
nand U9366 (N_9366,N_3529,N_1611);
and U9367 (N_9367,N_5614,N_445);
nand U9368 (N_9368,N_4632,N_4493);
nand U9369 (N_9369,N_2419,N_1818);
or U9370 (N_9370,N_1684,N_689);
nor U9371 (N_9371,N_1674,N_2136);
nor U9372 (N_9372,N_5835,N_4847);
nor U9373 (N_9373,N_6189,N_3026);
nand U9374 (N_9374,N_4556,N_4043);
nand U9375 (N_9375,N_1543,N_2749);
nor U9376 (N_9376,N_4920,N_5754);
or U9377 (N_9377,N_336,N_2745);
and U9378 (N_9378,N_3583,N_182);
nor U9379 (N_9379,N_5005,N_4683);
or U9380 (N_9380,N_253,N_2742);
and U9381 (N_9381,N_3321,N_4516);
nor U9382 (N_9382,N_465,N_683);
or U9383 (N_9383,N_2321,N_1527);
and U9384 (N_9384,N_4198,N_4861);
and U9385 (N_9385,N_740,N_6142);
nand U9386 (N_9386,N_361,N_492);
nor U9387 (N_9387,N_6152,N_4404);
nor U9388 (N_9388,N_5877,N_4527);
or U9389 (N_9389,N_2724,N_587);
and U9390 (N_9390,N_4921,N_1401);
nand U9391 (N_9391,N_5691,N_4995);
nor U9392 (N_9392,N_5773,N_1373);
nand U9393 (N_9393,N_4078,N_1595);
nor U9394 (N_9394,N_946,N_3454);
nand U9395 (N_9395,N_1301,N_1223);
or U9396 (N_9396,N_5365,N_2660);
nand U9397 (N_9397,N_4212,N_2029);
nor U9398 (N_9398,N_2859,N_692);
or U9399 (N_9399,N_1888,N_3129);
nand U9400 (N_9400,N_3333,N_4603);
xnor U9401 (N_9401,N_1871,N_3877);
nor U9402 (N_9402,N_843,N_4775);
xnor U9403 (N_9403,N_4408,N_1491);
nor U9404 (N_9404,N_476,N_969);
nand U9405 (N_9405,N_6216,N_5486);
nor U9406 (N_9406,N_6215,N_2277);
nor U9407 (N_9407,N_2220,N_3157);
or U9408 (N_9408,N_5934,N_5657);
and U9409 (N_9409,N_2471,N_4856);
and U9410 (N_9410,N_3167,N_4201);
nand U9411 (N_9411,N_61,N_1503);
nand U9412 (N_9412,N_2570,N_3630);
nand U9413 (N_9413,N_39,N_4095);
and U9414 (N_9414,N_4188,N_3352);
or U9415 (N_9415,N_5073,N_560);
or U9416 (N_9416,N_5438,N_5780);
nor U9417 (N_9417,N_2717,N_5431);
nor U9418 (N_9418,N_4378,N_4275);
nor U9419 (N_9419,N_1514,N_76);
and U9420 (N_9420,N_5038,N_3239);
and U9421 (N_9421,N_1447,N_4080);
or U9422 (N_9422,N_4565,N_5280);
nand U9423 (N_9423,N_5687,N_6120);
nand U9424 (N_9424,N_4335,N_3442);
or U9425 (N_9425,N_4694,N_5345);
and U9426 (N_9426,N_2524,N_2151);
and U9427 (N_9427,N_5110,N_2199);
nand U9428 (N_9428,N_4709,N_3016);
and U9429 (N_9429,N_3713,N_4696);
nand U9430 (N_9430,N_2502,N_4737);
nand U9431 (N_9431,N_4006,N_6091);
and U9432 (N_9432,N_1148,N_4525);
and U9433 (N_9433,N_2610,N_5866);
or U9434 (N_9434,N_5454,N_5299);
nor U9435 (N_9435,N_2103,N_77);
and U9436 (N_9436,N_3213,N_3290);
and U9437 (N_9437,N_5936,N_117);
or U9438 (N_9438,N_1779,N_1168);
nand U9439 (N_9439,N_1776,N_93);
nor U9440 (N_9440,N_5509,N_2101);
and U9441 (N_9441,N_769,N_4122);
and U9442 (N_9442,N_1237,N_3631);
nand U9443 (N_9443,N_465,N_1143);
or U9444 (N_9444,N_1058,N_3326);
or U9445 (N_9445,N_5422,N_62);
nand U9446 (N_9446,N_4533,N_1883);
or U9447 (N_9447,N_1020,N_184);
or U9448 (N_9448,N_1610,N_3358);
xor U9449 (N_9449,N_1765,N_3865);
nand U9450 (N_9450,N_5998,N_357);
nand U9451 (N_9451,N_4877,N_5465);
nand U9452 (N_9452,N_2162,N_4063);
nor U9453 (N_9453,N_4920,N_6084);
or U9454 (N_9454,N_1590,N_308);
or U9455 (N_9455,N_5388,N_3116);
or U9456 (N_9456,N_4346,N_1113);
nand U9457 (N_9457,N_4710,N_4728);
nand U9458 (N_9458,N_2812,N_4904);
nand U9459 (N_9459,N_2331,N_4323);
nand U9460 (N_9460,N_814,N_175);
or U9461 (N_9461,N_6104,N_3798);
or U9462 (N_9462,N_3062,N_5006);
nand U9463 (N_9463,N_732,N_3381);
and U9464 (N_9464,N_4855,N_5245);
and U9465 (N_9465,N_4619,N_5376);
or U9466 (N_9466,N_5322,N_3982);
nand U9467 (N_9467,N_1363,N_6245);
and U9468 (N_9468,N_5918,N_2985);
or U9469 (N_9469,N_5702,N_3930);
and U9470 (N_9470,N_974,N_4677);
nand U9471 (N_9471,N_665,N_2476);
nand U9472 (N_9472,N_1454,N_3849);
and U9473 (N_9473,N_1847,N_5479);
nor U9474 (N_9474,N_5493,N_3276);
or U9475 (N_9475,N_3877,N_5924);
nand U9476 (N_9476,N_3944,N_3327);
nor U9477 (N_9477,N_4998,N_4525);
and U9478 (N_9478,N_2412,N_5474);
nor U9479 (N_9479,N_2045,N_2184);
nor U9480 (N_9480,N_3875,N_4367);
nor U9481 (N_9481,N_62,N_5170);
and U9482 (N_9482,N_3415,N_2630);
nand U9483 (N_9483,N_1487,N_26);
nand U9484 (N_9484,N_5639,N_1784);
or U9485 (N_9485,N_3077,N_4080);
nand U9486 (N_9486,N_856,N_4922);
or U9487 (N_9487,N_2676,N_749);
or U9488 (N_9488,N_3934,N_1728);
nor U9489 (N_9489,N_4239,N_3506);
nor U9490 (N_9490,N_6102,N_630);
and U9491 (N_9491,N_713,N_4612);
nand U9492 (N_9492,N_4923,N_1129);
nand U9493 (N_9493,N_270,N_724);
and U9494 (N_9494,N_3466,N_112);
nor U9495 (N_9495,N_121,N_1288);
nand U9496 (N_9496,N_1500,N_794);
nor U9497 (N_9497,N_589,N_2976);
nand U9498 (N_9498,N_2746,N_5833);
or U9499 (N_9499,N_1858,N_5204);
nor U9500 (N_9500,N_1977,N_2036);
nand U9501 (N_9501,N_4550,N_3338);
and U9502 (N_9502,N_2113,N_3224);
nor U9503 (N_9503,N_4291,N_59);
nand U9504 (N_9504,N_821,N_5495);
nor U9505 (N_9505,N_750,N_4296);
nor U9506 (N_9506,N_5239,N_4164);
and U9507 (N_9507,N_2273,N_1860);
nor U9508 (N_9508,N_4369,N_1611);
and U9509 (N_9509,N_2722,N_3420);
or U9510 (N_9510,N_2147,N_73);
nor U9511 (N_9511,N_1131,N_5447);
nor U9512 (N_9512,N_297,N_4252);
nor U9513 (N_9513,N_4233,N_1600);
nor U9514 (N_9514,N_2062,N_5027);
or U9515 (N_9515,N_4783,N_4886);
and U9516 (N_9516,N_5471,N_3908);
nand U9517 (N_9517,N_5444,N_6136);
nor U9518 (N_9518,N_3392,N_6118);
or U9519 (N_9519,N_2796,N_1933);
and U9520 (N_9520,N_3774,N_82);
and U9521 (N_9521,N_712,N_177);
or U9522 (N_9522,N_3583,N_4000);
nor U9523 (N_9523,N_5177,N_5786);
or U9524 (N_9524,N_3441,N_6015);
nor U9525 (N_9525,N_1853,N_163);
nor U9526 (N_9526,N_5722,N_462);
or U9527 (N_9527,N_999,N_1097);
or U9528 (N_9528,N_4305,N_1319);
or U9529 (N_9529,N_5164,N_1143);
nand U9530 (N_9530,N_5504,N_235);
nor U9531 (N_9531,N_2762,N_4096);
and U9532 (N_9532,N_4465,N_74);
or U9533 (N_9533,N_482,N_1394);
nor U9534 (N_9534,N_3723,N_964);
or U9535 (N_9535,N_101,N_3453);
and U9536 (N_9536,N_4865,N_5369);
and U9537 (N_9537,N_339,N_1976);
nand U9538 (N_9538,N_3972,N_6134);
nor U9539 (N_9539,N_44,N_1410);
nand U9540 (N_9540,N_647,N_2345);
xnor U9541 (N_9541,N_1149,N_68);
or U9542 (N_9542,N_5481,N_5777);
or U9543 (N_9543,N_4065,N_6034);
nor U9544 (N_9544,N_2847,N_1624);
or U9545 (N_9545,N_5290,N_5210);
and U9546 (N_9546,N_1798,N_2481);
or U9547 (N_9547,N_4237,N_1979);
or U9548 (N_9548,N_3363,N_3789);
nor U9549 (N_9549,N_3209,N_1973);
nand U9550 (N_9550,N_3568,N_1672);
nor U9551 (N_9551,N_5652,N_444);
and U9552 (N_9552,N_615,N_2831);
and U9553 (N_9553,N_3986,N_4853);
nor U9554 (N_9554,N_5156,N_3532);
nor U9555 (N_9555,N_408,N_5193);
and U9556 (N_9556,N_2786,N_4290);
or U9557 (N_9557,N_2164,N_3917);
nand U9558 (N_9558,N_3947,N_1992);
xnor U9559 (N_9559,N_653,N_3586);
and U9560 (N_9560,N_3302,N_190);
or U9561 (N_9561,N_3042,N_3440);
or U9562 (N_9562,N_5876,N_3279);
nor U9563 (N_9563,N_5517,N_115);
nand U9564 (N_9564,N_6193,N_4262);
nor U9565 (N_9565,N_1522,N_4368);
or U9566 (N_9566,N_694,N_4106);
nor U9567 (N_9567,N_3427,N_1914);
xor U9568 (N_9568,N_2925,N_5145);
or U9569 (N_9569,N_4714,N_3448);
or U9570 (N_9570,N_3611,N_4351);
nor U9571 (N_9571,N_3649,N_3659);
or U9572 (N_9572,N_2220,N_4729);
nand U9573 (N_9573,N_3613,N_5091);
nand U9574 (N_9574,N_1170,N_4601);
nand U9575 (N_9575,N_4815,N_2002);
or U9576 (N_9576,N_4169,N_3953);
and U9577 (N_9577,N_5908,N_1054);
or U9578 (N_9578,N_2445,N_3175);
or U9579 (N_9579,N_1541,N_2286);
nor U9580 (N_9580,N_5931,N_4344);
nor U9581 (N_9581,N_1015,N_3814);
nand U9582 (N_9582,N_559,N_3184);
nand U9583 (N_9583,N_5239,N_3625);
or U9584 (N_9584,N_2247,N_2181);
and U9585 (N_9585,N_649,N_2598);
nand U9586 (N_9586,N_3601,N_5045);
nor U9587 (N_9587,N_4639,N_2858);
nand U9588 (N_9588,N_1644,N_3397);
nand U9589 (N_9589,N_4967,N_5253);
nand U9590 (N_9590,N_5255,N_847);
nor U9591 (N_9591,N_5406,N_348);
and U9592 (N_9592,N_5526,N_6129);
nor U9593 (N_9593,N_1958,N_1926);
and U9594 (N_9594,N_572,N_3617);
nand U9595 (N_9595,N_1032,N_4471);
nand U9596 (N_9596,N_4512,N_3706);
nor U9597 (N_9597,N_5730,N_1686);
or U9598 (N_9598,N_4558,N_3004);
nor U9599 (N_9599,N_4562,N_693);
nor U9600 (N_9600,N_2970,N_245);
and U9601 (N_9601,N_2972,N_4816);
nand U9602 (N_9602,N_3592,N_5466);
and U9603 (N_9603,N_4800,N_4044);
and U9604 (N_9604,N_597,N_5456);
and U9605 (N_9605,N_1891,N_373);
nand U9606 (N_9606,N_1721,N_5707);
nand U9607 (N_9607,N_91,N_1552);
and U9608 (N_9608,N_5645,N_1015);
nor U9609 (N_9609,N_1090,N_729);
nand U9610 (N_9610,N_3798,N_357);
and U9611 (N_9611,N_1850,N_88);
and U9612 (N_9612,N_5407,N_1823);
and U9613 (N_9613,N_1142,N_3872);
nor U9614 (N_9614,N_5785,N_5425);
nor U9615 (N_9615,N_3798,N_3289);
nor U9616 (N_9616,N_5368,N_2758);
and U9617 (N_9617,N_2225,N_73);
and U9618 (N_9618,N_1798,N_2289);
or U9619 (N_9619,N_3403,N_629);
nor U9620 (N_9620,N_2411,N_5596);
nand U9621 (N_9621,N_5084,N_5163);
nand U9622 (N_9622,N_367,N_3643);
and U9623 (N_9623,N_4951,N_910);
or U9624 (N_9624,N_4000,N_300);
nand U9625 (N_9625,N_1460,N_5062);
nor U9626 (N_9626,N_4915,N_5521);
and U9627 (N_9627,N_3911,N_4324);
or U9628 (N_9628,N_3639,N_27);
or U9629 (N_9629,N_6160,N_2901);
nor U9630 (N_9630,N_2056,N_4465);
nor U9631 (N_9631,N_676,N_3644);
nand U9632 (N_9632,N_1178,N_3098);
nor U9633 (N_9633,N_2627,N_4160);
or U9634 (N_9634,N_2024,N_1472);
nand U9635 (N_9635,N_834,N_5096);
nor U9636 (N_9636,N_4066,N_3515);
or U9637 (N_9637,N_4432,N_4948);
nor U9638 (N_9638,N_725,N_3989);
and U9639 (N_9639,N_4442,N_4708);
nor U9640 (N_9640,N_3648,N_3056);
or U9641 (N_9641,N_310,N_4228);
nor U9642 (N_9642,N_1133,N_4263);
nor U9643 (N_9643,N_5024,N_3934);
nor U9644 (N_9644,N_1667,N_3277);
nand U9645 (N_9645,N_3645,N_4939);
and U9646 (N_9646,N_2136,N_4685);
xnor U9647 (N_9647,N_3848,N_359);
or U9648 (N_9648,N_6187,N_4843);
nor U9649 (N_9649,N_5817,N_5680);
nor U9650 (N_9650,N_3119,N_2452);
and U9651 (N_9651,N_5902,N_5617);
or U9652 (N_9652,N_2476,N_2964);
nand U9653 (N_9653,N_5387,N_1990);
or U9654 (N_9654,N_5026,N_5574);
nor U9655 (N_9655,N_302,N_938);
nor U9656 (N_9656,N_4865,N_2266);
nand U9657 (N_9657,N_2971,N_5693);
nand U9658 (N_9658,N_1216,N_2849);
nor U9659 (N_9659,N_895,N_2814);
xor U9660 (N_9660,N_692,N_3222);
nand U9661 (N_9661,N_3051,N_3085);
or U9662 (N_9662,N_4928,N_3074);
nor U9663 (N_9663,N_4878,N_6135);
nor U9664 (N_9664,N_5981,N_2039);
and U9665 (N_9665,N_2129,N_5318);
and U9666 (N_9666,N_1960,N_171);
nand U9667 (N_9667,N_162,N_1302);
nor U9668 (N_9668,N_3238,N_1748);
nor U9669 (N_9669,N_3259,N_1684);
nand U9670 (N_9670,N_830,N_1144);
and U9671 (N_9671,N_2227,N_4512);
nand U9672 (N_9672,N_2281,N_5237);
or U9673 (N_9673,N_198,N_3636);
nand U9674 (N_9674,N_3066,N_118);
or U9675 (N_9675,N_1433,N_528);
nand U9676 (N_9676,N_5960,N_2048);
and U9677 (N_9677,N_3559,N_3796);
and U9678 (N_9678,N_2519,N_3391);
nand U9679 (N_9679,N_4570,N_111);
or U9680 (N_9680,N_5789,N_2765);
nor U9681 (N_9681,N_120,N_4596);
nor U9682 (N_9682,N_2456,N_1165);
and U9683 (N_9683,N_4355,N_2578);
and U9684 (N_9684,N_5959,N_4601);
and U9685 (N_9685,N_2241,N_1995);
or U9686 (N_9686,N_1610,N_4883);
and U9687 (N_9687,N_376,N_2194);
and U9688 (N_9688,N_5744,N_2822);
or U9689 (N_9689,N_1134,N_3740);
and U9690 (N_9690,N_5090,N_6040);
or U9691 (N_9691,N_6207,N_3146);
and U9692 (N_9692,N_5769,N_1929);
and U9693 (N_9693,N_3586,N_3413);
and U9694 (N_9694,N_1138,N_5639);
nor U9695 (N_9695,N_4734,N_5855);
and U9696 (N_9696,N_2029,N_122);
or U9697 (N_9697,N_2687,N_1035);
nand U9698 (N_9698,N_8,N_3330);
nand U9699 (N_9699,N_4589,N_5757);
and U9700 (N_9700,N_4174,N_3679);
nor U9701 (N_9701,N_1488,N_1547);
or U9702 (N_9702,N_1527,N_3470);
nor U9703 (N_9703,N_5592,N_5184);
and U9704 (N_9704,N_2680,N_5674);
and U9705 (N_9705,N_5323,N_4518);
or U9706 (N_9706,N_1181,N_1008);
or U9707 (N_9707,N_3633,N_1510);
nor U9708 (N_9708,N_2676,N_1714);
or U9709 (N_9709,N_4415,N_1590);
nor U9710 (N_9710,N_1261,N_1615);
nand U9711 (N_9711,N_639,N_5623);
and U9712 (N_9712,N_4288,N_1588);
nor U9713 (N_9713,N_3753,N_4622);
and U9714 (N_9714,N_1786,N_3921);
nand U9715 (N_9715,N_5259,N_2429);
nor U9716 (N_9716,N_3891,N_4657);
nor U9717 (N_9717,N_566,N_2764);
nor U9718 (N_9718,N_1107,N_563);
or U9719 (N_9719,N_1792,N_2826);
nor U9720 (N_9720,N_891,N_1529);
nor U9721 (N_9721,N_423,N_563);
nor U9722 (N_9722,N_2096,N_1287);
and U9723 (N_9723,N_4842,N_2707);
nand U9724 (N_9724,N_1459,N_1905);
or U9725 (N_9725,N_4999,N_5816);
nand U9726 (N_9726,N_5418,N_4546);
nor U9727 (N_9727,N_1860,N_2023);
nand U9728 (N_9728,N_1147,N_927);
or U9729 (N_9729,N_2225,N_3589);
nand U9730 (N_9730,N_824,N_5677);
nand U9731 (N_9731,N_1588,N_3578);
or U9732 (N_9732,N_3413,N_3151);
nor U9733 (N_9733,N_405,N_3501);
nor U9734 (N_9734,N_383,N_3308);
nor U9735 (N_9735,N_6106,N_6029);
nand U9736 (N_9736,N_752,N_920);
nor U9737 (N_9737,N_665,N_3224);
and U9738 (N_9738,N_1327,N_5068);
nor U9739 (N_9739,N_2360,N_4475);
or U9740 (N_9740,N_3500,N_3396);
and U9741 (N_9741,N_5038,N_4288);
or U9742 (N_9742,N_3907,N_4010);
or U9743 (N_9743,N_50,N_3567);
nor U9744 (N_9744,N_2726,N_2393);
nor U9745 (N_9745,N_4926,N_3830);
nor U9746 (N_9746,N_3507,N_4036);
nand U9747 (N_9747,N_1250,N_351);
or U9748 (N_9748,N_2926,N_4359);
nand U9749 (N_9749,N_2879,N_2404);
or U9750 (N_9750,N_2465,N_29);
nor U9751 (N_9751,N_51,N_2960);
or U9752 (N_9752,N_6177,N_5996);
nor U9753 (N_9753,N_2194,N_4805);
nor U9754 (N_9754,N_3406,N_2144);
nor U9755 (N_9755,N_1409,N_3242);
nor U9756 (N_9756,N_120,N_2337);
nor U9757 (N_9757,N_5502,N_1043);
or U9758 (N_9758,N_568,N_5818);
xor U9759 (N_9759,N_6188,N_5149);
and U9760 (N_9760,N_2895,N_4370);
or U9761 (N_9761,N_134,N_424);
or U9762 (N_9762,N_2150,N_3045);
or U9763 (N_9763,N_5225,N_290);
nand U9764 (N_9764,N_2912,N_465);
nor U9765 (N_9765,N_5415,N_2520);
nor U9766 (N_9766,N_5499,N_750);
nand U9767 (N_9767,N_5486,N_5944);
nand U9768 (N_9768,N_5238,N_543);
and U9769 (N_9769,N_360,N_1584);
nor U9770 (N_9770,N_1843,N_3221);
and U9771 (N_9771,N_3441,N_1033);
and U9772 (N_9772,N_5805,N_1971);
and U9773 (N_9773,N_2836,N_5064);
nor U9774 (N_9774,N_5766,N_781);
nand U9775 (N_9775,N_1884,N_5952);
nor U9776 (N_9776,N_3191,N_3981);
nand U9777 (N_9777,N_2884,N_5280);
nand U9778 (N_9778,N_1401,N_6100);
nand U9779 (N_9779,N_4482,N_2757);
nor U9780 (N_9780,N_2554,N_5560);
or U9781 (N_9781,N_2069,N_3795);
and U9782 (N_9782,N_1472,N_2538);
and U9783 (N_9783,N_1505,N_3038);
and U9784 (N_9784,N_4407,N_4755);
nor U9785 (N_9785,N_1743,N_4272);
nor U9786 (N_9786,N_5038,N_5569);
and U9787 (N_9787,N_2113,N_3989);
nand U9788 (N_9788,N_4500,N_4999);
and U9789 (N_9789,N_3088,N_1648);
or U9790 (N_9790,N_2145,N_6211);
and U9791 (N_9791,N_274,N_2818);
nand U9792 (N_9792,N_5426,N_5836);
or U9793 (N_9793,N_4960,N_4169);
and U9794 (N_9794,N_158,N_2352);
and U9795 (N_9795,N_5850,N_6078);
and U9796 (N_9796,N_4282,N_4901);
and U9797 (N_9797,N_3893,N_143);
or U9798 (N_9798,N_1378,N_4201);
and U9799 (N_9799,N_2667,N_2921);
nand U9800 (N_9800,N_3790,N_5566);
nor U9801 (N_9801,N_445,N_1817);
and U9802 (N_9802,N_1672,N_2636);
nand U9803 (N_9803,N_2105,N_2965);
and U9804 (N_9804,N_5364,N_1777);
nand U9805 (N_9805,N_3338,N_520);
nor U9806 (N_9806,N_710,N_5784);
nand U9807 (N_9807,N_1047,N_3100);
or U9808 (N_9808,N_93,N_697);
nor U9809 (N_9809,N_5929,N_4299);
or U9810 (N_9810,N_2481,N_3343);
or U9811 (N_9811,N_2763,N_1018);
nand U9812 (N_9812,N_2831,N_4152);
and U9813 (N_9813,N_3953,N_5661);
and U9814 (N_9814,N_4732,N_2286);
nor U9815 (N_9815,N_6042,N_1060);
nand U9816 (N_9816,N_1578,N_273);
nand U9817 (N_9817,N_1946,N_4291);
nand U9818 (N_9818,N_4345,N_2214);
nor U9819 (N_9819,N_4201,N_5814);
nor U9820 (N_9820,N_2092,N_2216);
and U9821 (N_9821,N_3204,N_4338);
nor U9822 (N_9822,N_4427,N_3227);
and U9823 (N_9823,N_4533,N_2029);
nor U9824 (N_9824,N_1003,N_5407);
nand U9825 (N_9825,N_2594,N_6055);
nor U9826 (N_9826,N_5935,N_596);
nand U9827 (N_9827,N_2083,N_5003);
nor U9828 (N_9828,N_5769,N_4428);
or U9829 (N_9829,N_5442,N_932);
or U9830 (N_9830,N_3676,N_1111);
and U9831 (N_9831,N_1324,N_5942);
nand U9832 (N_9832,N_2846,N_5458);
nor U9833 (N_9833,N_1019,N_3519);
nor U9834 (N_9834,N_3128,N_72);
or U9835 (N_9835,N_1128,N_2104);
or U9836 (N_9836,N_1970,N_5074);
or U9837 (N_9837,N_4485,N_2438);
nor U9838 (N_9838,N_6202,N_571);
or U9839 (N_9839,N_5591,N_3143);
nor U9840 (N_9840,N_5313,N_1);
nand U9841 (N_9841,N_4747,N_506);
nand U9842 (N_9842,N_4338,N_4256);
nor U9843 (N_9843,N_4153,N_713);
or U9844 (N_9844,N_3977,N_78);
nand U9845 (N_9845,N_4472,N_4096);
or U9846 (N_9846,N_3803,N_5550);
nor U9847 (N_9847,N_251,N_4435);
nand U9848 (N_9848,N_1215,N_1863);
or U9849 (N_9849,N_988,N_4810);
or U9850 (N_9850,N_2589,N_2304);
and U9851 (N_9851,N_972,N_5166);
or U9852 (N_9852,N_1854,N_4934);
or U9853 (N_9853,N_5432,N_532);
nor U9854 (N_9854,N_1004,N_1430);
or U9855 (N_9855,N_4920,N_4798);
or U9856 (N_9856,N_2121,N_166);
and U9857 (N_9857,N_3844,N_1972);
and U9858 (N_9858,N_5785,N_5009);
and U9859 (N_9859,N_6053,N_5432);
nor U9860 (N_9860,N_3342,N_3448);
nand U9861 (N_9861,N_4281,N_1798);
or U9862 (N_9862,N_975,N_4993);
nand U9863 (N_9863,N_5713,N_2747);
and U9864 (N_9864,N_1092,N_2953);
and U9865 (N_9865,N_5877,N_1523);
and U9866 (N_9866,N_1434,N_5186);
or U9867 (N_9867,N_2006,N_3301);
or U9868 (N_9868,N_2270,N_82);
or U9869 (N_9869,N_4639,N_4058);
nand U9870 (N_9870,N_1103,N_5439);
and U9871 (N_9871,N_5803,N_1995);
nand U9872 (N_9872,N_461,N_262);
nor U9873 (N_9873,N_76,N_319);
nor U9874 (N_9874,N_4916,N_3538);
or U9875 (N_9875,N_6086,N_4729);
and U9876 (N_9876,N_485,N_4416);
xnor U9877 (N_9877,N_4312,N_3905);
nor U9878 (N_9878,N_1246,N_4475);
or U9879 (N_9879,N_3175,N_3926);
or U9880 (N_9880,N_422,N_5196);
nand U9881 (N_9881,N_1954,N_2964);
and U9882 (N_9882,N_4007,N_3585);
nor U9883 (N_9883,N_4144,N_2058);
and U9884 (N_9884,N_2277,N_1835);
nand U9885 (N_9885,N_274,N_3895);
nand U9886 (N_9886,N_6060,N_1102);
and U9887 (N_9887,N_1970,N_958);
or U9888 (N_9888,N_1360,N_4669);
nand U9889 (N_9889,N_953,N_4946);
or U9890 (N_9890,N_333,N_5401);
nor U9891 (N_9891,N_3382,N_4958);
or U9892 (N_9892,N_4240,N_5283);
and U9893 (N_9893,N_299,N_1788);
and U9894 (N_9894,N_3307,N_5114);
and U9895 (N_9895,N_5287,N_1288);
nand U9896 (N_9896,N_4500,N_1607);
nand U9897 (N_9897,N_4116,N_3494);
nor U9898 (N_9898,N_1004,N_5227);
nor U9899 (N_9899,N_5119,N_2609);
nor U9900 (N_9900,N_6151,N_5544);
or U9901 (N_9901,N_4122,N_2811);
and U9902 (N_9902,N_3691,N_3036);
or U9903 (N_9903,N_1944,N_346);
and U9904 (N_9904,N_2909,N_4868);
nand U9905 (N_9905,N_1972,N_425);
nand U9906 (N_9906,N_4120,N_763);
xnor U9907 (N_9907,N_3169,N_4168);
and U9908 (N_9908,N_2170,N_4997);
or U9909 (N_9909,N_481,N_5121);
nor U9910 (N_9910,N_5910,N_3951);
or U9911 (N_9911,N_4629,N_4642);
nand U9912 (N_9912,N_1960,N_5879);
or U9913 (N_9913,N_4838,N_3978);
or U9914 (N_9914,N_2304,N_5977);
nand U9915 (N_9915,N_78,N_5019);
nand U9916 (N_9916,N_5203,N_3265);
nand U9917 (N_9917,N_6216,N_2175);
and U9918 (N_9918,N_5163,N_1206);
nor U9919 (N_9919,N_5686,N_2564);
and U9920 (N_9920,N_1253,N_2984);
nand U9921 (N_9921,N_3102,N_3608);
or U9922 (N_9922,N_2424,N_5135);
nor U9923 (N_9923,N_4530,N_1109);
nand U9924 (N_9924,N_2097,N_4429);
nand U9925 (N_9925,N_2396,N_299);
nand U9926 (N_9926,N_1331,N_4894);
nor U9927 (N_9927,N_2292,N_2736);
nor U9928 (N_9928,N_5737,N_892);
nand U9929 (N_9929,N_4413,N_3305);
and U9930 (N_9930,N_5062,N_4553);
nor U9931 (N_9931,N_4046,N_3557);
or U9932 (N_9932,N_4995,N_5554);
and U9933 (N_9933,N_4490,N_3074);
or U9934 (N_9934,N_1652,N_5126);
nand U9935 (N_9935,N_3686,N_2627);
nand U9936 (N_9936,N_4568,N_1668);
nand U9937 (N_9937,N_5599,N_4626);
and U9938 (N_9938,N_4854,N_5853);
or U9939 (N_9939,N_4678,N_1585);
nor U9940 (N_9940,N_5912,N_4851);
nand U9941 (N_9941,N_1702,N_472);
nor U9942 (N_9942,N_5424,N_3832);
and U9943 (N_9943,N_1704,N_3556);
or U9944 (N_9944,N_3958,N_4888);
or U9945 (N_9945,N_5950,N_3441);
or U9946 (N_9946,N_458,N_5487);
nor U9947 (N_9947,N_3484,N_1428);
and U9948 (N_9948,N_5974,N_5174);
or U9949 (N_9949,N_2057,N_794);
and U9950 (N_9950,N_476,N_6137);
nand U9951 (N_9951,N_332,N_934);
or U9952 (N_9952,N_1053,N_2762);
and U9953 (N_9953,N_3573,N_5294);
nand U9954 (N_9954,N_4794,N_160);
nand U9955 (N_9955,N_3282,N_478);
nor U9956 (N_9956,N_5976,N_3051);
nor U9957 (N_9957,N_5308,N_3550);
or U9958 (N_9958,N_4742,N_5842);
nand U9959 (N_9959,N_4497,N_1470);
nand U9960 (N_9960,N_5974,N_4192);
nor U9961 (N_9961,N_3309,N_1616);
or U9962 (N_9962,N_723,N_1613);
nor U9963 (N_9963,N_4960,N_2280);
xor U9964 (N_9964,N_5920,N_2374);
and U9965 (N_9965,N_6245,N_129);
nor U9966 (N_9966,N_4384,N_612);
nand U9967 (N_9967,N_239,N_2969);
and U9968 (N_9968,N_3413,N_3407);
or U9969 (N_9969,N_2502,N_5971);
and U9970 (N_9970,N_3522,N_601);
and U9971 (N_9971,N_2891,N_1990);
and U9972 (N_9972,N_6121,N_5124);
and U9973 (N_9973,N_4743,N_1646);
and U9974 (N_9974,N_4628,N_4415);
nor U9975 (N_9975,N_3822,N_3799);
nand U9976 (N_9976,N_4901,N_5435);
and U9977 (N_9977,N_3386,N_6150);
nor U9978 (N_9978,N_4837,N_3446);
xor U9979 (N_9979,N_2069,N_3759);
and U9980 (N_9980,N_648,N_0);
or U9981 (N_9981,N_3270,N_5691);
nor U9982 (N_9982,N_1617,N_3825);
and U9983 (N_9983,N_946,N_4186);
nor U9984 (N_9984,N_43,N_682);
nor U9985 (N_9985,N_945,N_5920);
or U9986 (N_9986,N_2370,N_3409);
nand U9987 (N_9987,N_3312,N_3339);
or U9988 (N_9988,N_3446,N_466);
and U9989 (N_9989,N_3721,N_933);
nand U9990 (N_9990,N_2336,N_2848);
nor U9991 (N_9991,N_4604,N_2357);
nor U9992 (N_9992,N_4889,N_3390);
nor U9993 (N_9993,N_1671,N_4100);
nor U9994 (N_9994,N_5085,N_81);
nand U9995 (N_9995,N_5284,N_4962);
or U9996 (N_9996,N_1546,N_2894);
and U9997 (N_9997,N_4000,N_5060);
and U9998 (N_9998,N_733,N_2868);
nor U9999 (N_9999,N_2825,N_3966);
nand U10000 (N_10000,N_3580,N_2992);
and U10001 (N_10001,N_2956,N_714);
or U10002 (N_10002,N_3353,N_901);
and U10003 (N_10003,N_4026,N_5723);
nand U10004 (N_10004,N_4114,N_430);
nand U10005 (N_10005,N_448,N_5011);
and U10006 (N_10006,N_1267,N_2957);
and U10007 (N_10007,N_514,N_5841);
nor U10008 (N_10008,N_1307,N_6189);
nor U10009 (N_10009,N_4780,N_5619);
nor U10010 (N_10010,N_4639,N_81);
or U10011 (N_10011,N_5724,N_997);
and U10012 (N_10012,N_4464,N_1541);
or U10013 (N_10013,N_425,N_6129);
nor U10014 (N_10014,N_2640,N_6188);
and U10015 (N_10015,N_4364,N_1999);
and U10016 (N_10016,N_5667,N_3917);
nand U10017 (N_10017,N_6161,N_2615);
nand U10018 (N_10018,N_1638,N_2423);
nand U10019 (N_10019,N_776,N_827);
nand U10020 (N_10020,N_392,N_6249);
nand U10021 (N_10021,N_5354,N_4771);
nor U10022 (N_10022,N_120,N_1520);
and U10023 (N_10023,N_3975,N_41);
or U10024 (N_10024,N_5595,N_2242);
nor U10025 (N_10025,N_2276,N_1170);
or U10026 (N_10026,N_2063,N_3669);
and U10027 (N_10027,N_5007,N_5217);
and U10028 (N_10028,N_2581,N_1865);
and U10029 (N_10029,N_1011,N_5023);
nand U10030 (N_10030,N_2368,N_4745);
or U10031 (N_10031,N_1062,N_1893);
and U10032 (N_10032,N_4381,N_2076);
nand U10033 (N_10033,N_3003,N_1077);
nand U10034 (N_10034,N_2396,N_5500);
nand U10035 (N_10035,N_871,N_2116);
nor U10036 (N_10036,N_396,N_1776);
and U10037 (N_10037,N_2010,N_3186);
or U10038 (N_10038,N_1234,N_206);
nand U10039 (N_10039,N_786,N_3824);
nor U10040 (N_10040,N_5844,N_2080);
or U10041 (N_10041,N_1265,N_5425);
and U10042 (N_10042,N_3954,N_2721);
and U10043 (N_10043,N_1739,N_2384);
nor U10044 (N_10044,N_5162,N_4150);
or U10045 (N_10045,N_5986,N_2793);
and U10046 (N_10046,N_3106,N_3989);
xnor U10047 (N_10047,N_1931,N_5395);
and U10048 (N_10048,N_3795,N_4452);
nand U10049 (N_10049,N_3244,N_4321);
nand U10050 (N_10050,N_2313,N_5425);
and U10051 (N_10051,N_2308,N_3994);
nor U10052 (N_10052,N_636,N_1576);
nand U10053 (N_10053,N_5673,N_825);
nor U10054 (N_10054,N_1916,N_3520);
nor U10055 (N_10055,N_4887,N_923);
nand U10056 (N_10056,N_3449,N_3662);
and U10057 (N_10057,N_3863,N_2145);
nand U10058 (N_10058,N_521,N_2374);
and U10059 (N_10059,N_3020,N_567);
nor U10060 (N_10060,N_4160,N_5841);
nand U10061 (N_10061,N_6048,N_3284);
nand U10062 (N_10062,N_1092,N_4092);
or U10063 (N_10063,N_5946,N_3803);
nor U10064 (N_10064,N_5921,N_5900);
and U10065 (N_10065,N_1811,N_4094);
or U10066 (N_10066,N_4646,N_3063);
nand U10067 (N_10067,N_1634,N_5201);
nand U10068 (N_10068,N_2167,N_368);
and U10069 (N_10069,N_4074,N_5784);
and U10070 (N_10070,N_4190,N_4596);
nand U10071 (N_10071,N_4867,N_1416);
and U10072 (N_10072,N_2057,N_4144);
nand U10073 (N_10073,N_268,N_1967);
and U10074 (N_10074,N_4695,N_2385);
or U10075 (N_10075,N_899,N_5391);
or U10076 (N_10076,N_4842,N_1982);
nand U10077 (N_10077,N_915,N_5701);
and U10078 (N_10078,N_3707,N_377);
nand U10079 (N_10079,N_2301,N_2566);
or U10080 (N_10080,N_5764,N_4556);
nor U10081 (N_10081,N_2391,N_5557);
and U10082 (N_10082,N_519,N_3507);
and U10083 (N_10083,N_5700,N_1200);
and U10084 (N_10084,N_3735,N_5015);
and U10085 (N_10085,N_4607,N_3843);
and U10086 (N_10086,N_1678,N_2417);
or U10087 (N_10087,N_319,N_4628);
nor U10088 (N_10088,N_3511,N_2779);
nor U10089 (N_10089,N_673,N_2245);
and U10090 (N_10090,N_1936,N_2789);
or U10091 (N_10091,N_4494,N_2883);
nand U10092 (N_10092,N_3660,N_2246);
nor U10093 (N_10093,N_973,N_5162);
nand U10094 (N_10094,N_3215,N_5177);
or U10095 (N_10095,N_821,N_2341);
or U10096 (N_10096,N_5969,N_800);
or U10097 (N_10097,N_2249,N_3048);
nor U10098 (N_10098,N_6205,N_2637);
or U10099 (N_10099,N_4656,N_1134);
nor U10100 (N_10100,N_3857,N_2726);
and U10101 (N_10101,N_2062,N_4873);
and U10102 (N_10102,N_6243,N_6235);
nand U10103 (N_10103,N_4235,N_596);
nor U10104 (N_10104,N_3789,N_4807);
or U10105 (N_10105,N_6120,N_1333);
nand U10106 (N_10106,N_2593,N_1242);
and U10107 (N_10107,N_4555,N_3726);
and U10108 (N_10108,N_2123,N_6194);
nand U10109 (N_10109,N_3019,N_3203);
or U10110 (N_10110,N_4347,N_4650);
nand U10111 (N_10111,N_5954,N_3778);
nand U10112 (N_10112,N_5336,N_6217);
and U10113 (N_10113,N_4105,N_1175);
nand U10114 (N_10114,N_6128,N_1519);
or U10115 (N_10115,N_2547,N_3930);
and U10116 (N_10116,N_5097,N_5912);
nand U10117 (N_10117,N_812,N_3190);
nor U10118 (N_10118,N_5292,N_4463);
and U10119 (N_10119,N_4812,N_5812);
or U10120 (N_10120,N_1882,N_1154);
or U10121 (N_10121,N_4023,N_4493);
nor U10122 (N_10122,N_860,N_95);
or U10123 (N_10123,N_2929,N_3343);
nor U10124 (N_10124,N_2377,N_3327);
nand U10125 (N_10125,N_895,N_449);
nor U10126 (N_10126,N_3409,N_2013);
nor U10127 (N_10127,N_3174,N_459);
or U10128 (N_10128,N_3508,N_101);
or U10129 (N_10129,N_2689,N_350);
nand U10130 (N_10130,N_2126,N_3810);
xnor U10131 (N_10131,N_5611,N_4515);
and U10132 (N_10132,N_1995,N_2655);
and U10133 (N_10133,N_429,N_3930);
or U10134 (N_10134,N_2051,N_507);
or U10135 (N_10135,N_4324,N_3409);
nor U10136 (N_10136,N_4519,N_440);
and U10137 (N_10137,N_2511,N_2826);
and U10138 (N_10138,N_5140,N_341);
nor U10139 (N_10139,N_5087,N_3101);
and U10140 (N_10140,N_448,N_2592);
nor U10141 (N_10141,N_1727,N_3359);
or U10142 (N_10142,N_1794,N_1541);
and U10143 (N_10143,N_6184,N_974);
and U10144 (N_10144,N_1007,N_3508);
nand U10145 (N_10145,N_2916,N_2806);
nand U10146 (N_10146,N_2695,N_2581);
nor U10147 (N_10147,N_6076,N_6194);
and U10148 (N_10148,N_800,N_5955);
nor U10149 (N_10149,N_1075,N_726);
or U10150 (N_10150,N_3461,N_3176);
nor U10151 (N_10151,N_5948,N_6183);
nand U10152 (N_10152,N_658,N_4538);
or U10153 (N_10153,N_5822,N_4297);
or U10154 (N_10154,N_2342,N_1719);
and U10155 (N_10155,N_5105,N_4425);
or U10156 (N_10156,N_5228,N_5651);
or U10157 (N_10157,N_614,N_4553);
and U10158 (N_10158,N_3258,N_5541);
or U10159 (N_10159,N_5783,N_2685);
nor U10160 (N_10160,N_2353,N_3031);
and U10161 (N_10161,N_5139,N_3523);
and U10162 (N_10162,N_3609,N_4983);
and U10163 (N_10163,N_4736,N_3436);
and U10164 (N_10164,N_1779,N_1594);
or U10165 (N_10165,N_5916,N_2387);
nand U10166 (N_10166,N_1427,N_2761);
or U10167 (N_10167,N_44,N_3544);
and U10168 (N_10168,N_2272,N_5456);
and U10169 (N_10169,N_5580,N_716);
or U10170 (N_10170,N_5099,N_1871);
nor U10171 (N_10171,N_3302,N_1512);
or U10172 (N_10172,N_6049,N_2058);
or U10173 (N_10173,N_5030,N_2937);
nand U10174 (N_10174,N_4105,N_3142);
nor U10175 (N_10175,N_2994,N_748);
and U10176 (N_10176,N_5060,N_4255);
and U10177 (N_10177,N_513,N_5601);
nand U10178 (N_10178,N_1769,N_5222);
nand U10179 (N_10179,N_1747,N_4179);
or U10180 (N_10180,N_1330,N_3458);
and U10181 (N_10181,N_5812,N_5106);
or U10182 (N_10182,N_6181,N_1059);
and U10183 (N_10183,N_694,N_4959);
or U10184 (N_10184,N_5950,N_4683);
nor U10185 (N_10185,N_5079,N_2055);
and U10186 (N_10186,N_1212,N_2856);
and U10187 (N_10187,N_1303,N_268);
nor U10188 (N_10188,N_6112,N_1100);
nor U10189 (N_10189,N_547,N_4265);
nand U10190 (N_10190,N_1361,N_5009);
or U10191 (N_10191,N_4519,N_766);
nand U10192 (N_10192,N_3952,N_2877);
nor U10193 (N_10193,N_192,N_4538);
or U10194 (N_10194,N_5032,N_480);
nand U10195 (N_10195,N_83,N_2915);
nor U10196 (N_10196,N_617,N_3171);
or U10197 (N_10197,N_2725,N_2906);
nand U10198 (N_10198,N_3027,N_3456);
or U10199 (N_10199,N_2511,N_4293);
or U10200 (N_10200,N_3951,N_4633);
nand U10201 (N_10201,N_0,N_4664);
or U10202 (N_10202,N_602,N_1645);
nand U10203 (N_10203,N_4795,N_3897);
and U10204 (N_10204,N_4993,N_4874);
and U10205 (N_10205,N_5895,N_2146);
and U10206 (N_10206,N_934,N_1254);
nand U10207 (N_10207,N_2466,N_2045);
nand U10208 (N_10208,N_4521,N_1089);
and U10209 (N_10209,N_4478,N_1218);
nand U10210 (N_10210,N_3768,N_4319);
xor U10211 (N_10211,N_3422,N_2181);
nand U10212 (N_10212,N_571,N_2567);
xor U10213 (N_10213,N_1902,N_3473);
nor U10214 (N_10214,N_2115,N_5656);
or U10215 (N_10215,N_5181,N_1102);
nor U10216 (N_10216,N_3790,N_2282);
nand U10217 (N_10217,N_6127,N_3860);
nor U10218 (N_10218,N_1273,N_1036);
nor U10219 (N_10219,N_2342,N_1715);
nand U10220 (N_10220,N_3253,N_3690);
nor U10221 (N_10221,N_1557,N_467);
nor U10222 (N_10222,N_1813,N_5379);
and U10223 (N_10223,N_2965,N_4658);
nand U10224 (N_10224,N_5980,N_2469);
and U10225 (N_10225,N_1848,N_4437);
or U10226 (N_10226,N_3102,N_3326);
and U10227 (N_10227,N_3838,N_5609);
nand U10228 (N_10228,N_1924,N_4464);
or U10229 (N_10229,N_4044,N_3844);
or U10230 (N_10230,N_3257,N_5011);
and U10231 (N_10231,N_4192,N_1251);
and U10232 (N_10232,N_5519,N_3369);
nor U10233 (N_10233,N_5957,N_4175);
and U10234 (N_10234,N_4327,N_860);
and U10235 (N_10235,N_2515,N_4079);
and U10236 (N_10236,N_4535,N_2285);
nand U10237 (N_10237,N_793,N_2191);
and U10238 (N_10238,N_5107,N_689);
or U10239 (N_10239,N_3679,N_5734);
and U10240 (N_10240,N_4503,N_4821);
and U10241 (N_10241,N_2736,N_2801);
or U10242 (N_10242,N_2477,N_4216);
nand U10243 (N_10243,N_2696,N_260);
nor U10244 (N_10244,N_2114,N_4730);
and U10245 (N_10245,N_1181,N_1492);
nor U10246 (N_10246,N_3917,N_5544);
nand U10247 (N_10247,N_3101,N_4215);
xnor U10248 (N_10248,N_5961,N_1124);
or U10249 (N_10249,N_5081,N_5519);
nor U10250 (N_10250,N_6208,N_1475);
nand U10251 (N_10251,N_0,N_1761);
and U10252 (N_10252,N_5348,N_4063);
nor U10253 (N_10253,N_4279,N_5898);
or U10254 (N_10254,N_4911,N_5551);
and U10255 (N_10255,N_4703,N_1241);
nand U10256 (N_10256,N_2533,N_604);
and U10257 (N_10257,N_1784,N_2551);
and U10258 (N_10258,N_4919,N_1160);
nor U10259 (N_10259,N_1842,N_76);
nand U10260 (N_10260,N_2811,N_1951);
and U10261 (N_10261,N_5390,N_462);
nand U10262 (N_10262,N_772,N_5905);
nand U10263 (N_10263,N_6155,N_5425);
or U10264 (N_10264,N_4034,N_5410);
and U10265 (N_10265,N_3335,N_3284);
or U10266 (N_10266,N_4314,N_4869);
or U10267 (N_10267,N_3140,N_4400);
nor U10268 (N_10268,N_488,N_6209);
or U10269 (N_10269,N_1577,N_531);
and U10270 (N_10270,N_5761,N_6203);
and U10271 (N_10271,N_5303,N_219);
nand U10272 (N_10272,N_670,N_802);
nor U10273 (N_10273,N_6032,N_2409);
nand U10274 (N_10274,N_2021,N_573);
nor U10275 (N_10275,N_2540,N_2444);
nand U10276 (N_10276,N_7,N_908);
or U10277 (N_10277,N_551,N_2985);
and U10278 (N_10278,N_1521,N_1871);
nor U10279 (N_10279,N_810,N_3277);
nand U10280 (N_10280,N_825,N_5397);
and U10281 (N_10281,N_220,N_1233);
and U10282 (N_10282,N_1822,N_85);
nor U10283 (N_10283,N_4118,N_3344);
nand U10284 (N_10284,N_1871,N_4331);
or U10285 (N_10285,N_2253,N_1117);
nand U10286 (N_10286,N_4358,N_918);
and U10287 (N_10287,N_3677,N_5790);
nor U10288 (N_10288,N_3388,N_2234);
and U10289 (N_10289,N_158,N_235);
nand U10290 (N_10290,N_4005,N_991);
and U10291 (N_10291,N_4339,N_5610);
nor U10292 (N_10292,N_4277,N_4999);
and U10293 (N_10293,N_4667,N_2587);
and U10294 (N_10294,N_2216,N_5549);
nor U10295 (N_10295,N_585,N_543);
and U10296 (N_10296,N_2745,N_5095);
nand U10297 (N_10297,N_1503,N_5652);
nor U10298 (N_10298,N_4321,N_4969);
nor U10299 (N_10299,N_5364,N_2944);
nand U10300 (N_10300,N_5145,N_912);
nor U10301 (N_10301,N_6212,N_1408);
or U10302 (N_10302,N_1263,N_1711);
or U10303 (N_10303,N_3691,N_6194);
nor U10304 (N_10304,N_3789,N_2423);
and U10305 (N_10305,N_1552,N_4259);
or U10306 (N_10306,N_6070,N_6084);
nand U10307 (N_10307,N_6113,N_5825);
nand U10308 (N_10308,N_2010,N_5707);
nand U10309 (N_10309,N_5137,N_5764);
and U10310 (N_10310,N_5402,N_6185);
nor U10311 (N_10311,N_4563,N_5874);
nand U10312 (N_10312,N_5891,N_4997);
nor U10313 (N_10313,N_3890,N_4501);
nor U10314 (N_10314,N_5554,N_1035);
or U10315 (N_10315,N_6128,N_839);
and U10316 (N_10316,N_2759,N_721);
nand U10317 (N_10317,N_2155,N_4010);
nor U10318 (N_10318,N_3403,N_2994);
nand U10319 (N_10319,N_3439,N_3627);
or U10320 (N_10320,N_5669,N_2703);
and U10321 (N_10321,N_5242,N_506);
or U10322 (N_10322,N_3370,N_2620);
or U10323 (N_10323,N_2186,N_4507);
nand U10324 (N_10324,N_5954,N_345);
or U10325 (N_10325,N_6201,N_2892);
nor U10326 (N_10326,N_6145,N_5730);
or U10327 (N_10327,N_6047,N_1450);
nor U10328 (N_10328,N_394,N_1403);
or U10329 (N_10329,N_462,N_1238);
and U10330 (N_10330,N_890,N_1442);
nor U10331 (N_10331,N_4343,N_1823);
and U10332 (N_10332,N_2484,N_3856);
and U10333 (N_10333,N_2169,N_4014);
or U10334 (N_10334,N_1007,N_3589);
and U10335 (N_10335,N_1912,N_3417);
and U10336 (N_10336,N_5927,N_5539);
nor U10337 (N_10337,N_3020,N_118);
nor U10338 (N_10338,N_4694,N_107);
or U10339 (N_10339,N_409,N_5089);
or U10340 (N_10340,N_3191,N_6113);
or U10341 (N_10341,N_1733,N_3494);
nand U10342 (N_10342,N_1320,N_1533);
and U10343 (N_10343,N_4404,N_5038);
nand U10344 (N_10344,N_5499,N_5523);
nor U10345 (N_10345,N_5986,N_3584);
and U10346 (N_10346,N_4552,N_959);
or U10347 (N_10347,N_816,N_3560);
or U10348 (N_10348,N_2032,N_916);
nand U10349 (N_10349,N_130,N_13);
nor U10350 (N_10350,N_2938,N_3203);
and U10351 (N_10351,N_6111,N_1820);
nor U10352 (N_10352,N_3603,N_3338);
or U10353 (N_10353,N_5025,N_14);
and U10354 (N_10354,N_1021,N_4064);
nor U10355 (N_10355,N_2987,N_3727);
or U10356 (N_10356,N_509,N_4870);
nand U10357 (N_10357,N_34,N_5047);
or U10358 (N_10358,N_3076,N_6152);
nor U10359 (N_10359,N_1466,N_5952);
and U10360 (N_10360,N_3856,N_3883);
nor U10361 (N_10361,N_4730,N_68);
or U10362 (N_10362,N_766,N_4620);
and U10363 (N_10363,N_1569,N_889);
nor U10364 (N_10364,N_1533,N_2304);
nor U10365 (N_10365,N_2845,N_1869);
nand U10366 (N_10366,N_4870,N_4621);
nand U10367 (N_10367,N_4456,N_1697);
nor U10368 (N_10368,N_4528,N_3645);
nand U10369 (N_10369,N_1947,N_4116);
and U10370 (N_10370,N_5639,N_1338);
nor U10371 (N_10371,N_2532,N_2666);
and U10372 (N_10372,N_4873,N_2037);
or U10373 (N_10373,N_2500,N_3533);
and U10374 (N_10374,N_4489,N_5103);
xor U10375 (N_10375,N_1509,N_5859);
nor U10376 (N_10376,N_3892,N_3324);
nand U10377 (N_10377,N_5266,N_3788);
or U10378 (N_10378,N_2993,N_1816);
and U10379 (N_10379,N_1281,N_1565);
or U10380 (N_10380,N_5390,N_5083);
nand U10381 (N_10381,N_1103,N_3377);
and U10382 (N_10382,N_5909,N_1687);
nor U10383 (N_10383,N_569,N_1818);
and U10384 (N_10384,N_2225,N_544);
or U10385 (N_10385,N_5976,N_3487);
and U10386 (N_10386,N_1943,N_1918);
nand U10387 (N_10387,N_1707,N_2967);
or U10388 (N_10388,N_5973,N_2856);
nor U10389 (N_10389,N_5729,N_3846);
and U10390 (N_10390,N_5867,N_2649);
nand U10391 (N_10391,N_3902,N_6193);
nand U10392 (N_10392,N_719,N_2989);
nor U10393 (N_10393,N_4847,N_2548);
nand U10394 (N_10394,N_259,N_1636);
and U10395 (N_10395,N_2961,N_2922);
nor U10396 (N_10396,N_1552,N_1398);
or U10397 (N_10397,N_3329,N_2901);
and U10398 (N_10398,N_4484,N_2443);
nor U10399 (N_10399,N_611,N_4671);
nor U10400 (N_10400,N_1205,N_4543);
nand U10401 (N_10401,N_2108,N_6141);
or U10402 (N_10402,N_3438,N_1126);
and U10403 (N_10403,N_4980,N_4096);
and U10404 (N_10404,N_3370,N_4365);
nor U10405 (N_10405,N_1067,N_3102);
nor U10406 (N_10406,N_3775,N_2340);
nor U10407 (N_10407,N_4995,N_3335);
and U10408 (N_10408,N_337,N_3313);
nor U10409 (N_10409,N_478,N_3943);
nand U10410 (N_10410,N_4688,N_3815);
or U10411 (N_10411,N_2307,N_5225);
and U10412 (N_10412,N_4083,N_2986);
nand U10413 (N_10413,N_1446,N_4474);
nor U10414 (N_10414,N_1522,N_4314);
nand U10415 (N_10415,N_5733,N_4269);
or U10416 (N_10416,N_1398,N_5745);
nor U10417 (N_10417,N_5928,N_5069);
and U10418 (N_10418,N_862,N_6035);
and U10419 (N_10419,N_668,N_4941);
nand U10420 (N_10420,N_50,N_5758);
nor U10421 (N_10421,N_2481,N_3639);
nand U10422 (N_10422,N_5911,N_1955);
nand U10423 (N_10423,N_1188,N_1538);
nand U10424 (N_10424,N_2102,N_655);
and U10425 (N_10425,N_6022,N_1494);
and U10426 (N_10426,N_149,N_3245);
nand U10427 (N_10427,N_4641,N_3014);
nor U10428 (N_10428,N_286,N_2420);
and U10429 (N_10429,N_6214,N_262);
nand U10430 (N_10430,N_3784,N_208);
or U10431 (N_10431,N_5329,N_2104);
nand U10432 (N_10432,N_3853,N_4921);
nor U10433 (N_10433,N_703,N_6054);
nand U10434 (N_10434,N_1436,N_2465);
nand U10435 (N_10435,N_6131,N_2741);
or U10436 (N_10436,N_5201,N_5271);
and U10437 (N_10437,N_2745,N_5709);
or U10438 (N_10438,N_5578,N_3338);
and U10439 (N_10439,N_5853,N_3918);
nand U10440 (N_10440,N_2064,N_5431);
and U10441 (N_10441,N_5054,N_1579);
and U10442 (N_10442,N_4635,N_1241);
and U10443 (N_10443,N_3625,N_309);
nor U10444 (N_10444,N_4944,N_5939);
or U10445 (N_10445,N_1767,N_4428);
nand U10446 (N_10446,N_4454,N_4484);
xnor U10447 (N_10447,N_2623,N_2863);
or U10448 (N_10448,N_3964,N_4136);
or U10449 (N_10449,N_4757,N_1042);
and U10450 (N_10450,N_4241,N_3374);
or U10451 (N_10451,N_2965,N_6148);
nor U10452 (N_10452,N_576,N_212);
nand U10453 (N_10453,N_1431,N_5374);
nor U10454 (N_10454,N_5994,N_765);
or U10455 (N_10455,N_2839,N_384);
and U10456 (N_10456,N_1890,N_3354);
nor U10457 (N_10457,N_844,N_1291);
or U10458 (N_10458,N_630,N_3490);
nand U10459 (N_10459,N_5261,N_4178);
nand U10460 (N_10460,N_2803,N_4662);
and U10461 (N_10461,N_4267,N_1049);
or U10462 (N_10462,N_5837,N_394);
or U10463 (N_10463,N_6187,N_177);
nand U10464 (N_10464,N_3205,N_1857);
or U10465 (N_10465,N_1598,N_4294);
nand U10466 (N_10466,N_2109,N_2587);
and U10467 (N_10467,N_292,N_5043);
nand U10468 (N_10468,N_1731,N_5879);
and U10469 (N_10469,N_5717,N_799);
nor U10470 (N_10470,N_1706,N_2379);
and U10471 (N_10471,N_4884,N_3094);
xor U10472 (N_10472,N_992,N_4132);
nor U10473 (N_10473,N_3088,N_3823);
nor U10474 (N_10474,N_1786,N_5978);
or U10475 (N_10475,N_2012,N_4200);
and U10476 (N_10476,N_3411,N_3239);
or U10477 (N_10477,N_3344,N_3366);
or U10478 (N_10478,N_4559,N_4626);
or U10479 (N_10479,N_1149,N_962);
and U10480 (N_10480,N_4145,N_2213);
nor U10481 (N_10481,N_851,N_5715);
or U10482 (N_10482,N_10,N_5277);
or U10483 (N_10483,N_4870,N_2755);
or U10484 (N_10484,N_5122,N_5162);
nor U10485 (N_10485,N_3071,N_1570);
nand U10486 (N_10486,N_2410,N_4608);
nor U10487 (N_10487,N_4723,N_34);
nand U10488 (N_10488,N_1521,N_5706);
nor U10489 (N_10489,N_1293,N_2652);
and U10490 (N_10490,N_5786,N_2019);
nand U10491 (N_10491,N_3346,N_872);
nor U10492 (N_10492,N_6223,N_6150);
nand U10493 (N_10493,N_5442,N_2044);
nand U10494 (N_10494,N_1772,N_350);
or U10495 (N_10495,N_935,N_1667);
and U10496 (N_10496,N_3584,N_3707);
and U10497 (N_10497,N_4994,N_5726);
and U10498 (N_10498,N_2772,N_3062);
or U10499 (N_10499,N_4677,N_385);
and U10500 (N_10500,N_2732,N_1175);
and U10501 (N_10501,N_6114,N_4142);
nand U10502 (N_10502,N_4056,N_2694);
nor U10503 (N_10503,N_5798,N_800);
nor U10504 (N_10504,N_5234,N_3284);
and U10505 (N_10505,N_4277,N_3072);
nand U10506 (N_10506,N_2177,N_5577);
nor U10507 (N_10507,N_4986,N_4713);
nand U10508 (N_10508,N_1334,N_2869);
or U10509 (N_10509,N_3355,N_2519);
nand U10510 (N_10510,N_3330,N_422);
and U10511 (N_10511,N_2659,N_2946);
or U10512 (N_10512,N_1479,N_1264);
and U10513 (N_10513,N_4741,N_6118);
nand U10514 (N_10514,N_4422,N_5595);
and U10515 (N_10515,N_4971,N_406);
and U10516 (N_10516,N_1548,N_1105);
and U10517 (N_10517,N_3677,N_3724);
and U10518 (N_10518,N_2428,N_4523);
nor U10519 (N_10519,N_1587,N_3347);
nand U10520 (N_10520,N_4550,N_4320);
nor U10521 (N_10521,N_4175,N_1418);
nand U10522 (N_10522,N_5262,N_5572);
or U10523 (N_10523,N_1394,N_6093);
and U10524 (N_10524,N_1593,N_1225);
and U10525 (N_10525,N_1249,N_5914);
or U10526 (N_10526,N_4101,N_3937);
and U10527 (N_10527,N_5795,N_1675);
nand U10528 (N_10528,N_3477,N_3274);
nor U10529 (N_10529,N_2582,N_5238);
or U10530 (N_10530,N_2967,N_1861);
nand U10531 (N_10531,N_2597,N_2916);
or U10532 (N_10532,N_889,N_1347);
and U10533 (N_10533,N_1339,N_6177);
or U10534 (N_10534,N_5852,N_5181);
nor U10535 (N_10535,N_1089,N_2255);
nor U10536 (N_10536,N_1909,N_810);
nand U10537 (N_10537,N_959,N_5529);
or U10538 (N_10538,N_5394,N_1345);
nand U10539 (N_10539,N_3640,N_4676);
or U10540 (N_10540,N_3459,N_3246);
and U10541 (N_10541,N_781,N_4487);
and U10542 (N_10542,N_679,N_5613);
nand U10543 (N_10543,N_1935,N_2181);
and U10544 (N_10544,N_4669,N_4044);
nand U10545 (N_10545,N_4355,N_1166);
nand U10546 (N_10546,N_4276,N_3969);
nor U10547 (N_10547,N_4083,N_3630);
nor U10548 (N_10548,N_2447,N_3377);
and U10549 (N_10549,N_863,N_5241);
or U10550 (N_10550,N_2712,N_3393);
or U10551 (N_10551,N_4034,N_1994);
nand U10552 (N_10552,N_5223,N_1115);
or U10553 (N_10553,N_2504,N_3477);
or U10554 (N_10554,N_674,N_2272);
or U10555 (N_10555,N_1196,N_924);
nand U10556 (N_10556,N_5447,N_1392);
or U10557 (N_10557,N_83,N_3171);
and U10558 (N_10558,N_5575,N_2423);
or U10559 (N_10559,N_876,N_4578);
or U10560 (N_10560,N_4004,N_4325);
nand U10561 (N_10561,N_3181,N_1028);
nand U10562 (N_10562,N_5052,N_5810);
nor U10563 (N_10563,N_1409,N_2063);
nand U10564 (N_10564,N_4544,N_3858);
or U10565 (N_10565,N_1632,N_3915);
and U10566 (N_10566,N_1437,N_4075);
nor U10567 (N_10567,N_3889,N_167);
and U10568 (N_10568,N_5452,N_1775);
nor U10569 (N_10569,N_5075,N_3913);
or U10570 (N_10570,N_5576,N_4299);
nor U10571 (N_10571,N_3971,N_5839);
nand U10572 (N_10572,N_5073,N_6249);
nand U10573 (N_10573,N_2685,N_5743);
or U10574 (N_10574,N_6074,N_3281);
and U10575 (N_10575,N_231,N_1220);
xor U10576 (N_10576,N_1879,N_801);
nand U10577 (N_10577,N_867,N_3222);
or U10578 (N_10578,N_961,N_5935);
nor U10579 (N_10579,N_120,N_4328);
and U10580 (N_10580,N_4565,N_3341);
or U10581 (N_10581,N_1122,N_3963);
and U10582 (N_10582,N_5851,N_4306);
nand U10583 (N_10583,N_4916,N_1022);
and U10584 (N_10584,N_3026,N_2738);
nand U10585 (N_10585,N_5471,N_1367);
and U10586 (N_10586,N_170,N_5049);
or U10587 (N_10587,N_4088,N_3070);
nand U10588 (N_10588,N_4251,N_5813);
and U10589 (N_10589,N_1000,N_699);
nand U10590 (N_10590,N_5492,N_2268);
or U10591 (N_10591,N_3089,N_4129);
nor U10592 (N_10592,N_1978,N_2993);
nor U10593 (N_10593,N_1080,N_1467);
nand U10594 (N_10594,N_2579,N_1859);
or U10595 (N_10595,N_1805,N_4826);
nand U10596 (N_10596,N_4260,N_3652);
nor U10597 (N_10597,N_2241,N_3822);
nor U10598 (N_10598,N_4952,N_5934);
and U10599 (N_10599,N_2774,N_1101);
and U10600 (N_10600,N_4203,N_4197);
nand U10601 (N_10601,N_2627,N_2217);
nor U10602 (N_10602,N_6103,N_285);
nor U10603 (N_10603,N_4971,N_2684);
or U10604 (N_10604,N_3015,N_2060);
and U10605 (N_10605,N_5984,N_1335);
nand U10606 (N_10606,N_1568,N_4541);
and U10607 (N_10607,N_400,N_3461);
nor U10608 (N_10608,N_3718,N_3067);
and U10609 (N_10609,N_312,N_746);
or U10610 (N_10610,N_6165,N_4577);
nand U10611 (N_10611,N_648,N_3085);
or U10612 (N_10612,N_1660,N_3488);
nor U10613 (N_10613,N_4217,N_76);
or U10614 (N_10614,N_6043,N_5911);
and U10615 (N_10615,N_3271,N_3619);
nand U10616 (N_10616,N_3058,N_5023);
nand U10617 (N_10617,N_1998,N_208);
and U10618 (N_10618,N_2580,N_1538);
nor U10619 (N_10619,N_2911,N_5970);
and U10620 (N_10620,N_6227,N_2935);
nor U10621 (N_10621,N_4111,N_12);
and U10622 (N_10622,N_158,N_4763);
nor U10623 (N_10623,N_4507,N_3269);
or U10624 (N_10624,N_5526,N_119);
nand U10625 (N_10625,N_5660,N_1732);
nor U10626 (N_10626,N_569,N_3177);
or U10627 (N_10627,N_2745,N_5861);
nor U10628 (N_10628,N_527,N_3267);
and U10629 (N_10629,N_2504,N_3179);
nand U10630 (N_10630,N_2938,N_177);
nand U10631 (N_10631,N_3513,N_6030);
and U10632 (N_10632,N_3232,N_2408);
or U10633 (N_10633,N_3841,N_2930);
or U10634 (N_10634,N_1971,N_5762);
nor U10635 (N_10635,N_4857,N_1922);
nor U10636 (N_10636,N_5723,N_4869);
nor U10637 (N_10637,N_778,N_5910);
and U10638 (N_10638,N_3892,N_1761);
nor U10639 (N_10639,N_715,N_5607);
nand U10640 (N_10640,N_5644,N_5614);
nand U10641 (N_10641,N_3921,N_4343);
and U10642 (N_10642,N_4555,N_6132);
or U10643 (N_10643,N_4780,N_1176);
and U10644 (N_10644,N_471,N_3944);
and U10645 (N_10645,N_4026,N_4128);
nor U10646 (N_10646,N_4094,N_5714);
nand U10647 (N_10647,N_3196,N_2570);
or U10648 (N_10648,N_2227,N_2052);
or U10649 (N_10649,N_1574,N_5521);
nand U10650 (N_10650,N_5054,N_4293);
and U10651 (N_10651,N_4271,N_2783);
and U10652 (N_10652,N_2446,N_5293);
and U10653 (N_10653,N_97,N_1698);
or U10654 (N_10654,N_353,N_5674);
or U10655 (N_10655,N_5828,N_3104);
nand U10656 (N_10656,N_1376,N_5222);
nor U10657 (N_10657,N_384,N_3768);
and U10658 (N_10658,N_5895,N_82);
nor U10659 (N_10659,N_4215,N_1174);
or U10660 (N_10660,N_4214,N_3813);
or U10661 (N_10661,N_5510,N_2492);
nor U10662 (N_10662,N_559,N_4787);
or U10663 (N_10663,N_3850,N_1956);
and U10664 (N_10664,N_972,N_5759);
nand U10665 (N_10665,N_2324,N_588);
xor U10666 (N_10666,N_1607,N_4730);
nand U10667 (N_10667,N_4572,N_4356);
nor U10668 (N_10668,N_340,N_553);
and U10669 (N_10669,N_5646,N_1345);
nor U10670 (N_10670,N_2042,N_932);
and U10671 (N_10671,N_5359,N_2586);
nand U10672 (N_10672,N_3265,N_2595);
and U10673 (N_10673,N_114,N_984);
or U10674 (N_10674,N_4812,N_4672);
nor U10675 (N_10675,N_1793,N_2117);
and U10676 (N_10676,N_5160,N_4648);
and U10677 (N_10677,N_3607,N_2058);
nor U10678 (N_10678,N_4622,N_867);
or U10679 (N_10679,N_3219,N_728);
or U10680 (N_10680,N_4341,N_1463);
nand U10681 (N_10681,N_4724,N_3419);
or U10682 (N_10682,N_4599,N_6184);
or U10683 (N_10683,N_1860,N_5322);
and U10684 (N_10684,N_4069,N_5378);
and U10685 (N_10685,N_2886,N_4327);
or U10686 (N_10686,N_1165,N_476);
nor U10687 (N_10687,N_5635,N_4045);
and U10688 (N_10688,N_723,N_4532);
nor U10689 (N_10689,N_5215,N_5493);
nor U10690 (N_10690,N_2743,N_5987);
nor U10691 (N_10691,N_1399,N_2521);
or U10692 (N_10692,N_1966,N_2558);
nand U10693 (N_10693,N_4047,N_3235);
nand U10694 (N_10694,N_5749,N_5688);
nor U10695 (N_10695,N_1357,N_4109);
nand U10696 (N_10696,N_1137,N_1361);
or U10697 (N_10697,N_2663,N_5210);
and U10698 (N_10698,N_164,N_4657);
or U10699 (N_10699,N_183,N_4229);
or U10700 (N_10700,N_4793,N_4936);
nand U10701 (N_10701,N_1705,N_2608);
or U10702 (N_10702,N_3875,N_2638);
and U10703 (N_10703,N_6027,N_733);
nor U10704 (N_10704,N_2290,N_6248);
or U10705 (N_10705,N_4274,N_1113);
nand U10706 (N_10706,N_1095,N_5588);
or U10707 (N_10707,N_627,N_2859);
nor U10708 (N_10708,N_2753,N_4725);
nand U10709 (N_10709,N_592,N_1228);
or U10710 (N_10710,N_4649,N_4933);
and U10711 (N_10711,N_2185,N_1296);
nand U10712 (N_10712,N_1878,N_3731);
nand U10713 (N_10713,N_5346,N_2304);
nand U10714 (N_10714,N_4767,N_473);
nand U10715 (N_10715,N_1865,N_840);
or U10716 (N_10716,N_484,N_4716);
and U10717 (N_10717,N_5480,N_4969);
and U10718 (N_10718,N_4850,N_5401);
or U10719 (N_10719,N_4073,N_1397);
nor U10720 (N_10720,N_2317,N_319);
nor U10721 (N_10721,N_3850,N_3275);
nor U10722 (N_10722,N_2395,N_309);
or U10723 (N_10723,N_389,N_747);
and U10724 (N_10724,N_2310,N_2192);
or U10725 (N_10725,N_508,N_2253);
and U10726 (N_10726,N_1994,N_4412);
nor U10727 (N_10727,N_783,N_1483);
and U10728 (N_10728,N_1994,N_1117);
nand U10729 (N_10729,N_2432,N_3677);
nor U10730 (N_10730,N_3515,N_1757);
or U10731 (N_10731,N_4814,N_2226);
or U10732 (N_10732,N_3810,N_984);
or U10733 (N_10733,N_5143,N_3169);
nand U10734 (N_10734,N_2060,N_4417);
nand U10735 (N_10735,N_127,N_60);
nor U10736 (N_10736,N_4187,N_5066);
nand U10737 (N_10737,N_6007,N_2558);
and U10738 (N_10738,N_5527,N_5668);
nand U10739 (N_10739,N_916,N_5083);
and U10740 (N_10740,N_5492,N_3408);
and U10741 (N_10741,N_5380,N_1831);
nor U10742 (N_10742,N_2019,N_1514);
and U10743 (N_10743,N_343,N_6037);
nor U10744 (N_10744,N_4462,N_1762);
and U10745 (N_10745,N_1452,N_2186);
nand U10746 (N_10746,N_6116,N_3370);
and U10747 (N_10747,N_5530,N_5290);
or U10748 (N_10748,N_1789,N_1590);
nand U10749 (N_10749,N_937,N_1521);
nand U10750 (N_10750,N_4864,N_6053);
nand U10751 (N_10751,N_2472,N_3223);
or U10752 (N_10752,N_1350,N_4097);
nand U10753 (N_10753,N_4741,N_4306);
or U10754 (N_10754,N_4794,N_3419);
and U10755 (N_10755,N_2070,N_2711);
nand U10756 (N_10756,N_2868,N_1067);
or U10757 (N_10757,N_221,N_3631);
and U10758 (N_10758,N_1113,N_4737);
or U10759 (N_10759,N_4409,N_3898);
and U10760 (N_10760,N_4352,N_160);
nand U10761 (N_10761,N_368,N_2214);
nor U10762 (N_10762,N_943,N_2305);
nor U10763 (N_10763,N_5904,N_2071);
and U10764 (N_10764,N_5222,N_3313);
or U10765 (N_10765,N_2755,N_4391);
or U10766 (N_10766,N_5596,N_544);
and U10767 (N_10767,N_804,N_6084);
nor U10768 (N_10768,N_5886,N_4215);
nand U10769 (N_10769,N_3072,N_5942);
nand U10770 (N_10770,N_2859,N_1849);
or U10771 (N_10771,N_4448,N_431);
and U10772 (N_10772,N_4903,N_1091);
nor U10773 (N_10773,N_3196,N_699);
nor U10774 (N_10774,N_154,N_2462);
and U10775 (N_10775,N_2535,N_4752);
and U10776 (N_10776,N_5915,N_5994);
nand U10777 (N_10777,N_3947,N_2009);
nand U10778 (N_10778,N_4801,N_3693);
or U10779 (N_10779,N_1629,N_6041);
or U10780 (N_10780,N_1265,N_4819);
nand U10781 (N_10781,N_5022,N_2051);
and U10782 (N_10782,N_5083,N_1667);
and U10783 (N_10783,N_1207,N_4350);
or U10784 (N_10784,N_295,N_3731);
and U10785 (N_10785,N_5480,N_5639);
or U10786 (N_10786,N_4276,N_5107);
nand U10787 (N_10787,N_576,N_2831);
and U10788 (N_10788,N_715,N_720);
or U10789 (N_10789,N_5250,N_4222);
nand U10790 (N_10790,N_4219,N_735);
or U10791 (N_10791,N_5082,N_518);
nor U10792 (N_10792,N_1642,N_3387);
nand U10793 (N_10793,N_5356,N_1169);
nor U10794 (N_10794,N_4758,N_3799);
nand U10795 (N_10795,N_4936,N_5072);
and U10796 (N_10796,N_59,N_3477);
or U10797 (N_10797,N_3011,N_4435);
xnor U10798 (N_10798,N_2521,N_5608);
nor U10799 (N_10799,N_546,N_2080);
nor U10800 (N_10800,N_5626,N_4022);
nand U10801 (N_10801,N_1381,N_1296);
and U10802 (N_10802,N_2010,N_2874);
nand U10803 (N_10803,N_5425,N_3395);
nand U10804 (N_10804,N_2048,N_2655);
and U10805 (N_10805,N_1294,N_1468);
and U10806 (N_10806,N_1539,N_2482);
and U10807 (N_10807,N_5659,N_6019);
nand U10808 (N_10808,N_4597,N_1065);
and U10809 (N_10809,N_4227,N_1456);
and U10810 (N_10810,N_5027,N_862);
or U10811 (N_10811,N_1697,N_3200);
nor U10812 (N_10812,N_3065,N_2252);
nand U10813 (N_10813,N_869,N_3614);
or U10814 (N_10814,N_4097,N_1346);
nand U10815 (N_10815,N_4999,N_2007);
nor U10816 (N_10816,N_5392,N_566);
nor U10817 (N_10817,N_2931,N_4656);
nor U10818 (N_10818,N_1974,N_501);
or U10819 (N_10819,N_369,N_2936);
nand U10820 (N_10820,N_3136,N_5059);
nand U10821 (N_10821,N_4067,N_522);
or U10822 (N_10822,N_3752,N_2365);
nand U10823 (N_10823,N_5185,N_4883);
or U10824 (N_10824,N_4670,N_5477);
or U10825 (N_10825,N_6135,N_3454);
and U10826 (N_10826,N_4917,N_9);
nand U10827 (N_10827,N_829,N_3231);
nand U10828 (N_10828,N_5300,N_3884);
nand U10829 (N_10829,N_578,N_5149);
nor U10830 (N_10830,N_5964,N_5823);
and U10831 (N_10831,N_4351,N_5045);
nand U10832 (N_10832,N_2896,N_5628);
nor U10833 (N_10833,N_4666,N_3657);
or U10834 (N_10834,N_4936,N_3360);
nand U10835 (N_10835,N_4846,N_5042);
and U10836 (N_10836,N_3253,N_5729);
and U10837 (N_10837,N_5393,N_4056);
or U10838 (N_10838,N_4105,N_3914);
nor U10839 (N_10839,N_6076,N_2974);
and U10840 (N_10840,N_5695,N_1575);
or U10841 (N_10841,N_3384,N_1436);
and U10842 (N_10842,N_3782,N_5759);
nor U10843 (N_10843,N_6235,N_977);
and U10844 (N_10844,N_3851,N_204);
and U10845 (N_10845,N_1452,N_5159);
and U10846 (N_10846,N_5996,N_796);
and U10847 (N_10847,N_4097,N_1924);
or U10848 (N_10848,N_3585,N_5849);
and U10849 (N_10849,N_2206,N_3458);
and U10850 (N_10850,N_3565,N_5289);
and U10851 (N_10851,N_3126,N_2284);
or U10852 (N_10852,N_3915,N_4320);
nand U10853 (N_10853,N_5576,N_751);
nand U10854 (N_10854,N_1711,N_2889);
or U10855 (N_10855,N_2440,N_2557);
and U10856 (N_10856,N_785,N_1876);
nand U10857 (N_10857,N_3201,N_3948);
nor U10858 (N_10858,N_3931,N_5201);
or U10859 (N_10859,N_1268,N_3635);
nand U10860 (N_10860,N_1310,N_4024);
or U10861 (N_10861,N_2106,N_3817);
and U10862 (N_10862,N_2829,N_1266);
and U10863 (N_10863,N_940,N_4219);
nor U10864 (N_10864,N_5311,N_5762);
or U10865 (N_10865,N_3783,N_48);
nand U10866 (N_10866,N_1416,N_5763);
and U10867 (N_10867,N_906,N_2205);
nor U10868 (N_10868,N_1175,N_1559);
nand U10869 (N_10869,N_2248,N_532);
nand U10870 (N_10870,N_1808,N_358);
nand U10871 (N_10871,N_167,N_5405);
or U10872 (N_10872,N_5863,N_1028);
or U10873 (N_10873,N_1714,N_758);
and U10874 (N_10874,N_159,N_4593);
or U10875 (N_10875,N_5283,N_333);
nand U10876 (N_10876,N_3623,N_905);
nand U10877 (N_10877,N_2893,N_11);
nor U10878 (N_10878,N_1372,N_4249);
or U10879 (N_10879,N_4096,N_5426);
nand U10880 (N_10880,N_1981,N_2314);
and U10881 (N_10881,N_214,N_1565);
nand U10882 (N_10882,N_4318,N_1374);
or U10883 (N_10883,N_5417,N_3865);
nor U10884 (N_10884,N_5734,N_4761);
or U10885 (N_10885,N_167,N_5986);
and U10886 (N_10886,N_2847,N_1282);
and U10887 (N_10887,N_5025,N_1645);
nand U10888 (N_10888,N_4926,N_1409);
or U10889 (N_10889,N_4891,N_2787);
nor U10890 (N_10890,N_5989,N_5704);
nor U10891 (N_10891,N_2559,N_5677);
xor U10892 (N_10892,N_4934,N_3037);
nand U10893 (N_10893,N_3478,N_5109);
nand U10894 (N_10894,N_2840,N_3556);
nor U10895 (N_10895,N_4058,N_6161);
and U10896 (N_10896,N_1496,N_4617);
or U10897 (N_10897,N_5764,N_387);
or U10898 (N_10898,N_3315,N_1421);
nand U10899 (N_10899,N_3430,N_2273);
or U10900 (N_10900,N_3596,N_1946);
and U10901 (N_10901,N_5705,N_2912);
nor U10902 (N_10902,N_2836,N_178);
nor U10903 (N_10903,N_5445,N_2924);
nor U10904 (N_10904,N_4797,N_5042);
or U10905 (N_10905,N_3137,N_268);
or U10906 (N_10906,N_448,N_5680);
or U10907 (N_10907,N_1914,N_1579);
nand U10908 (N_10908,N_4434,N_4875);
nand U10909 (N_10909,N_1265,N_4652);
nand U10910 (N_10910,N_2544,N_6082);
nor U10911 (N_10911,N_5044,N_5319);
and U10912 (N_10912,N_2020,N_2690);
nor U10913 (N_10913,N_3600,N_5252);
and U10914 (N_10914,N_4707,N_2584);
and U10915 (N_10915,N_1824,N_258);
and U10916 (N_10916,N_730,N_2610);
and U10917 (N_10917,N_4585,N_64);
nand U10918 (N_10918,N_3417,N_5896);
and U10919 (N_10919,N_1874,N_5165);
nand U10920 (N_10920,N_1267,N_5382);
nand U10921 (N_10921,N_462,N_2904);
or U10922 (N_10922,N_4167,N_1628);
and U10923 (N_10923,N_6182,N_3881);
or U10924 (N_10924,N_599,N_4094);
nand U10925 (N_10925,N_5734,N_2383);
nor U10926 (N_10926,N_5594,N_5522);
nor U10927 (N_10927,N_1030,N_477);
and U10928 (N_10928,N_2368,N_5069);
nor U10929 (N_10929,N_303,N_5273);
nor U10930 (N_10930,N_4812,N_3524);
nor U10931 (N_10931,N_4451,N_1326);
and U10932 (N_10932,N_862,N_596);
nor U10933 (N_10933,N_5189,N_3437);
nand U10934 (N_10934,N_5412,N_4573);
nor U10935 (N_10935,N_3717,N_2270);
or U10936 (N_10936,N_2598,N_1557);
or U10937 (N_10937,N_4478,N_3157);
xor U10938 (N_10938,N_223,N_5072);
and U10939 (N_10939,N_4822,N_3280);
and U10940 (N_10940,N_4921,N_4286);
and U10941 (N_10941,N_5992,N_1642);
or U10942 (N_10942,N_3418,N_4236);
or U10943 (N_10943,N_3258,N_4090);
or U10944 (N_10944,N_234,N_5254);
and U10945 (N_10945,N_3585,N_1292);
and U10946 (N_10946,N_6214,N_635);
and U10947 (N_10947,N_185,N_5312);
and U10948 (N_10948,N_4587,N_6226);
nand U10949 (N_10949,N_955,N_4721);
and U10950 (N_10950,N_5689,N_217);
or U10951 (N_10951,N_256,N_5530);
and U10952 (N_10952,N_1212,N_42);
nand U10953 (N_10953,N_3473,N_2099);
or U10954 (N_10954,N_4114,N_696);
and U10955 (N_10955,N_586,N_3839);
nand U10956 (N_10956,N_1230,N_2054);
and U10957 (N_10957,N_46,N_644);
nand U10958 (N_10958,N_4805,N_1752);
nand U10959 (N_10959,N_3590,N_3326);
or U10960 (N_10960,N_823,N_989);
nor U10961 (N_10961,N_5083,N_4842);
or U10962 (N_10962,N_1353,N_357);
nor U10963 (N_10963,N_5729,N_96);
or U10964 (N_10964,N_1471,N_4924);
nand U10965 (N_10965,N_149,N_870);
nand U10966 (N_10966,N_1602,N_1314);
or U10967 (N_10967,N_169,N_1547);
or U10968 (N_10968,N_2831,N_4350);
nand U10969 (N_10969,N_1887,N_2310);
or U10970 (N_10970,N_1837,N_279);
nand U10971 (N_10971,N_2903,N_6205);
or U10972 (N_10972,N_4112,N_2638);
nand U10973 (N_10973,N_4452,N_4359);
nand U10974 (N_10974,N_4458,N_800);
and U10975 (N_10975,N_1089,N_3182);
and U10976 (N_10976,N_622,N_3);
nor U10977 (N_10977,N_2200,N_4045);
and U10978 (N_10978,N_4363,N_5823);
or U10979 (N_10979,N_4284,N_3012);
nor U10980 (N_10980,N_117,N_2024);
or U10981 (N_10981,N_4217,N_2229);
nor U10982 (N_10982,N_3139,N_779);
nor U10983 (N_10983,N_2508,N_3440);
and U10984 (N_10984,N_4666,N_1274);
nand U10985 (N_10985,N_4162,N_1959);
nor U10986 (N_10986,N_1969,N_2957);
nand U10987 (N_10987,N_3481,N_455);
and U10988 (N_10988,N_5681,N_1198);
nor U10989 (N_10989,N_2053,N_3132);
and U10990 (N_10990,N_3749,N_4556);
nor U10991 (N_10991,N_321,N_3083);
or U10992 (N_10992,N_1001,N_1673);
nand U10993 (N_10993,N_4769,N_3824);
nor U10994 (N_10994,N_4822,N_844);
nand U10995 (N_10995,N_4149,N_5429);
nor U10996 (N_10996,N_5132,N_568);
nand U10997 (N_10997,N_2243,N_4296);
or U10998 (N_10998,N_2541,N_6182);
nor U10999 (N_10999,N_5729,N_5927);
and U11000 (N_11000,N_3470,N_927);
xnor U11001 (N_11001,N_1916,N_5062);
and U11002 (N_11002,N_1245,N_3391);
and U11003 (N_11003,N_4772,N_4190);
nand U11004 (N_11004,N_1845,N_4811);
nand U11005 (N_11005,N_1905,N_2158);
or U11006 (N_11006,N_4197,N_6092);
nor U11007 (N_11007,N_4227,N_5028);
nor U11008 (N_11008,N_248,N_925);
or U11009 (N_11009,N_4674,N_2933);
nor U11010 (N_11010,N_6042,N_1495);
and U11011 (N_11011,N_5535,N_3801);
and U11012 (N_11012,N_273,N_4569);
nand U11013 (N_11013,N_235,N_1706);
nor U11014 (N_11014,N_1211,N_1178);
nand U11015 (N_11015,N_1931,N_378);
and U11016 (N_11016,N_3951,N_852);
or U11017 (N_11017,N_4654,N_813);
nor U11018 (N_11018,N_3986,N_4622);
nand U11019 (N_11019,N_4450,N_3557);
xor U11020 (N_11020,N_6038,N_4405);
and U11021 (N_11021,N_1703,N_4339);
nand U11022 (N_11022,N_1821,N_6061);
and U11023 (N_11023,N_499,N_5087);
or U11024 (N_11024,N_4762,N_472);
nand U11025 (N_11025,N_1458,N_4810);
nand U11026 (N_11026,N_2288,N_3164);
and U11027 (N_11027,N_1259,N_2765);
and U11028 (N_11028,N_5745,N_3636);
xnor U11029 (N_11029,N_2172,N_450);
nand U11030 (N_11030,N_647,N_5661);
nor U11031 (N_11031,N_792,N_206);
nand U11032 (N_11032,N_2107,N_2147);
nor U11033 (N_11033,N_3240,N_5);
nor U11034 (N_11034,N_1752,N_774);
and U11035 (N_11035,N_4009,N_165);
and U11036 (N_11036,N_194,N_2961);
nor U11037 (N_11037,N_1118,N_2637);
or U11038 (N_11038,N_271,N_2146);
and U11039 (N_11039,N_4077,N_6170);
or U11040 (N_11040,N_2774,N_1785);
nand U11041 (N_11041,N_4416,N_3699);
nor U11042 (N_11042,N_5221,N_2973);
nand U11043 (N_11043,N_4036,N_5655);
and U11044 (N_11044,N_1500,N_420);
or U11045 (N_11045,N_1383,N_5187);
nand U11046 (N_11046,N_4871,N_4291);
nor U11047 (N_11047,N_5901,N_4021);
and U11048 (N_11048,N_5933,N_1362);
nor U11049 (N_11049,N_5687,N_17);
nor U11050 (N_11050,N_2386,N_2506);
nand U11051 (N_11051,N_2052,N_2183);
nor U11052 (N_11052,N_1776,N_1846);
nand U11053 (N_11053,N_3276,N_1794);
or U11054 (N_11054,N_2997,N_333);
or U11055 (N_11055,N_3400,N_3959);
nor U11056 (N_11056,N_4993,N_3010);
nor U11057 (N_11057,N_4960,N_3268);
and U11058 (N_11058,N_2670,N_1730);
or U11059 (N_11059,N_337,N_5337);
xnor U11060 (N_11060,N_1698,N_4515);
and U11061 (N_11061,N_3703,N_5131);
and U11062 (N_11062,N_4589,N_6098);
and U11063 (N_11063,N_1682,N_797);
and U11064 (N_11064,N_3568,N_592);
nor U11065 (N_11065,N_1410,N_4293);
nor U11066 (N_11066,N_3011,N_3504);
or U11067 (N_11067,N_2555,N_6175);
and U11068 (N_11068,N_3489,N_3440);
nor U11069 (N_11069,N_5911,N_3130);
and U11070 (N_11070,N_3859,N_4327);
or U11071 (N_11071,N_2986,N_3786);
and U11072 (N_11072,N_3230,N_591);
nand U11073 (N_11073,N_2491,N_5520);
or U11074 (N_11074,N_2252,N_4948);
nor U11075 (N_11075,N_4850,N_5701);
and U11076 (N_11076,N_1520,N_611);
or U11077 (N_11077,N_768,N_4818);
and U11078 (N_11078,N_654,N_105);
or U11079 (N_11079,N_2972,N_3197);
or U11080 (N_11080,N_129,N_2483);
nand U11081 (N_11081,N_4993,N_3383);
nand U11082 (N_11082,N_3993,N_4172);
nor U11083 (N_11083,N_3766,N_4703);
or U11084 (N_11084,N_5783,N_3244);
and U11085 (N_11085,N_5622,N_4985);
or U11086 (N_11086,N_5756,N_3435);
or U11087 (N_11087,N_2804,N_4226);
and U11088 (N_11088,N_5162,N_4550);
nand U11089 (N_11089,N_1573,N_768);
nand U11090 (N_11090,N_3318,N_370);
nor U11091 (N_11091,N_3544,N_4983);
nand U11092 (N_11092,N_1204,N_1833);
nor U11093 (N_11093,N_3458,N_2134);
and U11094 (N_11094,N_3666,N_5079);
or U11095 (N_11095,N_1180,N_318);
and U11096 (N_11096,N_1608,N_5890);
and U11097 (N_11097,N_5860,N_3499);
and U11098 (N_11098,N_5810,N_6212);
nor U11099 (N_11099,N_4848,N_5433);
and U11100 (N_11100,N_3379,N_2801);
and U11101 (N_11101,N_2185,N_244);
nor U11102 (N_11102,N_493,N_650);
nand U11103 (N_11103,N_1911,N_2497);
or U11104 (N_11104,N_4506,N_3083);
xor U11105 (N_11105,N_3786,N_5101);
or U11106 (N_11106,N_3571,N_3152);
nor U11107 (N_11107,N_2967,N_1494);
and U11108 (N_11108,N_4702,N_3579);
nand U11109 (N_11109,N_3761,N_2872);
nor U11110 (N_11110,N_6054,N_2720);
nand U11111 (N_11111,N_3356,N_4702);
nand U11112 (N_11112,N_989,N_3615);
nor U11113 (N_11113,N_2443,N_2592);
nor U11114 (N_11114,N_2929,N_4993);
nand U11115 (N_11115,N_3699,N_4341);
or U11116 (N_11116,N_674,N_3500);
or U11117 (N_11117,N_6154,N_5765);
and U11118 (N_11118,N_1772,N_6169);
nand U11119 (N_11119,N_486,N_1565);
nor U11120 (N_11120,N_3274,N_759);
nor U11121 (N_11121,N_5389,N_5824);
nand U11122 (N_11122,N_6089,N_418);
nor U11123 (N_11123,N_3188,N_5869);
nor U11124 (N_11124,N_1921,N_3490);
or U11125 (N_11125,N_4837,N_2332);
nand U11126 (N_11126,N_2574,N_5242);
nand U11127 (N_11127,N_885,N_2077);
or U11128 (N_11128,N_3995,N_1797);
and U11129 (N_11129,N_1220,N_4569);
and U11130 (N_11130,N_3927,N_3410);
nor U11131 (N_11131,N_3238,N_10);
nand U11132 (N_11132,N_934,N_2425);
or U11133 (N_11133,N_195,N_3270);
nor U11134 (N_11134,N_2180,N_4951);
nor U11135 (N_11135,N_1068,N_3427);
and U11136 (N_11136,N_2972,N_1651);
nand U11137 (N_11137,N_5561,N_5050);
and U11138 (N_11138,N_3070,N_5443);
or U11139 (N_11139,N_4407,N_1370);
nor U11140 (N_11140,N_2080,N_4972);
nand U11141 (N_11141,N_5758,N_3609);
nor U11142 (N_11142,N_3377,N_5313);
nand U11143 (N_11143,N_4421,N_374);
nor U11144 (N_11144,N_696,N_1226);
and U11145 (N_11145,N_1036,N_4438);
or U11146 (N_11146,N_6064,N_82);
or U11147 (N_11147,N_5165,N_2896);
nor U11148 (N_11148,N_5707,N_976);
or U11149 (N_11149,N_2250,N_5265);
nor U11150 (N_11150,N_4270,N_1811);
and U11151 (N_11151,N_4038,N_5725);
and U11152 (N_11152,N_129,N_181);
or U11153 (N_11153,N_551,N_1179);
nand U11154 (N_11154,N_5908,N_1754);
or U11155 (N_11155,N_2461,N_2954);
nor U11156 (N_11156,N_3130,N_864);
nor U11157 (N_11157,N_5366,N_4999);
nand U11158 (N_11158,N_4725,N_5400);
or U11159 (N_11159,N_2483,N_5792);
or U11160 (N_11160,N_5464,N_3213);
or U11161 (N_11161,N_2136,N_5108);
nor U11162 (N_11162,N_5032,N_5261);
nand U11163 (N_11163,N_4814,N_5574);
nor U11164 (N_11164,N_4434,N_2411);
nand U11165 (N_11165,N_1537,N_592);
nor U11166 (N_11166,N_4101,N_637);
or U11167 (N_11167,N_5476,N_270);
and U11168 (N_11168,N_2304,N_5183);
nand U11169 (N_11169,N_330,N_4136);
nor U11170 (N_11170,N_4733,N_5199);
nor U11171 (N_11171,N_4260,N_2678);
nor U11172 (N_11172,N_1817,N_45);
or U11173 (N_11173,N_3972,N_1027);
and U11174 (N_11174,N_140,N_61);
or U11175 (N_11175,N_5818,N_1506);
and U11176 (N_11176,N_5040,N_4493);
and U11177 (N_11177,N_2230,N_5943);
nand U11178 (N_11178,N_2469,N_5858);
nand U11179 (N_11179,N_5730,N_1302);
nand U11180 (N_11180,N_253,N_2206);
nand U11181 (N_11181,N_1470,N_1540);
or U11182 (N_11182,N_5374,N_862);
nor U11183 (N_11183,N_4475,N_3172);
and U11184 (N_11184,N_3922,N_608);
nor U11185 (N_11185,N_3496,N_137);
nor U11186 (N_11186,N_5565,N_3056);
nor U11187 (N_11187,N_1707,N_3292);
nor U11188 (N_11188,N_4490,N_965);
nor U11189 (N_11189,N_1935,N_2267);
and U11190 (N_11190,N_2128,N_4400);
and U11191 (N_11191,N_552,N_6000);
and U11192 (N_11192,N_2108,N_538);
and U11193 (N_11193,N_4202,N_4756);
or U11194 (N_11194,N_3359,N_3591);
or U11195 (N_11195,N_2124,N_2380);
nand U11196 (N_11196,N_6119,N_4553);
nor U11197 (N_11197,N_5492,N_144);
nor U11198 (N_11198,N_5399,N_5345);
nand U11199 (N_11199,N_4595,N_2274);
nand U11200 (N_11200,N_6192,N_2643);
and U11201 (N_11201,N_1732,N_2835);
or U11202 (N_11202,N_4207,N_5784);
and U11203 (N_11203,N_2176,N_909);
or U11204 (N_11204,N_4794,N_2285);
or U11205 (N_11205,N_3193,N_1794);
or U11206 (N_11206,N_5816,N_5299);
and U11207 (N_11207,N_5183,N_4148);
and U11208 (N_11208,N_4811,N_3029);
and U11209 (N_11209,N_5136,N_2577);
nor U11210 (N_11210,N_5763,N_1052);
nor U11211 (N_11211,N_2885,N_5426);
and U11212 (N_11212,N_2275,N_3995);
nor U11213 (N_11213,N_1890,N_777);
or U11214 (N_11214,N_4518,N_5256);
or U11215 (N_11215,N_516,N_802);
and U11216 (N_11216,N_1602,N_2182);
and U11217 (N_11217,N_1418,N_752);
and U11218 (N_11218,N_1763,N_4816);
or U11219 (N_11219,N_3634,N_3157);
nor U11220 (N_11220,N_175,N_1153);
nand U11221 (N_11221,N_2588,N_273);
and U11222 (N_11222,N_2730,N_103);
nor U11223 (N_11223,N_806,N_1463);
nor U11224 (N_11224,N_2958,N_5733);
or U11225 (N_11225,N_5953,N_3685);
nor U11226 (N_11226,N_3946,N_1498);
nand U11227 (N_11227,N_532,N_1840);
nand U11228 (N_11228,N_2294,N_669);
nor U11229 (N_11229,N_958,N_4540);
or U11230 (N_11230,N_1876,N_15);
and U11231 (N_11231,N_509,N_966);
nor U11232 (N_11232,N_2935,N_5458);
or U11233 (N_11233,N_222,N_3987);
xnor U11234 (N_11234,N_5034,N_2063);
nand U11235 (N_11235,N_3873,N_5565);
nor U11236 (N_11236,N_3467,N_1291);
nor U11237 (N_11237,N_4768,N_4188);
and U11238 (N_11238,N_3501,N_2763);
and U11239 (N_11239,N_131,N_4076);
nand U11240 (N_11240,N_1068,N_5111);
nand U11241 (N_11241,N_281,N_5049);
and U11242 (N_11242,N_2322,N_1518);
and U11243 (N_11243,N_1327,N_784);
and U11244 (N_11244,N_2322,N_2411);
or U11245 (N_11245,N_123,N_2614);
nor U11246 (N_11246,N_4322,N_4806);
nand U11247 (N_11247,N_3590,N_3860);
nand U11248 (N_11248,N_4387,N_591);
and U11249 (N_11249,N_357,N_2902);
or U11250 (N_11250,N_3050,N_46);
nand U11251 (N_11251,N_471,N_6162);
and U11252 (N_11252,N_1707,N_2555);
nor U11253 (N_11253,N_3498,N_5969);
nand U11254 (N_11254,N_540,N_2835);
and U11255 (N_11255,N_1551,N_2887);
nand U11256 (N_11256,N_2607,N_5368);
and U11257 (N_11257,N_5456,N_5040);
or U11258 (N_11258,N_2924,N_1775);
nand U11259 (N_11259,N_5228,N_1193);
or U11260 (N_11260,N_3138,N_5133);
nor U11261 (N_11261,N_5170,N_4843);
and U11262 (N_11262,N_6073,N_2856);
nand U11263 (N_11263,N_90,N_5471);
nand U11264 (N_11264,N_5658,N_3816);
and U11265 (N_11265,N_2111,N_3969);
or U11266 (N_11266,N_610,N_5919);
or U11267 (N_11267,N_2299,N_4282);
and U11268 (N_11268,N_2355,N_2194);
or U11269 (N_11269,N_684,N_2170);
or U11270 (N_11270,N_2702,N_5041);
nor U11271 (N_11271,N_1284,N_4784);
or U11272 (N_11272,N_4681,N_1868);
nand U11273 (N_11273,N_5601,N_2886);
and U11274 (N_11274,N_6058,N_1934);
nand U11275 (N_11275,N_5640,N_6231);
nand U11276 (N_11276,N_3853,N_2930);
and U11277 (N_11277,N_756,N_5517);
or U11278 (N_11278,N_45,N_100);
nor U11279 (N_11279,N_5401,N_2039);
nand U11280 (N_11280,N_3127,N_2537);
nor U11281 (N_11281,N_391,N_4599);
nor U11282 (N_11282,N_3415,N_1129);
nand U11283 (N_11283,N_982,N_349);
nand U11284 (N_11284,N_1242,N_3767);
and U11285 (N_11285,N_935,N_2607);
nand U11286 (N_11286,N_2268,N_2656);
nor U11287 (N_11287,N_6018,N_2286);
nor U11288 (N_11288,N_3690,N_1704);
and U11289 (N_11289,N_3918,N_4144);
and U11290 (N_11290,N_6239,N_3360);
or U11291 (N_11291,N_4701,N_2863);
or U11292 (N_11292,N_4312,N_2685);
and U11293 (N_11293,N_3339,N_3419);
nand U11294 (N_11294,N_1366,N_2498);
nand U11295 (N_11295,N_2124,N_3668);
or U11296 (N_11296,N_5079,N_2359);
nand U11297 (N_11297,N_335,N_5794);
and U11298 (N_11298,N_1255,N_5240);
nor U11299 (N_11299,N_1330,N_255);
nand U11300 (N_11300,N_3897,N_1852);
or U11301 (N_11301,N_569,N_2810);
nor U11302 (N_11302,N_1105,N_5313);
xnor U11303 (N_11303,N_281,N_1490);
nand U11304 (N_11304,N_2455,N_1977);
nor U11305 (N_11305,N_1981,N_5505);
and U11306 (N_11306,N_1875,N_860);
nor U11307 (N_11307,N_3671,N_6039);
and U11308 (N_11308,N_3071,N_2738);
nor U11309 (N_11309,N_2719,N_1128);
nor U11310 (N_11310,N_3410,N_3468);
and U11311 (N_11311,N_6181,N_291);
nor U11312 (N_11312,N_1175,N_4170);
and U11313 (N_11313,N_2458,N_419);
nor U11314 (N_11314,N_2386,N_767);
nand U11315 (N_11315,N_1779,N_4376);
and U11316 (N_11316,N_4268,N_6101);
nand U11317 (N_11317,N_3238,N_2298);
nand U11318 (N_11318,N_512,N_2000);
nor U11319 (N_11319,N_814,N_434);
and U11320 (N_11320,N_2868,N_3422);
nand U11321 (N_11321,N_2381,N_5264);
and U11322 (N_11322,N_4436,N_6234);
nor U11323 (N_11323,N_3302,N_877);
nand U11324 (N_11324,N_1950,N_122);
and U11325 (N_11325,N_3767,N_3948);
and U11326 (N_11326,N_414,N_2331);
nor U11327 (N_11327,N_3896,N_3735);
or U11328 (N_11328,N_153,N_1539);
nor U11329 (N_11329,N_1491,N_4690);
and U11330 (N_11330,N_3162,N_5241);
and U11331 (N_11331,N_2488,N_4440);
and U11332 (N_11332,N_1395,N_4341);
nand U11333 (N_11333,N_1836,N_4369);
nor U11334 (N_11334,N_2092,N_1850);
or U11335 (N_11335,N_4208,N_2955);
nand U11336 (N_11336,N_3883,N_4372);
or U11337 (N_11337,N_4223,N_2923);
or U11338 (N_11338,N_2115,N_5074);
nand U11339 (N_11339,N_840,N_4672);
and U11340 (N_11340,N_2652,N_3218);
or U11341 (N_11341,N_4375,N_1246);
nor U11342 (N_11342,N_4243,N_873);
or U11343 (N_11343,N_3227,N_1034);
nor U11344 (N_11344,N_6188,N_1310);
nor U11345 (N_11345,N_3218,N_3871);
and U11346 (N_11346,N_4644,N_6026);
or U11347 (N_11347,N_48,N_492);
nor U11348 (N_11348,N_2012,N_4099);
and U11349 (N_11349,N_5984,N_3148);
nand U11350 (N_11350,N_5458,N_1724);
and U11351 (N_11351,N_4408,N_2996);
nor U11352 (N_11352,N_4030,N_1907);
nand U11353 (N_11353,N_2394,N_5677);
nand U11354 (N_11354,N_5359,N_3580);
nand U11355 (N_11355,N_5084,N_827);
and U11356 (N_11356,N_3217,N_2739);
nor U11357 (N_11357,N_635,N_2037);
nor U11358 (N_11358,N_3167,N_6064);
nor U11359 (N_11359,N_395,N_1126);
and U11360 (N_11360,N_2611,N_4991);
and U11361 (N_11361,N_554,N_5288);
nand U11362 (N_11362,N_4495,N_660);
and U11363 (N_11363,N_3874,N_6111);
and U11364 (N_11364,N_4441,N_1435);
and U11365 (N_11365,N_1600,N_1700);
or U11366 (N_11366,N_132,N_1297);
and U11367 (N_11367,N_15,N_2908);
nand U11368 (N_11368,N_4079,N_1181);
nand U11369 (N_11369,N_1365,N_4340);
nor U11370 (N_11370,N_3990,N_6192);
or U11371 (N_11371,N_2414,N_646);
xnor U11372 (N_11372,N_3375,N_2790);
or U11373 (N_11373,N_5475,N_6032);
nand U11374 (N_11374,N_2098,N_49);
nor U11375 (N_11375,N_1856,N_5698);
or U11376 (N_11376,N_5713,N_1574);
and U11377 (N_11377,N_6131,N_5792);
and U11378 (N_11378,N_4346,N_5655);
nand U11379 (N_11379,N_264,N_3541);
nand U11380 (N_11380,N_784,N_3237);
nand U11381 (N_11381,N_1010,N_4457);
nand U11382 (N_11382,N_3296,N_507);
nand U11383 (N_11383,N_4079,N_2647);
nand U11384 (N_11384,N_5369,N_4949);
nand U11385 (N_11385,N_5549,N_623);
or U11386 (N_11386,N_1687,N_2244);
and U11387 (N_11387,N_2793,N_3244);
nor U11388 (N_11388,N_1537,N_1706);
or U11389 (N_11389,N_4906,N_3356);
or U11390 (N_11390,N_5145,N_5832);
and U11391 (N_11391,N_2041,N_5868);
nor U11392 (N_11392,N_4354,N_5210);
nor U11393 (N_11393,N_5960,N_4709);
nor U11394 (N_11394,N_5709,N_5852);
or U11395 (N_11395,N_3599,N_4081);
and U11396 (N_11396,N_3414,N_1918);
nand U11397 (N_11397,N_972,N_2304);
or U11398 (N_11398,N_6221,N_13);
or U11399 (N_11399,N_5969,N_4420);
nand U11400 (N_11400,N_1816,N_3242);
or U11401 (N_11401,N_4726,N_2601);
nor U11402 (N_11402,N_274,N_3247);
and U11403 (N_11403,N_717,N_492);
nor U11404 (N_11404,N_460,N_4792);
nand U11405 (N_11405,N_3099,N_6135);
and U11406 (N_11406,N_3098,N_6043);
or U11407 (N_11407,N_2060,N_4759);
and U11408 (N_11408,N_1900,N_520);
nand U11409 (N_11409,N_2250,N_2256);
nor U11410 (N_11410,N_164,N_1189);
and U11411 (N_11411,N_3968,N_4022);
and U11412 (N_11412,N_872,N_3755);
or U11413 (N_11413,N_1119,N_3588);
and U11414 (N_11414,N_177,N_1195);
nand U11415 (N_11415,N_1980,N_2780);
nor U11416 (N_11416,N_655,N_451);
or U11417 (N_11417,N_632,N_3396);
nor U11418 (N_11418,N_3835,N_5944);
and U11419 (N_11419,N_218,N_1328);
or U11420 (N_11420,N_5124,N_5962);
nor U11421 (N_11421,N_5251,N_4764);
nor U11422 (N_11422,N_832,N_115);
and U11423 (N_11423,N_4611,N_2449);
or U11424 (N_11424,N_755,N_2457);
and U11425 (N_11425,N_6048,N_1870);
or U11426 (N_11426,N_2091,N_4913);
nand U11427 (N_11427,N_2450,N_463);
nand U11428 (N_11428,N_2892,N_4471);
or U11429 (N_11429,N_3421,N_5655);
nor U11430 (N_11430,N_2374,N_646);
or U11431 (N_11431,N_3210,N_5617);
nand U11432 (N_11432,N_5420,N_2111);
nor U11433 (N_11433,N_5898,N_3880);
or U11434 (N_11434,N_2850,N_3890);
and U11435 (N_11435,N_3636,N_899);
or U11436 (N_11436,N_285,N_413);
and U11437 (N_11437,N_5417,N_1919);
nand U11438 (N_11438,N_1057,N_5924);
nand U11439 (N_11439,N_1899,N_828);
nor U11440 (N_11440,N_1280,N_1404);
and U11441 (N_11441,N_3937,N_3082);
and U11442 (N_11442,N_241,N_2359);
and U11443 (N_11443,N_4764,N_2453);
nor U11444 (N_11444,N_4280,N_750);
nor U11445 (N_11445,N_2843,N_6054);
and U11446 (N_11446,N_4926,N_2769);
nor U11447 (N_11447,N_2462,N_4425);
or U11448 (N_11448,N_1710,N_2243);
and U11449 (N_11449,N_2184,N_5005);
or U11450 (N_11450,N_1013,N_3302);
and U11451 (N_11451,N_1871,N_5119);
and U11452 (N_11452,N_1152,N_442);
nor U11453 (N_11453,N_2905,N_2904);
nor U11454 (N_11454,N_254,N_2478);
nor U11455 (N_11455,N_5016,N_3620);
nor U11456 (N_11456,N_4795,N_2040);
and U11457 (N_11457,N_947,N_5897);
nor U11458 (N_11458,N_1013,N_29);
and U11459 (N_11459,N_4254,N_2404);
nor U11460 (N_11460,N_2153,N_3507);
and U11461 (N_11461,N_5212,N_3308);
nor U11462 (N_11462,N_3625,N_1548);
or U11463 (N_11463,N_689,N_1730);
or U11464 (N_11464,N_2445,N_4828);
nand U11465 (N_11465,N_4142,N_240);
nor U11466 (N_11466,N_2337,N_5871);
nand U11467 (N_11467,N_6028,N_4249);
or U11468 (N_11468,N_351,N_2689);
and U11469 (N_11469,N_1282,N_3574);
or U11470 (N_11470,N_63,N_583);
nor U11471 (N_11471,N_5219,N_4313);
nand U11472 (N_11472,N_4184,N_4258);
and U11473 (N_11473,N_5,N_1252);
and U11474 (N_11474,N_495,N_3520);
or U11475 (N_11475,N_5575,N_6009);
or U11476 (N_11476,N_4011,N_4777);
nand U11477 (N_11477,N_5804,N_4714);
and U11478 (N_11478,N_3797,N_1638);
or U11479 (N_11479,N_3152,N_1628);
nor U11480 (N_11480,N_5656,N_4220);
nand U11481 (N_11481,N_761,N_5155);
nor U11482 (N_11482,N_6228,N_2839);
or U11483 (N_11483,N_3270,N_1211);
nand U11484 (N_11484,N_992,N_4205);
nor U11485 (N_11485,N_5537,N_2062);
nand U11486 (N_11486,N_5852,N_3160);
nand U11487 (N_11487,N_2724,N_1179);
nand U11488 (N_11488,N_3941,N_3182);
and U11489 (N_11489,N_2100,N_4594);
nand U11490 (N_11490,N_2424,N_2533);
and U11491 (N_11491,N_6087,N_2515);
or U11492 (N_11492,N_5567,N_3963);
nor U11493 (N_11493,N_399,N_1123);
or U11494 (N_11494,N_4671,N_2491);
nor U11495 (N_11495,N_4129,N_1502);
or U11496 (N_11496,N_553,N_4082);
or U11497 (N_11497,N_3369,N_405);
or U11498 (N_11498,N_1469,N_2862);
nor U11499 (N_11499,N_432,N_1479);
nand U11500 (N_11500,N_1228,N_2340);
and U11501 (N_11501,N_6139,N_5512);
nand U11502 (N_11502,N_3348,N_903);
and U11503 (N_11503,N_5017,N_5371);
or U11504 (N_11504,N_2985,N_1436);
nor U11505 (N_11505,N_1580,N_6159);
nand U11506 (N_11506,N_4109,N_4890);
nor U11507 (N_11507,N_2818,N_5089);
nor U11508 (N_11508,N_1347,N_5542);
nor U11509 (N_11509,N_666,N_2124);
and U11510 (N_11510,N_903,N_1636);
or U11511 (N_11511,N_3751,N_4108);
or U11512 (N_11512,N_3181,N_2926);
nand U11513 (N_11513,N_2476,N_3629);
or U11514 (N_11514,N_5460,N_75);
nor U11515 (N_11515,N_1351,N_3641);
or U11516 (N_11516,N_3358,N_47);
and U11517 (N_11517,N_4788,N_3078);
or U11518 (N_11518,N_5628,N_5453);
or U11519 (N_11519,N_3342,N_1592);
nor U11520 (N_11520,N_451,N_3886);
or U11521 (N_11521,N_1224,N_1150);
nor U11522 (N_11522,N_997,N_4169);
and U11523 (N_11523,N_1707,N_819);
nor U11524 (N_11524,N_4870,N_1298);
nor U11525 (N_11525,N_1673,N_4002);
or U11526 (N_11526,N_76,N_3192);
nor U11527 (N_11527,N_46,N_2166);
nor U11528 (N_11528,N_1735,N_1533);
nand U11529 (N_11529,N_928,N_2737);
xor U11530 (N_11530,N_5586,N_4191);
and U11531 (N_11531,N_4046,N_2727);
or U11532 (N_11532,N_5686,N_2582);
or U11533 (N_11533,N_3508,N_1480);
or U11534 (N_11534,N_1789,N_1033);
and U11535 (N_11535,N_199,N_3795);
and U11536 (N_11536,N_1362,N_5178);
and U11537 (N_11537,N_4470,N_5953);
or U11538 (N_11538,N_3793,N_3193);
or U11539 (N_11539,N_2000,N_5105);
nand U11540 (N_11540,N_1126,N_1995);
or U11541 (N_11541,N_3308,N_3367);
and U11542 (N_11542,N_1470,N_66);
and U11543 (N_11543,N_1886,N_2883);
nand U11544 (N_11544,N_3832,N_1314);
or U11545 (N_11545,N_3635,N_1884);
or U11546 (N_11546,N_4319,N_4845);
or U11547 (N_11547,N_1423,N_4361);
nand U11548 (N_11548,N_5420,N_75);
nor U11549 (N_11549,N_2384,N_1316);
and U11550 (N_11550,N_1401,N_265);
and U11551 (N_11551,N_3545,N_2295);
or U11552 (N_11552,N_965,N_4227);
nand U11553 (N_11553,N_3029,N_5898);
or U11554 (N_11554,N_3441,N_149);
nor U11555 (N_11555,N_2872,N_3286);
and U11556 (N_11556,N_2576,N_2974);
and U11557 (N_11557,N_525,N_2335);
and U11558 (N_11558,N_2584,N_3222);
or U11559 (N_11559,N_6140,N_5650);
nor U11560 (N_11560,N_6229,N_3751);
nor U11561 (N_11561,N_4892,N_390);
or U11562 (N_11562,N_1567,N_325);
or U11563 (N_11563,N_3311,N_960);
nand U11564 (N_11564,N_1776,N_81);
nand U11565 (N_11565,N_2603,N_6230);
nand U11566 (N_11566,N_1122,N_2978);
or U11567 (N_11567,N_1673,N_867);
or U11568 (N_11568,N_6210,N_3084);
xor U11569 (N_11569,N_5455,N_5709);
nand U11570 (N_11570,N_2052,N_5905);
nand U11571 (N_11571,N_5751,N_4363);
nand U11572 (N_11572,N_3154,N_638);
nand U11573 (N_11573,N_2865,N_3327);
or U11574 (N_11574,N_4635,N_3199);
or U11575 (N_11575,N_798,N_2474);
nor U11576 (N_11576,N_288,N_701);
or U11577 (N_11577,N_1853,N_6034);
or U11578 (N_11578,N_5605,N_2173);
nand U11579 (N_11579,N_654,N_2062);
and U11580 (N_11580,N_4834,N_3919);
nand U11581 (N_11581,N_2068,N_3429);
nand U11582 (N_11582,N_1570,N_5435);
and U11583 (N_11583,N_3161,N_3432);
nand U11584 (N_11584,N_3155,N_1423);
and U11585 (N_11585,N_5034,N_1158);
nor U11586 (N_11586,N_1669,N_3511);
nand U11587 (N_11587,N_78,N_5911);
or U11588 (N_11588,N_2632,N_2437);
nand U11589 (N_11589,N_3003,N_634);
or U11590 (N_11590,N_5453,N_3740);
nor U11591 (N_11591,N_1066,N_120);
nand U11592 (N_11592,N_4242,N_3942);
nor U11593 (N_11593,N_5022,N_5130);
or U11594 (N_11594,N_2594,N_1911);
and U11595 (N_11595,N_4472,N_5987);
nand U11596 (N_11596,N_1278,N_3038);
nor U11597 (N_11597,N_2115,N_142);
and U11598 (N_11598,N_3965,N_3577);
nor U11599 (N_11599,N_745,N_3635);
and U11600 (N_11600,N_4707,N_1598);
or U11601 (N_11601,N_3848,N_4440);
nand U11602 (N_11602,N_3833,N_6117);
nand U11603 (N_11603,N_932,N_5049);
nand U11604 (N_11604,N_2725,N_1358);
nor U11605 (N_11605,N_1597,N_5038);
and U11606 (N_11606,N_5575,N_1019);
nor U11607 (N_11607,N_726,N_5757);
nor U11608 (N_11608,N_2228,N_2154);
nor U11609 (N_11609,N_4687,N_4111);
or U11610 (N_11610,N_1702,N_3095);
and U11611 (N_11611,N_3074,N_5910);
and U11612 (N_11612,N_4680,N_3736);
or U11613 (N_11613,N_224,N_3505);
nor U11614 (N_11614,N_2506,N_383);
nor U11615 (N_11615,N_1677,N_3125);
nand U11616 (N_11616,N_346,N_1526);
and U11617 (N_11617,N_3556,N_346);
nand U11618 (N_11618,N_5861,N_256);
or U11619 (N_11619,N_4090,N_4623);
and U11620 (N_11620,N_3361,N_1603);
and U11621 (N_11621,N_4031,N_4772);
or U11622 (N_11622,N_3472,N_5595);
nor U11623 (N_11623,N_888,N_4215);
nor U11624 (N_11624,N_4548,N_5718);
nand U11625 (N_11625,N_6004,N_2675);
nor U11626 (N_11626,N_391,N_116);
and U11627 (N_11627,N_4538,N_4022);
nand U11628 (N_11628,N_5412,N_3139);
nor U11629 (N_11629,N_1239,N_2376);
nand U11630 (N_11630,N_2040,N_926);
nand U11631 (N_11631,N_178,N_3892);
and U11632 (N_11632,N_3851,N_5593);
nor U11633 (N_11633,N_1985,N_1380);
nand U11634 (N_11634,N_3788,N_6157);
nor U11635 (N_11635,N_5982,N_3023);
and U11636 (N_11636,N_3157,N_1674);
nand U11637 (N_11637,N_4318,N_677);
nand U11638 (N_11638,N_1867,N_5591);
or U11639 (N_11639,N_5858,N_584);
and U11640 (N_11640,N_5436,N_3133);
or U11641 (N_11641,N_5131,N_2400);
nand U11642 (N_11642,N_2513,N_4593);
nor U11643 (N_11643,N_4638,N_2897);
and U11644 (N_11644,N_4194,N_3628);
or U11645 (N_11645,N_2939,N_64);
nor U11646 (N_11646,N_260,N_4081);
and U11647 (N_11647,N_5047,N_4114);
or U11648 (N_11648,N_2662,N_4924);
nor U11649 (N_11649,N_3679,N_2592);
nor U11650 (N_11650,N_4132,N_4209);
nor U11651 (N_11651,N_228,N_2832);
and U11652 (N_11652,N_1558,N_3690);
and U11653 (N_11653,N_5623,N_3650);
nor U11654 (N_11654,N_3455,N_5876);
nand U11655 (N_11655,N_200,N_875);
nand U11656 (N_11656,N_1203,N_4378);
and U11657 (N_11657,N_4165,N_1207);
or U11658 (N_11658,N_2275,N_3247);
nor U11659 (N_11659,N_447,N_1566);
or U11660 (N_11660,N_1129,N_1528);
nor U11661 (N_11661,N_5833,N_6089);
nand U11662 (N_11662,N_241,N_5290);
and U11663 (N_11663,N_4956,N_1140);
nand U11664 (N_11664,N_3108,N_2506);
nand U11665 (N_11665,N_1624,N_565);
nor U11666 (N_11666,N_4311,N_4183);
or U11667 (N_11667,N_918,N_5032);
or U11668 (N_11668,N_122,N_206);
or U11669 (N_11669,N_3880,N_3316);
and U11670 (N_11670,N_5623,N_1913);
or U11671 (N_11671,N_6103,N_5084);
nand U11672 (N_11672,N_4261,N_5236);
nor U11673 (N_11673,N_2715,N_5391);
nand U11674 (N_11674,N_361,N_5726);
and U11675 (N_11675,N_4696,N_885);
or U11676 (N_11676,N_4006,N_4032);
or U11677 (N_11677,N_4270,N_2903);
or U11678 (N_11678,N_1396,N_4019);
or U11679 (N_11679,N_1380,N_3981);
or U11680 (N_11680,N_3320,N_3791);
and U11681 (N_11681,N_5247,N_4851);
nor U11682 (N_11682,N_20,N_4529);
or U11683 (N_11683,N_152,N_2179);
nand U11684 (N_11684,N_3037,N_2095);
or U11685 (N_11685,N_5158,N_6065);
or U11686 (N_11686,N_1354,N_4762);
nand U11687 (N_11687,N_2478,N_3945);
or U11688 (N_11688,N_1681,N_4198);
nand U11689 (N_11689,N_895,N_1803);
nand U11690 (N_11690,N_5549,N_5857);
nor U11691 (N_11691,N_2159,N_5594);
nand U11692 (N_11692,N_1112,N_2654);
or U11693 (N_11693,N_2820,N_2876);
or U11694 (N_11694,N_5158,N_4352);
nand U11695 (N_11695,N_277,N_4753);
nor U11696 (N_11696,N_51,N_5556);
nand U11697 (N_11697,N_1009,N_6006);
nor U11698 (N_11698,N_297,N_2507);
or U11699 (N_11699,N_2279,N_2903);
nand U11700 (N_11700,N_4480,N_3083);
nand U11701 (N_11701,N_5819,N_4025);
nand U11702 (N_11702,N_3559,N_1553);
nand U11703 (N_11703,N_3576,N_5446);
and U11704 (N_11704,N_2826,N_3991);
nand U11705 (N_11705,N_4445,N_2420);
or U11706 (N_11706,N_1063,N_803);
or U11707 (N_11707,N_2773,N_4288);
and U11708 (N_11708,N_2553,N_3541);
and U11709 (N_11709,N_687,N_5284);
and U11710 (N_11710,N_5952,N_3068);
and U11711 (N_11711,N_5026,N_6068);
nor U11712 (N_11712,N_6081,N_3010);
and U11713 (N_11713,N_1411,N_2307);
nor U11714 (N_11714,N_3452,N_3463);
or U11715 (N_11715,N_4601,N_1681);
and U11716 (N_11716,N_4844,N_2853);
or U11717 (N_11717,N_6065,N_5487);
or U11718 (N_11718,N_1941,N_985);
nor U11719 (N_11719,N_5781,N_4838);
and U11720 (N_11720,N_5823,N_1659);
and U11721 (N_11721,N_1275,N_414);
or U11722 (N_11722,N_457,N_4135);
nor U11723 (N_11723,N_6062,N_1202);
nor U11724 (N_11724,N_2019,N_821);
and U11725 (N_11725,N_5048,N_1614);
nand U11726 (N_11726,N_3233,N_6020);
nor U11727 (N_11727,N_1429,N_931);
nand U11728 (N_11728,N_2632,N_2917);
nand U11729 (N_11729,N_4071,N_5646);
or U11730 (N_11730,N_2079,N_119);
nor U11731 (N_11731,N_5825,N_5931);
nand U11732 (N_11732,N_2478,N_3728);
nor U11733 (N_11733,N_5092,N_6222);
or U11734 (N_11734,N_3481,N_2468);
or U11735 (N_11735,N_1276,N_1137);
or U11736 (N_11736,N_1264,N_3385);
and U11737 (N_11737,N_4744,N_6032);
nand U11738 (N_11738,N_3112,N_5624);
nand U11739 (N_11739,N_4939,N_3575);
and U11740 (N_11740,N_1705,N_3082);
nor U11741 (N_11741,N_1979,N_5);
and U11742 (N_11742,N_3864,N_3771);
and U11743 (N_11743,N_3284,N_902);
nand U11744 (N_11744,N_4157,N_2348);
or U11745 (N_11745,N_3022,N_2203);
nor U11746 (N_11746,N_5921,N_675);
nor U11747 (N_11747,N_1674,N_5854);
or U11748 (N_11748,N_6045,N_5697);
nand U11749 (N_11749,N_1136,N_117);
or U11750 (N_11750,N_6132,N_5634);
nand U11751 (N_11751,N_4187,N_1794);
or U11752 (N_11752,N_1272,N_2176);
nor U11753 (N_11753,N_3355,N_274);
and U11754 (N_11754,N_2290,N_4060);
or U11755 (N_11755,N_4911,N_3562);
nor U11756 (N_11756,N_1409,N_1393);
or U11757 (N_11757,N_2317,N_1021);
nand U11758 (N_11758,N_5121,N_4063);
nor U11759 (N_11759,N_3848,N_5674);
nand U11760 (N_11760,N_2531,N_4483);
nand U11761 (N_11761,N_1395,N_3884);
nand U11762 (N_11762,N_3528,N_1026);
and U11763 (N_11763,N_1664,N_706);
nor U11764 (N_11764,N_422,N_595);
nand U11765 (N_11765,N_2674,N_5322);
nor U11766 (N_11766,N_3923,N_972);
or U11767 (N_11767,N_1021,N_2849);
or U11768 (N_11768,N_5158,N_1532);
and U11769 (N_11769,N_1200,N_1874);
nor U11770 (N_11770,N_1443,N_3225);
or U11771 (N_11771,N_4727,N_1721);
nand U11772 (N_11772,N_3701,N_1757);
nor U11773 (N_11773,N_778,N_250);
and U11774 (N_11774,N_176,N_279);
or U11775 (N_11775,N_157,N_2251);
nand U11776 (N_11776,N_4775,N_4007);
or U11777 (N_11777,N_2604,N_2018);
and U11778 (N_11778,N_223,N_1710);
or U11779 (N_11779,N_395,N_1589);
or U11780 (N_11780,N_1501,N_3497);
nand U11781 (N_11781,N_2163,N_3011);
or U11782 (N_11782,N_5165,N_581);
nand U11783 (N_11783,N_5261,N_791);
nor U11784 (N_11784,N_3079,N_4931);
and U11785 (N_11785,N_4060,N_2456);
or U11786 (N_11786,N_5344,N_4304);
nor U11787 (N_11787,N_423,N_3642);
and U11788 (N_11788,N_6140,N_383);
nand U11789 (N_11789,N_3607,N_2339);
xor U11790 (N_11790,N_5176,N_4844);
and U11791 (N_11791,N_11,N_5295);
xnor U11792 (N_11792,N_114,N_764);
xnor U11793 (N_11793,N_3845,N_3558);
nand U11794 (N_11794,N_1303,N_972);
or U11795 (N_11795,N_4797,N_294);
or U11796 (N_11796,N_3457,N_3917);
nand U11797 (N_11797,N_1707,N_2093);
and U11798 (N_11798,N_6231,N_2325);
nor U11799 (N_11799,N_2952,N_978);
nand U11800 (N_11800,N_1595,N_5412);
nor U11801 (N_11801,N_612,N_2262);
or U11802 (N_11802,N_2295,N_3808);
and U11803 (N_11803,N_3480,N_4145);
and U11804 (N_11804,N_5606,N_1147);
and U11805 (N_11805,N_3492,N_709);
or U11806 (N_11806,N_2679,N_2776);
nor U11807 (N_11807,N_3576,N_4265);
or U11808 (N_11808,N_4248,N_5832);
and U11809 (N_11809,N_3403,N_135);
or U11810 (N_11810,N_3810,N_4435);
nor U11811 (N_11811,N_5611,N_445);
or U11812 (N_11812,N_3294,N_1474);
nor U11813 (N_11813,N_435,N_719);
nand U11814 (N_11814,N_1534,N_4552);
nor U11815 (N_11815,N_558,N_293);
or U11816 (N_11816,N_2063,N_5226);
nor U11817 (N_11817,N_4245,N_3137);
nand U11818 (N_11818,N_5443,N_1127);
or U11819 (N_11819,N_1885,N_2808);
or U11820 (N_11820,N_2825,N_1696);
nor U11821 (N_11821,N_1801,N_826);
nand U11822 (N_11822,N_3589,N_208);
nand U11823 (N_11823,N_3019,N_6126);
nand U11824 (N_11824,N_6191,N_578);
nand U11825 (N_11825,N_2744,N_4189);
or U11826 (N_11826,N_5456,N_465);
or U11827 (N_11827,N_5768,N_1323);
and U11828 (N_11828,N_1939,N_962);
nand U11829 (N_11829,N_5723,N_2552);
nand U11830 (N_11830,N_547,N_336);
nand U11831 (N_11831,N_5933,N_954);
nor U11832 (N_11832,N_5296,N_2187);
and U11833 (N_11833,N_536,N_6215);
or U11834 (N_11834,N_2635,N_3137);
or U11835 (N_11835,N_1755,N_5078);
and U11836 (N_11836,N_3829,N_4115);
nor U11837 (N_11837,N_3249,N_3326);
or U11838 (N_11838,N_264,N_3378);
or U11839 (N_11839,N_2996,N_4783);
xor U11840 (N_11840,N_4500,N_1755);
nand U11841 (N_11841,N_5226,N_4820);
nor U11842 (N_11842,N_3662,N_2418);
nand U11843 (N_11843,N_5476,N_1120);
nor U11844 (N_11844,N_1437,N_3340);
nand U11845 (N_11845,N_368,N_61);
nand U11846 (N_11846,N_2975,N_2711);
or U11847 (N_11847,N_3905,N_4917);
or U11848 (N_11848,N_5781,N_1391);
nand U11849 (N_11849,N_1768,N_987);
nand U11850 (N_11850,N_874,N_99);
or U11851 (N_11851,N_2380,N_4855);
nand U11852 (N_11852,N_595,N_2805);
nor U11853 (N_11853,N_1047,N_2264);
nand U11854 (N_11854,N_4048,N_4292);
nand U11855 (N_11855,N_310,N_2507);
nand U11856 (N_11856,N_1970,N_2885);
or U11857 (N_11857,N_1677,N_2316);
xor U11858 (N_11858,N_4551,N_1390);
or U11859 (N_11859,N_4530,N_5143);
nor U11860 (N_11860,N_3277,N_2774);
nand U11861 (N_11861,N_276,N_2770);
or U11862 (N_11862,N_574,N_5130);
nor U11863 (N_11863,N_5963,N_321);
nor U11864 (N_11864,N_5804,N_3931);
and U11865 (N_11865,N_3758,N_6177);
or U11866 (N_11866,N_3782,N_455);
nand U11867 (N_11867,N_5288,N_5349);
and U11868 (N_11868,N_2295,N_418);
nor U11869 (N_11869,N_5133,N_3632);
and U11870 (N_11870,N_5727,N_1643);
nor U11871 (N_11871,N_4,N_554);
or U11872 (N_11872,N_5481,N_3351);
or U11873 (N_11873,N_5814,N_4075);
or U11874 (N_11874,N_1984,N_2859);
nand U11875 (N_11875,N_305,N_451);
and U11876 (N_11876,N_3191,N_1825);
nand U11877 (N_11877,N_2597,N_4879);
nor U11878 (N_11878,N_2438,N_4698);
nand U11879 (N_11879,N_6051,N_1894);
or U11880 (N_11880,N_1873,N_3413);
or U11881 (N_11881,N_4426,N_1070);
nor U11882 (N_11882,N_2458,N_2074);
nor U11883 (N_11883,N_788,N_3969);
or U11884 (N_11884,N_4804,N_2240);
nand U11885 (N_11885,N_4327,N_5156);
nand U11886 (N_11886,N_1661,N_2886);
and U11887 (N_11887,N_5986,N_1151);
or U11888 (N_11888,N_106,N_2984);
nor U11889 (N_11889,N_5663,N_746);
or U11890 (N_11890,N_3344,N_431);
and U11891 (N_11891,N_596,N_217);
nor U11892 (N_11892,N_5852,N_543);
or U11893 (N_11893,N_6171,N_3621);
nand U11894 (N_11894,N_1592,N_4483);
and U11895 (N_11895,N_4964,N_2862);
and U11896 (N_11896,N_974,N_2266);
and U11897 (N_11897,N_2334,N_5824);
or U11898 (N_11898,N_2384,N_2094);
xnor U11899 (N_11899,N_5253,N_1632);
nor U11900 (N_11900,N_3465,N_1940);
or U11901 (N_11901,N_4257,N_4460);
nor U11902 (N_11902,N_5458,N_2507);
nand U11903 (N_11903,N_1286,N_3912);
nand U11904 (N_11904,N_3156,N_5943);
nor U11905 (N_11905,N_5633,N_4279);
and U11906 (N_11906,N_354,N_1218);
nor U11907 (N_11907,N_2658,N_4660);
nor U11908 (N_11908,N_346,N_2599);
or U11909 (N_11909,N_1396,N_4975);
nand U11910 (N_11910,N_364,N_5495);
nand U11911 (N_11911,N_4087,N_3527);
nor U11912 (N_11912,N_4285,N_4985);
nor U11913 (N_11913,N_5135,N_4615);
nor U11914 (N_11914,N_3049,N_883);
nand U11915 (N_11915,N_3390,N_1730);
nand U11916 (N_11916,N_470,N_3364);
nor U11917 (N_11917,N_2051,N_3672);
nor U11918 (N_11918,N_4608,N_3261);
and U11919 (N_11919,N_3470,N_435);
nor U11920 (N_11920,N_5417,N_198);
xnor U11921 (N_11921,N_3274,N_3373);
or U11922 (N_11922,N_1312,N_1380);
nor U11923 (N_11923,N_1604,N_1939);
and U11924 (N_11924,N_6169,N_2471);
or U11925 (N_11925,N_556,N_1915);
and U11926 (N_11926,N_4575,N_4881);
nand U11927 (N_11927,N_5643,N_4543);
and U11928 (N_11928,N_1693,N_356);
nor U11929 (N_11929,N_1874,N_1350);
and U11930 (N_11930,N_569,N_4694);
nand U11931 (N_11931,N_6075,N_1421);
or U11932 (N_11932,N_5766,N_5937);
nor U11933 (N_11933,N_4489,N_1081);
nand U11934 (N_11934,N_2654,N_5935);
or U11935 (N_11935,N_491,N_2505);
nor U11936 (N_11936,N_6185,N_3953);
or U11937 (N_11937,N_4685,N_2479);
nor U11938 (N_11938,N_1204,N_5344);
nand U11939 (N_11939,N_1306,N_336);
or U11940 (N_11940,N_5988,N_4050);
or U11941 (N_11941,N_1751,N_5052);
nor U11942 (N_11942,N_2123,N_397);
nor U11943 (N_11943,N_5080,N_701);
and U11944 (N_11944,N_238,N_5081);
and U11945 (N_11945,N_3399,N_3838);
nand U11946 (N_11946,N_3219,N_3378);
and U11947 (N_11947,N_2259,N_4777);
nor U11948 (N_11948,N_222,N_4525);
or U11949 (N_11949,N_4041,N_1384);
nand U11950 (N_11950,N_5317,N_1734);
nor U11951 (N_11951,N_642,N_3531);
and U11952 (N_11952,N_1979,N_2362);
nand U11953 (N_11953,N_5144,N_1628);
or U11954 (N_11954,N_992,N_994);
nand U11955 (N_11955,N_6138,N_2885);
nand U11956 (N_11956,N_3966,N_5779);
nor U11957 (N_11957,N_2748,N_1568);
and U11958 (N_11958,N_4335,N_2663);
and U11959 (N_11959,N_5964,N_5418);
and U11960 (N_11960,N_1166,N_1823);
and U11961 (N_11961,N_5247,N_5673);
and U11962 (N_11962,N_3596,N_1580);
or U11963 (N_11963,N_4841,N_4453);
and U11964 (N_11964,N_4901,N_2642);
nor U11965 (N_11965,N_1932,N_3511);
and U11966 (N_11966,N_5269,N_2240);
or U11967 (N_11967,N_970,N_4683);
nand U11968 (N_11968,N_4522,N_4384);
or U11969 (N_11969,N_3065,N_5857);
nor U11970 (N_11970,N_3662,N_2335);
or U11971 (N_11971,N_4281,N_4728);
nor U11972 (N_11972,N_4799,N_5272);
or U11973 (N_11973,N_2933,N_5348);
and U11974 (N_11974,N_5427,N_5737);
nor U11975 (N_11975,N_4316,N_506);
nand U11976 (N_11976,N_145,N_6052);
nor U11977 (N_11977,N_4602,N_6015);
or U11978 (N_11978,N_2822,N_75);
or U11979 (N_11979,N_4975,N_2262);
nand U11980 (N_11980,N_1362,N_4848);
nor U11981 (N_11981,N_1169,N_3083);
or U11982 (N_11982,N_5324,N_1115);
and U11983 (N_11983,N_4319,N_4587);
and U11984 (N_11984,N_2875,N_843);
nor U11985 (N_11985,N_3550,N_1476);
or U11986 (N_11986,N_2054,N_497);
or U11987 (N_11987,N_5672,N_2507);
or U11988 (N_11988,N_3411,N_3731);
nor U11989 (N_11989,N_3670,N_2602);
and U11990 (N_11990,N_3371,N_2024);
nor U11991 (N_11991,N_5970,N_2375);
nand U11992 (N_11992,N_696,N_164);
and U11993 (N_11993,N_3860,N_3232);
nor U11994 (N_11994,N_5273,N_3443);
nor U11995 (N_11995,N_1369,N_2447);
nand U11996 (N_11996,N_2418,N_4506);
or U11997 (N_11997,N_271,N_3422);
nor U11998 (N_11998,N_5544,N_4629);
or U11999 (N_11999,N_4452,N_4626);
nand U12000 (N_12000,N_240,N_1417);
nor U12001 (N_12001,N_4011,N_1314);
nand U12002 (N_12002,N_2156,N_1259);
and U12003 (N_12003,N_508,N_1074);
nor U12004 (N_12004,N_59,N_3886);
and U12005 (N_12005,N_3866,N_822);
or U12006 (N_12006,N_5696,N_1668);
nor U12007 (N_12007,N_2886,N_3972);
or U12008 (N_12008,N_751,N_48);
nor U12009 (N_12009,N_5870,N_4531);
nor U12010 (N_12010,N_5829,N_254);
nor U12011 (N_12011,N_2935,N_795);
nor U12012 (N_12012,N_130,N_4811);
and U12013 (N_12013,N_2766,N_1743);
nor U12014 (N_12014,N_1207,N_4315);
nand U12015 (N_12015,N_1607,N_5456);
nor U12016 (N_12016,N_3057,N_1667);
nand U12017 (N_12017,N_111,N_1198);
nor U12018 (N_12018,N_4739,N_525);
or U12019 (N_12019,N_5133,N_3244);
nor U12020 (N_12020,N_2974,N_4593);
nor U12021 (N_12021,N_4935,N_786);
and U12022 (N_12022,N_1935,N_3604);
or U12023 (N_12023,N_86,N_1643);
nor U12024 (N_12024,N_119,N_1816);
nor U12025 (N_12025,N_2551,N_5938);
nor U12026 (N_12026,N_2183,N_2705);
or U12027 (N_12027,N_4817,N_1422);
xnor U12028 (N_12028,N_3484,N_4038);
and U12029 (N_12029,N_6217,N_4819);
and U12030 (N_12030,N_5930,N_1573);
or U12031 (N_12031,N_5199,N_1731);
and U12032 (N_12032,N_1674,N_5125);
and U12033 (N_12033,N_785,N_5405);
nor U12034 (N_12034,N_4286,N_1234);
or U12035 (N_12035,N_2617,N_5951);
nand U12036 (N_12036,N_5341,N_4000);
nand U12037 (N_12037,N_1130,N_5007);
nor U12038 (N_12038,N_2217,N_5765);
nor U12039 (N_12039,N_3410,N_369);
and U12040 (N_12040,N_4083,N_1947);
and U12041 (N_12041,N_2044,N_989);
nand U12042 (N_12042,N_3898,N_1220);
nor U12043 (N_12043,N_4922,N_2300);
or U12044 (N_12044,N_5720,N_184);
nand U12045 (N_12045,N_3757,N_5130);
nor U12046 (N_12046,N_4712,N_1244);
nand U12047 (N_12047,N_2545,N_3717);
and U12048 (N_12048,N_3940,N_4);
and U12049 (N_12049,N_5903,N_4719);
or U12050 (N_12050,N_884,N_5792);
or U12051 (N_12051,N_4661,N_3610);
nor U12052 (N_12052,N_4979,N_1699);
nand U12053 (N_12053,N_1183,N_1533);
nor U12054 (N_12054,N_4373,N_446);
nor U12055 (N_12055,N_453,N_2918);
and U12056 (N_12056,N_4124,N_6240);
nor U12057 (N_12057,N_3156,N_1037);
nor U12058 (N_12058,N_3485,N_562);
nor U12059 (N_12059,N_3280,N_1952);
nand U12060 (N_12060,N_222,N_4180);
nand U12061 (N_12061,N_3362,N_599);
and U12062 (N_12062,N_4864,N_196);
nand U12063 (N_12063,N_389,N_5724);
nor U12064 (N_12064,N_767,N_3430);
nor U12065 (N_12065,N_2445,N_235);
nor U12066 (N_12066,N_730,N_1933);
or U12067 (N_12067,N_3216,N_132);
nand U12068 (N_12068,N_4,N_4550);
nand U12069 (N_12069,N_5297,N_2555);
nand U12070 (N_12070,N_3460,N_1423);
or U12071 (N_12071,N_5634,N_1915);
nor U12072 (N_12072,N_3230,N_6142);
or U12073 (N_12073,N_842,N_1677);
or U12074 (N_12074,N_1443,N_2461);
nand U12075 (N_12075,N_1974,N_3976);
or U12076 (N_12076,N_1795,N_3026);
nand U12077 (N_12077,N_203,N_867);
nor U12078 (N_12078,N_6138,N_1352);
nor U12079 (N_12079,N_511,N_4305);
and U12080 (N_12080,N_5924,N_1928);
and U12081 (N_12081,N_5648,N_2231);
and U12082 (N_12082,N_4899,N_2568);
and U12083 (N_12083,N_5054,N_5449);
or U12084 (N_12084,N_1695,N_4936);
or U12085 (N_12085,N_3433,N_3735);
nor U12086 (N_12086,N_3857,N_3345);
nor U12087 (N_12087,N_5920,N_2322);
and U12088 (N_12088,N_4003,N_3021);
nor U12089 (N_12089,N_3182,N_2705);
and U12090 (N_12090,N_5634,N_4996);
and U12091 (N_12091,N_2339,N_198);
nand U12092 (N_12092,N_6207,N_2821);
nand U12093 (N_12093,N_5548,N_901);
nand U12094 (N_12094,N_5177,N_281);
or U12095 (N_12095,N_4326,N_5211);
nand U12096 (N_12096,N_5116,N_5670);
and U12097 (N_12097,N_5595,N_5067);
xor U12098 (N_12098,N_3572,N_5864);
nand U12099 (N_12099,N_5324,N_5645);
nand U12100 (N_12100,N_3914,N_4494);
and U12101 (N_12101,N_4883,N_1381);
and U12102 (N_12102,N_4970,N_607);
nand U12103 (N_12103,N_4342,N_4540);
nand U12104 (N_12104,N_2163,N_1984);
nand U12105 (N_12105,N_1291,N_712);
nand U12106 (N_12106,N_1297,N_3841);
and U12107 (N_12107,N_6063,N_1702);
and U12108 (N_12108,N_2922,N_2024);
and U12109 (N_12109,N_4793,N_679);
and U12110 (N_12110,N_1781,N_1474);
or U12111 (N_12111,N_283,N_3151);
and U12112 (N_12112,N_1223,N_197);
nand U12113 (N_12113,N_4473,N_2347);
nand U12114 (N_12114,N_1697,N_6118);
or U12115 (N_12115,N_6013,N_2104);
nor U12116 (N_12116,N_1530,N_4927);
nor U12117 (N_12117,N_1708,N_4086);
nor U12118 (N_12118,N_5627,N_5991);
nand U12119 (N_12119,N_4211,N_5784);
and U12120 (N_12120,N_314,N_5366);
and U12121 (N_12121,N_2164,N_4102);
and U12122 (N_12122,N_3995,N_4071);
nand U12123 (N_12123,N_3796,N_3372);
nand U12124 (N_12124,N_4065,N_1309);
and U12125 (N_12125,N_2898,N_897);
or U12126 (N_12126,N_3314,N_4541);
nand U12127 (N_12127,N_61,N_3892);
and U12128 (N_12128,N_906,N_5613);
and U12129 (N_12129,N_2394,N_3219);
nand U12130 (N_12130,N_4535,N_1488);
and U12131 (N_12131,N_559,N_3276);
or U12132 (N_12132,N_500,N_4832);
nand U12133 (N_12133,N_5114,N_3471);
and U12134 (N_12134,N_137,N_307);
or U12135 (N_12135,N_3878,N_3285);
and U12136 (N_12136,N_4364,N_3888);
nand U12137 (N_12137,N_1359,N_237);
nor U12138 (N_12138,N_5148,N_901);
nor U12139 (N_12139,N_5207,N_434);
and U12140 (N_12140,N_687,N_5243);
nor U12141 (N_12141,N_4994,N_237);
or U12142 (N_12142,N_3535,N_5994);
nand U12143 (N_12143,N_2421,N_3468);
nor U12144 (N_12144,N_5805,N_1416);
nor U12145 (N_12145,N_1973,N_5637);
and U12146 (N_12146,N_2363,N_5874);
nor U12147 (N_12147,N_1995,N_2754);
nand U12148 (N_12148,N_4772,N_4788);
nor U12149 (N_12149,N_5788,N_2749);
or U12150 (N_12150,N_2138,N_5012);
nor U12151 (N_12151,N_3153,N_6210);
and U12152 (N_12152,N_6068,N_4014);
nor U12153 (N_12153,N_5803,N_4441);
and U12154 (N_12154,N_2771,N_612);
nand U12155 (N_12155,N_3177,N_5193);
nor U12156 (N_12156,N_2691,N_5431);
or U12157 (N_12157,N_5327,N_3123);
and U12158 (N_12158,N_1051,N_2501);
nand U12159 (N_12159,N_1986,N_3345);
nand U12160 (N_12160,N_1170,N_113);
nand U12161 (N_12161,N_219,N_3808);
nand U12162 (N_12162,N_267,N_2095);
nor U12163 (N_12163,N_1311,N_3814);
nor U12164 (N_12164,N_2693,N_5023);
and U12165 (N_12165,N_5531,N_1692);
nor U12166 (N_12166,N_3109,N_884);
nand U12167 (N_12167,N_5270,N_1009);
or U12168 (N_12168,N_2785,N_3849);
nand U12169 (N_12169,N_2996,N_458);
nor U12170 (N_12170,N_930,N_3929);
nor U12171 (N_12171,N_1955,N_4053);
nor U12172 (N_12172,N_4636,N_4478);
nor U12173 (N_12173,N_3773,N_5057);
or U12174 (N_12174,N_4807,N_6229);
nor U12175 (N_12175,N_1917,N_1065);
nand U12176 (N_12176,N_2974,N_5911);
and U12177 (N_12177,N_847,N_252);
and U12178 (N_12178,N_5051,N_4853);
nand U12179 (N_12179,N_4720,N_5618);
nor U12180 (N_12180,N_4947,N_3987);
nor U12181 (N_12181,N_2586,N_1408);
xor U12182 (N_12182,N_4637,N_1578);
nand U12183 (N_12183,N_5211,N_2577);
or U12184 (N_12184,N_5072,N_4037);
nor U12185 (N_12185,N_4323,N_5128);
and U12186 (N_12186,N_4242,N_3519);
nor U12187 (N_12187,N_835,N_3717);
nor U12188 (N_12188,N_4671,N_5584);
nand U12189 (N_12189,N_4328,N_1409);
nand U12190 (N_12190,N_6012,N_532);
nand U12191 (N_12191,N_325,N_2776);
or U12192 (N_12192,N_5439,N_1137);
and U12193 (N_12193,N_3949,N_2147);
nand U12194 (N_12194,N_4794,N_5571);
and U12195 (N_12195,N_3490,N_1109);
and U12196 (N_12196,N_5766,N_1064);
nand U12197 (N_12197,N_1936,N_2852);
nand U12198 (N_12198,N_4760,N_5677);
or U12199 (N_12199,N_1217,N_6004);
nand U12200 (N_12200,N_2272,N_3364);
nor U12201 (N_12201,N_1275,N_1425);
or U12202 (N_12202,N_2216,N_4956);
and U12203 (N_12203,N_6143,N_3639);
nor U12204 (N_12204,N_4641,N_4695);
nand U12205 (N_12205,N_3035,N_5895);
nor U12206 (N_12206,N_1784,N_3411);
or U12207 (N_12207,N_5765,N_6051);
nand U12208 (N_12208,N_1874,N_3513);
and U12209 (N_12209,N_5071,N_5503);
and U12210 (N_12210,N_269,N_3183);
nand U12211 (N_12211,N_5049,N_2367);
nand U12212 (N_12212,N_4018,N_776);
or U12213 (N_12213,N_4503,N_3279);
and U12214 (N_12214,N_4632,N_3331);
and U12215 (N_12215,N_5245,N_3556);
or U12216 (N_12216,N_5994,N_4578);
nand U12217 (N_12217,N_5873,N_5840);
and U12218 (N_12218,N_1336,N_69);
and U12219 (N_12219,N_1414,N_1965);
and U12220 (N_12220,N_5362,N_6125);
nand U12221 (N_12221,N_2,N_3188);
nand U12222 (N_12222,N_3681,N_2248);
nor U12223 (N_12223,N_3481,N_7);
or U12224 (N_12224,N_935,N_5884);
or U12225 (N_12225,N_5397,N_4709);
nand U12226 (N_12226,N_831,N_2819);
and U12227 (N_12227,N_3638,N_1540);
nand U12228 (N_12228,N_4747,N_2862);
nor U12229 (N_12229,N_1338,N_1283);
nor U12230 (N_12230,N_6210,N_27);
nor U12231 (N_12231,N_5201,N_4077);
nor U12232 (N_12232,N_5231,N_635);
and U12233 (N_12233,N_2067,N_1739);
nand U12234 (N_12234,N_4953,N_3369);
nor U12235 (N_12235,N_5963,N_3988);
nor U12236 (N_12236,N_3588,N_5609);
nand U12237 (N_12237,N_3596,N_2667);
or U12238 (N_12238,N_1577,N_2821);
nor U12239 (N_12239,N_6082,N_839);
or U12240 (N_12240,N_389,N_4441);
nor U12241 (N_12241,N_5290,N_2796);
nor U12242 (N_12242,N_2968,N_3693);
and U12243 (N_12243,N_1739,N_2423);
and U12244 (N_12244,N_3110,N_3243);
and U12245 (N_12245,N_6065,N_2204);
nand U12246 (N_12246,N_4178,N_5670);
nor U12247 (N_12247,N_4968,N_5370);
nand U12248 (N_12248,N_2096,N_2683);
nand U12249 (N_12249,N_1426,N_3966);
nor U12250 (N_12250,N_3657,N_4081);
nor U12251 (N_12251,N_5743,N_3946);
and U12252 (N_12252,N_290,N_697);
and U12253 (N_12253,N_4567,N_6045);
nand U12254 (N_12254,N_5237,N_4083);
or U12255 (N_12255,N_5929,N_2055);
nor U12256 (N_12256,N_3604,N_3209);
nor U12257 (N_12257,N_1273,N_2227);
or U12258 (N_12258,N_5526,N_4067);
nor U12259 (N_12259,N_719,N_5863);
nand U12260 (N_12260,N_845,N_6090);
or U12261 (N_12261,N_1085,N_4820);
or U12262 (N_12262,N_2600,N_3356);
nor U12263 (N_12263,N_1214,N_5771);
and U12264 (N_12264,N_1114,N_159);
and U12265 (N_12265,N_2131,N_2221);
and U12266 (N_12266,N_1146,N_4009);
or U12267 (N_12267,N_1228,N_1782);
or U12268 (N_12268,N_5897,N_2179);
nor U12269 (N_12269,N_1655,N_6183);
or U12270 (N_12270,N_1868,N_250);
nor U12271 (N_12271,N_134,N_2281);
nor U12272 (N_12272,N_3058,N_553);
or U12273 (N_12273,N_2931,N_1094);
nand U12274 (N_12274,N_3071,N_3839);
and U12275 (N_12275,N_4976,N_5972);
nand U12276 (N_12276,N_3934,N_2074);
nor U12277 (N_12277,N_579,N_501);
nand U12278 (N_12278,N_2988,N_3634);
or U12279 (N_12279,N_2157,N_303);
nor U12280 (N_12280,N_5188,N_2605);
nand U12281 (N_12281,N_5992,N_3273);
nand U12282 (N_12282,N_1508,N_3806);
or U12283 (N_12283,N_1133,N_2845);
nor U12284 (N_12284,N_3179,N_1962);
nor U12285 (N_12285,N_2565,N_4646);
or U12286 (N_12286,N_3303,N_2069);
and U12287 (N_12287,N_4728,N_3371);
nand U12288 (N_12288,N_5228,N_4715);
or U12289 (N_12289,N_255,N_1873);
nand U12290 (N_12290,N_3128,N_6161);
nand U12291 (N_12291,N_50,N_3014);
or U12292 (N_12292,N_1612,N_889);
or U12293 (N_12293,N_4549,N_1398);
or U12294 (N_12294,N_3041,N_808);
nand U12295 (N_12295,N_1782,N_1199);
or U12296 (N_12296,N_2019,N_2129);
and U12297 (N_12297,N_4954,N_5365);
nor U12298 (N_12298,N_3215,N_1884);
or U12299 (N_12299,N_3147,N_1351);
nand U12300 (N_12300,N_1760,N_3927);
or U12301 (N_12301,N_1762,N_1966);
or U12302 (N_12302,N_5242,N_3282);
nor U12303 (N_12303,N_487,N_2706);
or U12304 (N_12304,N_4409,N_1175);
or U12305 (N_12305,N_5716,N_2103);
nor U12306 (N_12306,N_2490,N_4904);
and U12307 (N_12307,N_4856,N_1520);
and U12308 (N_12308,N_1252,N_4674);
and U12309 (N_12309,N_4060,N_2861);
nor U12310 (N_12310,N_2056,N_1889);
xor U12311 (N_12311,N_1530,N_1520);
or U12312 (N_12312,N_4573,N_2855);
or U12313 (N_12313,N_1021,N_743);
nand U12314 (N_12314,N_4517,N_3442);
and U12315 (N_12315,N_4446,N_3110);
nor U12316 (N_12316,N_23,N_1625);
and U12317 (N_12317,N_1221,N_3277);
or U12318 (N_12318,N_132,N_2322);
nor U12319 (N_12319,N_5890,N_4742);
and U12320 (N_12320,N_912,N_2396);
nor U12321 (N_12321,N_3370,N_171);
xnor U12322 (N_12322,N_3200,N_4793);
or U12323 (N_12323,N_3874,N_6132);
nor U12324 (N_12324,N_1058,N_2185);
nor U12325 (N_12325,N_3388,N_1481);
or U12326 (N_12326,N_1430,N_4637);
or U12327 (N_12327,N_6144,N_3232);
or U12328 (N_12328,N_2248,N_1410);
or U12329 (N_12329,N_1840,N_1884);
xnor U12330 (N_12330,N_3367,N_2210);
or U12331 (N_12331,N_5497,N_237);
nand U12332 (N_12332,N_1021,N_2752);
nand U12333 (N_12333,N_813,N_1533);
and U12334 (N_12334,N_4467,N_5916);
nand U12335 (N_12335,N_5914,N_2791);
nand U12336 (N_12336,N_2476,N_223);
and U12337 (N_12337,N_1083,N_4812);
and U12338 (N_12338,N_3513,N_4435);
and U12339 (N_12339,N_2395,N_613);
and U12340 (N_12340,N_350,N_3473);
and U12341 (N_12341,N_5787,N_5179);
nand U12342 (N_12342,N_4240,N_502);
or U12343 (N_12343,N_1686,N_1889);
nor U12344 (N_12344,N_3578,N_1620);
and U12345 (N_12345,N_2986,N_2707);
and U12346 (N_12346,N_418,N_3390);
nor U12347 (N_12347,N_5037,N_193);
and U12348 (N_12348,N_2946,N_1512);
or U12349 (N_12349,N_1465,N_2579);
and U12350 (N_12350,N_2216,N_6120);
nor U12351 (N_12351,N_2237,N_3603);
or U12352 (N_12352,N_3487,N_4802);
nand U12353 (N_12353,N_3846,N_1368);
nor U12354 (N_12354,N_4848,N_2451);
and U12355 (N_12355,N_2771,N_2388);
or U12356 (N_12356,N_4234,N_4765);
nor U12357 (N_12357,N_5391,N_405);
nand U12358 (N_12358,N_2282,N_5608);
nor U12359 (N_12359,N_3151,N_6019);
nand U12360 (N_12360,N_3685,N_4152);
nor U12361 (N_12361,N_5330,N_1061);
or U12362 (N_12362,N_4559,N_4807);
and U12363 (N_12363,N_2679,N_4187);
nand U12364 (N_12364,N_1258,N_1191);
nand U12365 (N_12365,N_4182,N_4509);
nand U12366 (N_12366,N_2559,N_640);
nand U12367 (N_12367,N_0,N_3031);
and U12368 (N_12368,N_2694,N_3472);
or U12369 (N_12369,N_2861,N_3699);
nor U12370 (N_12370,N_669,N_1140);
nand U12371 (N_12371,N_1629,N_681);
nand U12372 (N_12372,N_1599,N_4022);
nand U12373 (N_12373,N_5934,N_1605);
and U12374 (N_12374,N_4115,N_5964);
nor U12375 (N_12375,N_471,N_5634);
or U12376 (N_12376,N_5415,N_2252);
or U12377 (N_12377,N_5060,N_3434);
nor U12378 (N_12378,N_4579,N_4373);
and U12379 (N_12379,N_5736,N_1036);
or U12380 (N_12380,N_4665,N_5190);
and U12381 (N_12381,N_5862,N_5063);
nand U12382 (N_12382,N_1122,N_3608);
and U12383 (N_12383,N_5401,N_1748);
nor U12384 (N_12384,N_304,N_5746);
nand U12385 (N_12385,N_6006,N_2479);
xor U12386 (N_12386,N_2071,N_1237);
nor U12387 (N_12387,N_857,N_2381);
nand U12388 (N_12388,N_5204,N_1286);
and U12389 (N_12389,N_4760,N_1580);
or U12390 (N_12390,N_3250,N_4640);
nor U12391 (N_12391,N_579,N_4982);
or U12392 (N_12392,N_4213,N_413);
nor U12393 (N_12393,N_1550,N_1385);
or U12394 (N_12394,N_3172,N_45);
or U12395 (N_12395,N_382,N_5602);
nor U12396 (N_12396,N_2520,N_6172);
nand U12397 (N_12397,N_3796,N_3869);
nor U12398 (N_12398,N_3580,N_4353);
nor U12399 (N_12399,N_5105,N_1447);
nor U12400 (N_12400,N_3209,N_242);
nand U12401 (N_12401,N_423,N_2551);
nand U12402 (N_12402,N_2792,N_4049);
nor U12403 (N_12403,N_1286,N_3242);
and U12404 (N_12404,N_4568,N_364);
nor U12405 (N_12405,N_4744,N_4290);
nand U12406 (N_12406,N_5782,N_826);
nor U12407 (N_12407,N_4406,N_4053);
or U12408 (N_12408,N_4426,N_4422);
or U12409 (N_12409,N_3637,N_1916);
or U12410 (N_12410,N_2411,N_3089);
or U12411 (N_12411,N_5757,N_1455);
nand U12412 (N_12412,N_5853,N_5816);
and U12413 (N_12413,N_608,N_5534);
nand U12414 (N_12414,N_3136,N_3904);
nand U12415 (N_12415,N_1998,N_2201);
nor U12416 (N_12416,N_2689,N_212);
nand U12417 (N_12417,N_1581,N_5200);
or U12418 (N_12418,N_2264,N_125);
or U12419 (N_12419,N_3516,N_2341);
nor U12420 (N_12420,N_4058,N_1233);
nand U12421 (N_12421,N_5480,N_3401);
and U12422 (N_12422,N_763,N_4489);
nor U12423 (N_12423,N_4866,N_5207);
nand U12424 (N_12424,N_3234,N_5644);
or U12425 (N_12425,N_3190,N_513);
and U12426 (N_12426,N_1678,N_5783);
nand U12427 (N_12427,N_1515,N_4594);
and U12428 (N_12428,N_1172,N_1254);
and U12429 (N_12429,N_2758,N_2866);
and U12430 (N_12430,N_329,N_3320);
nor U12431 (N_12431,N_687,N_2625);
nand U12432 (N_12432,N_232,N_3062);
and U12433 (N_12433,N_3863,N_5256);
and U12434 (N_12434,N_4260,N_5377);
nor U12435 (N_12435,N_1391,N_5702);
and U12436 (N_12436,N_4312,N_1171);
nand U12437 (N_12437,N_4546,N_943);
nand U12438 (N_12438,N_3356,N_1810);
nand U12439 (N_12439,N_5730,N_2335);
nand U12440 (N_12440,N_50,N_4331);
and U12441 (N_12441,N_6204,N_4433);
and U12442 (N_12442,N_6106,N_2655);
nor U12443 (N_12443,N_777,N_1056);
or U12444 (N_12444,N_2677,N_4013);
and U12445 (N_12445,N_3732,N_1787);
nor U12446 (N_12446,N_3527,N_3169);
nand U12447 (N_12447,N_4336,N_5878);
nor U12448 (N_12448,N_5479,N_4210);
nand U12449 (N_12449,N_3966,N_2049);
nand U12450 (N_12450,N_5358,N_1882);
nand U12451 (N_12451,N_554,N_5584);
and U12452 (N_12452,N_1649,N_3089);
nand U12453 (N_12453,N_5664,N_1666);
and U12454 (N_12454,N_3604,N_1640);
nor U12455 (N_12455,N_3887,N_4648);
nor U12456 (N_12456,N_4017,N_2782);
nor U12457 (N_12457,N_4788,N_5616);
and U12458 (N_12458,N_2453,N_1050);
or U12459 (N_12459,N_1540,N_1150);
xor U12460 (N_12460,N_6242,N_1426);
nand U12461 (N_12461,N_2862,N_1984);
nor U12462 (N_12462,N_1171,N_5401);
nand U12463 (N_12463,N_2393,N_3641);
or U12464 (N_12464,N_165,N_4144);
and U12465 (N_12465,N_452,N_2982);
nor U12466 (N_12466,N_1989,N_3994);
nor U12467 (N_12467,N_1828,N_5742);
nand U12468 (N_12468,N_1667,N_4949);
and U12469 (N_12469,N_4135,N_5418);
nor U12470 (N_12470,N_3178,N_4069);
nand U12471 (N_12471,N_6125,N_1847);
or U12472 (N_12472,N_4714,N_3827);
or U12473 (N_12473,N_5855,N_2264);
nor U12474 (N_12474,N_5464,N_693);
or U12475 (N_12475,N_4961,N_198);
nand U12476 (N_12476,N_3559,N_4269);
or U12477 (N_12477,N_1560,N_1201);
and U12478 (N_12478,N_4963,N_4267);
or U12479 (N_12479,N_4203,N_299);
and U12480 (N_12480,N_1275,N_1400);
nand U12481 (N_12481,N_6205,N_3680);
xor U12482 (N_12482,N_795,N_2259);
nand U12483 (N_12483,N_1173,N_1848);
and U12484 (N_12484,N_5341,N_51);
and U12485 (N_12485,N_3403,N_3192);
or U12486 (N_12486,N_3833,N_4700);
or U12487 (N_12487,N_487,N_1135);
nand U12488 (N_12488,N_4126,N_3521);
nor U12489 (N_12489,N_5634,N_2324);
or U12490 (N_12490,N_4703,N_4550);
nor U12491 (N_12491,N_4185,N_3075);
nor U12492 (N_12492,N_1870,N_4642);
xnor U12493 (N_12493,N_4975,N_4347);
and U12494 (N_12494,N_3710,N_2578);
or U12495 (N_12495,N_4147,N_1685);
nor U12496 (N_12496,N_2800,N_2439);
nor U12497 (N_12497,N_5088,N_1059);
nor U12498 (N_12498,N_3448,N_2050);
nor U12499 (N_12499,N_1439,N_1921);
or U12500 (N_12500,N_6835,N_8351);
and U12501 (N_12501,N_6978,N_11220);
nor U12502 (N_12502,N_11570,N_11985);
or U12503 (N_12503,N_9990,N_11502);
nor U12504 (N_12504,N_11568,N_9751);
nand U12505 (N_12505,N_7697,N_8771);
or U12506 (N_12506,N_12156,N_11745);
nand U12507 (N_12507,N_8969,N_11298);
nor U12508 (N_12508,N_8499,N_11226);
nor U12509 (N_12509,N_11749,N_8739);
and U12510 (N_12510,N_11256,N_12296);
or U12511 (N_12511,N_8719,N_11402);
and U12512 (N_12512,N_7449,N_7988);
and U12513 (N_12513,N_10830,N_9583);
or U12514 (N_12514,N_12030,N_11931);
nand U12515 (N_12515,N_10054,N_11387);
or U12516 (N_12516,N_9523,N_10484);
and U12517 (N_12517,N_10632,N_7848);
nand U12518 (N_12518,N_9397,N_12134);
and U12519 (N_12519,N_10396,N_8444);
nor U12520 (N_12520,N_11529,N_9882);
nor U12521 (N_12521,N_8293,N_11815);
nand U12522 (N_12522,N_9134,N_10862);
nor U12523 (N_12523,N_9365,N_9889);
and U12524 (N_12524,N_11277,N_10113);
nand U12525 (N_12525,N_6665,N_9071);
nor U12526 (N_12526,N_12300,N_8019);
nand U12527 (N_12527,N_9166,N_9822);
and U12528 (N_12528,N_12153,N_11487);
nand U12529 (N_12529,N_11305,N_6683);
or U12530 (N_12530,N_8613,N_7524);
or U12531 (N_12531,N_9775,N_6760);
or U12532 (N_12532,N_7700,N_9031);
and U12533 (N_12533,N_12363,N_10633);
or U12534 (N_12534,N_9307,N_9434);
nand U12535 (N_12535,N_9262,N_9660);
and U12536 (N_12536,N_11788,N_6552);
nand U12537 (N_12537,N_8225,N_7289);
or U12538 (N_12538,N_6253,N_10886);
or U12539 (N_12539,N_8948,N_11349);
or U12540 (N_12540,N_9180,N_8508);
nand U12541 (N_12541,N_6932,N_6620);
nor U12542 (N_12542,N_6447,N_11944);
or U12543 (N_12543,N_10177,N_8909);
and U12544 (N_12544,N_7963,N_9511);
or U12545 (N_12545,N_7896,N_8375);
nor U12546 (N_12546,N_8610,N_7716);
or U12547 (N_12547,N_11857,N_8215);
xnor U12548 (N_12548,N_6561,N_10142);
nand U12549 (N_12549,N_10023,N_8116);
nor U12550 (N_12550,N_8320,N_9518);
nor U12551 (N_12551,N_7266,N_7993);
and U12552 (N_12552,N_10731,N_8946);
or U12553 (N_12553,N_7547,N_9119);
nor U12554 (N_12554,N_12341,N_12447);
or U12555 (N_12555,N_6714,N_9426);
and U12556 (N_12556,N_9162,N_7117);
or U12557 (N_12557,N_6369,N_9924);
and U12558 (N_12558,N_10323,N_6356);
nand U12559 (N_12559,N_11526,N_7960);
or U12560 (N_12560,N_9536,N_9576);
or U12561 (N_12561,N_8652,N_9627);
and U12562 (N_12562,N_9984,N_11683);
nor U12563 (N_12563,N_11284,N_11520);
and U12564 (N_12564,N_8608,N_10454);
and U12565 (N_12565,N_10612,N_10656);
nand U12566 (N_12566,N_12490,N_8891);
and U12567 (N_12567,N_8330,N_7044);
nand U12568 (N_12568,N_11562,N_8653);
nor U12569 (N_12569,N_12294,N_7277);
nand U12570 (N_12570,N_8047,N_7548);
or U12571 (N_12571,N_10541,N_12204);
and U12572 (N_12572,N_11746,N_6581);
nor U12573 (N_12573,N_9604,N_7638);
nor U12574 (N_12574,N_6686,N_7225);
and U12575 (N_12575,N_11968,N_6777);
or U12576 (N_12576,N_11177,N_9324);
or U12577 (N_12577,N_9163,N_6934);
or U12578 (N_12578,N_10451,N_9338);
and U12579 (N_12579,N_12269,N_6700);
nor U12580 (N_12580,N_9081,N_10893);
or U12581 (N_12581,N_8140,N_6399);
nor U12582 (N_12582,N_9326,N_9546);
or U12583 (N_12583,N_10006,N_11820);
nand U12584 (N_12584,N_7982,N_9645);
and U12585 (N_12585,N_9044,N_6646);
and U12586 (N_12586,N_12462,N_6829);
nor U12587 (N_12587,N_7345,N_12349);
and U12588 (N_12588,N_11433,N_7417);
or U12589 (N_12589,N_6555,N_7240);
or U12590 (N_12590,N_6264,N_7897);
nor U12591 (N_12591,N_11830,N_8014);
nor U12592 (N_12592,N_12351,N_8033);
nand U12593 (N_12593,N_7410,N_7967);
and U12594 (N_12594,N_8382,N_7713);
nand U12595 (N_12595,N_6342,N_11891);
nand U12596 (N_12596,N_6305,N_8677);
nand U12597 (N_12597,N_11583,N_9383);
nand U12598 (N_12598,N_12141,N_11948);
nor U12599 (N_12599,N_10179,N_10292);
nand U12600 (N_12600,N_9104,N_8241);
nor U12601 (N_12601,N_8711,N_8656);
nor U12602 (N_12602,N_8311,N_12177);
and U12603 (N_12603,N_6675,N_9605);
or U12604 (N_12604,N_9690,N_7696);
nand U12605 (N_12605,N_6973,N_9347);
or U12606 (N_12606,N_8478,N_10297);
or U12607 (N_12607,N_11086,N_11032);
nor U12608 (N_12608,N_6506,N_10393);
nand U12609 (N_12609,N_7540,N_8841);
nand U12610 (N_12610,N_8319,N_9580);
and U12611 (N_12611,N_7767,N_9143);
nor U12612 (N_12612,N_9149,N_10132);
nor U12613 (N_12613,N_12012,N_8349);
nor U12614 (N_12614,N_8437,N_8269);
nor U12615 (N_12615,N_7204,N_11597);
nor U12616 (N_12616,N_11862,N_7118);
nand U12617 (N_12617,N_8815,N_12347);
and U12618 (N_12618,N_10681,N_10997);
or U12619 (N_12619,N_9320,N_10324);
or U12620 (N_12620,N_8883,N_8257);
and U12621 (N_12621,N_7925,N_7274);
nand U12622 (N_12622,N_8045,N_9389);
and U12623 (N_12623,N_8229,N_8192);
or U12624 (N_12624,N_8171,N_9670);
nor U12625 (N_12625,N_8724,N_9493);
nand U12626 (N_12626,N_11809,N_7581);
nand U12627 (N_12627,N_10486,N_12352);
or U12628 (N_12628,N_9284,N_7336);
and U12629 (N_12629,N_10707,N_8826);
nand U12630 (N_12630,N_10709,N_7811);
or U12631 (N_12631,N_7920,N_8957);
nand U12632 (N_12632,N_8600,N_10895);
and U12633 (N_12633,N_7987,N_10404);
or U12634 (N_12634,N_11818,N_10090);
and U12635 (N_12635,N_8298,N_9209);
or U12636 (N_12636,N_7416,N_11093);
nor U12637 (N_12637,N_8121,N_9745);
nand U12638 (N_12638,N_7671,N_10987);
and U12639 (N_12639,N_10599,N_9728);
or U12640 (N_12640,N_7455,N_11539);
nand U12641 (N_12641,N_8895,N_10028);
and U12642 (N_12642,N_10473,N_10435);
nor U12643 (N_12643,N_6458,N_8642);
or U12644 (N_12644,N_12094,N_8956);
and U12645 (N_12645,N_10736,N_11447);
nor U12646 (N_12646,N_10410,N_11538);
or U12647 (N_12647,N_8862,N_10316);
nor U12648 (N_12648,N_12354,N_7698);
or U12649 (N_12649,N_7728,N_6509);
nand U12650 (N_12650,N_10346,N_9385);
nand U12651 (N_12651,N_8119,N_6761);
nand U12652 (N_12652,N_6940,N_10180);
nor U12653 (N_12653,N_7928,N_11950);
xor U12654 (N_12654,N_10207,N_7699);
nand U12655 (N_12655,N_10703,N_10252);
nor U12656 (N_12656,N_8494,N_11789);
or U12657 (N_12657,N_7487,N_12144);
and U12658 (N_12658,N_12223,N_9086);
or U12659 (N_12659,N_10982,N_9483);
nand U12660 (N_12660,N_8186,N_12365);
nor U12661 (N_12661,N_12053,N_7677);
nand U12662 (N_12662,N_9520,N_8503);
nand U12663 (N_12663,N_11849,N_10691);
nand U12664 (N_12664,N_12113,N_7043);
and U12665 (N_12665,N_6582,N_6560);
nor U12666 (N_12666,N_7961,N_11922);
and U12667 (N_12667,N_12398,N_6601);
nor U12668 (N_12668,N_11676,N_8052);
and U12669 (N_12669,N_7860,N_6907);
or U12670 (N_12670,N_10885,N_11601);
nand U12671 (N_12671,N_11420,N_8143);
or U12672 (N_12672,N_6698,N_7629);
nand U12673 (N_12673,N_11840,N_9563);
nand U12674 (N_12674,N_9159,N_9155);
nor U12675 (N_12675,N_9746,N_7862);
nand U12676 (N_12676,N_11154,N_6833);
or U12677 (N_12677,N_9894,N_8367);
or U12678 (N_12678,N_9409,N_8604);
nand U12679 (N_12679,N_10569,N_7907);
nor U12680 (N_12680,N_9261,N_6810);
and U12681 (N_12681,N_11358,N_9363);
nor U12682 (N_12682,N_9063,N_9758);
nor U12683 (N_12683,N_7892,N_7795);
nand U12684 (N_12684,N_9457,N_9016);
and U12685 (N_12685,N_6598,N_11659);
nand U12686 (N_12686,N_10212,N_7190);
nand U12687 (N_12687,N_10872,N_9350);
and U12688 (N_12688,N_9931,N_9288);
nand U12689 (N_12689,N_7506,N_9800);
and U12690 (N_12690,N_7932,N_7396);
or U12691 (N_12691,N_8778,N_10072);
or U12692 (N_12692,N_10235,N_11832);
and U12693 (N_12693,N_10881,N_8445);
and U12694 (N_12694,N_7634,N_8369);
or U12695 (N_12695,N_9755,N_6470);
and U12696 (N_12696,N_11991,N_10930);
nand U12697 (N_12697,N_9242,N_7496);
and U12698 (N_12698,N_10593,N_6652);
and U12699 (N_12699,N_7992,N_10337);
xnor U12700 (N_12700,N_10947,N_10099);
and U12701 (N_12701,N_11463,N_10539);
nor U12702 (N_12702,N_10327,N_7591);
nand U12703 (N_12703,N_7062,N_8168);
and U12704 (N_12704,N_6604,N_8864);
or U12705 (N_12705,N_10036,N_9172);
nor U12706 (N_12706,N_6728,N_10827);
nor U12707 (N_12707,N_6405,N_7006);
and U12708 (N_12708,N_10136,N_10077);
or U12709 (N_12709,N_8422,N_11466);
or U12710 (N_12710,N_11039,N_7531);
nand U12711 (N_12711,N_11636,N_12071);
nor U12712 (N_12712,N_10956,N_11231);
nor U12713 (N_12713,N_8383,N_11361);
nand U12714 (N_12714,N_8871,N_8731);
nor U12715 (N_12715,N_8718,N_10230);
and U12716 (N_12716,N_6637,N_11351);
nor U12717 (N_12717,N_6417,N_11312);
or U12718 (N_12718,N_8307,N_8828);
nor U12719 (N_12719,N_10777,N_6880);
nor U12720 (N_12720,N_11962,N_7420);
and U12721 (N_12721,N_9617,N_9628);
nor U12722 (N_12722,N_10066,N_8408);
or U12723 (N_12723,N_7340,N_9414);
and U12724 (N_12724,N_10138,N_7317);
and U12725 (N_12725,N_9183,N_10260);
and U12726 (N_12726,N_6712,N_6296);
or U12727 (N_12727,N_9140,N_11582);
or U12728 (N_12728,N_7285,N_7426);
and U12729 (N_12729,N_12493,N_8843);
nand U12730 (N_12730,N_9561,N_10994);
nor U12731 (N_12731,N_9814,N_11490);
nor U12732 (N_12732,N_12492,N_8686);
nand U12733 (N_12733,N_11814,N_9689);
and U12734 (N_12734,N_12456,N_8262);
nand U12735 (N_12735,N_8451,N_9494);
or U12736 (N_12736,N_7724,N_6870);
or U12737 (N_12737,N_11059,N_9080);
or U12738 (N_12738,N_8616,N_9132);
and U12739 (N_12739,N_10915,N_12416);
nand U12740 (N_12740,N_9188,N_9330);
and U12741 (N_12741,N_9379,N_12389);
or U12742 (N_12742,N_6431,N_8628);
nor U12743 (N_12743,N_7397,N_11096);
nand U12744 (N_12744,N_12115,N_7181);
or U12745 (N_12745,N_6953,N_7816);
or U12746 (N_12746,N_11031,N_7511);
nand U12747 (N_12747,N_8285,N_7628);
and U12748 (N_12748,N_7352,N_10283);
nand U12749 (N_12749,N_8625,N_7199);
nand U12750 (N_12750,N_12298,N_9366);
or U12751 (N_12751,N_8425,N_10456);
or U12752 (N_12752,N_11495,N_8190);
and U12753 (N_12753,N_10576,N_7942);
and U12754 (N_12754,N_6867,N_11035);
nor U12755 (N_12755,N_7380,N_12087);
nand U12756 (N_12756,N_12104,N_12185);
and U12757 (N_12757,N_8372,N_10798);
nand U12758 (N_12758,N_9572,N_9684);
nor U12759 (N_12759,N_12034,N_8714);
xor U12760 (N_12760,N_7849,N_10874);
xnor U12761 (N_12761,N_7906,N_9396);
nand U12762 (N_12762,N_12186,N_8811);
or U12763 (N_12763,N_7479,N_8991);
or U12764 (N_12764,N_8857,N_10465);
nor U12765 (N_12765,N_8031,N_7284);
and U12766 (N_12766,N_7606,N_9908);
nand U12767 (N_12767,N_6877,N_7840);
or U12768 (N_12768,N_11537,N_10095);
nand U12769 (N_12769,N_11384,N_9671);
or U12770 (N_12770,N_11374,N_11533);
nor U12771 (N_12771,N_10556,N_9023);
xnor U12772 (N_12772,N_11721,N_9232);
nor U12773 (N_12773,N_10332,N_6545);
and U12774 (N_12774,N_10358,N_11038);
or U12775 (N_12775,N_8315,N_9423);
nor U12776 (N_12776,N_10640,N_8709);
or U12777 (N_12777,N_8475,N_12078);
nand U12778 (N_12778,N_7601,N_11262);
or U12779 (N_12779,N_7176,N_7279);
nor U12780 (N_12780,N_7879,N_9404);
or U12781 (N_12781,N_8465,N_9880);
nor U12782 (N_12782,N_9972,N_9007);
nand U12783 (N_12783,N_8107,N_9226);
nand U12784 (N_12784,N_8187,N_9705);
nor U12785 (N_12785,N_6947,N_9272);
nand U12786 (N_12786,N_10502,N_7807);
xor U12787 (N_12787,N_11665,N_8887);
nor U12788 (N_12788,N_11345,N_12457);
nor U12789 (N_12789,N_10610,N_8943);
and U12790 (N_12790,N_9344,N_12208);
or U12791 (N_12791,N_8491,N_7275);
nor U12792 (N_12792,N_9106,N_8310);
nand U12793 (N_12793,N_11354,N_10903);
nor U12794 (N_12794,N_7105,N_10091);
and U12795 (N_12795,N_11506,N_9308);
and U12796 (N_12796,N_10365,N_9555);
or U12797 (N_12797,N_6388,N_8550);
nor U12798 (N_12798,N_10457,N_8687);
and U12799 (N_12799,N_7950,N_7883);
and U12800 (N_12800,N_6954,N_9051);
nor U12801 (N_12801,N_7758,N_11939);
xor U12802 (N_12802,N_12148,N_6852);
or U12803 (N_12803,N_12130,N_8081);
and U12804 (N_12804,N_8230,N_9150);
nand U12805 (N_12805,N_9834,N_6471);
nor U12806 (N_12806,N_8384,N_9060);
or U12807 (N_12807,N_9939,N_8644);
nor U12808 (N_12808,N_12449,N_10354);
nand U12809 (N_12809,N_8231,N_9817);
nand U12810 (N_12810,N_6721,N_6386);
nor U12811 (N_12811,N_10050,N_9102);
nor U12812 (N_12812,N_12424,N_11435);
or U12813 (N_12813,N_6812,N_7528);
and U12814 (N_12814,N_8313,N_11839);
nor U12815 (N_12815,N_10437,N_9443);
or U12816 (N_12816,N_10149,N_11916);
nor U12817 (N_12817,N_8865,N_9754);
or U12818 (N_12818,N_6278,N_8403);
nand U12819 (N_12819,N_11450,N_11586);
or U12820 (N_12820,N_9360,N_6363);
nand U12821 (N_12821,N_6772,N_10755);
nand U12822 (N_12822,N_10712,N_10168);
and U12823 (N_12823,N_6821,N_9146);
nand U12824 (N_12824,N_9790,N_7341);
and U12825 (N_12825,N_10559,N_9400);
and U12826 (N_12826,N_7566,N_9903);
or U12827 (N_12827,N_6496,N_11474);
nor U12828 (N_12828,N_11011,N_7908);
nand U12829 (N_12829,N_10127,N_9210);
nor U12830 (N_12830,N_7372,N_11851);
or U12831 (N_12831,N_10772,N_6962);
and U12832 (N_12832,N_9005,N_6690);
nand U12833 (N_12833,N_11760,N_10514);
or U12834 (N_12834,N_7298,N_6883);
nand U12835 (N_12835,N_7159,N_7823);
and U12836 (N_12836,N_9100,N_8777);
nand U12837 (N_12837,N_7440,N_8779);
nand U12838 (N_12838,N_10469,N_9057);
or U12839 (N_12839,N_9652,N_10905);
or U12840 (N_12840,N_10756,N_8222);
or U12841 (N_12841,N_11124,N_8048);
and U12842 (N_12842,N_12473,N_10550);
nand U12843 (N_12843,N_10685,N_6890);
nor U12844 (N_12844,N_7989,N_10421);
nand U12845 (N_12845,N_7246,N_10290);
nand U12846 (N_12846,N_9448,N_6519);
or U12847 (N_12847,N_7639,N_12353);
and U12848 (N_12848,N_7088,N_8025);
and U12849 (N_12849,N_12461,N_12238);
nor U12850 (N_12850,N_6446,N_7565);
nand U12851 (N_12851,N_10866,N_7291);
and U12852 (N_12852,N_6924,N_10374);
nand U12853 (N_12853,N_6271,N_6437);
or U12854 (N_12854,N_7363,N_6332);
nor U12855 (N_12855,N_10345,N_7166);
nor U12856 (N_12856,N_10934,N_10578);
xor U12857 (N_12857,N_9666,N_11322);
or U12858 (N_12858,N_8660,N_8717);
nor U12859 (N_12859,N_7708,N_8833);
and U12860 (N_12860,N_6977,N_6827);
or U12861 (N_12861,N_9571,N_7114);
and U12862 (N_12862,N_9152,N_7448);
nor U12863 (N_12863,N_12033,N_6902);
nand U12864 (N_12864,N_10797,N_6532);
xnor U12865 (N_12865,N_6935,N_8200);
or U12866 (N_12866,N_7796,N_12463);
or U12867 (N_12867,N_11373,N_9439);
nor U12868 (N_12868,N_8510,N_11368);
or U12869 (N_12869,N_7308,N_12045);
or U12870 (N_12870,N_8481,N_10119);
nor U12871 (N_12871,N_7733,N_8501);
nand U12872 (N_12872,N_10543,N_9487);
nand U12873 (N_12873,N_10892,N_7342);
or U12874 (N_12874,N_11855,N_7598);
nor U12875 (N_12875,N_11097,N_8623);
and U12876 (N_12876,N_9227,N_10496);
and U12877 (N_12877,N_9851,N_10686);
or U12878 (N_12878,N_6494,N_7149);
nand U12879 (N_12879,N_7456,N_11195);
or U12880 (N_12880,N_11221,N_7666);
nor U12881 (N_12881,N_10694,N_12011);
and U12882 (N_12882,N_8825,N_11873);
nor U12883 (N_12883,N_9127,N_10482);
or U12884 (N_12884,N_9663,N_11692);
nand U12885 (N_12885,N_8654,N_12301);
and U12886 (N_12886,N_6438,N_7517);
nor U12887 (N_12887,N_10553,N_6265);
nand U12888 (N_12888,N_8577,N_11217);
and U12889 (N_12889,N_10644,N_7061);
nor U12890 (N_12890,N_9356,N_7624);
nand U12891 (N_12891,N_12304,N_9773);
and U12892 (N_12892,N_11489,N_11165);
and U12893 (N_12893,N_9374,N_6487);
nor U12894 (N_12894,N_9316,N_10989);
nand U12895 (N_12895,N_7099,N_7066);
and U12896 (N_12896,N_10926,N_9378);
nor U12897 (N_12897,N_10720,N_7838);
or U12898 (N_12898,N_6457,N_8409);
or U12899 (N_12899,N_6988,N_7136);
or U12900 (N_12900,N_9954,N_7331);
nand U12901 (N_12901,N_7025,N_6539);
and U12902 (N_12902,N_12357,N_9273);
nor U12903 (N_12903,N_10745,N_9793);
or U12904 (N_12904,N_10370,N_10222);
nand U12905 (N_12905,N_8632,N_7570);
and U12906 (N_12906,N_11107,N_12433);
and U12907 (N_12907,N_6345,N_6644);
nand U12908 (N_12908,N_7916,N_10174);
nor U12909 (N_12909,N_9535,N_8939);
nor U12910 (N_12910,N_6694,N_8587);
nor U12911 (N_12911,N_12391,N_7371);
nand U12912 (N_12912,N_9805,N_6389);
and U12913 (N_12913,N_7450,N_10846);
nand U12914 (N_12914,N_9749,N_12097);
nor U12915 (N_12915,N_12236,N_10342);
nand U12916 (N_12916,N_8721,N_7194);
or U12917 (N_12917,N_6705,N_10737);
and U12918 (N_12918,N_11933,N_11941);
and U12919 (N_12919,N_9642,N_11075);
or U12920 (N_12920,N_10999,N_8162);
or U12921 (N_12921,N_6856,N_8922);
or U12922 (N_12922,N_7490,N_8633);
and U12923 (N_12923,N_10536,N_10206);
and U12924 (N_12924,N_8504,N_8804);
or U12925 (N_12925,N_12276,N_11112);
or U12926 (N_12926,N_9190,N_9274);
nand U12927 (N_12927,N_8339,N_11359);
nand U12928 (N_12928,N_6486,N_6882);
nand U12929 (N_12929,N_8688,N_9915);
and U12930 (N_12930,N_8264,N_6400);
nand U12931 (N_12931,N_11792,N_11268);
nand U12932 (N_12932,N_8356,N_9622);
nand U12933 (N_12933,N_8994,N_11067);
and U12934 (N_12934,N_11085,N_7922);
nand U12935 (N_12935,N_6570,N_8363);
nor U12936 (N_12936,N_10340,N_7924);
and U12937 (N_12937,N_7021,N_10778);
and U12938 (N_12938,N_9176,N_6781);
nand U12939 (N_12939,N_11653,N_10696);
nand U12940 (N_12940,N_9997,N_11657);
xor U12941 (N_12941,N_6307,N_8332);
nor U12942 (N_12942,N_11691,N_9646);
and U12943 (N_12943,N_9437,N_9711);
nand U12944 (N_12944,N_7832,N_11541);
nor U12945 (N_12945,N_12451,N_10019);
nor U12946 (N_12946,N_9926,N_11662);
or U12947 (N_12947,N_11591,N_11943);
nor U12948 (N_12948,N_6915,N_7281);
nor U12949 (N_12949,N_7974,N_9407);
nand U12950 (N_12950,N_10082,N_12388);
or U12951 (N_12951,N_10657,N_11751);
nand U12952 (N_12952,N_6943,N_6685);
or U12953 (N_12953,N_9737,N_10980);
or U12954 (N_12954,N_7884,N_7818);
nor U12955 (N_12955,N_10010,N_10996);
or U12956 (N_12956,N_11119,N_9394);
and U12957 (N_12957,N_10250,N_8505);
nand U12958 (N_12958,N_7693,N_6792);
nor U12959 (N_12959,N_10900,N_10652);
nand U12960 (N_12960,N_6270,N_9070);
or U12961 (N_12961,N_10475,N_7923);
nor U12962 (N_12962,N_11297,N_9083);
or U12963 (N_12963,N_10757,N_11010);
or U12964 (N_12964,N_7474,N_10181);
nor U12965 (N_12965,N_10913,N_9507);
nand U12966 (N_12966,N_6499,N_10427);
and U12967 (N_12967,N_9042,N_7355);
nand U12968 (N_12968,N_10616,N_8390);
or U12969 (N_12969,N_9818,N_11468);
or U12970 (N_12970,N_8745,N_12394);
and U12971 (N_12971,N_6252,N_7749);
or U12972 (N_12972,N_11030,N_8364);
nor U12973 (N_12973,N_8018,N_9381);
nand U12974 (N_12974,N_10746,N_6450);
and U12975 (N_12975,N_11560,N_10075);
nor U12976 (N_12976,N_9205,N_8884);
nand U12977 (N_12977,N_11757,N_11584);
or U12978 (N_12978,N_7541,N_11904);
or U12979 (N_12979,N_7615,N_8044);
nor U12980 (N_12980,N_9144,N_7940);
and U12981 (N_12981,N_12047,N_8598);
or U12982 (N_12982,N_8509,N_11281);
or U12983 (N_12983,N_10390,N_10600);
nand U12984 (N_12984,N_11151,N_9126);
and U12985 (N_12985,N_11323,N_7354);
nor U12986 (N_12986,N_8430,N_10574);
nor U12987 (N_12987,N_10840,N_8899);
and U12988 (N_12988,N_6351,N_6480);
and U12989 (N_12989,N_10984,N_8536);
or U12990 (N_12990,N_11684,N_11673);
or U12991 (N_12991,N_7134,N_10969);
nand U12992 (N_12992,N_12495,N_7734);
and U12993 (N_12993,N_11725,N_7673);
nor U12994 (N_12994,N_10405,N_8785);
and U12995 (N_12995,N_6502,N_6735);
or U12996 (N_12996,N_10057,N_11465);
or U12997 (N_12997,N_11767,N_9545);
nand U12998 (N_12998,N_11342,N_8017);
and U12999 (N_12999,N_9113,N_9852);
or U13000 (N_13000,N_6460,N_10619);
nand U13001 (N_13001,N_8157,N_9390);
or U13002 (N_13002,N_7217,N_6376);
and U13003 (N_13003,N_7357,N_10498);
or U13004 (N_13004,N_11810,N_7502);
and U13005 (N_13005,N_9469,N_11720);
nand U13006 (N_13006,N_10089,N_10279);
and U13007 (N_13007,N_9647,N_12323);
or U13008 (N_13008,N_9956,N_11174);
or U13009 (N_13009,N_9771,N_7241);
and U13010 (N_13010,N_12418,N_11385);
or U13011 (N_13011,N_7330,N_9677);
nor U13012 (N_13012,N_9743,N_7071);
xnor U13013 (N_13013,N_12412,N_6622);
nor U13014 (N_13014,N_12029,N_9524);
nand U13015 (N_13015,N_10339,N_9309);
and U13016 (N_13016,N_9003,N_9573);
nand U13017 (N_13017,N_10429,N_7781);
nand U13018 (N_13018,N_9436,N_6708);
xnor U13019 (N_13019,N_9593,N_9447);
and U13020 (N_13020,N_9768,N_7579);
or U13021 (N_13021,N_10397,N_10165);
nand U13022 (N_13022,N_12103,N_10237);
and U13023 (N_13023,N_8513,N_6908);
nor U13024 (N_13024,N_12225,N_9673);
or U13025 (N_13025,N_9683,N_12399);
nand U13026 (N_13026,N_6364,N_12214);
and U13027 (N_13027,N_9079,N_12263);
nand U13028 (N_13028,N_7023,N_8179);
nand U13029 (N_13029,N_10336,N_9154);
nor U13030 (N_13030,N_11303,N_10570);
nor U13031 (N_13031,N_11408,N_8129);
or U13032 (N_13032,N_9450,N_10007);
and U13033 (N_13033,N_10668,N_9577);
nand U13034 (N_13034,N_6930,N_11170);
nor U13035 (N_13035,N_6283,N_10051);
or U13036 (N_13036,N_9870,N_10045);
nor U13037 (N_13037,N_8152,N_8457);
and U13038 (N_13038,N_10304,N_6393);
or U13039 (N_13039,N_8112,N_7300);
nor U13040 (N_13040,N_7249,N_7829);
or U13041 (N_13041,N_6981,N_12282);
nor U13042 (N_13042,N_12261,N_9621);
and U13043 (N_13043,N_8767,N_8735);
xnor U13044 (N_13044,N_8885,N_10244);
nor U13045 (N_13045,N_8631,N_12197);
nand U13046 (N_13046,N_9293,N_11079);
nand U13047 (N_13047,N_8153,N_8428);
and U13048 (N_13048,N_9502,N_10937);
nand U13049 (N_13049,N_10972,N_8954);
nand U13050 (N_13050,N_10583,N_8933);
nand U13051 (N_13051,N_9987,N_10959);
or U13052 (N_13052,N_8461,N_8211);
and U13053 (N_13053,N_8882,N_8593);
and U13054 (N_13054,N_9492,N_8808);
nor U13055 (N_13055,N_11834,N_10992);
or U13056 (N_13056,N_7748,N_9836);
nand U13057 (N_13057,N_6803,N_6951);
nand U13058 (N_13058,N_9971,N_7686);
and U13059 (N_13059,N_10510,N_6731);
nand U13060 (N_13060,N_8636,N_6788);
nor U13061 (N_13061,N_9402,N_11234);
nand U13062 (N_13062,N_6628,N_8280);
nor U13063 (N_13063,N_11769,N_7076);
nand U13064 (N_13064,N_9674,N_8324);
or U13065 (N_13065,N_10192,N_6495);
and U13066 (N_13066,N_11971,N_7964);
nor U13067 (N_13067,N_7467,N_11599);
and U13068 (N_13068,N_11776,N_8358);
and U13069 (N_13069,N_6590,N_10938);
and U13070 (N_13070,N_12278,N_10790);
nand U13071 (N_13071,N_12243,N_10154);
nor U13072 (N_13072,N_11069,N_8122);
and U13073 (N_13073,N_10814,N_6613);
and U13074 (N_13074,N_12292,N_8174);
nand U13075 (N_13075,N_11740,N_9056);
and U13076 (N_13076,N_8712,N_10148);
nor U13077 (N_13077,N_8265,N_12120);
and U13078 (N_13078,N_6906,N_12219);
or U13079 (N_13079,N_9228,N_10499);
and U13080 (N_13080,N_9776,N_11928);
nand U13081 (N_13081,N_10618,N_11615);
or U13082 (N_13082,N_8689,N_10479);
nand U13083 (N_13083,N_11847,N_8055);
nand U13084 (N_13084,N_8658,N_6588);
nand U13085 (N_13085,N_8580,N_10585);
or U13086 (N_13086,N_11340,N_7384);
nand U13087 (N_13087,N_8073,N_8988);
and U13088 (N_13088,N_7198,N_10487);
nor U13089 (N_13089,N_11409,N_8923);
nor U13090 (N_13090,N_10897,N_10760);
nor U13091 (N_13091,N_7383,N_10740);
and U13092 (N_13092,N_9804,N_11821);
and U13093 (N_13093,N_9762,N_11765);
or U13094 (N_13094,N_12230,N_11652);
nand U13095 (N_13095,N_9013,N_10831);
nand U13096 (N_13096,N_7774,N_10927);
nor U13097 (N_13097,N_8710,N_6762);
nor U13098 (N_13098,N_6591,N_8130);
nand U13099 (N_13099,N_11355,N_7222);
nand U13100 (N_13100,N_10871,N_12382);
or U13101 (N_13101,N_9276,N_7681);
nand U13102 (N_13102,N_10748,N_10800);
or U13103 (N_13103,N_11321,N_12333);
nor U13104 (N_13104,N_6891,N_7662);
nand U13105 (N_13105,N_11421,N_9497);
or U13106 (N_13106,N_7348,N_9479);
nor U13107 (N_13107,N_7007,N_10501);
nand U13108 (N_13108,N_6854,N_8892);
nor U13109 (N_13109,N_7962,N_8694);
or U13110 (N_13110,N_7431,N_7670);
and U13111 (N_13111,N_6479,N_6492);
nand U13112 (N_13112,N_12482,N_8083);
nor U13113 (N_13113,N_8263,N_6896);
or U13114 (N_13114,N_8072,N_9682);
nand U13115 (N_13115,N_11915,N_7203);
nor U13116 (N_13116,N_8426,N_12004);
or U13117 (N_13117,N_11452,N_11448);
or U13118 (N_13118,N_6571,N_9281);
or U13119 (N_13119,N_10284,N_7418);
nor U13120 (N_13120,N_12093,N_12248);
nand U13121 (N_13121,N_8102,N_8879);
or U13122 (N_13122,N_12157,N_8877);
nand U13123 (N_13123,N_7889,N_9137);
nand U13124 (N_13124,N_8070,N_6799);
and U13125 (N_13125,N_11306,N_8463);
nand U13126 (N_13126,N_10223,N_10280);
and U13127 (N_13127,N_7715,N_6901);
xnor U13128 (N_13128,N_8223,N_7239);
nor U13129 (N_13129,N_8764,N_7861);
or U13130 (N_13130,N_7169,N_8648);
nor U13131 (N_13131,N_11733,N_9946);
nand U13132 (N_13132,N_11006,N_11869);
and U13133 (N_13133,N_10156,N_9959);
and U13134 (N_13134,N_6989,N_10449);
nor U13135 (N_13135,N_12064,N_6404);
nor U13136 (N_13136,N_9530,N_9556);
or U13137 (N_13137,N_6673,N_9780);
or U13138 (N_13138,N_6655,N_9268);
or U13139 (N_13139,N_10598,N_10275);
nor U13140 (N_13140,N_7870,N_8697);
nand U13141 (N_13141,N_8549,N_6839);
or U13142 (N_13142,N_10084,N_12477);
and U13143 (N_13143,N_8834,N_6900);
and U13144 (N_13144,N_10602,N_8051);
or U13145 (N_13145,N_8377,N_12009);
nor U13146 (N_13146,N_10955,N_11958);
nor U13147 (N_13147,N_9672,N_8860);
nand U13148 (N_13148,N_9562,N_7742);
and U13149 (N_13149,N_11642,N_6963);
nor U13150 (N_13150,N_10545,N_10824);
nor U13151 (N_13151,N_10779,N_9802);
nor U13152 (N_13152,N_9062,N_12014);
or U13153 (N_13153,N_9271,N_7912);
nor U13154 (N_13154,N_9343,N_12023);
nand U13155 (N_13155,N_8023,N_7267);
nor U13156 (N_13156,N_7777,N_6726);
nor U13157 (N_13157,N_8271,N_7148);
nand U13158 (N_13158,N_9355,N_10933);
or U13159 (N_13159,N_6568,N_9600);
nand U13160 (N_13160,N_11407,N_7337);
nor U13161 (N_13161,N_9280,N_6748);
and U13162 (N_13162,N_6968,N_11161);
nor U13163 (N_13163,N_8960,N_9819);
nor U13164 (N_13164,N_9964,N_10303);
or U13165 (N_13165,N_7424,N_8316);
and U13166 (N_13166,N_8415,N_10864);
nor U13167 (N_13167,N_8462,N_10863);
or U13168 (N_13168,N_10508,N_9777);
and U13169 (N_13169,N_9504,N_8683);
nand U13170 (N_13170,N_9239,N_8566);
and U13171 (N_13171,N_11341,N_9734);
nor U13172 (N_13172,N_11129,N_11222);
and U13173 (N_13173,N_9362,N_9982);
nor U13174 (N_13174,N_10577,N_9618);
and U13175 (N_13175,N_9721,N_6764);
or U13176 (N_13176,N_7558,N_10481);
nand U13177 (N_13177,N_6703,N_10815);
and U13178 (N_13178,N_12207,N_10439);
nand U13179 (N_13179,N_11146,N_11577);
or U13180 (N_13180,N_9124,N_6273);
nand U13181 (N_13181,N_11796,N_7094);
nor U13182 (N_13182,N_11054,N_10641);
nor U13183 (N_13183,N_12480,N_9490);
nor U13184 (N_13184,N_8576,N_10912);
or U13185 (N_13185,N_10254,N_11744);
nand U13186 (N_13186,N_8289,N_10935);
nor U13187 (N_13187,N_8432,N_6903);
nand U13188 (N_13188,N_7847,N_10945);
or U13189 (N_13189,N_9371,N_11248);
nand U13190 (N_13190,N_7817,N_11947);
nand U13191 (N_13191,N_10344,N_11289);
nor U13192 (N_13192,N_6941,N_7143);
nor U13193 (N_13193,N_10704,N_12193);
and U13194 (N_13194,N_6489,N_10557);
nor U13195 (N_13195,N_12364,N_6595);
or U13196 (N_13196,N_11525,N_8720);
and U13197 (N_13197,N_7948,N_9428);
nand U13198 (N_13198,N_6636,N_7868);
and U13199 (N_13199,N_11622,N_7464);
and U13200 (N_13200,N_9848,N_8173);
and U13201 (N_13201,N_11911,N_10453);
or U13202 (N_13202,N_10718,N_10233);
and U13203 (N_13203,N_7966,N_11270);
nand U13204 (N_13204,N_12182,N_8920);
nand U13205 (N_13205,N_8203,N_11475);
nor U13206 (N_13206,N_8236,N_6544);
nand U13207 (N_13207,N_12348,N_7468);
nor U13208 (N_13208,N_11004,N_9747);
nand U13209 (N_13209,N_8973,N_9807);
nand U13210 (N_13210,N_8791,N_9796);
nand U13211 (N_13211,N_12397,N_11717);
and U13212 (N_13212,N_9349,N_9096);
and U13213 (N_13213,N_7188,N_9843);
nand U13214 (N_13214,N_11315,N_11632);
or U13215 (N_13215,N_11476,N_8479);
or U13216 (N_13216,N_11508,N_7841);
and U13217 (N_13217,N_6990,N_7265);
nand U13218 (N_13218,N_11587,N_9878);
or U13219 (N_13219,N_10812,N_8245);
nor U13220 (N_13220,N_8246,N_8220);
nor U13221 (N_13221,N_11392,N_10782);
nand U13222 (N_13222,N_11181,N_10112);
or U13223 (N_13223,N_12498,N_6831);
nor U13224 (N_13224,N_7789,N_12017);
or U13225 (N_13225,N_8728,N_8128);
or U13226 (N_13226,N_11109,N_9021);
nor U13227 (N_13227,N_7016,N_9049);
nor U13228 (N_13228,N_9858,N_6320);
and U13229 (N_13229,N_11422,N_10594);
nand U13230 (N_13230,N_10713,N_9168);
and U13231 (N_13231,N_11617,N_9321);
nand U13232 (N_13232,N_10957,N_6657);
and U13233 (N_13233,N_7347,N_10042);
or U13234 (N_13234,N_9047,N_7048);
nor U13235 (N_13235,N_10343,N_12264);
nor U13236 (N_13236,N_8678,N_6274);
nor U13237 (N_13237,N_8346,N_6767);
or U13238 (N_13238,N_9501,N_10787);
nor U13239 (N_13239,N_7731,N_6451);
and U13240 (N_13240,N_12340,N_11896);
and U13241 (N_13241,N_11972,N_12035);
nor U13242 (N_13242,N_12205,N_8559);
and U13243 (N_13243,N_7050,N_7000);
and U13244 (N_13244,N_10158,N_9421);
or U13245 (N_13245,N_11390,N_11172);
and U13246 (N_13246,N_12133,N_7057);
and U13247 (N_13247,N_8750,N_12306);
nor U13248 (N_13248,N_6779,N_6308);
nor U13249 (N_13249,N_12109,N_8630);
and U13250 (N_13250,N_10504,N_6878);
and U13251 (N_13251,N_10631,N_7475);
and U13252 (N_13252,N_11702,N_10369);
nand U13253 (N_13253,N_10650,N_10916);
nand U13254 (N_13254,N_10382,N_8065);
or U13255 (N_13255,N_8830,N_6952);
nor U13256 (N_13256,N_11527,N_8441);
nor U13257 (N_13257,N_10725,N_10518);
and U13258 (N_13258,N_7218,N_9066);
nor U13259 (N_13259,N_9175,N_10689);
or U13260 (N_13260,N_10604,N_8195);
or U13261 (N_13261,N_6795,N_8004);
or U13262 (N_13262,N_9788,N_10967);
and U13263 (N_13263,N_7192,N_8790);
and U13264 (N_13264,N_6971,N_6372);
nand U13265 (N_13265,N_6785,N_11817);
nand U13266 (N_13266,N_11099,N_9893);
and U13267 (N_13267,N_10817,N_7572);
or U13268 (N_13268,N_12426,N_12265);
nor U13269 (N_13269,N_9292,N_8053);
nor U13270 (N_13270,N_12429,N_7311);
or U13271 (N_13271,N_12172,N_9472);
or U13272 (N_13272,N_9499,N_7790);
and U13273 (N_13273,N_6348,N_12284);
nand U13274 (N_13274,N_12164,N_7119);
nand U13275 (N_13275,N_8866,N_7839);
and U13276 (N_13276,N_12076,N_8748);
nor U13277 (N_13277,N_8650,N_9329);
nand U13278 (N_13278,N_9753,N_7196);
or U13279 (N_13279,N_12489,N_6586);
nand U13280 (N_13280,N_9715,N_10122);
and U13281 (N_13281,N_11588,N_6583);
xor U13282 (N_13282,N_8156,N_11787);
and U13283 (N_13283,N_10491,N_10888);
or U13284 (N_13284,N_9170,N_9941);
nor U13285 (N_13285,N_10029,N_7746);
nand U13286 (N_13286,N_10044,N_8176);
and U13287 (N_13287,N_8793,N_8692);
nor U13288 (N_13288,N_9476,N_9539);
or U13289 (N_13289,N_11661,N_9869);
nor U13290 (N_13290,N_11446,N_12290);
nand U13291 (N_13291,N_11073,N_9778);
nand U13292 (N_13292,N_11317,N_8821);
nor U13293 (N_13293,N_6851,N_10059);
nor U13294 (N_13294,N_12135,N_11909);
nand U13295 (N_13295,N_8480,N_8333);
or U13296 (N_13296,N_10677,N_7985);
nor U13297 (N_13297,N_10739,N_12048);
and U13298 (N_13298,N_9578,N_9470);
nand U13299 (N_13299,N_10415,N_8464);
or U13300 (N_13300,N_12092,N_9783);
nand U13301 (N_13301,N_12222,N_8133);
or U13302 (N_13302,N_11879,N_10017);
or U13303 (N_13303,N_8302,N_9333);
and U13304 (N_13304,N_7211,N_11996);
nand U13305 (N_13305,N_8869,N_8569);
and U13306 (N_13306,N_11871,N_12334);
and U13307 (N_13307,N_10129,N_6353);
nand U13308 (N_13308,N_7367,N_8639);
nand U13309 (N_13309,N_10133,N_9656);
or U13310 (N_13310,N_7676,N_7387);
and U13311 (N_13311,N_10333,N_7600);
nor U13312 (N_13312,N_8529,N_7026);
nor U13313 (N_13313,N_12289,N_10515);
and U13314 (N_13314,N_8123,N_9398);
nand U13315 (N_13315,N_7828,N_10914);
nor U13316 (N_13316,N_10108,N_10452);
nand U13317 (N_13317,N_10282,N_6377);
nor U13318 (N_13318,N_9820,N_11987);
nand U13319 (N_13319,N_12010,N_9632);
and U13320 (N_13320,N_11403,N_12467);
and U13321 (N_13321,N_11679,N_8288);
nor U13322 (N_13322,N_8690,N_9097);
and U13323 (N_13323,N_8617,N_11558);
or U13324 (N_13324,N_9258,N_10248);
and U13325 (N_13325,N_10419,N_6876);
xor U13326 (N_13326,N_11274,N_6649);
and U13327 (N_13327,N_11444,N_7377);
nand U13328 (N_13328,N_12446,N_10672);
nor U13329 (N_13329,N_9131,N_11727);
nor U13330 (N_13330,N_10021,N_9020);
nor U13331 (N_13331,N_10985,N_8522);
or U13332 (N_13332,N_8235,N_9075);
or U13333 (N_13333,N_12438,N_6378);
and U13334 (N_13334,N_8902,N_11299);
or U13335 (N_13335,N_8942,N_9216);
or U13336 (N_13336,N_7498,N_6986);
and U13337 (N_13337,N_9221,N_10743);
nor U13338 (N_13338,N_7151,N_11556);
and U13339 (N_13339,N_7304,N_8674);
or U13340 (N_13340,N_7954,N_8874);
nand U13341 (N_13341,N_10232,N_10488);
nand U13342 (N_13342,N_10000,N_9002);
and U13343 (N_13343,N_6719,N_9553);
or U13344 (N_13344,N_9173,N_11964);
or U13345 (N_13345,N_6603,N_10540);
and U13346 (N_13346,N_9375,N_9099);
or U13347 (N_13347,N_12147,N_7836);
nand U13348 (N_13348,N_8987,N_6553);
nand U13349 (N_13349,N_8729,N_7425);
or U13350 (N_13350,N_8676,N_6668);
nor U13351 (N_13351,N_11051,N_11750);
and U13352 (N_13352,N_8472,N_8407);
and U13353 (N_13353,N_8418,N_11375);
or U13354 (N_13354,N_10626,N_6254);
and U13355 (N_13355,N_10267,N_10711);
and U13356 (N_13356,N_6478,N_7469);
or U13357 (N_13357,N_9700,N_11713);
nor U13358 (N_13358,N_11646,N_11369);
or U13359 (N_13359,N_11802,N_11580);
and U13360 (N_13360,N_10189,N_7253);
nor U13361 (N_13361,N_6868,N_8131);
nand U13362 (N_13362,N_12221,N_6409);
or U13363 (N_13363,N_8596,N_12410);
or U13364 (N_13364,N_8890,N_10398);
nand U13365 (N_13365,N_8740,N_9050);
and U13366 (N_13366,N_10901,N_8844);
and U13367 (N_13367,N_9392,N_11437);
nor U13368 (N_13368,N_10159,N_9305);
nor U13369 (N_13369,N_8500,N_9314);
nand U13370 (N_13370,N_7865,N_7578);
or U13371 (N_13371,N_12212,N_10167);
nand U13372 (N_13372,N_11544,N_8809);
or U13373 (N_13373,N_6944,N_12319);
xor U13374 (N_13374,N_12170,N_11250);
nand U13375 (N_13375,N_7002,N_6627);
and U13376 (N_13376,N_10265,N_8947);
nand U13377 (N_13377,N_12339,N_8071);
xnor U13378 (N_13378,N_8624,N_10990);
and U13379 (N_13379,N_8546,N_10783);
nor U13380 (N_13380,N_8455,N_7160);
nand U13381 (N_13381,N_8213,N_8544);
or U13382 (N_13382,N_8557,N_10328);
nor U13383 (N_13383,N_9694,N_12108);
or U13384 (N_13384,N_6964,N_6548);
nand U13385 (N_13385,N_7710,N_11371);
nand U13386 (N_13386,N_12355,N_8889);
nor U13387 (N_13387,N_10651,N_9636);
nor U13388 (N_13388,N_10561,N_7812);
and U13389 (N_13389,N_9303,N_7135);
nor U13390 (N_13390,N_7179,N_10944);
or U13391 (N_13391,N_9525,N_8855);
nand U13392 (N_13392,N_10011,N_8115);
xor U13393 (N_13393,N_11123,N_6577);
nor U13394 (N_13394,N_10771,N_9467);
nand U13395 (N_13395,N_7527,N_11429);
nand U13396 (N_13396,N_11705,N_6390);
or U13397 (N_13397,N_10706,N_7022);
nand U13398 (N_13398,N_6757,N_12370);
nor U13399 (N_13399,N_9528,N_10271);
nor U13400 (N_13400,N_9174,N_9996);
nand U13401 (N_13401,N_6609,N_11856);
or U13402 (N_13402,N_8137,N_9862);
or U13403 (N_13403,N_9500,N_12199);
and U13404 (N_13404,N_8338,N_8368);
nand U13405 (N_13405,N_6979,N_12286);
nand U13406 (N_13406,N_6836,N_10952);
or U13407 (N_13407,N_8575,N_7428);
nand U13408 (N_13408,N_7349,N_7293);
nand U13409 (N_13409,N_11706,N_7523);
or U13410 (N_13410,N_10200,N_6380);
nand U13411 (N_13411,N_8404,N_11132);
or U13412 (N_13412,N_9357,N_11548);
or U13413 (N_13413,N_7688,N_10025);
or U13414 (N_13414,N_11704,N_11907);
or U13415 (N_13415,N_11157,N_10822);
nor U13416 (N_13416,N_11464,N_11142);
nand U13417 (N_13417,N_7797,N_9064);
or U13418 (N_13418,N_12079,N_8706);
nand U13419 (N_13419,N_10946,N_9048);
nor U13420 (N_13420,N_10140,N_7986);
nor U13421 (N_13421,N_10873,N_9965);
and U13422 (N_13422,N_8801,N_8820);
nand U13423 (N_13423,N_11942,N_6398);
or U13424 (N_13424,N_12385,N_10693);
and U13425 (N_13425,N_10236,N_6333);
or U13426 (N_13426,N_6965,N_11243);
nand U13427 (N_13427,N_10414,N_12431);
nor U13428 (N_13428,N_7381,N_9710);
nor U13429 (N_13429,N_7419,N_7312);
nor U13430 (N_13430,N_6626,N_10128);
or U13431 (N_13431,N_11275,N_10318);
nor U13432 (N_13432,N_6942,N_7375);
nor U13433 (N_13433,N_8665,N_7368);
nor U13434 (N_13434,N_10107,N_7555);
nor U13435 (N_13435,N_9028,N_10310);
or U13436 (N_13436,N_7827,N_9707);
nor U13437 (N_13437,N_12151,N_7971);
or U13438 (N_13438,N_6679,N_6738);
or U13439 (N_13439,N_6518,N_10995);
nand U13440 (N_13440,N_6543,N_10172);
nand U13441 (N_13441,N_7882,N_10171);
nand U13442 (N_13442,N_11982,N_11728);
and U13443 (N_13443,N_7202,N_11191);
or U13444 (N_13444,N_8543,N_9234);
or U13445 (N_13445,N_11913,N_6869);
nor U13446 (N_13446,N_10750,N_6732);
nand U13447 (N_13447,N_12436,N_7060);
nand U13448 (N_13448,N_10884,N_6961);
or U13449 (N_13449,N_6670,N_10920);
nand U13450 (N_13450,N_6415,N_9369);
nor U13451 (N_13451,N_8919,N_9902);
nand U13452 (N_13452,N_7978,N_11040);
and U13453 (N_13453,N_10436,N_9942);
nor U13454 (N_13454,N_7518,N_8166);
and U13455 (N_13455,N_9269,N_12237);
nand U13456 (N_13456,N_9243,N_8274);
nor U13457 (N_13457,N_9812,N_6326);
nor U13458 (N_13458,N_9891,N_10909);
or U13459 (N_13459,N_7825,N_8562);
nor U13460 (N_13460,N_9803,N_6493);
or U13461 (N_13461,N_11926,N_7941);
or U13462 (N_13462,N_7584,N_7583);
and U13463 (N_13463,N_10579,N_6754);
and U13464 (N_13464,N_6858,N_11350);
nor U13465 (N_13465,N_6671,N_11701);
nor U13466 (N_13466,N_7738,N_7703);
nand U13467 (N_13467,N_6521,N_10671);
or U13468 (N_13468,N_10921,N_12213);
and U13469 (N_13469,N_7709,N_10351);
nand U13470 (N_13470,N_7904,N_10255);
nor U13471 (N_13471,N_11203,N_12442);
nand U13472 (N_13472,N_11861,N_9609);
and U13473 (N_13473,N_8181,N_8204);
and U13474 (N_13474,N_9425,N_11168);
or U13475 (N_13475,N_7727,N_7147);
nor U13476 (N_13476,N_7732,N_8272);
and U13477 (N_13477,N_9290,N_11685);
nand U13478 (N_13478,N_12056,N_10931);
nor U13479 (N_13479,N_7003,N_6344);
or U13480 (N_13480,N_9975,N_11829);
nand U13481 (N_13481,N_10161,N_10507);
and U13482 (N_13482,N_8847,N_10919);
or U13483 (N_13483,N_8661,N_10426);
and U13484 (N_13484,N_8074,N_10418);
nor U13485 (N_13485,N_8913,N_12050);
nand U13486 (N_13486,N_8420,N_8530);
and U13487 (N_13487,N_6482,N_6472);
and U13488 (N_13488,N_10981,N_9877);
nor U13489 (N_13489,N_7001,N_6594);
nand U13490 (N_13490,N_6267,N_9827);
or U13491 (N_13491,N_10792,N_10018);
nand U13492 (N_13492,N_9974,N_8286);
nand U13493 (N_13493,N_6563,N_6259);
and U13494 (N_13494,N_9367,N_7142);
or U13495 (N_13495,N_6403,N_7113);
nand U13496 (N_13496,N_11131,N_7549);
and U13497 (N_13497,N_9488,N_11106);
and U13498 (N_13498,N_11304,N_10807);
nand U13499 (N_13499,N_10533,N_6801);
nand U13500 (N_13500,N_6406,N_10575);
nor U13501 (N_13501,N_11894,N_7215);
nand U13502 (N_13502,N_12283,N_10891);
or U13503 (N_13503,N_9386,N_12227);
or U13504 (N_13504,N_11546,N_7559);
and U13505 (N_13505,N_7934,N_8822);
nand U13506 (N_13506,N_9238,N_10917);
and U13507 (N_13507,N_12069,N_11654);
nand U13508 (N_13508,N_7663,N_8266);
nor U13509 (N_13509,N_11288,N_7366);
xnor U13510 (N_13510,N_11185,N_9719);
or U13511 (N_13511,N_10988,N_10076);
nand U13512 (N_13512,N_9213,N_6709);
nor U13513 (N_13513,N_7213,N_7563);
and U13514 (N_13514,N_7472,N_9638);
nand U13515 (N_13515,N_7183,N_9001);
or U13516 (N_13516,N_11367,N_6866);
nor U13517 (N_13517,N_6542,N_6638);
nand U13518 (N_13518,N_9445,N_11995);
nor U13519 (N_13519,N_11026,N_6540);
or U13520 (N_13520,N_8961,N_11910);
nand U13521 (N_13521,N_12209,N_9928);
nand U13522 (N_13522,N_7752,N_11844);
and U13523 (N_13523,N_8555,N_11534);
nand U13524 (N_13524,N_7020,N_12287);
or U13525 (N_13525,N_8589,N_10716);
nor U13526 (N_13526,N_6811,N_7407);
or U13527 (N_13527,N_12200,N_9738);
and U13528 (N_13528,N_6881,N_7463);
or U13529 (N_13529,N_7376,N_6580);
and U13530 (N_13530,N_7509,N_6407);
nand U13531 (N_13531,N_9953,N_10932);
nor U13532 (N_13532,N_10629,N_11711);
nor U13533 (N_13533,N_10389,N_7785);
and U13534 (N_13534,N_7901,N_6557);
and U13535 (N_13535,N_9599,N_6608);
or U13536 (N_13536,N_11223,N_10249);
or U13537 (N_13537,N_9112,N_11889);
nand U13538 (N_13538,N_12251,N_9481);
and U13539 (N_13539,N_7098,N_12437);
or U13540 (N_13540,N_8651,N_9592);
and U13541 (N_13541,N_10227,N_12054);
nor U13542 (N_13542,N_12176,N_11090);
nand U13543 (N_13543,N_8846,N_10700);
or U13544 (N_13544,N_7434,N_11563);
and U13545 (N_13545,N_6391,N_6987);
nand U13546 (N_13546,N_11723,N_11505);
nand U13547 (N_13547,N_7438,N_10853);
nand U13548 (N_13548,N_11455,N_7520);
and U13549 (N_13549,N_6725,N_7880);
nand U13550 (N_13550,N_11551,N_8468);
nor U13551 (N_13551,N_6573,N_7853);
nor U13552 (N_13552,N_9844,N_12258);
and U13553 (N_13553,N_12360,N_9039);
nor U13554 (N_13554,N_8573,N_8411);
nor U13555 (N_13555,N_9736,N_10584);
or U13556 (N_13556,N_6257,N_8662);
nor U13557 (N_13557,N_11667,N_6911);
and U13558 (N_13558,N_8049,N_10855);
or U13559 (N_13559,N_8968,N_7182);
or U13560 (N_13560,N_7459,N_10093);
or U13561 (N_13561,N_8798,N_7965);
nand U13562 (N_13562,N_10198,N_9109);
and U13563 (N_13563,N_12448,N_11756);
nor U13564 (N_13564,N_10329,N_12211);
and U13565 (N_13565,N_7402,N_9735);
nand U13566 (N_13566,N_9534,N_6723);
and U13567 (N_13567,N_12393,N_11137);
nand U13568 (N_13568,N_12039,N_7819);
and U13569 (N_13569,N_7373,N_11781);
nand U13570 (N_13570,N_6632,N_10754);
and U13571 (N_13571,N_9969,N_11956);
or U13572 (N_13572,N_7364,N_9419);
nor U13573 (N_13573,N_8827,N_11399);
nand U13574 (N_13574,N_11083,N_7834);
nand U13575 (N_13575,N_6395,N_6938);
and U13576 (N_13576,N_8908,N_8193);
nor U13577 (N_13577,N_6528,N_10899);
nor U13578 (N_13578,N_11698,N_8517);
and U13579 (N_13579,N_10489,N_11227);
or U13580 (N_13580,N_8741,N_9791);
or U13581 (N_13581,N_9265,N_10837);
nand U13582 (N_13582,N_9198,N_10789);
and U13583 (N_13583,N_10620,N_8242);
nor U13584 (N_13584,N_10326,N_8578);
and U13585 (N_13585,N_12008,N_12254);
and U13586 (N_13586,N_9240,N_12231);
and U13587 (N_13587,N_11118,N_10073);
or U13588 (N_13588,N_8296,N_10865);
or U13589 (N_13589,N_9331,N_11753);
or U13590 (N_13590,N_8757,N_7979);
nand U13591 (N_13591,N_11439,N_10183);
nor U13592 (N_13592,N_7163,N_7201);
or U13593 (N_13593,N_10699,N_9084);
nor U13594 (N_13594,N_10468,N_6310);
and U13595 (N_13595,N_6660,N_6937);
and U13596 (N_13596,N_11128,N_8932);
or U13597 (N_13597,N_6357,N_9263);
or U13598 (N_13598,N_9035,N_12112);
nand U13599 (N_13599,N_7320,N_9794);
and U13600 (N_13600,N_8144,N_6863);
or U13601 (N_13601,N_7740,N_6702);
nor U13602 (N_13602,N_10169,N_6782);
nor U13603 (N_13603,N_10462,N_6682);
nor U13604 (N_13604,N_6992,N_8216);
and U13605 (N_13605,N_8794,N_12291);
nand U13606 (N_13606,N_6418,N_7792);
or U13607 (N_13607,N_9352,N_6606);
or U13608 (N_13608,N_10751,N_7756);
or U13609 (N_13609,N_10842,N_8322);
nand U13610 (N_13610,N_9192,N_9076);
nand U13611 (N_13611,N_11842,N_6473);
or U13612 (N_13612,N_8560,N_6718);
nor U13613 (N_13613,N_6864,N_10562);
nor U13614 (N_13614,N_11724,N_7791);
nor U13615 (N_13615,N_9961,N_10296);
nor U13616 (N_13616,N_11870,N_9090);
nand U13617 (N_13617,N_11470,N_11405);
nand U13618 (N_13618,N_10411,N_11404);
and U13619 (N_13619,N_10478,N_8917);
or U13620 (N_13620,N_11133,N_7435);
nor U13621 (N_13621,N_11951,N_6651);
or U13622 (N_13622,N_7983,N_9899);
and U13623 (N_13623,N_9998,N_11927);
nor U13624 (N_13624,N_7939,N_7205);
nor U13625 (N_13625,N_10277,N_11716);
or U13626 (N_13626,N_11990,N_11370);
nand U13627 (N_13627,N_9370,N_9709);
and U13628 (N_13628,N_10978,N_7943);
nand U13629 (N_13629,N_8136,N_7682);
and U13630 (N_13630,N_12143,N_11573);
and U13631 (N_13631,N_8572,N_7894);
and U13632 (N_13632,N_11812,N_10312);
nor U13633 (N_13633,N_9247,N_9406);
nand U13634 (N_13634,N_6258,N_11616);
nor U13635 (N_13635,N_9311,N_8077);
or U13636 (N_13636,N_8214,N_6662);
or U13637 (N_13637,N_6537,N_9784);
or U13638 (N_13638,N_8670,N_12337);
nand U13639 (N_13639,N_11328,N_7616);
or U13640 (N_13640,N_12273,N_11254);
nor U13641 (N_13641,N_8797,N_9611);
and U13642 (N_13642,N_10114,N_8000);
nand U13643 (N_13643,N_6658,N_8244);
and U13644 (N_13644,N_9704,N_7388);
or U13645 (N_13645,N_7718,N_8103);
or U13646 (N_13646,N_8371,N_6323);
nand U13647 (N_13647,N_9950,N_10764);
and U13648 (N_13648,N_8905,N_8561);
and U13649 (N_13649,N_10622,N_11811);
nand U13650 (N_13650,N_10976,N_10247);
nor U13651 (N_13651,N_8406,N_6260);
nor U13652 (N_13652,N_12021,N_12136);
nor U13653 (N_13653,N_11522,N_8945);
or U13654 (N_13654,N_7486,N_11398);
nand U13655 (N_13655,N_7324,N_9384);
xor U13656 (N_13656,N_8267,N_7243);
or U13657 (N_13657,N_7744,N_6411);
and U13658 (N_13658,N_10965,N_12366);
nor U13659 (N_13659,N_9929,N_10015);
and U13660 (N_13660,N_10321,N_11246);
nand U13661 (N_13661,N_11535,N_6432);
nand U13662 (N_13662,N_10749,N_11521);
and U13663 (N_13663,N_11893,N_10053);
nand U13664 (N_13664,N_10288,N_11273);
and U13665 (N_13665,N_11513,N_6530);
nand U13666 (N_13666,N_11953,N_9602);
or U13667 (N_13667,N_10199,N_8671);
nor U13668 (N_13668,N_11219,N_8185);
nor U13669 (N_13669,N_11325,N_12332);
or U13670 (N_13670,N_12089,N_11329);
and U13671 (N_13671,N_7820,N_8867);
or U13672 (N_13672,N_10020,N_10056);
nand U13673 (N_13673,N_9298,N_11860);
nand U13674 (N_13674,N_8641,N_9919);
nor U13675 (N_13675,N_9098,N_11053);
nor U13676 (N_13676,N_7503,N_6551);
nor U13677 (N_13677,N_6771,N_7391);
or U13678 (N_13678,N_12313,N_7784);
nor U13679 (N_13679,N_11145,N_6787);
nand U13680 (N_13680,N_7672,N_9988);
and U13681 (N_13681,N_11639,N_12066);
or U13682 (N_13682,N_9692,N_8345);
or U13683 (N_13683,N_11612,N_8512);
or U13684 (N_13684,N_8219,N_11175);
nor U13685 (N_13685,N_7885,N_9199);
and U13686 (N_13686,N_7115,N_9432);
or U13687 (N_13687,N_10366,N_7180);
and U13688 (N_13688,N_8620,N_9927);
and U13689 (N_13689,N_8819,N_8297);
nand U13690 (N_13690,N_10202,N_10907);
nor U13691 (N_13691,N_8202,N_10096);
or U13692 (N_13692,N_8534,N_11515);
nand U13693 (N_13693,N_6319,N_10103);
nand U13694 (N_13694,N_7635,N_11255);
or U13695 (N_13695,N_7745,N_11018);
nor U13696 (N_13696,N_12027,N_7220);
nand U13697 (N_13697,N_10875,N_9821);
and U13698 (N_13698,N_11135,N_6434);
and U13699 (N_13699,N_7398,N_10780);
or U13700 (N_13700,N_6793,N_9337);
or U13701 (N_13701,N_11600,N_7207);
and U13702 (N_13702,N_6893,N_10120);
nor U13703 (N_13703,N_7956,N_7018);
and U13704 (N_13704,N_11000,N_10829);
or U13705 (N_13705,N_8893,N_11737);
and U13706 (N_13706,N_12317,N_12028);
nand U13707 (N_13707,N_9897,N_11606);
or U13708 (N_13708,N_6321,N_11578);
or U13709 (N_13709,N_8520,N_9195);
nor U13710 (N_13710,N_6800,N_6823);
and U13711 (N_13711,N_10472,N_10371);
nand U13712 (N_13712,N_6433,N_9161);
nor U13713 (N_13713,N_7261,N_7833);
and U13714 (N_13714,N_8483,N_10925);
nand U13715 (N_13715,N_6920,N_6419);
or U13716 (N_13716,N_6846,N_10047);
nand U13717 (N_13717,N_6498,N_8667);
or U13718 (N_13718,N_9082,N_9052);
and U13719 (N_13719,N_9920,N_9245);
nand U13720 (N_13720,N_8261,N_7936);
or U13721 (N_13721,N_8786,N_10971);
and U13722 (N_13722,N_9531,N_10753);
nand U13723 (N_13723,N_9277,N_10240);
and U13724 (N_13724,N_12486,N_8998);
or U13725 (N_13725,N_11311,N_12165);
and U13726 (N_13726,N_10335,N_7855);
and U13727 (N_13727,N_7573,N_11978);
nor U13728 (N_13728,N_8158,N_12499);
or U13729 (N_13729,N_8419,N_7567);
nor U13730 (N_13730,N_11634,N_6840);
and U13731 (N_13731,N_8966,N_10476);
nand U13732 (N_13732,N_9514,N_7533);
or U13733 (N_13733,N_7717,N_7597);
nor U13734 (N_13734,N_9703,N_10221);
nand U13735 (N_13735,N_8117,N_6848);
or U13736 (N_13736,N_9887,N_7726);
nor U13737 (N_13737,N_6804,N_8622);
nor U13738 (N_13738,N_7484,N_12375);
or U13739 (N_13739,N_11778,N_9206);
nand U13740 (N_13740,N_9270,N_12068);
nor U13741 (N_13741,N_10825,N_10635);
and U13742 (N_13742,N_11741,N_11853);
nor U13743 (N_13743,N_7692,N_6991);
nor U13744 (N_13744,N_7128,N_9995);
nand U13745 (N_13745,N_10034,N_8036);
nand U13746 (N_13746,N_8466,N_11759);
or U13747 (N_13747,N_6366,N_11155);
and U13748 (N_13748,N_11799,N_8421);
or U13749 (N_13749,N_11009,N_11900);
nand U13750 (N_13750,N_7276,N_7537);
nor U13751 (N_13751,N_10734,N_11386);
and U13752 (N_13752,N_8744,N_8273);
nand U13753 (N_13753,N_7984,N_10839);
nand U13754 (N_13754,N_7185,N_11207);
or U13755 (N_13755,N_9541,N_8303);
nor U13756 (N_13756,N_11604,N_12439);
nand U13757 (N_13757,N_6427,N_8554);
and U13758 (N_13758,N_7067,N_6291);
nor U13759 (N_13759,N_9720,N_11708);
or U13760 (N_13760,N_8502,N_7305);
nor U13761 (N_13761,N_11674,N_6834);
nand U13762 (N_13762,N_6729,N_8986);
or U13763 (N_13763,N_9759,N_8995);
or U13764 (N_13764,N_11678,N_10139);
nor U13765 (N_13765,N_10195,N_11089);
nor U13766 (N_13766,N_10256,N_10074);
xor U13767 (N_13767,N_8118,N_9380);
nor U13768 (N_13768,N_6784,N_10196);
and U13769 (N_13769,N_8780,N_9092);
nand U13770 (N_13770,N_6324,N_6957);
or U13771 (N_13771,N_10729,N_7725);
or U13772 (N_13772,N_11635,N_7030);
or U13773 (N_13773,N_8755,N_6567);
nor U13774 (N_13774,N_8148,N_8515);
nor U13775 (N_13775,N_12372,N_8397);
and U13776 (N_13776,N_11650,N_10876);
or U13777 (N_13777,N_11641,N_6749);
or U13778 (N_13778,N_11845,N_8279);
or U13779 (N_13779,N_6250,N_8886);
nor U13780 (N_13780,N_7691,N_10461);
nand U13781 (N_13781,N_9267,N_7189);
and U13782 (N_13782,N_6449,N_9055);
nor U13783 (N_13783,N_6661,N_11360);
and U13784 (N_13784,N_8132,N_12158);
nand U13785 (N_13785,N_12373,N_10214);
or U13786 (N_13786,N_10208,N_8495);
nand U13787 (N_13787,N_6822,N_12198);
nor U13788 (N_13788,N_10445,N_8110);
or U13789 (N_13789,N_7483,N_7519);
nand U13790 (N_13790,N_11326,N_6420);
nor U13791 (N_13791,N_8433,N_7386);
nand U13792 (N_13792,N_6816,N_9415);
nand U13793 (N_13793,N_10217,N_9351);
nand U13794 (N_13794,N_10979,N_11598);
or U13795 (N_13795,N_12229,N_10038);
and U13796 (N_13796,N_10766,N_12441);
nand U13797 (N_13797,N_10964,N_8459);
and U13798 (N_13798,N_7171,N_7307);
and U13799 (N_13799,N_6693,N_10786);
nor U13800 (N_13800,N_9698,N_9459);
nor U13801 (N_13801,N_8894,N_10104);
and U13802 (N_13802,N_9069,N_8159);
nor U13803 (N_13803,N_11022,N_11618);
and U13804 (N_13804,N_8605,N_10658);
nor U13805 (N_13805,N_11983,N_9933);
nand U13806 (N_13806,N_10268,N_8301);
or U13807 (N_13807,N_6355,N_7077);
and U13808 (N_13808,N_10611,N_8446);
and U13809 (N_13809,N_11013,N_12419);
nand U13810 (N_13810,N_11206,N_6974);
nand U13811 (N_13811,N_9151,N_8290);
nand U13812 (N_13812,N_7580,N_6379);
or U13813 (N_13813,N_10603,N_6416);
nand U13814 (N_13814,N_11482,N_7083);
and U13815 (N_13815,N_11766,N_11790);
nor U13816 (N_13816,N_9077,N_8594);
nand U13817 (N_13817,N_6533,N_12404);
and U13818 (N_13818,N_11627,N_11314);
nor U13819 (N_13819,N_7476,N_7913);
and U13820 (N_13820,N_9873,N_10520);
and U13821 (N_13821,N_12262,N_12073);
or U13822 (N_13822,N_9829,N_8567);
nand U13823 (N_13823,N_10573,N_8328);
nor U13824 (N_13824,N_11516,N_11917);
and U13825 (N_13825,N_11686,N_12255);
and U13826 (N_13826,N_11782,N_11046);
nand U13827 (N_13827,N_10032,N_11074);
nand U13828 (N_13828,N_11492,N_8336);
nand U13829 (N_13829,N_7421,N_6753);
nor U13830 (N_13830,N_11589,N_6759);
or U13831 (N_13831,N_10688,N_8097);
nand U13832 (N_13832,N_8240,N_9503);
nor U13833 (N_13833,N_11062,N_10773);
nand U13834 (N_13834,N_7086,N_6808);
nand U13835 (N_13835,N_8868,N_7152);
nand U13836 (N_13836,N_11457,N_8876);
nor U13837 (N_13837,N_7636,N_10531);
or U13838 (N_13838,N_12070,N_8001);
and U13839 (N_13839,N_8518,N_8022);
nor U13840 (N_13840,N_9291,N_7322);
nor U13841 (N_13841,N_8066,N_8911);
nor U13842 (N_13842,N_6359,N_9983);
nor U13843 (N_13843,N_10991,N_10163);
nor U13844 (N_13844,N_6465,N_10647);
nand U13845 (N_13845,N_11210,N_9978);
and U13846 (N_13846,N_6913,N_8249);
nor U13847 (N_13847,N_7333,N_7244);
or U13848 (N_13848,N_11594,N_9795);
or U13849 (N_13849,N_8675,N_12342);
xor U13850 (N_13850,N_7711,N_11264);
nor U13851 (N_13851,N_11828,N_8060);
and U13852 (N_13852,N_12458,N_6737);
nand U13853 (N_13853,N_11579,N_9960);
nor U13854 (N_13854,N_11019,N_9513);
nor U13855 (N_13855,N_11974,N_6780);
nor U13856 (N_13856,N_7830,N_8366);
nand U13857 (N_13857,N_8101,N_12485);
nand U13858 (N_13858,N_6750,N_10145);
nor U13859 (N_13859,N_6912,N_7757);
nor U13860 (N_13860,N_9065,N_12369);
or U13861 (N_13861,N_11607,N_8682);
nor U13862 (N_13862,N_9125,N_7874);
and U13863 (N_13863,N_11383,N_11888);
nand U13864 (N_13864,N_10215,N_7078);
nor U13865 (N_13865,N_11629,N_7675);
and U13866 (N_13866,N_11876,N_11117);
nor U13867 (N_13867,N_11703,N_11624);
and U13868 (N_13868,N_7569,N_7915);
or U13869 (N_13869,N_6922,N_9158);
or U13870 (N_13870,N_8196,N_8393);
or U13871 (N_13871,N_10922,N_9117);
nor U13872 (N_13872,N_11055,N_6774);
nand U13873 (N_13873,N_8521,N_10193);
and U13874 (N_13874,N_11481,N_8638);
nand U13875 (N_13875,N_12117,N_11017);
nor U13876 (N_13876,N_9973,N_7102);
nand U13877 (N_13877,N_6488,N_10784);
and U13878 (N_13878,N_6279,N_9727);
nand U13879 (N_13879,N_8783,N_11092);
and U13880 (N_13880,N_9823,N_10816);
or U13881 (N_13881,N_7660,N_10820);
and U13882 (N_13882,N_10266,N_8098);
nor U13883 (N_13883,N_7800,N_6615);
and U13884 (N_13884,N_7251,N_8585);
or U13885 (N_13885,N_6534,N_11564);
or U13886 (N_13886,N_9420,N_6337);
nand U13887 (N_13887,N_7631,N_11143);
nor U13888 (N_13888,N_11919,N_6412);
and U13889 (N_13889,N_7085,N_8907);
and U13890 (N_13890,N_7564,N_10121);
nor U13891 (N_13891,N_9526,N_10458);
nand U13892 (N_13892,N_7562,N_12440);
nor U13893 (N_13893,N_9560,N_7013);
and U13894 (N_13894,N_11536,N_7252);
nor U13895 (N_13895,N_7209,N_7130);
or U13896 (N_13896,N_12038,N_7485);
nor U13897 (N_13897,N_11228,N_11194);
xor U13898 (N_13898,N_11419,N_6928);
nand U13899 (N_13899,N_6776,N_9842);
nor U13900 (N_13900,N_9115,N_7852);
or U13901 (N_13901,N_7092,N_9387);
or U13902 (N_13902,N_12173,N_9860);
nor U13903 (N_13903,N_8443,N_9696);
nand U13904 (N_13904,N_12285,N_9233);
or U13905 (N_13905,N_11554,N_10224);
or U13906 (N_13906,N_6328,N_10334);
or U13907 (N_13907,N_11485,N_11843);
and U13908 (N_13908,N_11835,N_8696);
or U13909 (N_13909,N_10546,N_11029);
nand U13910 (N_13910,N_10251,N_7886);
or U13911 (N_13911,N_9287,N_11783);
or U13912 (N_13912,N_10464,N_7231);
or U13913 (N_13913,N_7980,N_6350);
or U13914 (N_13914,N_8880,N_9991);
nor U13915 (N_13915,N_7859,N_9219);
nor U13916 (N_13916,N_6531,N_12280);
or U13917 (N_13917,N_11127,N_11283);
or U13918 (N_13918,N_11722,N_9197);
nand U13919 (N_13919,N_9516,N_9976);
or U13920 (N_13920,N_11784,N_9454);
or U13921 (N_13921,N_6371,N_12122);
nand U13922 (N_13922,N_10497,N_10188);
nor U13923 (N_13923,N_7321,N_10176);
nor U13924 (N_13924,N_7432,N_6696);
and U13925 (N_13925,N_6462,N_10490);
nand U13926 (N_13926,N_7611,N_7101);
nand U13927 (N_13927,N_8737,N_8681);
and U13928 (N_13928,N_6664,N_6717);
nor U13929 (N_13929,N_6597,N_9766);
and U13930 (N_13930,N_9046,N_9482);
nand U13931 (N_13931,N_9519,N_8175);
nand U13932 (N_13932,N_7011,N_6424);
and U13933 (N_13933,N_8149,N_10660);
and U13934 (N_13934,N_10027,N_7741);
or U13935 (N_13935,N_7702,N_9139);
or U13936 (N_13936,N_12140,N_9839);
or U13937 (N_13937,N_12077,N_8370);
nand U13938 (N_13938,N_8453,N_10506);
and U13939 (N_13939,N_10940,N_10683);
or U13940 (N_13940,N_11929,N_8990);
or U13941 (N_13941,N_10403,N_7494);
or U13942 (N_13942,N_6263,N_9011);
or U13943 (N_13943,N_6295,N_7689);
nand U13944 (N_13944,N_10563,N_7761);
or U13945 (N_13945,N_8965,N_10399);
nor U13946 (N_13946,N_9693,N_6444);
and U13947 (N_13947,N_7478,N_7361);
or U13948 (N_13948,N_7116,N_11682);
and U13949 (N_13949,N_8570,N_10102);
or U13950 (N_13950,N_9626,N_11731);
nor U13951 (N_13951,N_12302,N_10357);
and U13952 (N_13952,N_10315,N_11072);
nand U13953 (N_13953,N_9958,N_8221);
or U13954 (N_13954,N_9108,N_10954);
and U13955 (N_13955,N_8746,N_9416);
or U13956 (N_13956,N_11774,N_10425);
nand U13957 (N_13957,N_9442,N_10033);
nor U13958 (N_13958,N_10854,N_11819);
and U13959 (N_13959,N_6304,N_7462);
nand U13960 (N_13960,N_10664,N_8194);
nand U13961 (N_13961,N_6904,N_9781);
nor U13962 (N_13962,N_7875,N_11088);
nand U13963 (N_13963,N_9458,N_8306);
or U13964 (N_13964,N_9037,N_9888);
nor U13965 (N_13965,N_7034,N_11761);
nand U13966 (N_13966,N_11066,N_11147);
nand U13967 (N_13967,N_8255,N_9847);
nor U13968 (N_13968,N_10904,N_8953);
nand U13969 (N_13969,N_8396,N_6430);
nand U13970 (N_13970,N_11472,N_8085);
nor U13971 (N_13971,N_10298,N_8251);
or U13972 (N_13972,N_7005,N_10765);
and U13973 (N_13973,N_6327,N_9087);
nand U13974 (N_13974,N_10270,N_8612);
nand U13975 (N_13975,N_8295,N_8026);
or U13976 (N_13976,N_10347,N_8109);
nand U13977 (N_13977,N_7027,N_8568);
xor U13978 (N_13978,N_10320,N_6475);
nor U13979 (N_13979,N_11914,N_6550);
nor U13980 (N_13980,N_12202,N_11253);
nand U13981 (N_13981,N_9009,N_9312);
nand U13982 (N_13982,N_11967,N_10834);
nor U13983 (N_13983,N_7866,N_6692);
and U13984 (N_13984,N_7701,N_7096);
or U13985 (N_13985,N_11868,N_8283);
nand U13986 (N_13986,N_10503,N_12247);
or U13987 (N_13987,N_11352,N_7310);
nor U13988 (N_13988,N_11362,N_8627);
or U13989 (N_13989,N_7257,N_12450);
and U13990 (N_13990,N_6589,N_11901);
nor U13991 (N_13991,N_8163,N_7654);
nor U13992 (N_13992,N_7369,N_8489);
nor U13993 (N_13993,N_11762,N_10586);
or U13994 (N_13994,N_7605,N_7042);
nor U13995 (N_13995,N_9548,N_8976);
nand U13996 (N_13996,N_9225,N_10269);
and U13997 (N_13997,N_6442,N_7619);
or U13998 (N_13998,N_7245,N_8312);
or U13999 (N_13999,N_8058,N_6894);
or U14000 (N_14000,N_9651,N_6443);
nand U14001 (N_14001,N_9811,N_6874);
nor U14002 (N_14002,N_8352,N_11816);
or U14003 (N_14003,N_10117,N_6280);
or U14004 (N_14004,N_10190,N_10627);
or U14005 (N_14005,N_11738,N_10164);
nor U14006 (N_14006,N_12022,N_6566);
nand U14007 (N_14007,N_9181,N_10674);
nor U14008 (N_14008,N_10692,N_7110);
nor U14009 (N_14009,N_10705,N_8975);
and U14010 (N_14010,N_11640,N_6680);
and U14011 (N_14011,N_10606,N_11559);
or U14012 (N_14012,N_6909,N_7303);
and U14013 (N_14013,N_10495,N_9412);
nor U14014 (N_14014,N_7453,N_10847);
and U14015 (N_14015,N_10413,N_10614);
and U14016 (N_14016,N_10378,N_10673);
and U14017 (N_14017,N_8329,N_10131);
nor U14018 (N_14018,N_9461,N_8629);
and U14019 (N_14019,N_9229,N_10527);
or U14020 (N_14020,N_10918,N_11918);
or U14021 (N_14021,N_8318,N_9121);
or U14022 (N_14022,N_8206,N_12049);
and U14023 (N_14023,N_6505,N_8497);
and U14024 (N_14024,N_10717,N_9441);
or U14025 (N_14025,N_10175,N_6939);
nand U14026 (N_14026,N_7414,N_6751);
and U14027 (N_14027,N_6616,N_10377);
nor U14028 (N_14028,N_11801,N_9678);
nand U14029 (N_14029,N_8381,N_11357);
xnor U14030 (N_14030,N_12405,N_6358);
xnor U14031 (N_14031,N_9417,N_12019);
nand U14032 (N_14032,N_10331,N_11001);
or U14033 (N_14033,N_10587,N_9620);
nor U14034 (N_14034,N_11241,N_12277);
or U14035 (N_14035,N_7808,N_8127);
nand U14036 (N_14036,N_9061,N_10134);
nand U14037 (N_14037,N_10278,N_9000);
nand U14038 (N_14038,N_9451,N_7296);
nor U14039 (N_14039,N_10680,N_11795);
nand U14040 (N_14040,N_6339,N_7640);
or U14041 (N_14041,N_12107,N_10623);
nor U14042 (N_14042,N_11095,N_11899);
nand U14043 (N_14043,N_6976,N_11258);
nor U14044 (N_14044,N_8853,N_10639);
and U14045 (N_14045,N_9769,N_11575);
or U14046 (N_14046,N_10528,N_11966);
nand U14047 (N_14047,N_9837,N_9748);
nand U14048 (N_14048,N_10301,N_6650);
and U14049 (N_14049,N_6873,N_10213);
nor U14050 (N_14050,N_12383,N_9861);
nor U14051 (N_14051,N_11056,N_11413);
nor U14052 (N_14052,N_6459,N_12037);
and U14053 (N_14053,N_11130,N_10446);
nor U14054 (N_14054,N_7609,N_8831);
or U14055 (N_14055,N_9785,N_11171);
and U14056 (N_14056,N_6569,N_12413);
nand U14057 (N_14057,N_8030,N_6436);
nor U14058 (N_14058,N_9765,N_10970);
or U14059 (N_14059,N_8291,N_6592);
nor U14060 (N_14060,N_10535,N_11863);
nor U14061 (N_14061,N_10191,N_8927);
xnor U14062 (N_14062,N_7433,N_11081);
nand U14063 (N_14063,N_11344,N_11179);
nor U14064 (N_14064,N_9403,N_12020);
nand U14065 (N_14065,N_11479,N_11235);
and U14066 (N_14066,N_7423,N_9187);
and U14067 (N_14067,N_11748,N_7084);
nand U14068 (N_14068,N_9932,N_9015);
and U14069 (N_14069,N_10286,N_12425);
nand U14070 (N_14070,N_11633,N_6724);
and U14071 (N_14071,N_8078,N_7645);
and U14072 (N_14072,N_11504,N_6556);
or U14073 (N_14073,N_11050,N_11730);
and U14074 (N_14074,N_10285,N_12051);
and U14075 (N_14075,N_8075,N_6535);
and U14076 (N_14076,N_9322,N_6734);
nand U14077 (N_14077,N_7242,N_9041);
nand U14078 (N_14078,N_8647,N_6722);
nor U14079 (N_14079,N_8858,N_9088);
and U14080 (N_14080,N_6312,N_9279);
or U14081 (N_14081,N_10742,N_6562);
and U14082 (N_14082,N_12387,N_8896);
or U14083 (N_14083,N_11934,N_12217);
or U14084 (N_14084,N_7156,N_6517);
or U14085 (N_14085,N_11445,N_11309);
or U14086 (N_14086,N_9667,N_12220);
and U14087 (N_14087,N_11644,N_9918);
nor U14088 (N_14088,N_7873,N_10094);
or U14089 (N_14089,N_8057,N_6261);
nor U14090 (N_14090,N_12408,N_11205);
nand U14091 (N_14091,N_8254,N_11994);
or U14092 (N_14092,N_9453,N_6538);
nand U14093 (N_14093,N_10532,N_12001);
nor U14094 (N_14094,N_12232,N_8950);
or U14095 (N_14095,N_8967,N_8659);
nand U14096 (N_14096,N_9757,N_11743);
nor U14097 (N_14097,N_7379,N_11695);
and U14098 (N_14098,N_8595,N_9864);
nor U14099 (N_14099,N_10941,N_6421);
nor U14100 (N_14100,N_9944,N_10463);
or U14101 (N_14101,N_6276,N_12058);
nor U14102 (N_14102,N_11672,N_8091);
nand U14103 (N_14103,N_6367,N_7794);
nand U14104 (N_14104,N_10118,N_10317);
or U14105 (N_14105,N_6576,N_7976);
or U14106 (N_14106,N_7338,N_7683);
nor U14107 (N_14107,N_7146,N_10596);
or U14108 (N_14108,N_11012,N_12464);
and U14109 (N_14109,N_6958,N_12274);
or U14110 (N_14110,N_9934,N_8284);
nand U14111 (N_14111,N_10811,N_7447);
or U14112 (N_14112,N_12149,N_8964);
nor U14113 (N_14113,N_9597,N_11214);
and U14114 (N_14114,N_9521,N_9250);
and U14115 (N_14115,N_7068,N_6773);
or U14116 (N_14116,N_10762,N_7910);
or U14117 (N_14117,N_7221,N_12346);
and U14118 (N_14118,N_8548,N_12102);
or U14119 (N_14119,N_7762,N_7779);
nor U14120 (N_14120,N_9364,N_11566);
nor U14121 (N_14121,N_9224,N_11712);
nor U14122 (N_14122,N_7651,N_6889);
nand U14123 (N_14123,N_10857,N_12381);
or U14124 (N_14124,N_11596,N_11626);
and U14125 (N_14125,N_9557,N_10819);
nand U14126 (N_14126,N_10100,N_10494);
nor U14127 (N_14127,N_6485,N_7937);
or U14128 (N_14128,N_11425,N_10962);
nand U14129 (N_14129,N_7056,N_8134);
and U14130 (N_14130,N_10953,N_9701);
or U14131 (N_14131,N_10097,N_8565);
or U14132 (N_14132,N_12075,N_10581);
or U14133 (N_14133,N_12189,N_11970);
nor U14134 (N_14134,N_8308,N_11973);
or U14135 (N_14135,N_11507,N_12203);
and U14136 (N_14136,N_11337,N_7051);
or U14137 (N_14137,N_10804,N_10835);
nor U14138 (N_14138,N_6875,N_10654);
and U14139 (N_14139,N_9408,N_12281);
and U14140 (N_14140,N_9462,N_10662);
nor U14141 (N_14141,N_7290,N_7574);
or U14142 (N_14142,N_8738,N_9485);
and U14143 (N_14143,N_7233,N_11196);
nand U14144 (N_14144,N_12316,N_6546);
and U14145 (N_14145,N_10080,N_8715);
nand U14146 (N_14146,N_7154,N_8863);
nor U14147 (N_14147,N_11057,N_6423);
nor U14148 (N_14148,N_10738,N_10314);
xor U14149 (N_14149,N_7751,N_9477);
or U14150 (N_14150,N_10723,N_9489);
or U14151 (N_14151,N_11047,N_6865);
xnor U14152 (N_14152,N_6413,N_11838);
nor U14153 (N_14153,N_8054,N_9129);
and U14154 (N_14154,N_10306,N_7891);
xnor U14155 (N_14155,N_10160,N_6746);
nand U14156 (N_14156,N_8256,N_11822);
or U14157 (N_14157,N_7460,N_10124);
or U14158 (N_14158,N_7064,N_11892);
xnor U14159 (N_14159,N_6802,N_10661);
nor U14160 (N_14160,N_7235,N_7069);
or U14161 (N_14161,N_12320,N_6791);
nor U14162 (N_14162,N_8376,N_9059);
or U14163 (N_14163,N_8247,N_7175);
or U14164 (N_14164,N_7184,N_10048);
nor U14165 (N_14165,N_9943,N_11015);
and U14166 (N_14166,N_10272,N_9533);
nand U14167 (N_14167,N_6659,N_11431);
nor U14168 (N_14168,N_11094,N_10243);
nor U14169 (N_14169,N_8093,N_9085);
and U14170 (N_14170,N_6917,N_10628);
and U14171 (N_14171,N_8649,N_11666);
nor U14172 (N_14172,N_6672,N_7439);
nor U14173 (N_14173,N_7542,N_6727);
nand U14174 (N_14174,N_11308,N_11530);
nand U14175 (N_14175,N_12483,N_9697);
and U14176 (N_14176,N_6666,N_7492);
or U14177 (N_14177,N_6667,N_10485);
nor U14178 (N_14178,N_9045,N_10447);
and U14179 (N_14179,N_8619,N_8487);
nand U14180 (N_14180,N_9072,N_9318);
nor U14181 (N_14181,N_7714,N_8275);
and U14182 (N_14182,N_7626,N_7427);
or U14183 (N_14183,N_8842,N_6933);
and U14184 (N_14184,N_7256,N_7515);
and U14185 (N_14185,N_10046,N_9741);
or U14186 (N_14186,N_6491,N_12100);
nor U14187 (N_14187,N_12305,N_6629);
nor U14188 (N_14188,N_8449,N_9376);
xor U14189 (N_14189,N_6599,N_11669);
nor U14190 (N_14190,N_10519,N_7112);
or U14191 (N_14191,N_8287,N_11365);
nor U14192 (N_14192,N_8835,N_10035);
nor U14193 (N_14193,N_7680,N_9787);
and U14194 (N_14194,N_9435,N_7786);
nor U14195 (N_14195,N_12307,N_9947);
nand U14196 (N_14196,N_9191,N_7946);
nor U14197 (N_14197,N_6798,N_11116);
and U14198 (N_14198,N_9981,N_12154);
or U14199 (N_14199,N_9302,N_10526);
nor U14200 (N_14200,N_7646,N_10898);
nand U14201 (N_14201,N_7975,N_9949);
nand U14202 (N_14202,N_9491,N_7106);
and U14203 (N_14203,N_9336,N_6897);
and U14204 (N_14204,N_6919,N_7191);
nand U14205 (N_14205,N_11058,N_8142);
xor U14206 (N_14206,N_11091,N_7014);
and U14207 (N_14207,N_8456,N_11658);
nand U14208 (N_14208,N_9838,N_10867);
or U14209 (N_14209,N_11201,N_7144);
nand U14210 (N_14210,N_6819,N_9714);
and U14211 (N_14211,N_8806,N_6385);
and U14212 (N_14212,N_9222,N_9568);
or U14213 (N_14213,N_8918,N_10259);
or U14214 (N_14214,N_11034,N_7382);
nor U14215 (N_14215,N_9712,N_7035);
and U14216 (N_14216,N_9612,N_11423);
and U14217 (N_14217,N_8010,N_6950);
and U14218 (N_14218,N_12192,N_7931);
and U14219 (N_14219,N_9323,N_10625);
or U14220 (N_14220,N_9296,N_10511);
and U14221 (N_14221,N_11945,N_11952);
nor U14222 (N_14222,N_10785,N_7406);
or U14223 (N_14223,N_11296,N_8469);
nor U14224 (N_14224,N_8900,N_10420);
or U14225 (N_14225,N_8540,N_7443);
or U14226 (N_14226,N_8197,N_11020);
nand U14227 (N_14227,N_9496,N_12445);
nand U14228 (N_14228,N_10116,N_11229);
nand U14229 (N_14229,N_11471,N_11260);
nand U14230 (N_14230,N_11620,N_12392);
xnor U14231 (N_14231,N_7878,N_8028);
nor U14232 (N_14232,N_8523,N_12018);
and U14233 (N_14233,N_10385,N_11981);
nor U14234 (N_14234,N_10801,N_9806);
and U14235 (N_14235,N_7863,N_8067);
or U14236 (N_14236,N_11680,N_10538);
or U14237 (N_14237,N_11883,N_8232);
or U14238 (N_14238,N_11932,N_11141);
and U14239 (N_14239,N_8959,N_7620);
and U14240 (N_14240,N_10055,N_8248);
nor U14241 (N_14241,N_10111,N_10769);
xor U14242 (N_14242,N_7457,N_9006);
nand U14243 (N_14243,N_9317,N_11980);
nand U14244 (N_14244,N_8727,N_7058);
or U14245 (N_14245,N_9909,N_7586);
or U14246 (N_14246,N_7545,N_8716);
nor U14247 (N_14247,N_11885,N_11491);
and U14248 (N_14248,N_9510,N_9550);
or U14249 (N_14249,N_10791,N_8829);
and U14250 (N_14250,N_7493,N_11153);
and U14251 (N_14251,N_7286,N_9653);
or U14252 (N_14252,N_10220,N_11906);
nor U14253 (N_14253,N_6635,N_6362);
or U14254 (N_14254,N_11825,N_7033);
nor U14255 (N_14255,N_10253,N_11619);
nand U14256 (N_14256,N_12060,N_6713);
nand U14257 (N_14257,N_6677,N_10062);
or U14258 (N_14258,N_7029,N_10665);
and U14259 (N_14259,N_7047,N_9471);
nor U14260 (N_14260,N_10642,N_11592);
or U14261 (N_14261,N_9922,N_7353);
or U14262 (N_14262,N_11391,N_9248);
and U14263 (N_14263,N_10993,N_12171);
nand U14264 (N_14264,N_11376,N_8282);
nor U14265 (N_14265,N_12315,N_8029);
and U14266 (N_14266,N_9537,N_8872);
or U14267 (N_14267,N_12297,N_9824);
nor U14268 (N_14268,N_8564,N_12129);
nand U14269 (N_14269,N_10492,N_10551);
and U14270 (N_14270,N_11438,N_8440);
nor U14271 (N_14271,N_8807,N_8096);
nor U14272 (N_14272,N_7729,N_7576);
or U14273 (N_14273,N_8234,N_10774);
and U14274 (N_14274,N_10869,N_12057);
or U14275 (N_14275,N_9906,N_9237);
or U14276 (N_14276,N_8268,N_11014);
and U14277 (N_14277,N_11923,N_10030);
nand U14278 (N_14278,N_6500,N_11347);
or U14279 (N_14279,N_10942,N_8929);
nor U14280 (N_14280,N_6392,N_8359);
and U14281 (N_14281,N_7316,N_12063);
nor U14282 (N_14282,N_11152,N_11348);
or U14283 (N_14283,N_11793,N_12275);
or U14284 (N_14284,N_8762,N_10548);
nand U14285 (N_14285,N_6755,N_7899);
or U14286 (N_14286,N_9662,N_7851);
or U14287 (N_14287,N_12488,N_8439);
and U14288 (N_14288,N_10412,N_7326);
and U14289 (N_14289,N_11459,N_10387);
and U14290 (N_14290,N_8606,N_11808);
xor U14291 (N_14291,N_8698,N_11167);
and U14292 (N_14292,N_7505,N_11569);
nand U14293 (N_14293,N_12210,N_11183);
nor U14294 (N_14294,N_7292,N_10444);
nor U14295 (N_14295,N_8996,N_8813);
nand U14296 (N_14296,N_8416,N_12427);
and U14297 (N_14297,N_8353,N_10513);
nor U14298 (N_14298,N_9828,N_9264);
and U14299 (N_14299,N_9480,N_10194);
and U14300 (N_14300,N_6515,N_8581);
nand U14301 (N_14301,N_6956,N_7799);
nor U14302 (N_14302,N_8039,N_11500);
or U14303 (N_14303,N_11908,N_10975);
or U14304 (N_14304,N_8172,N_6452);
and U14305 (N_14305,N_11687,N_8579);
nand U14306 (N_14306,N_6859,N_7608);
nor U14307 (N_14307,N_9659,N_10795);
nor U14308 (N_14308,N_12321,N_6464);
nor U14309 (N_14309,N_12256,N_11412);
nor U14310 (N_14310,N_9460,N_6648);
or U14311 (N_14311,N_10770,N_12013);
nor U14312 (N_14312,N_12002,N_10368);
nand U14313 (N_14313,N_6370,N_7996);
nor U14314 (N_14314,N_9444,N_12312);
nor U14315 (N_14315,N_8016,N_12328);
and U14316 (N_14316,N_8201,N_8903);
nand U14317 (N_14317,N_8635,N_8597);
nor U14318 (N_14318,N_7046,N_10287);
nand U14319 (N_14319,N_7530,N_12465);
and U14320 (N_14320,N_10126,N_11319);
and U14321 (N_14321,N_11574,N_8861);
nand U14322 (N_14322,N_10241,N_8621);
nand U14323 (N_14323,N_8713,N_7481);
and U14324 (N_14324,N_11330,N_10362);
nand U14325 (N_14325,N_8177,N_6397);
or U14326 (N_14326,N_9010,N_11997);
nand U14327 (N_14327,N_7399,N_6292);
nor U14328 (N_14328,N_7195,N_6945);
or U14329 (N_14329,N_7753,N_9184);
nand U14330 (N_14330,N_11148,N_10376);
nor U14331 (N_14331,N_8958,N_6849);
and U14332 (N_14332,N_11631,N_6298);
nand U14333 (N_14333,N_11346,N_9885);
or U14334 (N_14334,N_9655,N_12099);
nor U14335 (N_14335,N_7801,N_11023);
nand U14336 (N_14336,N_11166,N_11276);
nand U14337 (N_14337,N_9630,N_10242);
and U14338 (N_14338,N_6301,N_6805);
or U14339 (N_14339,N_10493,N_10809);
and U14340 (N_14340,N_10026,N_11965);
and U14341 (N_14341,N_8944,N_11824);
nor U14342 (N_14342,N_12168,N_10338);
and U14343 (N_14343,N_10998,N_8707);
nand U14344 (N_14344,N_12423,N_9623);
or U14345 (N_14345,N_11156,N_10823);
or U14346 (N_14346,N_7210,N_9142);
nor U14347 (N_14347,N_7958,N_11126);
or U14348 (N_14348,N_7644,N_7526);
nand U14349 (N_14349,N_8373,N_11895);
and U14350 (N_14350,N_11803,N_11960);
or U14351 (N_14351,N_12271,N_9554);
nor U14352 (N_14352,N_10949,N_10808);
or U14353 (N_14353,N_7826,N_9881);
xor U14354 (N_14354,N_6936,N_12159);
or U14355 (N_14355,N_7411,N_6272);
and U14356 (N_14356,N_7236,N_9218);
or U14357 (N_14357,N_8326,N_10204);
nand U14358 (N_14358,N_8531,N_11754);
and U14359 (N_14359,N_9253,N_8506);
and U14360 (N_14360,N_11609,N_6998);
or U14361 (N_14361,N_11372,N_9992);
nor U14362 (N_14362,N_7087,N_8170);
and U14363 (N_14363,N_7126,N_6600);
or U14364 (N_14364,N_10238,N_6463);
and U14365 (N_14365,N_12178,N_12234);
nand U14366 (N_14366,N_10643,N_7856);
and U14367 (N_14367,N_11294,N_7846);
or U14368 (N_14368,N_8164,N_9898);
nor U14369 (N_14369,N_7773,N_7612);
or U14370 (N_14370,N_11561,N_12005);
nor U14371 (N_14371,N_6879,N_11063);
or U14372 (N_14372,N_6578,N_10069);
nand U14373 (N_14373,N_11087,N_7603);
or U14374 (N_14374,N_9388,N_12046);
nand U14375 (N_14375,N_12096,N_6384);
nor U14376 (N_14376,N_12266,N_8150);
nand U14377 (N_14377,N_9986,N_8556);
and U14378 (N_14378,N_9846,N_12293);
or U14379 (N_14379,N_11440,N_7497);
nor U14380 (N_14380,N_8852,N_8984);
nor U14381 (N_14381,N_11805,N_9786);
nor U14382 (N_14382,N_7080,N_7804);
and U14383 (N_14383,N_7610,N_6653);
or U14384 (N_14384,N_12371,N_10002);
nor U14385 (N_14385,N_8228,N_11016);
and U14386 (N_14386,N_9685,N_11140);
or U14387 (N_14387,N_10928,N_10313);
nand U14388 (N_14388,N_8982,N_8198);
or U14389 (N_14389,N_9968,N_7095);
or U14390 (N_14390,N_12272,N_10714);
or U14391 (N_14391,N_8796,N_7446);
nand U14392 (N_14392,N_8399,N_9054);
nand U14393 (N_14393,N_12407,N_10392);
or U14394 (N_14394,N_11186,N_9478);
nand U14395 (N_14395,N_11225,N_8672);
and U14396 (N_14396,N_11292,N_9211);
or U14397 (N_14397,N_7028,N_8800);
nor U14398 (N_14398,N_6453,N_8208);
nand U14399 (N_14399,N_11078,N_11651);
nand U14400 (N_14400,N_6984,N_6314);
nor U14401 (N_14401,N_8609,N_8218);
nor U14402 (N_14402,N_6621,N_7815);
or U14403 (N_14403,N_7124,N_9921);
nor U14404 (N_14404,N_7655,N_10882);
nor U14405 (N_14405,N_9220,N_9465);
and U14406 (N_14406,N_10428,N_9506);
nor U14407 (N_14407,N_7649,N_10307);
nor U14408 (N_14408,N_8708,N_7669);
nand U14409 (N_14409,N_8079,N_8553);
nor U14410 (N_14410,N_10309,N_11864);
nand U14411 (N_14411,N_6921,N_10013);
or U14412 (N_14412,N_11729,N_9648);
nor U14413 (N_14413,N_12081,N_12474);
and U14414 (N_14414,N_9446,N_6547);
or U14415 (N_14415,N_11158,N_7070);
nor U14416 (N_14416,N_10613,N_11874);
or U14417 (N_14417,N_11393,N_11603);
nor U14418 (N_14418,N_11742,N_11102);
or U14419 (N_14419,N_6716,N_7918);
and U14420 (N_14420,N_11428,N_11200);
or U14421 (N_14421,N_11416,N_7613);
or U14422 (N_14422,N_9644,N_9304);
nor U14423 (N_14423,N_8145,N_6503);
and U14424 (N_14424,N_9649,N_12215);
nor U14425 (N_14425,N_7627,N_11406);
or U14426 (N_14426,N_8938,N_11930);
nand U14427 (N_14427,N_11122,N_11836);
nor U14428 (N_14428,N_10406,N_9413);
or U14429 (N_14429,N_7674,N_6287);
and U14430 (N_14430,N_7970,N_6745);
or U14431 (N_14431,N_10961,N_10234);
nand U14432 (N_14432,N_9750,N_10589);
nor U14433 (N_14433,N_9993,N_12127);
or U14434 (N_14434,N_10564,N_11045);
or U14435 (N_14435,N_7269,N_12326);
and U14436 (N_14436,N_12331,N_11388);
xnor U14437 (N_14437,N_6862,N_9641);
and U14438 (N_14438,N_9074,N_8591);
or U14439 (N_14439,N_8299,N_10524);
or U14440 (N_14440,N_10424,N_10879);
and U14441 (N_14441,N_10744,N_8588);
nor U14442 (N_14442,N_12314,N_9440);
or U14443 (N_14443,N_7560,N_8012);
nor U14444 (N_14444,N_11736,N_11238);
nor U14445 (N_14445,N_10106,N_9215);
or U14446 (N_14446,N_6527,N_7539);
xnor U14447 (N_14447,N_9418,N_9538);
nand U14448 (N_14448,N_8634,N_10560);
nand U14449 (N_14449,N_11846,N_12386);
nand U14450 (N_14450,N_7694,N_11925);
and U14451 (N_14451,N_7921,N_10608);
nor U14452 (N_14452,N_12123,N_6306);
nor U14453 (N_14453,N_10887,N_11139);
xnor U14454 (N_14454,N_6720,N_9912);
nand U14455 (N_14455,N_11663,N_8292);
and U14456 (N_14456,N_10698,N_11204);
and U14457 (N_14457,N_8011,N_8816);
nand U14458 (N_14458,N_9813,N_6303);
nor U14459 (N_14459,N_8552,N_7595);
nor U14460 (N_14460,N_9345,N_11150);
and U14461 (N_14461,N_9498,N_8664);
nand U14462 (N_14462,N_11044,N_8126);
and U14463 (N_14463,N_6317,N_11379);
and U14464 (N_14464,N_11550,N_12110);
or U14465 (N_14465,N_8916,N_9774);
or U14466 (N_14466,N_6955,N_12494);
and U14467 (N_14467,N_6669,N_8270);
or U14468 (N_14468,N_6688,N_8442);
nor U14469 (N_14469,N_9613,N_8747);
nand U14470 (N_14470,N_9353,N_10730);
or U14471 (N_14471,N_10060,N_11293);
or U14472 (N_14472,N_6747,N_9359);
nor U14473 (N_14473,N_7705,N_10416);
and U14474 (N_14474,N_11239,N_12041);
and U14475 (N_14475,N_8848,N_10157);
and U14476 (N_14476,N_9742,N_10274);
nor U14477 (N_14477,N_9914,N_7055);
or U14478 (N_14478,N_7329,N_9859);
and U14479 (N_14479,N_9687,N_11212);
nand U14480 (N_14480,N_11567,N_6918);
nand U14481 (N_14481,N_7504,N_10851);
or U14482 (N_14482,N_7429,N_11364);
or U14483 (N_14483,N_8931,N_12497);
nor U14484 (N_14484,N_12259,N_7957);
nor U14485 (N_14485,N_7905,N_9713);
and U14486 (N_14486,N_11867,N_9635);
and U14487 (N_14487,N_9871,N_8493);
and U14488 (N_14488,N_6481,N_9722);
nand U14489 (N_14489,N_9967,N_8304);
nor U14490 (N_14490,N_11694,N_7529);
nor U14491 (N_14491,N_9979,N_11689);
nor U14492 (N_14492,N_7343,N_7544);
nor U14493 (N_14493,N_8169,N_11048);
nor U14494 (N_14494,N_8643,N_6634);
and U14495 (N_14495,N_9185,N_6262);
nor U14496 (N_14496,N_12084,N_8076);
nand U14497 (N_14497,N_6783,N_11461);
nand U14498 (N_14498,N_8901,N_7973);
xnor U14499 (N_14499,N_6969,N_11434);
nor U14500 (N_14500,N_6895,N_7109);
or U14501 (N_14501,N_11976,N_6946);
and U14502 (N_14502,N_10648,N_7690);
or U14503 (N_14503,N_7445,N_7877);
or U14504 (N_14504,N_9886,N_7178);
xor U14505 (N_14505,N_6559,N_7100);
nand U14506 (N_14506,N_12218,N_9203);
or U14507 (N_14507,N_10595,N_6269);
nor U14508 (N_14508,N_7010,N_11184);
nor U14509 (N_14509,N_11105,N_7959);
or U14510 (N_14510,N_8850,N_10710);
and U14511 (N_14511,N_7262,N_10767);
or U14512 (N_14512,N_11553,N_8839);
and U14513 (N_14513,N_7798,N_8663);
nor U14514 (N_14514,N_6691,N_8781);
and U14515 (N_14515,N_7845,N_10474);
and U14516 (N_14516,N_10467,N_12491);
nor U14517 (N_14517,N_9952,N_8278);
nor U14518 (N_14518,N_9078,N_10430);
and U14519 (N_14519,N_7521,N_11611);
or U14520 (N_14520,N_7271,N_9128);
and U14521 (N_14521,N_8183,N_9855);
nor U14522 (N_14522,N_9116,N_7351);
and U14523 (N_14523,N_10402,N_9865);
or U14524 (N_14524,N_12121,N_10695);
nand U14525 (N_14525,N_10806,N_9845);
or U14526 (N_14526,N_8024,N_10666);
nor U14527 (N_14527,N_11411,N_11065);
or U14528 (N_14528,N_11806,N_6817);
nand U14529 (N_14529,N_7264,N_7723);
nor U14530 (N_14530,N_11523,N_12118);
or U14531 (N_14531,N_12303,N_11192);
or U14532 (N_14532,N_8427,N_11719);
or U14533 (N_14533,N_8533,N_12043);
or U14534 (N_14534,N_6277,N_12246);
nand U14535 (N_14535,N_8669,N_9955);
nor U14536 (N_14536,N_7909,N_9810);
and U14537 (N_14537,N_10209,N_7643);
nand U14538 (N_14538,N_10566,N_7968);
and U14539 (N_14539,N_9313,N_7232);
and U14540 (N_14540,N_9551,N_7822);
nand U14541 (N_14541,N_9182,N_6813);
and U14542 (N_14542,N_7325,N_10646);
nand U14543 (N_14543,N_6786,N_10064);
and U14544 (N_14544,N_10455,N_7059);
and U14545 (N_14545,N_11496,N_8702);
and U14546 (N_14546,N_8357,N_11771);
or U14547 (N_14547,N_9809,N_8657);
and U14548 (N_14548,N_9565,N_11881);
or U14549 (N_14549,N_9830,N_12279);
or U14550 (N_14550,N_11998,N_8108);
nor U14551 (N_14551,N_10521,N_11903);
nor U14552 (N_14552,N_11777,N_11441);
nor U14553 (N_14553,N_7436,N_9431);
nand U14554 (N_14554,N_11036,N_12072);
and U14555 (N_14555,N_11310,N_6584);
nor U14556 (N_14556,N_7695,N_6886);
nand U14557 (N_14557,N_7168,N_11655);
or U14558 (N_14558,N_11473,N_6704);
nor U14559 (N_14559,N_9135,N_10150);
nor U14560 (N_14560,N_11021,N_8233);
nor U14561 (N_14561,N_10609,N_10257);
or U14562 (N_14562,N_12338,N_6375);
nand U14563 (N_14563,N_10308,N_10211);
nor U14564 (N_14564,N_10597,N_9892);
nor U14565 (N_14565,N_8086,N_9171);
nor U14566 (N_14566,N_12327,N_7633);
nor U14567 (N_14567,N_6830,N_11509);
or U14568 (N_14568,N_6381,N_11605);
nand U14569 (N_14569,N_8355,N_11453);
nor U14570 (N_14570,N_6402,N_8528);
or U14571 (N_14571,N_11670,N_10687);
and U14572 (N_14572,N_8212,N_10963);
nor U14573 (N_14573,N_6476,N_11912);
or U14574 (N_14574,N_11197,N_10776);
or U14575 (N_14575,N_11389,N_6549);
nor U14576 (N_14576,N_9985,N_11510);
and U14577 (N_14577,N_7821,N_10239);
nand U14578 (N_14578,N_8772,N_8524);
and U14579 (N_14579,N_8124,N_8840);
and U14580 (N_14580,N_6966,N_10024);
nand U14581 (N_14581,N_6843,N_10821);
and U14582 (N_14582,N_9522,N_10205);
and U14583 (N_14583,N_10291,N_9484);
nand U14584 (N_14584,N_8178,N_7415);
nand U14585 (N_14585,N_7556,N_9283);
or U14586 (N_14586,N_12175,N_9866);
or U14587 (N_14587,N_7719,N_6441);
and U14588 (N_14588,N_9368,N_6593);
and U14589 (N_14589,N_7571,N_11936);
nand U14590 (N_14590,N_10571,N_11710);
or U14591 (N_14591,N_7365,N_7514);
and U14592 (N_14592,N_10350,N_8558);
nor U14593 (N_14593,N_6923,N_11576);
nand U14594 (N_14594,N_11780,N_10229);
nor U14595 (N_14595,N_7079,N_10670);
or U14596 (N_14596,N_10186,N_9358);
nor U14597 (N_14597,N_7739,N_12040);
nand U14598 (N_14598,N_9236,N_10747);
nor U14599 (N_14599,N_11111,N_10722);
nand U14600 (N_14600,N_8910,N_11875);
and U14601 (N_14601,N_8845,N_6967);
or U14602 (N_14602,N_8898,N_10384);
and U14603 (N_14603,N_10356,N_6739);
nand U14604 (N_14604,N_11005,N_10637);
nor U14605 (N_14605,N_10702,N_7665);
nor U14606 (N_14606,N_11543,N_7193);
or U14607 (N_14607,N_6656,N_11176);
or U14608 (N_14608,N_12468,N_6522);
nand U14609 (N_14609,N_11410,N_10178);
xnor U14610 (N_14610,N_7770,N_6439);
nor U14611 (N_14611,N_9669,N_9999);
nor U14612 (N_14612,N_8599,N_7283);
nand U14613 (N_14613,N_8759,N_8042);
and U14614 (N_14614,N_6996,N_6618);
nor U14615 (N_14615,N_7513,N_8836);
and U14616 (N_14616,N_7234,N_11989);
nor U14617 (N_14617,N_9029,N_11865);
nor U14618 (N_14618,N_11935,N_10372);
or U14619 (N_14619,N_7653,N_10170);
nand U14620 (N_14620,N_9266,N_10554);
nor U14621 (N_14621,N_11252,N_11002);
or U14622 (N_14622,N_7876,N_11984);
nor U14623 (N_14623,N_8685,N_10151);
or U14624 (N_14624,N_7153,N_11833);
and U14625 (N_14625,N_9558,N_6837);
nand U14626 (N_14626,N_6625,N_10542);
and U14627 (N_14627,N_9879,N_6361);
nand U14628 (N_14628,N_7554,N_8805);
nor U14629 (N_14629,N_11498,N_9911);
or U14630 (N_14630,N_11823,N_11549);
nor U14631 (N_14631,N_11773,N_7592);
nand U14632 (N_14632,N_9512,N_8725);
nor U14633 (N_14633,N_7588,N_7052);
nand U14634 (N_14634,N_10450,N_10228);
and U14635 (N_14635,N_11859,N_7491);
or U14636 (N_14636,N_9856,N_7622);
nand U14637 (N_14637,N_10838,N_9940);
or U14638 (N_14638,N_7389,N_11557);
and U14639 (N_14639,N_7730,N_11630);
and U14640 (N_14640,N_10109,N_7535);
and U14641 (N_14641,N_11103,N_9103);
nor U14642 (N_14642,N_7081,N_6926);
and U14643 (N_14643,N_6346,N_9373);
nor U14644 (N_14644,N_9624,N_11800);
nand U14645 (N_14645,N_7585,N_6483);
or U14646 (N_14646,N_8963,N_12299);
nand U14647 (N_14647,N_10470,N_11585);
nand U14648 (N_14648,N_6347,N_9782);
or U14649 (N_14649,N_8205,N_10262);
and U14650 (N_14650,N_9405,N_12088);
or U14651 (N_14651,N_10617,N_10948);
nand U14652 (N_14652,N_11897,N_7768);
nor U14653 (N_14653,N_9027,N_11514);
nor U14654 (N_14654,N_9595,N_7313);
and U14655 (N_14655,N_11519,N_11791);
nand U14656 (N_14656,N_10868,N_9633);
nand U14657 (N_14657,N_11886,N_9640);
or U14658 (N_14658,N_12150,N_7577);
and U14659 (N_14659,N_7362,N_9789);
nor U14660 (N_14660,N_6639,N_12295);
nor U14661 (N_14661,N_10061,N_9101);
nand U14662 (N_14662,N_7501,N_11547);
nor U14663 (N_14663,N_10906,N_7935);
and U14664 (N_14664,N_10649,N_6892);
nor U14665 (N_14665,N_8940,N_10319);
nor U14666 (N_14666,N_11726,N_8814);
and U14667 (N_14667,N_7012,N_7659);
nor U14668 (N_14668,N_8111,N_9564);
or U14669 (N_14669,N_10443,N_10182);
and U14670 (N_14670,N_8458,N_6825);
and U14671 (N_14671,N_8547,N_12455);
or U14672 (N_14672,N_11353,N_8360);
or U14673 (N_14673,N_8410,N_10373);
nand U14674 (N_14674,N_9569,N_7103);
nor U14675 (N_14675,N_8094,N_11338);
nor U14676 (N_14676,N_9043,N_7409);
or U14677 (N_14677,N_7810,N_11280);
nor U14678 (N_14678,N_8063,N_8323);
nand U14679 (N_14679,N_8482,N_11108);
nor U14680 (N_14680,N_12128,N_6766);
and U14681 (N_14681,N_8034,N_7668);
and U14682 (N_14682,N_8970,N_7473);
and U14683 (N_14683,N_10037,N_7704);
or U14684 (N_14684,N_9723,N_8915);
or U14685 (N_14685,N_11764,N_7652);
nand U14686 (N_14686,N_7776,N_6523);
nor U14687 (N_14687,N_10009,N_7165);
or U14688 (N_14688,N_7412,N_6422);
and U14689 (N_14689,N_6554,N_11295);
nand U14690 (N_14690,N_11028,N_9631);
nor U14691 (N_14691,N_10068,N_8751);
xor U14692 (N_14692,N_8069,N_9495);
and U14693 (N_14693,N_11084,N_11397);
nor U14694 (N_14694,N_6365,N_8154);
and U14695 (N_14695,N_9584,N_9772);
nand U14696 (N_14696,N_6861,N_8799);
nand U14697 (N_14697,N_10678,N_7282);
xnor U14698 (N_14698,N_11451,N_11208);
and U14699 (N_14699,N_8962,N_10391);
or U14700 (N_14700,N_7512,N_9286);
or U14701 (N_14701,N_6985,N_11478);
nand U14702 (N_14702,N_8227,N_9549);
and U14703 (N_14703,N_6297,N_7842);
nand U14704 (N_14704,N_10849,N_9840);
or U14705 (N_14705,N_7522,N_6466);
nand U14706 (N_14706,N_6425,N_7039);
nand U14707 (N_14707,N_7173,N_11497);
or U14708 (N_14708,N_10216,N_7927);
nor U14709 (N_14709,N_12454,N_9301);
or U14710 (N_14710,N_8538,N_8769);
nand U14711 (N_14711,N_8337,N_6733);
and U14712 (N_14712,N_9977,N_10386);
nand U14713 (N_14713,N_12471,N_8331);
and U14714 (N_14714,N_11625,N_9256);
nor U14715 (N_14715,N_11581,N_11827);
xor U14716 (N_14716,N_6640,N_6820);
and U14717 (N_14717,N_12345,N_12350);
and U14718 (N_14718,N_8760,N_11963);
nand U14719 (N_14719,N_9708,N_9377);
nand U14720 (N_14720,N_9026,N_6282);
nor U14721 (N_14721,N_11324,N_7888);
and U14722 (N_14722,N_9657,N_9178);
or U14723 (N_14723,N_7887,N_6541);
nor U14724 (N_14724,N_10733,N_10910);
nor U14725 (N_14725,N_6268,N_7536);
and U14726 (N_14726,N_11417,N_7089);
nor U14727 (N_14727,N_10088,N_7065);
or U14728 (N_14728,N_10768,N_11699);
nand U14729 (N_14729,N_12226,N_8344);
or U14730 (N_14730,N_10850,N_11494);
nand U14731 (N_14731,N_9300,N_9177);
and U14732 (N_14732,N_6575,N_9591);
or U14733 (N_14733,N_9994,N_8754);
or U14734 (N_14734,N_6884,N_7430);
and U14735 (N_14735,N_8490,N_12114);
nor U14736 (N_14736,N_11202,N_8776);
or U14737 (N_14737,N_8673,N_9589);
xnor U14738 (N_14738,N_9395,N_10682);
or U14739 (N_14739,N_11218,N_12411);
nor U14740 (N_14740,N_6294,N_9850);
or U14741 (N_14741,N_10081,N_12308);
nor U14742 (N_14742,N_9872,N_12478);
and U14743 (N_14743,N_12253,N_10525);
and U14744 (N_14744,N_9610,N_11424);
nand U14745 (N_14745,N_7461,N_7335);
nand U14746 (N_14746,N_7507,N_8059);
nor U14747 (N_14747,N_12196,N_7599);
and U14748 (N_14748,N_6335,N_7759);
nand U14749 (N_14749,N_8391,N_12252);
and U14750 (N_14750,N_10759,N_12288);
or U14751 (N_14751,N_8854,N_6474);
and U14752 (N_14752,N_9008,N_7091);
or U14753 (N_14753,N_10582,N_9105);
or U14754 (N_14754,N_7806,N_9189);
and U14755 (N_14755,N_9876,N_7735);
nand U14756 (N_14756,N_11163,N_10580);
or U14757 (N_14757,N_7813,N_10848);
and U14758 (N_14758,N_6336,N_9214);
and U14759 (N_14759,N_10796,N_7637);
nand U14760 (N_14760,N_8120,N_7248);
nor U14761 (N_14761,N_11668,N_9033);
nor U14762 (N_14762,N_8379,N_7765);
nand U14763 (N_14763,N_10908,N_10826);
or U14764 (N_14764,N_10894,N_9058);
and U14765 (N_14765,N_8699,N_7837);
xor U14766 (N_14766,N_7230,N_11327);
or U14767 (N_14767,N_10676,N_9527);
and U14768 (N_14768,N_7228,N_11443);
and U14769 (N_14769,N_7350,N_7929);
nand U14770 (N_14770,N_10184,N_11488);
or U14771 (N_14771,N_11988,N_7226);
nand U14772 (N_14772,N_9486,N_8050);
or U14773 (N_14773,N_9410,N_9884);
nor U14774 (N_14774,N_10137,N_11249);
and U14775 (N_14775,N_7356,N_10726);
and U14776 (N_14776,N_11645,N_6428);
nor U14777 (N_14777,N_9608,N_7072);
nand U14778 (N_14778,N_7073,N_8810);
nor U14779 (N_14779,N_9254,N_6972);
and U14780 (N_14780,N_6809,N_12414);
and U14781 (N_14781,N_6959,N_7625);
nand U14782 (N_14782,N_8789,N_7132);
nor U14783 (N_14783,N_10355,N_7712);
or U14784 (N_14784,N_6654,N_10400);
nor U14785 (N_14785,N_10086,N_10115);
nand U14786 (N_14786,N_8398,N_12174);
nor U14787 (N_14787,N_11024,N_11244);
or U14788 (N_14788,N_9596,N_10690);
xor U14789 (N_14789,N_9169,N_6516);
nor U14790 (N_14790,N_6741,N_9980);
and U14791 (N_14791,N_12152,N_6975);
or U14792 (N_14792,N_10530,N_6818);
and U14793 (N_14793,N_11739,N_8015);
nor U14794 (N_14794,N_11213,N_6982);
nand U14795 (N_14795,N_11187,N_8603);
nand U14796 (N_14796,N_11043,N_8788);
and U14797 (N_14797,N_11671,N_12098);
nand U14798 (N_14798,N_12470,N_10555);
and U14799 (N_14799,N_9957,N_9724);
nor U14800 (N_14800,N_7641,N_9208);
and U14801 (N_14801,N_9508,N_7164);
nand U14802 (N_14802,N_8259,N_8450);
nor U14803 (N_14803,N_7543,N_9196);
or U14804 (N_14804,N_10441,N_10273);
or U14805 (N_14805,N_8210,N_11866);
or U14806 (N_14806,N_11484,N_8354);
and U14807 (N_14807,N_10432,N_6507);
nor U14808 (N_14808,N_12378,N_10201);
nand U14809 (N_14809,N_8773,N_9799);
or U14810 (N_14810,N_8161,N_8488);
nor U14811 (N_14811,N_10950,N_6794);
and U14812 (N_14812,N_9989,N_9217);
nor U14813 (N_14813,N_7857,N_10655);
nand U14814 (N_14814,N_8722,N_8182);
and U14815 (N_14815,N_9547,N_7263);
or U14816 (N_14816,N_10939,N_9455);
or U14817 (N_14817,N_12311,N_9310);
or U14818 (N_14818,N_12119,N_6980);
or U14819 (N_14819,N_6842,N_9833);
and U14820 (N_14820,N_9275,N_6318);
nand U14821 (N_14821,N_11301,N_11077);
xnor U14822 (N_14822,N_12067,N_6281);
nor U14823 (N_14823,N_8602,N_6796);
or U14824 (N_14824,N_11427,N_7871);
or U14825 (N_14825,N_10041,N_12132);
nand U14826 (N_14826,N_10512,N_7787);
nand U14827 (N_14827,N_6288,N_8770);
or U14828 (N_14828,N_6290,N_8921);
and U14829 (N_14829,N_9122,N_12106);
nand U14830 (N_14830,N_10141,N_8334);
and U14831 (N_14831,N_6769,N_6429);
nand U14832 (N_14832,N_7998,N_9730);
and U14833 (N_14833,N_11335,N_6871);
or U14834 (N_14834,N_10173,N_12183);
or U14835 (N_14835,N_11307,N_7259);
and U14836 (N_14836,N_11356,N_10409);
nand U14837 (N_14837,N_6681,N_7495);
and U14838 (N_14838,N_10732,N_11572);
nand U14839 (N_14839,N_8584,N_10388);
nand U14840 (N_14840,N_7618,N_11071);
nor U14841 (N_14841,N_8141,N_11794);
nand U14842 (N_14842,N_11700,N_9361);
nand U14843 (N_14843,N_11850,N_11198);
or U14844 (N_14844,N_7466,N_10601);
nand U14845 (N_14845,N_10679,N_11768);
or U14846 (N_14846,N_8765,N_10813);
or U14847 (N_14847,N_7844,N_9585);
and U14848 (N_14848,N_11949,N_11590);
nand U14849 (N_14849,N_8485,N_7139);
nor U14850 (N_14850,N_6331,N_9017);
nand U14851 (N_14851,N_10870,N_8258);
and U14852 (N_14852,N_6605,N_8414);
or U14853 (N_14853,N_8977,N_11318);
nor U14854 (N_14854,N_8217,N_8239);
nor U14855 (N_14855,N_10105,N_9327);
and U14856 (N_14856,N_11690,N_11278);
nand U14857 (N_14857,N_11436,N_11921);
and U14858 (N_14858,N_9863,N_11336);
or U14859 (N_14859,N_11884,N_8684);
nor U14860 (N_14860,N_6997,N_8492);
nand U14861 (N_14861,N_7053,N_8496);
and U14862 (N_14862,N_8038,N_10407);
nand U14863 (N_14863,N_6596,N_7550);
nor U14864 (N_14864,N_7401,N_10708);
nor U14865 (N_14865,N_8532,N_7177);
or U14866 (N_14866,N_8640,N_11697);
nor U14867 (N_14867,N_9706,N_8527);
nand U14868 (N_14868,N_7187,N_7890);
or U14869 (N_14869,N_10101,N_10878);
nand U14870 (N_14870,N_11162,N_7104);
nor U14871 (N_14871,N_11415,N_7843);
or U14872 (N_14872,N_11852,N_8484);
nand U14873 (N_14873,N_11060,N_12344);
nor U14874 (N_14874,N_9201,N_6914);
nor U14875 (N_14875,N_11621,N_8726);
nand U14876 (N_14876,N_10728,N_9699);
or U14877 (N_14877,N_9598,N_12228);
or U14878 (N_14878,N_8167,N_8507);
and U14879 (N_14879,N_8803,N_8614);
or U14880 (N_14880,N_10986,N_7037);
or U14881 (N_14881,N_10078,N_7131);
and U14882 (N_14882,N_11571,N_6855);
and U14883 (N_14883,N_7237,N_8188);
nand U14884 (N_14884,N_7782,N_10276);
nor U14885 (N_14885,N_9616,N_12052);
or U14886 (N_14886,N_9594,N_8519);
and U14887 (N_14887,N_7525,N_7778);
or U14888 (N_14888,N_6742,N_12239);
and U14889 (N_14889,N_9022,N_8189);
or U14890 (N_14890,N_11331,N_12025);
and U14891 (N_14891,N_10923,N_8974);
and U14892 (N_14892,N_8832,N_11677);
nand U14893 (N_14893,N_9835,N_10721);
nand U14894 (N_14894,N_10924,N_9923);
nand U14895 (N_14895,N_10802,N_9532);
nand U14896 (N_14896,N_10197,N_6684);
nand U14897 (N_14897,N_11290,N_8043);
nor U14898 (N_14898,N_11613,N_7867);
nor U14899 (N_14899,N_7471,N_9335);
nand U14900 (N_14900,N_9543,N_10083);
or U14901 (N_14901,N_12083,N_6806);
nand U14902 (N_14902,N_11240,N_9004);
and U14903 (N_14903,N_7895,N_11282);
nand U14904 (N_14904,N_7991,N_7755);
or U14905 (N_14905,N_9160,N_8949);
and U14906 (N_14906,N_8434,N_9962);
nand U14907 (N_14907,N_6322,N_10001);
or U14908 (N_14908,N_7287,N_10433);
nor U14909 (N_14909,N_6284,N_6826);
nand U14910 (N_14910,N_9832,N_10803);
nand U14911 (N_14911,N_11542,N_6960);
and U14912 (N_14912,N_9916,N_7422);
or U14913 (N_14913,N_6300,N_10568);
and U14914 (N_14914,N_8535,N_6504);
or U14915 (N_14915,N_11552,N_7400);
and U14916 (N_14916,N_8730,N_9905);
and U14917 (N_14917,N_11233,N_8056);
nand U14918 (N_14918,N_8361,N_8693);
and U14919 (N_14919,N_11110,N_11042);
nor U14920 (N_14920,N_11432,N_8412);
nor U14921 (N_14921,N_6674,N_10264);
nand U14922 (N_14922,N_10883,N_9433);
nor U14923 (N_14923,N_7743,N_9815);
nand U14924 (N_14924,N_8454,N_8583);
and U14925 (N_14925,N_9179,N_6490);
or U14926 (N_14926,N_7864,N_12452);
nor U14927 (N_14927,N_11113,N_10719);
nand U14928 (N_14928,N_12310,N_10630);
nor U14929 (N_14929,N_7953,N_8281);
nand U14930 (N_14930,N_10135,N_8009);
nor U14931 (N_14931,N_8008,N_7339);
and U14932 (N_14932,N_7911,N_11025);
or U14933 (N_14933,N_9570,N_11493);
nor U14934 (N_14934,N_6315,N_7247);
nor U14935 (N_14935,N_11499,N_8937);
nor U14936 (N_14936,N_9053,N_8766);
nor U14937 (N_14937,N_12146,N_10890);
nand U14938 (N_14938,N_10958,N_7150);
nor U14939 (N_14939,N_7881,N_7145);
nor U14940 (N_14940,N_11807,N_8925);
nor U14941 (N_14941,N_8092,N_6770);
or U14942 (N_14942,N_8936,N_6642);
nor U14943 (N_14943,N_10394,N_6285);
and U14944 (N_14944,N_11902,N_8252);
nor U14945 (N_14945,N_9259,N_9468);
and U14946 (N_14946,N_10225,N_10818);
nand U14947 (N_14947,N_9566,N_11380);
nand U14948 (N_14948,N_7780,N_11813);
or U14949 (N_14949,N_8753,N_11224);
nor U14950 (N_14950,N_9951,N_9890);
and U14951 (N_14951,N_6352,N_6445);
and U14952 (N_14952,N_11199,N_7395);
nor U14953 (N_14953,N_11878,N_7272);
or U14954 (N_14954,N_7926,N_7437);
nand U14955 (N_14955,N_9231,N_12160);
nand U14956 (N_14956,N_12036,N_10936);
or U14957 (N_14957,N_7238,N_11136);
nor U14958 (N_14958,N_6857,N_10022);
nor U14959 (N_14959,N_11115,N_7206);
or U14960 (N_14960,N_6343,N_11517);
nor U14961 (N_14961,N_12257,N_9717);
nand U14962 (N_14962,N_10295,N_6340);
and U14963 (N_14963,N_8511,N_9204);
or U14964 (N_14964,N_11693,N_12379);
and U14965 (N_14965,N_7952,N_11396);
and U14966 (N_14966,N_10152,N_9668);
nand U14967 (N_14967,N_9167,N_10877);
nand U14968 (N_14968,N_8191,N_10016);
nor U14969 (N_14969,N_8516,N_10547);
nand U14970 (N_14970,N_8756,N_10845);
or U14971 (N_14971,N_9767,N_9779);
nor U14972 (N_14972,N_10522,N_11763);
or U14973 (N_14973,N_9294,N_9354);
or U14974 (N_14974,N_8041,N_7309);
nand U14975 (N_14975,N_6293,N_10143);
nor U14976 (N_14976,N_8294,N_11477);
and U14977 (N_14977,N_9731,N_7900);
nand U14978 (N_14978,N_7994,N_12417);
nor U14979 (N_14979,N_9297,N_11382);
nand U14980 (N_14980,N_8325,N_6373);
nor U14981 (N_14981,N_12195,N_7687);
and U14982 (N_14982,N_12245,N_11887);
or U14983 (N_14983,N_8784,N_11880);
and U14984 (N_14984,N_10348,N_7684);
xor U14985 (N_14985,N_11216,N_9966);
nor U14986 (N_14986,N_9801,N_6815);
or U14987 (N_14987,N_9474,N_6845);
nor U14988 (N_14988,N_11938,N_12330);
xnor U14989 (N_14989,N_8645,N_12336);
and U14990 (N_14990,N_11454,N_10245);
nand U14991 (N_14991,N_11524,N_8539);
or U14992 (N_14992,N_9120,N_7258);
nand U14993 (N_14993,N_10087,N_9246);
nor U14994 (N_14994,N_6778,N_7090);
and U14995 (N_14995,N_12095,N_8935);
nand U14996 (N_14996,N_7219,N_7590);
nor U14997 (N_14997,N_10667,N_10070);
nor U14998 (N_14998,N_11979,N_12260);
or U14999 (N_14999,N_9136,N_7589);
nor U15000 (N_15000,N_11339,N_9854);
and U15001 (N_15001,N_8930,N_10065);
or U15002 (N_15002,N_9540,N_8335);
and U15003 (N_15003,N_11511,N_7186);
nand U15004 (N_15004,N_12194,N_8106);
and U15005 (N_15005,N_11188,N_12016);
nor U15006 (N_15006,N_8417,N_6744);
or U15007 (N_15007,N_10880,N_7075);
or U15008 (N_15008,N_12443,N_10477);
or U15009 (N_15009,N_11068,N_12138);
nor U15010 (N_15010,N_10004,N_12145);
nor U15011 (N_15011,N_11501,N_8125);
or U15012 (N_15012,N_8749,N_10841);
or U15013 (N_15013,N_6512,N_8005);
nor U15014 (N_15014,N_10592,N_9857);
or U15015 (N_15015,N_9091,N_10615);
nor U15016 (N_15016,N_10092,N_9118);
nand U15017 (N_15017,N_9018,N_11041);
or U15018 (N_15018,N_9138,N_8062);
nor U15019 (N_15019,N_9348,N_10353);
nand U15020 (N_15020,N_11614,N_8473);
and U15021 (N_15021,N_10805,N_7334);
nor U15022 (N_15022,N_12402,N_6524);
or U15023 (N_15023,N_9816,N_9165);
nor U15024 (N_15024,N_9895,N_9252);
or U15025 (N_15025,N_9739,N_7898);
and U15026 (N_15026,N_9907,N_7358);
and U15027 (N_15027,N_7482,N_7208);
and U15028 (N_15028,N_8095,N_7858);
nor U15029 (N_15029,N_7155,N_7172);
and U15030 (N_15030,N_8582,N_9328);
or U15031 (N_15031,N_11180,N_7480);
or U15032 (N_15032,N_8068,N_8243);
nor U15033 (N_15033,N_11378,N_10360);
nand U15034 (N_15034,N_9691,N_7108);
xnor U15035 (N_15035,N_9601,N_6758);
and U15036 (N_15036,N_7444,N_9664);
nor U15037 (N_15037,N_11189,N_6396);
and U15038 (N_15038,N_8276,N_9505);
or U15039 (N_15039,N_9257,N_6612);
and U15040 (N_15040,N_10012,N_10085);
nor U15041 (N_15041,N_10110,N_12400);
or U15042 (N_15042,N_7678,N_10517);
or U15043 (N_15043,N_6850,N_10258);
nor U15044 (N_15044,N_7552,N_6455);
nand U15045 (N_15045,N_10968,N_8590);
and U15046 (N_15046,N_7161,N_11715);
nor U15047 (N_15047,N_9466,N_8680);
nor U15048 (N_15048,N_10155,N_9945);
nand U15049 (N_15049,N_9438,N_7642);
nand U15050 (N_15050,N_12026,N_9153);
nand U15051 (N_15051,N_10293,N_6949);
nand U15052 (N_15052,N_12137,N_6910);
nand U15053 (N_15053,N_10741,N_6426);
or U15054 (N_15054,N_6256,N_7452);
or U15055 (N_15055,N_11064,N_11149);
nand U15056 (N_15056,N_11940,N_8646);
nor U15057 (N_15057,N_11430,N_8873);
nor U15058 (N_15058,N_7319,N_8139);
and U15059 (N_15059,N_7933,N_7656);
or U15060 (N_15060,N_12430,N_9729);
nor U15061 (N_15061,N_12184,N_11173);
or U15062 (N_15062,N_11320,N_10565);
nor U15063 (N_15063,N_10794,N_10005);
nand U15064 (N_15064,N_9260,N_11302);
nor U15065 (N_15065,N_11469,N_8537);
and U15066 (N_15066,N_11681,N_10380);
nand U15067 (N_15067,N_9925,N_10125);
or U15068 (N_15068,N_7442,N_10289);
and U15069 (N_15069,N_8758,N_6440);
nand U15070 (N_15070,N_8040,N_12126);
nor U15071 (N_15071,N_9756,N_7831);
nand U15072 (N_15072,N_8037,N_8165);
nor U15073 (N_15073,N_6374,N_6468);
or U15074 (N_15074,N_7063,N_9429);
and U15075 (N_15075,N_11696,N_8926);
nor U15076 (N_15076,N_7534,N_11251);
and U15077 (N_15077,N_12479,N_9582);
nor U15078 (N_15078,N_8774,N_12475);
nor U15079 (N_15079,N_12459,N_11920);
and U15080 (N_15080,N_8787,N_7614);
nor U15081 (N_15081,N_9295,N_7557);
nand U15082 (N_15082,N_8870,N_8374);
nor U15083 (N_15083,N_8743,N_11779);
or U15084 (N_15084,N_7332,N_12435);
and U15085 (N_15085,N_12015,N_6993);
and U15086 (N_15086,N_9917,N_6614);
nor U15087 (N_15087,N_9141,N_12367);
nand U15088 (N_15088,N_9463,N_12335);
and U15089 (N_15089,N_11518,N_6706);
nand U15090 (N_15090,N_7122,N_8147);
nand U15091 (N_15091,N_9695,N_8402);
or U15092 (N_15092,N_8146,N_12384);
or U15093 (N_15093,N_9679,N_6970);
nor U15094 (N_15094,N_8997,N_9299);
nor U15095 (N_15095,N_12329,N_8035);
and U15096 (N_15096,N_9156,N_10960);
nor U15097 (N_15097,N_11602,N_10383);
nand U15098 (N_15098,N_8637,N_8317);
nor U15099 (N_15099,N_10735,N_7661);
and U15100 (N_15100,N_8327,N_11313);
and U15101 (N_15101,N_9193,N_7041);
nand U15102 (N_15102,N_10408,N_9340);
or U15103 (N_15103,N_8429,N_9654);
nor U15104 (N_15104,N_12325,N_9716);
nand U15105 (N_15105,N_12105,N_8611);
and U15106 (N_15106,N_12362,N_11798);
and U15107 (N_15107,N_7314,N_9567);
nand U15108 (N_15108,N_9935,N_11209);
or U15109 (N_15109,N_11937,N_11458);
nor U15110 (N_15110,N_10187,N_9874);
or U15111 (N_15111,N_7093,N_10322);
and U15112 (N_15112,N_11797,N_7032);
nor U15113 (N_15113,N_10440,N_10675);
nor U15114 (N_15114,N_9579,N_11993);
nand U15115 (N_15115,N_6536,N_7306);
or U15116 (N_15116,N_10008,N_8924);
and U15117 (N_15117,N_8837,N_9202);
nor U15118 (N_15118,N_11259,N_8705);
nand U15119 (N_15119,N_10146,N_7229);
nand U15120 (N_15120,N_6824,N_11955);
or U15121 (N_15121,N_10663,N_6394);
nand U15122 (N_15122,N_9883,N_10210);
or U15123 (N_15123,N_6687,N_8237);
nor U15124 (N_15124,N_12006,N_10359);
xor U15125 (N_15125,N_7318,N_9970);
and U15126 (N_15126,N_6255,N_6710);
or U15127 (N_15127,N_11648,N_11531);
or U15128 (N_15128,N_9515,N_6828);
and U15129 (N_15129,N_9733,N_11992);
nand U15130 (N_15130,N_11076,N_12139);
and U15131 (N_15131,N_9529,N_7111);
or U15132 (N_15132,N_6645,N_8348);
nor U15133 (N_15133,N_12061,N_7174);
or U15134 (N_15134,N_9718,N_7107);
and U15135 (N_15135,N_11316,N_9430);
nand U15136 (N_15136,N_10761,N_6501);
nor U15137 (N_15137,N_6368,N_9332);
and U15138 (N_15138,N_11027,N_11082);
or U15139 (N_15139,N_6927,N_12090);
or U15140 (N_15140,N_11061,N_10294);
and U15141 (N_15141,N_7036,N_7650);
nand U15142 (N_15142,N_7999,N_9841);
and U15143 (N_15143,N_9223,N_9614);
or U15144 (N_15144,N_10858,N_9658);
xor U15145 (N_15145,N_6995,N_10844);
and U15146 (N_15146,N_10537,N_11732);
or U15147 (N_15147,N_11242,N_6611);
or U15148 (N_15148,N_10605,N_8881);
nor U15149 (N_15149,N_7378,N_8021);
nand U15150 (N_15150,N_8752,N_11480);
or U15151 (N_15151,N_6520,N_11343);
nand U15152 (N_15152,N_9740,N_12091);
nand U15153 (N_15153,N_12080,N_8856);
nand U15154 (N_15154,N_11872,N_6633);
xnor U15155 (N_15155,N_7054,N_8823);
and U15156 (N_15156,N_8470,N_11230);
or U15157 (N_15157,N_6775,N_11462);
or U15158 (N_15158,N_8734,N_6872);
and U15159 (N_15159,N_9581,N_9427);
nor U15160 (N_15160,N_9251,N_7393);
or U15161 (N_15161,N_6707,N_8695);
or U15162 (N_15162,N_7630,N_7621);
nand U15163 (N_15163,N_7667,N_7157);
nor U15164 (N_15164,N_11890,N_8906);
and U15165 (N_15165,N_8979,N_6643);
or U15166 (N_15166,N_9725,N_11263);
nor U15167 (N_15167,N_11098,N_9073);
or U15168 (N_15168,N_7969,N_9559);
or U15169 (N_15169,N_6929,N_10098);
and U15170 (N_15170,N_8424,N_12358);
or U15171 (N_15171,N_8104,N_6484);
nand U15172 (N_15172,N_7568,N_7602);
nor U15173 (N_15173,N_10147,N_10793);
and U15174 (N_15174,N_10130,N_11770);
nor U15175 (N_15175,N_9110,N_11008);
nand U15176 (N_15176,N_6847,N_6898);
and U15177 (N_15177,N_6697,N_6330);
or U15178 (N_15178,N_10049,N_7685);
nand U15179 (N_15179,N_9849,N_10014);
nor U15180 (N_15180,N_11772,N_8775);
nand U15181 (N_15181,N_12420,N_11688);
and U15182 (N_15182,N_11565,N_11266);
and U15183 (N_15183,N_11272,N_11593);
and U15184 (N_15184,N_7344,N_6574);
and U15185 (N_15185,N_12241,N_9036);
or U15186 (N_15186,N_7408,N_8300);
nor U15187 (N_15187,N_12368,N_8679);
nor U15188 (N_15188,N_7955,N_9249);
nand U15189 (N_15189,N_11961,N_6526);
nor U15190 (N_15190,N_6610,N_7775);
nand U15191 (N_15191,N_8394,N_7299);
nor U15192 (N_15192,N_8668,N_7938);
nor U15193 (N_15193,N_10836,N_9586);
and U15194 (N_15194,N_6763,N_7031);
and U15195 (N_15195,N_10367,N_7750);
nand U15196 (N_15196,N_9194,N_6354);
nor U15197 (N_15197,N_10261,N_7664);
nor U15198 (N_15198,N_6299,N_11714);
nor U15199 (N_15199,N_8099,N_11532);
or U15200 (N_15200,N_8792,N_7294);
nand U15201 (N_15201,N_8006,N_12031);
or U15202 (N_15202,N_11969,N_11734);
nand U15203 (N_15203,N_9681,N_12318);
nand U15204 (N_15204,N_12167,N_7947);
and U15205 (N_15205,N_10364,N_12086);
nand U15206 (N_15206,N_12406,N_9038);
and U15207 (N_15207,N_8027,N_8477);
and U15208 (N_15208,N_7945,N_7903);
nor U15209 (N_15209,N_11977,N_7990);
and U15210 (N_15210,N_8253,N_9763);
xnor U15211 (N_15211,N_10040,N_6983);
nor U15212 (N_15212,N_6302,N_8180);
xor U15213 (N_15213,N_6329,N_6558);
nand U15214 (N_15214,N_8392,N_7301);
nand U15215 (N_15215,N_10361,N_9230);
nor U15216 (N_15216,N_6701,N_12111);
nor U15217 (N_15217,N_8838,N_12233);
nor U15218 (N_15218,N_7607,N_9853);
or U15219 (N_15219,N_8486,N_6497);
or U15220 (N_15220,N_8184,N_8736);
nand U15221 (N_15221,N_10471,N_6948);
nor U15222 (N_15222,N_8084,N_9034);
or U15223 (N_15223,N_7593,N_8989);
nand U15224 (N_15224,N_7850,N_12401);
nor U15225 (N_15225,N_8090,N_6630);
nor U15226 (N_15226,N_9130,N_6994);
or U15227 (N_15227,N_12376,N_10375);
and U15228 (N_15228,N_8435,N_11959);
and U15229 (N_15229,N_7981,N_11707);
and U15230 (N_15230,N_7657,N_6408);
nor U15231 (N_15231,N_8386,N_12356);
xnor U15232 (N_15232,N_10659,N_10572);
or U15233 (N_15233,N_9207,N_7510);
or U15234 (N_15234,N_6931,N_7747);
nor U15235 (N_15235,N_12390,N_7754);
nor U15236 (N_15236,N_10395,N_12216);
xnor U15237 (N_15237,N_6383,N_12249);
and U15238 (N_15238,N_7197,N_9937);
and U15239 (N_15239,N_9686,N_7170);
and U15240 (N_15240,N_11660,N_6587);
nor U15241 (N_15241,N_8380,N_8467);
nand U15242 (N_15242,N_10788,N_8742);
nand U15243 (N_15243,N_12322,N_11215);
nand U15244 (N_15244,N_11854,N_9030);
nand U15245 (N_15245,N_10591,N_6619);
and U15246 (N_15246,N_9200,N_10052);
nor U15247 (N_15247,N_8563,N_6925);
and U15248 (N_15248,N_8209,N_11125);
and U15249 (N_15249,N_8003,N_12361);
or U15250 (N_15250,N_6289,N_9913);
or U15251 (N_15251,N_7835,N_10071);
or U15252 (N_15252,N_11363,N_9726);
nand U15253 (N_15253,N_6313,N_10300);
or U15254 (N_15254,N_9391,N_10828);
nand U15255 (N_15255,N_9241,N_7721);
nor U15256 (N_15256,N_8542,N_7214);
and U15257 (N_15257,N_8385,N_8723);
nor U15258 (N_15258,N_7255,N_10896);
or U15259 (N_15259,N_9575,N_11975);
or U15260 (N_15260,N_8812,N_9285);
nor U15261 (N_15261,N_8448,N_10638);
and U15262 (N_15262,N_7049,N_10299);
nor U15263 (N_15263,N_9372,N_8343);
or U15264 (N_15264,N_8526,N_8545);
nand U15265 (N_15265,N_9114,N_7167);
or U15266 (N_15266,N_12131,N_10727);
nand U15267 (N_15267,N_10889,N_8818);
and U15268 (N_15268,N_11456,N_11747);
nor U15269 (N_15269,N_6641,N_11656);
nand U15270 (N_15270,N_9808,N_11381);
and U15271 (N_15271,N_11555,N_6752);
and U15272 (N_15272,N_6887,N_10902);
and U15273 (N_15273,N_11332,N_10379);
nor U15274 (N_15274,N_8160,N_6860);
or U15275 (N_15275,N_8761,N_8277);
nand U15276 (N_15276,N_6341,N_11138);
nand U15277 (N_15277,N_10544,N_11718);
and U15278 (N_15278,N_7278,N_8978);
nor U15279 (N_15279,N_12250,N_11442);
or U15280 (N_15280,N_10843,N_6765);
nand U15281 (N_15281,N_7392,N_7223);
or U15282 (N_15282,N_11101,N_12453);
nor U15283 (N_15283,N_8795,N_12074);
and U15284 (N_15284,N_12409,N_7009);
nand U15285 (N_15285,N_7995,N_8340);
nand U15286 (N_15286,N_8704,N_11924);
nand U15287 (N_15287,N_8981,N_7802);
or U15288 (N_15288,N_9422,N_8452);
and U15289 (N_15289,N_11752,N_7707);
nor U15290 (N_15290,N_11414,N_11159);
nand U15291 (N_15291,N_10153,N_10607);
nor U15292 (N_15292,N_9382,N_8912);
and U15293 (N_15293,N_10505,N_8551);
nor U15294 (N_15294,N_8618,N_11164);
nand U15295 (N_15295,N_10509,N_12267);
and U15296 (N_15296,N_11460,N_6572);
nand U15297 (N_15297,N_9282,N_7914);
and U15298 (N_15298,N_8972,N_12484);
nor U15299 (N_15299,N_12082,N_11483);
or U15300 (N_15300,N_10431,N_8400);
or U15301 (N_15301,N_8250,N_7138);
or U15302 (N_15302,N_7385,N_7854);
or U15303 (N_15303,N_8574,N_7893);
or U15304 (N_15304,N_7647,N_10166);
or U15305 (N_15305,N_11100,N_11954);
nor U15306 (N_15306,N_10860,N_7390);
or U15307 (N_15307,N_8782,N_11675);
nor U15308 (N_15308,N_9452,N_8626);
nor U15309 (N_15309,N_6414,N_7260);
and U15310 (N_15310,N_6585,N_6565);
or U15311 (N_15311,N_7532,N_6564);
nor U15312 (N_15312,N_6508,N_9702);
and U15313 (N_15313,N_10063,N_8305);
nor U15314 (N_15314,N_8824,N_10123);
or U15315 (N_15315,N_9424,N_10724);
nor U15316 (N_15316,N_10031,N_9289);
and U15317 (N_15317,N_11267,N_8032);
and U15318 (N_15318,N_11946,N_11858);
nor U15319 (N_15319,N_12242,N_9093);
or U15320 (N_15320,N_7125,N_9542);
or U15321 (N_15321,N_9089,N_10929);
nor U15322 (N_15322,N_8389,N_9341);
nor U15323 (N_15323,N_12055,N_10645);
nor U15324 (N_15324,N_9643,N_9339);
nor U15325 (N_15325,N_7370,N_7930);
and U15326 (N_15326,N_11070,N_7575);
nand U15327 (N_15327,N_10422,N_8875);
nor U15328 (N_15328,N_10466,N_10856);
nand U15329 (N_15329,N_6905,N_7477);
nand U15330 (N_15330,N_10852,N_11957);
nand U15331 (N_15331,N_8080,N_8607);
and U15332 (N_15332,N_11114,N_8525);
nand U15333 (N_15333,N_6730,N_7123);
nand U15334 (N_15334,N_10330,N_9040);
and U15335 (N_15335,N_11643,N_9744);
or U15336 (N_15336,N_12395,N_8113);
nand U15337 (N_15337,N_11628,N_6286);
nand U15338 (N_15338,N_12042,N_7772);
nand U15339 (N_15339,N_11882,N_9509);
or U15340 (N_15340,N_6790,N_12155);
or U15341 (N_15341,N_7004,N_11334);
or U15342 (N_15342,N_6410,N_12101);
and U15343 (N_15343,N_9067,N_7763);
and U15344 (N_15344,N_12466,N_8362);
and U15345 (N_15345,N_10459,N_12235);
nor U15346 (N_15346,N_8980,N_7760);
nor U15347 (N_15347,N_10758,N_7454);
and U15348 (N_15348,N_7227,N_8436);
and U15349 (N_15349,N_11512,N_7824);
nand U15350 (N_15350,N_10701,N_10973);
nand U15351 (N_15351,N_8732,N_10305);
nor U15352 (N_15352,N_10752,N_11080);
or U15353 (N_15353,N_7470,N_9319);
nand U15354 (N_15354,N_12270,N_7404);
nor U15355 (N_15355,N_9148,N_12179);
and U15356 (N_15356,N_9095,N_8904);
and U15357 (N_15357,N_7944,N_7803);
or U15358 (N_15358,N_8064,N_11287);
nand U15359 (N_15359,N_9896,N_9019);
or U15360 (N_15360,N_12415,N_11426);
or U15361 (N_15361,N_8100,N_8207);
nor U15362 (N_15362,N_12201,N_10516);
nand U15363 (N_15363,N_9212,N_10226);
xor U15364 (N_15364,N_8105,N_12324);
nor U15365 (N_15365,N_7972,N_6525);
and U15366 (N_15366,N_8971,N_7764);
nand U15367 (N_15367,N_6469,N_6461);
nor U15368 (N_15368,N_11735,N_12481);
nor U15369 (N_15369,N_7594,N_10231);
and U15370 (N_15370,N_8460,N_9680);
nand U15371 (N_15371,N_7997,N_9255);
nand U15372 (N_15372,N_8763,N_6456);
nor U15373 (N_15373,N_8914,N_12476);
or U15374 (N_15374,N_7516,N_11182);
or U15375 (N_15375,N_8476,N_9411);
or U15376 (N_15376,N_8955,N_6663);
and U15377 (N_15377,N_9456,N_7766);
or U15378 (N_15378,N_6454,N_9123);
or U15379 (N_15379,N_8897,N_10203);
nor U15380 (N_15380,N_11595,N_11211);
and U15381 (N_15381,N_7250,N_11608);
nor U15382 (N_15382,N_6360,N_12460);
and U15383 (N_15383,N_6435,N_6387);
nand U15384 (N_15384,N_8138,N_7346);
and U15385 (N_15385,N_10448,N_6678);
nor U15386 (N_15386,N_9107,N_11245);
nor U15387 (N_15387,N_9111,N_10951);
and U15388 (N_15388,N_9625,N_9650);
nand U15389 (N_15389,N_10219,N_10974);
nand U15390 (N_15390,N_9875,N_9761);
nand U15391 (N_15391,N_11503,N_6789);
nor U15392 (N_15392,N_12085,N_8046);
nand U15393 (N_15393,N_9590,N_10480);
nand U15394 (N_15394,N_6853,N_9145);
nand U15395 (N_15395,N_9475,N_9676);
and U15396 (N_15396,N_8199,N_10363);
nand U15397 (N_15397,N_7254,N_9552);
nor U15398 (N_15398,N_9910,N_6768);
and U15399 (N_15399,N_11279,N_6448);
and U15400 (N_15400,N_10833,N_8089);
and U15401 (N_15401,N_9629,N_12065);
nor U15402 (N_15402,N_9244,N_7587);
nand U15403 (N_15403,N_12059,N_9732);
or U15404 (N_15404,N_8405,N_8993);
or U15405 (N_15405,N_7465,N_10977);
and U15406 (N_15406,N_9661,N_11394);
or U15407 (N_15407,N_12166,N_9825);
or U15408 (N_15408,N_6382,N_7617);
or U15409 (N_15409,N_6349,N_12190);
and U15410 (N_15410,N_9025,N_11052);
nor U15411 (N_15411,N_7127,N_8592);
nand U15412 (N_15412,N_7374,N_12187);
or U15413 (N_15413,N_10460,N_11395);
and U15414 (N_15414,N_12125,N_11647);
and U15415 (N_15415,N_6807,N_12032);
nor U15416 (N_15416,N_6647,N_8135);
or U15417 (N_15417,N_7489,N_10861);
nand U15418 (N_15418,N_11400,N_6251);
nor U15419 (N_15419,N_12359,N_9792);
or U15420 (N_15420,N_10246,N_12428);
nand U15421 (N_15421,N_7359,N_7394);
nand U15422 (N_15422,N_8087,N_11837);
nor U15423 (N_15423,N_7623,N_6695);
or U15424 (N_15424,N_9517,N_12374);
or U15425 (N_15425,N_6711,N_7499);
and U15426 (N_15426,N_7441,N_10039);
or U15427 (N_15427,N_7706,N_8350);
nand U15428 (N_15428,N_7658,N_10067);
or U15429 (N_15429,N_7783,N_9464);
or U15430 (N_15430,N_12024,N_8002);
nor U15431 (N_15431,N_7917,N_11786);
or U15432 (N_15432,N_7315,N_6715);
and U15433 (N_15433,N_11758,N_10558);
nand U15434 (N_15434,N_10534,N_9831);
and U15435 (N_15435,N_7140,N_9588);
nor U15436 (N_15436,N_10715,N_11286);
and U15437 (N_15437,N_10349,N_11785);
or U15438 (N_15438,N_6689,N_6832);
or U15439 (N_15439,N_7632,N_7327);
and U15440 (N_15440,N_12244,N_8768);
nor U15441 (N_15441,N_11247,N_8733);
or U15442 (N_15442,N_11037,N_11486);
or U15443 (N_15443,N_7949,N_12309);
or U15444 (N_15444,N_12044,N_11049);
nand U15445 (N_15445,N_7141,N_12380);
or U15446 (N_15446,N_9797,N_7736);
and U15447 (N_15447,N_10003,N_10636);
nand U15448 (N_15448,N_12487,N_10523);
nand U15449 (N_15449,N_8238,N_7977);
or U15450 (N_15450,N_11826,N_6838);
and U15451 (N_15451,N_7551,N_7273);
and U15452 (N_15452,N_6316,N_11999);
nand U15453 (N_15453,N_11232,N_11664);
or U15454 (N_15454,N_9936,N_8388);
or U15455 (N_15455,N_12003,N_11285);
or U15456 (N_15456,N_7038,N_6510);
or U15457 (N_15457,N_12116,N_7951);
nor U15458 (N_15458,N_11120,N_8082);
or U15459 (N_15459,N_8431,N_10634);
or U15460 (N_15460,N_10281,N_9665);
nand U15461 (N_15461,N_11178,N_7216);
nor U15462 (N_15462,N_8691,N_8983);
and U15463 (N_15463,N_11401,N_12062);
and U15464 (N_15464,N_8802,N_10423);
and U15465 (N_15465,N_10943,N_10218);
nor U15466 (N_15466,N_6916,N_8347);
and U15467 (N_15467,N_7040,N_7133);
nand U15468 (N_15468,N_8601,N_7596);
nand U15469 (N_15469,N_12181,N_12191);
nor U15470 (N_15470,N_9948,N_11160);
nand U15471 (N_15471,N_9930,N_10043);
or U15472 (N_15472,N_11545,N_7323);
xnor U15473 (N_15473,N_10684,N_6885);
or U15474 (N_15474,N_7017,N_10438);
nor U15475 (N_15475,N_12206,N_6899);
and U15476 (N_15476,N_9147,N_11169);
nand U15477 (N_15477,N_11986,N_9306);
and U15478 (N_15478,N_10401,N_11300);
and U15479 (N_15479,N_6275,N_10381);
nor U15480 (N_15480,N_6699,N_6797);
nor U15481 (N_15481,N_10500,N_7297);
or U15482 (N_15482,N_9325,N_9639);
or U15483 (N_15483,N_11269,N_9278);
nand U15484 (N_15484,N_12224,N_8226);
nand U15485 (N_15485,N_7648,N_10799);
and U15486 (N_15486,N_8020,N_7679);
and U15487 (N_15487,N_10624,N_10669);
nor U15488 (N_15488,N_12434,N_8851);
xnor U15489 (N_15489,N_10185,N_10529);
or U15490 (N_15490,N_7737,N_9938);
nand U15491 (N_15491,N_10621,N_6607);
and U15492 (N_15492,N_9315,N_8700);
and U15493 (N_15493,N_11540,N_11804);
or U15494 (N_15494,N_9904,N_9473);
nand U15495 (N_15495,N_10144,N_7722);
nand U15496 (N_15496,N_7720,N_9637);
nand U15497 (N_15497,N_7771,N_8438);
nand U15498 (N_15498,N_11637,N_8941);
and U15499 (N_15499,N_10311,N_7162);
nor U15500 (N_15500,N_6311,N_9157);
nand U15501 (N_15501,N_10417,N_9606);
nand U15502 (N_15502,N_7074,N_10859);
nor U15503 (N_15503,N_10567,N_7268);
nor U15504 (N_15504,N_7097,N_11003);
nor U15505 (N_15505,N_7295,N_10588);
xor U15506 (N_15506,N_9068,N_9012);
nor U15507 (N_15507,N_7793,N_7488);
or U15508 (N_15508,N_6511,N_7129);
nor U15509 (N_15509,N_6338,N_9544);
nor U15510 (N_15510,N_7788,N_9798);
and U15511 (N_15511,N_9393,N_12163);
or U15512 (N_15512,N_8224,N_11877);
nand U15513 (N_15513,N_6736,N_8365);
and U15514 (N_15514,N_6844,N_8088);
nor U15515 (N_15515,N_10653,N_12396);
nor U15516 (N_15516,N_8571,N_10483);
nand U15517 (N_15517,N_10263,N_6325);
or U15518 (N_15518,N_11638,N_8934);
or U15519 (N_15519,N_11831,N_9752);
nand U15520 (N_15520,N_7458,N_8447);
or U15521 (N_15521,N_6676,N_7451);
nor U15522 (N_15522,N_11623,N_11007);
or U15523 (N_15523,N_9014,N_8114);
and U15524 (N_15524,N_11265,N_9634);
nand U15525 (N_15525,N_7137,N_8514);
or U15526 (N_15526,N_6623,N_12007);
nand U15527 (N_15527,N_10341,N_7553);
or U15528 (N_15528,N_8155,N_7328);
nor U15529 (N_15529,N_7120,N_12124);
and U15530 (N_15530,N_7008,N_8387);
nor U15531 (N_15531,N_8314,N_6513);
or U15532 (N_15532,N_10697,N_12180);
nand U15533 (N_15533,N_11257,N_7809);
or U15534 (N_15534,N_7224,N_9133);
nand U15535 (N_15535,N_7814,N_7405);
nor U15536 (N_15536,N_9094,N_10763);
nand U15537 (N_15537,N_11271,N_8655);
or U15538 (N_15538,N_11291,N_8061);
xnor U15539 (N_15539,N_8992,N_11905);
and U15540 (N_15540,N_9164,N_7158);
nand U15541 (N_15541,N_9574,N_7769);
or U15542 (N_15542,N_12432,N_8999);
nand U15543 (N_15543,N_11190,N_7212);
or U15544 (N_15544,N_6743,N_11898);
nand U15545 (N_15545,N_7045,N_11610);
nor U15546 (N_15546,N_10983,N_11709);
and U15547 (N_15547,N_8951,N_6624);
and U15548 (N_15548,N_7902,N_6841);
nor U15549 (N_15549,N_6617,N_11848);
and U15550 (N_15550,N_12377,N_7019);
nand U15551 (N_15551,N_10079,N_8666);
and U15552 (N_15552,N_8007,N_8378);
and U15553 (N_15553,N_7919,N_11528);
or U15554 (N_15554,N_10325,N_6999);
and U15555 (N_15555,N_9963,N_11333);
nor U15556 (N_15556,N_6401,N_8615);
or U15557 (N_15557,N_8423,N_8151);
or U15558 (N_15558,N_10352,N_10781);
or U15559 (N_15559,N_12403,N_12496);
or U15560 (N_15560,N_7280,N_9619);
nor U15561 (N_15561,N_6309,N_9764);
nor U15562 (N_15562,N_8498,N_11193);
nor U15563 (N_15563,N_7015,N_7538);
nor U15564 (N_15564,N_7270,N_7500);
nor U15565 (N_15565,N_11841,N_10442);
nand U15566 (N_15566,N_8342,N_9346);
or U15567 (N_15567,N_10549,N_9760);
nor U15568 (N_15568,N_11236,N_8888);
and U15569 (N_15569,N_8878,N_9901);
or U15570 (N_15570,N_12421,N_12343);
or U15571 (N_15571,N_10832,N_6631);
nand U15572 (N_15572,N_9607,N_8586);
nand U15573 (N_15573,N_7561,N_8260);
nand U15574 (N_15574,N_8309,N_9826);
nor U15575 (N_15575,N_7869,N_9688);
and U15576 (N_15576,N_12142,N_10552);
or U15577 (N_15577,N_7288,N_6467);
or U15578 (N_15578,N_8013,N_6514);
or U15579 (N_15579,N_11261,N_11366);
or U15580 (N_15580,N_10162,N_6814);
and U15581 (N_15581,N_9342,N_12161);
or U15582 (N_15582,N_12469,N_6602);
nor U15583 (N_15583,N_8703,N_9770);
or U15584 (N_15584,N_8701,N_11134);
or U15585 (N_15585,N_9401,N_10966);
and U15586 (N_15586,N_11467,N_11237);
or U15587 (N_15587,N_9024,N_6579);
nand U15588 (N_15588,N_8952,N_10058);
and U15589 (N_15589,N_9900,N_10775);
and U15590 (N_15590,N_12444,N_8541);
nor U15591 (N_15591,N_11755,N_11104);
nor U15592 (N_15592,N_9867,N_12472);
and U15593 (N_15593,N_9587,N_11121);
nor U15594 (N_15594,N_11449,N_8401);
nand U15595 (N_15595,N_7302,N_6334);
nand U15596 (N_15596,N_7121,N_7024);
or U15597 (N_15597,N_7805,N_6477);
or U15598 (N_15598,N_11649,N_8341);
or U15599 (N_15599,N_9603,N_6266);
nor U15600 (N_15600,N_7413,N_11033);
and U15601 (N_15601,N_11144,N_8985);
or U15602 (N_15602,N_6529,N_12162);
and U15603 (N_15603,N_8474,N_9032);
or U15604 (N_15604,N_7360,N_7508);
nand U15605 (N_15605,N_10434,N_9235);
and U15606 (N_15606,N_7403,N_10911);
and U15607 (N_15607,N_8928,N_7872);
and U15608 (N_15608,N_7582,N_8817);
nand U15609 (N_15609,N_9449,N_7082);
nor U15610 (N_15610,N_6888,N_11377);
and U15611 (N_15611,N_8849,N_7200);
or U15612 (N_15612,N_9334,N_10302);
xnor U15613 (N_15613,N_8395,N_7604);
nand U15614 (N_15614,N_10810,N_6740);
nand U15615 (N_15615,N_9399,N_9186);
and U15616 (N_15616,N_7546,N_8471);
nor U15617 (N_15617,N_9868,N_12240);
nor U15618 (N_15618,N_11418,N_12169);
nor U15619 (N_15619,N_12188,N_9615);
or U15620 (N_15620,N_12000,N_12422);
nor U15621 (N_15621,N_10590,N_12268);
and U15622 (N_15622,N_8859,N_8413);
nor U15623 (N_15623,N_11775,N_6756);
nand U15624 (N_15624,N_8321,N_9675);
and U15625 (N_15625,N_6425,N_6293);
and U15626 (N_15626,N_6529,N_11148);
nand U15627 (N_15627,N_11375,N_7766);
or U15628 (N_15628,N_11206,N_6882);
and U15629 (N_15629,N_11747,N_6365);
nor U15630 (N_15630,N_10384,N_8520);
nand U15631 (N_15631,N_7444,N_7525);
or U15632 (N_15632,N_6827,N_8078);
nor U15633 (N_15633,N_8883,N_11928);
or U15634 (N_15634,N_6943,N_6433);
nor U15635 (N_15635,N_7877,N_8747);
nor U15636 (N_15636,N_10330,N_12376);
and U15637 (N_15637,N_7089,N_7258);
and U15638 (N_15638,N_9890,N_6636);
and U15639 (N_15639,N_11212,N_10782);
or U15640 (N_15640,N_9468,N_8235);
and U15641 (N_15641,N_10439,N_11337);
nand U15642 (N_15642,N_8153,N_6671);
or U15643 (N_15643,N_9750,N_12271);
and U15644 (N_15644,N_12483,N_9172);
nor U15645 (N_15645,N_9599,N_6890);
nor U15646 (N_15646,N_12346,N_7012);
nand U15647 (N_15647,N_11836,N_8147);
nor U15648 (N_15648,N_8556,N_10357);
and U15649 (N_15649,N_7419,N_10780);
or U15650 (N_15650,N_11820,N_9597);
and U15651 (N_15651,N_11586,N_12073);
nand U15652 (N_15652,N_12124,N_10057);
nand U15653 (N_15653,N_7516,N_8658);
nor U15654 (N_15654,N_12112,N_12293);
and U15655 (N_15655,N_6366,N_7055);
or U15656 (N_15656,N_6839,N_12048);
or U15657 (N_15657,N_9206,N_9363);
nor U15658 (N_15658,N_11976,N_8050);
nand U15659 (N_15659,N_11209,N_11390);
nand U15660 (N_15660,N_10942,N_11875);
or U15661 (N_15661,N_7689,N_8234);
and U15662 (N_15662,N_11447,N_9398);
nor U15663 (N_15663,N_6820,N_10125);
and U15664 (N_15664,N_7594,N_7918);
nor U15665 (N_15665,N_10510,N_6345);
and U15666 (N_15666,N_10333,N_12320);
nor U15667 (N_15667,N_12438,N_9883);
nand U15668 (N_15668,N_9444,N_8921);
or U15669 (N_15669,N_7791,N_8813);
nand U15670 (N_15670,N_8066,N_11214);
or U15671 (N_15671,N_11667,N_12150);
or U15672 (N_15672,N_10003,N_9806);
or U15673 (N_15673,N_9950,N_7092);
nand U15674 (N_15674,N_8253,N_9190);
nor U15675 (N_15675,N_11897,N_10197);
or U15676 (N_15676,N_9205,N_8428);
or U15677 (N_15677,N_7627,N_8237);
or U15678 (N_15678,N_10121,N_9118);
nor U15679 (N_15679,N_6355,N_6683);
or U15680 (N_15680,N_7687,N_10941);
nor U15681 (N_15681,N_9273,N_7369);
nand U15682 (N_15682,N_10922,N_9059);
nand U15683 (N_15683,N_9010,N_9508);
or U15684 (N_15684,N_11344,N_11901);
and U15685 (N_15685,N_10179,N_8151);
nor U15686 (N_15686,N_7175,N_10807);
nand U15687 (N_15687,N_9805,N_10304);
nor U15688 (N_15688,N_10595,N_11798);
nor U15689 (N_15689,N_6825,N_9480);
or U15690 (N_15690,N_8636,N_10998);
nor U15691 (N_15691,N_9013,N_9190);
nor U15692 (N_15692,N_8189,N_8668);
nor U15693 (N_15693,N_7184,N_10252);
nor U15694 (N_15694,N_6514,N_9255);
nor U15695 (N_15695,N_8857,N_11177);
or U15696 (N_15696,N_10844,N_6282);
or U15697 (N_15697,N_10278,N_12166);
and U15698 (N_15698,N_9166,N_6330);
or U15699 (N_15699,N_8884,N_8409);
nand U15700 (N_15700,N_6990,N_7146);
nand U15701 (N_15701,N_11570,N_11419);
nand U15702 (N_15702,N_11958,N_12306);
or U15703 (N_15703,N_8802,N_8765);
and U15704 (N_15704,N_12266,N_9508);
nor U15705 (N_15705,N_7304,N_7009);
nand U15706 (N_15706,N_6653,N_9757);
or U15707 (N_15707,N_8434,N_6965);
or U15708 (N_15708,N_10406,N_10166);
or U15709 (N_15709,N_7057,N_10451);
nor U15710 (N_15710,N_7658,N_8002);
nor U15711 (N_15711,N_7222,N_6297);
nor U15712 (N_15712,N_6795,N_8113);
or U15713 (N_15713,N_7436,N_9712);
nor U15714 (N_15714,N_12060,N_6654);
and U15715 (N_15715,N_7424,N_10979);
and U15716 (N_15716,N_7827,N_9386);
nor U15717 (N_15717,N_7693,N_10515);
nand U15718 (N_15718,N_9425,N_11166);
or U15719 (N_15719,N_7789,N_10324);
nand U15720 (N_15720,N_6699,N_11338);
and U15721 (N_15721,N_11206,N_11071);
nor U15722 (N_15722,N_7756,N_10508);
nand U15723 (N_15723,N_10084,N_7732);
nand U15724 (N_15724,N_8333,N_10111);
nand U15725 (N_15725,N_7373,N_11146);
or U15726 (N_15726,N_7448,N_8261);
nand U15727 (N_15727,N_6545,N_12097);
nor U15728 (N_15728,N_10208,N_11952);
and U15729 (N_15729,N_9342,N_9762);
nand U15730 (N_15730,N_6298,N_7100);
nor U15731 (N_15731,N_8854,N_8320);
or U15732 (N_15732,N_11785,N_7541);
nor U15733 (N_15733,N_11808,N_11177);
or U15734 (N_15734,N_7724,N_7343);
and U15735 (N_15735,N_9186,N_10026);
and U15736 (N_15736,N_6297,N_7624);
nor U15737 (N_15737,N_9819,N_12421);
or U15738 (N_15738,N_9302,N_7842);
nand U15739 (N_15739,N_10190,N_8495);
nand U15740 (N_15740,N_10271,N_6698);
or U15741 (N_15741,N_7425,N_8203);
nand U15742 (N_15742,N_6362,N_10351);
or U15743 (N_15743,N_8905,N_9144);
and U15744 (N_15744,N_10503,N_9140);
nor U15745 (N_15745,N_7068,N_10840);
nor U15746 (N_15746,N_12213,N_8745);
nand U15747 (N_15747,N_9706,N_10994);
and U15748 (N_15748,N_9884,N_8649);
nor U15749 (N_15749,N_9941,N_8141);
and U15750 (N_15750,N_8960,N_12164);
nand U15751 (N_15751,N_6579,N_10199);
nand U15752 (N_15752,N_10968,N_10417);
or U15753 (N_15753,N_8684,N_6884);
nand U15754 (N_15754,N_6394,N_11645);
nor U15755 (N_15755,N_10736,N_6909);
nor U15756 (N_15756,N_6293,N_6587);
nor U15757 (N_15757,N_11939,N_8985);
nand U15758 (N_15758,N_12024,N_10797);
or U15759 (N_15759,N_8310,N_11771);
and U15760 (N_15760,N_10139,N_7677);
and U15761 (N_15761,N_7303,N_12083);
nand U15762 (N_15762,N_9673,N_11961);
nand U15763 (N_15763,N_11627,N_12116);
or U15764 (N_15764,N_9414,N_12342);
nand U15765 (N_15765,N_8701,N_12027);
nand U15766 (N_15766,N_8208,N_9557);
nor U15767 (N_15767,N_8681,N_11890);
and U15768 (N_15768,N_7383,N_6690);
and U15769 (N_15769,N_10126,N_6358);
and U15770 (N_15770,N_12248,N_8692);
or U15771 (N_15771,N_9012,N_7716);
nand U15772 (N_15772,N_11416,N_9247);
or U15773 (N_15773,N_9078,N_9089);
nor U15774 (N_15774,N_10591,N_6707);
nand U15775 (N_15775,N_6836,N_10223);
nand U15776 (N_15776,N_9899,N_6567);
nand U15777 (N_15777,N_8315,N_8261);
and U15778 (N_15778,N_10961,N_9566);
nor U15779 (N_15779,N_9631,N_6939);
or U15780 (N_15780,N_7647,N_7197);
nand U15781 (N_15781,N_7180,N_12300);
nor U15782 (N_15782,N_10463,N_11238);
or U15783 (N_15783,N_10775,N_8482);
nand U15784 (N_15784,N_7228,N_10432);
or U15785 (N_15785,N_7326,N_11608);
and U15786 (N_15786,N_7561,N_7048);
nor U15787 (N_15787,N_10587,N_10076);
nand U15788 (N_15788,N_9328,N_11546);
nor U15789 (N_15789,N_7815,N_11871);
and U15790 (N_15790,N_9347,N_10592);
nand U15791 (N_15791,N_11266,N_10004);
or U15792 (N_15792,N_11312,N_6538);
nor U15793 (N_15793,N_8149,N_7711);
nand U15794 (N_15794,N_9691,N_8419);
nor U15795 (N_15795,N_9106,N_6861);
nor U15796 (N_15796,N_11196,N_10026);
or U15797 (N_15797,N_12165,N_7951);
nor U15798 (N_15798,N_11774,N_6409);
nor U15799 (N_15799,N_8001,N_11714);
nand U15800 (N_15800,N_6368,N_9767);
nand U15801 (N_15801,N_10154,N_10585);
or U15802 (N_15802,N_9252,N_6314);
nor U15803 (N_15803,N_9377,N_12094);
nor U15804 (N_15804,N_11287,N_12373);
and U15805 (N_15805,N_11209,N_12089);
nand U15806 (N_15806,N_8711,N_9881);
nor U15807 (N_15807,N_9552,N_10774);
nor U15808 (N_15808,N_11641,N_11219);
or U15809 (N_15809,N_6735,N_9587);
nand U15810 (N_15810,N_7975,N_7803);
or U15811 (N_15811,N_11543,N_9521);
or U15812 (N_15812,N_8655,N_8432);
and U15813 (N_15813,N_11284,N_12288);
nor U15814 (N_15814,N_8766,N_8690);
and U15815 (N_15815,N_7681,N_7411);
nor U15816 (N_15816,N_6736,N_6742);
nand U15817 (N_15817,N_7492,N_12017);
or U15818 (N_15818,N_9471,N_8776);
or U15819 (N_15819,N_11224,N_10954);
nor U15820 (N_15820,N_11766,N_11772);
nand U15821 (N_15821,N_6396,N_8486);
nand U15822 (N_15822,N_12218,N_6325);
nand U15823 (N_15823,N_11500,N_8769);
and U15824 (N_15824,N_11206,N_7130);
nor U15825 (N_15825,N_9804,N_9977);
and U15826 (N_15826,N_8004,N_11709);
nor U15827 (N_15827,N_8264,N_12315);
nor U15828 (N_15828,N_6264,N_11151);
nand U15829 (N_15829,N_9659,N_11125);
nand U15830 (N_15830,N_8460,N_9544);
nand U15831 (N_15831,N_7097,N_6961);
and U15832 (N_15832,N_12332,N_7245);
nor U15833 (N_15833,N_12172,N_10801);
nand U15834 (N_15834,N_8375,N_11730);
nor U15835 (N_15835,N_10492,N_7950);
nor U15836 (N_15836,N_10655,N_10198);
and U15837 (N_15837,N_9665,N_6552);
nand U15838 (N_15838,N_7463,N_10506);
or U15839 (N_15839,N_8909,N_9040);
nor U15840 (N_15840,N_11728,N_11875);
nand U15841 (N_15841,N_11433,N_12336);
nand U15842 (N_15842,N_11898,N_7043);
or U15843 (N_15843,N_7186,N_8341);
nor U15844 (N_15844,N_10307,N_8867);
or U15845 (N_15845,N_11283,N_10127);
or U15846 (N_15846,N_11101,N_10984);
nor U15847 (N_15847,N_7800,N_10242);
nand U15848 (N_15848,N_8510,N_10286);
and U15849 (N_15849,N_8104,N_8460);
nand U15850 (N_15850,N_9877,N_12043);
or U15851 (N_15851,N_10875,N_8034);
nand U15852 (N_15852,N_8091,N_10519);
and U15853 (N_15853,N_9539,N_11849);
nand U15854 (N_15854,N_8901,N_8908);
and U15855 (N_15855,N_9136,N_12362);
or U15856 (N_15856,N_11899,N_10928);
or U15857 (N_15857,N_11146,N_11662);
nor U15858 (N_15858,N_9821,N_9434);
nand U15859 (N_15859,N_11785,N_10601);
nor U15860 (N_15860,N_9521,N_11132);
or U15861 (N_15861,N_10848,N_7090);
and U15862 (N_15862,N_6480,N_9088);
or U15863 (N_15863,N_8327,N_6921);
xnor U15864 (N_15864,N_10455,N_6417);
nand U15865 (N_15865,N_10551,N_11788);
nor U15866 (N_15866,N_9092,N_8004);
and U15867 (N_15867,N_9982,N_9062);
nand U15868 (N_15868,N_9421,N_11451);
nand U15869 (N_15869,N_11837,N_10349);
and U15870 (N_15870,N_10340,N_10197);
nand U15871 (N_15871,N_10262,N_6779);
or U15872 (N_15872,N_8506,N_9606);
and U15873 (N_15873,N_9973,N_11588);
and U15874 (N_15874,N_7896,N_9520);
nand U15875 (N_15875,N_12407,N_11742);
and U15876 (N_15876,N_7052,N_10482);
and U15877 (N_15877,N_10374,N_9503);
or U15878 (N_15878,N_8001,N_8576);
or U15879 (N_15879,N_7693,N_9639);
and U15880 (N_15880,N_9343,N_6752);
or U15881 (N_15881,N_10174,N_9808);
or U15882 (N_15882,N_12457,N_11379);
and U15883 (N_15883,N_6294,N_10794);
nor U15884 (N_15884,N_8339,N_11850);
and U15885 (N_15885,N_7732,N_9020);
nor U15886 (N_15886,N_7874,N_12216);
and U15887 (N_15887,N_6508,N_9543);
nand U15888 (N_15888,N_11366,N_12351);
or U15889 (N_15889,N_11406,N_6827);
nor U15890 (N_15890,N_12388,N_11974);
or U15891 (N_15891,N_12119,N_11042);
nand U15892 (N_15892,N_10459,N_10705);
or U15893 (N_15893,N_10005,N_11771);
and U15894 (N_15894,N_9681,N_7788);
and U15895 (N_15895,N_12364,N_7151);
and U15896 (N_15896,N_7489,N_8347);
and U15897 (N_15897,N_10969,N_12085);
nor U15898 (N_15898,N_7500,N_10781);
or U15899 (N_15899,N_9511,N_10322);
or U15900 (N_15900,N_9063,N_10635);
or U15901 (N_15901,N_10649,N_9324);
nand U15902 (N_15902,N_8742,N_6423);
and U15903 (N_15903,N_8216,N_10568);
nor U15904 (N_15904,N_6765,N_9376);
nand U15905 (N_15905,N_11123,N_9254);
or U15906 (N_15906,N_11342,N_12278);
nor U15907 (N_15907,N_10160,N_6533);
nor U15908 (N_15908,N_9882,N_6908);
nand U15909 (N_15909,N_7778,N_8757);
nor U15910 (N_15910,N_8746,N_8254);
nor U15911 (N_15911,N_7968,N_10727);
and U15912 (N_15912,N_11601,N_8611);
nor U15913 (N_15913,N_8212,N_7403);
or U15914 (N_15914,N_11476,N_7958);
nand U15915 (N_15915,N_6738,N_6858);
nor U15916 (N_15916,N_10920,N_10026);
or U15917 (N_15917,N_11916,N_12156);
and U15918 (N_15918,N_11215,N_11432);
or U15919 (N_15919,N_8926,N_11792);
or U15920 (N_15920,N_10327,N_10287);
nand U15921 (N_15921,N_7253,N_10562);
nor U15922 (N_15922,N_9374,N_10892);
nor U15923 (N_15923,N_7416,N_6257);
nor U15924 (N_15924,N_9882,N_6522);
nor U15925 (N_15925,N_9284,N_6544);
and U15926 (N_15926,N_7096,N_11859);
nand U15927 (N_15927,N_10644,N_7983);
nor U15928 (N_15928,N_9874,N_10589);
or U15929 (N_15929,N_11221,N_9629);
or U15930 (N_15930,N_9814,N_7271);
and U15931 (N_15931,N_9427,N_8017);
nor U15932 (N_15932,N_9174,N_11768);
nand U15933 (N_15933,N_6551,N_7165);
and U15934 (N_15934,N_9410,N_10381);
nand U15935 (N_15935,N_11040,N_6428);
nand U15936 (N_15936,N_11257,N_11571);
nand U15937 (N_15937,N_8642,N_9672);
nand U15938 (N_15938,N_10473,N_7598);
and U15939 (N_15939,N_10536,N_11536);
or U15940 (N_15940,N_7919,N_7790);
and U15941 (N_15941,N_7466,N_10327);
and U15942 (N_15942,N_8484,N_7289);
nor U15943 (N_15943,N_11757,N_11458);
nor U15944 (N_15944,N_12257,N_11829);
nor U15945 (N_15945,N_9618,N_7068);
nand U15946 (N_15946,N_11345,N_7046);
nand U15947 (N_15947,N_6431,N_9805);
nor U15948 (N_15948,N_11714,N_9340);
or U15949 (N_15949,N_9075,N_7546);
nor U15950 (N_15950,N_8330,N_11428);
nor U15951 (N_15951,N_12099,N_7337);
nor U15952 (N_15952,N_10884,N_7098);
nor U15953 (N_15953,N_9620,N_10999);
nor U15954 (N_15954,N_6787,N_12031);
nand U15955 (N_15955,N_9778,N_10960);
or U15956 (N_15956,N_8347,N_11951);
nor U15957 (N_15957,N_12093,N_11753);
nor U15958 (N_15958,N_11475,N_9249);
and U15959 (N_15959,N_11163,N_7165);
nor U15960 (N_15960,N_8530,N_12322);
nand U15961 (N_15961,N_10643,N_8360);
nor U15962 (N_15962,N_11058,N_6662);
nor U15963 (N_15963,N_8940,N_11038);
nor U15964 (N_15964,N_7097,N_9229);
nand U15965 (N_15965,N_7176,N_8203);
nor U15966 (N_15966,N_8579,N_8598);
nor U15967 (N_15967,N_7166,N_9628);
nand U15968 (N_15968,N_8290,N_11555);
or U15969 (N_15969,N_6819,N_9395);
nor U15970 (N_15970,N_8563,N_9072);
nor U15971 (N_15971,N_7674,N_10911);
nand U15972 (N_15972,N_11289,N_11755);
nor U15973 (N_15973,N_7416,N_10067);
nor U15974 (N_15974,N_11122,N_8483);
nand U15975 (N_15975,N_7606,N_8410);
and U15976 (N_15976,N_9322,N_9794);
or U15977 (N_15977,N_10818,N_11471);
or U15978 (N_15978,N_11554,N_9828);
nor U15979 (N_15979,N_7260,N_8777);
and U15980 (N_15980,N_11623,N_11655);
or U15981 (N_15981,N_9597,N_9427);
nor U15982 (N_15982,N_6642,N_9799);
nand U15983 (N_15983,N_9923,N_11541);
nor U15984 (N_15984,N_9549,N_8139);
and U15985 (N_15985,N_11033,N_7930);
nand U15986 (N_15986,N_9914,N_12334);
or U15987 (N_15987,N_11265,N_8829);
or U15988 (N_15988,N_11536,N_11421);
nand U15989 (N_15989,N_9662,N_10020);
or U15990 (N_15990,N_12467,N_8102);
nor U15991 (N_15991,N_11353,N_8685);
nand U15992 (N_15992,N_11594,N_11629);
or U15993 (N_15993,N_10989,N_11915);
or U15994 (N_15994,N_7508,N_7363);
or U15995 (N_15995,N_8559,N_10931);
nand U15996 (N_15996,N_10070,N_8024);
nand U15997 (N_15997,N_10548,N_6572);
nor U15998 (N_15998,N_6565,N_11062);
and U15999 (N_15999,N_10082,N_11788);
or U16000 (N_16000,N_12155,N_11481);
and U16001 (N_16001,N_6930,N_7176);
nor U16002 (N_16002,N_11013,N_9190);
nand U16003 (N_16003,N_7679,N_7579);
and U16004 (N_16004,N_12132,N_9385);
xnor U16005 (N_16005,N_11097,N_9180);
and U16006 (N_16006,N_6654,N_11539);
and U16007 (N_16007,N_9827,N_10328);
and U16008 (N_16008,N_8816,N_9416);
and U16009 (N_16009,N_10611,N_11337);
nor U16010 (N_16010,N_11306,N_11906);
nand U16011 (N_16011,N_12359,N_10800);
nand U16012 (N_16012,N_7750,N_8752);
nor U16013 (N_16013,N_7151,N_9587);
or U16014 (N_16014,N_10394,N_6834);
or U16015 (N_16015,N_9982,N_9746);
or U16016 (N_16016,N_7572,N_6492);
nand U16017 (N_16017,N_11507,N_11179);
and U16018 (N_16018,N_10352,N_9043);
and U16019 (N_16019,N_8883,N_8168);
nor U16020 (N_16020,N_8421,N_10664);
nor U16021 (N_16021,N_9168,N_11083);
nor U16022 (N_16022,N_6329,N_9675);
or U16023 (N_16023,N_8927,N_10319);
and U16024 (N_16024,N_10487,N_6555);
nor U16025 (N_16025,N_8144,N_7064);
nand U16026 (N_16026,N_6835,N_9576);
and U16027 (N_16027,N_10589,N_7470);
or U16028 (N_16028,N_8960,N_8299);
or U16029 (N_16029,N_8083,N_6906);
and U16030 (N_16030,N_11521,N_10673);
or U16031 (N_16031,N_11803,N_8481);
nor U16032 (N_16032,N_10681,N_6312);
nor U16033 (N_16033,N_9109,N_7079);
or U16034 (N_16034,N_9302,N_7278);
nand U16035 (N_16035,N_7598,N_8716);
or U16036 (N_16036,N_12381,N_10630);
and U16037 (N_16037,N_8694,N_6500);
or U16038 (N_16038,N_10358,N_10277);
or U16039 (N_16039,N_7327,N_10586);
and U16040 (N_16040,N_7258,N_12274);
nand U16041 (N_16041,N_9728,N_8617);
nand U16042 (N_16042,N_11941,N_7556);
nand U16043 (N_16043,N_7040,N_7933);
nand U16044 (N_16044,N_8294,N_6816);
nor U16045 (N_16045,N_11477,N_10434);
nor U16046 (N_16046,N_9762,N_7207);
and U16047 (N_16047,N_8272,N_10849);
nor U16048 (N_16048,N_12294,N_8966);
nor U16049 (N_16049,N_9568,N_8433);
nand U16050 (N_16050,N_11161,N_8754);
nand U16051 (N_16051,N_7893,N_7172);
or U16052 (N_16052,N_10144,N_7122);
and U16053 (N_16053,N_12365,N_9784);
nand U16054 (N_16054,N_6362,N_6639);
or U16055 (N_16055,N_7527,N_10133);
and U16056 (N_16056,N_11851,N_9603);
or U16057 (N_16057,N_6996,N_8284);
xor U16058 (N_16058,N_10128,N_11196);
or U16059 (N_16059,N_9052,N_9583);
nand U16060 (N_16060,N_6436,N_7453);
nand U16061 (N_16061,N_7196,N_10474);
and U16062 (N_16062,N_12169,N_10176);
nand U16063 (N_16063,N_10430,N_11961);
nor U16064 (N_16064,N_11372,N_10770);
or U16065 (N_16065,N_9350,N_9869);
nand U16066 (N_16066,N_11226,N_7318);
nand U16067 (N_16067,N_7344,N_6369);
or U16068 (N_16068,N_7056,N_10358);
nand U16069 (N_16069,N_10710,N_10735);
nand U16070 (N_16070,N_10530,N_12499);
nand U16071 (N_16071,N_10108,N_11302);
nand U16072 (N_16072,N_11448,N_7202);
and U16073 (N_16073,N_8731,N_11240);
and U16074 (N_16074,N_10403,N_11391);
nor U16075 (N_16075,N_10678,N_10819);
and U16076 (N_16076,N_9191,N_11394);
nor U16077 (N_16077,N_6441,N_9773);
or U16078 (N_16078,N_9819,N_10593);
nor U16079 (N_16079,N_10662,N_12007);
nor U16080 (N_16080,N_8473,N_8988);
nor U16081 (N_16081,N_7968,N_11543);
and U16082 (N_16082,N_7124,N_11529);
and U16083 (N_16083,N_8206,N_7342);
nor U16084 (N_16084,N_9131,N_8804);
nor U16085 (N_16085,N_9610,N_11759);
or U16086 (N_16086,N_6309,N_6278);
and U16087 (N_16087,N_12175,N_10465);
nor U16088 (N_16088,N_10900,N_10816);
or U16089 (N_16089,N_12410,N_10200);
nor U16090 (N_16090,N_7142,N_11054);
nand U16091 (N_16091,N_6944,N_9681);
and U16092 (N_16092,N_7405,N_12155);
nor U16093 (N_16093,N_6352,N_9001);
nand U16094 (N_16094,N_11074,N_7780);
nor U16095 (N_16095,N_10435,N_10087);
nand U16096 (N_16096,N_6685,N_10694);
or U16097 (N_16097,N_10012,N_9802);
or U16098 (N_16098,N_6863,N_10073);
or U16099 (N_16099,N_7867,N_11799);
nand U16100 (N_16100,N_12483,N_6886);
nor U16101 (N_16101,N_10611,N_6590);
nand U16102 (N_16102,N_6883,N_11039);
nor U16103 (N_16103,N_9522,N_11342);
or U16104 (N_16104,N_7926,N_10012);
nand U16105 (N_16105,N_10416,N_10177);
nand U16106 (N_16106,N_9215,N_7108);
nor U16107 (N_16107,N_9680,N_10968);
nand U16108 (N_16108,N_9506,N_9570);
nor U16109 (N_16109,N_10749,N_9489);
nand U16110 (N_16110,N_7722,N_9305);
nand U16111 (N_16111,N_6805,N_11391);
nand U16112 (N_16112,N_11494,N_9651);
nand U16113 (N_16113,N_9611,N_7499);
nor U16114 (N_16114,N_6257,N_11084);
nor U16115 (N_16115,N_10432,N_10573);
nor U16116 (N_16116,N_8810,N_6728);
nor U16117 (N_16117,N_9013,N_8252);
nor U16118 (N_16118,N_10013,N_10537);
or U16119 (N_16119,N_10284,N_8211);
or U16120 (N_16120,N_7195,N_10297);
xor U16121 (N_16121,N_10112,N_7121);
and U16122 (N_16122,N_11395,N_7828);
nand U16123 (N_16123,N_6937,N_9813);
nor U16124 (N_16124,N_7461,N_7797);
nor U16125 (N_16125,N_10672,N_11724);
nor U16126 (N_16126,N_11004,N_7637);
nand U16127 (N_16127,N_11245,N_10234);
and U16128 (N_16128,N_9594,N_11407);
nand U16129 (N_16129,N_7222,N_7540);
and U16130 (N_16130,N_6393,N_6482);
or U16131 (N_16131,N_7703,N_9098);
nor U16132 (N_16132,N_11295,N_9586);
nor U16133 (N_16133,N_8634,N_12474);
nor U16134 (N_16134,N_6529,N_12312);
nor U16135 (N_16135,N_11223,N_7081);
or U16136 (N_16136,N_11726,N_6764);
nand U16137 (N_16137,N_10993,N_9684);
and U16138 (N_16138,N_7573,N_9000);
nand U16139 (N_16139,N_10878,N_6583);
nand U16140 (N_16140,N_7973,N_9731);
and U16141 (N_16141,N_9623,N_10157);
or U16142 (N_16142,N_9589,N_10840);
and U16143 (N_16143,N_11942,N_6861);
and U16144 (N_16144,N_8534,N_7450);
or U16145 (N_16145,N_7723,N_7784);
or U16146 (N_16146,N_9319,N_7282);
nor U16147 (N_16147,N_7001,N_8359);
nor U16148 (N_16148,N_9957,N_9538);
or U16149 (N_16149,N_7259,N_8479);
or U16150 (N_16150,N_9768,N_11538);
and U16151 (N_16151,N_10049,N_9977);
and U16152 (N_16152,N_10115,N_6716);
and U16153 (N_16153,N_6523,N_12455);
or U16154 (N_16154,N_7499,N_8427);
nor U16155 (N_16155,N_6638,N_10286);
or U16156 (N_16156,N_8830,N_11105);
or U16157 (N_16157,N_7934,N_6770);
or U16158 (N_16158,N_7017,N_11347);
or U16159 (N_16159,N_7111,N_10201);
nor U16160 (N_16160,N_6659,N_9024);
and U16161 (N_16161,N_8145,N_11310);
nand U16162 (N_16162,N_11381,N_8231);
and U16163 (N_16163,N_10185,N_11053);
or U16164 (N_16164,N_7353,N_6522);
and U16165 (N_16165,N_11351,N_9790);
nand U16166 (N_16166,N_7689,N_8843);
nor U16167 (N_16167,N_8957,N_11371);
nor U16168 (N_16168,N_10462,N_11834);
nand U16169 (N_16169,N_8852,N_11178);
nand U16170 (N_16170,N_6259,N_7370);
nand U16171 (N_16171,N_10018,N_8820);
and U16172 (N_16172,N_10937,N_10327);
nand U16173 (N_16173,N_10445,N_10793);
nand U16174 (N_16174,N_11178,N_12278);
nand U16175 (N_16175,N_9435,N_11922);
or U16176 (N_16176,N_11413,N_12252);
nand U16177 (N_16177,N_7184,N_8656);
nor U16178 (N_16178,N_11198,N_8472);
and U16179 (N_16179,N_11822,N_6818);
nand U16180 (N_16180,N_8220,N_7025);
nor U16181 (N_16181,N_12037,N_6839);
or U16182 (N_16182,N_6680,N_9725);
nor U16183 (N_16183,N_9150,N_10872);
or U16184 (N_16184,N_12456,N_6417);
and U16185 (N_16185,N_8288,N_12272);
nand U16186 (N_16186,N_9954,N_9767);
nand U16187 (N_16187,N_8253,N_7000);
nor U16188 (N_16188,N_9625,N_7020);
nand U16189 (N_16189,N_10029,N_10290);
or U16190 (N_16190,N_9417,N_6609);
nor U16191 (N_16191,N_8244,N_6409);
or U16192 (N_16192,N_11743,N_10578);
or U16193 (N_16193,N_9553,N_11603);
or U16194 (N_16194,N_11571,N_8250);
and U16195 (N_16195,N_7967,N_12154);
or U16196 (N_16196,N_9619,N_7842);
or U16197 (N_16197,N_8962,N_9024);
or U16198 (N_16198,N_7713,N_11271);
nand U16199 (N_16199,N_6424,N_9268);
and U16200 (N_16200,N_6639,N_8380);
nor U16201 (N_16201,N_7081,N_12428);
nor U16202 (N_16202,N_7107,N_6884);
and U16203 (N_16203,N_6293,N_11382);
nand U16204 (N_16204,N_6286,N_11138);
nor U16205 (N_16205,N_8402,N_9267);
nor U16206 (N_16206,N_8887,N_10553);
and U16207 (N_16207,N_7289,N_10814);
nor U16208 (N_16208,N_9217,N_8900);
and U16209 (N_16209,N_6520,N_6289);
nor U16210 (N_16210,N_9610,N_6357);
nor U16211 (N_16211,N_6799,N_11346);
nand U16212 (N_16212,N_10931,N_6827);
nand U16213 (N_16213,N_9098,N_9320);
and U16214 (N_16214,N_11512,N_11014);
nand U16215 (N_16215,N_11035,N_11896);
nand U16216 (N_16216,N_11000,N_11656);
nor U16217 (N_16217,N_12131,N_6515);
or U16218 (N_16218,N_6276,N_9149);
nand U16219 (N_16219,N_7685,N_9646);
nor U16220 (N_16220,N_9156,N_9921);
and U16221 (N_16221,N_11651,N_9186);
or U16222 (N_16222,N_6629,N_10643);
nand U16223 (N_16223,N_10453,N_6883);
nor U16224 (N_16224,N_7541,N_11866);
or U16225 (N_16225,N_9058,N_12131);
nand U16226 (N_16226,N_6692,N_11429);
nand U16227 (N_16227,N_6529,N_8530);
and U16228 (N_16228,N_7532,N_11392);
nand U16229 (N_16229,N_10073,N_10311);
and U16230 (N_16230,N_6544,N_9874);
nor U16231 (N_16231,N_7785,N_10113);
and U16232 (N_16232,N_7059,N_12381);
nor U16233 (N_16233,N_9636,N_7412);
and U16234 (N_16234,N_6404,N_7097);
nand U16235 (N_16235,N_7785,N_6760);
or U16236 (N_16236,N_7804,N_9706);
nor U16237 (N_16237,N_6885,N_7468);
nor U16238 (N_16238,N_9679,N_12291);
xnor U16239 (N_16239,N_9425,N_10922);
nand U16240 (N_16240,N_12338,N_11788);
nor U16241 (N_16241,N_7537,N_10679);
or U16242 (N_16242,N_11838,N_12176);
and U16243 (N_16243,N_12006,N_10800);
nor U16244 (N_16244,N_7104,N_9945);
and U16245 (N_16245,N_12255,N_8723);
xor U16246 (N_16246,N_6769,N_8236);
and U16247 (N_16247,N_11573,N_7430);
and U16248 (N_16248,N_11084,N_10677);
nand U16249 (N_16249,N_8204,N_7057);
nand U16250 (N_16250,N_11378,N_10541);
and U16251 (N_16251,N_12196,N_10126);
nand U16252 (N_16252,N_11071,N_7261);
and U16253 (N_16253,N_10934,N_6510);
or U16254 (N_16254,N_8599,N_8037);
nor U16255 (N_16255,N_8363,N_6302);
and U16256 (N_16256,N_12099,N_7600);
nand U16257 (N_16257,N_6387,N_10149);
nor U16258 (N_16258,N_6998,N_6636);
and U16259 (N_16259,N_7339,N_6281);
or U16260 (N_16260,N_6621,N_12464);
and U16261 (N_16261,N_8773,N_11213);
nor U16262 (N_16262,N_10824,N_6967);
and U16263 (N_16263,N_10207,N_7183);
nor U16264 (N_16264,N_8242,N_6997);
nor U16265 (N_16265,N_7948,N_7775);
and U16266 (N_16266,N_7771,N_9752);
xor U16267 (N_16267,N_11559,N_7730);
nor U16268 (N_16268,N_9083,N_9593);
nand U16269 (N_16269,N_7105,N_8336);
or U16270 (N_16270,N_7050,N_12357);
and U16271 (N_16271,N_6962,N_7746);
nor U16272 (N_16272,N_12400,N_8263);
nand U16273 (N_16273,N_10416,N_11619);
or U16274 (N_16274,N_6768,N_12155);
and U16275 (N_16275,N_6903,N_8008);
nand U16276 (N_16276,N_11210,N_7793);
xnor U16277 (N_16277,N_9264,N_11217);
nor U16278 (N_16278,N_9855,N_10484);
nor U16279 (N_16279,N_11816,N_8006);
and U16280 (N_16280,N_7175,N_8868);
or U16281 (N_16281,N_10860,N_7672);
and U16282 (N_16282,N_6887,N_6895);
and U16283 (N_16283,N_8273,N_7062);
or U16284 (N_16284,N_11056,N_9223);
nor U16285 (N_16285,N_11882,N_11137);
or U16286 (N_16286,N_12372,N_11464);
and U16287 (N_16287,N_12376,N_6542);
and U16288 (N_16288,N_6874,N_6663);
nor U16289 (N_16289,N_8738,N_9423);
and U16290 (N_16290,N_10310,N_8130);
or U16291 (N_16291,N_6763,N_12098);
nor U16292 (N_16292,N_12399,N_6798);
nor U16293 (N_16293,N_7496,N_10973);
or U16294 (N_16294,N_11761,N_6371);
nor U16295 (N_16295,N_6861,N_7372);
nor U16296 (N_16296,N_10687,N_10440);
and U16297 (N_16297,N_9024,N_10188);
and U16298 (N_16298,N_9869,N_10140);
nor U16299 (N_16299,N_6914,N_10044);
or U16300 (N_16300,N_8112,N_10232);
or U16301 (N_16301,N_8932,N_12289);
and U16302 (N_16302,N_12329,N_11464);
or U16303 (N_16303,N_8544,N_10486);
nor U16304 (N_16304,N_11703,N_8351);
or U16305 (N_16305,N_9610,N_9629);
or U16306 (N_16306,N_8936,N_12056);
nor U16307 (N_16307,N_9470,N_8873);
and U16308 (N_16308,N_9661,N_9412);
nand U16309 (N_16309,N_8008,N_6724);
nor U16310 (N_16310,N_6632,N_9373);
and U16311 (N_16311,N_8488,N_6752);
nor U16312 (N_16312,N_11319,N_10343);
nor U16313 (N_16313,N_10161,N_11146);
nor U16314 (N_16314,N_6787,N_8413);
or U16315 (N_16315,N_12150,N_7073);
and U16316 (N_16316,N_8629,N_9833);
and U16317 (N_16317,N_7871,N_6875);
nand U16318 (N_16318,N_8894,N_12452);
nand U16319 (N_16319,N_9816,N_6569);
or U16320 (N_16320,N_10562,N_6480);
nor U16321 (N_16321,N_8683,N_9440);
nor U16322 (N_16322,N_9638,N_10929);
nor U16323 (N_16323,N_11294,N_10599);
nor U16324 (N_16324,N_11058,N_7287);
or U16325 (N_16325,N_9136,N_10749);
nor U16326 (N_16326,N_11447,N_8003);
nand U16327 (N_16327,N_10074,N_7918);
and U16328 (N_16328,N_6692,N_10931);
nand U16329 (N_16329,N_7587,N_8368);
nand U16330 (N_16330,N_11277,N_7918);
nor U16331 (N_16331,N_10000,N_9369);
and U16332 (N_16332,N_10265,N_8909);
nor U16333 (N_16333,N_6824,N_10614);
and U16334 (N_16334,N_10765,N_7981);
and U16335 (N_16335,N_11786,N_8384);
nand U16336 (N_16336,N_6464,N_9388);
nand U16337 (N_16337,N_8364,N_7059);
nor U16338 (N_16338,N_11931,N_10523);
and U16339 (N_16339,N_9284,N_10687);
nand U16340 (N_16340,N_12041,N_6366);
or U16341 (N_16341,N_11310,N_9424);
nand U16342 (N_16342,N_8007,N_8644);
nor U16343 (N_16343,N_11661,N_8055);
or U16344 (N_16344,N_7306,N_7247);
and U16345 (N_16345,N_8208,N_6474);
and U16346 (N_16346,N_11614,N_10800);
nand U16347 (N_16347,N_10695,N_9276);
and U16348 (N_16348,N_9779,N_8237);
and U16349 (N_16349,N_11989,N_6356);
or U16350 (N_16350,N_8807,N_10747);
nand U16351 (N_16351,N_8675,N_10006);
nor U16352 (N_16352,N_12459,N_7284);
nand U16353 (N_16353,N_12160,N_6948);
and U16354 (N_16354,N_6717,N_10617);
nand U16355 (N_16355,N_12106,N_10249);
nor U16356 (N_16356,N_11622,N_8227);
nor U16357 (N_16357,N_9129,N_9824);
nand U16358 (N_16358,N_6265,N_11228);
or U16359 (N_16359,N_6487,N_8585);
or U16360 (N_16360,N_6652,N_10140);
nor U16361 (N_16361,N_10705,N_7449);
or U16362 (N_16362,N_12277,N_11660);
and U16363 (N_16363,N_10629,N_11381);
nor U16364 (N_16364,N_8658,N_9784);
nor U16365 (N_16365,N_10025,N_9896);
and U16366 (N_16366,N_10489,N_7963);
xnor U16367 (N_16367,N_7884,N_9936);
nor U16368 (N_16368,N_6275,N_12264);
nor U16369 (N_16369,N_7855,N_7765);
or U16370 (N_16370,N_10689,N_11132);
nand U16371 (N_16371,N_6812,N_9087);
nand U16372 (N_16372,N_6601,N_9186);
nor U16373 (N_16373,N_6448,N_12336);
xnor U16374 (N_16374,N_6561,N_6450);
nor U16375 (N_16375,N_10860,N_8327);
and U16376 (N_16376,N_9194,N_7387);
or U16377 (N_16377,N_9079,N_6655);
nand U16378 (N_16378,N_7249,N_9481);
nand U16379 (N_16379,N_8658,N_10022);
nand U16380 (N_16380,N_10231,N_11967);
nand U16381 (N_16381,N_6437,N_10326);
nor U16382 (N_16382,N_12111,N_11982);
and U16383 (N_16383,N_11879,N_12137);
nand U16384 (N_16384,N_12293,N_7379);
or U16385 (N_16385,N_10364,N_8571);
nand U16386 (N_16386,N_8536,N_10911);
and U16387 (N_16387,N_7398,N_12014);
or U16388 (N_16388,N_6281,N_7687);
and U16389 (N_16389,N_6407,N_7688);
or U16390 (N_16390,N_9385,N_6992);
and U16391 (N_16391,N_11448,N_10887);
nand U16392 (N_16392,N_9157,N_10331);
nor U16393 (N_16393,N_9433,N_7385);
nand U16394 (N_16394,N_9179,N_11282);
and U16395 (N_16395,N_12063,N_8829);
and U16396 (N_16396,N_6360,N_8566);
nand U16397 (N_16397,N_11563,N_10124);
nand U16398 (N_16398,N_6789,N_9194);
nand U16399 (N_16399,N_8996,N_10387);
nand U16400 (N_16400,N_6640,N_11993);
or U16401 (N_16401,N_10511,N_9705);
nor U16402 (N_16402,N_9282,N_11949);
nand U16403 (N_16403,N_7839,N_12041);
nand U16404 (N_16404,N_10930,N_8447);
or U16405 (N_16405,N_11549,N_8948);
nand U16406 (N_16406,N_10509,N_10123);
or U16407 (N_16407,N_11117,N_7820);
and U16408 (N_16408,N_8291,N_8605);
and U16409 (N_16409,N_9129,N_8192);
nand U16410 (N_16410,N_10530,N_8157);
nor U16411 (N_16411,N_7400,N_11582);
nand U16412 (N_16412,N_10290,N_10047);
nand U16413 (N_16413,N_11283,N_12076);
or U16414 (N_16414,N_10303,N_9473);
and U16415 (N_16415,N_12218,N_6867);
nor U16416 (N_16416,N_7261,N_8357);
or U16417 (N_16417,N_10596,N_12285);
nor U16418 (N_16418,N_11396,N_9760);
nand U16419 (N_16419,N_10359,N_10946);
and U16420 (N_16420,N_11992,N_7915);
nor U16421 (N_16421,N_11472,N_8050);
and U16422 (N_16422,N_11637,N_6404);
nor U16423 (N_16423,N_8438,N_7954);
nor U16424 (N_16424,N_12337,N_12329);
or U16425 (N_16425,N_11703,N_11443);
nand U16426 (N_16426,N_10993,N_10553);
nor U16427 (N_16427,N_11265,N_7930);
nand U16428 (N_16428,N_6639,N_6373);
and U16429 (N_16429,N_12300,N_7275);
and U16430 (N_16430,N_8069,N_10162);
and U16431 (N_16431,N_9591,N_7438);
nor U16432 (N_16432,N_11687,N_9469);
and U16433 (N_16433,N_12040,N_11887);
or U16434 (N_16434,N_10495,N_11445);
or U16435 (N_16435,N_10044,N_7181);
and U16436 (N_16436,N_6917,N_7829);
and U16437 (N_16437,N_8303,N_9225);
xor U16438 (N_16438,N_10275,N_8708);
nor U16439 (N_16439,N_11484,N_7290);
or U16440 (N_16440,N_11236,N_9437);
nor U16441 (N_16441,N_7489,N_8273);
or U16442 (N_16442,N_7925,N_8641);
nor U16443 (N_16443,N_10646,N_9478);
nand U16444 (N_16444,N_10674,N_7702);
nand U16445 (N_16445,N_10675,N_9587);
and U16446 (N_16446,N_11193,N_8996);
or U16447 (N_16447,N_11473,N_6680);
nor U16448 (N_16448,N_9316,N_7556);
and U16449 (N_16449,N_8701,N_11404);
and U16450 (N_16450,N_10728,N_7522);
and U16451 (N_16451,N_6511,N_10491);
and U16452 (N_16452,N_11630,N_10116);
or U16453 (N_16453,N_6526,N_10790);
xor U16454 (N_16454,N_11098,N_8616);
and U16455 (N_16455,N_7462,N_9332);
and U16456 (N_16456,N_8581,N_8144);
or U16457 (N_16457,N_9714,N_8677);
nand U16458 (N_16458,N_7986,N_9129);
nand U16459 (N_16459,N_8235,N_9227);
nand U16460 (N_16460,N_7995,N_10811);
nand U16461 (N_16461,N_10684,N_7907);
nand U16462 (N_16462,N_6275,N_9104);
or U16463 (N_16463,N_9654,N_9767);
nand U16464 (N_16464,N_9605,N_8620);
or U16465 (N_16465,N_9661,N_11122);
nor U16466 (N_16466,N_11907,N_11244);
nor U16467 (N_16467,N_11885,N_11763);
nor U16468 (N_16468,N_7284,N_11865);
nand U16469 (N_16469,N_8395,N_6577);
nor U16470 (N_16470,N_8433,N_8336);
xor U16471 (N_16471,N_12157,N_12499);
and U16472 (N_16472,N_8615,N_6421);
or U16473 (N_16473,N_12314,N_9277);
or U16474 (N_16474,N_10021,N_6790);
nor U16475 (N_16475,N_12147,N_11391);
nor U16476 (N_16476,N_9966,N_7173);
nor U16477 (N_16477,N_8624,N_11179);
nand U16478 (N_16478,N_6810,N_6624);
nor U16479 (N_16479,N_11086,N_8803);
and U16480 (N_16480,N_8809,N_11390);
nand U16481 (N_16481,N_6675,N_7387);
and U16482 (N_16482,N_11783,N_10139);
nor U16483 (N_16483,N_7191,N_9131);
nor U16484 (N_16484,N_8431,N_7800);
nand U16485 (N_16485,N_7590,N_10649);
or U16486 (N_16486,N_10864,N_10516);
nor U16487 (N_16487,N_9909,N_9376);
nor U16488 (N_16488,N_7124,N_8978);
nand U16489 (N_16489,N_11017,N_9267);
and U16490 (N_16490,N_8092,N_6286);
or U16491 (N_16491,N_11539,N_8026);
and U16492 (N_16492,N_10967,N_7610);
and U16493 (N_16493,N_6543,N_11289);
nor U16494 (N_16494,N_10517,N_6782);
and U16495 (N_16495,N_7547,N_7846);
nor U16496 (N_16496,N_10956,N_7023);
nor U16497 (N_16497,N_9720,N_6723);
nand U16498 (N_16498,N_10102,N_11603);
nand U16499 (N_16499,N_8087,N_9619);
and U16500 (N_16500,N_10348,N_11764);
or U16501 (N_16501,N_7106,N_12032);
nor U16502 (N_16502,N_7642,N_11936);
and U16503 (N_16503,N_10264,N_6950);
and U16504 (N_16504,N_8091,N_9234);
nor U16505 (N_16505,N_11532,N_7419);
xnor U16506 (N_16506,N_12125,N_9633);
nand U16507 (N_16507,N_10858,N_9520);
and U16508 (N_16508,N_7877,N_8398);
or U16509 (N_16509,N_8499,N_8672);
and U16510 (N_16510,N_9104,N_10991);
nand U16511 (N_16511,N_8620,N_12294);
or U16512 (N_16512,N_8046,N_9608);
or U16513 (N_16513,N_11692,N_12372);
nand U16514 (N_16514,N_12360,N_11172);
nand U16515 (N_16515,N_8948,N_11123);
and U16516 (N_16516,N_7945,N_6983);
or U16517 (N_16517,N_11264,N_9971);
or U16518 (N_16518,N_8496,N_10203);
nor U16519 (N_16519,N_8492,N_10667);
or U16520 (N_16520,N_10482,N_6737);
or U16521 (N_16521,N_9508,N_7003);
nand U16522 (N_16522,N_8865,N_10149);
or U16523 (N_16523,N_11617,N_11931);
and U16524 (N_16524,N_9412,N_8803);
nand U16525 (N_16525,N_10368,N_7351);
or U16526 (N_16526,N_8424,N_6489);
or U16527 (N_16527,N_6575,N_6312);
or U16528 (N_16528,N_8162,N_9249);
or U16529 (N_16529,N_7023,N_10212);
nand U16530 (N_16530,N_10827,N_11926);
or U16531 (N_16531,N_11933,N_11313);
nor U16532 (N_16532,N_9142,N_11280);
or U16533 (N_16533,N_12407,N_10084);
nor U16534 (N_16534,N_11100,N_9810);
and U16535 (N_16535,N_6725,N_12414);
nor U16536 (N_16536,N_6735,N_10443);
nor U16537 (N_16537,N_10156,N_11102);
and U16538 (N_16538,N_10225,N_11949);
nor U16539 (N_16539,N_7198,N_10640);
or U16540 (N_16540,N_8492,N_9613);
nor U16541 (N_16541,N_11693,N_9612);
and U16542 (N_16542,N_7832,N_6981);
nor U16543 (N_16543,N_11564,N_8866);
nor U16544 (N_16544,N_8929,N_6844);
or U16545 (N_16545,N_7825,N_6874);
or U16546 (N_16546,N_11508,N_8070);
and U16547 (N_16547,N_12331,N_7402);
and U16548 (N_16548,N_11999,N_10619);
nand U16549 (N_16549,N_9069,N_8456);
nand U16550 (N_16550,N_9938,N_10846);
and U16551 (N_16551,N_8810,N_9951);
or U16552 (N_16552,N_11032,N_8140);
nand U16553 (N_16553,N_12320,N_11645);
nor U16554 (N_16554,N_10176,N_7755);
and U16555 (N_16555,N_8811,N_10906);
and U16556 (N_16556,N_7925,N_10969);
nor U16557 (N_16557,N_11166,N_11133);
xor U16558 (N_16558,N_6731,N_6726);
or U16559 (N_16559,N_11208,N_10595);
nor U16560 (N_16560,N_10117,N_11333);
nor U16561 (N_16561,N_12483,N_8021);
and U16562 (N_16562,N_8112,N_10770);
nand U16563 (N_16563,N_8213,N_11222);
or U16564 (N_16564,N_11627,N_6340);
nor U16565 (N_16565,N_11712,N_11459);
xnor U16566 (N_16566,N_9738,N_8098);
or U16567 (N_16567,N_11669,N_11159);
and U16568 (N_16568,N_7845,N_6505);
or U16569 (N_16569,N_12434,N_8430);
nor U16570 (N_16570,N_8630,N_10248);
nand U16571 (N_16571,N_8520,N_9317);
nor U16572 (N_16572,N_11296,N_10553);
and U16573 (N_16573,N_7289,N_7031);
or U16574 (N_16574,N_10675,N_9669);
or U16575 (N_16575,N_12423,N_11962);
xor U16576 (N_16576,N_6403,N_7869);
nand U16577 (N_16577,N_11029,N_7189);
nor U16578 (N_16578,N_9632,N_11439);
nand U16579 (N_16579,N_6430,N_9876);
and U16580 (N_16580,N_8788,N_7024);
or U16581 (N_16581,N_8896,N_11089);
nand U16582 (N_16582,N_9880,N_11481);
or U16583 (N_16583,N_7037,N_6668);
nand U16584 (N_16584,N_11649,N_8913);
nand U16585 (N_16585,N_8658,N_7661);
or U16586 (N_16586,N_9173,N_7344);
nor U16587 (N_16587,N_8008,N_11048);
nand U16588 (N_16588,N_11129,N_9518);
or U16589 (N_16589,N_12142,N_8822);
nor U16590 (N_16590,N_9446,N_8151);
or U16591 (N_16591,N_11297,N_10084);
nor U16592 (N_16592,N_10816,N_10003);
nor U16593 (N_16593,N_7957,N_9876);
or U16594 (N_16594,N_7108,N_8991);
nor U16595 (N_16595,N_10986,N_9387);
nand U16596 (N_16596,N_9326,N_9409);
or U16597 (N_16597,N_12090,N_10319);
nor U16598 (N_16598,N_9843,N_8799);
nand U16599 (N_16599,N_6802,N_8718);
or U16600 (N_16600,N_11409,N_10089);
or U16601 (N_16601,N_7967,N_6963);
or U16602 (N_16602,N_6816,N_8222);
and U16603 (N_16603,N_9431,N_8595);
nor U16604 (N_16604,N_10334,N_7138);
or U16605 (N_16605,N_7257,N_8928);
nand U16606 (N_16606,N_6255,N_9677);
or U16607 (N_16607,N_8677,N_11711);
or U16608 (N_16608,N_12047,N_9408);
and U16609 (N_16609,N_7176,N_7002);
and U16610 (N_16610,N_8454,N_10551);
nand U16611 (N_16611,N_12188,N_8084);
or U16612 (N_16612,N_6938,N_10588);
and U16613 (N_16613,N_6812,N_12194);
nor U16614 (N_16614,N_8167,N_9118);
xnor U16615 (N_16615,N_11421,N_10220);
and U16616 (N_16616,N_11975,N_10421);
nand U16617 (N_16617,N_9519,N_7900);
nor U16618 (N_16618,N_9058,N_10720);
nand U16619 (N_16619,N_11854,N_10672);
and U16620 (N_16620,N_6297,N_7880);
nor U16621 (N_16621,N_8957,N_10051);
nand U16622 (N_16622,N_11804,N_9796);
nor U16623 (N_16623,N_9915,N_8926);
nor U16624 (N_16624,N_11626,N_9903);
nor U16625 (N_16625,N_12285,N_7428);
and U16626 (N_16626,N_8430,N_6820);
nor U16627 (N_16627,N_11740,N_11032);
and U16628 (N_16628,N_6756,N_7961);
nor U16629 (N_16629,N_8174,N_9182);
or U16630 (N_16630,N_8943,N_7702);
xor U16631 (N_16631,N_10908,N_12161);
nand U16632 (N_16632,N_10317,N_8459);
or U16633 (N_16633,N_11107,N_12063);
nand U16634 (N_16634,N_7677,N_10552);
nand U16635 (N_16635,N_11692,N_10431);
nand U16636 (N_16636,N_9303,N_10582);
and U16637 (N_16637,N_8033,N_9137);
or U16638 (N_16638,N_10925,N_6627);
and U16639 (N_16639,N_11172,N_7851);
nor U16640 (N_16640,N_7101,N_12460);
nor U16641 (N_16641,N_12296,N_9015);
nand U16642 (N_16642,N_9306,N_7464);
nor U16643 (N_16643,N_9764,N_9169);
and U16644 (N_16644,N_9328,N_11729);
or U16645 (N_16645,N_7498,N_8560);
and U16646 (N_16646,N_8039,N_6814);
and U16647 (N_16647,N_11577,N_12307);
nand U16648 (N_16648,N_9741,N_8511);
nand U16649 (N_16649,N_9299,N_8618);
nor U16650 (N_16650,N_6329,N_10228);
nor U16651 (N_16651,N_8272,N_12250);
or U16652 (N_16652,N_6927,N_6438);
nor U16653 (N_16653,N_9496,N_10157);
nor U16654 (N_16654,N_8624,N_6723);
nor U16655 (N_16655,N_7280,N_7199);
nor U16656 (N_16656,N_7601,N_6419);
and U16657 (N_16657,N_10119,N_11396);
and U16658 (N_16658,N_7398,N_7718);
or U16659 (N_16659,N_10480,N_8968);
nor U16660 (N_16660,N_7677,N_12017);
and U16661 (N_16661,N_9040,N_6426);
nand U16662 (N_16662,N_6284,N_8116);
nand U16663 (N_16663,N_9897,N_11475);
and U16664 (N_16664,N_10393,N_6771);
nor U16665 (N_16665,N_8490,N_11408);
and U16666 (N_16666,N_9162,N_9897);
nor U16667 (N_16667,N_6371,N_6740);
or U16668 (N_16668,N_10310,N_8550);
or U16669 (N_16669,N_6812,N_10671);
nor U16670 (N_16670,N_6564,N_7092);
nor U16671 (N_16671,N_10631,N_9175);
or U16672 (N_16672,N_8005,N_6473);
nand U16673 (N_16673,N_9371,N_8264);
nand U16674 (N_16674,N_10222,N_7440);
xor U16675 (N_16675,N_6602,N_12053);
and U16676 (N_16676,N_9235,N_7514);
xnor U16677 (N_16677,N_10564,N_11115);
and U16678 (N_16678,N_11166,N_7695);
nor U16679 (N_16679,N_8242,N_8090);
and U16680 (N_16680,N_8567,N_8821);
nor U16681 (N_16681,N_10416,N_9000);
or U16682 (N_16682,N_8384,N_7180);
and U16683 (N_16683,N_8844,N_9346);
nand U16684 (N_16684,N_9389,N_9119);
or U16685 (N_16685,N_10356,N_9003);
and U16686 (N_16686,N_6914,N_8479);
nand U16687 (N_16687,N_11278,N_10331);
nor U16688 (N_16688,N_6278,N_8437);
nand U16689 (N_16689,N_9316,N_6955);
or U16690 (N_16690,N_11101,N_6562);
or U16691 (N_16691,N_7860,N_10780);
or U16692 (N_16692,N_6371,N_10384);
and U16693 (N_16693,N_7688,N_11853);
nor U16694 (N_16694,N_9919,N_7873);
and U16695 (N_16695,N_7157,N_6714);
or U16696 (N_16696,N_7072,N_7739);
nor U16697 (N_16697,N_10897,N_10662);
and U16698 (N_16698,N_11501,N_12335);
nor U16699 (N_16699,N_7252,N_8672);
and U16700 (N_16700,N_6908,N_7785);
nand U16701 (N_16701,N_10704,N_6617);
and U16702 (N_16702,N_12163,N_12300);
nand U16703 (N_16703,N_10455,N_7948);
nand U16704 (N_16704,N_8809,N_12042);
nor U16705 (N_16705,N_7558,N_7954);
nand U16706 (N_16706,N_7047,N_6265);
nor U16707 (N_16707,N_11885,N_8855);
and U16708 (N_16708,N_7047,N_6579);
nand U16709 (N_16709,N_7661,N_11482);
nor U16710 (N_16710,N_7029,N_7464);
nor U16711 (N_16711,N_9590,N_10822);
or U16712 (N_16712,N_10793,N_11335);
xnor U16713 (N_16713,N_12063,N_7602);
and U16714 (N_16714,N_7462,N_6795);
nor U16715 (N_16715,N_10191,N_11765);
nand U16716 (N_16716,N_7581,N_11631);
nor U16717 (N_16717,N_11789,N_6406);
or U16718 (N_16718,N_10563,N_8939);
nand U16719 (N_16719,N_8775,N_9223);
nor U16720 (N_16720,N_8830,N_9386);
nand U16721 (N_16721,N_11669,N_7321);
nor U16722 (N_16722,N_10023,N_7280);
or U16723 (N_16723,N_10478,N_9374);
and U16724 (N_16724,N_7001,N_9959);
and U16725 (N_16725,N_6793,N_10362);
and U16726 (N_16726,N_11851,N_8798);
nand U16727 (N_16727,N_11637,N_6993);
and U16728 (N_16728,N_9690,N_12146);
and U16729 (N_16729,N_6335,N_10914);
or U16730 (N_16730,N_9721,N_9435);
nor U16731 (N_16731,N_7712,N_10907);
or U16732 (N_16732,N_11278,N_11380);
nand U16733 (N_16733,N_8590,N_12392);
xor U16734 (N_16734,N_9885,N_10407);
and U16735 (N_16735,N_6926,N_12311);
nand U16736 (N_16736,N_10301,N_6631);
nor U16737 (N_16737,N_8713,N_9561);
nand U16738 (N_16738,N_8230,N_7948);
nand U16739 (N_16739,N_9913,N_12302);
and U16740 (N_16740,N_11854,N_12363);
or U16741 (N_16741,N_11279,N_8748);
nand U16742 (N_16742,N_6784,N_8162);
nor U16743 (N_16743,N_6689,N_7218);
and U16744 (N_16744,N_11812,N_12367);
nand U16745 (N_16745,N_10328,N_8984);
nand U16746 (N_16746,N_9496,N_9901);
nor U16747 (N_16747,N_9160,N_8422);
and U16748 (N_16748,N_9232,N_11653);
nand U16749 (N_16749,N_9340,N_10687);
and U16750 (N_16750,N_8968,N_8779);
nand U16751 (N_16751,N_11907,N_7853);
nor U16752 (N_16752,N_8750,N_11085);
nor U16753 (N_16753,N_10092,N_9474);
nand U16754 (N_16754,N_8418,N_11907);
nor U16755 (N_16755,N_11744,N_10459);
or U16756 (N_16756,N_10116,N_12078);
xnor U16757 (N_16757,N_9187,N_10239);
or U16758 (N_16758,N_7132,N_7043);
xnor U16759 (N_16759,N_9286,N_9616);
or U16760 (N_16760,N_9931,N_9945);
and U16761 (N_16761,N_9297,N_11318);
or U16762 (N_16762,N_7553,N_8848);
nand U16763 (N_16763,N_10987,N_12166);
and U16764 (N_16764,N_11367,N_7309);
nand U16765 (N_16765,N_12390,N_7529);
and U16766 (N_16766,N_10488,N_9100);
nor U16767 (N_16767,N_11661,N_11534);
nand U16768 (N_16768,N_10860,N_7931);
and U16769 (N_16769,N_8426,N_6629);
and U16770 (N_16770,N_11407,N_11753);
nor U16771 (N_16771,N_7954,N_10573);
and U16772 (N_16772,N_9658,N_8189);
and U16773 (N_16773,N_8756,N_11326);
xnor U16774 (N_16774,N_11293,N_8380);
or U16775 (N_16775,N_12187,N_9252);
nand U16776 (N_16776,N_10846,N_11502);
nor U16777 (N_16777,N_7181,N_9144);
nand U16778 (N_16778,N_7094,N_11968);
and U16779 (N_16779,N_8951,N_6910);
and U16780 (N_16780,N_6934,N_7377);
nor U16781 (N_16781,N_8054,N_12147);
or U16782 (N_16782,N_10586,N_7836);
nor U16783 (N_16783,N_12462,N_10173);
or U16784 (N_16784,N_8150,N_8637);
nand U16785 (N_16785,N_8557,N_9412);
nand U16786 (N_16786,N_7257,N_8549);
and U16787 (N_16787,N_7175,N_6386);
or U16788 (N_16788,N_11779,N_9571);
nand U16789 (N_16789,N_8722,N_10386);
and U16790 (N_16790,N_11526,N_10125);
or U16791 (N_16791,N_11595,N_7199);
nand U16792 (N_16792,N_6518,N_8855);
and U16793 (N_16793,N_9879,N_8803);
nor U16794 (N_16794,N_8758,N_7781);
nor U16795 (N_16795,N_10662,N_11955);
nor U16796 (N_16796,N_6324,N_11130);
nand U16797 (N_16797,N_9214,N_8729);
nor U16798 (N_16798,N_6407,N_12093);
or U16799 (N_16799,N_7009,N_10579);
or U16800 (N_16800,N_7302,N_9433);
and U16801 (N_16801,N_9756,N_6283);
nand U16802 (N_16802,N_8661,N_10968);
or U16803 (N_16803,N_8124,N_8250);
or U16804 (N_16804,N_6868,N_10616);
nor U16805 (N_16805,N_8065,N_7117);
nor U16806 (N_16806,N_7944,N_12334);
and U16807 (N_16807,N_11829,N_9207);
or U16808 (N_16808,N_11869,N_11390);
nand U16809 (N_16809,N_11127,N_7370);
or U16810 (N_16810,N_12378,N_6321);
nand U16811 (N_16811,N_10379,N_8320);
or U16812 (N_16812,N_12437,N_8308);
or U16813 (N_16813,N_6869,N_7207);
and U16814 (N_16814,N_9828,N_9646);
and U16815 (N_16815,N_11009,N_6933);
nor U16816 (N_16816,N_10122,N_11536);
and U16817 (N_16817,N_11898,N_11588);
nand U16818 (N_16818,N_8395,N_10734);
nand U16819 (N_16819,N_7838,N_12195);
and U16820 (N_16820,N_8843,N_8875);
and U16821 (N_16821,N_7463,N_10016);
and U16822 (N_16822,N_7485,N_10655);
or U16823 (N_16823,N_11690,N_6867);
nor U16824 (N_16824,N_12217,N_6278);
or U16825 (N_16825,N_7713,N_11113);
or U16826 (N_16826,N_8892,N_10481);
or U16827 (N_16827,N_7901,N_10934);
nor U16828 (N_16828,N_12160,N_11834);
and U16829 (N_16829,N_10162,N_8787);
nor U16830 (N_16830,N_6517,N_6561);
or U16831 (N_16831,N_11446,N_11391);
nand U16832 (N_16832,N_6306,N_7363);
nand U16833 (N_16833,N_9487,N_11158);
nand U16834 (N_16834,N_9069,N_8519);
nor U16835 (N_16835,N_11863,N_11871);
nand U16836 (N_16836,N_7651,N_12336);
nor U16837 (N_16837,N_7788,N_10708);
nand U16838 (N_16838,N_9956,N_12298);
and U16839 (N_16839,N_8412,N_10363);
nor U16840 (N_16840,N_10420,N_7469);
or U16841 (N_16841,N_9284,N_10633);
nor U16842 (N_16842,N_11694,N_9066);
nand U16843 (N_16843,N_9271,N_9805);
and U16844 (N_16844,N_7430,N_11138);
or U16845 (N_16845,N_10467,N_9190);
and U16846 (N_16846,N_8894,N_8946);
nor U16847 (N_16847,N_8015,N_9648);
nand U16848 (N_16848,N_10572,N_6991);
nand U16849 (N_16849,N_8829,N_10166);
or U16850 (N_16850,N_11863,N_11872);
nor U16851 (N_16851,N_7333,N_8099);
nor U16852 (N_16852,N_6355,N_10543);
nand U16853 (N_16853,N_7369,N_11595);
nor U16854 (N_16854,N_7777,N_7721);
nand U16855 (N_16855,N_8843,N_8546);
nand U16856 (N_16856,N_9606,N_8428);
nor U16857 (N_16857,N_10003,N_9908);
nand U16858 (N_16858,N_7492,N_10345);
nor U16859 (N_16859,N_6312,N_7529);
nor U16860 (N_16860,N_8931,N_7342);
or U16861 (N_16861,N_12241,N_7116);
or U16862 (N_16862,N_9002,N_10003);
or U16863 (N_16863,N_8802,N_10688);
or U16864 (N_16864,N_8778,N_11693);
or U16865 (N_16865,N_11390,N_10256);
nand U16866 (N_16866,N_6705,N_10954);
nor U16867 (N_16867,N_9774,N_9349);
and U16868 (N_16868,N_7776,N_10011);
or U16869 (N_16869,N_6407,N_12266);
nand U16870 (N_16870,N_11246,N_11440);
nor U16871 (N_16871,N_8487,N_9006);
or U16872 (N_16872,N_9845,N_7368);
nor U16873 (N_16873,N_12455,N_8510);
or U16874 (N_16874,N_10911,N_7027);
or U16875 (N_16875,N_6465,N_8965);
and U16876 (N_16876,N_6974,N_6744);
or U16877 (N_16877,N_10404,N_8881);
or U16878 (N_16878,N_7577,N_9583);
or U16879 (N_16879,N_11009,N_7341);
nor U16880 (N_16880,N_11480,N_7156);
or U16881 (N_16881,N_11102,N_7270);
and U16882 (N_16882,N_11981,N_12227);
nand U16883 (N_16883,N_9831,N_8803);
or U16884 (N_16884,N_9422,N_7710);
nor U16885 (N_16885,N_9142,N_9961);
or U16886 (N_16886,N_8137,N_7967);
nor U16887 (N_16887,N_10688,N_11286);
or U16888 (N_16888,N_12408,N_12058);
nand U16889 (N_16889,N_10366,N_8115);
nand U16890 (N_16890,N_11183,N_11335);
nand U16891 (N_16891,N_8436,N_11618);
nor U16892 (N_16892,N_7859,N_11300);
nand U16893 (N_16893,N_6965,N_7337);
nand U16894 (N_16894,N_10083,N_6278);
or U16895 (N_16895,N_12311,N_8731);
and U16896 (N_16896,N_12158,N_7915);
nand U16897 (N_16897,N_10578,N_8140);
nor U16898 (N_16898,N_12012,N_10630);
nand U16899 (N_16899,N_7898,N_7388);
nand U16900 (N_16900,N_9659,N_9053);
nand U16901 (N_16901,N_8129,N_9394);
nor U16902 (N_16902,N_9386,N_7635);
nand U16903 (N_16903,N_11912,N_12172);
nor U16904 (N_16904,N_11972,N_11691);
nand U16905 (N_16905,N_9661,N_10110);
nor U16906 (N_16906,N_12230,N_7680);
nor U16907 (N_16907,N_11302,N_7157);
nor U16908 (N_16908,N_10261,N_6976);
and U16909 (N_16909,N_10147,N_8282);
or U16910 (N_16910,N_10629,N_9268);
nand U16911 (N_16911,N_11637,N_7848);
or U16912 (N_16912,N_10769,N_8328);
xor U16913 (N_16913,N_9274,N_10064);
or U16914 (N_16914,N_7218,N_6721);
or U16915 (N_16915,N_7281,N_7029);
nor U16916 (N_16916,N_7255,N_11081);
nand U16917 (N_16917,N_10181,N_10148);
and U16918 (N_16918,N_7666,N_9354);
or U16919 (N_16919,N_8932,N_7997);
nor U16920 (N_16920,N_11321,N_9170);
nor U16921 (N_16921,N_11433,N_12449);
and U16922 (N_16922,N_7688,N_7603);
and U16923 (N_16923,N_10992,N_12212);
nor U16924 (N_16924,N_6570,N_8097);
or U16925 (N_16925,N_8524,N_6901);
nor U16926 (N_16926,N_6870,N_6405);
and U16927 (N_16927,N_9225,N_8801);
or U16928 (N_16928,N_12495,N_12372);
and U16929 (N_16929,N_10929,N_8642);
nor U16930 (N_16930,N_6868,N_8720);
and U16931 (N_16931,N_6433,N_9011);
and U16932 (N_16932,N_8310,N_6586);
and U16933 (N_16933,N_11528,N_8191);
nand U16934 (N_16934,N_6448,N_12012);
nor U16935 (N_16935,N_8953,N_9229);
or U16936 (N_16936,N_11727,N_6743);
or U16937 (N_16937,N_10104,N_8430);
or U16938 (N_16938,N_6278,N_8394);
nor U16939 (N_16939,N_9348,N_7187);
nand U16940 (N_16940,N_8724,N_8622);
nand U16941 (N_16941,N_10127,N_9572);
or U16942 (N_16942,N_6354,N_11524);
or U16943 (N_16943,N_10022,N_7946);
nor U16944 (N_16944,N_11562,N_9708);
nor U16945 (N_16945,N_8535,N_7560);
or U16946 (N_16946,N_9118,N_10104);
nor U16947 (N_16947,N_9768,N_11349);
and U16948 (N_16948,N_10767,N_7836);
or U16949 (N_16949,N_6984,N_10439);
or U16950 (N_16950,N_9154,N_10732);
or U16951 (N_16951,N_11113,N_6637);
nor U16952 (N_16952,N_8747,N_7769);
nand U16953 (N_16953,N_8895,N_12018);
nand U16954 (N_16954,N_11472,N_10573);
and U16955 (N_16955,N_10898,N_9362);
nand U16956 (N_16956,N_7211,N_8096);
nand U16957 (N_16957,N_10273,N_6758);
or U16958 (N_16958,N_10152,N_6913);
nand U16959 (N_16959,N_6411,N_10530);
or U16960 (N_16960,N_9673,N_11126);
nand U16961 (N_16961,N_9596,N_10700);
and U16962 (N_16962,N_7561,N_10185);
and U16963 (N_16963,N_9274,N_8555);
and U16964 (N_16964,N_9223,N_8197);
nor U16965 (N_16965,N_11971,N_11106);
nor U16966 (N_16966,N_9188,N_7278);
and U16967 (N_16967,N_8599,N_8956);
and U16968 (N_16968,N_7182,N_10832);
and U16969 (N_16969,N_11419,N_11510);
nand U16970 (N_16970,N_6261,N_7604);
nand U16971 (N_16971,N_8236,N_6691);
and U16972 (N_16972,N_6583,N_10237);
nor U16973 (N_16973,N_9070,N_8471);
and U16974 (N_16974,N_9343,N_10620);
or U16975 (N_16975,N_10229,N_11966);
nand U16976 (N_16976,N_9831,N_7557);
nor U16977 (N_16977,N_9612,N_11448);
nand U16978 (N_16978,N_6262,N_9177);
or U16979 (N_16979,N_11479,N_10050);
and U16980 (N_16980,N_10657,N_6770);
nor U16981 (N_16981,N_8463,N_11933);
and U16982 (N_16982,N_6389,N_7015);
or U16983 (N_16983,N_9877,N_8945);
and U16984 (N_16984,N_10828,N_11811);
and U16985 (N_16985,N_6505,N_11237);
nor U16986 (N_16986,N_10408,N_8528);
nor U16987 (N_16987,N_7220,N_9869);
nor U16988 (N_16988,N_8866,N_8453);
and U16989 (N_16989,N_7868,N_7503);
or U16990 (N_16990,N_9078,N_9875);
or U16991 (N_16991,N_8397,N_7601);
and U16992 (N_16992,N_8253,N_8382);
xnor U16993 (N_16993,N_8896,N_8160);
or U16994 (N_16994,N_8094,N_9502);
nor U16995 (N_16995,N_6847,N_11015);
or U16996 (N_16996,N_12374,N_8579);
and U16997 (N_16997,N_8308,N_6646);
nand U16998 (N_16998,N_11241,N_9129);
or U16999 (N_16999,N_6402,N_7686);
nor U17000 (N_17000,N_9071,N_11728);
nor U17001 (N_17001,N_9448,N_9185);
and U17002 (N_17002,N_12175,N_7697);
xnor U17003 (N_17003,N_10659,N_7825);
nand U17004 (N_17004,N_8950,N_10261);
and U17005 (N_17005,N_11876,N_9966);
nand U17006 (N_17006,N_10485,N_11245);
nor U17007 (N_17007,N_6402,N_10632);
nor U17008 (N_17008,N_8881,N_7253);
nor U17009 (N_17009,N_10301,N_9906);
or U17010 (N_17010,N_12032,N_8177);
nor U17011 (N_17011,N_8867,N_6801);
nor U17012 (N_17012,N_7861,N_11049);
nand U17013 (N_17013,N_6870,N_8265);
nand U17014 (N_17014,N_7381,N_11316);
nor U17015 (N_17015,N_8295,N_7534);
nor U17016 (N_17016,N_6950,N_6572);
nand U17017 (N_17017,N_10304,N_6953);
and U17018 (N_17018,N_7937,N_9257);
or U17019 (N_17019,N_8574,N_9469);
nor U17020 (N_17020,N_10336,N_7765);
nand U17021 (N_17021,N_8324,N_6987);
and U17022 (N_17022,N_11316,N_7554);
nor U17023 (N_17023,N_10111,N_7553);
nor U17024 (N_17024,N_10116,N_6409);
or U17025 (N_17025,N_8135,N_9487);
and U17026 (N_17026,N_9860,N_8386);
nor U17027 (N_17027,N_11576,N_6349);
or U17028 (N_17028,N_8298,N_8744);
nor U17029 (N_17029,N_9166,N_8771);
or U17030 (N_17030,N_9614,N_8818);
nor U17031 (N_17031,N_9305,N_7008);
or U17032 (N_17032,N_10438,N_7910);
and U17033 (N_17033,N_7387,N_7728);
and U17034 (N_17034,N_7959,N_10778);
nor U17035 (N_17035,N_7213,N_11513);
nand U17036 (N_17036,N_7739,N_11938);
and U17037 (N_17037,N_11302,N_9593);
or U17038 (N_17038,N_8625,N_8548);
and U17039 (N_17039,N_8546,N_11117);
and U17040 (N_17040,N_12036,N_11344);
nor U17041 (N_17041,N_11611,N_7476);
nand U17042 (N_17042,N_8573,N_11520);
and U17043 (N_17043,N_8522,N_8141);
and U17044 (N_17044,N_8984,N_6457);
and U17045 (N_17045,N_7090,N_8230);
or U17046 (N_17046,N_7704,N_6820);
nor U17047 (N_17047,N_6756,N_9988);
nand U17048 (N_17048,N_6577,N_11839);
and U17049 (N_17049,N_11755,N_11016);
nor U17050 (N_17050,N_8471,N_6805);
and U17051 (N_17051,N_10181,N_12375);
or U17052 (N_17052,N_8594,N_12369);
nand U17053 (N_17053,N_11907,N_6795);
nor U17054 (N_17054,N_6281,N_8674);
or U17055 (N_17055,N_10871,N_7501);
nand U17056 (N_17056,N_6418,N_6357);
nor U17057 (N_17057,N_9605,N_11041);
or U17058 (N_17058,N_6770,N_10853);
and U17059 (N_17059,N_8341,N_8646);
nor U17060 (N_17060,N_8194,N_7254);
nor U17061 (N_17061,N_7319,N_7608);
or U17062 (N_17062,N_10904,N_10711);
nor U17063 (N_17063,N_11329,N_7379);
and U17064 (N_17064,N_9631,N_7125);
and U17065 (N_17065,N_7549,N_6350);
nand U17066 (N_17066,N_10794,N_6343);
or U17067 (N_17067,N_9857,N_9174);
nand U17068 (N_17068,N_8298,N_7356);
and U17069 (N_17069,N_8021,N_11364);
and U17070 (N_17070,N_9377,N_11542);
or U17071 (N_17071,N_9893,N_10562);
or U17072 (N_17072,N_11318,N_11511);
nor U17073 (N_17073,N_6345,N_10840);
and U17074 (N_17074,N_11821,N_12106);
nand U17075 (N_17075,N_9175,N_11219);
or U17076 (N_17076,N_10177,N_7805);
or U17077 (N_17077,N_8432,N_10739);
nand U17078 (N_17078,N_8325,N_10155);
and U17079 (N_17079,N_6972,N_10465);
or U17080 (N_17080,N_9976,N_9517);
and U17081 (N_17081,N_9261,N_6537);
or U17082 (N_17082,N_7558,N_10029);
and U17083 (N_17083,N_7535,N_11354);
nand U17084 (N_17084,N_6547,N_8998);
or U17085 (N_17085,N_7989,N_7128);
and U17086 (N_17086,N_9802,N_8004);
nor U17087 (N_17087,N_8205,N_7673);
and U17088 (N_17088,N_9543,N_8144);
and U17089 (N_17089,N_9849,N_12398);
nand U17090 (N_17090,N_11729,N_12467);
nand U17091 (N_17091,N_12334,N_11287);
nand U17092 (N_17092,N_6746,N_11593);
and U17093 (N_17093,N_11073,N_7075);
and U17094 (N_17094,N_8779,N_10669);
nor U17095 (N_17095,N_7298,N_9399);
nor U17096 (N_17096,N_10075,N_6506);
nor U17097 (N_17097,N_11945,N_6739);
nor U17098 (N_17098,N_7074,N_10416);
or U17099 (N_17099,N_11179,N_7371);
nand U17100 (N_17100,N_11002,N_7095);
and U17101 (N_17101,N_10328,N_10922);
and U17102 (N_17102,N_7632,N_6272);
nand U17103 (N_17103,N_10817,N_9438);
nand U17104 (N_17104,N_10310,N_11779);
and U17105 (N_17105,N_9443,N_6950);
or U17106 (N_17106,N_9837,N_11226);
nand U17107 (N_17107,N_7891,N_7162);
and U17108 (N_17108,N_11999,N_11249);
nor U17109 (N_17109,N_6612,N_10209);
and U17110 (N_17110,N_10617,N_8595);
nor U17111 (N_17111,N_8953,N_12494);
or U17112 (N_17112,N_10844,N_10073);
nor U17113 (N_17113,N_6738,N_9103);
and U17114 (N_17114,N_8994,N_10562);
or U17115 (N_17115,N_7493,N_9542);
and U17116 (N_17116,N_10715,N_9107);
nor U17117 (N_17117,N_9395,N_6371);
nor U17118 (N_17118,N_8111,N_11899);
nand U17119 (N_17119,N_8435,N_7315);
or U17120 (N_17120,N_11041,N_6602);
or U17121 (N_17121,N_9935,N_9958);
and U17122 (N_17122,N_7698,N_12477);
or U17123 (N_17123,N_7698,N_8555);
and U17124 (N_17124,N_7072,N_7374);
nand U17125 (N_17125,N_7986,N_11730);
nand U17126 (N_17126,N_12243,N_10351);
nor U17127 (N_17127,N_8434,N_11769);
or U17128 (N_17128,N_7152,N_9130);
and U17129 (N_17129,N_10936,N_8420);
nor U17130 (N_17130,N_7343,N_7761);
nand U17131 (N_17131,N_8857,N_6625);
or U17132 (N_17132,N_6875,N_10928);
nor U17133 (N_17133,N_6578,N_12409);
nand U17134 (N_17134,N_12489,N_8996);
and U17135 (N_17135,N_6480,N_8976);
nand U17136 (N_17136,N_6703,N_7292);
and U17137 (N_17137,N_12065,N_7683);
or U17138 (N_17138,N_8161,N_6514);
nand U17139 (N_17139,N_8719,N_8789);
or U17140 (N_17140,N_10926,N_10930);
nand U17141 (N_17141,N_11546,N_7074);
nor U17142 (N_17142,N_6732,N_9170);
nor U17143 (N_17143,N_10140,N_12123);
and U17144 (N_17144,N_12192,N_7815);
nand U17145 (N_17145,N_8005,N_10592);
nand U17146 (N_17146,N_9295,N_11837);
nor U17147 (N_17147,N_8188,N_7410);
or U17148 (N_17148,N_10376,N_8806);
and U17149 (N_17149,N_12016,N_12049);
nand U17150 (N_17150,N_10261,N_11138);
nor U17151 (N_17151,N_8106,N_10286);
or U17152 (N_17152,N_7341,N_7247);
nand U17153 (N_17153,N_10306,N_9732);
and U17154 (N_17154,N_9443,N_7969);
nor U17155 (N_17155,N_8124,N_6471);
nor U17156 (N_17156,N_10908,N_12036);
nand U17157 (N_17157,N_11402,N_9296);
or U17158 (N_17158,N_11136,N_10734);
nor U17159 (N_17159,N_6323,N_10189);
nor U17160 (N_17160,N_12115,N_7221);
nor U17161 (N_17161,N_6455,N_9958);
nor U17162 (N_17162,N_11353,N_7537);
nor U17163 (N_17163,N_9175,N_10764);
nor U17164 (N_17164,N_10394,N_7842);
nor U17165 (N_17165,N_12216,N_11110);
or U17166 (N_17166,N_10006,N_12292);
or U17167 (N_17167,N_9544,N_6614);
nor U17168 (N_17168,N_9819,N_8423);
or U17169 (N_17169,N_10797,N_9768);
or U17170 (N_17170,N_9420,N_7959);
and U17171 (N_17171,N_9369,N_6600);
or U17172 (N_17172,N_9264,N_9093);
or U17173 (N_17173,N_11816,N_11793);
nor U17174 (N_17174,N_7742,N_10136);
nor U17175 (N_17175,N_9060,N_7957);
nor U17176 (N_17176,N_10047,N_12213);
nor U17177 (N_17177,N_10114,N_7794);
nand U17178 (N_17178,N_9089,N_9040);
nor U17179 (N_17179,N_7938,N_10943);
nand U17180 (N_17180,N_10779,N_7290);
and U17181 (N_17181,N_9063,N_11273);
nor U17182 (N_17182,N_8010,N_12185);
nand U17183 (N_17183,N_7978,N_12166);
nor U17184 (N_17184,N_8274,N_7619);
nor U17185 (N_17185,N_6684,N_8818);
or U17186 (N_17186,N_10491,N_10651);
nor U17187 (N_17187,N_8168,N_7167);
or U17188 (N_17188,N_10896,N_8371);
or U17189 (N_17189,N_7196,N_8972);
and U17190 (N_17190,N_11281,N_10154);
or U17191 (N_17191,N_11818,N_11276);
nand U17192 (N_17192,N_8436,N_7824);
or U17193 (N_17193,N_11611,N_12486);
or U17194 (N_17194,N_11499,N_12474);
nor U17195 (N_17195,N_6690,N_8835);
nand U17196 (N_17196,N_9823,N_7638);
and U17197 (N_17197,N_11764,N_9702);
and U17198 (N_17198,N_7260,N_11314);
nor U17199 (N_17199,N_8530,N_6758);
or U17200 (N_17200,N_9391,N_6640);
nor U17201 (N_17201,N_7213,N_8452);
or U17202 (N_17202,N_6442,N_9159);
and U17203 (N_17203,N_7536,N_12139);
or U17204 (N_17204,N_10622,N_11186);
or U17205 (N_17205,N_9341,N_10989);
or U17206 (N_17206,N_9813,N_10298);
and U17207 (N_17207,N_9126,N_8064);
nor U17208 (N_17208,N_8682,N_8388);
nand U17209 (N_17209,N_7186,N_10356);
or U17210 (N_17210,N_8923,N_10123);
nand U17211 (N_17211,N_9414,N_9928);
or U17212 (N_17212,N_7462,N_7287);
nand U17213 (N_17213,N_8778,N_7748);
and U17214 (N_17214,N_8081,N_9175);
nand U17215 (N_17215,N_11517,N_11392);
nand U17216 (N_17216,N_8229,N_7932);
or U17217 (N_17217,N_12246,N_12469);
nor U17218 (N_17218,N_12127,N_10672);
nor U17219 (N_17219,N_10423,N_12344);
nor U17220 (N_17220,N_8449,N_7684);
nor U17221 (N_17221,N_8355,N_11639);
nand U17222 (N_17222,N_9777,N_6681);
or U17223 (N_17223,N_9750,N_7609);
and U17224 (N_17224,N_10298,N_6598);
nand U17225 (N_17225,N_9256,N_8958);
and U17226 (N_17226,N_7066,N_12467);
or U17227 (N_17227,N_9655,N_10180);
nor U17228 (N_17228,N_12322,N_10514);
and U17229 (N_17229,N_11907,N_7419);
and U17230 (N_17230,N_9902,N_6357);
nand U17231 (N_17231,N_10552,N_9518);
nand U17232 (N_17232,N_9495,N_7528);
nand U17233 (N_17233,N_12395,N_9551);
or U17234 (N_17234,N_9793,N_10514);
and U17235 (N_17235,N_9210,N_6699);
nand U17236 (N_17236,N_7459,N_6302);
and U17237 (N_17237,N_11745,N_9259);
nor U17238 (N_17238,N_7956,N_10827);
nor U17239 (N_17239,N_7953,N_12232);
nor U17240 (N_17240,N_9909,N_8405);
and U17241 (N_17241,N_10548,N_7313);
nand U17242 (N_17242,N_6306,N_6784);
or U17243 (N_17243,N_9322,N_7617);
and U17244 (N_17244,N_7296,N_9941);
and U17245 (N_17245,N_10897,N_8491);
nand U17246 (N_17246,N_9258,N_6676);
nor U17247 (N_17247,N_6493,N_6710);
nor U17248 (N_17248,N_11969,N_11598);
or U17249 (N_17249,N_7655,N_6488);
nand U17250 (N_17250,N_8479,N_8007);
nor U17251 (N_17251,N_9998,N_11186);
or U17252 (N_17252,N_12297,N_6621);
nand U17253 (N_17253,N_6353,N_7467);
or U17254 (N_17254,N_10445,N_7825);
and U17255 (N_17255,N_6357,N_7032);
nand U17256 (N_17256,N_8272,N_8428);
and U17257 (N_17257,N_11115,N_9517);
and U17258 (N_17258,N_10634,N_8409);
nor U17259 (N_17259,N_10830,N_11639);
or U17260 (N_17260,N_9967,N_9263);
nor U17261 (N_17261,N_7708,N_7629);
nor U17262 (N_17262,N_8850,N_7041);
and U17263 (N_17263,N_7364,N_11845);
or U17264 (N_17264,N_11322,N_10759);
or U17265 (N_17265,N_9316,N_7834);
and U17266 (N_17266,N_11282,N_7026);
xnor U17267 (N_17267,N_10313,N_11468);
nand U17268 (N_17268,N_11310,N_10799);
or U17269 (N_17269,N_9396,N_9993);
and U17270 (N_17270,N_8659,N_8465);
and U17271 (N_17271,N_7199,N_12454);
or U17272 (N_17272,N_7584,N_7593);
or U17273 (N_17273,N_8929,N_7017);
or U17274 (N_17274,N_10232,N_8092);
nand U17275 (N_17275,N_9400,N_8540);
and U17276 (N_17276,N_8780,N_8390);
nand U17277 (N_17277,N_9930,N_8592);
or U17278 (N_17278,N_12462,N_10854);
and U17279 (N_17279,N_7590,N_7906);
or U17280 (N_17280,N_9951,N_10392);
nand U17281 (N_17281,N_9602,N_8090);
or U17282 (N_17282,N_8870,N_10886);
nand U17283 (N_17283,N_8764,N_8817);
and U17284 (N_17284,N_8433,N_7194);
or U17285 (N_17285,N_11823,N_9195);
and U17286 (N_17286,N_8798,N_7816);
nand U17287 (N_17287,N_10954,N_7403);
or U17288 (N_17288,N_8530,N_10268);
and U17289 (N_17289,N_10780,N_7673);
or U17290 (N_17290,N_11948,N_9502);
nor U17291 (N_17291,N_7254,N_12178);
and U17292 (N_17292,N_12003,N_11543);
nand U17293 (N_17293,N_8914,N_12345);
nand U17294 (N_17294,N_11983,N_10698);
nand U17295 (N_17295,N_8178,N_7331);
and U17296 (N_17296,N_9559,N_10521);
or U17297 (N_17297,N_6791,N_10194);
or U17298 (N_17298,N_10426,N_8433);
nand U17299 (N_17299,N_6966,N_12479);
nand U17300 (N_17300,N_12295,N_12261);
nand U17301 (N_17301,N_7778,N_7071);
or U17302 (N_17302,N_6311,N_11613);
or U17303 (N_17303,N_8286,N_10540);
nor U17304 (N_17304,N_9127,N_9737);
nand U17305 (N_17305,N_11770,N_10144);
nand U17306 (N_17306,N_7662,N_10045);
or U17307 (N_17307,N_9997,N_9820);
nand U17308 (N_17308,N_10721,N_8067);
nor U17309 (N_17309,N_11761,N_6560);
and U17310 (N_17310,N_9504,N_10877);
nor U17311 (N_17311,N_9012,N_10002);
nand U17312 (N_17312,N_6834,N_7463);
or U17313 (N_17313,N_7396,N_9595);
or U17314 (N_17314,N_6268,N_9625);
or U17315 (N_17315,N_8024,N_12163);
and U17316 (N_17316,N_11467,N_9414);
nor U17317 (N_17317,N_12064,N_11074);
or U17318 (N_17318,N_9522,N_7419);
nand U17319 (N_17319,N_6606,N_10327);
or U17320 (N_17320,N_9587,N_8557);
nor U17321 (N_17321,N_9475,N_10173);
nor U17322 (N_17322,N_8224,N_8774);
and U17323 (N_17323,N_6996,N_9288);
nand U17324 (N_17324,N_8330,N_12427);
nand U17325 (N_17325,N_9581,N_11615);
nand U17326 (N_17326,N_10622,N_9823);
nor U17327 (N_17327,N_9161,N_8151);
and U17328 (N_17328,N_6989,N_7942);
nand U17329 (N_17329,N_10903,N_6597);
nand U17330 (N_17330,N_8960,N_9635);
and U17331 (N_17331,N_10087,N_10601);
nor U17332 (N_17332,N_12384,N_11534);
or U17333 (N_17333,N_12350,N_10369);
nand U17334 (N_17334,N_9085,N_9693);
nor U17335 (N_17335,N_10461,N_6370);
nand U17336 (N_17336,N_11150,N_9297);
and U17337 (N_17337,N_9493,N_8284);
and U17338 (N_17338,N_12209,N_7488);
nor U17339 (N_17339,N_10530,N_8737);
and U17340 (N_17340,N_10956,N_6673);
and U17341 (N_17341,N_11263,N_7696);
and U17342 (N_17342,N_10827,N_10466);
nor U17343 (N_17343,N_12388,N_9384);
nand U17344 (N_17344,N_8056,N_11881);
nand U17345 (N_17345,N_8262,N_11739);
and U17346 (N_17346,N_8274,N_11370);
nor U17347 (N_17347,N_11240,N_7672);
xnor U17348 (N_17348,N_6938,N_9063);
nor U17349 (N_17349,N_10844,N_7297);
nand U17350 (N_17350,N_6751,N_9360);
nand U17351 (N_17351,N_7152,N_8951);
and U17352 (N_17352,N_12393,N_8328);
xor U17353 (N_17353,N_9647,N_11328);
and U17354 (N_17354,N_6820,N_7690);
or U17355 (N_17355,N_10834,N_10183);
or U17356 (N_17356,N_7914,N_6776);
nor U17357 (N_17357,N_6318,N_8658);
nor U17358 (N_17358,N_9810,N_9082);
nor U17359 (N_17359,N_9990,N_9966);
or U17360 (N_17360,N_8097,N_8346);
nand U17361 (N_17361,N_10782,N_7412);
nor U17362 (N_17362,N_7492,N_11606);
or U17363 (N_17363,N_9362,N_10828);
nor U17364 (N_17364,N_11735,N_10884);
nor U17365 (N_17365,N_9007,N_7955);
and U17366 (N_17366,N_10135,N_6871);
and U17367 (N_17367,N_6847,N_7372);
or U17368 (N_17368,N_9025,N_10539);
nand U17369 (N_17369,N_10705,N_8678);
or U17370 (N_17370,N_10815,N_6742);
nand U17371 (N_17371,N_6973,N_9779);
and U17372 (N_17372,N_11274,N_8671);
nand U17373 (N_17373,N_12324,N_8249);
or U17374 (N_17374,N_11905,N_9058);
or U17375 (N_17375,N_6494,N_8160);
nor U17376 (N_17376,N_6886,N_8880);
or U17377 (N_17377,N_6669,N_12389);
or U17378 (N_17378,N_7908,N_12286);
nand U17379 (N_17379,N_9411,N_6905);
or U17380 (N_17380,N_10624,N_8150);
nand U17381 (N_17381,N_11181,N_9586);
and U17382 (N_17382,N_9161,N_6594);
and U17383 (N_17383,N_8793,N_6867);
nand U17384 (N_17384,N_10410,N_7766);
nor U17385 (N_17385,N_11271,N_9945);
nand U17386 (N_17386,N_11249,N_11910);
or U17387 (N_17387,N_10640,N_10277);
nor U17388 (N_17388,N_7093,N_11868);
and U17389 (N_17389,N_6714,N_11629);
nor U17390 (N_17390,N_6956,N_7939);
or U17391 (N_17391,N_12367,N_7293);
nor U17392 (N_17392,N_10730,N_8909);
or U17393 (N_17393,N_8327,N_6487);
or U17394 (N_17394,N_12476,N_11860);
or U17395 (N_17395,N_7638,N_11755);
nand U17396 (N_17396,N_8534,N_11440);
nor U17397 (N_17397,N_10264,N_10761);
or U17398 (N_17398,N_11226,N_9285);
nand U17399 (N_17399,N_6971,N_12062);
and U17400 (N_17400,N_11512,N_12236);
nor U17401 (N_17401,N_10546,N_9900);
nor U17402 (N_17402,N_10252,N_6441);
or U17403 (N_17403,N_11200,N_9616);
nor U17404 (N_17404,N_8039,N_10170);
or U17405 (N_17405,N_9441,N_7799);
nor U17406 (N_17406,N_7755,N_9402);
and U17407 (N_17407,N_7669,N_10000);
and U17408 (N_17408,N_12391,N_9694);
and U17409 (N_17409,N_9956,N_6808);
nand U17410 (N_17410,N_6982,N_10083);
nor U17411 (N_17411,N_8689,N_12462);
nor U17412 (N_17412,N_10054,N_6664);
nand U17413 (N_17413,N_11544,N_9786);
nor U17414 (N_17414,N_11262,N_11128);
and U17415 (N_17415,N_9982,N_11073);
nand U17416 (N_17416,N_7521,N_6599);
nand U17417 (N_17417,N_11847,N_9980);
nand U17418 (N_17418,N_8242,N_7190);
nand U17419 (N_17419,N_7151,N_11960);
nand U17420 (N_17420,N_9318,N_6327);
nand U17421 (N_17421,N_11059,N_7131);
and U17422 (N_17422,N_8466,N_6803);
and U17423 (N_17423,N_7633,N_9081);
and U17424 (N_17424,N_10250,N_9283);
nand U17425 (N_17425,N_11703,N_8235);
or U17426 (N_17426,N_9079,N_11076);
nor U17427 (N_17427,N_11891,N_8892);
and U17428 (N_17428,N_10037,N_6529);
and U17429 (N_17429,N_11818,N_12060);
and U17430 (N_17430,N_8643,N_11788);
nand U17431 (N_17431,N_8438,N_7099);
nor U17432 (N_17432,N_11612,N_8513);
nand U17433 (N_17433,N_10205,N_9289);
and U17434 (N_17434,N_7244,N_10419);
and U17435 (N_17435,N_8361,N_6631);
nor U17436 (N_17436,N_10538,N_11974);
xor U17437 (N_17437,N_8693,N_10152);
and U17438 (N_17438,N_11632,N_10039);
nand U17439 (N_17439,N_9533,N_10937);
and U17440 (N_17440,N_12394,N_12383);
nand U17441 (N_17441,N_6309,N_9249);
or U17442 (N_17442,N_12247,N_8551);
nand U17443 (N_17443,N_6459,N_9592);
and U17444 (N_17444,N_8547,N_9748);
nor U17445 (N_17445,N_7209,N_11986);
and U17446 (N_17446,N_12475,N_9905);
nor U17447 (N_17447,N_11658,N_9445);
and U17448 (N_17448,N_8538,N_6630);
nand U17449 (N_17449,N_8176,N_10030);
or U17450 (N_17450,N_9552,N_11623);
and U17451 (N_17451,N_11497,N_8359);
nor U17452 (N_17452,N_8299,N_9076);
nor U17453 (N_17453,N_7146,N_7734);
or U17454 (N_17454,N_7366,N_9128);
nor U17455 (N_17455,N_8799,N_11645);
or U17456 (N_17456,N_12340,N_8038);
or U17457 (N_17457,N_8158,N_9272);
and U17458 (N_17458,N_8993,N_9987);
nor U17459 (N_17459,N_9075,N_10182);
nor U17460 (N_17460,N_6314,N_11755);
nand U17461 (N_17461,N_9352,N_10386);
nor U17462 (N_17462,N_7739,N_10590);
xor U17463 (N_17463,N_9990,N_9114);
nor U17464 (N_17464,N_9885,N_8516);
nand U17465 (N_17465,N_6428,N_8035);
nand U17466 (N_17466,N_11007,N_7792);
or U17467 (N_17467,N_6397,N_11886);
or U17468 (N_17468,N_12112,N_11158);
nor U17469 (N_17469,N_11190,N_9952);
and U17470 (N_17470,N_10933,N_11868);
nand U17471 (N_17471,N_9499,N_6314);
or U17472 (N_17472,N_10813,N_11014);
nand U17473 (N_17473,N_11079,N_11178);
nand U17474 (N_17474,N_8141,N_6978);
and U17475 (N_17475,N_6554,N_8008);
nand U17476 (N_17476,N_6273,N_6608);
nand U17477 (N_17477,N_9754,N_7011);
and U17478 (N_17478,N_9919,N_7707);
or U17479 (N_17479,N_9792,N_9800);
nor U17480 (N_17480,N_8083,N_6577);
nand U17481 (N_17481,N_11694,N_9437);
and U17482 (N_17482,N_11415,N_9332);
and U17483 (N_17483,N_6525,N_9294);
and U17484 (N_17484,N_10067,N_9193);
or U17485 (N_17485,N_10696,N_10328);
nand U17486 (N_17486,N_8481,N_8929);
and U17487 (N_17487,N_12408,N_7681);
nand U17488 (N_17488,N_11988,N_7473);
nor U17489 (N_17489,N_6465,N_11705);
nand U17490 (N_17490,N_8471,N_6826);
nand U17491 (N_17491,N_11217,N_6876);
nand U17492 (N_17492,N_6845,N_10663);
nor U17493 (N_17493,N_8925,N_8797);
or U17494 (N_17494,N_8423,N_10239);
and U17495 (N_17495,N_6908,N_10986);
nor U17496 (N_17496,N_7485,N_9613);
nor U17497 (N_17497,N_7977,N_6274);
and U17498 (N_17498,N_8275,N_9597);
or U17499 (N_17499,N_8525,N_9697);
nand U17500 (N_17500,N_6924,N_12026);
and U17501 (N_17501,N_8670,N_10317);
nor U17502 (N_17502,N_10445,N_7949);
or U17503 (N_17503,N_6666,N_8412);
nor U17504 (N_17504,N_12283,N_10640);
nand U17505 (N_17505,N_7463,N_8080);
nor U17506 (N_17506,N_7811,N_10367);
nand U17507 (N_17507,N_8180,N_6598);
xor U17508 (N_17508,N_12316,N_8837);
nor U17509 (N_17509,N_6526,N_7060);
nand U17510 (N_17510,N_10253,N_7104);
and U17511 (N_17511,N_8251,N_8290);
nand U17512 (N_17512,N_8543,N_7607);
or U17513 (N_17513,N_8104,N_11223);
nor U17514 (N_17514,N_6973,N_6873);
nor U17515 (N_17515,N_10741,N_8355);
and U17516 (N_17516,N_9662,N_9758);
or U17517 (N_17517,N_7258,N_10570);
or U17518 (N_17518,N_6594,N_10094);
and U17519 (N_17519,N_7268,N_12438);
nand U17520 (N_17520,N_10559,N_11060);
or U17521 (N_17521,N_6692,N_9648);
and U17522 (N_17522,N_9916,N_9607);
nor U17523 (N_17523,N_12144,N_8996);
or U17524 (N_17524,N_12259,N_8284);
nand U17525 (N_17525,N_7093,N_6250);
and U17526 (N_17526,N_9255,N_9233);
and U17527 (N_17527,N_10794,N_11441);
and U17528 (N_17528,N_10129,N_7258);
or U17529 (N_17529,N_9162,N_12177);
or U17530 (N_17530,N_11791,N_11637);
or U17531 (N_17531,N_7427,N_11565);
or U17532 (N_17532,N_9272,N_11324);
or U17533 (N_17533,N_10877,N_6256);
and U17534 (N_17534,N_11937,N_7102);
and U17535 (N_17535,N_11223,N_6830);
nand U17536 (N_17536,N_7837,N_7298);
or U17537 (N_17537,N_6366,N_11045);
nand U17538 (N_17538,N_11394,N_7007);
nor U17539 (N_17539,N_12270,N_8539);
nor U17540 (N_17540,N_11380,N_7399);
or U17541 (N_17541,N_11837,N_10370);
nand U17542 (N_17542,N_9909,N_11380);
nor U17543 (N_17543,N_8948,N_9497);
and U17544 (N_17544,N_9327,N_7829);
nor U17545 (N_17545,N_10312,N_7300);
nand U17546 (N_17546,N_6794,N_11504);
nand U17547 (N_17547,N_6873,N_6507);
nand U17548 (N_17548,N_8932,N_8677);
or U17549 (N_17549,N_9471,N_12231);
nand U17550 (N_17550,N_7285,N_7564);
nand U17551 (N_17551,N_10853,N_6678);
nor U17552 (N_17552,N_6259,N_10615);
nand U17553 (N_17553,N_9800,N_10251);
xor U17554 (N_17554,N_9408,N_8292);
nand U17555 (N_17555,N_6467,N_8871);
nand U17556 (N_17556,N_6836,N_12300);
or U17557 (N_17557,N_10948,N_9877);
nand U17558 (N_17558,N_11910,N_7047);
nor U17559 (N_17559,N_10078,N_8246);
xnor U17560 (N_17560,N_8176,N_6684);
or U17561 (N_17561,N_10771,N_7643);
nand U17562 (N_17562,N_11691,N_10925);
and U17563 (N_17563,N_11199,N_7064);
and U17564 (N_17564,N_7919,N_8538);
and U17565 (N_17565,N_11710,N_11091);
nor U17566 (N_17566,N_12204,N_9178);
and U17567 (N_17567,N_10951,N_8325);
xor U17568 (N_17568,N_9300,N_11249);
and U17569 (N_17569,N_9655,N_10913);
nand U17570 (N_17570,N_10486,N_6643);
and U17571 (N_17571,N_7121,N_9726);
and U17572 (N_17572,N_10422,N_10256);
or U17573 (N_17573,N_6671,N_9779);
nand U17574 (N_17574,N_8591,N_9986);
and U17575 (N_17575,N_11786,N_8502);
or U17576 (N_17576,N_8063,N_8469);
or U17577 (N_17577,N_8244,N_6929);
nand U17578 (N_17578,N_12358,N_10657);
and U17579 (N_17579,N_8182,N_6841);
and U17580 (N_17580,N_12086,N_11347);
or U17581 (N_17581,N_9012,N_11688);
nor U17582 (N_17582,N_10577,N_11497);
and U17583 (N_17583,N_11185,N_7991);
nand U17584 (N_17584,N_10045,N_6416);
and U17585 (N_17585,N_10826,N_8500);
and U17586 (N_17586,N_7449,N_12102);
and U17587 (N_17587,N_10202,N_9789);
or U17588 (N_17588,N_11075,N_11232);
nor U17589 (N_17589,N_11855,N_11290);
nor U17590 (N_17590,N_7456,N_11631);
nand U17591 (N_17591,N_7035,N_8739);
nand U17592 (N_17592,N_8814,N_8272);
or U17593 (N_17593,N_7648,N_9377);
or U17594 (N_17594,N_6321,N_7839);
and U17595 (N_17595,N_10846,N_12468);
nand U17596 (N_17596,N_12201,N_7852);
or U17597 (N_17597,N_12467,N_9808);
nor U17598 (N_17598,N_6989,N_6893);
nand U17599 (N_17599,N_6380,N_12488);
nand U17600 (N_17600,N_8146,N_8384);
nand U17601 (N_17601,N_9838,N_8225);
nor U17602 (N_17602,N_12351,N_10216);
or U17603 (N_17603,N_12323,N_11919);
and U17604 (N_17604,N_10889,N_10785);
nor U17605 (N_17605,N_7913,N_10913);
nand U17606 (N_17606,N_10314,N_12057);
or U17607 (N_17607,N_10783,N_11720);
and U17608 (N_17608,N_11457,N_7323);
nor U17609 (N_17609,N_8358,N_7505);
nand U17610 (N_17610,N_9124,N_11850);
nor U17611 (N_17611,N_10447,N_10575);
and U17612 (N_17612,N_12221,N_9622);
and U17613 (N_17613,N_8047,N_8835);
and U17614 (N_17614,N_9239,N_6796);
nor U17615 (N_17615,N_10700,N_10741);
or U17616 (N_17616,N_7382,N_6452);
and U17617 (N_17617,N_10682,N_10547);
or U17618 (N_17618,N_10192,N_11619);
or U17619 (N_17619,N_11408,N_8300);
and U17620 (N_17620,N_10277,N_7551);
and U17621 (N_17621,N_12060,N_10784);
nand U17622 (N_17622,N_7522,N_7616);
and U17623 (N_17623,N_10145,N_9404);
nor U17624 (N_17624,N_11791,N_11845);
and U17625 (N_17625,N_8984,N_9843);
or U17626 (N_17626,N_6831,N_7344);
nand U17627 (N_17627,N_10659,N_6430);
nor U17628 (N_17628,N_7603,N_6450);
or U17629 (N_17629,N_10889,N_11713);
and U17630 (N_17630,N_11861,N_12363);
nand U17631 (N_17631,N_9076,N_9936);
or U17632 (N_17632,N_11218,N_10571);
and U17633 (N_17633,N_11576,N_12316);
nor U17634 (N_17634,N_9675,N_11394);
nand U17635 (N_17635,N_11240,N_9524);
nand U17636 (N_17636,N_10878,N_8072);
nand U17637 (N_17637,N_7083,N_12012);
and U17638 (N_17638,N_12100,N_8889);
or U17639 (N_17639,N_6978,N_7538);
and U17640 (N_17640,N_11598,N_8888);
or U17641 (N_17641,N_10746,N_10896);
and U17642 (N_17642,N_9997,N_7528);
and U17643 (N_17643,N_8419,N_7554);
nand U17644 (N_17644,N_7924,N_9007);
nor U17645 (N_17645,N_7266,N_11112);
and U17646 (N_17646,N_10566,N_10909);
nand U17647 (N_17647,N_7740,N_6830);
and U17648 (N_17648,N_12132,N_10670);
or U17649 (N_17649,N_8241,N_12000);
or U17650 (N_17650,N_8942,N_10843);
nand U17651 (N_17651,N_10624,N_11973);
or U17652 (N_17652,N_7969,N_6654);
or U17653 (N_17653,N_6947,N_8518);
and U17654 (N_17654,N_6304,N_9112);
or U17655 (N_17655,N_9416,N_7637);
or U17656 (N_17656,N_8836,N_12252);
and U17657 (N_17657,N_7309,N_10984);
nor U17658 (N_17658,N_11014,N_12223);
and U17659 (N_17659,N_6699,N_12208);
nor U17660 (N_17660,N_9015,N_11020);
nor U17661 (N_17661,N_7769,N_10907);
or U17662 (N_17662,N_9957,N_12216);
and U17663 (N_17663,N_9028,N_7203);
nand U17664 (N_17664,N_9690,N_9976);
or U17665 (N_17665,N_8840,N_7777);
nand U17666 (N_17666,N_9280,N_7993);
and U17667 (N_17667,N_9723,N_11747);
and U17668 (N_17668,N_8793,N_11034);
nand U17669 (N_17669,N_10094,N_12196);
and U17670 (N_17670,N_12251,N_7663);
nor U17671 (N_17671,N_12412,N_10960);
nand U17672 (N_17672,N_9039,N_8869);
nand U17673 (N_17673,N_6546,N_8959);
and U17674 (N_17674,N_12219,N_9192);
nor U17675 (N_17675,N_8746,N_10498);
or U17676 (N_17676,N_12034,N_8573);
and U17677 (N_17677,N_9201,N_8431);
and U17678 (N_17678,N_8622,N_6798);
and U17679 (N_17679,N_6587,N_11849);
or U17680 (N_17680,N_11719,N_10922);
or U17681 (N_17681,N_6992,N_11640);
nor U17682 (N_17682,N_10963,N_10713);
nor U17683 (N_17683,N_11987,N_7233);
and U17684 (N_17684,N_12169,N_10369);
or U17685 (N_17685,N_11120,N_6281);
and U17686 (N_17686,N_11005,N_8772);
and U17687 (N_17687,N_10467,N_6353);
or U17688 (N_17688,N_9670,N_8937);
nor U17689 (N_17689,N_10644,N_9446);
and U17690 (N_17690,N_12008,N_10333);
and U17691 (N_17691,N_11962,N_8745);
and U17692 (N_17692,N_8485,N_9922);
and U17693 (N_17693,N_9558,N_8219);
nor U17694 (N_17694,N_9924,N_12320);
or U17695 (N_17695,N_11369,N_8825);
or U17696 (N_17696,N_10481,N_7110);
and U17697 (N_17697,N_10604,N_8230);
or U17698 (N_17698,N_6854,N_10745);
nand U17699 (N_17699,N_6895,N_10351);
nand U17700 (N_17700,N_11234,N_11227);
or U17701 (N_17701,N_10394,N_8618);
nor U17702 (N_17702,N_10569,N_11405);
and U17703 (N_17703,N_8951,N_11145);
nand U17704 (N_17704,N_8345,N_9451);
nor U17705 (N_17705,N_9723,N_10461);
xor U17706 (N_17706,N_10563,N_7544);
and U17707 (N_17707,N_10426,N_7762);
nor U17708 (N_17708,N_9638,N_11248);
nor U17709 (N_17709,N_6312,N_7138);
nand U17710 (N_17710,N_12215,N_7997);
or U17711 (N_17711,N_11083,N_8620);
nand U17712 (N_17712,N_10671,N_11115);
nand U17713 (N_17713,N_11607,N_7633);
or U17714 (N_17714,N_9739,N_11188);
nand U17715 (N_17715,N_7278,N_6334);
nor U17716 (N_17716,N_10944,N_10154);
nor U17717 (N_17717,N_6547,N_9331);
and U17718 (N_17718,N_8887,N_6934);
nor U17719 (N_17719,N_12334,N_10260);
and U17720 (N_17720,N_11626,N_12106);
or U17721 (N_17721,N_9747,N_10631);
nor U17722 (N_17722,N_10528,N_8977);
nor U17723 (N_17723,N_8323,N_7767);
xor U17724 (N_17724,N_10365,N_10320);
and U17725 (N_17725,N_8625,N_8072);
nand U17726 (N_17726,N_6386,N_7225);
nor U17727 (N_17727,N_8880,N_8306);
nand U17728 (N_17728,N_10193,N_7675);
nand U17729 (N_17729,N_10829,N_6535);
or U17730 (N_17730,N_7405,N_11717);
and U17731 (N_17731,N_6756,N_11550);
nand U17732 (N_17732,N_9661,N_9306);
nand U17733 (N_17733,N_10730,N_9726);
nand U17734 (N_17734,N_8529,N_7566);
xnor U17735 (N_17735,N_8139,N_8021);
nand U17736 (N_17736,N_7640,N_9017);
nor U17737 (N_17737,N_11080,N_9946);
or U17738 (N_17738,N_6671,N_9579);
nor U17739 (N_17739,N_11981,N_12082);
nor U17740 (N_17740,N_11868,N_7148);
nand U17741 (N_17741,N_6715,N_8855);
nor U17742 (N_17742,N_8217,N_12141);
and U17743 (N_17743,N_8126,N_10686);
nor U17744 (N_17744,N_8844,N_9153);
nor U17745 (N_17745,N_11360,N_10743);
or U17746 (N_17746,N_7007,N_9668);
nor U17747 (N_17747,N_8910,N_9427);
or U17748 (N_17748,N_9177,N_11290);
nand U17749 (N_17749,N_11737,N_6530);
nor U17750 (N_17750,N_8813,N_8803);
xor U17751 (N_17751,N_10505,N_7843);
and U17752 (N_17752,N_6586,N_11184);
nand U17753 (N_17753,N_9967,N_8004);
or U17754 (N_17754,N_7168,N_9242);
or U17755 (N_17755,N_7314,N_6649);
and U17756 (N_17756,N_7330,N_9730);
nand U17757 (N_17757,N_6438,N_9409);
xor U17758 (N_17758,N_11972,N_12191);
or U17759 (N_17759,N_6529,N_7290);
or U17760 (N_17760,N_12217,N_7983);
nor U17761 (N_17761,N_10131,N_8389);
nand U17762 (N_17762,N_7699,N_9869);
nand U17763 (N_17763,N_11024,N_9413);
nand U17764 (N_17764,N_11977,N_11831);
and U17765 (N_17765,N_10264,N_9968);
and U17766 (N_17766,N_9362,N_8460);
and U17767 (N_17767,N_11354,N_9534);
and U17768 (N_17768,N_8476,N_12345);
nor U17769 (N_17769,N_11799,N_11334);
or U17770 (N_17770,N_8136,N_12214);
nor U17771 (N_17771,N_10216,N_9025);
or U17772 (N_17772,N_10056,N_11676);
nor U17773 (N_17773,N_8762,N_9637);
nand U17774 (N_17774,N_11915,N_9394);
and U17775 (N_17775,N_8516,N_6654);
or U17776 (N_17776,N_10067,N_8310);
nand U17777 (N_17777,N_12184,N_12257);
nand U17778 (N_17778,N_11926,N_12260);
or U17779 (N_17779,N_8802,N_7814);
or U17780 (N_17780,N_8062,N_10800);
nor U17781 (N_17781,N_10506,N_7067);
or U17782 (N_17782,N_9159,N_9352);
and U17783 (N_17783,N_11369,N_9776);
nor U17784 (N_17784,N_9326,N_11979);
nand U17785 (N_17785,N_11089,N_12112);
nand U17786 (N_17786,N_11179,N_10353);
and U17787 (N_17787,N_11743,N_10820);
and U17788 (N_17788,N_6810,N_11888);
nor U17789 (N_17789,N_8435,N_8328);
and U17790 (N_17790,N_12343,N_7445);
nor U17791 (N_17791,N_7871,N_8165);
nor U17792 (N_17792,N_7660,N_8404);
and U17793 (N_17793,N_9571,N_10496);
or U17794 (N_17794,N_8850,N_7839);
or U17795 (N_17795,N_9031,N_7061);
nand U17796 (N_17796,N_6630,N_10371);
or U17797 (N_17797,N_7821,N_12357);
nor U17798 (N_17798,N_9048,N_7145);
and U17799 (N_17799,N_8790,N_6570);
nor U17800 (N_17800,N_9305,N_10604);
or U17801 (N_17801,N_7451,N_9443);
and U17802 (N_17802,N_7172,N_6567);
or U17803 (N_17803,N_12494,N_10557);
nand U17804 (N_17804,N_6621,N_11129);
or U17805 (N_17805,N_6576,N_12410);
and U17806 (N_17806,N_9270,N_10861);
and U17807 (N_17807,N_9844,N_9486);
nand U17808 (N_17808,N_9434,N_12039);
and U17809 (N_17809,N_12158,N_9221);
nor U17810 (N_17810,N_11352,N_9419);
nand U17811 (N_17811,N_11127,N_8388);
nor U17812 (N_17812,N_8994,N_11743);
and U17813 (N_17813,N_11804,N_7268);
nor U17814 (N_17814,N_8212,N_9904);
and U17815 (N_17815,N_9181,N_8744);
nor U17816 (N_17816,N_11942,N_11556);
nand U17817 (N_17817,N_8684,N_8406);
nand U17818 (N_17818,N_9669,N_10579);
and U17819 (N_17819,N_9524,N_11936);
and U17820 (N_17820,N_9459,N_10408);
nor U17821 (N_17821,N_6327,N_8277);
nor U17822 (N_17822,N_8760,N_8654);
nor U17823 (N_17823,N_8931,N_9660);
nor U17824 (N_17824,N_9752,N_12233);
and U17825 (N_17825,N_9286,N_8376);
or U17826 (N_17826,N_9461,N_10426);
nand U17827 (N_17827,N_10273,N_10735);
nand U17828 (N_17828,N_8233,N_9590);
nor U17829 (N_17829,N_11377,N_9758);
nand U17830 (N_17830,N_10776,N_10169);
or U17831 (N_17831,N_9798,N_12278);
nor U17832 (N_17832,N_7545,N_12284);
nand U17833 (N_17833,N_7329,N_8821);
nand U17834 (N_17834,N_11462,N_8606);
nor U17835 (N_17835,N_7882,N_6555);
nand U17836 (N_17836,N_12158,N_7135);
or U17837 (N_17837,N_11682,N_6438);
nor U17838 (N_17838,N_8558,N_7715);
nand U17839 (N_17839,N_10203,N_10589);
nor U17840 (N_17840,N_9019,N_10762);
nor U17841 (N_17841,N_6655,N_9420);
and U17842 (N_17842,N_7416,N_9713);
and U17843 (N_17843,N_8638,N_10323);
nand U17844 (N_17844,N_8185,N_11583);
or U17845 (N_17845,N_7529,N_7135);
or U17846 (N_17846,N_11879,N_9645);
and U17847 (N_17847,N_9545,N_9527);
nand U17848 (N_17848,N_7791,N_12002);
nand U17849 (N_17849,N_8422,N_10215);
and U17850 (N_17850,N_10935,N_8867);
or U17851 (N_17851,N_9362,N_11099);
or U17852 (N_17852,N_9997,N_11120);
or U17853 (N_17853,N_11905,N_7673);
and U17854 (N_17854,N_10359,N_11193);
nand U17855 (N_17855,N_9715,N_10968);
nand U17856 (N_17856,N_7206,N_9496);
nand U17857 (N_17857,N_7064,N_9759);
xnor U17858 (N_17858,N_9320,N_8041);
nand U17859 (N_17859,N_6589,N_7326);
and U17860 (N_17860,N_7482,N_11851);
nor U17861 (N_17861,N_11972,N_7964);
or U17862 (N_17862,N_9029,N_7073);
nand U17863 (N_17863,N_9378,N_6562);
and U17864 (N_17864,N_7641,N_6700);
nand U17865 (N_17865,N_8038,N_10502);
nand U17866 (N_17866,N_11450,N_8605);
nand U17867 (N_17867,N_6587,N_8615);
and U17868 (N_17868,N_10374,N_11671);
nand U17869 (N_17869,N_8030,N_8137);
nor U17870 (N_17870,N_11561,N_6646);
nand U17871 (N_17871,N_8834,N_12336);
nand U17872 (N_17872,N_10923,N_11827);
or U17873 (N_17873,N_10412,N_9467);
nand U17874 (N_17874,N_9850,N_11992);
nand U17875 (N_17875,N_8177,N_11459);
or U17876 (N_17876,N_9858,N_7589);
nand U17877 (N_17877,N_12424,N_8566);
or U17878 (N_17878,N_9275,N_7722);
xor U17879 (N_17879,N_12143,N_9566);
and U17880 (N_17880,N_6703,N_8715);
or U17881 (N_17881,N_9527,N_9850);
and U17882 (N_17882,N_11046,N_10947);
or U17883 (N_17883,N_10115,N_8879);
nand U17884 (N_17884,N_7391,N_10347);
or U17885 (N_17885,N_7837,N_8223);
nor U17886 (N_17886,N_12345,N_10160);
nor U17887 (N_17887,N_7974,N_6355);
or U17888 (N_17888,N_8322,N_11552);
or U17889 (N_17889,N_10195,N_8185);
or U17890 (N_17890,N_8312,N_7434);
and U17891 (N_17891,N_8214,N_9947);
or U17892 (N_17892,N_10855,N_11274);
nor U17893 (N_17893,N_8847,N_7490);
nand U17894 (N_17894,N_12157,N_11899);
nand U17895 (N_17895,N_11651,N_6843);
and U17896 (N_17896,N_11541,N_9673);
and U17897 (N_17897,N_7185,N_6942);
nand U17898 (N_17898,N_10706,N_10337);
or U17899 (N_17899,N_9094,N_12261);
nor U17900 (N_17900,N_7539,N_8388);
nor U17901 (N_17901,N_6262,N_10343);
nor U17902 (N_17902,N_6346,N_8725);
nand U17903 (N_17903,N_10313,N_8275);
nand U17904 (N_17904,N_7260,N_8789);
nand U17905 (N_17905,N_11269,N_10982);
and U17906 (N_17906,N_6959,N_8384);
and U17907 (N_17907,N_11206,N_8368);
xnor U17908 (N_17908,N_7973,N_8232);
or U17909 (N_17909,N_10496,N_6610);
nand U17910 (N_17910,N_12299,N_8828);
nor U17911 (N_17911,N_6269,N_8591);
nand U17912 (N_17912,N_8228,N_8131);
or U17913 (N_17913,N_11430,N_11678);
nor U17914 (N_17914,N_11242,N_8037);
or U17915 (N_17915,N_8238,N_11628);
or U17916 (N_17916,N_7137,N_10374);
and U17917 (N_17917,N_6474,N_7433);
and U17918 (N_17918,N_10230,N_8499);
or U17919 (N_17919,N_11759,N_10624);
nand U17920 (N_17920,N_8696,N_9690);
or U17921 (N_17921,N_9828,N_10100);
nand U17922 (N_17922,N_6296,N_7385);
or U17923 (N_17923,N_10273,N_11534);
nor U17924 (N_17924,N_8066,N_7148);
nand U17925 (N_17925,N_8323,N_8291);
nand U17926 (N_17926,N_12062,N_12085);
nor U17927 (N_17927,N_9309,N_10575);
nand U17928 (N_17928,N_10301,N_8441);
and U17929 (N_17929,N_9528,N_11896);
nand U17930 (N_17930,N_7277,N_7673);
or U17931 (N_17931,N_12462,N_10648);
or U17932 (N_17932,N_8450,N_8641);
and U17933 (N_17933,N_11069,N_12078);
and U17934 (N_17934,N_11744,N_7227);
and U17935 (N_17935,N_10436,N_7249);
and U17936 (N_17936,N_7286,N_9350);
or U17937 (N_17937,N_7900,N_9091);
nor U17938 (N_17938,N_7114,N_7065);
nor U17939 (N_17939,N_7094,N_8220);
nor U17940 (N_17940,N_9165,N_8225);
nor U17941 (N_17941,N_8981,N_8997);
or U17942 (N_17942,N_7986,N_12291);
or U17943 (N_17943,N_11269,N_12220);
and U17944 (N_17944,N_12366,N_10425);
nand U17945 (N_17945,N_10360,N_11698);
or U17946 (N_17946,N_9712,N_8368);
and U17947 (N_17947,N_11958,N_11215);
and U17948 (N_17948,N_8943,N_9757);
nand U17949 (N_17949,N_9103,N_9819);
or U17950 (N_17950,N_11313,N_9210);
and U17951 (N_17951,N_12474,N_6570);
or U17952 (N_17952,N_7847,N_9091);
and U17953 (N_17953,N_12309,N_10575);
and U17954 (N_17954,N_8305,N_6684);
nor U17955 (N_17955,N_6830,N_11895);
nor U17956 (N_17956,N_11000,N_10859);
and U17957 (N_17957,N_9496,N_11572);
nand U17958 (N_17958,N_11296,N_11376);
or U17959 (N_17959,N_6563,N_10196);
nor U17960 (N_17960,N_11923,N_11043);
and U17961 (N_17961,N_10081,N_6895);
nor U17962 (N_17962,N_7105,N_8251);
nand U17963 (N_17963,N_8813,N_10743);
or U17964 (N_17964,N_11359,N_11404);
and U17965 (N_17965,N_12101,N_9433);
nand U17966 (N_17966,N_7515,N_7009);
xnor U17967 (N_17967,N_11449,N_10441);
or U17968 (N_17968,N_9075,N_9466);
nand U17969 (N_17969,N_10024,N_9530);
or U17970 (N_17970,N_7687,N_9724);
nand U17971 (N_17971,N_11690,N_7232);
nand U17972 (N_17972,N_8081,N_8575);
and U17973 (N_17973,N_9165,N_8735);
and U17974 (N_17974,N_10280,N_8839);
and U17975 (N_17975,N_7790,N_6315);
and U17976 (N_17976,N_10705,N_10985);
or U17977 (N_17977,N_11219,N_11581);
nor U17978 (N_17978,N_10677,N_11233);
and U17979 (N_17979,N_8006,N_8013);
and U17980 (N_17980,N_8927,N_8676);
nor U17981 (N_17981,N_6842,N_7723);
or U17982 (N_17982,N_8981,N_10550);
nor U17983 (N_17983,N_9450,N_7708);
nor U17984 (N_17984,N_11038,N_8156);
nand U17985 (N_17985,N_6493,N_8491);
nor U17986 (N_17986,N_10488,N_12246);
nand U17987 (N_17987,N_9956,N_11066);
nor U17988 (N_17988,N_8424,N_6432);
and U17989 (N_17989,N_7882,N_11548);
or U17990 (N_17990,N_7539,N_9007);
or U17991 (N_17991,N_8431,N_6293);
nor U17992 (N_17992,N_11425,N_9933);
nor U17993 (N_17993,N_10529,N_10367);
nor U17994 (N_17994,N_7341,N_12065);
or U17995 (N_17995,N_11801,N_11118);
nand U17996 (N_17996,N_8902,N_10112);
nor U17997 (N_17997,N_9054,N_11479);
nor U17998 (N_17998,N_10097,N_6946);
and U17999 (N_17999,N_11766,N_7773);
or U18000 (N_18000,N_9222,N_12413);
nor U18001 (N_18001,N_10619,N_9753);
or U18002 (N_18002,N_8029,N_8663);
and U18003 (N_18003,N_6764,N_9038);
or U18004 (N_18004,N_9479,N_6392);
nand U18005 (N_18005,N_12191,N_8633);
or U18006 (N_18006,N_10212,N_8626);
nand U18007 (N_18007,N_9761,N_10090);
nand U18008 (N_18008,N_7685,N_6910);
nor U18009 (N_18009,N_12459,N_7190);
nor U18010 (N_18010,N_11308,N_10459);
nand U18011 (N_18011,N_7585,N_11734);
nor U18012 (N_18012,N_12059,N_7380);
or U18013 (N_18013,N_12255,N_11337);
and U18014 (N_18014,N_11854,N_12479);
nand U18015 (N_18015,N_7390,N_7995);
nand U18016 (N_18016,N_8511,N_8348);
nand U18017 (N_18017,N_6259,N_12425);
nand U18018 (N_18018,N_11571,N_7248);
or U18019 (N_18019,N_8365,N_9193);
nand U18020 (N_18020,N_6908,N_10410);
or U18021 (N_18021,N_10323,N_7772);
or U18022 (N_18022,N_6377,N_11059);
nor U18023 (N_18023,N_7448,N_11473);
or U18024 (N_18024,N_10042,N_7035);
or U18025 (N_18025,N_7942,N_8035);
or U18026 (N_18026,N_8503,N_11254);
or U18027 (N_18027,N_9094,N_12395);
nand U18028 (N_18028,N_8074,N_9926);
or U18029 (N_18029,N_7736,N_7212);
or U18030 (N_18030,N_7998,N_10315);
or U18031 (N_18031,N_10113,N_6993);
or U18032 (N_18032,N_6636,N_10729);
xor U18033 (N_18033,N_6313,N_11337);
nor U18034 (N_18034,N_10333,N_9309);
nor U18035 (N_18035,N_7346,N_6438);
nand U18036 (N_18036,N_7102,N_12190);
nand U18037 (N_18037,N_10608,N_11182);
or U18038 (N_18038,N_10234,N_8926);
or U18039 (N_18039,N_12384,N_8027);
nor U18040 (N_18040,N_7428,N_10284);
nand U18041 (N_18041,N_8875,N_10112);
or U18042 (N_18042,N_9626,N_10521);
or U18043 (N_18043,N_7622,N_6260);
nand U18044 (N_18044,N_6806,N_12227);
nand U18045 (N_18045,N_11977,N_11454);
or U18046 (N_18046,N_9116,N_11669);
nor U18047 (N_18047,N_7517,N_10482);
nand U18048 (N_18048,N_8726,N_7394);
nor U18049 (N_18049,N_10463,N_11127);
nand U18050 (N_18050,N_11655,N_9368);
or U18051 (N_18051,N_9275,N_6872);
or U18052 (N_18052,N_11270,N_11876);
nor U18053 (N_18053,N_10430,N_9605);
and U18054 (N_18054,N_6906,N_8260);
nand U18055 (N_18055,N_7454,N_8027);
nor U18056 (N_18056,N_9575,N_10403);
and U18057 (N_18057,N_9793,N_10197);
or U18058 (N_18058,N_6944,N_9285);
and U18059 (N_18059,N_10742,N_9961);
or U18060 (N_18060,N_7329,N_11643);
and U18061 (N_18061,N_11953,N_7449);
or U18062 (N_18062,N_11177,N_9214);
nor U18063 (N_18063,N_10555,N_11993);
nand U18064 (N_18064,N_8751,N_12244);
nor U18065 (N_18065,N_6477,N_11518);
nor U18066 (N_18066,N_8530,N_10040);
or U18067 (N_18067,N_6796,N_6627);
or U18068 (N_18068,N_9781,N_11457);
nor U18069 (N_18069,N_7539,N_12389);
and U18070 (N_18070,N_7943,N_9007);
nor U18071 (N_18071,N_10007,N_11077);
or U18072 (N_18072,N_6632,N_7583);
and U18073 (N_18073,N_11377,N_8848);
nor U18074 (N_18074,N_8751,N_11999);
or U18075 (N_18075,N_12367,N_8041);
or U18076 (N_18076,N_11953,N_9756);
or U18077 (N_18077,N_7358,N_9008);
nand U18078 (N_18078,N_10924,N_11251);
nand U18079 (N_18079,N_8123,N_7764);
nand U18080 (N_18080,N_9193,N_10911);
or U18081 (N_18081,N_10832,N_11268);
or U18082 (N_18082,N_9304,N_11295);
or U18083 (N_18083,N_6356,N_6360);
or U18084 (N_18084,N_10302,N_8011);
nand U18085 (N_18085,N_6696,N_7202);
and U18086 (N_18086,N_6887,N_12233);
or U18087 (N_18087,N_6644,N_12292);
nor U18088 (N_18088,N_9593,N_10552);
nor U18089 (N_18089,N_10660,N_12011);
or U18090 (N_18090,N_6865,N_11821);
nor U18091 (N_18091,N_9485,N_12215);
nor U18092 (N_18092,N_7865,N_11519);
nor U18093 (N_18093,N_8424,N_11862);
nor U18094 (N_18094,N_8656,N_8114);
nand U18095 (N_18095,N_7402,N_7983);
nand U18096 (N_18096,N_9843,N_8065);
and U18097 (N_18097,N_11419,N_9958);
or U18098 (N_18098,N_7706,N_7833);
and U18099 (N_18099,N_8385,N_7975);
nor U18100 (N_18100,N_10324,N_7684);
nand U18101 (N_18101,N_6769,N_11298);
nor U18102 (N_18102,N_11568,N_10697);
and U18103 (N_18103,N_8238,N_12453);
and U18104 (N_18104,N_7255,N_9091);
nand U18105 (N_18105,N_12372,N_10445);
or U18106 (N_18106,N_10196,N_6690);
or U18107 (N_18107,N_9277,N_8898);
nor U18108 (N_18108,N_12303,N_8940);
nor U18109 (N_18109,N_7801,N_11139);
nor U18110 (N_18110,N_7342,N_8048);
nor U18111 (N_18111,N_8858,N_12346);
nand U18112 (N_18112,N_6558,N_7433);
nor U18113 (N_18113,N_12278,N_8800);
nor U18114 (N_18114,N_10712,N_8093);
and U18115 (N_18115,N_8458,N_12468);
or U18116 (N_18116,N_10888,N_9395);
nand U18117 (N_18117,N_8934,N_11554);
or U18118 (N_18118,N_8631,N_6709);
nor U18119 (N_18119,N_10057,N_9290);
or U18120 (N_18120,N_6413,N_10801);
or U18121 (N_18121,N_8694,N_7650);
nand U18122 (N_18122,N_12238,N_6397);
and U18123 (N_18123,N_12462,N_8249);
or U18124 (N_18124,N_9739,N_10008);
and U18125 (N_18125,N_6404,N_8596);
nor U18126 (N_18126,N_7815,N_9141);
nor U18127 (N_18127,N_7881,N_12353);
or U18128 (N_18128,N_6267,N_7615);
nor U18129 (N_18129,N_8946,N_11752);
nor U18130 (N_18130,N_7040,N_12315);
and U18131 (N_18131,N_9461,N_7578);
nand U18132 (N_18132,N_11130,N_6855);
nand U18133 (N_18133,N_10143,N_6717);
nand U18134 (N_18134,N_11063,N_10579);
nand U18135 (N_18135,N_12078,N_10163);
nor U18136 (N_18136,N_9826,N_6942);
and U18137 (N_18137,N_6779,N_8487);
and U18138 (N_18138,N_12240,N_8826);
or U18139 (N_18139,N_9918,N_7265);
nor U18140 (N_18140,N_7296,N_8330);
or U18141 (N_18141,N_8377,N_6474);
nor U18142 (N_18142,N_8139,N_10737);
nand U18143 (N_18143,N_9056,N_7616);
and U18144 (N_18144,N_9982,N_11774);
xnor U18145 (N_18145,N_7154,N_10964);
and U18146 (N_18146,N_7954,N_7915);
and U18147 (N_18147,N_10035,N_12199);
and U18148 (N_18148,N_6645,N_9975);
nand U18149 (N_18149,N_11671,N_11854);
nand U18150 (N_18150,N_6391,N_9388);
nand U18151 (N_18151,N_11201,N_6477);
and U18152 (N_18152,N_11871,N_9420);
nor U18153 (N_18153,N_9119,N_6591);
nand U18154 (N_18154,N_11752,N_6768);
and U18155 (N_18155,N_7674,N_11898);
nand U18156 (N_18156,N_11228,N_12448);
and U18157 (N_18157,N_8318,N_8243);
nor U18158 (N_18158,N_11737,N_8195);
or U18159 (N_18159,N_11259,N_10482);
nor U18160 (N_18160,N_8066,N_10345);
or U18161 (N_18161,N_9419,N_7355);
and U18162 (N_18162,N_8473,N_6295);
and U18163 (N_18163,N_6584,N_8283);
nor U18164 (N_18164,N_10343,N_11911);
and U18165 (N_18165,N_9260,N_10027);
nand U18166 (N_18166,N_10290,N_8434);
nand U18167 (N_18167,N_8355,N_7304);
and U18168 (N_18168,N_10692,N_9481);
or U18169 (N_18169,N_8977,N_11287);
and U18170 (N_18170,N_6253,N_11377);
nand U18171 (N_18171,N_7749,N_7268);
nor U18172 (N_18172,N_9589,N_9444);
nor U18173 (N_18173,N_9581,N_11741);
or U18174 (N_18174,N_10967,N_8659);
or U18175 (N_18175,N_10622,N_8487);
or U18176 (N_18176,N_11998,N_11967);
and U18177 (N_18177,N_9707,N_12192);
or U18178 (N_18178,N_11854,N_7405);
and U18179 (N_18179,N_11999,N_8821);
nor U18180 (N_18180,N_11011,N_7766);
and U18181 (N_18181,N_7366,N_11108);
or U18182 (N_18182,N_10259,N_7914);
or U18183 (N_18183,N_10462,N_7393);
nor U18184 (N_18184,N_12099,N_10741);
or U18185 (N_18185,N_8957,N_10524);
xnor U18186 (N_18186,N_12016,N_6629);
or U18187 (N_18187,N_9737,N_8265);
nand U18188 (N_18188,N_8280,N_8933);
and U18189 (N_18189,N_11355,N_10524);
or U18190 (N_18190,N_8939,N_6363);
nand U18191 (N_18191,N_7398,N_9815);
or U18192 (N_18192,N_7158,N_9825);
and U18193 (N_18193,N_6561,N_11261);
nor U18194 (N_18194,N_8468,N_11727);
nor U18195 (N_18195,N_8140,N_10868);
nand U18196 (N_18196,N_8953,N_9623);
nand U18197 (N_18197,N_10015,N_10202);
or U18198 (N_18198,N_8212,N_7098);
nand U18199 (N_18199,N_7121,N_10940);
or U18200 (N_18200,N_10476,N_8289);
nand U18201 (N_18201,N_7852,N_12489);
nand U18202 (N_18202,N_6712,N_11103);
nor U18203 (N_18203,N_10350,N_9142);
or U18204 (N_18204,N_10963,N_6546);
or U18205 (N_18205,N_7172,N_10330);
nand U18206 (N_18206,N_7965,N_10410);
or U18207 (N_18207,N_9204,N_10204);
or U18208 (N_18208,N_7220,N_6776);
nand U18209 (N_18209,N_8613,N_7729);
nand U18210 (N_18210,N_9763,N_6827);
nand U18211 (N_18211,N_10985,N_6816);
or U18212 (N_18212,N_11969,N_12215);
and U18213 (N_18213,N_8717,N_12276);
and U18214 (N_18214,N_10682,N_10693);
or U18215 (N_18215,N_8844,N_6395);
nor U18216 (N_18216,N_7170,N_12357);
nand U18217 (N_18217,N_11118,N_12025);
nand U18218 (N_18218,N_8406,N_8320);
nor U18219 (N_18219,N_7008,N_9223);
nand U18220 (N_18220,N_10700,N_11571);
nand U18221 (N_18221,N_8438,N_8220);
nand U18222 (N_18222,N_7032,N_10049);
nor U18223 (N_18223,N_10514,N_7610);
nor U18224 (N_18224,N_11542,N_11377);
and U18225 (N_18225,N_8332,N_7900);
and U18226 (N_18226,N_11930,N_12073);
and U18227 (N_18227,N_6310,N_9683);
or U18228 (N_18228,N_9990,N_11527);
nand U18229 (N_18229,N_7468,N_11231);
nor U18230 (N_18230,N_9269,N_7995);
or U18231 (N_18231,N_12065,N_6466);
nand U18232 (N_18232,N_8579,N_12352);
xnor U18233 (N_18233,N_12349,N_10293);
nand U18234 (N_18234,N_7155,N_8308);
nand U18235 (N_18235,N_8573,N_6304);
or U18236 (N_18236,N_8940,N_6746);
or U18237 (N_18237,N_6593,N_10563);
xnor U18238 (N_18238,N_7127,N_10539);
nand U18239 (N_18239,N_7844,N_10278);
nand U18240 (N_18240,N_6599,N_11460);
or U18241 (N_18241,N_6659,N_12316);
nand U18242 (N_18242,N_8166,N_7593);
nand U18243 (N_18243,N_8257,N_9038);
nor U18244 (N_18244,N_10791,N_8951);
nand U18245 (N_18245,N_10334,N_12282);
nand U18246 (N_18246,N_6716,N_10228);
nand U18247 (N_18247,N_7189,N_7641);
or U18248 (N_18248,N_7508,N_11799);
or U18249 (N_18249,N_7940,N_10214);
or U18250 (N_18250,N_8652,N_10931);
nand U18251 (N_18251,N_6668,N_10936);
or U18252 (N_18252,N_12395,N_11589);
and U18253 (N_18253,N_11591,N_7105);
or U18254 (N_18254,N_7887,N_9238);
nand U18255 (N_18255,N_9315,N_7353);
or U18256 (N_18256,N_11177,N_11295);
nand U18257 (N_18257,N_6464,N_9458);
and U18258 (N_18258,N_9965,N_9913);
or U18259 (N_18259,N_7817,N_10376);
and U18260 (N_18260,N_11932,N_11904);
nand U18261 (N_18261,N_10932,N_6254);
nand U18262 (N_18262,N_7825,N_11909);
nand U18263 (N_18263,N_6766,N_8620);
and U18264 (N_18264,N_12266,N_11998);
nor U18265 (N_18265,N_11825,N_7555);
nand U18266 (N_18266,N_9934,N_11734);
and U18267 (N_18267,N_11967,N_11210);
nand U18268 (N_18268,N_12382,N_8580);
or U18269 (N_18269,N_9241,N_11724);
nand U18270 (N_18270,N_12296,N_10562);
nand U18271 (N_18271,N_8988,N_11060);
or U18272 (N_18272,N_9901,N_8848);
and U18273 (N_18273,N_11532,N_11371);
nor U18274 (N_18274,N_8107,N_11378);
nand U18275 (N_18275,N_9689,N_8290);
or U18276 (N_18276,N_9517,N_10819);
or U18277 (N_18277,N_6850,N_6727);
and U18278 (N_18278,N_9868,N_10845);
and U18279 (N_18279,N_10005,N_9288);
or U18280 (N_18280,N_7947,N_11187);
and U18281 (N_18281,N_9909,N_11277);
nand U18282 (N_18282,N_10531,N_8680);
and U18283 (N_18283,N_9073,N_11255);
and U18284 (N_18284,N_8430,N_8710);
nand U18285 (N_18285,N_7389,N_9827);
and U18286 (N_18286,N_7835,N_7235);
xnor U18287 (N_18287,N_11230,N_10195);
or U18288 (N_18288,N_9754,N_7867);
nand U18289 (N_18289,N_9929,N_9955);
or U18290 (N_18290,N_12304,N_12007);
or U18291 (N_18291,N_9798,N_11798);
nand U18292 (N_18292,N_11326,N_9540);
or U18293 (N_18293,N_12329,N_8365);
or U18294 (N_18294,N_8041,N_7220);
or U18295 (N_18295,N_7554,N_10720);
and U18296 (N_18296,N_6575,N_7736);
or U18297 (N_18297,N_6977,N_12262);
nor U18298 (N_18298,N_7460,N_12421);
or U18299 (N_18299,N_8712,N_7705);
or U18300 (N_18300,N_10385,N_10548);
or U18301 (N_18301,N_9994,N_10942);
or U18302 (N_18302,N_7239,N_8530);
nor U18303 (N_18303,N_11678,N_9209);
nor U18304 (N_18304,N_12406,N_6760);
nand U18305 (N_18305,N_7872,N_9221);
and U18306 (N_18306,N_7806,N_11555);
nand U18307 (N_18307,N_10691,N_7594);
or U18308 (N_18308,N_11810,N_12410);
nor U18309 (N_18309,N_8387,N_10313);
or U18310 (N_18310,N_7783,N_12251);
or U18311 (N_18311,N_6697,N_11465);
and U18312 (N_18312,N_10928,N_10801);
nor U18313 (N_18313,N_11687,N_11712);
nor U18314 (N_18314,N_11182,N_8778);
nor U18315 (N_18315,N_10854,N_6438);
nor U18316 (N_18316,N_7443,N_10781);
nor U18317 (N_18317,N_9524,N_12496);
nand U18318 (N_18318,N_9053,N_10803);
and U18319 (N_18319,N_10866,N_6807);
or U18320 (N_18320,N_11508,N_12491);
and U18321 (N_18321,N_9679,N_11503);
or U18322 (N_18322,N_10997,N_11406);
xor U18323 (N_18323,N_11978,N_7160);
or U18324 (N_18324,N_10774,N_12393);
nand U18325 (N_18325,N_10566,N_6821);
and U18326 (N_18326,N_7113,N_7861);
and U18327 (N_18327,N_11259,N_11349);
nand U18328 (N_18328,N_11281,N_10250);
nand U18329 (N_18329,N_6348,N_10497);
nand U18330 (N_18330,N_10860,N_9749);
nand U18331 (N_18331,N_10823,N_7088);
nand U18332 (N_18332,N_11152,N_11586);
nand U18333 (N_18333,N_9512,N_6291);
or U18334 (N_18334,N_9027,N_9820);
or U18335 (N_18335,N_11218,N_7041);
nor U18336 (N_18336,N_10834,N_8217);
nor U18337 (N_18337,N_10090,N_11296);
nand U18338 (N_18338,N_8068,N_8471);
or U18339 (N_18339,N_9944,N_11265);
nor U18340 (N_18340,N_9618,N_10379);
nor U18341 (N_18341,N_7002,N_10081);
and U18342 (N_18342,N_7639,N_6769);
nand U18343 (N_18343,N_9230,N_8143);
or U18344 (N_18344,N_10659,N_11862);
nand U18345 (N_18345,N_7404,N_8371);
nor U18346 (N_18346,N_10882,N_11306);
and U18347 (N_18347,N_10065,N_10448);
nand U18348 (N_18348,N_9233,N_10245);
or U18349 (N_18349,N_11551,N_11860);
nand U18350 (N_18350,N_7276,N_8775);
nor U18351 (N_18351,N_9868,N_6329);
and U18352 (N_18352,N_11735,N_10301);
and U18353 (N_18353,N_9836,N_8401);
or U18354 (N_18354,N_10702,N_8765);
or U18355 (N_18355,N_8564,N_9661);
nor U18356 (N_18356,N_9951,N_7729);
nor U18357 (N_18357,N_11709,N_6883);
nand U18358 (N_18358,N_10279,N_11502);
nand U18359 (N_18359,N_6462,N_11720);
nor U18360 (N_18360,N_11191,N_7588);
nand U18361 (N_18361,N_12067,N_12320);
or U18362 (N_18362,N_12220,N_7479);
nor U18363 (N_18363,N_11889,N_6810);
nand U18364 (N_18364,N_8879,N_9905);
nand U18365 (N_18365,N_11544,N_6913);
nor U18366 (N_18366,N_7229,N_9103);
nand U18367 (N_18367,N_8109,N_7999);
nand U18368 (N_18368,N_8495,N_11639);
or U18369 (N_18369,N_9489,N_6451);
nor U18370 (N_18370,N_11160,N_7030);
nand U18371 (N_18371,N_7025,N_11277);
nand U18372 (N_18372,N_8422,N_6913);
nor U18373 (N_18373,N_10112,N_10240);
or U18374 (N_18374,N_9576,N_9695);
and U18375 (N_18375,N_11204,N_11878);
xnor U18376 (N_18376,N_7609,N_12356);
nand U18377 (N_18377,N_10347,N_10461);
or U18378 (N_18378,N_11722,N_7699);
nor U18379 (N_18379,N_12267,N_12381);
nand U18380 (N_18380,N_8229,N_11516);
or U18381 (N_18381,N_10260,N_7216);
or U18382 (N_18382,N_7883,N_9069);
and U18383 (N_18383,N_8770,N_6895);
and U18384 (N_18384,N_9508,N_11619);
and U18385 (N_18385,N_6271,N_6274);
or U18386 (N_18386,N_8806,N_8620);
nor U18387 (N_18387,N_11986,N_9754);
nor U18388 (N_18388,N_8595,N_7321);
nor U18389 (N_18389,N_6460,N_10570);
nand U18390 (N_18390,N_12068,N_8069);
or U18391 (N_18391,N_12479,N_6351);
nor U18392 (N_18392,N_10160,N_9169);
nand U18393 (N_18393,N_10375,N_10248);
or U18394 (N_18394,N_7368,N_10643);
nor U18395 (N_18395,N_9271,N_11569);
nand U18396 (N_18396,N_11738,N_8190);
or U18397 (N_18397,N_9149,N_11808);
or U18398 (N_18398,N_6825,N_7718);
nand U18399 (N_18399,N_12326,N_7917);
nor U18400 (N_18400,N_7171,N_6594);
xnor U18401 (N_18401,N_8601,N_9463);
nand U18402 (N_18402,N_9889,N_9795);
nand U18403 (N_18403,N_10512,N_6879);
or U18404 (N_18404,N_10729,N_7274);
nor U18405 (N_18405,N_10829,N_8586);
nand U18406 (N_18406,N_9500,N_10013);
nor U18407 (N_18407,N_6272,N_8388);
or U18408 (N_18408,N_9321,N_6516);
or U18409 (N_18409,N_7282,N_11175);
and U18410 (N_18410,N_9329,N_10584);
nand U18411 (N_18411,N_11545,N_9256);
or U18412 (N_18412,N_9911,N_8577);
nand U18413 (N_18413,N_7845,N_11566);
or U18414 (N_18414,N_7314,N_8284);
and U18415 (N_18415,N_7740,N_7898);
nor U18416 (N_18416,N_10100,N_7624);
nand U18417 (N_18417,N_9333,N_10293);
and U18418 (N_18418,N_11231,N_7394);
nor U18419 (N_18419,N_7880,N_11138);
or U18420 (N_18420,N_6785,N_6403);
or U18421 (N_18421,N_12448,N_8404);
or U18422 (N_18422,N_9670,N_10695);
or U18423 (N_18423,N_10122,N_12334);
nand U18424 (N_18424,N_9036,N_9400);
and U18425 (N_18425,N_11871,N_9763);
nand U18426 (N_18426,N_11224,N_7078);
xor U18427 (N_18427,N_10063,N_12456);
nor U18428 (N_18428,N_8016,N_7629);
nor U18429 (N_18429,N_11785,N_8819);
nor U18430 (N_18430,N_7692,N_10527);
or U18431 (N_18431,N_6692,N_10655);
nor U18432 (N_18432,N_8861,N_7328);
nor U18433 (N_18433,N_9909,N_9466);
nand U18434 (N_18434,N_6722,N_8972);
or U18435 (N_18435,N_10317,N_9563);
or U18436 (N_18436,N_10569,N_7893);
or U18437 (N_18437,N_10710,N_7366);
nand U18438 (N_18438,N_10489,N_8335);
and U18439 (N_18439,N_11967,N_11788);
nand U18440 (N_18440,N_6512,N_9503);
nand U18441 (N_18441,N_6465,N_11695);
nor U18442 (N_18442,N_9975,N_7584);
or U18443 (N_18443,N_11653,N_10399);
nor U18444 (N_18444,N_9828,N_8819);
nor U18445 (N_18445,N_10441,N_7609);
nor U18446 (N_18446,N_10098,N_11802);
or U18447 (N_18447,N_11431,N_7191);
nor U18448 (N_18448,N_10773,N_7520);
or U18449 (N_18449,N_9718,N_12072);
nor U18450 (N_18450,N_7329,N_10016);
nor U18451 (N_18451,N_10707,N_11087);
nand U18452 (N_18452,N_6351,N_12055);
and U18453 (N_18453,N_7551,N_6987);
nand U18454 (N_18454,N_9921,N_10915);
or U18455 (N_18455,N_9291,N_8724);
nand U18456 (N_18456,N_10523,N_9902);
or U18457 (N_18457,N_7465,N_8188);
and U18458 (N_18458,N_6320,N_11661);
nor U18459 (N_18459,N_12034,N_12431);
nor U18460 (N_18460,N_6580,N_8151);
nand U18461 (N_18461,N_6542,N_8928);
and U18462 (N_18462,N_11419,N_6900);
nand U18463 (N_18463,N_7779,N_6672);
nand U18464 (N_18464,N_10360,N_10708);
nor U18465 (N_18465,N_11223,N_9702);
nand U18466 (N_18466,N_7897,N_12240);
and U18467 (N_18467,N_7506,N_8383);
or U18468 (N_18468,N_7085,N_7201);
or U18469 (N_18469,N_9064,N_8573);
and U18470 (N_18470,N_12325,N_7657);
nor U18471 (N_18471,N_10939,N_9827);
and U18472 (N_18472,N_7186,N_8583);
and U18473 (N_18473,N_8243,N_8542);
or U18474 (N_18474,N_7567,N_8778);
or U18475 (N_18475,N_7967,N_9909);
or U18476 (N_18476,N_10460,N_10629);
nand U18477 (N_18477,N_12266,N_11080);
and U18478 (N_18478,N_9269,N_11355);
or U18479 (N_18479,N_8553,N_10252);
nand U18480 (N_18480,N_6589,N_9421);
nand U18481 (N_18481,N_6600,N_12078);
or U18482 (N_18482,N_9930,N_8758);
and U18483 (N_18483,N_11165,N_11997);
or U18484 (N_18484,N_8059,N_8522);
nand U18485 (N_18485,N_7840,N_10230);
or U18486 (N_18486,N_9574,N_7879);
and U18487 (N_18487,N_10638,N_9192);
and U18488 (N_18488,N_8549,N_9626);
nand U18489 (N_18489,N_9308,N_9921);
nor U18490 (N_18490,N_7032,N_8387);
and U18491 (N_18491,N_11112,N_9086);
and U18492 (N_18492,N_10881,N_9070);
and U18493 (N_18493,N_8817,N_7510);
and U18494 (N_18494,N_6829,N_11016);
or U18495 (N_18495,N_6417,N_11140);
or U18496 (N_18496,N_7649,N_7841);
nand U18497 (N_18497,N_8023,N_8154);
and U18498 (N_18498,N_8529,N_6543);
or U18499 (N_18499,N_11525,N_12272);
nand U18500 (N_18500,N_6275,N_11308);
nor U18501 (N_18501,N_10750,N_10216);
nand U18502 (N_18502,N_10586,N_9755);
or U18503 (N_18503,N_10991,N_7498);
and U18504 (N_18504,N_11713,N_6543);
or U18505 (N_18505,N_11199,N_6388);
nor U18506 (N_18506,N_7822,N_7268);
and U18507 (N_18507,N_8212,N_9253);
nor U18508 (N_18508,N_8244,N_11793);
and U18509 (N_18509,N_10801,N_12111);
and U18510 (N_18510,N_10741,N_9617);
and U18511 (N_18511,N_9211,N_9221);
nor U18512 (N_18512,N_11279,N_10646);
xnor U18513 (N_18513,N_8469,N_6954);
nand U18514 (N_18514,N_10718,N_10889);
or U18515 (N_18515,N_10294,N_12043);
nand U18516 (N_18516,N_10198,N_10459);
and U18517 (N_18517,N_7812,N_7585);
or U18518 (N_18518,N_9828,N_8856);
and U18519 (N_18519,N_6552,N_10834);
nand U18520 (N_18520,N_8357,N_8865);
nor U18521 (N_18521,N_11629,N_10792);
nor U18522 (N_18522,N_7017,N_11283);
or U18523 (N_18523,N_8261,N_10550);
nor U18524 (N_18524,N_9983,N_8680);
and U18525 (N_18525,N_12250,N_7056);
nand U18526 (N_18526,N_11667,N_10345);
nand U18527 (N_18527,N_9305,N_7629);
and U18528 (N_18528,N_7695,N_10163);
and U18529 (N_18529,N_10004,N_9531);
and U18530 (N_18530,N_7336,N_7271);
xnor U18531 (N_18531,N_6279,N_6581);
or U18532 (N_18532,N_12226,N_10106);
and U18533 (N_18533,N_10700,N_8878);
nor U18534 (N_18534,N_9492,N_6567);
or U18535 (N_18535,N_6260,N_11856);
nor U18536 (N_18536,N_8868,N_11287);
and U18537 (N_18537,N_10756,N_6933);
or U18538 (N_18538,N_7467,N_7523);
nor U18539 (N_18539,N_11870,N_8820);
and U18540 (N_18540,N_7431,N_10960);
nand U18541 (N_18541,N_9642,N_7536);
nand U18542 (N_18542,N_10382,N_11165);
or U18543 (N_18543,N_11357,N_9282);
and U18544 (N_18544,N_10210,N_6570);
or U18545 (N_18545,N_10128,N_7168);
or U18546 (N_18546,N_8868,N_8985);
nand U18547 (N_18547,N_8548,N_12020);
nand U18548 (N_18548,N_12381,N_9087);
nor U18549 (N_18549,N_11998,N_11346);
and U18550 (N_18550,N_11731,N_9953);
nand U18551 (N_18551,N_6934,N_11185);
nor U18552 (N_18552,N_11537,N_8133);
nor U18553 (N_18553,N_12069,N_9647);
or U18554 (N_18554,N_11022,N_6887);
nor U18555 (N_18555,N_10375,N_6727);
and U18556 (N_18556,N_11516,N_10021);
or U18557 (N_18557,N_11803,N_7068);
nand U18558 (N_18558,N_9176,N_10084);
nor U18559 (N_18559,N_11653,N_11721);
and U18560 (N_18560,N_8613,N_9381);
nand U18561 (N_18561,N_7049,N_11980);
nand U18562 (N_18562,N_12379,N_10393);
and U18563 (N_18563,N_11753,N_8408);
or U18564 (N_18564,N_9557,N_11237);
nand U18565 (N_18565,N_11249,N_11356);
xor U18566 (N_18566,N_8456,N_11788);
nor U18567 (N_18567,N_11149,N_10839);
or U18568 (N_18568,N_7756,N_11570);
nand U18569 (N_18569,N_10122,N_10816);
nor U18570 (N_18570,N_11125,N_8474);
nor U18571 (N_18571,N_9350,N_6353);
or U18572 (N_18572,N_8659,N_10715);
or U18573 (N_18573,N_6844,N_6792);
or U18574 (N_18574,N_10218,N_8103);
nor U18575 (N_18575,N_11598,N_12378);
nand U18576 (N_18576,N_8474,N_11491);
and U18577 (N_18577,N_11148,N_7387);
nand U18578 (N_18578,N_8053,N_7870);
xnor U18579 (N_18579,N_12297,N_7637);
or U18580 (N_18580,N_9970,N_10064);
xor U18581 (N_18581,N_9035,N_10321);
nor U18582 (N_18582,N_10024,N_8008);
or U18583 (N_18583,N_12246,N_12280);
or U18584 (N_18584,N_8196,N_9434);
or U18585 (N_18585,N_11390,N_11570);
nor U18586 (N_18586,N_12338,N_7887);
nand U18587 (N_18587,N_7937,N_12289);
and U18588 (N_18588,N_11672,N_7607);
nand U18589 (N_18589,N_6478,N_9074);
and U18590 (N_18590,N_9372,N_7097);
nor U18591 (N_18591,N_8132,N_8432);
nor U18592 (N_18592,N_9848,N_10316);
xor U18593 (N_18593,N_11373,N_10509);
nand U18594 (N_18594,N_7922,N_10241);
nand U18595 (N_18595,N_11692,N_11963);
and U18596 (N_18596,N_7946,N_10068);
and U18597 (N_18597,N_10429,N_11915);
nor U18598 (N_18598,N_11603,N_10199);
nor U18599 (N_18599,N_8666,N_10384);
nand U18600 (N_18600,N_8421,N_12181);
nand U18601 (N_18601,N_8223,N_9202);
and U18602 (N_18602,N_6308,N_7595);
nor U18603 (N_18603,N_6828,N_11126);
or U18604 (N_18604,N_9749,N_9138);
nand U18605 (N_18605,N_6981,N_11374);
nor U18606 (N_18606,N_11797,N_10534);
nand U18607 (N_18607,N_8408,N_7464);
and U18608 (N_18608,N_11272,N_6837);
or U18609 (N_18609,N_10700,N_11073);
and U18610 (N_18610,N_10494,N_12402);
nor U18611 (N_18611,N_10317,N_6628);
or U18612 (N_18612,N_11235,N_10545);
nor U18613 (N_18613,N_11656,N_10489);
nor U18614 (N_18614,N_12383,N_8534);
nor U18615 (N_18615,N_6741,N_12017);
nor U18616 (N_18616,N_6385,N_9573);
nor U18617 (N_18617,N_11312,N_11103);
nand U18618 (N_18618,N_9721,N_12088);
nand U18619 (N_18619,N_7039,N_12139);
and U18620 (N_18620,N_6925,N_12297);
and U18621 (N_18621,N_7311,N_8474);
xnor U18622 (N_18622,N_11799,N_9683);
nor U18623 (N_18623,N_8792,N_11890);
and U18624 (N_18624,N_7971,N_7016);
and U18625 (N_18625,N_10403,N_8137);
nand U18626 (N_18626,N_8643,N_11384);
and U18627 (N_18627,N_9943,N_12196);
nand U18628 (N_18628,N_9149,N_10375);
or U18629 (N_18629,N_9564,N_11171);
and U18630 (N_18630,N_10357,N_11721);
and U18631 (N_18631,N_7158,N_7436);
nor U18632 (N_18632,N_7474,N_9481);
or U18633 (N_18633,N_12309,N_12430);
or U18634 (N_18634,N_8158,N_9475);
or U18635 (N_18635,N_11406,N_7415);
nor U18636 (N_18636,N_11595,N_12208);
nand U18637 (N_18637,N_7980,N_6680);
or U18638 (N_18638,N_9834,N_9670);
nor U18639 (N_18639,N_8013,N_8281);
and U18640 (N_18640,N_7313,N_10397);
and U18641 (N_18641,N_8138,N_6576);
or U18642 (N_18642,N_7284,N_7111);
and U18643 (N_18643,N_6422,N_8433);
nand U18644 (N_18644,N_9312,N_9883);
and U18645 (N_18645,N_8165,N_8110);
nand U18646 (N_18646,N_11780,N_9149);
nand U18647 (N_18647,N_10008,N_7318);
nand U18648 (N_18648,N_9046,N_11567);
nor U18649 (N_18649,N_9233,N_10556);
and U18650 (N_18650,N_11996,N_7634);
and U18651 (N_18651,N_8838,N_9466);
nor U18652 (N_18652,N_8051,N_12067);
and U18653 (N_18653,N_8599,N_9501);
nor U18654 (N_18654,N_9151,N_8045);
or U18655 (N_18655,N_7773,N_8349);
and U18656 (N_18656,N_11900,N_6812);
nand U18657 (N_18657,N_6979,N_11762);
and U18658 (N_18658,N_12374,N_12195);
or U18659 (N_18659,N_8196,N_10530);
nand U18660 (N_18660,N_10026,N_12064);
nor U18661 (N_18661,N_6937,N_10343);
or U18662 (N_18662,N_9473,N_7623);
nand U18663 (N_18663,N_11383,N_10955);
nand U18664 (N_18664,N_7345,N_11070);
nand U18665 (N_18665,N_6446,N_11228);
nand U18666 (N_18666,N_7819,N_11734);
nand U18667 (N_18667,N_7269,N_12141);
nor U18668 (N_18668,N_7379,N_7920);
nand U18669 (N_18669,N_7516,N_11731);
or U18670 (N_18670,N_8962,N_6509);
nand U18671 (N_18671,N_12276,N_7229);
or U18672 (N_18672,N_8687,N_11385);
nor U18673 (N_18673,N_10327,N_6278);
or U18674 (N_18674,N_11098,N_7977);
and U18675 (N_18675,N_9627,N_11481);
nor U18676 (N_18676,N_11518,N_9477);
or U18677 (N_18677,N_6419,N_9796);
and U18678 (N_18678,N_7625,N_6651);
nor U18679 (N_18679,N_10884,N_10417);
and U18680 (N_18680,N_8054,N_9935);
and U18681 (N_18681,N_7855,N_11487);
nand U18682 (N_18682,N_7061,N_12324);
and U18683 (N_18683,N_11806,N_11842);
or U18684 (N_18684,N_6860,N_10220);
nand U18685 (N_18685,N_8004,N_11147);
and U18686 (N_18686,N_8780,N_11439);
or U18687 (N_18687,N_6623,N_8871);
and U18688 (N_18688,N_10739,N_10512);
nor U18689 (N_18689,N_9802,N_8214);
nor U18690 (N_18690,N_8376,N_7228);
nand U18691 (N_18691,N_7921,N_7785);
and U18692 (N_18692,N_7039,N_10965);
nand U18693 (N_18693,N_7026,N_11271);
xor U18694 (N_18694,N_8555,N_10621);
nand U18695 (N_18695,N_7590,N_7629);
and U18696 (N_18696,N_7095,N_6744);
nor U18697 (N_18697,N_10119,N_8715);
or U18698 (N_18698,N_11623,N_10443);
nand U18699 (N_18699,N_9666,N_11636);
nor U18700 (N_18700,N_6361,N_12305);
or U18701 (N_18701,N_10451,N_9351);
nor U18702 (N_18702,N_11489,N_9039);
nand U18703 (N_18703,N_10397,N_6533);
and U18704 (N_18704,N_8698,N_11254);
nor U18705 (N_18705,N_10330,N_7604);
or U18706 (N_18706,N_10557,N_10186);
and U18707 (N_18707,N_9146,N_9873);
nand U18708 (N_18708,N_10828,N_11791);
nand U18709 (N_18709,N_7571,N_11888);
nor U18710 (N_18710,N_6686,N_7029);
or U18711 (N_18711,N_12207,N_11075);
and U18712 (N_18712,N_10521,N_7838);
nand U18713 (N_18713,N_11509,N_6371);
or U18714 (N_18714,N_10546,N_10439);
or U18715 (N_18715,N_10173,N_6529);
and U18716 (N_18716,N_12306,N_12149);
or U18717 (N_18717,N_12457,N_9260);
and U18718 (N_18718,N_11280,N_6837);
nor U18719 (N_18719,N_10374,N_8298);
nor U18720 (N_18720,N_9031,N_12189);
nor U18721 (N_18721,N_7712,N_12442);
nor U18722 (N_18722,N_9619,N_11247);
or U18723 (N_18723,N_8535,N_9152);
and U18724 (N_18724,N_6421,N_9100);
or U18725 (N_18725,N_10882,N_8579);
nor U18726 (N_18726,N_6606,N_8623);
nand U18727 (N_18727,N_8063,N_12403);
or U18728 (N_18728,N_11788,N_8638);
nand U18729 (N_18729,N_7178,N_11723);
and U18730 (N_18730,N_9131,N_6427);
or U18731 (N_18731,N_6348,N_12040);
or U18732 (N_18732,N_11209,N_11838);
nor U18733 (N_18733,N_12009,N_8075);
and U18734 (N_18734,N_11024,N_10430);
nand U18735 (N_18735,N_7307,N_8163);
nor U18736 (N_18736,N_8422,N_9236);
or U18737 (N_18737,N_8062,N_11956);
or U18738 (N_18738,N_8123,N_10506);
nor U18739 (N_18739,N_10227,N_7550);
and U18740 (N_18740,N_7908,N_10392);
nor U18741 (N_18741,N_11162,N_11858);
or U18742 (N_18742,N_12161,N_10038);
or U18743 (N_18743,N_9090,N_12200);
nand U18744 (N_18744,N_6668,N_7576);
and U18745 (N_18745,N_8134,N_7068);
or U18746 (N_18746,N_10184,N_8174);
nand U18747 (N_18747,N_10736,N_9489);
nor U18748 (N_18748,N_12492,N_11782);
nand U18749 (N_18749,N_9902,N_9408);
nor U18750 (N_18750,N_14066,N_13363);
nor U18751 (N_18751,N_14097,N_13564);
nor U18752 (N_18752,N_18509,N_13780);
nor U18753 (N_18753,N_13736,N_14899);
and U18754 (N_18754,N_18383,N_13813);
nand U18755 (N_18755,N_12530,N_16687);
nand U18756 (N_18756,N_18610,N_18555);
or U18757 (N_18757,N_17894,N_12686);
nor U18758 (N_18758,N_12715,N_14669);
or U18759 (N_18759,N_17153,N_13580);
or U18760 (N_18760,N_17168,N_14302);
nor U18761 (N_18761,N_13196,N_12734);
and U18762 (N_18762,N_15746,N_13300);
or U18763 (N_18763,N_18408,N_17193);
and U18764 (N_18764,N_17981,N_15939);
nor U18765 (N_18765,N_14436,N_15732);
nand U18766 (N_18766,N_17347,N_18121);
nor U18767 (N_18767,N_16221,N_15264);
and U18768 (N_18768,N_17989,N_18184);
and U18769 (N_18769,N_14390,N_14083);
and U18770 (N_18770,N_15821,N_18377);
and U18771 (N_18771,N_16938,N_16219);
and U18772 (N_18772,N_17539,N_15598);
or U18773 (N_18773,N_13815,N_15488);
or U18774 (N_18774,N_12835,N_14008);
nand U18775 (N_18775,N_17964,N_18692);
nand U18776 (N_18776,N_18251,N_18000);
nor U18777 (N_18777,N_15270,N_13814);
and U18778 (N_18778,N_14359,N_18313);
nand U18779 (N_18779,N_18083,N_15786);
or U18780 (N_18780,N_16532,N_18059);
nand U18781 (N_18781,N_17351,N_17979);
xnor U18782 (N_18782,N_16502,N_17505);
nand U18783 (N_18783,N_16740,N_14857);
nor U18784 (N_18784,N_12839,N_14307);
or U18785 (N_18785,N_13180,N_18673);
nor U18786 (N_18786,N_17320,N_16737);
nand U18787 (N_18787,N_14033,N_13922);
and U18788 (N_18788,N_15183,N_12905);
or U18789 (N_18789,N_13956,N_18286);
nor U18790 (N_18790,N_18245,N_13174);
nand U18791 (N_18791,N_17341,N_16739);
and U18792 (N_18792,N_14349,N_17866);
and U18793 (N_18793,N_15458,N_17840);
nand U18794 (N_18794,N_12860,N_15966);
or U18795 (N_18795,N_13468,N_14306);
and U18796 (N_18796,N_13404,N_14563);
or U18797 (N_18797,N_14023,N_14181);
and U18798 (N_18798,N_17234,N_14754);
nand U18799 (N_18799,N_14274,N_18566);
and U18800 (N_18800,N_13089,N_15872);
and U18801 (N_18801,N_17358,N_14922);
or U18802 (N_18802,N_14262,N_17547);
nor U18803 (N_18803,N_14670,N_13154);
or U18804 (N_18804,N_15906,N_16040);
nand U18805 (N_18805,N_15856,N_14575);
and U18806 (N_18806,N_16696,N_16885);
or U18807 (N_18807,N_14744,N_16478);
nand U18808 (N_18808,N_17674,N_14743);
nor U18809 (N_18809,N_16634,N_15589);
nor U18810 (N_18810,N_15835,N_16330);
or U18811 (N_18811,N_13985,N_17160);
nand U18812 (N_18812,N_17939,N_18367);
and U18813 (N_18813,N_18553,N_15690);
nor U18814 (N_18814,N_13103,N_14682);
or U18815 (N_18815,N_15641,N_12829);
or U18816 (N_18816,N_18291,N_16184);
and U18817 (N_18817,N_15235,N_15283);
and U18818 (N_18818,N_18015,N_17764);
nor U18819 (N_18819,N_15627,N_12675);
nor U18820 (N_18820,N_15797,N_13545);
or U18821 (N_18821,N_16389,N_15278);
or U18822 (N_18822,N_13137,N_18329);
nor U18823 (N_18823,N_16760,N_17060);
or U18824 (N_18824,N_17633,N_15206);
nor U18825 (N_18825,N_16793,N_15505);
nor U18826 (N_18826,N_13717,N_15764);
nor U18827 (N_18827,N_15637,N_18572);
or U18828 (N_18828,N_13573,N_18434);
nor U18829 (N_18829,N_13806,N_17728);
nor U18830 (N_18830,N_13658,N_15405);
nor U18831 (N_18831,N_12730,N_12856);
nor U18832 (N_18832,N_14467,N_13537);
and U18833 (N_18833,N_14363,N_12576);
or U18834 (N_18834,N_17555,N_17739);
nand U18835 (N_18835,N_13969,N_15360);
nand U18836 (N_18836,N_17807,N_12944);
nor U18837 (N_18837,N_17285,N_14965);
or U18838 (N_18838,N_12643,N_13816);
and U18839 (N_18839,N_18139,N_14718);
and U18840 (N_18840,N_14497,N_15429);
nor U18841 (N_18841,N_14408,N_16937);
nor U18842 (N_18842,N_16287,N_17540);
or U18843 (N_18843,N_15704,N_15813);
nand U18844 (N_18844,N_17877,N_14045);
nand U18845 (N_18845,N_12722,N_15408);
and U18846 (N_18846,N_15179,N_15995);
nand U18847 (N_18847,N_13737,N_14056);
nand U18848 (N_18848,N_17130,N_14425);
and U18849 (N_18849,N_14297,N_15684);
or U18850 (N_18850,N_12701,N_12747);
and U18851 (N_18851,N_17299,N_16597);
and U18852 (N_18852,N_15734,N_17693);
and U18853 (N_18853,N_13826,N_15387);
or U18854 (N_18854,N_13407,N_17819);
nand U18855 (N_18855,N_15897,N_13710);
and U18856 (N_18856,N_17617,N_15852);
and U18857 (N_18857,N_18220,N_15290);
and U18858 (N_18858,N_15067,N_17650);
and U18859 (N_18859,N_13641,N_16365);
xor U18860 (N_18860,N_16875,N_14044);
and U18861 (N_18861,N_13220,N_16032);
nand U18862 (N_18862,N_18538,N_18520);
or U18863 (N_18863,N_16583,N_14533);
nor U18864 (N_18864,N_14423,N_12574);
nand U18865 (N_18865,N_14879,N_18160);
or U18866 (N_18866,N_16311,N_18525);
nor U18867 (N_18867,N_18544,N_12610);
nand U18868 (N_18868,N_15147,N_18400);
and U18869 (N_18869,N_17105,N_17369);
nor U18870 (N_18870,N_13097,N_17996);
or U18871 (N_18871,N_17647,N_14574);
nor U18872 (N_18872,N_17533,N_18308);
or U18873 (N_18873,N_16526,N_14554);
nor U18874 (N_18874,N_14263,N_14671);
or U18875 (N_18875,N_15004,N_16637);
or U18876 (N_18876,N_12975,N_13524);
nor U18877 (N_18877,N_13324,N_14404);
or U18878 (N_18878,N_18310,N_17361);
nand U18879 (N_18879,N_15203,N_13712);
and U18880 (N_18880,N_14600,N_12503);
nor U18881 (N_18881,N_17554,N_15048);
or U18882 (N_18882,N_13534,N_16312);
nand U18883 (N_18883,N_17587,N_14878);
or U18884 (N_18884,N_12685,N_14143);
nor U18885 (N_18885,N_18445,N_17391);
nand U18886 (N_18886,N_14199,N_14295);
nor U18887 (N_18887,N_18606,N_16440);
nor U18888 (N_18888,N_15355,N_16870);
or U18889 (N_18889,N_13749,N_16578);
or U18890 (N_18890,N_18479,N_14915);
nand U18891 (N_18891,N_16404,N_12621);
or U18892 (N_18892,N_16611,N_13606);
nor U18893 (N_18893,N_18195,N_14875);
or U18894 (N_18894,N_12876,N_14060);
nand U18895 (N_18895,N_14004,N_13971);
and U18896 (N_18896,N_17576,N_16987);
and U18897 (N_18897,N_14544,N_12815);
nand U18898 (N_18898,N_13551,N_13568);
nor U18899 (N_18899,N_15624,N_17604);
and U18900 (N_18900,N_14132,N_17519);
nand U18901 (N_18901,N_14805,N_13833);
and U18902 (N_18902,N_17305,N_18249);
nor U18903 (N_18903,N_13898,N_15857);
nand U18904 (N_18904,N_15537,N_14643);
and U18905 (N_18905,N_13998,N_13374);
nand U18906 (N_18906,N_16301,N_12716);
xor U18907 (N_18907,N_13062,N_18266);
or U18908 (N_18908,N_18001,N_18393);
nor U18909 (N_18909,N_13491,N_14590);
and U18910 (N_18910,N_17883,N_17805);
and U18911 (N_18911,N_15791,N_16631);
nand U18912 (N_18912,N_13155,N_18109);
or U18913 (N_18913,N_16707,N_15366);
or U18914 (N_18914,N_18593,N_16347);
and U18915 (N_18915,N_14852,N_18186);
and U18916 (N_18916,N_16999,N_17700);
and U18917 (N_18917,N_16897,N_15053);
and U18918 (N_18918,N_12859,N_15007);
nor U18919 (N_18919,N_16280,N_15105);
nand U18920 (N_18920,N_13275,N_17499);
or U18921 (N_18921,N_13613,N_16797);
xnor U18922 (N_18922,N_17366,N_15879);
and U18923 (N_18923,N_16399,N_12587);
and U18924 (N_18924,N_14821,N_14789);
nor U18925 (N_18925,N_15097,N_15487);
nand U18926 (N_18926,N_16249,N_14940);
nor U18927 (N_18927,N_16736,N_17681);
or U18928 (N_18928,N_13330,N_13336);
and U18929 (N_18929,N_14516,N_15417);
and U18930 (N_18930,N_13988,N_14429);
nor U18931 (N_18931,N_18158,N_16203);
nor U18932 (N_18932,N_15755,N_13775);
nor U18933 (N_18933,N_18685,N_17476);
nor U18934 (N_18934,N_12752,N_17084);
nand U18935 (N_18935,N_15463,N_16603);
and U18936 (N_18936,N_15483,N_14779);
and U18937 (N_18937,N_18017,N_15626);
xor U18938 (N_18938,N_12708,N_15436);
or U18939 (N_18939,N_14187,N_18091);
nor U18940 (N_18940,N_13065,N_16428);
and U18941 (N_18941,N_12939,N_16930);
or U18942 (N_18942,N_16756,N_17003);
nor U18943 (N_18943,N_14774,N_18484);
or U18944 (N_18944,N_17182,N_14732);
xor U18945 (N_18945,N_17240,N_18315);
or U18946 (N_18946,N_17441,N_13785);
nand U18947 (N_18947,N_17659,N_14361);
nor U18948 (N_18948,N_14142,N_15378);
nor U18949 (N_18949,N_13555,N_18737);
nor U18950 (N_18950,N_14714,N_13250);
nor U18951 (N_18951,N_13596,N_14511);
or U18952 (N_18952,N_13740,N_16016);
and U18953 (N_18953,N_17909,N_14335);
nor U18954 (N_18954,N_17304,N_16935);
and U18955 (N_18955,N_17280,N_18153);
nand U18956 (N_18956,N_14287,N_17638);
nand U18957 (N_18957,N_18543,N_18114);
nand U18958 (N_18958,N_17745,N_13305);
or U18959 (N_18959,N_18702,N_17814);
nand U18960 (N_18960,N_13413,N_18202);
or U18961 (N_18961,N_15272,N_14583);
and U18962 (N_18962,N_17772,N_16346);
and U18963 (N_18963,N_17402,N_16601);
nor U18964 (N_18964,N_12510,N_18200);
nand U18965 (N_18965,N_12799,N_12899);
nand U18966 (N_18966,N_18292,N_15014);
nand U18967 (N_18967,N_14947,N_17312);
nor U18968 (N_18968,N_15792,N_17662);
nand U18969 (N_18969,N_16796,N_13756);
or U18970 (N_18970,N_17691,N_15774);
nor U18971 (N_18971,N_16645,N_17356);
nand U18972 (N_18972,N_12853,N_13367);
or U18973 (N_18973,N_14186,N_14726);
or U18974 (N_18974,N_16952,N_13027);
nor U18975 (N_18975,N_13990,N_14339);
nand U18976 (N_18976,N_18345,N_15807);
or U18977 (N_18977,N_14636,N_12571);
and U18978 (N_18978,N_15107,N_13805);
or U18979 (N_18979,N_16821,N_18029);
or U18980 (N_18980,N_12569,N_14084);
or U18981 (N_18981,N_14498,N_17790);
nor U18982 (N_18982,N_15396,N_13008);
or U18983 (N_18983,N_18020,N_15834);
nand U18984 (N_18984,N_17118,N_13049);
or U18985 (N_18985,N_18055,N_13381);
nor U18986 (N_18986,N_16263,N_18006);
and U18987 (N_18987,N_13777,N_15259);
or U18988 (N_18988,N_13124,N_14639);
or U18989 (N_18989,N_14820,N_18070);
nor U18990 (N_18990,N_17574,N_14730);
or U18991 (N_18991,N_18682,N_17594);
and U18992 (N_18992,N_16860,N_18574);
nor U18993 (N_18993,N_17159,N_12872);
nor U18994 (N_18994,N_18027,N_15265);
and U18995 (N_18995,N_14047,N_14546);
and U18996 (N_18996,N_13256,N_16564);
and U18997 (N_18997,N_17085,N_17117);
nor U18998 (N_18998,N_15023,N_18644);
nand U18999 (N_18999,N_17449,N_17238);
or U19000 (N_19000,N_17844,N_15016);
nand U19001 (N_19001,N_17020,N_14281);
nand U19002 (N_19002,N_17876,N_13999);
and U19003 (N_19003,N_17599,N_17173);
and U19004 (N_19004,N_13763,N_16027);
and U19005 (N_19005,N_17773,N_13301);
and U19006 (N_19006,N_13630,N_13132);
nor U19007 (N_19007,N_13398,N_17392);
or U19008 (N_19008,N_15291,N_15351);
or U19009 (N_19009,N_13681,N_16717);
nand U19010 (N_19010,N_13197,N_16521);
and U19011 (N_19011,N_13422,N_17925);
or U19012 (N_19012,N_17446,N_18639);
nor U19013 (N_19013,N_18468,N_18043);
nand U19014 (N_19014,N_12992,N_13688);
or U19015 (N_19015,N_14489,N_17463);
nand U19016 (N_19016,N_16486,N_18085);
or U19017 (N_19017,N_15033,N_16361);
or U19018 (N_19018,N_14793,N_16618);
and U19019 (N_19019,N_14316,N_12877);
nor U19020 (N_19020,N_16001,N_14322);
xnor U19021 (N_19021,N_17690,N_12970);
nor U19022 (N_19022,N_15092,N_17958);
and U19023 (N_19023,N_13632,N_16491);
or U19024 (N_19024,N_15032,N_13703);
and U19025 (N_19025,N_18728,N_16528);
nand U19026 (N_19026,N_16841,N_14381);
nand U19027 (N_19027,N_15006,N_16956);
xnor U19028 (N_19028,N_13726,N_17873);
nor U19029 (N_19029,N_17157,N_14421);
nand U19030 (N_19030,N_14571,N_14104);
nand U19031 (N_19031,N_16196,N_17218);
or U19032 (N_19032,N_18011,N_17059);
or U19033 (N_19033,N_17683,N_14487);
and U19034 (N_19034,N_17052,N_12502);
nor U19035 (N_19035,N_18429,N_18233);
and U19036 (N_19036,N_14666,N_18670);
or U19037 (N_19037,N_18415,N_12583);
and U19038 (N_19038,N_14503,N_17453);
nand U19039 (N_19039,N_17217,N_18129);
nor U19040 (N_19040,N_13742,N_12573);
and U19041 (N_19041,N_17077,N_16066);
or U19042 (N_19042,N_17957,N_14891);
nand U19043 (N_19043,N_12867,N_13648);
or U19044 (N_19044,N_14581,N_15026);
nand U19045 (N_19045,N_16883,N_14450);
nor U19046 (N_19046,N_17777,N_14254);
or U19047 (N_19047,N_13809,N_12606);
nor U19048 (N_19048,N_14502,N_15655);
and U19049 (N_19049,N_18330,N_12971);
nand U19050 (N_19050,N_12828,N_13018);
nand U19051 (N_19051,N_14887,N_17559);
or U19052 (N_19052,N_16051,N_14317);
nor U19053 (N_19053,N_18744,N_18361);
and U19054 (N_19054,N_17542,N_14723);
and U19055 (N_19055,N_16406,N_16520);
nor U19056 (N_19056,N_13760,N_15126);
nor U19057 (N_19057,N_17897,N_17144);
nand U19058 (N_19058,N_17213,N_14746);
nand U19059 (N_19059,N_16238,N_13267);
or U19060 (N_19060,N_13676,N_15754);
nor U19061 (N_19061,N_13393,N_17868);
and U19062 (N_19062,N_13045,N_15043);
xnor U19063 (N_19063,N_17705,N_12847);
nor U19064 (N_19064,N_12816,N_18643);
or U19065 (N_19065,N_16501,N_18013);
nand U19066 (N_19066,N_17724,N_17704);
or U19067 (N_19067,N_17001,N_16672);
nor U19068 (N_19068,N_18050,N_17028);
nor U19069 (N_19069,N_17349,N_16150);
or U19070 (N_19070,N_16158,N_14838);
xnor U19071 (N_19071,N_15199,N_15213);
nor U19072 (N_19072,N_15996,N_14768);
and U19073 (N_19073,N_18080,N_16147);
and U19074 (N_19074,N_18503,N_17265);
or U19075 (N_19075,N_18311,N_18549);
nor U19076 (N_19076,N_18470,N_16338);
nor U19077 (N_19077,N_12743,N_16002);
or U19078 (N_19078,N_16480,N_15343);
nor U19079 (N_19079,N_16137,N_16206);
or U19080 (N_19080,N_17846,N_16622);
or U19081 (N_19081,N_14163,N_14631);
or U19082 (N_19082,N_13497,N_17222);
nand U19083 (N_19083,N_17904,N_15570);
nand U19084 (N_19084,N_15441,N_17603);
nor U19085 (N_19085,N_14379,N_18036);
or U19086 (N_19086,N_15500,N_15325);
nand U19087 (N_19087,N_18480,N_15143);
and U19088 (N_19088,N_15938,N_14606);
nand U19089 (N_19089,N_13773,N_17270);
nor U19090 (N_19090,N_13327,N_15494);
nor U19091 (N_19091,N_16344,N_13872);
nor U19092 (N_19092,N_16554,N_18684);
and U19093 (N_19093,N_14983,N_14996);
and U19094 (N_19094,N_14245,N_18556);
or U19095 (N_19095,N_18634,N_16418);
or U19096 (N_19096,N_14742,N_18414);
or U19097 (N_19097,N_16214,N_13184);
nand U19098 (N_19098,N_13920,N_16921);
nand U19099 (N_19099,N_14035,N_12881);
nor U19100 (N_19100,N_13601,N_14909);
and U19101 (N_19101,N_16457,N_17889);
nand U19102 (N_19102,N_16102,N_14847);
nor U19103 (N_19103,N_15468,N_14266);
or U19104 (N_19104,N_14180,N_15548);
or U19105 (N_19105,N_15082,N_14395);
nor U19106 (N_19106,N_17988,N_15731);
nor U19107 (N_19107,N_15660,N_13923);
xor U19108 (N_19108,N_13099,N_13216);
nand U19109 (N_19109,N_14889,N_13080);
and U19110 (N_19110,N_17634,N_17692);
and U19111 (N_19111,N_13368,N_18689);
nand U19112 (N_19112,N_17324,N_13347);
and U19113 (N_19113,N_13280,N_14505);
nand U19114 (N_19114,N_13957,N_16430);
and U19115 (N_19115,N_17590,N_15733);
and U19116 (N_19116,N_17608,N_18740);
and U19117 (N_19117,N_16615,N_14913);
and U19118 (N_19118,N_18280,N_14595);
and U19119 (N_19119,N_17335,N_18583);
nor U19120 (N_19120,N_12626,N_17830);
and U19121 (N_19121,N_16610,N_14464);
nor U19122 (N_19122,N_17671,N_14515);
and U19123 (N_19123,N_15973,N_12957);
and U19124 (N_19124,N_16007,N_18726);
and U19125 (N_19125,N_13035,N_16630);
or U19126 (N_19126,N_14698,N_16979);
nand U19127 (N_19127,N_14610,N_15565);
or U19128 (N_19128,N_18481,N_14905);
and U19129 (N_19129,N_15956,N_15763);
and U19130 (N_19130,N_16977,N_14230);
and U19131 (N_19131,N_17415,N_16161);
nand U19132 (N_19132,N_18743,N_18223);
xor U19133 (N_19133,N_13536,N_15703);
nor U19134 (N_19134,N_16705,N_18483);
and U19135 (N_19135,N_17562,N_14396);
nor U19136 (N_19136,N_14668,N_15578);
nand U19137 (N_19137,N_13786,N_16036);
or U19138 (N_19138,N_13528,N_14435);
nor U19139 (N_19139,N_14347,N_14030);
nor U19140 (N_19140,N_16257,N_15386);
nor U19141 (N_19141,N_17624,N_16391);
or U19142 (N_19142,N_17276,N_12884);
nor U19143 (N_19143,N_18508,N_16211);
nor U19144 (N_19144,N_13748,N_15568);
or U19145 (N_19145,N_15263,N_18487);
nor U19146 (N_19146,N_16386,N_12919);
or U19147 (N_19147,N_14759,N_17763);
or U19148 (N_19148,N_15022,N_18355);
nor U19149 (N_19149,N_14693,N_12733);
nor U19150 (N_19150,N_12711,N_14329);
nor U19151 (N_19151,N_13510,N_15839);
or U19152 (N_19152,N_12796,N_12914);
or U19153 (N_19153,N_14334,N_17256);
or U19154 (N_19154,N_15768,N_16733);
and U19155 (N_19155,N_17307,N_15708);
and U19156 (N_19156,N_12917,N_16209);
and U19157 (N_19157,N_13211,N_12967);
nor U19158 (N_19158,N_17570,N_16019);
nor U19159 (N_19159,N_16185,N_16684);
nor U19160 (N_19160,N_13364,N_12618);
or U19161 (N_19161,N_17960,N_14021);
and U19162 (N_19162,N_15375,N_13447);
nor U19163 (N_19163,N_14969,N_16484);
and U19164 (N_19164,N_13457,N_13512);
nand U19165 (N_19165,N_18265,N_18530);
nand U19166 (N_19166,N_14434,N_17629);
and U19167 (N_19167,N_16111,N_12608);
nand U19168 (N_19168,N_16006,N_15659);
or U19169 (N_19169,N_14757,N_16332);
and U19170 (N_19170,N_16172,N_16500);
and U19171 (N_19171,N_17104,N_12582);
or U19172 (N_19172,N_13732,N_14330);
and U19173 (N_19173,N_16121,N_15280);
nor U19174 (N_19174,N_15510,N_13012);
nor U19175 (N_19175,N_13500,N_13001);
nor U19176 (N_19176,N_18394,N_13126);
and U19177 (N_19177,N_12516,N_15148);
and U19178 (N_19178,N_17615,N_17491);
and U19179 (N_19179,N_16131,N_15306);
nand U19180 (N_19180,N_15108,N_12789);
nor U19181 (N_19181,N_17040,N_12861);
nand U19182 (N_19182,N_16152,N_14304);
nand U19183 (N_19183,N_16068,N_13662);
or U19184 (N_19184,N_17195,N_18648);
nand U19185 (N_19185,N_15224,N_16809);
or U19186 (N_19186,N_16425,N_15432);
nor U19187 (N_19187,N_13506,N_18038);
nand U19188 (N_19188,N_18626,N_14537);
nand U19189 (N_19189,N_13005,N_16671);
nand U19190 (N_19190,N_15083,N_16288);
and U19191 (N_19191,N_15124,N_13711);
nor U19192 (N_19192,N_14433,N_15762);
nor U19193 (N_19193,N_15055,N_16779);
nor U19194 (N_19194,N_16792,N_12520);
and U19195 (N_19195,N_18459,N_18053);
and U19196 (N_19196,N_13191,N_14265);
nand U19197 (N_19197,N_17373,N_18357);
and U19198 (N_19198,N_17906,N_17716);
and U19199 (N_19199,N_12792,N_14228);
or U19200 (N_19200,N_13276,N_16980);
or U19201 (N_19201,N_16397,N_14767);
nor U19202 (N_19202,N_13303,N_15584);
or U19203 (N_19203,N_15489,N_13770);
nor U19204 (N_19204,N_14208,N_13808);
or U19205 (N_19205,N_13122,N_13618);
or U19206 (N_19206,N_16023,N_17431);
nor U19207 (N_19207,N_14658,N_17506);
or U19208 (N_19208,N_15931,N_14242);
nor U19209 (N_19209,N_16826,N_17826);
nand U19210 (N_19210,N_17246,N_13169);
or U19211 (N_19211,N_17058,N_17186);
or U19212 (N_19212,N_13257,N_18102);
or U19213 (N_19213,N_16237,N_17272);
or U19214 (N_19214,N_17689,N_15649);
nor U19215 (N_19215,N_13961,N_15036);
and U19216 (N_19216,N_12945,N_15312);
nand U19217 (N_19217,N_14618,N_18067);
and U19218 (N_19218,N_18034,N_14234);
nand U19219 (N_19219,N_16799,N_15593);
nor U19220 (N_19220,N_17991,N_14482);
and U19221 (N_19221,N_14911,N_14432);
nand U19222 (N_19222,N_16376,N_14865);
and U19223 (N_19223,N_18569,N_14129);
or U19224 (N_19224,N_15622,N_17541);
nand U19225 (N_19225,N_15061,N_16827);
and U19226 (N_19226,N_18523,N_17239);
and U19227 (N_19227,N_18524,N_18476);
and U19228 (N_19228,N_13698,N_16207);
nor U19229 (N_19229,N_13247,N_17072);
nand U19230 (N_19230,N_15020,N_14437);
and U19231 (N_19231,N_16644,N_16182);
and U19232 (N_19232,N_12960,N_14810);
nor U19233 (N_19233,N_17236,N_14098);
or U19234 (N_19234,N_13819,N_15576);
xnor U19235 (N_19235,N_16354,N_18533);
nand U19236 (N_19236,N_16924,N_17284);
and U19237 (N_19237,N_16616,N_13863);
and U19238 (N_19238,N_14534,N_12611);
nand U19239 (N_19239,N_13302,N_16636);
or U19240 (N_19240,N_17433,N_13899);
nand U19241 (N_19241,N_16818,N_15529);
or U19242 (N_19242,N_14738,N_14828);
and U19243 (N_19243,N_17189,N_12525);
xnor U19244 (N_19244,N_12763,N_17743);
nor U19245 (N_19245,N_14599,N_15042);
nand U19246 (N_19246,N_16983,N_13262);
or U19247 (N_19247,N_17303,N_17413);
nor U19248 (N_19248,N_18430,N_16334);
or U19249 (N_19249,N_17708,N_13337);
nand U19250 (N_19250,N_14917,N_17825);
nand U19251 (N_19251,N_13289,N_15884);
nor U19252 (N_19252,N_16157,N_15089);
xor U19253 (N_19253,N_16804,N_12717);
nor U19254 (N_19254,N_16427,N_13362);
and U19255 (N_19255,N_16268,N_13040);
xnor U19256 (N_19256,N_15910,N_15688);
nand U19257 (N_19257,N_18211,N_16026);
and U19258 (N_19258,N_15794,N_14291);
or U19259 (N_19259,N_15916,N_17838);
nor U19260 (N_19260,N_16115,N_16299);
nand U19261 (N_19261,N_16762,N_13160);
and U19262 (N_19262,N_16042,N_12756);
and U19263 (N_19263,N_15181,N_16505);
nor U19264 (N_19264,N_14413,N_17009);
and U19265 (N_19265,N_16227,N_17436);
nor U19266 (N_19266,N_13572,N_16949);
nor U19267 (N_19267,N_15120,N_18285);
and U19268 (N_19268,N_13840,N_17025);
nand U19269 (N_19269,N_16982,N_15738);
nand U19270 (N_19270,N_14679,N_14125);
and U19271 (N_19271,N_12667,N_15069);
and U19272 (N_19272,N_16713,N_16327);
nor U19273 (N_19273,N_16906,N_16384);
xor U19274 (N_19274,N_14382,N_14586);
or U19275 (N_19275,N_17480,N_17139);
nand U19276 (N_19276,N_15327,N_15767);
nand U19277 (N_19277,N_12737,N_13881);
and U19278 (N_19278,N_16517,N_17994);
nand U19279 (N_19279,N_15072,N_14428);
or U19280 (N_19280,N_16188,N_16642);
nand U19281 (N_19281,N_18446,N_17385);
or U19282 (N_19282,N_16744,N_13539);
or U19283 (N_19283,N_12553,N_15694);
nand U19284 (N_19284,N_17401,N_12915);
or U19285 (N_19285,N_15698,N_14276);
nor U19286 (N_19286,N_13950,N_17818);
nor U19287 (N_19287,N_15997,N_16351);
nor U19288 (N_19288,N_15434,N_15223);
nand U19289 (N_19289,N_12691,N_17126);
and U19290 (N_19290,N_13679,N_17933);
nor U19291 (N_19291,N_16881,N_18193);
or U19292 (N_19292,N_14018,N_17682);
nor U19293 (N_19293,N_15379,N_14736);
nor U19294 (N_19294,N_17282,N_14806);
nand U19295 (N_19295,N_16395,N_17170);
and U19296 (N_19296,N_14861,N_14691);
nand U19297 (N_19297,N_13862,N_18352);
or U19298 (N_19298,N_17423,N_14565);
nor U19299 (N_19299,N_13494,N_17398);
or U19300 (N_19300,N_17998,N_17835);
nand U19301 (N_19301,N_15854,N_14486);
nor U19302 (N_19302,N_13997,N_15971);
or U19303 (N_19303,N_18664,N_15985);
and U19304 (N_19304,N_18507,N_16604);
nand U19305 (N_19305,N_15262,N_18284);
or U19306 (N_19306,N_15365,N_14734);
nand U19307 (N_19307,N_15535,N_12993);
and U19308 (N_19308,N_12668,N_14271);
nor U19309 (N_19309,N_12921,N_16048);
nor U19310 (N_19310,N_16393,N_18264);
and U19311 (N_19311,N_13970,N_16621);
and U19312 (N_19312,N_16558,N_15934);
and U19313 (N_19313,N_16193,N_13032);
nor U19314 (N_19314,N_16902,N_16010);
or U19315 (N_19315,N_12515,N_13294);
xnor U19316 (N_19316,N_15513,N_15796);
nand U19317 (N_19317,N_12837,N_18004);
or U19318 (N_19318,N_13514,N_12559);
or U19319 (N_19319,N_16800,N_15743);
nand U19320 (N_19320,N_12911,N_15476);
and U19321 (N_19321,N_15296,N_16362);
or U19322 (N_19322,N_12927,N_13416);
or U19323 (N_19323,N_15328,N_15948);
and U19324 (N_19324,N_16101,N_18505);
nand U19325 (N_19325,N_13574,N_17949);
nand U19326 (N_19326,N_16751,N_18542);
nor U19327 (N_19327,N_16489,N_15000);
nand U19328 (N_19328,N_15845,N_15070);
nand U19329 (N_19329,N_17512,N_17592);
nand U19330 (N_19330,N_13513,N_15984);
nor U19331 (N_19331,N_17093,N_13285);
or U19332 (N_19332,N_16820,N_13832);
and U19333 (N_19333,N_18427,N_15758);
or U19334 (N_19334,N_15722,N_14243);
or U19335 (N_19335,N_13480,N_17810);
nand U19336 (N_19336,N_14531,N_18498);
nand U19337 (N_19337,N_14484,N_14357);
nor U19338 (N_19338,N_14403,N_13475);
nand U19339 (N_19339,N_13473,N_13215);
and U19340 (N_19340,N_16967,N_12521);
nand U19341 (N_19341,N_12956,N_17326);
nor U19342 (N_19342,N_16005,N_13781);
nor U19343 (N_19343,N_15433,N_12898);
nor U19344 (N_19344,N_18100,N_13823);
and U19345 (N_19345,N_14870,N_16625);
and U19346 (N_19346,N_12783,N_18680);
and U19347 (N_19347,N_13292,N_16819);
or U19348 (N_19348,N_17231,N_17678);
and U19349 (N_19349,N_17253,N_17161);
nor U19350 (N_19350,N_17612,N_15936);
xor U19351 (N_19351,N_15766,N_15986);
or U19352 (N_19352,N_15718,N_13868);
nor U19353 (N_19353,N_17178,N_13745);
and U19354 (N_19354,N_16774,N_14513);
and U19355 (N_19355,N_16547,N_18155);
nand U19356 (N_19356,N_16396,N_17696);
or U19357 (N_19357,N_17523,N_13236);
and U19358 (N_19358,N_13629,N_12538);
nand U19359 (N_19359,N_16195,N_17621);
or U19360 (N_19360,N_14777,N_15341);
nor U19361 (N_19361,N_17527,N_18044);
or U19362 (N_19362,N_13900,N_16348);
nand U19363 (N_19363,N_17224,N_14337);
and U19364 (N_19364,N_18250,N_13892);
and U19365 (N_19365,N_15546,N_18418);
xor U19366 (N_19366,N_17333,N_15150);
and U19367 (N_19367,N_15154,N_17442);
nand U19368 (N_19368,N_12999,N_14448);
and U19369 (N_19369,N_15301,N_16627);
nor U19370 (N_19370,N_18686,N_12846);
nand U19371 (N_19371,N_14924,N_13668);
nor U19372 (N_19372,N_16889,N_12836);
nor U19373 (N_19373,N_17416,N_16531);
and U19374 (N_19374,N_17279,N_17399);
or U19375 (N_19375,N_13522,N_18189);
and U19376 (N_19376,N_16091,N_15748);
nand U19377 (N_19377,N_14722,N_14703);
nor U19378 (N_19378,N_15846,N_17639);
and U19379 (N_19379,N_15621,N_13691);
or U19380 (N_19380,N_16283,N_16488);
nand U19381 (N_19381,N_18318,N_17345);
or U19382 (N_19382,N_13263,N_14880);
nor U19383 (N_19383,N_16224,N_18552);
nor U19384 (N_19384,N_13231,N_15282);
or U19385 (N_19385,N_17427,N_17495);
nor U19386 (N_19386,N_13401,N_14923);
nand U19387 (N_19387,N_15196,N_16493);
nand U19388 (N_19388,N_14567,N_13746);
and U19389 (N_19389,N_12712,N_13427);
and U19390 (N_19390,N_13210,N_15582);
or U19391 (N_19391,N_14350,N_13237);
or U19392 (N_19392,N_17622,N_15404);
or U19393 (N_19393,N_14570,N_18110);
nor U19394 (N_19394,N_15059,N_14000);
and U19395 (N_19395,N_15521,N_17046);
or U19396 (N_19396,N_15220,N_17912);
nand U19397 (N_19397,N_16436,N_12969);
and U19398 (N_19398,N_16693,N_17517);
or U19399 (N_19399,N_18609,N_15112);
and U19400 (N_19400,N_16919,N_15744);
nand U19401 (N_19401,N_17852,N_15060);
and U19402 (N_19402,N_16252,N_15972);
or U19403 (N_19403,N_12695,N_13382);
nand U19404 (N_19404,N_14442,N_15099);
and U19405 (N_19405,N_15957,N_17411);
and U19406 (N_19406,N_17987,N_18494);
and U19407 (N_19407,N_14106,N_12632);
and U19408 (N_19408,N_18496,N_13450);
nand U19409 (N_19409,N_13794,N_13951);
and U19410 (N_19410,N_13476,N_12933);
or U19411 (N_19411,N_16757,N_16931);
nor U19412 (N_19412,N_15602,N_15974);
nor U19413 (N_19413,N_15180,N_16509);
nor U19414 (N_19414,N_13209,N_13287);
nor U19415 (N_19415,N_17437,N_12584);
nor U19416 (N_19416,N_15219,N_16225);
nor U19417 (N_19417,N_13412,N_12823);
or U19418 (N_19418,N_16098,N_18420);
or U19419 (N_19419,N_18698,N_14303);
nand U19420 (N_19420,N_18699,N_13558);
nor U19421 (N_19421,N_18312,N_16579);
and U19422 (N_19422,N_12544,N_14762);
nand U19423 (N_19423,N_15779,N_13842);
nand U19424 (N_19424,N_13259,N_16812);
and U19425 (N_19425,N_13791,N_17532);
nor U19426 (N_19426,N_18437,N_17755);
nor U19427 (N_19427,N_14010,N_18271);
or U19428 (N_19428,N_16117,N_16473);
or U19429 (N_19429,N_14523,N_17010);
or U19430 (N_19430,N_13615,N_16112);
or U19431 (N_19431,N_17032,N_16300);
nand U19432 (N_19432,N_17741,N_15319);
nand U19433 (N_19433,N_13397,N_13979);
or U19434 (N_19434,N_12681,N_18281);
nand U19435 (N_19435,N_12594,N_14372);
or U19436 (N_19436,N_15075,N_16816);
and U19437 (N_19437,N_13252,N_17531);
or U19438 (N_19438,N_14519,N_17753);
nor U19439 (N_19439,N_14739,N_14391);
nand U19440 (N_19440,N_14930,N_13581);
and U19441 (N_19441,N_13801,N_13017);
or U19442 (N_19442,N_16871,N_14118);
nor U19443 (N_19443,N_16660,N_18712);
nand U19444 (N_19444,N_14708,N_16593);
and U19445 (N_19445,N_13718,N_13058);
nand U19446 (N_19446,N_16720,N_13642);
nand U19447 (N_19447,N_15929,N_12640);
nand U19448 (N_19448,N_17098,N_14543);
nor U19449 (N_19449,N_18199,N_15527);
or U19450 (N_19450,N_14415,N_18201);
nor U19451 (N_19451,N_14264,N_13334);
nor U19452 (N_19452,N_18068,N_14623);
and U19453 (N_19453,N_14578,N_13917);
and U19454 (N_19454,N_18638,N_16160);
nand U19455 (N_19455,N_13521,N_14314);
and U19456 (N_19456,N_16379,N_15686);
nand U19457 (N_19457,N_16518,N_18518);
and U19458 (N_19458,N_17859,N_12631);
nor U19459 (N_19459,N_15121,N_17103);
nand U19460 (N_19460,N_14026,N_12713);
and U19461 (N_19461,N_17275,N_14277);
nor U19462 (N_19462,N_18419,N_15243);
or U19463 (N_19463,N_13217,N_14090);
or U19464 (N_19464,N_12868,N_15629);
and U19465 (N_19465,N_13024,N_13493);
or U19466 (N_19466,N_16097,N_14560);
and U19467 (N_19467,N_13954,N_15990);
nor U19468 (N_19468,N_16144,N_13636);
nor U19469 (N_19469,N_12536,N_12636);
nor U19470 (N_19470,N_15693,N_18031);
or U19471 (N_19471,N_16653,N_13249);
and U19472 (N_19472,N_16132,N_14815);
or U19473 (N_19473,N_17426,N_12776);
nand U19474 (N_19474,N_17625,N_13709);
or U19475 (N_19475,N_17905,N_14680);
and U19476 (N_19476,N_12988,N_18216);
nand U19477 (N_19477,N_13798,N_17357);
and U19478 (N_19478,N_17021,N_14598);
and U19479 (N_19479,N_13807,N_15141);
and U19480 (N_19480,N_14568,N_14978);
or U19481 (N_19481,N_14202,N_13383);
nand U19482 (N_19482,N_14811,N_18136);
and U19483 (N_19483,N_13942,N_17493);
xor U19484 (N_19484,N_12539,N_14094);
or U19485 (N_19485,N_14127,N_13835);
nand U19486 (N_19486,N_17731,N_16292);
nand U19487 (N_19487,N_16516,N_12775);
nor U19488 (N_19488,N_15829,N_12814);
nand U19489 (N_19489,N_16345,N_13050);
nand U19490 (N_19490,N_12809,N_13091);
and U19491 (N_19491,N_15613,N_15347);
and U19492 (N_19492,N_17172,N_16950);
nor U19493 (N_19493,N_14493,N_18116);
and U19494 (N_19494,N_15525,N_12736);
or U19495 (N_19495,N_17274,N_17951);
nand U19496 (N_19496,N_12968,N_18597);
or U19497 (N_19497,N_16594,N_16553);
nor U19498 (N_19498,N_13308,N_13467);
nand U19499 (N_19499,N_17997,N_17013);
nor U19500 (N_19500,N_17583,N_16942);
or U19501 (N_19501,N_17405,N_18618);
nand U19502 (N_19502,N_13517,N_17005);
and U19503 (N_19503,N_17525,N_15551);
or U19504 (N_19504,N_17990,N_17535);
nand U19505 (N_19505,N_12929,N_16228);
nand U19506 (N_19506,N_15080,N_17334);
nor U19507 (N_19507,N_13731,N_18625);
nand U19508 (N_19508,N_13133,N_14500);
nor U19509 (N_19509,N_15853,N_13912);
nor U19510 (N_19510,N_14207,N_16894);
or U19511 (N_19511,N_12512,N_18347);
nand U19512 (N_19512,N_17567,N_13079);
or U19513 (N_19513,N_17063,N_18714);
nand U19514 (N_19514,N_18431,N_14377);
nor U19515 (N_19515,N_15166,N_16701);
nor U19516 (N_19516,N_12901,N_13550);
nand U19517 (N_19517,N_16763,N_17522);
nand U19518 (N_19518,N_15446,N_12761);
or U19519 (N_19519,N_13266,N_15239);
nor U19520 (N_19520,N_13733,N_13896);
or U19521 (N_19521,N_17931,N_16014);
or U19522 (N_19522,N_18584,N_18599);
nand U19523 (N_19523,N_17744,N_14706);
nand U19524 (N_19524,N_17096,N_16202);
or U19525 (N_19525,N_16022,N_16153);
nand U19526 (N_19526,N_14149,N_17572);
or U19527 (N_19527,N_13628,N_18204);
and U19528 (N_19528,N_13795,N_15249);
and U19529 (N_19529,N_17450,N_18715);
nand U19530 (N_19530,N_17551,N_13719);
and U19531 (N_19531,N_17137,N_13023);
and U19532 (N_19532,N_15982,N_14219);
and U19533 (N_19533,N_17249,N_17740);
nand U19534 (N_19534,N_16367,N_13373);
or U19535 (N_19535,N_13559,N_14078);
nor U19536 (N_19536,N_18301,N_13385);
or U19537 (N_19537,N_13083,N_12578);
and U19538 (N_19538,N_18526,N_18667);
nand U19539 (N_19539,N_17806,N_15185);
and U19540 (N_19540,N_12858,N_13825);
nor U19541 (N_19541,N_16973,N_14412);
nand U19542 (N_19542,N_13159,N_13150);
and U19543 (N_19543,N_13784,N_12700);
nand U19544 (N_19544,N_14960,N_14673);
or U19545 (N_19545,N_16990,N_17607);
nor U19546 (N_19546,N_14853,N_17589);
and U19547 (N_19547,N_14630,N_15011);
nor U19548 (N_19548,N_16941,N_16953);
nor U19549 (N_19549,N_14088,N_13976);
or U19550 (N_19550,N_14416,N_18069);
and U19551 (N_19551,N_13271,N_15998);
nor U19552 (N_19552,N_15480,N_16815);
nand U19553 (N_19553,N_16957,N_14710);
and U19554 (N_19554,N_17380,N_16898);
or U19555 (N_19555,N_15811,N_17961);
and U19556 (N_19556,N_16256,N_14555);
nand U19557 (N_19557,N_16993,N_16328);
nand U19558 (N_19558,N_14165,N_16274);
nand U19559 (N_19559,N_17770,N_18150);
and U19560 (N_19560,N_13669,N_16204);
and U19561 (N_19561,N_18477,N_15942);
nand U19562 (N_19562,N_16507,N_17129);
or U19563 (N_19563,N_17636,N_18406);
nor U19564 (N_19564,N_14225,N_15776);
nand U19565 (N_19565,N_15256,N_13505);
nand U19566 (N_19566,N_15711,N_15585);
or U19567 (N_19567,N_17338,N_14772);
nand U19568 (N_19568,N_18585,N_14705);
nand U19569 (N_19569,N_12527,N_14509);
or U19570 (N_19570,N_16697,N_16913);
and U19571 (N_19571,N_15747,N_16208);
or U19572 (N_19572,N_18179,N_16514);
or U19573 (N_19573,N_16899,N_16069);
and U19574 (N_19574,N_17215,N_14650);
or U19575 (N_19575,N_17561,N_16534);
and U19576 (N_19576,N_17220,N_15424);
nor U19577 (N_19577,N_14054,N_18243);
or U19578 (N_19578,N_17087,N_18192);
and U19579 (N_19579,N_18725,N_15189);
and U19580 (N_19580,N_16468,N_15297);
and U19581 (N_19581,N_18212,N_16410);
nand U19582 (N_19582,N_14877,N_13858);
nor U19583 (N_19583,N_13949,N_16745);
and U19584 (N_19584,N_17917,N_13288);
nor U19585 (N_19585,N_18614,N_17023);
nand U19586 (N_19586,N_13861,N_17655);
nand U19587 (N_19587,N_15781,N_13357);
and U19588 (N_19588,N_13038,N_18079);
nand U19589 (N_19589,N_18337,N_15473);
nor U19590 (N_19590,N_15859,N_13621);
and U19591 (N_19591,N_13650,N_16248);
nand U19592 (N_19592,N_15056,N_14344);
nor U19593 (N_19593,N_17125,N_14833);
and U19594 (N_19594,N_14756,N_17619);
or U19595 (N_19595,N_15750,N_14627);
nand U19596 (N_19596,N_17210,N_16456);
and U19597 (N_19597,N_13127,N_14677);
nand U19598 (N_19598,N_13195,N_18086);
and U19599 (N_19599,N_17377,N_15157);
and U19600 (N_19600,N_18090,N_15419);
nand U19601 (N_19601,N_13782,N_13875);
nand U19602 (N_19602,N_18094,N_16859);
and U19603 (N_19603,N_15287,N_14999);
and U19604 (N_19604,N_15787,N_18622);
nor U19605 (N_19605,N_12504,N_16035);
xnor U19606 (N_19606,N_15675,N_14982);
nor U19607 (N_19607,N_14944,N_16896);
and U19608 (N_19608,N_18448,N_18188);
nor U19609 (N_19609,N_18316,N_13379);
nor U19610 (N_19610,N_15427,N_18575);
nor U19611 (N_19611,N_18252,N_17837);
and U19612 (N_19612,N_16038,N_15876);
and U19613 (N_19613,N_17243,N_15286);
nor U19614 (N_19614,N_15975,N_14153);
nand U19615 (N_19615,N_12509,N_15040);
xnor U19616 (N_19616,N_17507,N_13325);
and U19617 (N_19617,N_17856,N_13081);
nor U19618 (N_19618,N_14053,N_17513);
nor U19619 (N_19619,N_15601,N_15908);
nor U19620 (N_19620,N_13405,N_12529);
nor U19621 (N_19621,N_17839,N_18269);
nand U19622 (N_19622,N_12731,N_14849);
nand U19623 (N_19623,N_18424,N_13812);
or U19624 (N_19624,N_18323,N_13188);
nand U19625 (N_19625,N_13311,N_16453);
nor U19626 (N_19626,N_14244,N_17288);
nand U19627 (N_19627,N_15887,N_13074);
or U19628 (N_19628,N_17471,N_12647);
and U19629 (N_19629,N_16704,N_14928);
or U19630 (N_19630,N_15222,N_13645);
nand U19631 (N_19631,N_13471,N_14150);
or U19632 (N_19632,N_16319,N_17613);
nor U19633 (N_19633,N_17111,N_14155);
and U19634 (N_19634,N_17194,N_16149);
nand U19635 (N_19635,N_13052,N_13919);
nor U19636 (N_19636,N_13571,N_17120);
nor U19637 (N_19637,N_15692,N_12523);
nand U19638 (N_19638,N_18382,N_18461);
nor U19639 (N_19639,N_14629,N_16619);
nor U19640 (N_19640,N_17330,N_15579);
nor U19641 (N_19641,N_18348,N_14984);
nor U19642 (N_19642,N_15639,N_14397);
nor U19643 (N_19643,N_14501,N_18156);
nand U19644 (N_19644,N_13678,N_12545);
nor U19645 (N_19645,N_12940,N_15805);
and U19646 (N_19646,N_17119,N_17640);
nand U19647 (N_19647,N_18054,N_16912);
nand U19648 (N_19648,N_14495,N_15332);
nand U19649 (N_19649,N_13495,N_18325);
nand U19650 (N_19650,N_18262,N_14884);
nor U19651 (N_19651,N_18198,N_14617);
or U19652 (N_19652,N_13562,N_14446);
or U19653 (N_19653,N_15285,N_13867);
nor U19654 (N_19654,N_18591,N_13044);
or U19655 (N_19655,N_13435,N_14521);
nand U19656 (N_19656,N_13624,N_18295);
nand U19657 (N_19657,N_17793,N_13502);
and U19658 (N_19658,N_15571,N_15586);
nand U19659 (N_19659,N_13649,N_12601);
and U19660 (N_19660,N_14921,N_13163);
and U19661 (N_19661,N_17116,N_16070);
xor U19662 (N_19662,N_13859,N_14032);
nand U19663 (N_19663,N_16850,N_16015);
or U19664 (N_19664,N_15825,N_16085);
or U19665 (N_19665,N_14387,N_17630);
and U19666 (N_19666,N_15607,N_13509);
and U19667 (N_19667,N_17732,N_14380);
nor U19668 (N_19668,N_12563,N_17954);
and U19669 (N_19669,N_13878,N_12723);
or U19670 (N_19670,N_13696,N_13030);
nand U19671 (N_19671,N_12628,N_13750);
and U19672 (N_19672,N_14788,N_13414);
or U19673 (N_19673,N_12875,N_12813);
or U19674 (N_19674,N_15820,N_14260);
or U19675 (N_19675,N_17027,N_16998);
or U19676 (N_19676,N_14200,N_17646);
nand U19677 (N_19677,N_16681,N_18168);
or U19678 (N_19678,N_16535,N_14831);
nand U19679 (N_19679,N_16629,N_16079);
or U19680 (N_19680,N_13909,N_17296);
or U19681 (N_19681,N_17549,N_17474);
or U19682 (N_19682,N_14882,N_17586);
xor U19683 (N_19683,N_14313,N_13192);
or U19684 (N_19684,N_15822,N_12622);
or U19685 (N_19685,N_15798,N_17051);
or U19686 (N_19686,N_17771,N_15479);
or U19687 (N_19687,N_12500,N_15540);
and U19688 (N_19688,N_14608,N_13887);
and U19689 (N_19689,N_16758,N_14562);
and U19690 (N_19690,N_16305,N_18425);
nand U19691 (N_19691,N_17715,N_14108);
and U19692 (N_19692,N_15524,N_16853);
and U19693 (N_19693,N_14524,N_16524);
and U19694 (N_19694,N_14748,N_14787);
nand U19695 (N_19695,N_18032,N_15697);
nand U19696 (N_19696,N_13067,N_14981);
nor U19697 (N_19697,N_12589,N_16966);
nand U19698 (N_19698,N_17393,N_17199);
or U19699 (N_19699,N_15144,N_15683);
and U19700 (N_19700,N_12770,N_13057);
nand U19701 (N_19701,N_18082,N_15195);
nor U19702 (N_19702,N_12900,N_16617);
nor U19703 (N_19703,N_18441,N_15516);
and U19704 (N_19704,N_14048,N_16753);
nor U19705 (N_19705,N_16877,N_17203);
or U19706 (N_19706,N_12833,N_17526);
nand U19707 (N_19707,N_14951,N_13421);
and U19708 (N_19708,N_16848,N_17368);
or U19709 (N_19709,N_16063,N_16659);
nor U19710 (N_19710,N_13064,N_15625);
and U19711 (N_19711,N_13205,N_17314);
nor U19712 (N_19712,N_14886,N_12658);
and U19713 (N_19713,N_12930,N_15241);
and U19714 (N_19714,N_18242,N_12548);
and U19715 (N_19715,N_14711,N_12942);
nor U19716 (N_19716,N_12534,N_13151);
or U19717 (N_19717,N_13272,N_18384);
nand U19718 (N_19718,N_13472,N_17887);
nand U19719 (N_19719,N_18235,N_16282);
and U19720 (N_19720,N_18703,N_13992);
nand U19721 (N_19721,N_16721,N_18534);
nor U19722 (N_19722,N_16903,N_14015);
or U19723 (N_19723,N_14473,N_18152);
or U19724 (N_19724,N_15309,N_15567);
nand U19725 (N_19725,N_14058,N_16174);
xnor U19726 (N_19726,N_16892,N_15164);
or U19727 (N_19727,N_17885,N_17290);
nand U19728 (N_19728,N_15497,N_16405);
nor U19729 (N_19729,N_16324,N_18581);
or U19730 (N_19730,N_14475,N_17543);
or U19731 (N_19731,N_14091,N_16242);
nor U19732 (N_19732,N_15850,N_15969);
nor U19733 (N_19733,N_13685,N_14019);
or U19734 (N_19734,N_12787,N_14525);
nor U19735 (N_19735,N_16110,N_17202);
nor U19736 (N_19736,N_13498,N_16273);
nand U19737 (N_19737,N_16220,N_13335);
nand U19738 (N_19738,N_13315,N_17774);
or U19739 (N_19739,N_14817,N_15561);
nand U19740 (N_19740,N_15824,N_18023);
and U19741 (N_19741,N_12966,N_16472);
and U19742 (N_19742,N_16695,N_15869);
and U19743 (N_19743,N_12937,N_16310);
or U19744 (N_19744,N_18219,N_17836);
or U19745 (N_19745,N_12630,N_17664);
nand U19746 (N_19746,N_14468,N_16285);
and U19747 (N_19747,N_17673,N_17212);
nor U19748 (N_19748,N_15700,N_17047);
nand U19749 (N_19749,N_13705,N_18302);
or U19750 (N_19750,N_15921,N_17110);
or U19751 (N_19751,N_15961,N_13879);
or U19752 (N_19752,N_15832,N_15911);
and U19753 (N_19753,N_16475,N_13474);
and U19754 (N_19754,N_14463,N_14761);
nand U19755 (N_19755,N_17145,N_16829);
nand U19756 (N_19756,N_12874,N_18731);
xnor U19757 (N_19757,N_13848,N_16343);
or U19758 (N_19758,N_15466,N_17382);
or U19759 (N_19759,N_14701,N_16691);
and U19760 (N_19760,N_17928,N_13479);
nor U19761 (N_19761,N_14807,N_15554);
nand U19762 (N_19762,N_13119,N_15782);
or U19763 (N_19763,N_15354,N_15090);
and U19764 (N_19764,N_14352,N_16212);
nor U19765 (N_19765,N_18196,N_14809);
or U19766 (N_19766,N_12995,N_17626);
or U19767 (N_19767,N_14102,N_15848);
and U19768 (N_19768,N_14721,N_14968);
or U19769 (N_19769,N_13113,N_13125);
nor U19770 (N_19770,N_18660,N_14139);
nand U19771 (N_19771,N_17322,N_14393);
and U19772 (N_19772,N_18322,N_15710);
nand U19773 (N_19773,N_15114,N_14741);
nand U19774 (N_19774,N_14764,N_18127);
nand U19775 (N_19775,N_17786,N_16276);
or U19776 (N_19776,N_16984,N_16955);
xnor U19777 (N_19777,N_17181,N_14690);
or U19778 (N_19778,N_13403,N_15052);
xor U19779 (N_19779,N_13792,N_15010);
nand U19780 (N_19780,N_13831,N_15292);
or U19781 (N_19781,N_17999,N_17097);
and U19782 (N_19782,N_17115,N_16217);
nor U19783 (N_19783,N_13070,N_17348);
or U19784 (N_19784,N_15155,N_18539);
and U19785 (N_19785,N_17294,N_17242);
and U19786 (N_19786,N_18205,N_14842);
and U19787 (N_19787,N_12866,N_13652);
nor U19788 (N_19788,N_13241,N_15415);
nor U19789 (N_19789,N_14695,N_15590);
nor U19790 (N_19790,N_17853,N_17900);
and U19791 (N_19791,N_14386,N_17410);
and U19792 (N_19792,N_18389,N_12755);
or U19793 (N_19793,N_18651,N_14237);
nor U19794 (N_19794,N_16725,N_16571);
nand U19795 (N_19795,N_14649,N_17167);
or U19796 (N_19796,N_16471,N_17950);
nand U19797 (N_19797,N_14204,N_13286);
and U19798 (N_19798,N_14740,N_18493);
nand U19799 (N_19799,N_18736,N_17271);
and U19800 (N_19800,N_16567,N_16135);
and U19801 (N_19801,N_15818,N_17534);
or U19802 (N_19802,N_17910,N_12984);
or U19803 (N_19803,N_12656,N_13317);
and U19804 (N_19804,N_16154,N_18294);
and U19805 (N_19805,N_18475,N_12535);
and U19806 (N_19806,N_17190,N_14585);
and U19807 (N_19807,N_13797,N_16151);
and U19808 (N_19808,N_12740,N_14845);
and U19809 (N_19809,N_17484,N_15533);
nor U19810 (N_19810,N_13085,N_16749);
nor U19811 (N_19811,N_14538,N_17438);
or U19812 (N_19812,N_15418,N_14311);
nand U19813 (N_19813,N_18306,N_18253);
nor U19814 (N_19814,N_13947,N_15172);
nor U19815 (N_19815,N_12849,N_16349);
nor U19816 (N_19816,N_18577,N_13721);
nand U19817 (N_19817,N_14717,N_13295);
and U19818 (N_19818,N_18221,N_16232);
nand U19819 (N_19819,N_15604,N_15907);
nand U19820 (N_19820,N_14953,N_16083);
or U19821 (N_19821,N_16265,N_14418);
or U19822 (N_19822,N_13531,N_16960);
and U19823 (N_19823,N_12615,N_18489);
nand U19824 (N_19824,N_13561,N_16722);
and U19825 (N_19825,N_17482,N_13240);
nand U19826 (N_19826,N_18364,N_14369);
and U19827 (N_19827,N_17154,N_14133);
or U19828 (N_19828,N_14479,N_13116);
or U19829 (N_19829,N_15802,N_16612);
and U19830 (N_19830,N_16947,N_18040);
nand U19831 (N_19831,N_15129,N_12842);
nor U19832 (N_19832,N_18748,N_12893);
nor U19833 (N_19833,N_17736,N_15979);
nor U19834 (N_19834,N_18621,N_16092);
nand U19835 (N_19835,N_15176,N_14961);
and U19836 (N_19836,N_13829,N_13053);
or U19837 (N_19837,N_15399,N_18104);
xnor U19838 (N_19838,N_15716,N_15937);
nor U19839 (N_19839,N_13556,N_15242);
nor U19840 (N_19840,N_13485,N_15945);
and U19841 (N_19841,N_17313,N_15131);
nand U19842 (N_19842,N_16469,N_18320);
and U19843 (N_19843,N_17381,N_13852);
and U19844 (N_19844,N_16732,N_12834);
nor U19845 (N_19845,N_13442,N_13194);
and U19846 (N_19846,N_15491,N_18469);
nor U19847 (N_19847,N_13727,N_18128);
and U19848 (N_19848,N_13677,N_13783);
or U19849 (N_19849,N_17553,N_17983);
nor U19850 (N_19850,N_17090,N_13088);
nand U19851 (N_19851,N_15865,N_18541);
nor U19852 (N_19852,N_14967,N_12908);
or U19853 (N_19853,N_17762,N_13520);
nor U19854 (N_19854,N_17751,N_18041);
or U19855 (N_19855,N_17197,N_16989);
nand U19856 (N_19856,N_16253,N_18668);
nor U19857 (N_19857,N_14573,N_13730);
and U19858 (N_19858,N_18273,N_14976);
and U19859 (N_19859,N_12607,N_16462);
nand U19860 (N_19860,N_17329,N_14601);
and U19861 (N_19861,N_13123,N_16962);
nand U19862 (N_19862,N_13077,N_17323);
and U19863 (N_19863,N_13511,N_16789);
and U19864 (N_19864,N_14986,N_13989);
and U19865 (N_19865,N_17390,N_15573);
and U19866 (N_19866,N_16331,N_18733);
nor U19867 (N_19867,N_15706,N_17895);
nor U19868 (N_19868,N_15751,N_18594);
nand U19869 (N_19869,N_15368,N_14221);
and U19870 (N_19870,N_15519,N_15981);
or U19871 (N_19871,N_12926,N_13229);
nor U19872 (N_19872,N_14931,N_15840);
nand U19873 (N_19873,N_13765,N_13565);
or U19874 (N_19874,N_16446,N_13094);
and U19875 (N_19875,N_17223,N_15316);
nand U19876 (N_19876,N_12604,N_13131);
or U19877 (N_19877,N_18690,N_17726);
or U19878 (N_19878,N_18277,N_13332);
nor U19879 (N_19879,N_18132,N_18611);
or U19880 (N_19880,N_14926,N_16540);
nand U19881 (N_19881,N_12649,N_18647);
or U19882 (N_19882,N_15863,N_15729);
nand U19883 (N_19883,N_14251,N_14247);
or U19884 (N_19884,N_16381,N_18563);
and U19885 (N_19885,N_15514,N_14119);
or U19886 (N_19886,N_15765,N_15502);
nand U19887 (N_19887,N_12703,N_13420);
or U19888 (N_19888,N_18140,N_18288);
and U19889 (N_19889,N_15313,N_18561);
nand U19890 (N_19890,N_12613,N_13073);
and U19891 (N_19891,N_13738,N_18372);
or U19892 (N_19892,N_18073,N_13321);
and U19893 (N_19893,N_13007,N_17371);
nand U19894 (N_19894,N_18047,N_15338);
and U19895 (N_19895,N_12669,N_13326);
nor U19896 (N_19896,N_17277,N_16200);
nand U19897 (N_19897,N_17663,N_16371);
and U19898 (N_19898,N_13980,N_14093);
and U19899 (N_19899,N_16934,N_16556);
and U19900 (N_19900,N_13519,N_13640);
nor U19901 (N_19901,N_16759,N_16833);
nand U19902 (N_19902,N_16223,N_16096);
and U19903 (N_19903,N_16357,N_14072);
or U19904 (N_19904,N_14064,N_16416);
nand U19905 (N_19905,N_13410,N_12744);
or U19906 (N_19906,N_17665,N_12603);
or U19907 (N_19907,N_15498,N_13890);
nor U19908 (N_19908,N_13361,N_16433);
nand U19909 (N_19909,N_17444,N_17569);
nor U19910 (N_19910,N_18254,N_17089);
nand U19911 (N_19911,N_18573,N_17854);
nand U19912 (N_19912,N_13543,N_15344);
nand U19913 (N_19913,N_14068,N_13345);
or U19914 (N_19914,N_17867,N_15753);
nand U19915 (N_19915,N_17460,N_18165);
nor U19916 (N_19916,N_16726,N_17174);
or U19917 (N_19917,N_12955,N_14183);
nand U19918 (N_19918,N_17874,N_16511);
and U19919 (N_19919,N_13078,N_13820);
and U19920 (N_19920,N_15817,N_12511);
nor U19921 (N_19921,N_18362,N_15946);
or U19922 (N_19922,N_14520,N_15191);
nor U19923 (N_19923,N_17457,N_18675);
xor U19924 (N_19924,N_13166,N_15198);
xor U19925 (N_19925,N_16790,N_16808);
or U19926 (N_19926,N_16728,N_15658);
or U19927 (N_19927,N_14233,N_15915);
and U19928 (N_19928,N_17214,N_18727);
nor U19929 (N_19929,N_13353,N_15530);
and U19930 (N_19930,N_13482,N_13323);
nor U19931 (N_19931,N_16699,N_13548);
nor U19932 (N_19932,N_12785,N_12781);
or U19933 (N_19933,N_15723,N_16711);
and U19934 (N_19934,N_18747,N_13423);
or U19935 (N_19935,N_12522,N_13608);
and U19936 (N_19936,N_14160,N_12779);
and U19937 (N_19937,N_15739,N_15230);
or U19938 (N_19938,N_15362,N_14871);
or U19939 (N_19939,N_15603,N_13893);
nor U19940 (N_19940,N_17445,N_15646);
and U19941 (N_19941,N_15870,N_14566);
and U19942 (N_19942,N_12772,N_16761);
nor U19943 (N_19943,N_17041,N_13943);
or U19944 (N_19944,N_15630,N_17291);
and U19945 (N_19945,N_12935,N_13456);
and U19946 (N_19946,N_17473,N_17907);
and U19947 (N_19947,N_17725,N_18488);
nand U19948 (N_19948,N_18658,N_18270);
nor U19949 (N_19949,N_13002,N_17785);
nand U19950 (N_19950,N_16607,N_13905);
or U19951 (N_19951,N_14217,N_12943);
or U19952 (N_19952,N_13546,N_16056);
and U19953 (N_19953,N_15238,N_18485);
nand U19954 (N_19954,N_16120,N_13371);
or U19955 (N_19955,N_14506,N_18387);
and U19956 (N_19956,N_13981,N_15632);
nand U19957 (N_19957,N_18642,N_12825);
nand U19958 (N_19958,N_16544,N_18363);
and U19959 (N_19959,N_16046,N_16169);
nor U19960 (N_19960,N_13389,N_16712);
nor U19961 (N_19961,N_16865,N_15517);
or U19962 (N_19962,N_12827,N_14002);
nand U19963 (N_19963,N_15460,N_15701);
or U19964 (N_19964,N_15790,N_13884);
and U19965 (N_19965,N_13069,N_18521);
nand U19966 (N_19966,N_14235,N_14289);
nor U19967 (N_19967,N_15559,N_17342);
or U19968 (N_19968,N_17915,N_17529);
nand U19969 (N_19969,N_14012,N_16976);
nor U19970 (N_19970,N_18603,N_12557);
nand U19971 (N_19971,N_13212,N_17245);
nor U19972 (N_19972,N_15318,N_17575);
nor U19973 (N_19973,N_13631,N_13244);
nor U19974 (N_19974,N_15719,N_15359);
nand U19975 (N_19975,N_14232,N_14399);
and U19976 (N_19976,N_16443,N_15522);
and U19977 (N_19977,N_18161,N_17050);
or U19978 (N_19978,N_18145,N_14934);
and U19979 (N_19979,N_15486,N_13176);
or U19980 (N_19980,N_16229,N_17515);
and U19981 (N_19981,N_14747,N_15599);
and U19982 (N_19982,N_12838,N_18026);
nand U19983 (N_19983,N_17000,N_16922);
or U19984 (N_19984,N_17686,N_16747);
and U19985 (N_19985,N_17229,N_15085);
or U19986 (N_19986,N_16123,N_16125);
and U19987 (N_19987,N_15371,N_17896);
xor U19988 (N_19988,N_12575,N_14324);
or U19989 (N_19989,N_14196,N_14211);
nor U19990 (N_19990,N_18500,N_13384);
nand U19991 (N_19991,N_15717,N_13518);
and U19992 (N_19992,N_18010,N_16830);
nand U19993 (N_19993,N_13043,N_17579);
and U19994 (N_19994,N_16358,N_14282);
nor U19995 (N_19995,N_16768,N_16951);
nor U19996 (N_19996,N_13433,N_18438);
or U19997 (N_19997,N_16805,N_16568);
nand U19998 (N_19998,N_13599,N_17822);
or U19999 (N_19999,N_15363,N_14854);
nor U20000 (N_20000,N_14559,N_14733);
nand U20001 (N_20001,N_17881,N_18081);
or U20002 (N_20002,N_14542,N_14803);
nor U20003 (N_20003,N_16155,N_17289);
nand U20004 (N_20004,N_15587,N_16814);
and U20005 (N_20005,N_18096,N_16963);
nand U20006 (N_20006,N_15891,N_17564);
and U20007 (N_20007,N_14009,N_12567);
nor U20008 (N_20008,N_13598,N_16450);
and U20009 (N_20009,N_17121,N_17187);
nor U20010 (N_20010,N_18338,N_14681);
nand U20011 (N_20011,N_16801,N_13175);
or U20012 (N_20012,N_17706,N_16064);
or U20013 (N_20013,N_12707,N_14145);
and U20014 (N_20014,N_17106,N_18332);
nor U20015 (N_20015,N_14226,N_13051);
or U20016 (N_20016,N_18123,N_15204);
nor U20017 (N_20017,N_14876,N_13880);
or U20018 (N_20018,N_17738,N_18351);
or U20019 (N_20019,N_15631,N_14096);
nand U20020 (N_20020,N_13915,N_14791);
nor U20021 (N_20021,N_16074,N_14355);
and U20022 (N_20022,N_14963,N_15305);
nor U20023 (N_20023,N_14702,N_14634);
nor U20024 (N_20024,N_15177,N_12680);
and U20025 (N_20025,N_15348,N_16783);
nand U20026 (N_20026,N_18317,N_13841);
nand U20027 (N_20027,N_13619,N_17791);
or U20028 (N_20028,N_13183,N_18261);
nor U20029 (N_20029,N_15511,N_18022);
nor U20030 (N_20030,N_14481,N_12951);
or U20031 (N_20031,N_14729,N_16703);
or U20032 (N_20032,N_15896,N_17141);
or U20033 (N_20033,N_12549,N_17038);
or U20034 (N_20034,N_14851,N_16991);
or U20035 (N_20035,N_13204,N_17045);
and U20036 (N_20036,N_15076,N_12888);
nand U20037 (N_20037,N_16970,N_17571);
nor U20038 (N_20038,N_18471,N_17711);
and U20039 (N_20039,N_14162,N_16352);
nor U20040 (N_20040,N_15923,N_16936);
nor U20041 (N_20041,N_18135,N_13466);
nand U20042 (N_20042,N_18274,N_18213);
nor U20043 (N_20043,N_12803,N_13096);
nor U20044 (N_20044,N_15581,N_12965);
or U20045 (N_20045,N_12880,N_13066);
nand U20046 (N_20046,N_12665,N_16080);
nand U20047 (N_20047,N_15421,N_13946);
and U20048 (N_20048,N_17099,N_13945);
nor U20049 (N_20049,N_13764,N_17344);
nor U20050 (N_20050,N_14356,N_16551);
or U20051 (N_20051,N_16148,N_16434);
or U20052 (N_20052,N_15214,N_15566);
and U20053 (N_20053,N_15912,N_17364);
nand U20054 (N_20054,N_17972,N_13757);
nor U20055 (N_20055,N_14001,N_15978);
nor U20056 (N_20056,N_16944,N_14158);
or U20057 (N_20057,N_18457,N_16777);
or U20058 (N_20058,N_18051,N_16862);
nand U20059 (N_20059,N_16840,N_14873);
nor U20060 (N_20060,N_17902,N_17015);
nor U20061 (N_20061,N_15456,N_18624);
nand U20062 (N_20062,N_14507,N_15132);
nand U20063 (N_20063,N_13355,N_13646);
and U20064 (N_20064,N_17992,N_18707);
nor U20065 (N_20065,N_16295,N_12961);
nand U20066 (N_20066,N_16585,N_16166);
or U20067 (N_20067,N_16570,N_15261);
and U20068 (N_20068,N_16661,N_17752);
xnor U20069 (N_20069,N_12588,N_14699);
nand U20070 (N_20070,N_16213,N_18590);
nand U20071 (N_20071,N_15216,N_15275);
and U20072 (N_20072,N_14185,N_13022);
nand U20073 (N_20073,N_16128,N_17439);
nand U20074 (N_20074,N_14938,N_17974);
or U20075 (N_20075,N_14368,N_16543);
nand U20076 (N_20076,N_13439,N_13644);
or U20077 (N_20077,N_17191,N_17086);
and U20078 (N_20078,N_13754,N_14239);
or U20079 (N_20079,N_14644,N_18177);
and U20080 (N_20080,N_13637,N_13228);
and U20081 (N_20081,N_13161,N_13029);
or U20082 (N_20082,N_14952,N_14645);
nor U20083 (N_20083,N_16197,N_18334);
and U20084 (N_20084,N_18492,N_16652);
or U20085 (N_20085,N_17733,N_17179);
nand U20086 (N_20086,N_14348,N_14813);
nand U20087 (N_20087,N_16548,N_16437);
nand U20088 (N_20088,N_18287,N_18122);
and U20089 (N_20089,N_14808,N_14823);
nand U20090 (N_20090,N_17984,N_16766);
nand U20091 (N_20091,N_13333,N_13702);
or U20092 (N_20092,N_17544,N_13540);
nor U20093 (N_20093,N_16127,N_16557);
and U20094 (N_20094,N_17631,N_17458);
or U20095 (N_20095,N_14103,N_14214);
nor U20096 (N_20096,N_12863,N_12854);
and U20097 (N_20097,N_18166,N_14812);
or U20098 (N_20098,N_13185,N_13895);
nor U20099 (N_20099,N_13213,N_15260);
or U20100 (N_20100,N_13882,N_15438);
nor U20101 (N_20101,N_15868,N_18148);
nor U20102 (N_20102,N_13690,N_14948);
nor U20103 (N_20103,N_16588,N_14974);
nand U20104 (N_20104,N_15008,N_12683);
and U20105 (N_20105,N_14602,N_16895);
and U20106 (N_20106,N_13973,N_13399);
and U20107 (N_20107,N_15109,N_14624);
nand U20108 (N_20108,N_13449,N_17798);
nand U20109 (N_20109,N_17372,N_13725);
nand U20110 (N_20110,N_18157,N_14117);
or U20111 (N_20111,N_13932,N_17394);
and U20112 (N_20112,N_14037,N_16454);
nor U20113 (N_20113,N_17435,N_14942);
nor U20114 (N_20114,N_16000,N_15406);
nor U20115 (N_20115,N_15833,N_12879);
nand U20116 (N_20116,N_14997,N_15062);
nand U20117 (N_20117,N_15078,N_16506);
and U20118 (N_20118,N_13490,N_17766);
nor U20119 (N_20119,N_16879,N_15930);
xor U20120 (N_20120,N_14402,N_15720);
nand U20121 (N_20121,N_14024,N_15310);
and U20122 (N_20122,N_16278,N_16824);
nor U20123 (N_20123,N_17404,N_15367);
and U20124 (N_20124,N_15389,N_15851);
and U20125 (N_20125,N_18103,N_14038);
nor U20126 (N_20126,N_15187,N_17878);
nor U20127 (N_20127,N_13800,N_16303);
nor U20128 (N_20128,N_16118,N_17073);
and U20129 (N_20129,N_16624,N_14231);
and U20130 (N_20130,N_13310,N_14407);
nand U20131 (N_20131,N_14508,N_15989);
or U20132 (N_20132,N_12739,N_16743);
nand U20133 (N_20133,N_13747,N_15759);
and U20134 (N_20134,N_17095,N_14490);
nand U20135 (N_20135,N_16187,N_12558);
nor U20136 (N_20136,N_18486,N_14062);
or U20137 (N_20137,N_13297,N_12972);
nand U20138 (N_20138,N_13274,N_17483);
and U20139 (N_20139,N_13341,N_18278);
nand U20140 (N_20140,N_16398,N_16522);
nand U20141 (N_20141,N_13189,N_15689);
or U20142 (N_20142,N_18559,N_13734);
xor U20143 (N_20143,N_13218,N_14626);
nor U20144 (N_20144,N_16700,N_17472);
nand U20145 (N_20145,N_16715,N_12597);
and U20146 (N_20146,N_14687,N_14488);
nand U20147 (N_20147,N_17497,N_17669);
nand U20148 (N_20148,N_13496,N_12678);
or U20149 (N_20149,N_14483,N_13318);
nand U20150 (N_20150,N_17088,N_16284);
and U20151 (N_20151,N_15652,N_13265);
and U20152 (N_20152,N_16403,N_18665);
and U20153 (N_20153,N_18111,N_15866);
nor U20154 (N_20154,N_14478,N_17645);
nor U20155 (N_20155,N_18646,N_18499);
or U20156 (N_20156,N_14100,N_12598);
nand U20157 (N_20157,N_15741,N_14253);
or U20158 (N_20158,N_13084,N_15788);
or U20159 (N_20159,N_14069,N_13395);
or U20160 (N_20160,N_16271,N_13121);
nor U20161 (N_20161,N_16291,N_17462);
nor U20162 (N_20162,N_18571,N_15208);
nand U20163 (N_20163,N_14034,N_17292);
and U20164 (N_20164,N_17944,N_13006);
and U20165 (N_20165,N_14109,N_15771);
or U20166 (N_20166,N_14027,N_17789);
nor U20167 (N_20167,N_18296,N_15248);
nand U20168 (N_20168,N_16974,N_14619);
or U20169 (N_20169,N_16011,N_18421);
nand U20170 (N_20170,N_17901,N_14210);
and U20171 (N_20171,N_17467,N_14474);
and U20172 (N_20172,N_16981,N_16176);
or U20173 (N_20173,N_15009,N_14115);
and U20174 (N_20174,N_15162,N_18239);
nor U20175 (N_20175,N_18435,N_12925);
and U20176 (N_20176,N_18374,N_14724);
nand U20177 (N_20177,N_12820,N_14731);
and U20178 (N_20178,N_18596,N_12887);
nor U20179 (N_20179,N_16538,N_13016);
or U20180 (N_20180,N_15165,N_13874);
or U20181 (N_20181,N_14547,N_17180);
nor U20182 (N_20182,N_16267,N_18695);
nor U20183 (N_20183,N_15146,N_18227);
and U20184 (N_20184,N_14175,N_13147);
nand U20185 (N_20185,N_18551,N_15127);
nand U20186 (N_20186,N_17748,N_14309);
nor U20187 (N_20187,N_14751,N_18694);
nand U20188 (N_20188,N_14195,N_14962);
nand U20189 (N_20189,N_16099,N_18222);
nand U20190 (N_20190,N_12948,N_14063);
nand U20191 (N_20191,N_17056,N_15197);
nor U20192 (N_20192,N_16623,N_17709);
or U20193 (N_20193,N_13589,N_14454);
and U20194 (N_20194,N_17412,N_17848);
nand U20195 (N_20195,N_13100,N_15501);
nand U20196 (N_20196,N_17548,N_15862);
nand U20197 (N_20197,N_17503,N_15925);
nand U20198 (N_20198,N_14939,N_17152);
nor U20199 (N_20199,N_13866,N_18403);
or U20200 (N_20200,N_17521,N_15864);
or U20201 (N_20201,N_17301,N_17970);
nand U20202 (N_20202,N_14332,N_16515);
nand U20203 (N_20203,N_17560,N_15454);
nor U20204 (N_20204,N_14444,N_15543);
nand U20205 (N_20205,N_14178,N_16904);
nor U20206 (N_20206,N_13402,N_14527);
nand U20207 (N_20207,N_15721,N_13162);
and U20208 (N_20208,N_15271,N_17781);
nor U20209 (N_20209,N_15648,N_17107);
and U20210 (N_20210,N_13944,N_12958);
nand U20211 (N_20211,N_13766,N_16423);
nand U20212 (N_20212,N_14536,N_17016);
and U20213 (N_20213,N_13799,N_13788);
xor U20214 (N_20214,N_14374,N_17501);
nor U20215 (N_20215,N_13921,N_16483);
nor U20216 (N_20216,N_15361,N_15633);
and U20217 (N_20217,N_16477,N_18098);
nor U20218 (N_20218,N_15320,N_14925);
nor U20219 (N_20219,N_16741,N_13010);
and U20220 (N_20220,N_17475,N_12784);
nor U20221 (N_20221,N_12729,N_15801);
nor U20222 (N_20222,N_13142,N_14301);
and U20223 (N_20223,N_16047,N_17227);
and U20224 (N_20224,N_14937,N_13093);
nand U20225 (N_20225,N_18661,N_14652);
nand U20226 (N_20226,N_18093,N_14971);
nand U20227 (N_20227,N_15125,N_15944);
nor U20228 (N_20228,N_18709,N_14151);
xnor U20229 (N_20229,N_14584,N_18627);
nor U20230 (N_20230,N_16559,N_17652);
nand U20231 (N_20231,N_13469,N_12710);
or U20232 (N_20232,N_17875,N_17008);
or U20233 (N_20233,N_12778,N_13714);
or U20234 (N_20234,N_18412,N_17816);
or U20235 (N_20235,N_13365,N_12938);
nand U20236 (N_20236,N_14227,N_14130);
and U20237 (N_20237,N_12767,N_13625);
nor U20238 (N_20238,N_15443,N_13802);
nand U20239 (N_20239,N_13021,N_15970);
or U20240 (N_20240,N_15449,N_12705);
and U20241 (N_20241,N_15699,N_18101);
nand U20242 (N_20242,N_13222,N_14893);
and U20243 (N_20243,N_12653,N_14760);
or U20244 (N_20244,N_15001,N_18191);
or U20245 (N_20245,N_16407,N_13665);
or U20246 (N_20246,N_12666,N_17355);
nor U20247 (N_20247,N_17332,N_14906);
or U20248 (N_20248,N_16314,N_14727);
and U20249 (N_20249,N_15904,N_13901);
or U20250 (N_20250,N_16591,N_14371);
or U20251 (N_20251,N_17456,N_18515);
and U20252 (N_20252,N_17061,N_12570);
and U20253 (N_20253,N_13282,N_18021);
and U20254 (N_20254,N_16178,N_18495);
or U20255 (N_20255,N_15941,N_17452);
or U20256 (N_20256,N_14916,N_18512);
and U20257 (N_20257,N_14189,N_13845);
nor U20258 (N_20258,N_14697,N_15336);
or U20259 (N_20259,N_17101,N_15212);
nor U20260 (N_20260,N_14299,N_16893);
nand U20261 (N_20261,N_15654,N_15158);
or U20262 (N_20262,N_13934,N_12619);
nor U20263 (N_20263,N_15311,N_14020);
and U20264 (N_20264,N_12528,N_13759);
or U20265 (N_20265,N_17226,N_15992);
or U20266 (N_20266,N_15608,N_15569);
or U20267 (N_20267,N_13082,N_14661);
and U20268 (N_20268,N_12547,N_16785);
nor U20269 (N_20269,N_18380,N_16834);
nor U20270 (N_20270,N_14919,N_13104);
nand U20271 (N_20271,N_14569,N_13953);
and U20272 (N_20272,N_13955,N_15098);
nor U20273 (N_20273,N_16058,N_18513);
and U20274 (N_20274,N_16138,N_17923);
nand U20275 (N_20275,N_17932,N_14075);
or U20276 (N_20276,N_12795,N_15668);
nor U20277 (N_20277,N_16573,N_13269);
xor U20278 (N_20278,N_14819,N_15667);
or U20279 (N_20279,N_18386,N_17872);
and U20280 (N_20280,N_13735,N_13042);
or U20281 (N_20281,N_16948,N_16071);
or U20282 (N_20282,N_14146,N_18579);
or U20283 (N_20283,N_13554,N_13888);
and U20284 (N_20284,N_18214,N_13567);
or U20285 (N_20285,N_16605,N_16972);
nor U20286 (N_20286,N_12556,N_15952);
or U20287 (N_20287,N_15785,N_17065);
or U20288 (N_20288,N_17721,N_16552);
and U20289 (N_20289,N_18567,N_13428);
nor U20290 (N_20290,N_16613,N_14465);
and U20291 (N_20291,N_14686,N_16887);
or U20292 (N_20292,N_13741,N_18659);
nand U20293 (N_20293,N_16954,N_14888);
or U20294 (N_20294,N_13817,N_18360);
or U20295 (N_20295,N_15401,N_16459);
nand U20296 (N_20296,N_18467,N_16542);
nand U20297 (N_20297,N_14684,N_12638);
nand U20298 (N_20298,N_13138,N_13593);
nand U20299 (N_20299,N_15215,N_14637);
nor U20300 (N_20300,N_14176,N_17884);
nor U20301 (N_20301,N_13684,N_12542);
or U20302 (N_20302,N_13239,N_14814);
nor U20303 (N_20303,N_14476,N_14614);
nand U20304 (N_20304,N_13720,N_16943);
and U20305 (N_20305,N_14280,N_17759);
nand U20306 (N_20306,N_12616,N_13092);
and U20307 (N_20307,N_15073,N_17565);
nor U20308 (N_20308,N_12869,N_18035);
and U20309 (N_20309,N_14095,N_13120);
nor U20310 (N_20310,N_12934,N_16024);
nand U20311 (N_20311,N_13015,N_15358);
nand U20312 (N_20312,N_14949,N_17429);
and U20313 (N_20313,N_14834,N_15823);
nand U20314 (N_20314,N_13172,N_13933);
and U20315 (N_20315,N_18118,N_16003);
nand U20316 (N_20316,N_13037,N_15836);
and U20317 (N_20317,N_18176,N_13523);
and U20318 (N_20318,N_14031,N_17530);
or U20319 (N_20319,N_13697,N_13891);
nor U20320 (N_20320,N_14070,N_13307);
xnor U20321 (N_20321,N_15031,N_17833);
nor U20322 (N_20322,N_17746,N_13902);
nor U20323 (N_20323,N_12633,N_15705);
nor U20324 (N_20324,N_15288,N_16986);
nand U20325 (N_20325,N_15827,N_17899);
nor U20326 (N_20326,N_15398,N_16323);
nor U20327 (N_20327,N_15381,N_12890);
nand U20328 (N_20328,N_14134,N_14770);
or U20329 (N_20329,N_15303,N_14822);
nand U20330 (N_20330,N_15134,N_14628);
nand U20331 (N_20331,N_15390,N_13430);
and U20332 (N_20332,N_15531,N_12902);
nand U20333 (N_20333,N_18705,N_17941);
nor U20334 (N_20334,N_14620,N_16854);
or U20335 (N_20335,N_17012,N_16246);
nand U20336 (N_20336,N_15321,N_16798);
nor U20337 (N_20337,N_13928,N_15207);
and U20338 (N_20338,N_18065,N_14837);
nor U20339 (N_20339,N_13025,N_16835);
nand U20340 (N_20340,N_15819,N_17911);
and U20341 (N_20341,N_18042,N_18710);
nand U20342 (N_20342,N_14438,N_13109);
or U20343 (N_20343,N_13140,N_18056);
nor U20344 (N_20344,N_18447,N_14783);
nor U20345 (N_20345,N_14752,N_17605);
and U20346 (N_20346,N_17632,N_18595);
and U20347 (N_20347,N_16363,N_13692);
nor U20348 (N_20348,N_15289,N_14036);
nand U20349 (N_20349,N_17228,N_16576);
nor U20350 (N_20350,N_16180,N_15252);
nand U20351 (N_20351,N_15276,N_17360);
and U20352 (N_20352,N_15588,N_18491);
or U20353 (N_20353,N_12577,N_15229);
xnor U20354 (N_20354,N_13525,N_12994);
xor U20355 (N_20355,N_17485,N_17637);
nor U20356 (N_20356,N_14343,N_13994);
nor U20357 (N_20357,N_17030,N_14285);
nand U20358 (N_20358,N_17591,N_16104);
nor U20359 (N_20359,N_13202,N_17310);
nor U20360 (N_20360,N_17695,N_17325);
nand U20361 (N_20361,N_13507,N_18578);
nand U20362 (N_20362,N_12818,N_16141);
and U20363 (N_20363,N_15130,N_18012);
or U20364 (N_20364,N_14959,N_12600);
nand U20365 (N_20365,N_13261,N_13107);
and U20366 (N_20366,N_13227,N_13290);
and U20367 (N_20367,N_13004,N_15471);
nand U20368 (N_20368,N_13391,N_14640);
and U20369 (N_20369,N_14051,N_12947);
nand U20370 (N_20370,N_13145,N_15534);
nand U20371 (N_20371,N_15267,N_16302);
or U20372 (N_20372,N_14579,N_14737);
and U20373 (N_20373,N_15873,N_14970);
nand U20374 (N_20374,N_15077,N_15269);
nor U20375 (N_20375,N_14267,N_12830);
nor U20376 (N_20376,N_14420,N_14526);
or U20377 (N_20377,N_13689,N_13432);
nand U20378 (N_20378,N_14113,N_14294);
and U20379 (N_20379,N_13009,N_16574);
and U20380 (N_20380,N_14895,N_14832);
and U20381 (N_20381,N_18028,N_18604);
or U20382 (N_20382,N_13483,N_15295);
nand U20383 (N_20383,N_16569,N_12997);
nor U20384 (N_20384,N_14941,N_14192);
nand U20385 (N_20385,N_18335,N_18416);
or U20386 (N_20386,N_14659,N_17114);
or U20387 (N_20387,N_16842,N_13547);
nor U20388 (N_20388,N_12892,N_17809);
nor U20389 (N_20389,N_17829,N_13281);
or U20390 (N_20390,N_14664,N_16031);
and U20391 (N_20391,N_15895,N_14310);
nor U20392 (N_20392,N_13903,N_16499);
or U20393 (N_20393,N_17049,N_16075);
and U20394 (N_20394,N_16388,N_14331);
nor U20395 (N_20395,N_16447,N_15902);
nor U20396 (N_20396,N_16325,N_14269);
nand U20397 (N_20397,N_17319,N_17658);
nor U20398 (N_20398,N_13931,N_18687);
nand U20399 (N_20399,N_16439,N_16218);
and U20400 (N_20400,N_14972,N_13974);
or U20401 (N_20401,N_16851,N_18548);
or U20402 (N_20402,N_15642,N_18637);
and U20403 (N_20403,N_16577,N_12924);
nand U20404 (N_20404,N_12596,N_13299);
nand U20405 (N_20405,N_18071,N_13060);
nand U20406 (N_20406,N_16374,N_14663);
nand U20407 (N_20407,N_15202,N_17536);
and U20408 (N_20408,N_14215,N_12555);
nand U20409 (N_20409,N_15447,N_18693);
xnor U20410 (N_20410,N_14790,N_16918);
nor U20411 (N_20411,N_18532,N_13278);
or U20412 (N_20412,N_13762,N_17158);
and U20413 (N_20413,N_17201,N_16039);
and U20414 (N_20414,N_15397,N_13839);
nand U20415 (N_20415,N_13541,N_17953);
nand U20416 (N_20416,N_16452,N_16928);
xnor U20417 (N_20417,N_15346,N_16095);
or U20418 (N_20418,N_14006,N_15255);
or U20419 (N_20419,N_16382,N_14504);
nor U20420 (N_20420,N_17150,N_13937);
nor U20421 (N_20421,N_15349,N_12644);
and U20422 (N_20422,N_18588,N_15773);
nand U20423 (N_20423,N_14384,N_13168);
or U20424 (N_20424,N_16081,N_15182);
or U20425 (N_20425,N_16108,N_15044);
nand U20426 (N_20426,N_17006,N_17812);
and U20427 (N_20427,N_15474,N_18077);
nand U20428 (N_20428,N_16336,N_17908);
and U20429 (N_20429,N_14364,N_16655);
and U20430 (N_20430,N_13415,N_12821);
xor U20431 (N_20431,N_16401,N_18735);
nor U20432 (N_20432,N_18247,N_17557);
and U20433 (N_20433,N_14016,N_13360);
and U20434 (N_20434,N_17775,N_16093);
nor U20435 (N_20435,N_17898,N_13927);
and U20436 (N_20436,N_17688,N_13708);
nor U20437 (N_20437,N_15558,N_16170);
nor U20438 (N_20438,N_18537,N_18005);
and U20439 (N_20439,N_13960,N_17880);
nand U20440 (N_20440,N_17204,N_17336);
and U20441 (N_20441,N_13298,N_13190);
or U20442 (N_20442,N_13653,N_14445);
nand U20443 (N_20443,N_16142,N_17053);
and U20444 (N_20444,N_13343,N_17293);
nand U20445 (N_20445,N_16529,N_16061);
nor U20446 (N_20446,N_17869,N_14462);
nor U20447 (N_20447,N_16240,N_14550);
and U20448 (N_20448,N_16191,N_18300);
or U20449 (N_20449,N_14753,N_14541);
nor U20450 (N_20450,N_14612,N_16198);
and U20451 (N_20451,N_16849,N_14826);
or U20452 (N_20452,N_17109,N_16536);
or U20453 (N_20453,N_13963,N_13846);
or U20454 (N_20454,N_18304,N_18696);
nand U20455 (N_20455,N_16911,N_15886);
or U20456 (N_20456,N_16669,N_14835);
or U20457 (N_20457,N_17903,N_14994);
nand U20458 (N_20458,N_16891,N_14958);
nor U20459 (N_20459,N_14336,N_14453);
nand U20460 (N_20460,N_18024,N_18440);
or U20461 (N_20461,N_17417,N_17036);
or U20462 (N_20462,N_16890,N_12862);
and U20463 (N_20463,N_18142,N_17260);
or U20464 (N_20464,N_15556,N_14973);
and U20465 (N_20465,N_16372,N_17920);
nor U20466 (N_20466,N_14140,N_17396);
nor U20467 (N_20467,N_15499,N_17490);
or U20468 (N_20468,N_15372,N_13818);
nor U20469 (N_20469,N_13279,N_12800);
nor U20470 (N_20470,N_18248,N_17803);
and U20471 (N_20471,N_16632,N_17198);
nor U20472 (N_20472,N_15560,N_12562);
nand U20473 (N_20473,N_12963,N_17584);
nand U20474 (N_20474,N_13855,N_13938);
and U20475 (N_20475,N_18141,N_17184);
and U20476 (N_20476,N_18681,N_15881);
nor U20477 (N_20477,N_13700,N_12609);
and U20478 (N_20478,N_17754,N_16831);
nand U20479 (N_20479,N_14112,N_14424);
or U20480 (N_20480,N_13489,N_14647);
nand U20481 (N_20481,N_12918,N_17966);
and U20482 (N_20482,N_15784,N_17842);
nand U20483 (N_20483,N_18602,N_15532);
nor U20484 (N_20484,N_14712,N_18410);
nor U20485 (N_20485,N_17183,N_17378);
and U20486 (N_20486,N_17841,N_15803);
or U20487 (N_20487,N_15104,N_18131);
or U20488 (N_20488,N_18133,N_17862);
nor U20489 (N_20489,N_13940,N_17383);
or U20490 (N_20490,N_15726,N_15096);
nor U20491 (N_20491,N_17935,N_17100);
or U20492 (N_20492,N_13657,N_18691);
and U20493 (N_20493,N_17176,N_17524);
nand U20494 (N_20494,N_15656,N_14700);
nor U20495 (N_20495,N_16492,N_14389);
and U20496 (N_20496,N_15591,N_17080);
or U20497 (N_20497,N_15983,N_16173);
or U20498 (N_20498,N_14451,N_16234);
or U20499 (N_20499,N_13576,N_17892);
nor U20500 (N_20500,N_15100,N_15268);
and U20501 (N_20501,N_14932,N_13234);
nand U20502 (N_20502,N_16320,N_17466);
and U20503 (N_20503,N_16329,N_16638);
xnor U20504 (N_20504,N_13803,N_17258);
or U20505 (N_20505,N_16408,N_14929);
or U20506 (N_20506,N_16939,N_14904);
and U20507 (N_20507,N_17758,N_12586);
and U20508 (N_20508,N_15575,N_15893);
nor U20509 (N_20509,N_12554,N_15133);
nand U20510 (N_20510,N_15209,N_17208);
and U20511 (N_20511,N_16342,N_15512);
nand U20512 (N_20512,N_17677,N_13224);
and U20513 (N_20513,N_14998,N_15894);
and U20514 (N_20514,N_14656,N_15435);
nor U20515 (N_20515,N_16772,N_12514);
or U20516 (N_20516,N_16364,N_16426);
nand U20517 (N_20517,N_18636,N_14410);
or U20518 (N_20518,N_13165,N_15493);
nand U20519 (N_20519,N_16675,N_18697);
nor U20520 (N_20520,N_13753,N_16377);
nand U20521 (N_20521,N_14159,N_14591);
nand U20522 (N_20522,N_15674,N_18207);
nor U20523 (N_20523,N_15826,N_18568);
nor U20524 (N_20524,N_14005,N_17076);
and U20525 (N_20525,N_17685,N_15218);
and U20526 (N_20526,N_15194,N_14830);
nor U20527 (N_20527,N_12750,N_17488);
nor U20528 (N_20528,N_18662,N_14358);
or U20529 (N_20529,N_12903,N_14716);
nor U20530 (N_20530,N_14979,N_14136);
or U20531 (N_20531,N_14046,N_12952);
nand U20532 (N_20532,N_13588,N_15453);
nand U20533 (N_20533,N_12916,N_15783);
xnor U20534 (N_20534,N_15071,N_13461);
or U20535 (N_20535,N_14171,N_16044);
nand U20536 (N_20536,N_16236,N_12749);
or U20537 (N_20537,N_15385,N_16296);
and U20538 (N_20538,N_15174,N_15217);
nand U20539 (N_20539,N_14270,N_18173);
and U20540 (N_20540,N_14869,N_17128);
nor U20541 (N_20541,N_18683,N_14017);
nand U20542 (N_20542,N_13380,N_15184);
nand U20543 (N_20543,N_15391,N_18724);
nor U20544 (N_20544,N_13844,N_13296);
nand U20545 (N_20545,N_15352,N_12985);
or U20546 (N_20546,N_16926,N_18562);
nor U20547 (N_20547,N_14867,N_12635);
nor U20548 (N_20548,N_14203,N_13101);
nand U20549 (N_20549,N_16417,N_18645);
nor U20550 (N_20550,N_15838,N_15068);
nor U20551 (N_20551,N_15116,N_17614);
nor U20552 (N_20552,N_13889,N_18640);
or U20553 (N_20553,N_16839,N_18309);
nand U20554 (N_20554,N_13072,N_16073);
nor U20555 (N_20555,N_12871,N_16482);
or U20556 (N_20556,N_13821,N_18401);
and U20557 (N_20557,N_12754,N_12894);
and U20558 (N_20558,N_15777,N_16686);
and U20559 (N_20559,N_13563,N_15640);
or U20560 (N_20560,N_14688,N_13246);
and U20561 (N_20561,N_12540,N_16387);
nand U20562 (N_20562,N_13219,N_18708);
nor U20563 (N_20563,N_12526,N_14296);
and U20564 (N_20564,N_12660,N_14179);
or U20565 (N_20565,N_14447,N_14715);
nand U20566 (N_20566,N_16882,N_14392);
and U20567 (N_20567,N_15909,N_14648);
or U20568 (N_20568,N_16965,N_18060);
nor U20569 (N_20569,N_18669,N_18629);
and U20570 (N_20570,N_13935,N_14472);
nor U20571 (N_20571,N_18206,N_15364);
nand U20572 (N_20572,N_14868,N_16422);
and U20573 (N_20573,N_12702,N_18560);
and U20574 (N_20574,N_13838,N_15490);
and U20575 (N_20575,N_16290,N_14050);
or U20576 (N_20576,N_18172,N_16018);
nor U20577 (N_20577,N_15638,N_13675);
and U20578 (N_20578,N_17606,N_16243);
and U20579 (N_20579,N_16788,N_12873);
and U20580 (N_20580,N_17936,N_13071);
or U20581 (N_20581,N_18215,N_17967);
or U20582 (N_20582,N_15115,N_15437);
or U20583 (N_20583,N_17108,N_13552);
and U20584 (N_20584,N_16216,N_14148);
nor U20585 (N_20585,N_12923,N_15959);
and U20586 (N_20586,N_15063,N_14582);
and U20587 (N_20587,N_14766,N_15903);
and U20588 (N_20588,N_16369,N_15695);
or U20589 (N_20589,N_12741,N_15324);
or U20590 (N_20590,N_15455,N_17496);
and U20591 (N_20591,N_18061,N_13667);
or U20592 (N_20592,N_17135,N_17520);
and U20593 (N_20593,N_18230,N_13011);
and U20594 (N_20594,N_17138,N_17712);
nand U20595 (N_20595,N_16175,N_16666);
nor U20596 (N_20596,N_17424,N_17965);
nand U20597 (N_20597,N_14872,N_15420);
and U20598 (N_20598,N_14605,N_14378);
and U20599 (N_20599,N_12762,N_17146);
and U20600 (N_20600,N_14128,N_12832);
nand U20601 (N_20601,N_16012,N_17403);
and U20602 (N_20602,N_16876,N_16392);
and U20603 (N_20603,N_16029,N_16415);
or U20604 (N_20604,N_14802,N_15079);
nand U20605 (N_20605,N_12508,N_18124);
and U20606 (N_20606,N_16413,N_17127);
and U20607 (N_20607,N_18397,N_18373);
nor U20608 (N_20608,N_17500,N_17849);
or U20609 (N_20609,N_17387,N_12546);
and U20610 (N_20610,N_15464,N_18246);
nor U20611 (N_20611,N_17566,N_16165);
and U20612 (N_20612,N_14342,N_12690);
nor U20613 (N_20613,N_17851,N_18739);
nand U20614 (N_20614,N_14292,N_13713);
nor U20615 (N_20615,N_15334,N_15900);
nor U20616 (N_20616,N_12641,N_15231);
and U20617 (N_20617,N_17982,N_14795);
or U20618 (N_20618,N_16009,N_16340);
or U20619 (N_20619,N_14613,N_14116);
nor U20620 (N_20620,N_16817,N_14138);
nor U20621 (N_20621,N_18164,N_13019);
nor U20622 (N_20622,N_15644,N_13687);
or U20623 (N_20623,N_17177,N_17952);
or U20624 (N_20624,N_16375,N_18417);
and U20625 (N_20625,N_12953,N_16445);
and U20626 (N_20626,N_16226,N_15380);
or U20627 (N_20627,N_15685,N_16657);
nand U20628 (N_20628,N_14771,N_18720);
nand U20629 (N_20629,N_18617,N_16685);
or U20630 (N_20630,N_14261,N_15678);
nand U20631 (N_20631,N_12676,N_15572);
nand U20632 (N_20632,N_14394,N_14469);
nor U20633 (N_20633,N_13751,N_15594);
nand U20634 (N_20634,N_16072,N_14548);
nand U20635 (N_20635,N_16908,N_12659);
nand U20636 (N_20636,N_16847,N_13438);
or U20637 (N_20637,N_17577,N_13492);
nand U20638 (N_20638,N_17014,N_15544);
and U20639 (N_20639,N_18224,N_15507);
nor U20640 (N_20640,N_13156,N_15882);
and U20641 (N_20641,N_14367,N_14685);
or U20642 (N_20642,N_14430,N_18504);
nor U20643 (N_20643,N_15403,N_18238);
or U20644 (N_20644,N_12766,N_13128);
nor U20645 (N_20645,N_16677,N_15167);
or U20646 (N_20646,N_17026,N_15102);
or U20647 (N_20647,N_13028,N_18734);
nor U20648 (N_20648,N_15874,N_13320);
and U20649 (N_20649,N_18501,N_17886);
or U20650 (N_20650,N_16043,N_12817);
and U20651 (N_20651,N_13152,N_12980);
nand U20652 (N_20652,N_16813,N_15110);
and U20653 (N_20653,N_16723,N_17864);
and U20654 (N_20654,N_16746,N_18545);
or U20655 (N_20655,N_17468,N_15034);
or U20656 (N_20656,N_15962,N_13245);
xor U20657 (N_20657,N_14406,N_18458);
and U20658 (N_20658,N_17124,N_18511);
nor U20659 (N_20659,N_16992,N_15999);
nand U20660 (N_20660,N_13201,N_13346);
xor U20661 (N_20661,N_16145,N_18217);
and U20662 (N_20662,N_18656,N_14439);
or U20663 (N_20663,N_16059,N_15138);
nand U20664 (N_20664,N_13778,N_14780);
and U20665 (N_20665,N_16090,N_13910);
nor U20666 (N_20666,N_17694,N_15113);
nor U20667 (N_20667,N_13463,N_16497);
or U20668 (N_20668,N_18704,N_14642);
or U20669 (N_20669,N_15550,N_17440);
nand U20670 (N_20670,N_13535,N_13586);
xor U20671 (N_20671,N_17927,N_16412);
nor U20672 (N_20672,N_15943,N_12977);
or U20673 (N_20673,N_17432,N_12532);
nor U20674 (N_20674,N_13699,N_17808);
nor U20675 (N_20675,N_14164,N_16628);
and U20676 (N_20676,N_13638,N_16917);
or U20677 (N_20677,N_17362,N_14405);
nor U20678 (N_20678,N_17221,N_18194);
and U20679 (N_20679,N_15555,N_14184);
or U20680 (N_20680,N_12698,N_16530);
or U20681 (N_20681,N_16689,N_16803);
nand U20682 (N_20682,N_16498,N_13221);
nand U20683 (N_20683,N_13429,N_17971);
nor U20684 (N_20684,N_18723,N_16650);
or U20685 (N_20685,N_15118,N_15337);
nand U20686 (N_20686,N_17082,N_17568);
and U20687 (N_20687,N_18678,N_17929);
and U20688 (N_20688,N_14061,N_14290);
and U20689 (N_20689,N_14459,N_17776);
nor U20690 (N_20690,N_13411,N_15775);
nor U20691 (N_20691,N_17595,N_18402);
or U20692 (N_20692,N_15225,N_14797);
nor U20693 (N_20693,N_14850,N_16738);
nand U20694 (N_20694,N_16888,N_17975);
nand U20695 (N_20695,N_13663,N_17597);
or U20696 (N_20696,N_16481,N_14625);
or U20697 (N_20697,N_16678,N_17823);
nor U20698 (N_20698,N_13434,N_18113);
nand U20699 (N_20699,N_14283,N_15843);
nor U20700 (N_20700,N_14778,N_17946);
nor U20701 (N_20701,N_14985,N_12852);
or U20702 (N_20702,N_14312,N_15370);
nand U20703 (N_20703,N_15152,N_17888);
nand U20704 (N_20704,N_17409,N_16940);
nand U20705 (N_20705,N_13031,N_14328);
xor U20706 (N_20706,N_13622,N_16109);
and U20707 (N_20707,N_18587,N_13857);
nor U20708 (N_20708,N_12922,N_12671);
nor U20709 (N_20709,N_18449,N_14657);
xnor U20710 (N_20710,N_15247,N_16269);
nand U20711 (N_20711,N_16368,N_14156);
nand U20712 (N_20712,N_15472,N_17066);
and U20713 (N_20713,N_16866,N_14323);
nor U20714 (N_20714,N_18598,N_13682);
and U20715 (N_20715,N_15018,N_17163);
and U20716 (N_20716,N_18546,N_17750);
or U20717 (N_20717,N_12841,N_15541);
nand U20718 (N_20718,N_17328,N_14414);
nand U20719 (N_20719,N_15885,N_18119);
or U20720 (N_20720,N_17778,N_12605);
and U20721 (N_20721,N_18371,N_17353);
nand U20722 (N_20722,N_17147,N_16688);
nand U20723 (N_20723,N_17259,N_17767);
nand U20724 (N_20724,N_18025,N_14076);
or U20725 (N_20725,N_17075,N_17546);
and U20726 (N_20726,N_17916,N_13179);
and U20727 (N_20727,N_13503,N_12771);
or U20728 (N_20728,N_14894,N_18455);
or U20729 (N_20729,N_14750,N_14426);
or U20730 (N_20730,N_13977,N_18095);
nand U20731 (N_20731,N_17389,N_17370);
nand U20732 (N_20732,N_14341,N_15770);
or U20733 (N_20733,N_15520,N_18510);
or U20734 (N_20734,N_13111,N_15250);
nor U20735 (N_20735,N_17309,N_15423);
nand U20736 (N_20736,N_16017,N_16004);
or U20737 (N_20737,N_13350,N_13409);
nand U20738 (N_20738,N_13529,N_13533);
nor U20739 (N_20739,N_14609,N_18298);
nand U20740 (N_20740,N_16964,N_15616);
nand U20741 (N_20741,N_16969,N_13059);
or U20742 (N_20742,N_18391,N_15200);
or U20743 (N_20743,N_15769,N_13936);
nand U20744 (N_20744,N_15600,N_16945);
or U20745 (N_20745,N_12662,N_15232);
nor U20746 (N_20746,N_14456,N_13918);
and U20747 (N_20747,N_16708,N_14370);
nand U20748 (N_20748,N_14209,N_17007);
and U20749 (N_20749,N_16676,N_16260);
or U20750 (N_20750,N_14655,N_14859);
or U20751 (N_20751,N_12694,N_16199);
nand U20752 (N_20752,N_18244,N_18390);
xnor U20753 (N_20753,N_15240,N_16590);
and U20754 (N_20754,N_16504,N_17735);
or U20755 (N_20755,N_18688,N_13136);
and U20756 (N_20756,N_14862,N_16262);
nand U20757 (N_20757,N_16116,N_16122);
nand U20758 (N_20758,N_18333,N_18399);
or U20759 (N_20759,N_17367,N_18497);
nand U20760 (N_20760,N_17339,N_17787);
nor U20761 (N_20761,N_13340,N_12673);
nor U20762 (N_20762,N_13372,N_17331);
and U20763 (N_20763,N_13715,N_14201);
or U20764 (N_20764,N_18713,N_14480);
and U20765 (N_20765,N_15035,N_14362);
nand U20766 (N_20766,N_17070,N_16495);
or U20767 (N_20767,N_15106,N_15669);
nand U20768 (N_20768,N_16598,N_12979);
nor U20769 (N_20769,N_12663,N_15210);
and U20770 (N_20770,N_12543,N_17995);
or U20771 (N_20771,N_17601,N_15657);
or U20772 (N_20772,N_16210,N_18411);
or U20773 (N_20773,N_15793,N_13771);
or U20774 (N_20774,N_15481,N_16823);
nor U20775 (N_20775,N_13755,N_15810);
nand U20776 (N_20776,N_17033,N_15440);
nor U20777 (N_20777,N_15161,N_15394);
nand U20778 (N_20778,N_13680,N_15159);
and U20779 (N_20779,N_17241,N_14353);
nand U20780 (N_20780,N_15445,N_14758);
nor U20781 (N_20781,N_13400,N_12726);
and U20782 (N_20782,N_16654,N_17801);
or U20783 (N_20783,N_15536,N_14499);
nand U20784 (N_20784,N_14989,N_16810);
xnor U20785 (N_20785,N_15444,N_18169);
nor U20786 (N_20786,N_18341,N_12897);
nor U20787 (N_20787,N_17890,N_17747);
nand U20788 (N_20788,N_16861,N_14169);
nand U20789 (N_20789,N_14319,N_13394);
or U20790 (N_20790,N_18344,N_17244);
nor U20791 (N_20791,N_14799,N_15245);
nand U20792 (N_20792,N_14082,N_16126);
and U20793 (N_20793,N_13787,N_15709);
or U20794 (N_20794,N_12850,N_12602);
and U20795 (N_20795,N_16049,N_12885);
and U20796 (N_20796,N_13313,N_16045);
and U20797 (N_20797,N_13034,N_18016);
and U20798 (N_20798,N_13603,N_15376);
or U20799 (N_20799,N_13199,N_13230);
nand U20800 (N_20800,N_14755,N_16844);
nand U20801 (N_20801,N_16251,N_13186);
or U20802 (N_20802,N_15329,N_12819);
nor U20803 (N_20803,N_16782,N_13370);
or U20804 (N_20804,N_16985,N_12564);
and U20805 (N_20805,N_15662,N_14881);
nor U20806 (N_20806,N_13779,N_18162);
or U20807 (N_20807,N_15465,N_13810);
or U20808 (N_20808,N_14077,N_12913);
or U20809 (N_20809,N_13651,N_17792);
nand U20810 (N_20810,N_16869,N_14540);
nand U20811 (N_20811,N_14170,N_12758);
nand U20812 (N_20812,N_14073,N_16033);
and U20813 (N_20813,N_14081,N_16586);
nor U20814 (N_20814,N_17298,N_16791);
or U20815 (N_20815,N_14043,N_14914);
nor U20816 (N_20816,N_13141,N_16028);
and U20817 (N_20817,N_14589,N_12748);
or U20818 (N_20818,N_15951,N_15855);
or U20819 (N_20819,N_15400,N_14315);
and U20820 (N_20820,N_14549,N_18092);
nand U20821 (N_20821,N_16806,N_14840);
and U20822 (N_20822,N_14360,N_13306);
or U20823 (N_20823,N_12735,N_18255);
nand U20824 (N_20824,N_16694,N_15005);
nor U20825 (N_20825,N_17461,N_15954);
nand U20826 (N_20826,N_12572,N_14124);
nand U20827 (N_20827,N_15066,N_13607);
nand U20828 (N_20828,N_17863,N_18259);
nor U20829 (N_20829,N_14558,N_14255);
nor U20830 (N_20830,N_14765,N_15871);
and U20831 (N_20831,N_17943,N_15388);
nor U20832 (N_20832,N_13701,N_13499);
nor U20833 (N_20833,N_13117,N_12693);
nand U20834 (N_20834,N_13659,N_13582);
nor U20835 (N_20835,N_12599,N_13849);
nor U20836 (N_20836,N_14964,N_14461);
and U20837 (N_20837,N_18228,N_15211);
nor U20838 (N_20838,N_13877,N_15326);
nand U20839 (N_20839,N_18527,N_16682);
nand U20840 (N_20840,N_15702,N_15383);
nor U20841 (N_20841,N_15153,N_15918);
and U20842 (N_20842,N_17871,N_14288);
nand U20843 (N_20843,N_18045,N_17969);
nand U20844 (N_20844,N_14839,N_15922);
nand U20845 (N_20845,N_17233,N_13926);
and U20846 (N_20846,N_16277,N_16863);
and U20847 (N_20847,N_16878,N_16235);
nand U20848 (N_20848,N_18321,N_17175);
nand U20849 (N_20849,N_18182,N_15875);
nor U20850 (N_20850,N_14346,N_14441);
or U20851 (N_20851,N_16767,N_16233);
and U20852 (N_20852,N_13991,N_12627);
or U20853 (N_20853,N_12878,N_15330);
and U20854 (N_20854,N_15428,N_17379);
nand U20855 (N_20855,N_18181,N_17287);
or U20856 (N_20856,N_17494,N_13843);
nand U20857 (N_20857,N_13722,N_17865);
or U20858 (N_20858,N_13225,N_16513);
nand U20859 (N_20859,N_15812,N_15304);
and U20860 (N_20860,N_18078,N_17802);
or U20861 (N_20861,N_15742,N_15411);
or U20862 (N_20862,N_17934,N_13242);
nor U20863 (N_20863,N_16561,N_15898);
nor U20864 (N_20864,N_14704,N_14022);
and U20865 (N_20865,N_17455,N_13544);
nand U20866 (N_20866,N_18008,N_16674);
nand U20867 (N_20867,N_15597,N_14980);
nor U20868 (N_20868,N_14539,N_16455);
and U20869 (N_20869,N_13853,N_12974);
or U20870 (N_20870,N_15021,N_13255);
and U20871 (N_20871,N_18529,N_15094);
or U20872 (N_20872,N_13772,N_18159);
nor U20873 (N_20873,N_15645,N_12910);
nor U20874 (N_20874,N_13214,N_16082);
or U20875 (N_20875,N_18473,N_16550);
and U20876 (N_20876,N_14954,N_18260);
and U20877 (N_20877,N_18482,N_17188);
nor U20878 (N_20878,N_16279,N_17257);
nand U20879 (N_20879,N_17196,N_16337);
nand U20880 (N_20880,N_14417,N_17162);
or U20881 (N_20881,N_14007,N_13793);
and U20882 (N_20882,N_17963,N_15877);
and U20883 (N_20883,N_17827,N_16770);
nand U20884 (N_20884,N_16656,N_13392);
nor U20885 (N_20885,N_16496,N_15057);
or U20886 (N_20886,N_17609,N_13143);
and U20887 (N_20887,N_16465,N_15814);
nand U20888 (N_20888,N_13098,N_15186);
or U20889 (N_20889,N_15461,N_18535);
nor U20890 (N_20890,N_15128,N_13647);
nand U20891 (N_20891,N_13331,N_12851);
nor U20892 (N_20892,N_13187,N_17406);
nor U20893 (N_20893,N_16086,N_16620);
or U20894 (N_20894,N_18138,N_16575);
or U20895 (N_20895,N_16836,N_13377);
nand U20896 (N_20896,N_15475,N_16545);
or U20897 (N_20897,N_16714,N_13827);
nor U20898 (N_20898,N_12982,N_13672);
or U20899 (N_20899,N_17627,N_15331);
and U20900 (N_20900,N_18616,N_17074);
or U20901 (N_20901,N_18426,N_17834);
nand U20902 (N_20902,N_16589,N_12505);
or U20903 (N_20903,N_16648,N_15914);
nand U20904 (N_20904,N_15673,N_18062);
nand U20905 (N_20905,N_16846,N_12826);
nor U20906 (N_20906,N_14135,N_16731);
nor U20907 (N_20907,N_15342,N_17185);
or U20908 (N_20908,N_18234,N_13488);
or U20909 (N_20909,N_16215,N_15679);
nand U20910 (N_20910,N_13243,N_14689);
nand U20911 (N_20911,N_16380,N_14131);
nor U20912 (N_20912,N_12757,N_15003);
nor U20913 (N_20913,N_16366,N_12941);
nor U20914 (N_20914,N_14308,N_14345);
and U20915 (N_20915,N_14427,N_13206);
nor U20916 (N_20916,N_18632,N_16129);
and U20917 (N_20917,N_14144,N_16668);
or U20918 (N_20918,N_17306,N_14398);
and U20919 (N_20919,N_12865,N_12912);
and U20920 (N_20920,N_15661,N_17420);
and U20921 (N_20921,N_16084,N_14071);
and U20922 (N_20922,N_18075,N_14252);
and U20923 (N_20923,N_13674,N_18565);
nand U20924 (N_20924,N_15977,N_18019);
and U20925 (N_20925,N_17148,N_14898);
nor U20926 (N_20926,N_18463,N_13406);
or U20927 (N_20927,N_17938,N_16304);
nand U20928 (N_20928,N_14672,N_16633);
nor U20929 (N_20929,N_14375,N_13158);
and U20930 (N_20930,N_14205,N_13270);
or U20931 (N_20931,N_13930,N_13344);
and U20932 (N_20932,N_14918,N_18178);
or U20933 (N_20933,N_15968,N_15425);
or U20934 (N_20934,N_18404,N_17454);
nor U20935 (N_20935,N_17618,N_16458);
nor U20936 (N_20936,N_12983,N_15924);
or U20937 (N_20937,N_17558,N_15691);
nor U20938 (N_20938,N_15899,N_17430);
and U20939 (N_20939,N_16259,N_17149);
nor U20940 (N_20940,N_12895,N_17071);
nor U20941 (N_20941,N_13419,N_13605);
xor U20942 (N_20942,N_15140,N_14216);
nor U20943 (N_20943,N_18366,N_13264);
and U20944 (N_20944,N_14241,N_14477);
nand U20945 (N_20945,N_12986,N_17511);
or U20946 (N_20946,N_18522,N_16146);
nor U20947 (N_20947,N_16546,N_12907);
nand U20948 (N_20948,N_14365,N_17352);
nand U20949 (N_20949,N_17552,N_17266);
or U20950 (N_20950,N_16359,N_13118);
and U20951 (N_20951,N_12651,N_16915);
nor U20952 (N_20952,N_15156,N_17283);
and U20953 (N_20953,N_18672,N_17593);
nor U20954 (N_20954,N_18108,N_15173);
nor U20955 (N_20955,N_12773,N_15892);
and U20956 (N_20956,N_17921,N_14920);
nor U20957 (N_20957,N_15226,N_12976);
nor U20958 (N_20958,N_17067,N_13789);
nor U20959 (N_20959,N_15707,N_13847);
nand U20960 (N_20960,N_16136,N_13508);
nand U20961 (N_20961,N_14683,N_13634);
or U20962 (N_20962,N_18163,N_18554);
nand U20963 (N_20963,N_15350,N_12909);
and U20964 (N_20964,N_12692,N_14653);
or U20965 (N_20965,N_16856,N_18052);
and U20966 (N_20966,N_15353,N_14843);
nand U20967 (N_20967,N_15574,N_17940);
or U20968 (N_20968,N_18407,N_17749);
or U20969 (N_20969,N_17761,N_15477);
nor U20970 (N_20970,N_13883,N_13486);
and U20971 (N_20971,N_18641,N_16318);
nand U20972 (N_20972,N_18232,N_17720);
or U20973 (N_20973,N_16872,N_15377);
nand U20974 (N_20974,N_16244,N_17850);
or U20975 (N_20975,N_17779,N_12679);
nor U20976 (N_20976,N_13309,N_13139);
nand U20977 (N_20977,N_14249,N_15139);
and U20978 (N_20978,N_17727,N_13268);
and U20979 (N_20979,N_12517,N_15547);
nand U20980 (N_20980,N_13436,N_14470);
nor U20981 (N_20981,N_14782,N_18125);
and U20982 (N_20982,N_18564,N_17628);
nor U20983 (N_20983,N_16609,N_12568);
nand U20984 (N_20984,N_18002,N_15136);
and U20985 (N_20985,N_12896,N_18385);
and U20986 (N_20986,N_12765,N_12870);
nor U20987 (N_20987,N_17955,N_16527);
and U20988 (N_20988,N_14223,N_17893);
nor U20989 (N_20989,N_18112,N_14220);
and U20990 (N_20990,N_17702,N_12727);
nor U20991 (N_20991,N_12906,N_18354);
nor U20992 (N_20992,N_13952,N_16541);
and U20993 (N_20993,N_16008,N_18087);
nand U20994 (N_20994,N_18146,N_16975);
nor U20995 (N_20995,N_15967,N_14126);
or U20996 (N_20996,N_16490,N_15374);
and U20997 (N_20997,N_13148,N_15515);
nand U20998 (N_20998,N_17281,N_15933);
nand U20999 (N_20999,N_13767,N_16566);
or U21000 (N_21000,N_17487,N_17843);
nand U21001 (N_21001,N_18711,N_16599);
nand U21002 (N_21002,N_17419,N_12855);
and U21003 (N_21003,N_17143,N_14455);
nand U21004 (N_21004,N_15671,N_14874);
or U21005 (N_21005,N_17600,N_18256);
xnor U21006 (N_21006,N_13354,N_14622);
nand U21007 (N_21007,N_17914,N_14099);
nor U21008 (N_21008,N_18106,N_15019);
nand U21009 (N_21009,N_18037,N_13907);
nor U21010 (N_21010,N_12791,N_16266);
nor U21011 (N_21011,N_17024,N_13458);
or U21012 (N_21012,N_12746,N_16133);
nor U21013 (N_21013,N_16886,N_18433);
or U21014 (N_21014,N_15612,N_15539);
nand U21015 (N_21015,N_13460,N_13673);
and U21016 (N_21016,N_12954,N_18324);
or U21017 (N_21017,N_18472,N_13585);
and U21018 (N_21018,N_15830,N_15058);
nand U21019 (N_21019,N_16560,N_15557);
and U21020 (N_21020,N_15672,N_12672);
or U21021 (N_21021,N_15298,N_14300);
nand U21022 (N_21022,N_15273,N_12889);
or U21023 (N_21023,N_16411,N_15905);
or U21024 (N_21024,N_16525,N_12661);
nor U21025 (N_21025,N_14326,N_13633);
nor U21026 (N_21026,N_15714,N_15439);
and U21027 (N_21027,N_12590,N_13993);
nand U21028 (N_21028,N_13112,N_18729);
nor U21029 (N_21029,N_15168,N_14248);
xor U21030 (N_21030,N_12624,N_17924);
and U21031 (N_21031,N_17037,N_14079);
nor U21032 (N_21032,N_17581,N_17350);
or U21033 (N_21033,N_16419,N_17302);
nand U21034 (N_21034,N_12978,N_15402);
nand U21035 (N_21035,N_14957,N_12625);
or U21036 (N_21036,N_15628,N_14660);
nor U21037 (N_21037,N_14588,N_18057);
or U21038 (N_21038,N_14177,N_14769);
nand U21039 (N_21039,N_18453,N_13418);
or U21040 (N_21040,N_12962,N_17573);
and U21041 (N_21041,N_15307,N_12798);
or U21042 (N_21042,N_16254,N_17048);
and U21043 (N_21043,N_14340,N_16400);
nand U21044 (N_21044,N_17616,N_13000);
and U21045 (N_21045,N_18240,N_17123);
and U21046 (N_21046,N_15027,N_17397);
nand U21047 (N_21047,N_15611,N_15619);
nand U21048 (N_21048,N_15393,N_16873);
or U21049 (N_21049,N_18677,N_15542);
and U21050 (N_21050,N_12777,N_15091);
nor U21051 (N_21051,N_13254,N_16100);
and U21052 (N_21052,N_17796,N_13284);
nor U21053 (N_21053,N_17002,N_17666);
or U21054 (N_21054,N_14086,N_15495);
and U21055 (N_21055,N_14863,N_18620);
or U21056 (N_21056,N_15017,N_18719);
nor U21057 (N_21057,N_13351,N_14551);
nor U21058 (N_21058,N_12928,N_17993);
nor U21059 (N_21059,N_17171,N_18076);
and U21060 (N_21060,N_17131,N_14229);
nor U21061 (N_21061,N_16735,N_17528);
and U21062 (N_21062,N_16089,N_15188);
nand U21063 (N_21063,N_14182,N_17039);
and U21064 (N_21064,N_13013,N_14040);
xor U21065 (N_21065,N_15086,N_14141);
nor U21066 (N_21066,N_18717,N_13996);
nor U21067 (N_21067,N_14286,N_17516);
nor U21068 (N_21068,N_17824,N_16786);
nand U21069 (N_21069,N_14816,N_13338);
or U21070 (N_21070,N_16222,N_18619);
and U21071 (N_21071,N_18174,N_17094);
or U21072 (N_21072,N_17232,N_13577);
and U21073 (N_21073,N_14385,N_12706);
nor U21074 (N_21074,N_18359,N_15927);
nand U21075 (N_21075,N_18701,N_14338);
and U21076 (N_21076,N_13804,N_17255);
nor U21077 (N_21077,N_17799,N_15045);
nor U21078 (N_21078,N_13448,N_16658);
nand U21079 (N_21079,N_17757,N_17278);
nor U21080 (N_21080,N_13583,N_15736);
nand U21081 (N_21081,N_12724,N_17985);
or U21082 (N_21082,N_17729,N_17644);
or U21083 (N_21083,N_15234,N_16832);
nand U21084 (N_21084,N_14594,N_16667);
nand U21085 (N_21085,N_13293,N_14279);
or U21086 (N_21086,N_18432,N_15170);
nor U21087 (N_21087,N_15237,N_18365);
and U21088 (N_21088,N_18307,N_15727);
and U21089 (N_21089,N_18151,N_14383);
or U21090 (N_21090,N_15595,N_18336);
nand U21091 (N_21091,N_13666,N_18436);
nor U21092 (N_21092,N_18187,N_15373);
nand U21093 (N_21093,N_16438,N_17297);
nand U21094 (N_21094,N_13108,N_18283);
or U21095 (N_21095,N_17962,N_12857);
nor U21096 (N_21096,N_16995,N_17327);
and U21097 (N_21097,N_14956,N_14674);
nand U21098 (N_21098,N_14191,N_18650);
or U21099 (N_21099,N_17211,N_14855);
and U21100 (N_21100,N_15392,N_13584);
nand U21101 (N_21101,N_15737,N_17891);
and U21102 (N_21102,N_15713,N_12891);
xor U21103 (N_21103,N_18679,N_15712);
or U21104 (N_21104,N_16241,N_15828);
and U21105 (N_21105,N_16245,N_17315);
nor U21106 (N_21106,N_17062,N_15258);
and U21107 (N_21107,N_13553,N_18197);
nor U21108 (N_21108,N_17760,N_12959);
or U21109 (N_21109,N_16494,N_12612);
and U21110 (N_21110,N_17134,N_18170);
and U21111 (N_21111,N_13578,N_17643);
nand U21112 (N_21112,N_16321,N_16442);
nor U21113 (N_21113,N_15761,N_14166);
nand U21114 (N_21114,N_16807,N_18072);
and U21115 (N_21115,N_17832,N_18456);
and U21116 (N_21116,N_16680,N_15041);
nor U21117 (N_21117,N_14471,N_18490);
or U21118 (N_21118,N_12550,N_13850);
nand U21119 (N_21119,N_17913,N_14528);
and U21120 (N_21120,N_17064,N_15634);
nand U21121 (N_21121,N_13356,N_16857);
nor U21122 (N_21122,N_14910,N_12804);
and U21123 (N_21123,N_13962,N_17019);
nand U21124 (N_21124,N_13595,N_18502);
nor U21125 (N_21125,N_15051,N_14692);
nand U21126 (N_21126,N_14275,N_16719);
nand U21127 (N_21127,N_16421,N_14327);
nand U21128 (N_21128,N_17486,N_13388);
nor U21129 (N_21129,N_18058,N_12519);
or U21130 (N_21130,N_13828,N_16837);
nor U21131 (N_21131,N_15715,N_15800);
or U21132 (N_21132,N_14014,N_16519);
and U21133 (N_21133,N_18267,N_17142);
nor U21134 (N_21134,N_13693,N_15749);
nor U21135 (N_21135,N_17620,N_18506);
nor U21136 (N_21136,N_12802,N_15111);
and U21137 (N_21137,N_15012,N_14987);
nand U21138 (N_21138,N_13656,N_16910);
nor U21139 (N_21139,N_17514,N_14896);
nand U21140 (N_21140,N_18279,N_17701);
nand U21141 (N_21141,N_15725,N_17598);
nand U21142 (N_21142,N_18340,N_18120);
nand U21143 (N_21143,N_16838,N_15687);
nand U21144 (N_21144,N_18605,N_14936);
nor U21145 (N_21145,N_14298,N_12848);
and U21146 (N_21146,N_17443,N_13445);
and U21147 (N_21147,N_17845,N_18210);
nor U21148 (N_21148,N_18392,N_17317);
nor U21149 (N_21149,N_13441,N_12513);
and U21150 (N_21150,N_14293,N_16858);
or U21151 (N_21151,N_16855,N_14908);
nor U21152 (N_21152,N_15151,N_17672);
nor U21153 (N_21153,N_13968,N_12931);
or U21154 (N_21154,N_16512,N_15119);
nand U21155 (N_21155,N_13253,N_16581);
nor U21156 (N_21156,N_17676,N_16864);
nor U21157 (N_21157,N_16884,N_18613);
and U21158 (N_21158,N_12593,N_17768);
nand U21159 (N_21159,N_16177,N_13515);
nand U21160 (N_21160,N_15300,N_15093);
nor U21161 (N_21161,N_15526,N_15485);
and U21162 (N_21162,N_14443,N_14641);
nand U21163 (N_21163,N_18105,N_15842);
and U21164 (N_21164,N_15416,N_16094);
nand U21165 (N_21165,N_14388,N_15841);
or U21166 (N_21166,N_14604,N_14305);
nor U21167 (N_21167,N_14735,N_13600);
nor U21168 (N_21168,N_14927,N_16901);
and U21169 (N_21169,N_17980,N_17261);
nand U21170 (N_21170,N_18465,N_17602);
or U21171 (N_21171,N_18276,N_15950);
nand U21172 (N_21172,N_13916,N_17206);
and U21173 (N_21173,N_17821,N_16626);
nand U21174 (N_21174,N_14993,N_15620);
nor U21175 (N_21175,N_18746,N_15145);
nor U21176 (N_21176,N_13729,N_17400);
and U21177 (N_21177,N_14794,N_16383);
nor U21178 (N_21178,N_16880,N_13965);
nand U21179 (N_21179,N_15837,N_15294);
nand U21180 (N_21180,N_13020,N_17422);
nor U21181 (N_21181,N_14085,N_16013);
or U21182 (N_21182,N_17395,N_18375);
or U21183 (N_21183,N_16764,N_17354);
nor U21184 (N_21184,N_17386,N_13181);
nand U21185 (N_21185,N_14101,N_17794);
nand U21186 (N_21186,N_14676,N_16584);
nor U21187 (N_21187,N_13532,N_12551);
xor U21188 (N_21188,N_12720,N_16261);
or U21189 (N_21189,N_18289,N_16424);
nor U21190 (N_21190,N_14621,N_13959);
nor U21191 (N_21191,N_15013,N_13232);
and U21192 (N_21192,N_15431,N_16316);
nor U21193 (N_21193,N_16702,N_15847);
nand U21194 (N_21194,N_13869,N_15680);
and U21195 (N_21195,N_12751,N_14749);
or U21196 (N_21196,N_13612,N_18049);
and U21197 (N_21197,N_16078,N_13390);
or U21198 (N_21198,N_12634,N_17250);
and U21199 (N_21199,N_14860,N_16355);
and U21200 (N_21200,N_13620,N_13440);
or U21201 (N_21201,N_16230,N_13617);
nor U21202 (N_21202,N_18314,N_13277);
or U21203 (N_21203,N_15333,N_18379);
nor U21204 (N_21204,N_14572,N_16994);
and U21205 (N_21205,N_14517,N_12697);
nand U21206 (N_21206,N_15681,N_14272);
nor U21207 (N_21207,N_14720,N_15382);
and U21208 (N_21208,N_14975,N_16679);
nor U21209 (N_21209,N_17286,N_13716);
or U21210 (N_21210,N_14535,N_17968);
or U21211 (N_21211,N_13425,N_13076);
and U21212 (N_21212,N_15459,N_13707);
and U21213 (N_21213,N_12501,N_12642);
and U21214 (N_21214,N_15670,N_16748);
nor U21215 (N_21215,N_14707,N_13178);
nand U21216 (N_21216,N_13575,N_15919);
nand U21217 (N_21217,N_15412,N_12840);
or U21218 (N_21218,N_14110,N_15281);
or U21219 (N_21219,N_15760,N_15414);
and U21220 (N_21220,N_13375,N_18671);
nor U21221 (N_21221,N_15254,N_17133);
nor U21222 (N_21222,N_18208,N_15831);
nor U21223 (N_21223,N_16183,N_17252);
nand U21224 (N_21224,N_18654,N_16054);
nor U21225 (N_21225,N_13316,N_16113);
or U21226 (N_21226,N_13978,N_14646);
nor U21227 (N_21227,N_16308,N_15457);
nand U21228 (N_21228,N_14422,N_14603);
or U21229 (N_21229,N_12524,N_16606);
or U21230 (N_21230,N_15636,N_13322);
nor U21231 (N_21231,N_18444,N_12768);
nor U21232 (N_21232,N_15137,N_13964);
nor U21233 (N_21233,N_13886,N_12657);
or U21234 (N_21234,N_17782,N_15756);
or U21235 (N_21235,N_17976,N_13660);
nand U21236 (N_21236,N_18063,N_15025);
nor U21237 (N_21237,N_16771,N_16730);
nor U21238 (N_21238,N_15677,N_16905);
and U21239 (N_21239,N_17697,N_16057);
nor U21240 (N_21240,N_18396,N_14278);
nand U21241 (N_21241,N_12531,N_14449);
xnor U21242 (N_21242,N_13408,N_16335);
or U21243 (N_21243,N_14633,N_12812);
nand U21244 (N_21244,N_17926,N_17703);
nor U21245 (N_21245,N_13739,N_18117);
nand U21246 (N_21246,N_16444,N_14564);
nor U21247 (N_21247,N_16231,N_16181);
and U21248 (N_21248,N_13087,N_14885);
nor U21249 (N_21249,N_16716,N_17376);
nand U21250 (N_21250,N_16385,N_16390);
or U21251 (N_21251,N_18171,N_15663);
or U21252 (N_21252,N_18074,N_13924);
nand U21253 (N_21253,N_14123,N_14607);
and U21254 (N_21254,N_13167,N_13686);
nand U21255 (N_21255,N_13437,N_13654);
nor U21256 (N_21256,N_13939,N_17847);
nor U21257 (N_21257,N_17684,N_13376);
or U21258 (N_21258,N_12987,N_17882);
nand U21259 (N_21259,N_15553,N_15101);
nor U21260 (N_21260,N_18462,N_12794);
nor U21261 (N_21261,N_13424,N_13635);
nand U21262 (N_21262,N_14858,N_15623);
and U21263 (N_21263,N_15552,N_14059);
nor U21264 (N_21264,N_18331,N_15160);
or U21265 (N_21265,N_14966,N_16932);
nor U21266 (N_21266,N_17251,N_16946);
nand U21267 (N_21267,N_14400,N_15410);
and U21268 (N_21268,N_13134,N_18305);
nor U21269 (N_21269,N_17102,N_15484);
or U21270 (N_21270,N_13664,N_14654);
nor U21271 (N_21271,N_15205,N_13235);
nor U21272 (N_21272,N_12998,N_15735);
and U21273 (N_21273,N_16683,N_17713);
and U21274 (N_21274,N_16565,N_12831);
or U21275 (N_21275,N_16608,N_17205);
or U21276 (N_21276,N_14522,N_14883);
nor U21277 (N_21277,N_16239,N_16802);
nor U21278 (N_21278,N_13597,N_12579);
nor U21279 (N_21279,N_14013,N_12946);
nor U21280 (N_21280,N_13542,N_16020);
nand U21281 (N_21281,N_16537,N_17200);
and U21282 (N_21282,N_17464,N_13462);
nor U21283 (N_21283,N_17031,N_13260);
or U21284 (N_21284,N_12648,N_15469);
nor U21285 (N_21285,N_16402,N_15617);
or U21286 (N_21286,N_17267,N_18601);
nand U21287 (N_21287,N_16168,N_16781);
and U21288 (N_21288,N_14494,N_15889);
nand U21289 (N_21289,N_14167,N_15523);
nand U21290 (N_21290,N_12844,N_15492);
nor U21291 (N_21291,N_16190,N_16255);
and U21292 (N_21292,N_12745,N_14092);
nand U21293 (N_21293,N_14320,N_16037);
or U21294 (N_21294,N_17418,N_16562);
nand U21295 (N_21295,N_14401,N_16920);
and U21296 (N_21296,N_14197,N_17611);
and U21297 (N_21297,N_16077,N_17986);
nand U21298 (N_21298,N_16460,N_14995);
nor U21299 (N_21299,N_17930,N_14011);
and U21300 (N_21300,N_13527,N_14121);
nor U21301 (N_21301,N_14351,N_14057);
or U21302 (N_21302,N_18066,N_17343);
nand U21303 (N_21303,N_18450,N_15504);
nor U21304 (N_21304,N_12738,N_17247);
or U21305 (N_21305,N_13173,N_14719);
nor U21306 (N_21306,N_15920,N_14912);
and U21307 (N_21307,N_16159,N_13146);
nor U21308 (N_21308,N_17340,N_14990);
nand U21309 (N_21309,N_17029,N_12709);
or U21310 (N_21310,N_14900,N_15816);
and U21311 (N_21311,N_12805,N_13177);
nand U21312 (N_21312,N_16356,N_15935);
or U21313 (N_21313,N_13706,N_13036);
nand U21314 (N_21314,N_15369,N_18353);
nand U21315 (N_21315,N_12595,N_14049);
nor U21316 (N_21316,N_16670,N_15339);
nor U21317 (N_21317,N_18167,N_17363);
nor U21318 (N_21318,N_13526,N_17428);
nor U21319 (N_21319,N_15849,N_15201);
or U21320 (N_21320,N_17384,N_17054);
and U21321 (N_21321,N_14824,N_17112);
nand U21322 (N_21322,N_14491,N_17151);
and U21323 (N_21323,N_13972,N_15175);
nand U21324 (N_21324,N_16643,N_13834);
and U21325 (N_21325,N_14206,N_18225);
nor U21326 (N_21326,N_13319,N_17718);
and U21327 (N_21327,N_18154,N_18190);
nor U21328 (N_21328,N_18115,N_17675);
or U21329 (N_21329,N_18319,N_12932);
nor U21330 (N_21330,N_15251,N_12689);
and U21331 (N_21331,N_17230,N_13743);
nor U21332 (N_21332,N_18721,N_17225);
and U21333 (N_21333,N_13233,N_16822);
or U21334 (N_21334,N_18706,N_12506);
and U21335 (N_21335,N_13504,N_14530);
nor U21336 (N_21336,N_13090,N_18608);
nor U21337 (N_21337,N_18749,N_15192);
nor U21338 (N_21338,N_12769,N_15778);
or U21339 (N_21339,N_17508,N_12623);
or U21340 (N_21340,N_15448,N_14532);
and U21341 (N_21341,N_12991,N_16449);
and U21342 (N_21342,N_14366,N_15980);
and U21343 (N_21343,N_16596,N_13342);
nand U21344 (N_21344,N_15470,N_15844);
nor U21345 (N_21345,N_16580,N_18454);
xor U21346 (N_21346,N_17804,N_15430);
nor U21347 (N_21347,N_14458,N_16750);
nor U21348 (N_21348,N_17459,N_15618);
nand U21349 (N_21349,N_13041,N_16968);
nor U21350 (N_21350,N_13694,N_14991);
nand U21351 (N_21351,N_18536,N_12774);
and U21352 (N_21352,N_18460,N_15789);
or U21353 (N_21353,N_13105,N_17973);
and U21354 (N_21354,N_13614,N_18144);
nand U21355 (N_21355,N_12882,N_12845);
nand U21356 (N_21356,N_15799,N_18237);
nor U21357 (N_21357,N_15993,N_13054);
nor U21358 (N_21358,N_18258,N_18236);
nand U21359 (N_21359,N_17580,N_16286);
nand U21360 (N_21360,N_17043,N_16370);
and U21361 (N_21361,N_18356,N_17788);
nand U21362 (N_21362,N_17959,N_17156);
and U21363 (N_21363,N_18738,N_15257);
nand U21364 (N_21364,N_17942,N_13570);
nor U21365 (N_21365,N_16272,N_12684);
nor U21366 (N_21366,N_18623,N_17922);
or U21367 (N_21367,N_16435,N_14518);
or U21368 (N_21368,N_16088,N_14188);
and U21369 (N_21369,N_14168,N_13182);
nand U21370 (N_21370,N_13328,N_12721);
or U21371 (N_21371,N_14907,N_18423);
nor U21372 (N_21372,N_15564,N_17481);
or U21373 (N_21373,N_13594,N_15940);
and U21374 (N_21374,N_14157,N_14492);
or U21375 (N_21375,N_13446,N_18409);
or U21376 (N_21376,N_16651,N_13929);
and U21377 (N_21377,N_16350,N_15142);
nand U21378 (N_21378,N_18268,N_18218);
or U21379 (N_21379,N_15122,N_18631);
nand U21380 (N_21380,N_13048,N_14273);
nor U21381 (N_21381,N_13914,N_17780);
nor U21382 (N_21382,N_16709,N_17166);
and U21383 (N_21383,N_16959,N_13941);
and U21384 (N_21384,N_15024,N_16698);
and U21385 (N_21385,N_14651,N_17945);
nand U21386 (N_21386,N_14950,N_16795);
nand U21387 (N_21387,N_17235,N_18126);
or U21388 (N_21388,N_13366,N_14111);
nor U21389 (N_21389,N_18009,N_16635);
and U21390 (N_21390,N_16041,N_16164);
nand U21391 (N_21391,N_17113,N_16281);
nand U21392 (N_21392,N_12629,N_17262);
and U21393 (N_21393,N_13431,N_17680);
nand U21394 (N_21394,N_15103,N_13203);
and U21395 (N_21395,N_15563,N_13396);
nor U21396 (N_21396,N_16595,N_15407);
nor U21397 (N_21397,N_13995,N_14512);
and U21398 (N_21398,N_12654,N_18388);
nor U21399 (N_21399,N_12742,N_13369);
and U21400 (N_21400,N_18633,N_12864);
and U21401 (N_21401,N_13975,N_16294);
nor U21402 (N_21402,N_16690,N_18516);
nand U21403 (N_21403,N_13386,N_18282);
nor U21404 (N_21404,N_16205,N_16811);
and U21405 (N_21405,N_15804,N_17797);
or U21406 (N_21406,N_12552,N_13046);
nor U21407 (N_21407,N_15384,N_18742);
and U21408 (N_21408,N_18369,N_14856);
or U21409 (N_21409,N_16167,N_16852);
nor U21410 (N_21410,N_13623,N_14561);
nand U21411 (N_21411,N_16692,N_17596);
nand U21412 (N_21412,N_16874,N_13164);
nor U21413 (N_21413,N_16432,N_14829);
nor U21414 (N_21414,N_13153,N_15047);
or U21415 (N_21415,N_17937,N_18652);
or U21416 (N_21416,N_13068,N_13352);
or U21417 (N_21417,N_15335,N_16030);
or U21418 (N_21418,N_13207,N_13897);
nand U21419 (N_21419,N_15880,N_13661);
nor U21420 (N_21420,N_15643,N_16485);
nor U21421 (N_21421,N_14992,N_16907);
nor U21422 (N_21422,N_16021,N_12808);
or U21423 (N_21423,N_18700,N_16258);
and U21424 (N_21424,N_13610,N_14800);
nand U21425 (N_21425,N_18342,N_14945);
nor U21426 (N_21426,N_15780,N_14946);
nand U21427 (N_21427,N_13451,N_17209);
nand U21428 (N_21428,N_12883,N_17264);
or U21429 (N_21429,N_14792,N_14376);
and U21430 (N_21430,N_15171,N_14041);
nor U21431 (N_21431,N_13758,N_16971);
nor U21432 (N_21432,N_17122,N_16710);
and U21433 (N_21433,N_16441,N_17504);
and U21434 (N_21434,N_18558,N_13444);
or U21435 (N_21435,N_14713,N_13110);
nor U21436 (N_21436,N_16773,N_15482);
nand U21437 (N_21437,N_16775,N_15772);
nand U21438 (N_21438,N_17978,N_13459);
nand U21439 (N_21439,N_13790,N_16755);
and U21440 (N_21440,N_13639,N_16103);
nand U21441 (N_21441,N_13349,N_14457);
and U21442 (N_21442,N_17722,N_17057);
or U21443 (N_21443,N_17140,N_15149);
nand U21444 (N_21444,N_14029,N_15806);
or U21445 (N_21445,N_15745,N_15508);
nand U21446 (N_21446,N_18272,N_17509);
and U21447 (N_21447,N_18630,N_15308);
or U21448 (N_21448,N_15795,N_17578);
or U21449 (N_21449,N_17448,N_16461);
nor U21450 (N_21450,N_16729,N_15123);
or U21451 (N_21451,N_17192,N_16186);
nor U21452 (N_21452,N_16765,N_13339);
or U21453 (N_21453,N_13761,N_16105);
and U21454 (N_21454,N_15117,N_14419);
nor U21455 (N_21455,N_16503,N_17860);
nand U21456 (N_21456,N_14213,N_14055);
nor U21457 (N_21457,N_14943,N_17582);
nand U21458 (N_21458,N_13149,N_15065);
or U21459 (N_21459,N_12790,N_17654);
or U21460 (N_21460,N_18381,N_18376);
or U21461 (N_21461,N_18655,N_16143);
nor U21462 (N_21462,N_15963,N_16828);
nand U21463 (N_21463,N_17556,N_17407);
and U21464 (N_21464,N_14105,N_16640);
or U21465 (N_21465,N_17857,N_12764);
and U21466 (N_21466,N_13728,N_16463);
and U21467 (N_21467,N_15450,N_15545);
nor U21468 (N_21468,N_16649,N_14580);
nand U21469 (N_21469,N_16119,N_17207);
or U21470 (N_21470,N_18226,N_18180);
nand U21471 (N_21471,N_13452,N_16867);
nor U21472 (N_21472,N_17956,N_12565);
nand U21473 (N_21473,N_15605,N_16997);
nand U21474 (N_21474,N_17510,N_13626);
and U21475 (N_21475,N_17081,N_14667);
or U21476 (N_21476,N_16270,N_14638);
nand U21477 (N_21477,N_16060,N_16055);
nand U21478 (N_21478,N_17311,N_15081);
or U21479 (N_21479,N_14846,N_14238);
nor U21480 (N_21480,N_13061,N_15724);
nor U21481 (N_21481,N_16414,N_16156);
nand U21482 (N_21482,N_13591,N_15246);
nand U21483 (N_21483,N_17769,N_13129);
nor U21484 (N_21484,N_14174,N_14258);
and U21485 (N_21485,N_13314,N_17375);
nand U21486 (N_21486,N_17263,N_15193);
nand U21487 (N_21487,N_12807,N_15991);
and U21488 (N_21488,N_14553,N_13865);
or U21489 (N_21489,N_18326,N_15503);
nor U21490 (N_21490,N_18183,N_12782);
nand U21491 (N_21491,N_16140,N_18466);
or U21492 (N_21492,N_12950,N_14784);
nor U21493 (N_21493,N_15163,N_12561);
nand U21494 (N_21494,N_16641,N_14246);
and U21495 (N_21495,N_15317,N_15442);
and U21496 (N_21496,N_14977,N_13906);
and U21497 (N_21497,N_17815,N_17648);
nand U21498 (N_21498,N_12645,N_17811);
nor U21499 (N_21499,N_13047,N_12655);
and U21500 (N_21500,N_15279,N_14172);
and U21501 (N_21501,N_17414,N_16297);
and U21502 (N_21502,N_18185,N_17478);
and U21503 (N_21503,N_13768,N_14496);
or U21504 (N_21504,N_15029,N_18137);
nor U21505 (N_21505,N_13590,N_15583);
nor U21506 (N_21506,N_17714,N_18368);
nor U21507 (N_21507,N_15947,N_16727);
and U21508 (N_21508,N_18099,N_16373);
nand U21509 (N_21509,N_17408,N_18147);
or U21510 (N_21510,N_17479,N_16961);
or U21511 (N_21511,N_14120,N_17318);
and U21512 (N_21512,N_16933,N_18649);
nand U21513 (N_21513,N_15955,N_13655);
nor U21514 (N_21514,N_14556,N_18084);
and U21515 (N_21515,N_16639,N_14611);
or U21516 (N_21516,N_17092,N_12617);
and U21517 (N_21517,N_12964,N_15676);
and U21518 (N_21518,N_17661,N_13465);
nand U21519 (N_21519,N_14597,N_17042);
nand U21520 (N_21520,N_17044,N_18297);
nor U21521 (N_21521,N_13193,N_17068);
nand U21522 (N_21522,N_16646,N_18722);
or U21523 (N_21523,N_14935,N_16914);
or U21524 (N_21524,N_13417,N_16163);
nand U21525 (N_21525,N_15958,N_16062);
and U21526 (N_21526,N_16925,N_16313);
nor U21527 (N_21527,N_14257,N_12637);
nor U21528 (N_21528,N_17321,N_17477);
nor U21529 (N_21529,N_17855,N_15867);
and U21530 (N_21530,N_14452,N_15356);
or U21531 (N_21531,N_14025,N_16706);
nor U21532 (N_21532,N_18039,N_14218);
or U21533 (N_21533,N_18413,N_15227);
nand U21534 (N_21534,N_15284,N_13144);
and U21535 (N_21535,N_14259,N_16192);
nor U21536 (N_21536,N_18349,N_13948);
nand U21537 (N_21537,N_15221,N_13359);
or U21538 (N_21538,N_14678,N_14074);
and U21539 (N_21539,N_15462,N_15064);
nand U21540 (N_21540,N_14662,N_14557);
nand U21541 (N_21541,N_13114,N_18730);
or U21542 (N_21542,N_15917,N_13704);
and U21543 (N_21543,N_17649,N_15860);
or U21544 (N_21544,N_13822,N_12580);
nor U21545 (N_21545,N_17469,N_16134);
xnor U21546 (N_21546,N_15580,N_18370);
and U21547 (N_21547,N_13055,N_18663);
nand U21548 (N_21548,N_15861,N_14801);
nor U21549 (N_21549,N_18570,N_13986);
or U21550 (N_21550,N_13248,N_12664);
and U21551 (N_21551,N_15088,N_17434);
or U21552 (N_21552,N_13258,N_18589);
nand U21553 (N_21553,N_14892,N_15274);
nor U21554 (N_21554,N_18257,N_17365);
nor U21555 (N_21555,N_16510,N_12696);
or U21556 (N_21556,N_16769,N_15752);
nor U21557 (N_21557,N_12989,N_16752);
or U21558 (N_21558,N_15964,N_16317);
nand U21559 (N_21559,N_16843,N_17273);
and U21560 (N_21560,N_13238,N_17269);
and U21561 (N_21561,N_14190,N_15395);
nor U21562 (N_21562,N_15666,N_18528);
nor U21563 (N_21563,N_15506,N_17657);
and U21564 (N_21564,N_17489,N_17035);
and U21565 (N_21565,N_18657,N_13958);
nand U21566 (N_21566,N_17447,N_15302);
nor U21567 (N_21567,N_16194,N_12677);
nor U21568 (N_21568,N_14460,N_18582);
nand U21569 (N_21569,N_16787,N_16289);
nor U21570 (N_21570,N_13251,N_16247);
nand U21571 (N_21571,N_15994,N_15413);
nand U21572 (N_21572,N_18046,N_12592);
nand U21573 (N_21573,N_17670,N_18615);
nor U21574 (N_21574,N_14152,N_18398);
nand U21575 (N_21575,N_14067,N_15740);
or U21576 (N_21576,N_15244,N_14154);
nand U21577 (N_21577,N_13063,N_12518);
or U21578 (N_21578,N_13876,N_16996);
nor U21579 (N_21579,N_14864,N_17765);
nand U21580 (N_21580,N_18339,N_16429);
or U21581 (N_21581,N_12718,N_13904);
or U21582 (N_21582,N_14836,N_17425);
nor U21583 (N_21583,N_16868,N_14587);
or U21584 (N_21584,N_17858,N_14694);
nor U21585 (N_21585,N_12560,N_16353);
or U21586 (N_21586,N_16394,N_12810);
or U21587 (N_21587,N_12646,N_15233);
nor U21588 (N_21588,N_12581,N_18263);
or U21589 (N_21589,N_14321,N_14827);
nor U21590 (N_21590,N_13683,N_14003);
or U21591 (N_21591,N_18275,N_14325);
or U21592 (N_21592,N_15610,N_12780);
or U21593 (N_21593,N_12753,N_18030);
nand U21594 (N_21594,N_17710,N_13171);
and U21595 (N_21595,N_15190,N_14866);
or U21596 (N_21596,N_14903,N_18088);
nor U21597 (N_21597,N_15953,N_17004);
nor U21598 (N_21598,N_17660,N_17563);
and U21599 (N_21599,N_12793,N_16673);
nor U21600 (N_21600,N_16923,N_16663);
or U21601 (N_21601,N_16451,N_14411);
or U21602 (N_21602,N_15451,N_13616);
nand U21603 (N_21603,N_17316,N_18586);
nand U21604 (N_21604,N_13208,N_16474);
or U21605 (N_21605,N_12759,N_17717);
nand U21606 (N_21606,N_15883,N_15049);
and U21607 (N_21607,N_13611,N_12682);
nand U21608 (N_21608,N_14593,N_16025);
or U21609 (N_21609,N_13860,N_15467);
or U21610 (N_21610,N_12904,N_14147);
and U21611 (N_21611,N_15478,N_17300);
or U21612 (N_21612,N_18395,N_16050);
or U21613 (N_21613,N_12687,N_13776);
nand U21614 (N_21614,N_12949,N_16479);
or U21615 (N_21615,N_16339,N_17831);
nand U21616 (N_21616,N_16587,N_18229);
and U21617 (N_21617,N_15901,N_14844);
and U21618 (N_21618,N_18443,N_15577);
nor U21619 (N_21619,N_15039,N_18003);
or U21620 (N_21620,N_16275,N_16467);
or U21621 (N_21621,N_13966,N_16592);
nor U21622 (N_21622,N_15135,N_14268);
and U21623 (N_21623,N_13856,N_16106);
and U21624 (N_21624,N_17216,N_15518);
or U21625 (N_21625,N_14818,N_15596);
and U21626 (N_21626,N_15345,N_16448);
nor U21627 (N_21627,N_14796,N_13908);
nor U21628 (N_21628,N_16845,N_14786);
and U21629 (N_21629,N_17498,N_18576);
nand U21630 (N_21630,N_15878,N_16470);
or U21631 (N_21631,N_18107,N_15236);
nor U21632 (N_21632,N_14902,N_18134);
or U21633 (N_21633,N_13744,N_13003);
or U21634 (N_21634,N_12824,N_15730);
nand U21635 (N_21635,N_13291,N_12507);
nor U21636 (N_21636,N_15054,N_13837);
nor U21637 (N_21637,N_16309,N_14236);
or U21638 (N_21638,N_13983,N_14431);
nand U21639 (N_21639,N_16734,N_17164);
nand U21640 (N_21640,N_15426,N_18241);
or U21641 (N_21641,N_13487,N_15528);
nand U21642 (N_21642,N_16988,N_17518);
nor U21643 (N_21643,N_12822,N_12639);
nand U21644 (N_21644,N_16307,N_17783);
nor U21645 (N_21645,N_16360,N_13115);
or U21646 (N_21646,N_18653,N_13478);
nand U21647 (N_21647,N_18531,N_13501);
nor U21648 (N_21648,N_16315,N_13811);
or U21649 (N_21649,N_16409,N_17699);
or U21650 (N_21650,N_15562,N_18231);
or U21651 (N_21651,N_13348,N_15422);
nor U21652 (N_21652,N_14194,N_13464);
and U21653 (N_21653,N_15038,N_18464);
or U21654 (N_21654,N_14240,N_16293);
nand U21655 (N_21655,N_15050,N_18007);
or U21656 (N_21656,N_13086,N_14161);
nand U21657 (N_21657,N_17091,N_13443);
and U21658 (N_21658,N_17651,N_17870);
nand U21659 (N_21659,N_16107,N_13830);
nand U21660 (N_21660,N_17635,N_14552);
nor U21661 (N_21661,N_18442,N_15538);
or U21662 (N_21662,N_16523,N_14080);
and U21663 (N_21663,N_16189,N_13724);
nand U21664 (N_21664,N_15614,N_17165);
or U21665 (N_21665,N_13387,N_18557);
nand U21666 (N_21666,N_17079,N_14250);
nor U21667 (N_21667,N_15087,N_15650);
and U21668 (N_21668,N_13774,N_13609);
and U21669 (N_21669,N_16464,N_13135);
nor U21670 (N_21670,N_17641,N_18745);
nand U21671 (N_21671,N_14222,N_15609);
xnor U21672 (N_21672,N_17734,N_18378);
and U21673 (N_21673,N_17719,N_18328);
or U21674 (N_21674,N_13014,N_13226);
and U21675 (N_21675,N_15323,N_17538);
nor U21676 (N_21676,N_15028,N_14440);
and U21677 (N_21677,N_18048,N_14028);
nand U21678 (N_21678,N_14122,N_15452);
or U21679 (N_21679,N_14665,N_16916);
nor U21680 (N_21680,N_15074,N_17421);
nand U21681 (N_21681,N_13453,N_18600);
and U21682 (N_21682,N_17083,N_15913);
nand U21683 (N_21683,N_14825,N_17248);
nor U21684 (N_21684,N_12704,N_16466);
and U21685 (N_21685,N_12591,N_16431);
or U21686 (N_21686,N_18014,N_14804);
nor U21687 (N_21687,N_13602,N_16139);
and U21688 (N_21688,N_14616,N_14545);
or U21689 (N_21689,N_16298,N_16264);
nand U21690 (N_21690,N_14137,N_12843);
nand U21691 (N_21691,N_17919,N_15228);
nor U21692 (N_21692,N_12699,N_13569);
and U21693 (N_21693,N_12714,N_13378);
nor U21694 (N_21694,N_13312,N_18612);
nor U21695 (N_21695,N_13982,N_13967);
or U21696 (N_21696,N_16662,N_14675);
nand U21697 (N_21697,N_14052,N_14577);
and U21698 (N_21698,N_12920,N_13026);
and U21699 (N_21699,N_13592,N_18033);
nor U21700 (N_21700,N_13426,N_15635);
and U21701 (N_21701,N_18303,N_16825);
nand U21702 (N_21702,N_14592,N_13477);
nand U21703 (N_21703,N_13198,N_16549);
nand U21704 (N_21704,N_16665,N_14409);
nor U21705 (N_21705,N_18674,N_12541);
nor U21706 (N_21706,N_13670,N_16600);
or U21707 (N_21707,N_13796,N_15277);
and U21708 (N_21708,N_13106,N_17817);
nor U21709 (N_21709,N_16162,N_16322);
nor U21710 (N_21710,N_18514,N_18540);
or U21711 (N_21711,N_18547,N_18175);
or U21712 (N_21712,N_15808,N_16909);
or U21713 (N_21713,N_15728,N_12725);
nand U21714 (N_21714,N_13484,N_13579);
xnor U21715 (N_21715,N_17136,N_13304);
and U21716 (N_21716,N_15960,N_13223);
nor U21717 (N_21717,N_17374,N_16533);
or U21718 (N_21718,N_16420,N_14709);
and U21719 (N_21719,N_18018,N_18327);
or U21720 (N_21720,N_16326,N_13170);
nor U21721 (N_21721,N_13769,N_18550);
or U21722 (N_21722,N_15314,N_12650);
nor U21723 (N_21723,N_12973,N_16487);
or U21724 (N_21724,N_13885,N_13587);
and U21725 (N_21725,N_14725,N_15665);
and U21726 (N_21726,N_15651,N_13075);
and U21727 (N_21727,N_18666,N_16034);
or U21728 (N_21728,N_14798,N_17742);
nand U21729 (N_21729,N_13671,N_18299);
or U21730 (N_21730,N_12585,N_13516);
or U21731 (N_21731,N_17388,N_14955);
nor U21732 (N_21732,N_12728,N_15615);
xnor U21733 (N_21733,N_15653,N_13329);
nand U21734 (N_21734,N_12981,N_12786);
or U21735 (N_21735,N_14087,N_16929);
nor U21736 (N_21736,N_17268,N_12719);
nand U21737 (N_21737,N_14615,N_13836);
and U21738 (N_21738,N_15858,N_18405);
or U21739 (N_21739,N_17723,N_17668);
nand U21740 (N_21740,N_13643,N_16978);
and U21741 (N_21741,N_13470,N_14848);
or U21742 (N_21742,N_14373,N_13455);
nor U21743 (N_21743,N_15815,N_13095);
xnor U21744 (N_21744,N_14284,N_18635);
or U21745 (N_21745,N_16555,N_17295);
nand U21746 (N_21746,N_17069,N_13752);
nor U21747 (N_21747,N_17756,N_13056);
and U21748 (N_21748,N_14514,N_13538);
and U21749 (N_21749,N_15888,N_14333);
nand U21750 (N_21750,N_16718,N_12614);
nand U21751 (N_21751,N_13039,N_14193);
or U21752 (N_21752,N_17707,N_14763);
nor U21753 (N_21753,N_12688,N_16476);
nand U21754 (N_21754,N_14576,N_16114);
nor U21755 (N_21755,N_18676,N_17545);
nand U21756 (N_21756,N_17346,N_16124);
and U21757 (N_21757,N_18592,N_16179);
nor U21758 (N_21758,N_13824,N_17879);
or U21759 (N_21759,N_17155,N_13695);
and U21760 (N_21760,N_18358,N_18716);
nand U21761 (N_21761,N_16742,N_12936);
or U21762 (N_21762,N_13454,N_14841);
or U21763 (N_21763,N_18290,N_17308);
nor U21764 (N_21764,N_15757,N_12566);
nand U21765 (N_21765,N_12806,N_18519);
nor U21766 (N_21766,N_18064,N_17698);
nor U21767 (N_21767,N_18451,N_13358);
nor U21768 (N_21768,N_18350,N_17011);
and U21769 (N_21769,N_17465,N_16130);
or U21770 (N_21770,N_18346,N_15002);
or U21771 (N_21771,N_14107,N_12788);
or U21772 (N_21772,N_13273,N_13481);
nor U21773 (N_21773,N_17022,N_14632);
nand U21774 (N_21774,N_15037,N_17078);
or U21775 (N_21775,N_14256,N_13894);
or U21776 (N_21776,N_15315,N_12537);
nand U21777 (N_21777,N_15357,N_17820);
and U21778 (N_21778,N_17034,N_14039);
and U21779 (N_21779,N_14114,N_18439);
nor U21780 (N_21780,N_16582,N_14173);
nand U21781 (N_21781,N_14065,N_13283);
or U21782 (N_21782,N_14901,N_16201);
or U21783 (N_21783,N_13864,N_15809);
and U21784 (N_21784,N_15664,N_16563);
and U21785 (N_21785,N_17254,N_16052);
nor U21786 (N_21786,N_17492,N_15592);
or U21787 (N_21787,N_17861,N_12797);
or U21788 (N_21788,N_18203,N_18607);
and U21789 (N_21789,N_17359,N_18628);
and U21790 (N_21790,N_15266,N_17948);
nand U21791 (N_21791,N_14696,N_13549);
nand U21792 (N_21792,N_12620,N_15340);
and U21793 (N_21793,N_13870,N_14224);
nand U21794 (N_21794,N_14728,N_14596);
nor U21795 (N_21795,N_16778,N_15932);
and U21796 (N_21796,N_13925,N_13130);
or U21797 (N_21797,N_17169,N_18422);
and U21798 (N_21798,N_13557,N_17813);
or U21799 (N_21799,N_14775,N_13913);
nor U21800 (N_21800,N_12533,N_15987);
or U21801 (N_21801,N_17642,N_18209);
and U21802 (N_21802,N_17502,N_17588);
and U21803 (N_21803,N_13987,N_15696);
nor U21804 (N_21804,N_14773,N_16076);
or U21805 (N_21805,N_13604,N_15647);
nor U21806 (N_21806,N_18474,N_16958);
and U21807 (N_21807,N_16341,N_15322);
nand U21808 (N_21808,N_15965,N_18452);
xor U21809 (N_21809,N_12652,N_15928);
and U21810 (N_21810,N_12674,N_15084);
nand U21811 (N_21811,N_13723,N_14510);
nor U21812 (N_21812,N_13851,N_16508);
nor U21813 (N_21813,N_16602,N_13627);
nor U21814 (N_21814,N_16306,N_17737);
and U21815 (N_21815,N_14745,N_15606);
nor U21816 (N_21816,N_14988,N_16927);
nor U21817 (N_21817,N_15253,N_15095);
or U21818 (N_21818,N_15988,N_15926);
and U21819 (N_21819,N_17667,N_16664);
and U21820 (N_21820,N_17730,N_18149);
nand U21821 (N_21821,N_18718,N_16754);
and U21822 (N_21822,N_17610,N_17679);
nor U21823 (N_21823,N_15030,N_16572);
nor U21824 (N_21824,N_17947,N_12990);
or U21825 (N_21825,N_15046,N_15015);
and U21826 (N_21826,N_18517,N_18741);
and U21827 (N_21827,N_14890,N_13984);
nand U21828 (N_21828,N_15178,N_13873);
nand U21829 (N_21829,N_18089,N_17537);
nor U21830 (N_21830,N_15409,N_17623);
or U21831 (N_21831,N_12760,N_17451);
nand U21832 (N_21832,N_12886,N_16776);
nand U21833 (N_21833,N_14529,N_16087);
nand U21834 (N_21834,N_16333,N_13033);
or U21835 (N_21835,N_18428,N_15299);
nand U21836 (N_21836,N_14089,N_16053);
nand U21837 (N_21837,N_14212,N_13530);
and U21838 (N_21838,N_16780,N_15949);
or U21839 (N_21839,N_13566,N_16539);
nand U21840 (N_21840,N_17132,N_16784);
nor U21841 (N_21841,N_17653,N_12996);
and U21842 (N_21842,N_18343,N_13871);
and U21843 (N_21843,N_17470,N_14781);
nor U21844 (N_21844,N_14318,N_18143);
nand U21845 (N_21845,N_14485,N_18293);
or U21846 (N_21846,N_13200,N_18478);
and U21847 (N_21847,N_16250,N_17795);
or U21848 (N_21848,N_17800,N_16378);
nor U21849 (N_21849,N_13157,N_12732);
or U21850 (N_21850,N_15496,N_17550);
nand U21851 (N_21851,N_16067,N_17687);
or U21852 (N_21852,N_15549,N_16724);
nor U21853 (N_21853,N_16614,N_16171);
or U21854 (N_21854,N_15890,N_18097);
nor U21855 (N_21855,N_14933,N_12811);
nor U21856 (N_21856,N_17337,N_13102);
nand U21857 (N_21857,N_17018,N_18580);
and U21858 (N_21858,N_17219,N_17055);
and U21859 (N_21859,N_13854,N_14897);
nand U21860 (N_21860,N_15509,N_12670);
nand U21861 (N_21861,N_17918,N_16900);
and U21862 (N_21862,N_16065,N_17784);
or U21863 (N_21863,N_17828,N_14785);
and U21864 (N_21864,N_18732,N_12801);
nor U21865 (N_21865,N_13560,N_15293);
nand U21866 (N_21866,N_14198,N_17237);
nand U21867 (N_21867,N_17585,N_14042);
and U21868 (N_21868,N_16647,N_17656);
and U21869 (N_21869,N_16794,N_15682);
nand U21870 (N_21870,N_17017,N_14466);
or U21871 (N_21871,N_15976,N_15169);
nor U21872 (N_21872,N_14354,N_13911);
nand U21873 (N_21873,N_17977,N_14635);
nand U21874 (N_21874,N_14776,N_18130);
nand U21875 (N_21875,N_15374,N_13732);
nand U21876 (N_21876,N_16575,N_15970);
or U21877 (N_21877,N_18509,N_16448);
nor U21878 (N_21878,N_18156,N_17143);
or U21879 (N_21879,N_17484,N_13407);
nand U21880 (N_21880,N_17723,N_18251);
nor U21881 (N_21881,N_15891,N_18085);
nor U21882 (N_21882,N_18102,N_12883);
nand U21883 (N_21883,N_16454,N_17624);
nand U21884 (N_21884,N_17459,N_18265);
or U21885 (N_21885,N_12838,N_18290);
or U21886 (N_21886,N_18275,N_15690);
nor U21887 (N_21887,N_17781,N_17194);
or U21888 (N_21888,N_17056,N_13530);
or U21889 (N_21889,N_13644,N_12528);
and U21890 (N_21890,N_17059,N_14328);
or U21891 (N_21891,N_18499,N_16278);
and U21892 (N_21892,N_12505,N_17785);
nand U21893 (N_21893,N_14157,N_16762);
nand U21894 (N_21894,N_13931,N_15226);
or U21895 (N_21895,N_12520,N_16873);
or U21896 (N_21896,N_16195,N_14529);
or U21897 (N_21897,N_16312,N_16039);
or U21898 (N_21898,N_17787,N_13279);
nor U21899 (N_21899,N_13569,N_14308);
nand U21900 (N_21900,N_17744,N_17225);
nand U21901 (N_21901,N_14331,N_14995);
nand U21902 (N_21902,N_18478,N_12686);
or U21903 (N_21903,N_13256,N_14648);
nand U21904 (N_21904,N_13788,N_16014);
or U21905 (N_21905,N_16557,N_13281);
nand U21906 (N_21906,N_14096,N_14641);
nor U21907 (N_21907,N_15823,N_13070);
nor U21908 (N_21908,N_14142,N_18063);
and U21909 (N_21909,N_12951,N_15511);
nor U21910 (N_21910,N_18024,N_15070);
and U21911 (N_21911,N_17523,N_12777);
nor U21912 (N_21912,N_15248,N_14212);
nor U21913 (N_21913,N_18452,N_15798);
nand U21914 (N_21914,N_12742,N_18703);
nand U21915 (N_21915,N_13281,N_15770);
and U21916 (N_21916,N_18207,N_13196);
nand U21917 (N_21917,N_15412,N_14209);
or U21918 (N_21918,N_16781,N_17632);
nor U21919 (N_21919,N_18420,N_17532);
nand U21920 (N_21920,N_14322,N_14613);
and U21921 (N_21921,N_15553,N_16951);
and U21922 (N_21922,N_17688,N_17101);
nor U21923 (N_21923,N_13433,N_15566);
nand U21924 (N_21924,N_13493,N_16190);
or U21925 (N_21925,N_17866,N_16108);
nor U21926 (N_21926,N_13463,N_18520);
and U21927 (N_21927,N_14512,N_12940);
and U21928 (N_21928,N_15170,N_12883);
and U21929 (N_21929,N_18747,N_17720);
or U21930 (N_21930,N_17320,N_16238);
nor U21931 (N_21931,N_14211,N_17070);
nor U21932 (N_21932,N_16114,N_12852);
or U21933 (N_21933,N_14579,N_16600);
and U21934 (N_21934,N_15533,N_17243);
nand U21935 (N_21935,N_18123,N_14815);
nor U21936 (N_21936,N_15341,N_18443);
and U21937 (N_21937,N_13590,N_16234);
nor U21938 (N_21938,N_16607,N_13018);
nor U21939 (N_21939,N_13383,N_18178);
nand U21940 (N_21940,N_17682,N_16804);
and U21941 (N_21941,N_16081,N_13565);
nand U21942 (N_21942,N_15446,N_13652);
nand U21943 (N_21943,N_18567,N_14532);
nand U21944 (N_21944,N_16537,N_16141);
nand U21945 (N_21945,N_14813,N_15651);
nand U21946 (N_21946,N_17881,N_17897);
and U21947 (N_21947,N_17697,N_17662);
nand U21948 (N_21948,N_14507,N_17172);
or U21949 (N_21949,N_15784,N_12699);
and U21950 (N_21950,N_17136,N_17190);
and U21951 (N_21951,N_18028,N_13092);
nand U21952 (N_21952,N_17136,N_15245);
and U21953 (N_21953,N_14043,N_15567);
nor U21954 (N_21954,N_15145,N_17130);
nor U21955 (N_21955,N_15502,N_14849);
nor U21956 (N_21956,N_15672,N_16168);
and U21957 (N_21957,N_13811,N_15980);
and U21958 (N_21958,N_16883,N_13809);
and U21959 (N_21959,N_13739,N_12787);
nor U21960 (N_21960,N_15790,N_14818);
nor U21961 (N_21961,N_14551,N_14529);
and U21962 (N_21962,N_13072,N_17952);
nand U21963 (N_21963,N_15270,N_15786);
or U21964 (N_21964,N_18268,N_13357);
and U21965 (N_21965,N_15085,N_13829);
nand U21966 (N_21966,N_13525,N_12560);
or U21967 (N_21967,N_15472,N_18640);
and U21968 (N_21968,N_15096,N_18260);
or U21969 (N_21969,N_16711,N_12654);
xor U21970 (N_21970,N_18380,N_13609);
and U21971 (N_21971,N_15562,N_13982);
xor U21972 (N_21972,N_16708,N_16530);
nor U21973 (N_21973,N_17199,N_14014);
or U21974 (N_21974,N_16903,N_14416);
and U21975 (N_21975,N_15251,N_13928);
or U21976 (N_21976,N_17727,N_16852);
or U21977 (N_21977,N_17998,N_13498);
or U21978 (N_21978,N_16779,N_13797);
and U21979 (N_21979,N_16904,N_17390);
and U21980 (N_21980,N_14910,N_15648);
or U21981 (N_21981,N_13755,N_13006);
and U21982 (N_21982,N_13642,N_14900);
nor U21983 (N_21983,N_18298,N_16652);
or U21984 (N_21984,N_17587,N_14203);
nor U21985 (N_21985,N_13895,N_13552);
nand U21986 (N_21986,N_14258,N_18324);
or U21987 (N_21987,N_13695,N_14031);
nor U21988 (N_21988,N_14032,N_16790);
or U21989 (N_21989,N_15245,N_14236);
nor U21990 (N_21990,N_13429,N_13344);
and U21991 (N_21991,N_15322,N_18174);
or U21992 (N_21992,N_12658,N_18645);
and U21993 (N_21993,N_17813,N_12672);
nor U21994 (N_21994,N_14895,N_18710);
or U21995 (N_21995,N_15730,N_16371);
or U21996 (N_21996,N_16329,N_17862);
nor U21997 (N_21997,N_16806,N_14602);
or U21998 (N_21998,N_17844,N_14786);
or U21999 (N_21999,N_14835,N_15715);
and U22000 (N_22000,N_16068,N_16861);
nor U22001 (N_22001,N_16675,N_16751);
nor U22002 (N_22002,N_18511,N_17555);
nand U22003 (N_22003,N_18696,N_15676);
nor U22004 (N_22004,N_14941,N_13118);
or U22005 (N_22005,N_16871,N_15921);
or U22006 (N_22006,N_15722,N_18223);
and U22007 (N_22007,N_18584,N_14046);
and U22008 (N_22008,N_15354,N_13793);
nor U22009 (N_22009,N_16690,N_15950);
and U22010 (N_22010,N_14129,N_13150);
and U22011 (N_22011,N_14515,N_13013);
nand U22012 (N_22012,N_17079,N_18637);
nand U22013 (N_22013,N_13473,N_15443);
and U22014 (N_22014,N_18229,N_12952);
and U22015 (N_22015,N_14419,N_14247);
and U22016 (N_22016,N_18348,N_17478);
and U22017 (N_22017,N_17862,N_12833);
or U22018 (N_22018,N_14267,N_16424);
and U22019 (N_22019,N_13271,N_14684);
and U22020 (N_22020,N_14156,N_15793);
nand U22021 (N_22021,N_17647,N_12663);
nor U22022 (N_22022,N_15207,N_15857);
or U22023 (N_22023,N_16027,N_17003);
and U22024 (N_22024,N_13866,N_13786);
or U22025 (N_22025,N_12689,N_14802);
and U22026 (N_22026,N_18565,N_13309);
and U22027 (N_22027,N_17586,N_17763);
and U22028 (N_22028,N_12566,N_16243);
xnor U22029 (N_22029,N_14324,N_13825);
nor U22030 (N_22030,N_13518,N_14094);
or U22031 (N_22031,N_15494,N_15385);
and U22032 (N_22032,N_15303,N_13941);
or U22033 (N_22033,N_17536,N_16182);
nand U22034 (N_22034,N_15953,N_12622);
and U22035 (N_22035,N_16433,N_15135);
or U22036 (N_22036,N_18086,N_13266);
or U22037 (N_22037,N_18727,N_14951);
nand U22038 (N_22038,N_12737,N_12799);
nor U22039 (N_22039,N_13212,N_14901);
or U22040 (N_22040,N_17210,N_18508);
and U22041 (N_22041,N_18128,N_15552);
nand U22042 (N_22042,N_14988,N_15907);
and U22043 (N_22043,N_17740,N_17763);
or U22044 (N_22044,N_17230,N_15746);
or U22045 (N_22045,N_15350,N_14521);
xnor U22046 (N_22046,N_16943,N_16702);
nor U22047 (N_22047,N_18358,N_14435);
nand U22048 (N_22048,N_18073,N_14606);
nand U22049 (N_22049,N_12679,N_15936);
nor U22050 (N_22050,N_13705,N_13370);
and U22051 (N_22051,N_13472,N_18603);
nand U22052 (N_22052,N_13082,N_12694);
or U22053 (N_22053,N_18044,N_14991);
or U22054 (N_22054,N_12885,N_16334);
and U22055 (N_22055,N_18025,N_16468);
nand U22056 (N_22056,N_13212,N_16485);
or U22057 (N_22057,N_15645,N_17886);
and U22058 (N_22058,N_14332,N_13985);
nor U22059 (N_22059,N_16682,N_16343);
and U22060 (N_22060,N_13039,N_18741);
nand U22061 (N_22061,N_18063,N_14191);
or U22062 (N_22062,N_17113,N_13343);
and U22063 (N_22063,N_18218,N_13162);
nor U22064 (N_22064,N_16279,N_14104);
nand U22065 (N_22065,N_12712,N_13149);
and U22066 (N_22066,N_13459,N_16869);
or U22067 (N_22067,N_14760,N_14452);
nor U22068 (N_22068,N_17090,N_16290);
or U22069 (N_22069,N_17544,N_16142);
nand U22070 (N_22070,N_13662,N_13274);
or U22071 (N_22071,N_14189,N_17786);
nand U22072 (N_22072,N_13500,N_16337);
nor U22073 (N_22073,N_14787,N_13266);
nand U22074 (N_22074,N_17165,N_15741);
nor U22075 (N_22075,N_17225,N_13110);
nor U22076 (N_22076,N_12696,N_16475);
nand U22077 (N_22077,N_14456,N_17147);
or U22078 (N_22078,N_14506,N_14072);
and U22079 (N_22079,N_16461,N_16800);
and U22080 (N_22080,N_15235,N_13057);
nand U22081 (N_22081,N_16808,N_14856);
nand U22082 (N_22082,N_16797,N_13997);
nor U22083 (N_22083,N_13332,N_15859);
and U22084 (N_22084,N_17101,N_17548);
nand U22085 (N_22085,N_16607,N_17186);
and U22086 (N_22086,N_16065,N_17739);
nor U22087 (N_22087,N_17888,N_17426);
and U22088 (N_22088,N_16377,N_14137);
nand U22089 (N_22089,N_18262,N_18225);
or U22090 (N_22090,N_17377,N_16068);
nor U22091 (N_22091,N_15549,N_13639);
or U22092 (N_22092,N_16336,N_16185);
nor U22093 (N_22093,N_14278,N_15912);
nand U22094 (N_22094,N_16987,N_18674);
nand U22095 (N_22095,N_13932,N_18532);
and U22096 (N_22096,N_14378,N_14408);
and U22097 (N_22097,N_16701,N_16168);
nor U22098 (N_22098,N_14132,N_16430);
nand U22099 (N_22099,N_17595,N_14592);
nor U22100 (N_22100,N_14175,N_17003);
nand U22101 (N_22101,N_16779,N_12591);
or U22102 (N_22102,N_12786,N_15358);
and U22103 (N_22103,N_13305,N_17706);
or U22104 (N_22104,N_18269,N_16408);
and U22105 (N_22105,N_17787,N_15005);
and U22106 (N_22106,N_14746,N_13597);
or U22107 (N_22107,N_17892,N_15651);
or U22108 (N_22108,N_16879,N_14801);
nor U22109 (N_22109,N_12773,N_15952);
and U22110 (N_22110,N_17726,N_13488);
nand U22111 (N_22111,N_12624,N_17951);
or U22112 (N_22112,N_18400,N_18270);
nand U22113 (N_22113,N_13985,N_16521);
and U22114 (N_22114,N_12664,N_13812);
nand U22115 (N_22115,N_15163,N_17194);
nand U22116 (N_22116,N_12823,N_13123);
or U22117 (N_22117,N_14220,N_14111);
nand U22118 (N_22118,N_15967,N_18664);
nand U22119 (N_22119,N_15468,N_13446);
nor U22120 (N_22120,N_15063,N_13109);
and U22121 (N_22121,N_17572,N_18394);
and U22122 (N_22122,N_18035,N_17856);
and U22123 (N_22123,N_17229,N_15617);
nor U22124 (N_22124,N_17238,N_15422);
nor U22125 (N_22125,N_17206,N_16289);
nor U22126 (N_22126,N_17951,N_18559);
nand U22127 (N_22127,N_14015,N_16563);
nor U22128 (N_22128,N_12523,N_13344);
or U22129 (N_22129,N_12725,N_14672);
and U22130 (N_22130,N_13310,N_16632);
nor U22131 (N_22131,N_17688,N_14621);
or U22132 (N_22132,N_13301,N_14369);
nand U22133 (N_22133,N_15050,N_13749);
and U22134 (N_22134,N_18197,N_14120);
or U22135 (N_22135,N_13698,N_18142);
or U22136 (N_22136,N_18205,N_18659);
nor U22137 (N_22137,N_16542,N_14324);
or U22138 (N_22138,N_17361,N_18471);
nand U22139 (N_22139,N_12617,N_14765);
nor U22140 (N_22140,N_16675,N_15615);
or U22141 (N_22141,N_15842,N_14476);
and U22142 (N_22142,N_18442,N_16567);
and U22143 (N_22143,N_14952,N_14292);
nand U22144 (N_22144,N_18070,N_16538);
nand U22145 (N_22145,N_14637,N_15984);
and U22146 (N_22146,N_17112,N_15871);
or U22147 (N_22147,N_15497,N_16054);
or U22148 (N_22148,N_16995,N_13345);
or U22149 (N_22149,N_16089,N_15338);
nor U22150 (N_22150,N_17859,N_17409);
nand U22151 (N_22151,N_13039,N_16400);
nand U22152 (N_22152,N_14367,N_18489);
and U22153 (N_22153,N_18474,N_15837);
and U22154 (N_22154,N_15896,N_13267);
or U22155 (N_22155,N_14698,N_17220);
and U22156 (N_22156,N_16681,N_15747);
or U22157 (N_22157,N_15182,N_12949);
nor U22158 (N_22158,N_16778,N_14508);
nand U22159 (N_22159,N_18267,N_15413);
nand U22160 (N_22160,N_16374,N_14770);
nand U22161 (N_22161,N_16792,N_16194);
or U22162 (N_22162,N_16953,N_13174);
nor U22163 (N_22163,N_16528,N_16442);
nand U22164 (N_22164,N_13540,N_14333);
or U22165 (N_22165,N_13173,N_16188);
or U22166 (N_22166,N_14999,N_17774);
nor U22167 (N_22167,N_13719,N_17627);
nor U22168 (N_22168,N_16137,N_14402);
or U22169 (N_22169,N_12923,N_16132);
nand U22170 (N_22170,N_16207,N_13628);
or U22171 (N_22171,N_16350,N_15529);
nand U22172 (N_22172,N_16954,N_17715);
or U22173 (N_22173,N_12746,N_14157);
nand U22174 (N_22174,N_16925,N_15709);
nand U22175 (N_22175,N_14114,N_16822);
nor U22176 (N_22176,N_14585,N_18454);
or U22177 (N_22177,N_16026,N_18394);
nor U22178 (N_22178,N_13423,N_17178);
nor U22179 (N_22179,N_16686,N_18610);
nand U22180 (N_22180,N_16198,N_16397);
and U22181 (N_22181,N_16253,N_16361);
nand U22182 (N_22182,N_13677,N_16155);
nand U22183 (N_22183,N_17989,N_13114);
and U22184 (N_22184,N_13249,N_18101);
nand U22185 (N_22185,N_14250,N_15888);
and U22186 (N_22186,N_15312,N_16410);
or U22187 (N_22187,N_13038,N_17108);
or U22188 (N_22188,N_13685,N_13274);
and U22189 (N_22189,N_16216,N_15400);
nand U22190 (N_22190,N_13918,N_13097);
nor U22191 (N_22191,N_17299,N_13670);
and U22192 (N_22192,N_17832,N_14148);
and U22193 (N_22193,N_12639,N_15597);
or U22194 (N_22194,N_18165,N_13481);
and U22195 (N_22195,N_14815,N_16643);
nand U22196 (N_22196,N_13175,N_18665);
nand U22197 (N_22197,N_13541,N_14308);
nand U22198 (N_22198,N_14552,N_13138);
or U22199 (N_22199,N_16496,N_14531);
nand U22200 (N_22200,N_12736,N_16127);
and U22201 (N_22201,N_17151,N_13940);
and U22202 (N_22202,N_14624,N_16268);
nor U22203 (N_22203,N_15985,N_15499);
nor U22204 (N_22204,N_13509,N_12648);
nand U22205 (N_22205,N_17122,N_15026);
and U22206 (N_22206,N_17830,N_13837);
or U22207 (N_22207,N_17703,N_18260);
nor U22208 (N_22208,N_16084,N_14234);
nor U22209 (N_22209,N_18465,N_14915);
nor U22210 (N_22210,N_16348,N_16620);
nor U22211 (N_22211,N_17427,N_14027);
xnor U22212 (N_22212,N_13817,N_15282);
or U22213 (N_22213,N_18121,N_13663);
or U22214 (N_22214,N_13576,N_14901);
xnor U22215 (N_22215,N_18709,N_14216);
nand U22216 (N_22216,N_16657,N_18744);
nor U22217 (N_22217,N_14128,N_15415);
or U22218 (N_22218,N_17484,N_15203);
nand U22219 (N_22219,N_16118,N_14571);
nand U22220 (N_22220,N_18637,N_17322);
nand U22221 (N_22221,N_16038,N_17741);
or U22222 (N_22222,N_17685,N_14825);
or U22223 (N_22223,N_16278,N_12718);
nor U22224 (N_22224,N_14805,N_13503);
or U22225 (N_22225,N_12953,N_17480);
or U22226 (N_22226,N_17470,N_18187);
and U22227 (N_22227,N_12959,N_14929);
nor U22228 (N_22228,N_14548,N_17766);
xnor U22229 (N_22229,N_14169,N_15820);
and U22230 (N_22230,N_14946,N_15406);
nor U22231 (N_22231,N_18518,N_16330);
or U22232 (N_22232,N_13840,N_16262);
nand U22233 (N_22233,N_16145,N_16729);
nor U22234 (N_22234,N_17614,N_16843);
nor U22235 (N_22235,N_13034,N_17539);
nor U22236 (N_22236,N_17199,N_17160);
or U22237 (N_22237,N_16419,N_12588);
or U22238 (N_22238,N_15565,N_15147);
xnor U22239 (N_22239,N_18000,N_12897);
nand U22240 (N_22240,N_14595,N_17447);
nand U22241 (N_22241,N_16232,N_14346);
or U22242 (N_22242,N_17777,N_17587);
nor U22243 (N_22243,N_12759,N_12954);
nor U22244 (N_22244,N_15389,N_15596);
nand U22245 (N_22245,N_15839,N_15631);
nor U22246 (N_22246,N_14262,N_16024);
or U22247 (N_22247,N_18542,N_16054);
and U22248 (N_22248,N_18195,N_15446);
nand U22249 (N_22249,N_15107,N_14125);
or U22250 (N_22250,N_15763,N_16362);
nand U22251 (N_22251,N_13272,N_17579);
and U22252 (N_22252,N_17609,N_18637);
or U22253 (N_22253,N_16329,N_17731);
nor U22254 (N_22254,N_18335,N_16102);
nor U22255 (N_22255,N_18007,N_14596);
nand U22256 (N_22256,N_14526,N_18323);
nand U22257 (N_22257,N_14108,N_18644);
or U22258 (N_22258,N_17380,N_16554);
nand U22259 (N_22259,N_12832,N_12944);
xor U22260 (N_22260,N_18185,N_13036);
or U22261 (N_22261,N_16104,N_14994);
nand U22262 (N_22262,N_18157,N_15410);
nor U22263 (N_22263,N_14254,N_16677);
nor U22264 (N_22264,N_16820,N_17267);
nor U22265 (N_22265,N_18740,N_14100);
nand U22266 (N_22266,N_18500,N_12663);
nand U22267 (N_22267,N_15933,N_18045);
nand U22268 (N_22268,N_13304,N_15027);
nand U22269 (N_22269,N_15746,N_16231);
or U22270 (N_22270,N_16172,N_16972);
nor U22271 (N_22271,N_14588,N_18682);
or U22272 (N_22272,N_14596,N_15954);
nand U22273 (N_22273,N_14261,N_16792);
or U22274 (N_22274,N_16118,N_13668);
nor U22275 (N_22275,N_14060,N_13218);
or U22276 (N_22276,N_16870,N_16121);
and U22277 (N_22277,N_14061,N_13509);
xor U22278 (N_22278,N_17106,N_16032);
and U22279 (N_22279,N_15026,N_13525);
and U22280 (N_22280,N_13441,N_14118);
nor U22281 (N_22281,N_16990,N_14468);
nor U22282 (N_22282,N_17655,N_15788);
nand U22283 (N_22283,N_15026,N_14851);
and U22284 (N_22284,N_13126,N_14893);
nand U22285 (N_22285,N_14032,N_16226);
or U22286 (N_22286,N_18672,N_17011);
or U22287 (N_22287,N_18205,N_17464);
nor U22288 (N_22288,N_15892,N_14589);
and U22289 (N_22289,N_17337,N_12809);
xor U22290 (N_22290,N_15942,N_13757);
nor U22291 (N_22291,N_14510,N_15033);
and U22292 (N_22292,N_15239,N_12649);
nor U22293 (N_22293,N_14888,N_15415);
and U22294 (N_22294,N_14611,N_18697);
nand U22295 (N_22295,N_14764,N_14593);
and U22296 (N_22296,N_13026,N_18052);
and U22297 (N_22297,N_18092,N_15323);
nand U22298 (N_22298,N_13842,N_15050);
or U22299 (N_22299,N_18682,N_12958);
or U22300 (N_22300,N_14526,N_14979);
nand U22301 (N_22301,N_13063,N_17350);
and U22302 (N_22302,N_14150,N_16832);
nand U22303 (N_22303,N_17862,N_14837);
xor U22304 (N_22304,N_14907,N_18686);
and U22305 (N_22305,N_18145,N_14290);
and U22306 (N_22306,N_14347,N_16617);
nand U22307 (N_22307,N_16131,N_14849);
or U22308 (N_22308,N_13954,N_17345);
nor U22309 (N_22309,N_14033,N_14596);
nor U22310 (N_22310,N_16152,N_12554);
nand U22311 (N_22311,N_18592,N_18510);
and U22312 (N_22312,N_17483,N_17880);
and U22313 (N_22313,N_13694,N_17145);
or U22314 (N_22314,N_14123,N_17150);
nand U22315 (N_22315,N_13925,N_13485);
or U22316 (N_22316,N_13204,N_14000);
and U22317 (N_22317,N_17467,N_14830);
or U22318 (N_22318,N_12858,N_18698);
or U22319 (N_22319,N_14855,N_17465);
and U22320 (N_22320,N_14704,N_14455);
nand U22321 (N_22321,N_18682,N_13027);
nand U22322 (N_22322,N_17034,N_16964);
and U22323 (N_22323,N_16971,N_13504);
nor U22324 (N_22324,N_15012,N_17487);
or U22325 (N_22325,N_13296,N_15787);
and U22326 (N_22326,N_16519,N_18248);
or U22327 (N_22327,N_14229,N_13160);
and U22328 (N_22328,N_14661,N_15541);
and U22329 (N_22329,N_14822,N_12673);
and U22330 (N_22330,N_15465,N_13691);
nor U22331 (N_22331,N_14521,N_13366);
nor U22332 (N_22332,N_17021,N_16285);
nand U22333 (N_22333,N_13823,N_13146);
or U22334 (N_22334,N_12725,N_14659);
nor U22335 (N_22335,N_14275,N_14199);
nand U22336 (N_22336,N_16357,N_15960);
and U22337 (N_22337,N_16628,N_17041);
and U22338 (N_22338,N_17435,N_14073);
and U22339 (N_22339,N_16168,N_14019);
nor U22340 (N_22340,N_17581,N_17336);
and U22341 (N_22341,N_16820,N_17838);
nand U22342 (N_22342,N_13592,N_14959);
and U22343 (N_22343,N_15550,N_16595);
and U22344 (N_22344,N_15994,N_16153);
nor U22345 (N_22345,N_14592,N_15809);
nor U22346 (N_22346,N_14980,N_14046);
or U22347 (N_22347,N_12928,N_18073);
and U22348 (N_22348,N_18333,N_16982);
nor U22349 (N_22349,N_16688,N_17960);
nand U22350 (N_22350,N_17237,N_18740);
nor U22351 (N_22351,N_17589,N_14702);
nand U22352 (N_22352,N_14335,N_15219);
or U22353 (N_22353,N_16945,N_17138);
nand U22354 (N_22354,N_12756,N_14296);
nor U22355 (N_22355,N_17281,N_15731);
nor U22356 (N_22356,N_12553,N_13821);
or U22357 (N_22357,N_18101,N_17252);
nand U22358 (N_22358,N_18096,N_12564);
or U22359 (N_22359,N_16208,N_13313);
and U22360 (N_22360,N_18320,N_16701);
and U22361 (N_22361,N_18450,N_12767);
and U22362 (N_22362,N_12768,N_18238);
nand U22363 (N_22363,N_13106,N_16513);
nand U22364 (N_22364,N_17969,N_17058);
nor U22365 (N_22365,N_12908,N_14266);
nor U22366 (N_22366,N_16872,N_12544);
nand U22367 (N_22367,N_15174,N_17047);
nor U22368 (N_22368,N_13898,N_18735);
nand U22369 (N_22369,N_15882,N_16088);
nor U22370 (N_22370,N_14518,N_14389);
nand U22371 (N_22371,N_17362,N_16661);
and U22372 (N_22372,N_15135,N_15349);
nor U22373 (N_22373,N_15289,N_17092);
nand U22374 (N_22374,N_17467,N_13601);
nand U22375 (N_22375,N_16235,N_13522);
nand U22376 (N_22376,N_14125,N_13512);
and U22377 (N_22377,N_15287,N_14803);
and U22378 (N_22378,N_13958,N_17434);
and U22379 (N_22379,N_18667,N_14864);
and U22380 (N_22380,N_14130,N_12504);
or U22381 (N_22381,N_12540,N_18339);
and U22382 (N_22382,N_14336,N_12557);
nor U22383 (N_22383,N_14466,N_15385);
nor U22384 (N_22384,N_14623,N_17077);
nand U22385 (N_22385,N_14422,N_16964);
nand U22386 (N_22386,N_16197,N_12636);
and U22387 (N_22387,N_16720,N_16902);
and U22388 (N_22388,N_12585,N_15261);
nor U22389 (N_22389,N_15256,N_18033);
nand U22390 (N_22390,N_17908,N_17338);
or U22391 (N_22391,N_14402,N_13520);
nand U22392 (N_22392,N_17051,N_14146);
nor U22393 (N_22393,N_13413,N_13574);
or U22394 (N_22394,N_13559,N_13796);
nor U22395 (N_22395,N_17280,N_16475);
or U22396 (N_22396,N_15050,N_14369);
or U22397 (N_22397,N_17606,N_15510);
or U22398 (N_22398,N_16209,N_14641);
nand U22399 (N_22399,N_15893,N_13813);
or U22400 (N_22400,N_15429,N_15036);
and U22401 (N_22401,N_17381,N_12727);
nand U22402 (N_22402,N_13412,N_13922);
nand U22403 (N_22403,N_17140,N_13368);
nand U22404 (N_22404,N_13264,N_15850);
nand U22405 (N_22405,N_16806,N_15223);
nand U22406 (N_22406,N_13918,N_15995);
nor U22407 (N_22407,N_13771,N_13687);
nand U22408 (N_22408,N_17384,N_17367);
nand U22409 (N_22409,N_12535,N_16042);
and U22410 (N_22410,N_16027,N_13197);
nand U22411 (N_22411,N_13850,N_12895);
nor U22412 (N_22412,N_12502,N_12824);
nor U22413 (N_22413,N_15211,N_17800);
nand U22414 (N_22414,N_15971,N_15092);
and U22415 (N_22415,N_17895,N_14981);
and U22416 (N_22416,N_16428,N_13735);
nand U22417 (N_22417,N_14503,N_18038);
nand U22418 (N_22418,N_17415,N_12809);
and U22419 (N_22419,N_13745,N_18473);
and U22420 (N_22420,N_13347,N_12505);
nor U22421 (N_22421,N_17417,N_17325);
or U22422 (N_22422,N_18451,N_18322);
nor U22423 (N_22423,N_15288,N_14827);
or U22424 (N_22424,N_14462,N_16196);
nand U22425 (N_22425,N_14111,N_13694);
and U22426 (N_22426,N_15582,N_14482);
or U22427 (N_22427,N_16079,N_15703);
nand U22428 (N_22428,N_12576,N_13984);
and U22429 (N_22429,N_14284,N_17168);
nor U22430 (N_22430,N_17895,N_17390);
or U22431 (N_22431,N_14494,N_16808);
xnor U22432 (N_22432,N_16389,N_12684);
nand U22433 (N_22433,N_16801,N_18024);
nand U22434 (N_22434,N_13284,N_15510);
and U22435 (N_22435,N_16433,N_14075);
nand U22436 (N_22436,N_14053,N_12749);
and U22437 (N_22437,N_14342,N_13509);
nor U22438 (N_22438,N_18491,N_14604);
nor U22439 (N_22439,N_15637,N_17487);
nor U22440 (N_22440,N_13738,N_13024);
nor U22441 (N_22441,N_12627,N_14111);
xor U22442 (N_22442,N_17932,N_15553);
and U22443 (N_22443,N_15634,N_14080);
and U22444 (N_22444,N_14289,N_13075);
nand U22445 (N_22445,N_15126,N_18744);
or U22446 (N_22446,N_13239,N_18630);
nand U22447 (N_22447,N_16333,N_13931);
or U22448 (N_22448,N_13454,N_13753);
nand U22449 (N_22449,N_16687,N_12520);
xor U22450 (N_22450,N_16120,N_17765);
or U22451 (N_22451,N_15995,N_16631);
and U22452 (N_22452,N_14302,N_16243);
or U22453 (N_22453,N_14766,N_13046);
or U22454 (N_22454,N_18057,N_18020);
nand U22455 (N_22455,N_15894,N_17661);
nand U22456 (N_22456,N_18432,N_15519);
nor U22457 (N_22457,N_17895,N_16698);
nor U22458 (N_22458,N_13964,N_13137);
and U22459 (N_22459,N_17091,N_16368);
and U22460 (N_22460,N_12657,N_17043);
and U22461 (N_22461,N_15670,N_13606);
nand U22462 (N_22462,N_17398,N_13963);
nor U22463 (N_22463,N_15282,N_13048);
and U22464 (N_22464,N_16760,N_17903);
xnor U22465 (N_22465,N_16159,N_14689);
or U22466 (N_22466,N_13175,N_16890);
nor U22467 (N_22467,N_15799,N_15481);
and U22468 (N_22468,N_15209,N_12894);
nand U22469 (N_22469,N_14497,N_18619);
nand U22470 (N_22470,N_13567,N_15344);
nand U22471 (N_22471,N_15607,N_16430);
nand U22472 (N_22472,N_16080,N_18326);
nor U22473 (N_22473,N_16715,N_16928);
or U22474 (N_22474,N_15087,N_13852);
and U22475 (N_22475,N_12691,N_17928);
nor U22476 (N_22476,N_15153,N_14530);
and U22477 (N_22477,N_13749,N_18483);
nand U22478 (N_22478,N_14962,N_18681);
nand U22479 (N_22479,N_12521,N_13477);
nand U22480 (N_22480,N_14944,N_16430);
nor U22481 (N_22481,N_13136,N_13075);
nor U22482 (N_22482,N_16537,N_13669);
nand U22483 (N_22483,N_15434,N_14950);
nor U22484 (N_22484,N_12790,N_17568);
and U22485 (N_22485,N_14363,N_15013);
nand U22486 (N_22486,N_17748,N_17382);
nor U22487 (N_22487,N_14253,N_16362);
and U22488 (N_22488,N_14663,N_16825);
or U22489 (N_22489,N_13062,N_17080);
nor U22490 (N_22490,N_13541,N_14280);
or U22491 (N_22491,N_14577,N_13892);
nor U22492 (N_22492,N_16561,N_16313);
nor U22493 (N_22493,N_15820,N_16217);
and U22494 (N_22494,N_18707,N_16608);
nand U22495 (N_22495,N_15229,N_14480);
and U22496 (N_22496,N_13428,N_17442);
and U22497 (N_22497,N_15942,N_13855);
nor U22498 (N_22498,N_16066,N_13322);
or U22499 (N_22499,N_18721,N_17256);
xnor U22500 (N_22500,N_17018,N_13637);
or U22501 (N_22501,N_15098,N_17092);
or U22502 (N_22502,N_12747,N_13021);
xnor U22503 (N_22503,N_16851,N_13996);
or U22504 (N_22504,N_13686,N_15982);
or U22505 (N_22505,N_17612,N_17637);
nor U22506 (N_22506,N_17687,N_15920);
nand U22507 (N_22507,N_17341,N_15277);
nand U22508 (N_22508,N_16304,N_18555);
or U22509 (N_22509,N_16611,N_18473);
nand U22510 (N_22510,N_14681,N_14149);
and U22511 (N_22511,N_18567,N_12583);
or U22512 (N_22512,N_15413,N_15405);
or U22513 (N_22513,N_14199,N_16985);
nor U22514 (N_22514,N_15212,N_12892);
nor U22515 (N_22515,N_17592,N_16255);
and U22516 (N_22516,N_14825,N_18564);
and U22517 (N_22517,N_13308,N_13477);
nor U22518 (N_22518,N_18051,N_14794);
and U22519 (N_22519,N_16575,N_18688);
nand U22520 (N_22520,N_17156,N_14446);
nand U22521 (N_22521,N_13199,N_12680);
nor U22522 (N_22522,N_16031,N_15488);
and U22523 (N_22523,N_12684,N_15523);
or U22524 (N_22524,N_17515,N_15010);
nor U22525 (N_22525,N_16058,N_15145);
or U22526 (N_22526,N_18740,N_12657);
nand U22527 (N_22527,N_16431,N_14300);
nand U22528 (N_22528,N_12990,N_13729);
or U22529 (N_22529,N_15137,N_17205);
or U22530 (N_22530,N_17485,N_15921);
or U22531 (N_22531,N_14432,N_13026);
or U22532 (N_22532,N_16899,N_12746);
and U22533 (N_22533,N_16590,N_17564);
and U22534 (N_22534,N_13224,N_16017);
and U22535 (N_22535,N_16099,N_15057);
nor U22536 (N_22536,N_18238,N_15337);
or U22537 (N_22537,N_17155,N_16446);
nor U22538 (N_22538,N_13292,N_13311);
or U22539 (N_22539,N_17366,N_14608);
nor U22540 (N_22540,N_15137,N_13356);
or U22541 (N_22541,N_13928,N_13251);
nand U22542 (N_22542,N_18519,N_18333);
and U22543 (N_22543,N_16941,N_18444);
nand U22544 (N_22544,N_17149,N_16727);
nor U22545 (N_22545,N_17892,N_17059);
nand U22546 (N_22546,N_16096,N_17279);
or U22547 (N_22547,N_17101,N_14855);
or U22548 (N_22548,N_18065,N_14628);
nor U22549 (N_22549,N_12659,N_12956);
nand U22550 (N_22550,N_13660,N_17610);
nor U22551 (N_22551,N_14917,N_16789);
nor U22552 (N_22552,N_16651,N_16890);
or U22553 (N_22553,N_18686,N_13980);
nand U22554 (N_22554,N_15919,N_13197);
or U22555 (N_22555,N_15394,N_15791);
or U22556 (N_22556,N_16476,N_16605);
or U22557 (N_22557,N_17398,N_17983);
and U22558 (N_22558,N_14047,N_14752);
nand U22559 (N_22559,N_18133,N_17231);
nor U22560 (N_22560,N_13774,N_13431);
nand U22561 (N_22561,N_12993,N_13731);
and U22562 (N_22562,N_14964,N_12926);
nand U22563 (N_22563,N_16263,N_15178);
or U22564 (N_22564,N_18611,N_15064);
or U22565 (N_22565,N_18181,N_16186);
nand U22566 (N_22566,N_15409,N_15612);
or U22567 (N_22567,N_17269,N_15151);
nand U22568 (N_22568,N_18513,N_15767);
and U22569 (N_22569,N_16536,N_14569);
nand U22570 (N_22570,N_15198,N_15327);
and U22571 (N_22571,N_13449,N_14825);
or U22572 (N_22572,N_13843,N_16984);
and U22573 (N_22573,N_18395,N_16560);
nand U22574 (N_22574,N_17680,N_13347);
nand U22575 (N_22575,N_13323,N_17419);
nand U22576 (N_22576,N_18512,N_14297);
nor U22577 (N_22577,N_13947,N_16796);
or U22578 (N_22578,N_16825,N_17061);
and U22579 (N_22579,N_15738,N_17594);
and U22580 (N_22580,N_17734,N_18032);
nand U22581 (N_22581,N_16913,N_16800);
or U22582 (N_22582,N_13278,N_14189);
and U22583 (N_22583,N_14745,N_16117);
nor U22584 (N_22584,N_18221,N_16278);
nand U22585 (N_22585,N_16395,N_14666);
and U22586 (N_22586,N_17452,N_18633);
nand U22587 (N_22587,N_14745,N_16669);
and U22588 (N_22588,N_17818,N_16197);
or U22589 (N_22589,N_16918,N_14194);
and U22590 (N_22590,N_16276,N_13048);
and U22591 (N_22591,N_18072,N_15346);
nand U22592 (N_22592,N_13068,N_16023);
nand U22593 (N_22593,N_14462,N_15488);
nand U22594 (N_22594,N_17533,N_13029);
and U22595 (N_22595,N_18301,N_17353);
nor U22596 (N_22596,N_17467,N_18701);
or U22597 (N_22597,N_13344,N_18682);
or U22598 (N_22598,N_16554,N_17793);
or U22599 (N_22599,N_15670,N_12881);
nand U22600 (N_22600,N_16457,N_13163);
and U22601 (N_22601,N_13512,N_17579);
and U22602 (N_22602,N_18435,N_14697);
or U22603 (N_22603,N_17557,N_14218);
and U22604 (N_22604,N_15414,N_18645);
or U22605 (N_22605,N_13724,N_17802);
nor U22606 (N_22606,N_13242,N_13023);
and U22607 (N_22607,N_15977,N_18485);
or U22608 (N_22608,N_16721,N_12751);
or U22609 (N_22609,N_13430,N_12732);
or U22610 (N_22610,N_14539,N_18511);
nand U22611 (N_22611,N_15728,N_17898);
or U22612 (N_22612,N_14857,N_12781);
nand U22613 (N_22613,N_14762,N_18309);
nand U22614 (N_22614,N_16498,N_15532);
or U22615 (N_22615,N_17957,N_13997);
nor U22616 (N_22616,N_14989,N_16331);
nor U22617 (N_22617,N_15981,N_13361);
or U22618 (N_22618,N_13833,N_13122);
nand U22619 (N_22619,N_17581,N_16487);
nand U22620 (N_22620,N_14267,N_18430);
nor U22621 (N_22621,N_16048,N_17301);
nor U22622 (N_22622,N_16699,N_14905);
nor U22623 (N_22623,N_17382,N_12677);
nor U22624 (N_22624,N_16079,N_16748);
and U22625 (N_22625,N_17140,N_18506);
nand U22626 (N_22626,N_13315,N_17648);
and U22627 (N_22627,N_17094,N_18123);
xor U22628 (N_22628,N_16386,N_14497);
and U22629 (N_22629,N_15281,N_16457);
or U22630 (N_22630,N_17269,N_15154);
and U22631 (N_22631,N_18152,N_15151);
or U22632 (N_22632,N_14406,N_12760);
and U22633 (N_22633,N_14964,N_15913);
nor U22634 (N_22634,N_15303,N_14190);
and U22635 (N_22635,N_13153,N_18717);
nor U22636 (N_22636,N_16716,N_18715);
and U22637 (N_22637,N_13760,N_13622);
nand U22638 (N_22638,N_16053,N_17771);
nand U22639 (N_22639,N_16598,N_17818);
nand U22640 (N_22640,N_17705,N_12544);
and U22641 (N_22641,N_15341,N_16682);
nor U22642 (N_22642,N_16214,N_12624);
or U22643 (N_22643,N_14719,N_13509);
nor U22644 (N_22644,N_17017,N_14368);
or U22645 (N_22645,N_14624,N_13529);
nor U22646 (N_22646,N_14547,N_16180);
nor U22647 (N_22647,N_17829,N_17859);
nand U22648 (N_22648,N_13008,N_12651);
or U22649 (N_22649,N_18132,N_14926);
nor U22650 (N_22650,N_18153,N_13504);
nor U22651 (N_22651,N_17861,N_16537);
nor U22652 (N_22652,N_15575,N_15945);
nand U22653 (N_22653,N_13452,N_14572);
or U22654 (N_22654,N_15462,N_14688);
or U22655 (N_22655,N_17360,N_16401);
nand U22656 (N_22656,N_17399,N_18140);
and U22657 (N_22657,N_13990,N_15605);
or U22658 (N_22658,N_15109,N_14455);
nand U22659 (N_22659,N_15412,N_13662);
or U22660 (N_22660,N_18619,N_17887);
nor U22661 (N_22661,N_15736,N_18260);
or U22662 (N_22662,N_13492,N_17589);
and U22663 (N_22663,N_14642,N_16554);
nor U22664 (N_22664,N_13441,N_16021);
nor U22665 (N_22665,N_15964,N_18019);
nor U22666 (N_22666,N_15592,N_18173);
or U22667 (N_22667,N_13456,N_14977);
and U22668 (N_22668,N_13379,N_12642);
or U22669 (N_22669,N_14807,N_13337);
nand U22670 (N_22670,N_16404,N_18629);
and U22671 (N_22671,N_13119,N_17205);
nor U22672 (N_22672,N_16941,N_12599);
and U22673 (N_22673,N_18226,N_14361);
nand U22674 (N_22674,N_14606,N_17286);
nand U22675 (N_22675,N_14262,N_15121);
or U22676 (N_22676,N_17485,N_17374);
nand U22677 (N_22677,N_17198,N_14005);
or U22678 (N_22678,N_17225,N_18541);
nand U22679 (N_22679,N_12506,N_13113);
nor U22680 (N_22680,N_14260,N_16688);
nor U22681 (N_22681,N_17106,N_15673);
or U22682 (N_22682,N_12794,N_16734);
nor U22683 (N_22683,N_16805,N_14655);
or U22684 (N_22684,N_14199,N_14741);
nor U22685 (N_22685,N_12520,N_14973);
nor U22686 (N_22686,N_16204,N_14878);
and U22687 (N_22687,N_18061,N_15525);
nand U22688 (N_22688,N_15028,N_15133);
or U22689 (N_22689,N_14690,N_16447);
and U22690 (N_22690,N_15582,N_16800);
nor U22691 (N_22691,N_12837,N_14069);
or U22692 (N_22692,N_14710,N_13336);
nor U22693 (N_22693,N_17782,N_15087);
nor U22694 (N_22694,N_13874,N_18683);
xnor U22695 (N_22695,N_12546,N_15254);
nor U22696 (N_22696,N_15124,N_12534);
xor U22697 (N_22697,N_12529,N_14786);
nand U22698 (N_22698,N_14450,N_16692);
nand U22699 (N_22699,N_15746,N_17154);
or U22700 (N_22700,N_13312,N_12559);
nor U22701 (N_22701,N_17434,N_13769);
nor U22702 (N_22702,N_14718,N_18371);
nor U22703 (N_22703,N_13232,N_13208);
nor U22704 (N_22704,N_16913,N_12581);
nor U22705 (N_22705,N_14239,N_18320);
nand U22706 (N_22706,N_14022,N_16150);
nand U22707 (N_22707,N_15883,N_13453);
and U22708 (N_22708,N_18635,N_16676);
nor U22709 (N_22709,N_18356,N_14428);
or U22710 (N_22710,N_13272,N_16205);
or U22711 (N_22711,N_15526,N_16272);
and U22712 (N_22712,N_14456,N_15184);
or U22713 (N_22713,N_14409,N_15585);
and U22714 (N_22714,N_15599,N_16146);
and U22715 (N_22715,N_12976,N_17624);
nor U22716 (N_22716,N_14291,N_18423);
nor U22717 (N_22717,N_13838,N_12954);
and U22718 (N_22718,N_13780,N_17898);
nand U22719 (N_22719,N_17714,N_17625);
nor U22720 (N_22720,N_18308,N_17076);
nand U22721 (N_22721,N_18273,N_16113);
or U22722 (N_22722,N_18214,N_15294);
nand U22723 (N_22723,N_12784,N_14855);
or U22724 (N_22724,N_15879,N_15478);
nor U22725 (N_22725,N_16518,N_13699);
or U22726 (N_22726,N_16399,N_16913);
nor U22727 (N_22727,N_13313,N_12844);
or U22728 (N_22728,N_14668,N_14241);
and U22729 (N_22729,N_14096,N_16421);
and U22730 (N_22730,N_13342,N_13666);
nor U22731 (N_22731,N_17119,N_16577);
nand U22732 (N_22732,N_14345,N_16403);
or U22733 (N_22733,N_18509,N_17652);
or U22734 (N_22734,N_18448,N_17326);
and U22735 (N_22735,N_12749,N_17207);
nand U22736 (N_22736,N_17069,N_15925);
and U22737 (N_22737,N_18578,N_12851);
nor U22738 (N_22738,N_18619,N_12912);
nand U22739 (N_22739,N_14990,N_18018);
nor U22740 (N_22740,N_12732,N_15408);
or U22741 (N_22741,N_13889,N_17246);
or U22742 (N_22742,N_13413,N_13668);
and U22743 (N_22743,N_17463,N_16772);
nor U22744 (N_22744,N_15980,N_18707);
or U22745 (N_22745,N_17284,N_17763);
nand U22746 (N_22746,N_14611,N_17625);
nand U22747 (N_22747,N_15278,N_13147);
nand U22748 (N_22748,N_17946,N_15832);
nand U22749 (N_22749,N_17142,N_13167);
or U22750 (N_22750,N_18743,N_18286);
and U22751 (N_22751,N_15444,N_14287);
nand U22752 (N_22752,N_13252,N_15170);
nor U22753 (N_22753,N_17665,N_15228);
or U22754 (N_22754,N_12728,N_16680);
and U22755 (N_22755,N_17517,N_16071);
nand U22756 (N_22756,N_17343,N_17060);
and U22757 (N_22757,N_18529,N_12723);
or U22758 (N_22758,N_13315,N_17626);
and U22759 (N_22759,N_13562,N_14584);
nand U22760 (N_22760,N_15788,N_14322);
nor U22761 (N_22761,N_18573,N_13129);
nand U22762 (N_22762,N_18743,N_18398);
and U22763 (N_22763,N_15542,N_15816);
and U22764 (N_22764,N_17111,N_17047);
nor U22765 (N_22765,N_17379,N_14742);
nand U22766 (N_22766,N_18190,N_18714);
nand U22767 (N_22767,N_17857,N_15053);
nor U22768 (N_22768,N_13984,N_15735);
nor U22769 (N_22769,N_15221,N_17995);
and U22770 (N_22770,N_13825,N_13567);
and U22771 (N_22771,N_15565,N_17932);
nor U22772 (N_22772,N_18012,N_16453);
and U22773 (N_22773,N_13280,N_12749);
nor U22774 (N_22774,N_13492,N_15337);
nand U22775 (N_22775,N_17887,N_13153);
nand U22776 (N_22776,N_17914,N_12912);
or U22777 (N_22777,N_18626,N_16239);
nand U22778 (N_22778,N_15378,N_14541);
and U22779 (N_22779,N_17395,N_18035);
or U22780 (N_22780,N_17877,N_17423);
or U22781 (N_22781,N_16855,N_12902);
and U22782 (N_22782,N_18039,N_16448);
nor U22783 (N_22783,N_14505,N_15548);
nand U22784 (N_22784,N_16358,N_16860);
nor U22785 (N_22785,N_13581,N_17445);
or U22786 (N_22786,N_16409,N_18251);
nor U22787 (N_22787,N_18117,N_16991);
nor U22788 (N_22788,N_15794,N_15245);
nor U22789 (N_22789,N_15468,N_18629);
or U22790 (N_22790,N_14867,N_18568);
and U22791 (N_22791,N_13776,N_13542);
or U22792 (N_22792,N_17145,N_15310);
nand U22793 (N_22793,N_16577,N_13557);
nand U22794 (N_22794,N_15311,N_12929);
and U22795 (N_22795,N_15694,N_16384);
or U22796 (N_22796,N_14974,N_15382);
nand U22797 (N_22797,N_17442,N_14160);
and U22798 (N_22798,N_17365,N_13938);
nor U22799 (N_22799,N_13665,N_18714);
nand U22800 (N_22800,N_13818,N_16386);
and U22801 (N_22801,N_18575,N_16955);
nand U22802 (N_22802,N_15750,N_16811);
nor U22803 (N_22803,N_13345,N_16278);
nor U22804 (N_22804,N_17543,N_16930);
or U22805 (N_22805,N_15524,N_17543);
and U22806 (N_22806,N_12568,N_16611);
or U22807 (N_22807,N_15984,N_13302);
nand U22808 (N_22808,N_12666,N_15729);
xor U22809 (N_22809,N_17146,N_17261);
or U22810 (N_22810,N_18024,N_17433);
nand U22811 (N_22811,N_13728,N_16507);
nor U22812 (N_22812,N_18392,N_13867);
and U22813 (N_22813,N_13868,N_12966);
and U22814 (N_22814,N_18071,N_16754);
and U22815 (N_22815,N_18162,N_14074);
nor U22816 (N_22816,N_17207,N_17650);
nand U22817 (N_22817,N_17139,N_16983);
and U22818 (N_22818,N_12828,N_13881);
nor U22819 (N_22819,N_15551,N_12923);
nand U22820 (N_22820,N_18717,N_14499);
or U22821 (N_22821,N_15151,N_14412);
and U22822 (N_22822,N_18703,N_17794);
nor U22823 (N_22823,N_13127,N_16866);
nor U22824 (N_22824,N_13189,N_13728);
and U22825 (N_22825,N_18105,N_17035);
or U22826 (N_22826,N_15446,N_17494);
and U22827 (N_22827,N_15301,N_18092);
and U22828 (N_22828,N_17167,N_17242);
nand U22829 (N_22829,N_17546,N_18155);
or U22830 (N_22830,N_15119,N_18499);
or U22831 (N_22831,N_17813,N_13842);
nand U22832 (N_22832,N_13545,N_13483);
and U22833 (N_22833,N_14680,N_17505);
and U22834 (N_22834,N_17080,N_17488);
nand U22835 (N_22835,N_16450,N_14029);
or U22836 (N_22836,N_14994,N_15871);
nand U22837 (N_22837,N_17081,N_14984);
nand U22838 (N_22838,N_16609,N_17620);
and U22839 (N_22839,N_14671,N_14338);
nor U22840 (N_22840,N_13774,N_16315);
nor U22841 (N_22841,N_14421,N_16570);
nand U22842 (N_22842,N_18574,N_16602);
and U22843 (N_22843,N_17361,N_16776);
and U22844 (N_22844,N_17161,N_17962);
and U22845 (N_22845,N_14369,N_12515);
nand U22846 (N_22846,N_14515,N_16755);
or U22847 (N_22847,N_15257,N_17804);
nor U22848 (N_22848,N_13158,N_14119);
xor U22849 (N_22849,N_13467,N_15579);
or U22850 (N_22850,N_13506,N_18173);
nor U22851 (N_22851,N_16058,N_12740);
and U22852 (N_22852,N_14021,N_15006);
nand U22853 (N_22853,N_16182,N_17912);
nor U22854 (N_22854,N_13354,N_18411);
or U22855 (N_22855,N_17075,N_14063);
or U22856 (N_22856,N_17408,N_16186);
nor U22857 (N_22857,N_13548,N_15423);
nand U22858 (N_22858,N_16440,N_12647);
nor U22859 (N_22859,N_17668,N_15371);
and U22860 (N_22860,N_18609,N_18188);
nor U22861 (N_22861,N_17026,N_16614);
and U22862 (N_22862,N_18514,N_14603);
or U22863 (N_22863,N_13735,N_16579);
or U22864 (N_22864,N_17462,N_14993);
or U22865 (N_22865,N_14813,N_17693);
nand U22866 (N_22866,N_18688,N_15818);
and U22867 (N_22867,N_17052,N_15435);
nand U22868 (N_22868,N_16397,N_16649);
and U22869 (N_22869,N_12992,N_12544);
and U22870 (N_22870,N_17911,N_18596);
and U22871 (N_22871,N_18644,N_12709);
and U22872 (N_22872,N_13740,N_13139);
or U22873 (N_22873,N_14004,N_18142);
and U22874 (N_22874,N_15680,N_12678);
nor U22875 (N_22875,N_14668,N_18389);
nor U22876 (N_22876,N_16620,N_13141);
nand U22877 (N_22877,N_17924,N_14162);
and U22878 (N_22878,N_14345,N_18676);
nor U22879 (N_22879,N_14784,N_16615);
nor U22880 (N_22880,N_14431,N_12619);
nand U22881 (N_22881,N_16189,N_14336);
or U22882 (N_22882,N_16690,N_17570);
or U22883 (N_22883,N_18113,N_13581);
or U22884 (N_22884,N_16614,N_17396);
and U22885 (N_22885,N_16297,N_14389);
nand U22886 (N_22886,N_17653,N_18423);
nand U22887 (N_22887,N_16372,N_17537);
nor U22888 (N_22888,N_16914,N_16463);
or U22889 (N_22889,N_18327,N_14740);
and U22890 (N_22890,N_13395,N_13869);
nand U22891 (N_22891,N_15425,N_18598);
xnor U22892 (N_22892,N_15809,N_16149);
and U22893 (N_22893,N_13405,N_12550);
nand U22894 (N_22894,N_14679,N_13009);
nor U22895 (N_22895,N_16103,N_15089);
nand U22896 (N_22896,N_13553,N_17085);
and U22897 (N_22897,N_18411,N_18379);
nand U22898 (N_22898,N_16541,N_14423);
nand U22899 (N_22899,N_14803,N_17329);
nand U22900 (N_22900,N_14215,N_16779);
and U22901 (N_22901,N_15667,N_18691);
or U22902 (N_22902,N_15847,N_12632);
or U22903 (N_22903,N_17900,N_16624);
nand U22904 (N_22904,N_14860,N_12782);
nand U22905 (N_22905,N_14259,N_13358);
nor U22906 (N_22906,N_14482,N_13985);
nor U22907 (N_22907,N_16864,N_14009);
and U22908 (N_22908,N_14318,N_16302);
and U22909 (N_22909,N_12722,N_15029);
and U22910 (N_22910,N_16491,N_15438);
and U22911 (N_22911,N_16994,N_13166);
or U22912 (N_22912,N_16482,N_13379);
or U22913 (N_22913,N_18115,N_14825);
or U22914 (N_22914,N_13953,N_16137);
or U22915 (N_22915,N_17370,N_14117);
nor U22916 (N_22916,N_12583,N_14500);
xor U22917 (N_22917,N_13757,N_13979);
nand U22918 (N_22918,N_17690,N_15918);
and U22919 (N_22919,N_15613,N_13522);
or U22920 (N_22920,N_13577,N_15013);
or U22921 (N_22921,N_17795,N_14555);
and U22922 (N_22922,N_18429,N_14845);
or U22923 (N_22923,N_15741,N_17126);
nor U22924 (N_22924,N_13570,N_18614);
nor U22925 (N_22925,N_14104,N_15271);
nor U22926 (N_22926,N_12580,N_13341);
or U22927 (N_22927,N_17835,N_18037);
nor U22928 (N_22928,N_15240,N_13698);
or U22929 (N_22929,N_17094,N_17633);
and U22930 (N_22930,N_15231,N_13732);
or U22931 (N_22931,N_17669,N_17343);
xnor U22932 (N_22932,N_17848,N_17849);
and U22933 (N_22933,N_18173,N_18224);
or U22934 (N_22934,N_12732,N_16216);
nor U22935 (N_22935,N_14266,N_14954);
nand U22936 (N_22936,N_12757,N_18656);
nand U22937 (N_22937,N_13064,N_14754);
and U22938 (N_22938,N_16869,N_12613);
or U22939 (N_22939,N_15197,N_12785);
or U22940 (N_22940,N_15418,N_13174);
or U22941 (N_22941,N_16821,N_18297);
nand U22942 (N_22942,N_14818,N_14950);
and U22943 (N_22943,N_18350,N_14635);
nand U22944 (N_22944,N_14020,N_17500);
and U22945 (N_22945,N_16684,N_17572);
nor U22946 (N_22946,N_12554,N_16159);
nand U22947 (N_22947,N_16360,N_14929);
or U22948 (N_22948,N_18723,N_13739);
and U22949 (N_22949,N_14588,N_17356);
nand U22950 (N_22950,N_13693,N_13912);
or U22951 (N_22951,N_13818,N_16312);
and U22952 (N_22952,N_17709,N_17356);
nor U22953 (N_22953,N_14924,N_12619);
or U22954 (N_22954,N_18292,N_15317);
and U22955 (N_22955,N_18464,N_17710);
nor U22956 (N_22956,N_15295,N_16510);
nor U22957 (N_22957,N_17564,N_16989);
nand U22958 (N_22958,N_18543,N_18541);
or U22959 (N_22959,N_17249,N_17758);
and U22960 (N_22960,N_18253,N_14400);
nor U22961 (N_22961,N_15740,N_14907);
nor U22962 (N_22962,N_15831,N_13271);
or U22963 (N_22963,N_14255,N_17841);
xnor U22964 (N_22964,N_17192,N_17877);
nand U22965 (N_22965,N_13690,N_14796);
xnor U22966 (N_22966,N_14636,N_15436);
nand U22967 (N_22967,N_14639,N_12863);
and U22968 (N_22968,N_13607,N_17903);
nor U22969 (N_22969,N_17638,N_15280);
and U22970 (N_22970,N_17192,N_15479);
nand U22971 (N_22971,N_18653,N_16642);
nand U22972 (N_22972,N_17246,N_18431);
nor U22973 (N_22973,N_17664,N_13178);
or U22974 (N_22974,N_14692,N_16645);
or U22975 (N_22975,N_13717,N_16562);
xor U22976 (N_22976,N_17208,N_15742);
nor U22977 (N_22977,N_13031,N_18179);
and U22978 (N_22978,N_12839,N_16682);
or U22979 (N_22979,N_16547,N_12896);
and U22980 (N_22980,N_17964,N_15999);
or U22981 (N_22981,N_16687,N_16954);
nand U22982 (N_22982,N_13635,N_15533);
and U22983 (N_22983,N_15454,N_16150);
nand U22984 (N_22984,N_15881,N_14565);
nor U22985 (N_22985,N_13133,N_14742);
or U22986 (N_22986,N_15596,N_14830);
nand U22987 (N_22987,N_17037,N_14230);
nor U22988 (N_22988,N_13870,N_16231);
or U22989 (N_22989,N_15646,N_17511);
nand U22990 (N_22990,N_16165,N_17661);
nand U22991 (N_22991,N_18016,N_14052);
nor U22992 (N_22992,N_13926,N_16685);
or U22993 (N_22993,N_13972,N_16157);
nor U22994 (N_22994,N_15931,N_14518);
nand U22995 (N_22995,N_13041,N_15350);
nand U22996 (N_22996,N_18201,N_16384);
nor U22997 (N_22997,N_13673,N_16303);
nand U22998 (N_22998,N_14027,N_15818);
and U22999 (N_22999,N_14190,N_14603);
or U23000 (N_23000,N_16595,N_14442);
nor U23001 (N_23001,N_14728,N_15904);
nor U23002 (N_23002,N_18009,N_13127);
or U23003 (N_23003,N_17480,N_14457);
and U23004 (N_23004,N_13894,N_14275);
and U23005 (N_23005,N_14265,N_18650);
or U23006 (N_23006,N_15921,N_18316);
and U23007 (N_23007,N_13763,N_18139);
nor U23008 (N_23008,N_18469,N_17232);
nand U23009 (N_23009,N_18530,N_15357);
and U23010 (N_23010,N_17931,N_16442);
nand U23011 (N_23011,N_17613,N_13473);
or U23012 (N_23012,N_16830,N_17537);
nor U23013 (N_23013,N_18177,N_17825);
nand U23014 (N_23014,N_12930,N_16229);
or U23015 (N_23015,N_16086,N_17094);
nor U23016 (N_23016,N_13043,N_13539);
or U23017 (N_23017,N_17871,N_18152);
or U23018 (N_23018,N_14761,N_15769);
nand U23019 (N_23019,N_12821,N_17920);
nand U23020 (N_23020,N_12769,N_17416);
or U23021 (N_23021,N_13788,N_14526);
nand U23022 (N_23022,N_18446,N_16730);
nor U23023 (N_23023,N_17965,N_17092);
and U23024 (N_23024,N_17519,N_18018);
nor U23025 (N_23025,N_16227,N_16369);
or U23026 (N_23026,N_17721,N_17120);
nor U23027 (N_23027,N_13232,N_15451);
and U23028 (N_23028,N_12673,N_13734);
and U23029 (N_23029,N_13897,N_16602);
or U23030 (N_23030,N_15367,N_12507);
and U23031 (N_23031,N_17524,N_15829);
or U23032 (N_23032,N_14450,N_12770);
or U23033 (N_23033,N_16159,N_18014);
nand U23034 (N_23034,N_15864,N_17069);
and U23035 (N_23035,N_17056,N_15295);
nand U23036 (N_23036,N_16562,N_14987);
or U23037 (N_23037,N_15888,N_14788);
and U23038 (N_23038,N_16934,N_14131);
or U23039 (N_23039,N_15239,N_16897);
nand U23040 (N_23040,N_17383,N_16625);
nand U23041 (N_23041,N_15077,N_14019);
nor U23042 (N_23042,N_17945,N_17244);
and U23043 (N_23043,N_16946,N_13013);
and U23044 (N_23044,N_13567,N_17187);
nor U23045 (N_23045,N_13177,N_13544);
or U23046 (N_23046,N_18371,N_15528);
nor U23047 (N_23047,N_12739,N_16506);
and U23048 (N_23048,N_18648,N_14302);
nor U23049 (N_23049,N_14387,N_14152);
nand U23050 (N_23050,N_15303,N_16085);
nand U23051 (N_23051,N_18308,N_14343);
and U23052 (N_23052,N_17889,N_15810);
nand U23053 (N_23053,N_15108,N_12844);
and U23054 (N_23054,N_16915,N_17707);
and U23055 (N_23055,N_13490,N_13683);
and U23056 (N_23056,N_14964,N_15694);
nand U23057 (N_23057,N_15837,N_16365);
or U23058 (N_23058,N_16177,N_16712);
or U23059 (N_23059,N_14397,N_18249);
nand U23060 (N_23060,N_18300,N_12746);
nor U23061 (N_23061,N_17680,N_18148);
or U23062 (N_23062,N_15184,N_15889);
nor U23063 (N_23063,N_14378,N_15009);
nand U23064 (N_23064,N_12673,N_14414);
and U23065 (N_23065,N_13248,N_18387);
or U23066 (N_23066,N_16043,N_14064);
or U23067 (N_23067,N_15454,N_16401);
nor U23068 (N_23068,N_16180,N_14212);
nor U23069 (N_23069,N_15357,N_18589);
nor U23070 (N_23070,N_17868,N_18426);
nor U23071 (N_23071,N_15633,N_16897);
nand U23072 (N_23072,N_13382,N_13807);
and U23073 (N_23073,N_13122,N_17229);
nor U23074 (N_23074,N_12972,N_16591);
and U23075 (N_23075,N_15428,N_14752);
nand U23076 (N_23076,N_15005,N_17457);
nor U23077 (N_23077,N_15666,N_14683);
nor U23078 (N_23078,N_17200,N_17632);
or U23079 (N_23079,N_14841,N_14874);
and U23080 (N_23080,N_15956,N_17421);
nor U23081 (N_23081,N_17502,N_16809);
or U23082 (N_23082,N_18524,N_14191);
and U23083 (N_23083,N_16122,N_17447);
and U23084 (N_23084,N_15303,N_15810);
nor U23085 (N_23085,N_15005,N_12746);
and U23086 (N_23086,N_14959,N_16174);
and U23087 (N_23087,N_13615,N_18034);
nor U23088 (N_23088,N_17433,N_18736);
nor U23089 (N_23089,N_14592,N_13413);
or U23090 (N_23090,N_16174,N_16200);
or U23091 (N_23091,N_15245,N_14956);
nand U23092 (N_23092,N_17508,N_16308);
nand U23093 (N_23093,N_18671,N_14313);
nand U23094 (N_23094,N_16486,N_16094);
or U23095 (N_23095,N_18505,N_16047);
nor U23096 (N_23096,N_15480,N_17463);
nand U23097 (N_23097,N_17083,N_15385);
nand U23098 (N_23098,N_17862,N_17578);
xnor U23099 (N_23099,N_12729,N_18629);
or U23100 (N_23100,N_16364,N_17254);
nand U23101 (N_23101,N_14458,N_18183);
nand U23102 (N_23102,N_15080,N_14159);
nor U23103 (N_23103,N_17354,N_16184);
nor U23104 (N_23104,N_13072,N_14539);
nand U23105 (N_23105,N_15121,N_14924);
or U23106 (N_23106,N_17117,N_18488);
or U23107 (N_23107,N_18182,N_15320);
or U23108 (N_23108,N_16904,N_16591);
and U23109 (N_23109,N_17229,N_13549);
nor U23110 (N_23110,N_15766,N_17807);
nor U23111 (N_23111,N_14216,N_13716);
nand U23112 (N_23112,N_18354,N_13781);
nor U23113 (N_23113,N_17520,N_17107);
xor U23114 (N_23114,N_17620,N_15766);
nand U23115 (N_23115,N_14066,N_16718);
nor U23116 (N_23116,N_18278,N_18218);
nand U23117 (N_23117,N_15577,N_16483);
nor U23118 (N_23118,N_16036,N_17140);
nor U23119 (N_23119,N_15330,N_12592);
and U23120 (N_23120,N_15448,N_14143);
or U23121 (N_23121,N_13358,N_15644);
nand U23122 (N_23122,N_16706,N_17921);
nand U23123 (N_23123,N_17463,N_17201);
and U23124 (N_23124,N_18634,N_13084);
and U23125 (N_23125,N_15623,N_14126);
nor U23126 (N_23126,N_15731,N_18017);
and U23127 (N_23127,N_13315,N_16855);
or U23128 (N_23128,N_15724,N_13749);
nand U23129 (N_23129,N_16477,N_14689);
nor U23130 (N_23130,N_16111,N_16762);
or U23131 (N_23131,N_15541,N_17381);
and U23132 (N_23132,N_18668,N_17160);
nand U23133 (N_23133,N_16352,N_16952);
or U23134 (N_23134,N_14076,N_12847);
or U23135 (N_23135,N_18347,N_18296);
nor U23136 (N_23136,N_16159,N_15011);
nand U23137 (N_23137,N_14498,N_18031);
and U23138 (N_23138,N_13340,N_14267);
nor U23139 (N_23139,N_17797,N_14078);
nor U23140 (N_23140,N_16950,N_18465);
and U23141 (N_23141,N_16181,N_15006);
nand U23142 (N_23142,N_15877,N_12897);
nand U23143 (N_23143,N_14730,N_15113);
nand U23144 (N_23144,N_14981,N_14563);
nand U23145 (N_23145,N_16783,N_15706);
and U23146 (N_23146,N_15352,N_14732);
or U23147 (N_23147,N_15968,N_15199);
nand U23148 (N_23148,N_16424,N_16360);
or U23149 (N_23149,N_18418,N_15923);
or U23150 (N_23150,N_15667,N_18515);
or U23151 (N_23151,N_17589,N_13493);
or U23152 (N_23152,N_16899,N_15934);
or U23153 (N_23153,N_18573,N_18234);
nand U23154 (N_23154,N_13823,N_12533);
nor U23155 (N_23155,N_16854,N_13196);
nand U23156 (N_23156,N_13642,N_16054);
or U23157 (N_23157,N_16698,N_13077);
nor U23158 (N_23158,N_15240,N_13578);
and U23159 (N_23159,N_15010,N_14332);
nor U23160 (N_23160,N_15351,N_13170);
and U23161 (N_23161,N_15895,N_16556);
or U23162 (N_23162,N_16234,N_14065);
and U23163 (N_23163,N_17835,N_17335);
and U23164 (N_23164,N_14372,N_16312);
or U23165 (N_23165,N_16450,N_17721);
nor U23166 (N_23166,N_14576,N_12640);
or U23167 (N_23167,N_12596,N_17951);
nor U23168 (N_23168,N_14060,N_18719);
nand U23169 (N_23169,N_15250,N_16675);
or U23170 (N_23170,N_12806,N_14720);
and U23171 (N_23171,N_16947,N_14033);
or U23172 (N_23172,N_18280,N_18086);
or U23173 (N_23173,N_18499,N_15325);
or U23174 (N_23174,N_14120,N_14590);
nand U23175 (N_23175,N_17070,N_17883);
or U23176 (N_23176,N_14656,N_17738);
or U23177 (N_23177,N_18228,N_15667);
nor U23178 (N_23178,N_16323,N_17885);
nand U23179 (N_23179,N_15116,N_12762);
or U23180 (N_23180,N_16664,N_12707);
and U23181 (N_23181,N_15999,N_18401);
nand U23182 (N_23182,N_15460,N_15896);
nand U23183 (N_23183,N_17507,N_13844);
or U23184 (N_23184,N_13151,N_13527);
or U23185 (N_23185,N_16838,N_17346);
nand U23186 (N_23186,N_16435,N_15801);
nor U23187 (N_23187,N_15919,N_17935);
or U23188 (N_23188,N_18397,N_16451);
and U23189 (N_23189,N_16397,N_16531);
or U23190 (N_23190,N_14926,N_17664);
nor U23191 (N_23191,N_16739,N_15911);
and U23192 (N_23192,N_17364,N_18441);
nor U23193 (N_23193,N_16149,N_12534);
or U23194 (N_23194,N_18438,N_14015);
nor U23195 (N_23195,N_17209,N_12588);
nand U23196 (N_23196,N_14364,N_15417);
and U23197 (N_23197,N_14116,N_15131);
or U23198 (N_23198,N_14451,N_14994);
nand U23199 (N_23199,N_15970,N_14155);
xor U23200 (N_23200,N_14265,N_17563);
and U23201 (N_23201,N_15154,N_16712);
nand U23202 (N_23202,N_17513,N_17163);
and U23203 (N_23203,N_18332,N_14250);
nand U23204 (N_23204,N_18208,N_16124);
or U23205 (N_23205,N_17205,N_18578);
nor U23206 (N_23206,N_16943,N_14925);
nand U23207 (N_23207,N_13551,N_17040);
or U23208 (N_23208,N_14139,N_17555);
and U23209 (N_23209,N_14479,N_13543);
nor U23210 (N_23210,N_13900,N_17687);
nand U23211 (N_23211,N_13489,N_14949);
nor U23212 (N_23212,N_15816,N_17745);
nor U23213 (N_23213,N_18552,N_12831);
and U23214 (N_23214,N_12673,N_18227);
nor U23215 (N_23215,N_17225,N_15779);
nand U23216 (N_23216,N_15251,N_14425);
nor U23217 (N_23217,N_15106,N_13882);
or U23218 (N_23218,N_12823,N_17017);
nor U23219 (N_23219,N_13550,N_17664);
nor U23220 (N_23220,N_13190,N_17350);
nand U23221 (N_23221,N_17563,N_16377);
nor U23222 (N_23222,N_16074,N_17660);
xor U23223 (N_23223,N_17933,N_12936);
and U23224 (N_23224,N_18083,N_15152);
nand U23225 (N_23225,N_14659,N_13325);
nor U23226 (N_23226,N_12728,N_16983);
nand U23227 (N_23227,N_14423,N_13691);
or U23228 (N_23228,N_12635,N_17983);
nand U23229 (N_23229,N_15375,N_14425);
nand U23230 (N_23230,N_15857,N_17419);
xor U23231 (N_23231,N_12546,N_17065);
nand U23232 (N_23232,N_13577,N_15323);
or U23233 (N_23233,N_13236,N_17900);
nor U23234 (N_23234,N_17153,N_13093);
and U23235 (N_23235,N_16912,N_16134);
nand U23236 (N_23236,N_14899,N_16873);
and U23237 (N_23237,N_12702,N_13902);
nand U23238 (N_23238,N_17580,N_17238);
and U23239 (N_23239,N_15333,N_12916);
nand U23240 (N_23240,N_12874,N_15901);
xor U23241 (N_23241,N_17325,N_13002);
nand U23242 (N_23242,N_17379,N_15861);
or U23243 (N_23243,N_13204,N_14087);
nor U23244 (N_23244,N_13300,N_14880);
nand U23245 (N_23245,N_17917,N_13036);
nand U23246 (N_23246,N_16437,N_15069);
and U23247 (N_23247,N_14932,N_17231);
or U23248 (N_23248,N_17729,N_12551);
or U23249 (N_23249,N_14643,N_15567);
and U23250 (N_23250,N_18099,N_14224);
and U23251 (N_23251,N_13062,N_14300);
or U23252 (N_23252,N_15414,N_15709);
and U23253 (N_23253,N_14096,N_17214);
nor U23254 (N_23254,N_13835,N_14510);
nand U23255 (N_23255,N_14830,N_14656);
and U23256 (N_23256,N_15449,N_17826);
or U23257 (N_23257,N_15999,N_17459);
and U23258 (N_23258,N_16551,N_17923);
nor U23259 (N_23259,N_17196,N_16557);
or U23260 (N_23260,N_18342,N_16878);
or U23261 (N_23261,N_13777,N_16198);
nor U23262 (N_23262,N_15188,N_13350);
and U23263 (N_23263,N_16088,N_18550);
or U23264 (N_23264,N_14129,N_15938);
nor U23265 (N_23265,N_16163,N_15859);
nand U23266 (N_23266,N_16640,N_17460);
and U23267 (N_23267,N_14813,N_15581);
nor U23268 (N_23268,N_15342,N_16414);
nand U23269 (N_23269,N_15457,N_13751);
nand U23270 (N_23270,N_13344,N_12963);
nand U23271 (N_23271,N_13160,N_14544);
nor U23272 (N_23272,N_17951,N_14119);
and U23273 (N_23273,N_17102,N_15990);
and U23274 (N_23274,N_16698,N_13147);
nor U23275 (N_23275,N_17621,N_12868);
nor U23276 (N_23276,N_13223,N_14559);
and U23277 (N_23277,N_12516,N_15055);
nor U23278 (N_23278,N_17363,N_17063);
and U23279 (N_23279,N_13735,N_13277);
and U23280 (N_23280,N_18391,N_13604);
or U23281 (N_23281,N_14812,N_13168);
nand U23282 (N_23282,N_18405,N_13603);
nor U23283 (N_23283,N_13552,N_12527);
nand U23284 (N_23284,N_14873,N_17653);
nor U23285 (N_23285,N_14170,N_18335);
nor U23286 (N_23286,N_17160,N_14294);
or U23287 (N_23287,N_17993,N_18682);
nand U23288 (N_23288,N_13397,N_18585);
nor U23289 (N_23289,N_16326,N_14711);
or U23290 (N_23290,N_15812,N_14227);
and U23291 (N_23291,N_15850,N_14794);
nor U23292 (N_23292,N_16042,N_14124);
nand U23293 (N_23293,N_12701,N_18742);
and U23294 (N_23294,N_17395,N_17268);
or U23295 (N_23295,N_17253,N_16926);
nor U23296 (N_23296,N_18097,N_15190);
and U23297 (N_23297,N_15694,N_18100);
or U23298 (N_23298,N_18118,N_15349);
or U23299 (N_23299,N_16202,N_14108);
and U23300 (N_23300,N_14223,N_16809);
nor U23301 (N_23301,N_15638,N_16646);
and U23302 (N_23302,N_13349,N_13177);
and U23303 (N_23303,N_16526,N_14496);
nor U23304 (N_23304,N_17064,N_16560);
nor U23305 (N_23305,N_14938,N_15274);
and U23306 (N_23306,N_18361,N_18572);
or U23307 (N_23307,N_16580,N_14172);
nand U23308 (N_23308,N_16719,N_14511);
nand U23309 (N_23309,N_15812,N_14295);
and U23310 (N_23310,N_12876,N_14310);
or U23311 (N_23311,N_15231,N_17101);
nor U23312 (N_23312,N_14351,N_17502);
xnor U23313 (N_23313,N_13302,N_15473);
or U23314 (N_23314,N_15958,N_17460);
or U23315 (N_23315,N_18155,N_13167);
nor U23316 (N_23316,N_14043,N_16884);
nand U23317 (N_23317,N_14278,N_14484);
or U23318 (N_23318,N_15644,N_15758);
nor U23319 (N_23319,N_14173,N_17807);
or U23320 (N_23320,N_18566,N_17646);
nand U23321 (N_23321,N_14519,N_18494);
or U23322 (N_23322,N_12548,N_17707);
or U23323 (N_23323,N_17406,N_16702);
nand U23324 (N_23324,N_12806,N_17601);
and U23325 (N_23325,N_16502,N_17967);
and U23326 (N_23326,N_17288,N_16111);
and U23327 (N_23327,N_16555,N_17210);
or U23328 (N_23328,N_14273,N_18542);
or U23329 (N_23329,N_15869,N_17399);
and U23330 (N_23330,N_14296,N_17201);
nand U23331 (N_23331,N_16626,N_16846);
nor U23332 (N_23332,N_16180,N_15551);
and U23333 (N_23333,N_18199,N_14098);
and U23334 (N_23334,N_18633,N_14538);
or U23335 (N_23335,N_17999,N_12804);
nor U23336 (N_23336,N_17527,N_16665);
and U23337 (N_23337,N_16244,N_15245);
or U23338 (N_23338,N_12548,N_18229);
nor U23339 (N_23339,N_16023,N_17367);
nand U23340 (N_23340,N_17782,N_18594);
nand U23341 (N_23341,N_16337,N_18258);
nor U23342 (N_23342,N_16988,N_17246);
or U23343 (N_23343,N_15631,N_13790);
nor U23344 (N_23344,N_17967,N_14043);
and U23345 (N_23345,N_17553,N_14037);
nand U23346 (N_23346,N_17155,N_15741);
and U23347 (N_23347,N_15888,N_12989);
nor U23348 (N_23348,N_15895,N_14230);
nor U23349 (N_23349,N_15684,N_13993);
or U23350 (N_23350,N_14194,N_13514);
or U23351 (N_23351,N_14861,N_18196);
or U23352 (N_23352,N_14456,N_18605);
and U23353 (N_23353,N_18384,N_14530);
and U23354 (N_23354,N_15302,N_18293);
nor U23355 (N_23355,N_17475,N_18374);
nor U23356 (N_23356,N_13924,N_17948);
and U23357 (N_23357,N_18579,N_13072);
nor U23358 (N_23358,N_14968,N_14237);
nor U23359 (N_23359,N_17373,N_13053);
or U23360 (N_23360,N_18710,N_17056);
or U23361 (N_23361,N_15054,N_16192);
nand U23362 (N_23362,N_17481,N_14431);
nor U23363 (N_23363,N_18674,N_18340);
and U23364 (N_23364,N_15750,N_13716);
nor U23365 (N_23365,N_15957,N_17634);
and U23366 (N_23366,N_13607,N_17157);
or U23367 (N_23367,N_13698,N_16549);
nand U23368 (N_23368,N_16659,N_16175);
or U23369 (N_23369,N_18620,N_17025);
nor U23370 (N_23370,N_16051,N_16236);
or U23371 (N_23371,N_15506,N_18238);
or U23372 (N_23372,N_14333,N_17221);
nor U23373 (N_23373,N_12632,N_14831);
and U23374 (N_23374,N_14539,N_13320);
and U23375 (N_23375,N_17432,N_13452);
or U23376 (N_23376,N_12602,N_15132);
nor U23377 (N_23377,N_17995,N_18257);
or U23378 (N_23378,N_16446,N_17855);
or U23379 (N_23379,N_17649,N_14113);
nor U23380 (N_23380,N_14288,N_14691);
and U23381 (N_23381,N_14848,N_14182);
nand U23382 (N_23382,N_18530,N_14744);
or U23383 (N_23383,N_15156,N_14790);
or U23384 (N_23384,N_14612,N_14331);
and U23385 (N_23385,N_12616,N_15606);
nor U23386 (N_23386,N_15385,N_17790);
and U23387 (N_23387,N_15593,N_16615);
or U23388 (N_23388,N_15719,N_15112);
nand U23389 (N_23389,N_13758,N_16566);
nand U23390 (N_23390,N_16289,N_15373);
nor U23391 (N_23391,N_15400,N_16854);
nor U23392 (N_23392,N_17449,N_16956);
or U23393 (N_23393,N_15843,N_17011);
nand U23394 (N_23394,N_17061,N_17050);
and U23395 (N_23395,N_14875,N_12972);
nor U23396 (N_23396,N_16341,N_15987);
nor U23397 (N_23397,N_13547,N_16019);
and U23398 (N_23398,N_14305,N_12967);
and U23399 (N_23399,N_12916,N_12904);
nand U23400 (N_23400,N_16676,N_14548);
nand U23401 (N_23401,N_17955,N_13388);
and U23402 (N_23402,N_17931,N_18149);
or U23403 (N_23403,N_13954,N_17694);
nor U23404 (N_23404,N_13574,N_15197);
nor U23405 (N_23405,N_18660,N_16677);
and U23406 (N_23406,N_15283,N_12604);
or U23407 (N_23407,N_18433,N_15200);
nor U23408 (N_23408,N_16460,N_17291);
nand U23409 (N_23409,N_13308,N_14412);
and U23410 (N_23410,N_13920,N_16085);
nor U23411 (N_23411,N_17507,N_16831);
nor U23412 (N_23412,N_14726,N_14880);
and U23413 (N_23413,N_18167,N_15949);
and U23414 (N_23414,N_18287,N_12771);
nand U23415 (N_23415,N_17058,N_15455);
nor U23416 (N_23416,N_13383,N_14181);
or U23417 (N_23417,N_13378,N_15642);
nor U23418 (N_23418,N_18275,N_16762);
nand U23419 (N_23419,N_14325,N_15676);
nand U23420 (N_23420,N_17675,N_17721);
nand U23421 (N_23421,N_17613,N_15244);
or U23422 (N_23422,N_15460,N_17133);
and U23423 (N_23423,N_14272,N_18674);
and U23424 (N_23424,N_15871,N_13175);
and U23425 (N_23425,N_12865,N_13387);
nor U23426 (N_23426,N_14465,N_17679);
nand U23427 (N_23427,N_18112,N_17119);
or U23428 (N_23428,N_13202,N_15389);
or U23429 (N_23429,N_12925,N_15818);
or U23430 (N_23430,N_14489,N_14441);
nor U23431 (N_23431,N_15681,N_12568);
or U23432 (N_23432,N_15833,N_12790);
nor U23433 (N_23433,N_13184,N_18417);
and U23434 (N_23434,N_18188,N_16198);
or U23435 (N_23435,N_14361,N_16187);
or U23436 (N_23436,N_16205,N_14202);
nor U23437 (N_23437,N_16924,N_15085);
or U23438 (N_23438,N_13394,N_18159);
and U23439 (N_23439,N_14996,N_14548);
nand U23440 (N_23440,N_17971,N_16842);
or U23441 (N_23441,N_17592,N_13984);
nand U23442 (N_23442,N_14632,N_15890);
and U23443 (N_23443,N_16908,N_13612);
nand U23444 (N_23444,N_15855,N_18671);
and U23445 (N_23445,N_17959,N_14134);
or U23446 (N_23446,N_15947,N_13914);
and U23447 (N_23447,N_12823,N_15671);
nand U23448 (N_23448,N_13237,N_15600);
or U23449 (N_23449,N_13670,N_12524);
nor U23450 (N_23450,N_13108,N_14167);
or U23451 (N_23451,N_13532,N_13876);
and U23452 (N_23452,N_13075,N_16031);
and U23453 (N_23453,N_16143,N_18354);
nand U23454 (N_23454,N_13288,N_12742);
nor U23455 (N_23455,N_15232,N_16701);
nor U23456 (N_23456,N_13522,N_14165);
xnor U23457 (N_23457,N_17914,N_15340);
nand U23458 (N_23458,N_13972,N_16245);
or U23459 (N_23459,N_18301,N_14194);
or U23460 (N_23460,N_17295,N_17261);
or U23461 (N_23461,N_17727,N_15720);
or U23462 (N_23462,N_17963,N_17748);
and U23463 (N_23463,N_17877,N_14825);
nand U23464 (N_23464,N_14308,N_14724);
and U23465 (N_23465,N_15649,N_15977);
or U23466 (N_23466,N_17512,N_17084);
and U23467 (N_23467,N_16021,N_15789);
or U23468 (N_23468,N_13695,N_15647);
or U23469 (N_23469,N_12593,N_17014);
nor U23470 (N_23470,N_14120,N_18104);
nor U23471 (N_23471,N_14999,N_17094);
nand U23472 (N_23472,N_16907,N_14019);
and U23473 (N_23473,N_15301,N_16851);
nand U23474 (N_23474,N_16173,N_17352);
or U23475 (N_23475,N_16066,N_16276);
nor U23476 (N_23476,N_13059,N_15844);
nor U23477 (N_23477,N_15363,N_14853);
nand U23478 (N_23478,N_13996,N_18184);
or U23479 (N_23479,N_12766,N_17616);
nor U23480 (N_23480,N_13712,N_16725);
or U23481 (N_23481,N_15822,N_16751);
nand U23482 (N_23482,N_13322,N_16738);
nand U23483 (N_23483,N_16334,N_12737);
and U23484 (N_23484,N_18397,N_17177);
and U23485 (N_23485,N_14397,N_12727);
nor U23486 (N_23486,N_15342,N_13523);
xnor U23487 (N_23487,N_17650,N_16916);
nand U23488 (N_23488,N_14611,N_15726);
or U23489 (N_23489,N_13896,N_14152);
or U23490 (N_23490,N_15775,N_12819);
nand U23491 (N_23491,N_13146,N_16823);
nor U23492 (N_23492,N_17009,N_18218);
and U23493 (N_23493,N_17679,N_17896);
nor U23494 (N_23494,N_16898,N_14178);
nand U23495 (N_23495,N_14777,N_13500);
and U23496 (N_23496,N_17742,N_13449);
nand U23497 (N_23497,N_13974,N_12615);
and U23498 (N_23498,N_14579,N_18042);
and U23499 (N_23499,N_15729,N_16320);
nand U23500 (N_23500,N_17216,N_16958);
or U23501 (N_23501,N_13826,N_12611);
nor U23502 (N_23502,N_18340,N_13187);
or U23503 (N_23503,N_16043,N_16698);
and U23504 (N_23504,N_14234,N_14654);
nor U23505 (N_23505,N_13215,N_15240);
or U23506 (N_23506,N_17202,N_16787);
nand U23507 (N_23507,N_16967,N_15867);
or U23508 (N_23508,N_14553,N_13223);
or U23509 (N_23509,N_15812,N_13977);
nor U23510 (N_23510,N_15842,N_16023);
nor U23511 (N_23511,N_13954,N_17924);
nand U23512 (N_23512,N_16226,N_17799);
nor U23513 (N_23513,N_15284,N_18675);
nand U23514 (N_23514,N_14753,N_13344);
nand U23515 (N_23515,N_16332,N_17017);
and U23516 (N_23516,N_15474,N_14452);
and U23517 (N_23517,N_14450,N_16334);
or U23518 (N_23518,N_14016,N_16385);
and U23519 (N_23519,N_17757,N_13905);
nand U23520 (N_23520,N_16501,N_13831);
nand U23521 (N_23521,N_15612,N_17972);
and U23522 (N_23522,N_18153,N_17201);
nand U23523 (N_23523,N_14035,N_15183);
nand U23524 (N_23524,N_14959,N_13601);
or U23525 (N_23525,N_12815,N_12859);
nand U23526 (N_23526,N_17067,N_16807);
nor U23527 (N_23527,N_14787,N_16318);
nand U23528 (N_23528,N_15876,N_13493);
and U23529 (N_23529,N_12724,N_17389);
or U23530 (N_23530,N_14669,N_12964);
nor U23531 (N_23531,N_17517,N_14539);
nand U23532 (N_23532,N_17463,N_16992);
or U23533 (N_23533,N_16315,N_16198);
nor U23534 (N_23534,N_13955,N_12506);
and U23535 (N_23535,N_16412,N_15027);
nor U23536 (N_23536,N_13840,N_18088);
or U23537 (N_23537,N_17848,N_17997);
nand U23538 (N_23538,N_13068,N_17030);
and U23539 (N_23539,N_14384,N_13734);
nor U23540 (N_23540,N_14193,N_14610);
or U23541 (N_23541,N_18125,N_13058);
nor U23542 (N_23542,N_18228,N_13224);
nor U23543 (N_23543,N_15273,N_15597);
or U23544 (N_23544,N_13810,N_18472);
and U23545 (N_23545,N_14817,N_16787);
nand U23546 (N_23546,N_17844,N_15650);
nand U23547 (N_23547,N_14256,N_17084);
nand U23548 (N_23548,N_18534,N_14642);
nand U23549 (N_23549,N_14276,N_13969);
and U23550 (N_23550,N_16103,N_17218);
nor U23551 (N_23551,N_15106,N_16350);
nor U23552 (N_23552,N_14492,N_16903);
or U23553 (N_23553,N_18221,N_15364);
nor U23554 (N_23554,N_14591,N_13039);
nor U23555 (N_23555,N_14413,N_18282);
nand U23556 (N_23556,N_17593,N_17008);
or U23557 (N_23557,N_13420,N_13581);
nand U23558 (N_23558,N_18235,N_18672);
nor U23559 (N_23559,N_15925,N_12638);
and U23560 (N_23560,N_15295,N_16852);
nor U23561 (N_23561,N_17662,N_16124);
or U23562 (N_23562,N_16653,N_18728);
xnor U23563 (N_23563,N_18652,N_16369);
or U23564 (N_23564,N_12874,N_16945);
nor U23565 (N_23565,N_12814,N_13790);
nand U23566 (N_23566,N_12819,N_13982);
or U23567 (N_23567,N_14195,N_17074);
nor U23568 (N_23568,N_18348,N_16404);
or U23569 (N_23569,N_15292,N_12876);
nand U23570 (N_23570,N_15119,N_17251);
and U23571 (N_23571,N_16815,N_13638);
and U23572 (N_23572,N_16531,N_15675);
or U23573 (N_23573,N_14863,N_17632);
nor U23574 (N_23574,N_14974,N_13519);
or U23575 (N_23575,N_14235,N_17154);
or U23576 (N_23576,N_16820,N_18557);
nor U23577 (N_23577,N_17745,N_15154);
and U23578 (N_23578,N_13819,N_13630);
nor U23579 (N_23579,N_12534,N_18676);
nor U23580 (N_23580,N_17318,N_17495);
nor U23581 (N_23581,N_16181,N_15123);
nor U23582 (N_23582,N_18593,N_16223);
nand U23583 (N_23583,N_18364,N_13459);
and U23584 (N_23584,N_18606,N_15536);
nand U23585 (N_23585,N_18275,N_17637);
and U23586 (N_23586,N_17280,N_14023);
xor U23587 (N_23587,N_18415,N_15051);
xor U23588 (N_23588,N_17418,N_14486);
nand U23589 (N_23589,N_12825,N_15759);
and U23590 (N_23590,N_13026,N_17042);
and U23591 (N_23591,N_13552,N_16014);
nand U23592 (N_23592,N_12777,N_18216);
or U23593 (N_23593,N_15971,N_14873);
nand U23594 (N_23594,N_12923,N_13389);
and U23595 (N_23595,N_13805,N_15573);
and U23596 (N_23596,N_15793,N_16214);
nor U23597 (N_23597,N_15660,N_16821);
nor U23598 (N_23598,N_13831,N_16669);
nor U23599 (N_23599,N_18589,N_13147);
and U23600 (N_23600,N_18387,N_17086);
and U23601 (N_23601,N_13168,N_14174);
and U23602 (N_23602,N_17338,N_13915);
nor U23603 (N_23603,N_16119,N_16341);
and U23604 (N_23604,N_16572,N_14997);
nand U23605 (N_23605,N_14053,N_18175);
nor U23606 (N_23606,N_13343,N_16541);
and U23607 (N_23607,N_13074,N_17686);
or U23608 (N_23608,N_18438,N_16116);
nor U23609 (N_23609,N_16592,N_17886);
and U23610 (N_23610,N_13254,N_16938);
or U23611 (N_23611,N_13359,N_16276);
and U23612 (N_23612,N_16201,N_13843);
nor U23613 (N_23613,N_16866,N_14246);
xor U23614 (N_23614,N_13690,N_13183);
nor U23615 (N_23615,N_13277,N_17568);
and U23616 (N_23616,N_15417,N_17738);
nor U23617 (N_23617,N_18595,N_16141);
nand U23618 (N_23618,N_13730,N_18706);
or U23619 (N_23619,N_16773,N_14437);
nor U23620 (N_23620,N_13073,N_12968);
nand U23621 (N_23621,N_15411,N_18082);
nor U23622 (N_23622,N_17544,N_15830);
nand U23623 (N_23623,N_15767,N_18589);
and U23624 (N_23624,N_12714,N_15706);
or U23625 (N_23625,N_14623,N_16422);
and U23626 (N_23626,N_13768,N_18619);
nor U23627 (N_23627,N_14477,N_13644);
nand U23628 (N_23628,N_18405,N_17334);
nor U23629 (N_23629,N_13723,N_18261);
or U23630 (N_23630,N_14375,N_18117);
nand U23631 (N_23631,N_16046,N_15648);
nand U23632 (N_23632,N_14970,N_16355);
or U23633 (N_23633,N_17616,N_16065);
nand U23634 (N_23634,N_14321,N_16493);
nor U23635 (N_23635,N_18469,N_13066);
or U23636 (N_23636,N_15943,N_14893);
nor U23637 (N_23637,N_13620,N_16770);
and U23638 (N_23638,N_16209,N_13017);
and U23639 (N_23639,N_13906,N_12671);
and U23640 (N_23640,N_15609,N_14079);
nand U23641 (N_23641,N_14701,N_14736);
nand U23642 (N_23642,N_14961,N_12584);
and U23643 (N_23643,N_14268,N_17416);
and U23644 (N_23644,N_17164,N_14657);
nor U23645 (N_23645,N_16734,N_15951);
nor U23646 (N_23646,N_15156,N_12949);
nand U23647 (N_23647,N_16638,N_14926);
or U23648 (N_23648,N_13843,N_15609);
nor U23649 (N_23649,N_14602,N_15939);
nor U23650 (N_23650,N_15863,N_18615);
or U23651 (N_23651,N_16162,N_18249);
and U23652 (N_23652,N_14007,N_13458);
or U23653 (N_23653,N_13020,N_16604);
nand U23654 (N_23654,N_14042,N_12961);
nand U23655 (N_23655,N_18049,N_12508);
or U23656 (N_23656,N_16101,N_18510);
xnor U23657 (N_23657,N_16821,N_14057);
nor U23658 (N_23658,N_16022,N_17462);
and U23659 (N_23659,N_16934,N_17786);
or U23660 (N_23660,N_14828,N_18511);
and U23661 (N_23661,N_14533,N_18488);
xnor U23662 (N_23662,N_14045,N_12519);
or U23663 (N_23663,N_18629,N_14747);
and U23664 (N_23664,N_15457,N_14001);
nand U23665 (N_23665,N_18303,N_15315);
or U23666 (N_23666,N_17453,N_14149);
or U23667 (N_23667,N_15791,N_17947);
nor U23668 (N_23668,N_14611,N_14875);
or U23669 (N_23669,N_13522,N_16529);
or U23670 (N_23670,N_13469,N_12554);
and U23671 (N_23671,N_12914,N_17235);
nand U23672 (N_23672,N_17392,N_17815);
or U23673 (N_23673,N_17642,N_15968);
or U23674 (N_23674,N_17504,N_14887);
or U23675 (N_23675,N_14520,N_12508);
nor U23676 (N_23676,N_16493,N_14446);
nor U23677 (N_23677,N_14775,N_17020);
and U23678 (N_23678,N_13449,N_15093);
nand U23679 (N_23679,N_13944,N_16576);
nor U23680 (N_23680,N_13979,N_13122);
nor U23681 (N_23681,N_15920,N_15430);
nand U23682 (N_23682,N_13814,N_18638);
nor U23683 (N_23683,N_15234,N_13886);
and U23684 (N_23684,N_13931,N_15317);
and U23685 (N_23685,N_17572,N_17249);
nand U23686 (N_23686,N_18564,N_15199);
and U23687 (N_23687,N_18224,N_12682);
nand U23688 (N_23688,N_12593,N_15524);
nand U23689 (N_23689,N_17809,N_17642);
nand U23690 (N_23690,N_13731,N_13695);
or U23691 (N_23691,N_12907,N_16159);
nand U23692 (N_23692,N_17714,N_12843);
and U23693 (N_23693,N_18386,N_17211);
or U23694 (N_23694,N_12737,N_14767);
nand U23695 (N_23695,N_16840,N_14630);
and U23696 (N_23696,N_12957,N_14789);
nor U23697 (N_23697,N_13620,N_16358);
xor U23698 (N_23698,N_13451,N_15764);
nor U23699 (N_23699,N_15233,N_13583);
nand U23700 (N_23700,N_16086,N_17470);
nor U23701 (N_23701,N_13527,N_17721);
nand U23702 (N_23702,N_15560,N_16354);
or U23703 (N_23703,N_16215,N_15223);
nand U23704 (N_23704,N_12961,N_18633);
nand U23705 (N_23705,N_12922,N_15332);
or U23706 (N_23706,N_13209,N_13403);
nor U23707 (N_23707,N_18265,N_18250);
and U23708 (N_23708,N_15226,N_14481);
nand U23709 (N_23709,N_15285,N_14471);
nor U23710 (N_23710,N_18072,N_16250);
nor U23711 (N_23711,N_16981,N_12817);
nor U23712 (N_23712,N_12756,N_16617);
and U23713 (N_23713,N_18249,N_14800);
and U23714 (N_23714,N_18039,N_14232);
nand U23715 (N_23715,N_12618,N_13029);
or U23716 (N_23716,N_16412,N_17381);
nor U23717 (N_23717,N_14595,N_15049);
nand U23718 (N_23718,N_18133,N_17299);
or U23719 (N_23719,N_17360,N_18365);
nand U23720 (N_23720,N_17377,N_12966);
and U23721 (N_23721,N_13790,N_13463);
or U23722 (N_23722,N_12738,N_17614);
nand U23723 (N_23723,N_18077,N_13030);
nor U23724 (N_23724,N_13327,N_13148);
nand U23725 (N_23725,N_13961,N_17446);
and U23726 (N_23726,N_15461,N_14979);
and U23727 (N_23727,N_12901,N_13205);
or U23728 (N_23728,N_17470,N_16303);
or U23729 (N_23729,N_14802,N_12817);
nand U23730 (N_23730,N_17298,N_17383);
nor U23731 (N_23731,N_16384,N_14545);
nand U23732 (N_23732,N_16586,N_12729);
nor U23733 (N_23733,N_17835,N_13409);
nor U23734 (N_23734,N_16968,N_15641);
nand U23735 (N_23735,N_15779,N_16306);
nor U23736 (N_23736,N_16475,N_16054);
or U23737 (N_23737,N_15947,N_12560);
and U23738 (N_23738,N_14673,N_16338);
nor U23739 (N_23739,N_13920,N_16900);
and U23740 (N_23740,N_13152,N_16577);
and U23741 (N_23741,N_16943,N_17628);
nor U23742 (N_23742,N_14131,N_18567);
nand U23743 (N_23743,N_17525,N_17218);
or U23744 (N_23744,N_15860,N_13410);
or U23745 (N_23745,N_16824,N_13222);
nand U23746 (N_23746,N_15845,N_14788);
nor U23747 (N_23747,N_17470,N_17570);
nor U23748 (N_23748,N_15836,N_17612);
nor U23749 (N_23749,N_18718,N_14912);
or U23750 (N_23750,N_18041,N_17215);
or U23751 (N_23751,N_15816,N_15765);
or U23752 (N_23752,N_14899,N_18240);
or U23753 (N_23753,N_16315,N_13134);
or U23754 (N_23754,N_14567,N_18309);
nor U23755 (N_23755,N_17613,N_13048);
and U23756 (N_23756,N_14333,N_15665);
or U23757 (N_23757,N_16580,N_13941);
and U23758 (N_23758,N_13304,N_14603);
nor U23759 (N_23759,N_18060,N_13365);
or U23760 (N_23760,N_18002,N_14800);
nor U23761 (N_23761,N_16895,N_16474);
or U23762 (N_23762,N_14631,N_15234);
or U23763 (N_23763,N_18004,N_16029);
or U23764 (N_23764,N_17070,N_14424);
and U23765 (N_23765,N_18499,N_13664);
and U23766 (N_23766,N_13521,N_14391);
nand U23767 (N_23767,N_13722,N_17183);
and U23768 (N_23768,N_17618,N_14121);
nor U23769 (N_23769,N_16243,N_13066);
nand U23770 (N_23770,N_14467,N_16018);
or U23771 (N_23771,N_14349,N_18085);
or U23772 (N_23772,N_18459,N_13515);
nor U23773 (N_23773,N_14946,N_15320);
nand U23774 (N_23774,N_13304,N_13271);
nor U23775 (N_23775,N_14938,N_18704);
nand U23776 (N_23776,N_15203,N_17611);
nor U23777 (N_23777,N_17272,N_16039);
and U23778 (N_23778,N_14854,N_16083);
nand U23779 (N_23779,N_17441,N_15424);
nor U23780 (N_23780,N_13100,N_16159);
or U23781 (N_23781,N_14118,N_14861);
or U23782 (N_23782,N_13566,N_16536);
nand U23783 (N_23783,N_18341,N_15063);
nand U23784 (N_23784,N_18531,N_18200);
nor U23785 (N_23785,N_17578,N_12757);
and U23786 (N_23786,N_17558,N_18366);
or U23787 (N_23787,N_15960,N_16341);
and U23788 (N_23788,N_15042,N_18138);
and U23789 (N_23789,N_18150,N_14444);
nand U23790 (N_23790,N_12687,N_14748);
nor U23791 (N_23791,N_14193,N_12563);
and U23792 (N_23792,N_12566,N_18641);
or U23793 (N_23793,N_17279,N_18625);
nand U23794 (N_23794,N_14116,N_15548);
or U23795 (N_23795,N_17078,N_16160);
nand U23796 (N_23796,N_15643,N_13791);
nand U23797 (N_23797,N_15967,N_13672);
or U23798 (N_23798,N_16255,N_17263);
or U23799 (N_23799,N_17920,N_16872);
or U23800 (N_23800,N_18507,N_12611);
and U23801 (N_23801,N_13735,N_15454);
nor U23802 (N_23802,N_16335,N_17577);
nand U23803 (N_23803,N_17074,N_13989);
nor U23804 (N_23804,N_14860,N_14643);
and U23805 (N_23805,N_18122,N_17413);
and U23806 (N_23806,N_16312,N_18389);
and U23807 (N_23807,N_15699,N_12816);
and U23808 (N_23808,N_12722,N_12508);
and U23809 (N_23809,N_15369,N_12517);
nor U23810 (N_23810,N_14459,N_13830);
and U23811 (N_23811,N_12717,N_17966);
nor U23812 (N_23812,N_15895,N_13996);
or U23813 (N_23813,N_15755,N_12814);
or U23814 (N_23814,N_14738,N_15157);
and U23815 (N_23815,N_14531,N_12674);
or U23816 (N_23816,N_15052,N_18293);
nor U23817 (N_23817,N_18372,N_15701);
nand U23818 (N_23818,N_16494,N_18106);
or U23819 (N_23819,N_12747,N_14570);
nor U23820 (N_23820,N_12983,N_16027);
xor U23821 (N_23821,N_18466,N_13654);
and U23822 (N_23822,N_17541,N_13794);
or U23823 (N_23823,N_14269,N_13415);
nor U23824 (N_23824,N_16940,N_16544);
nand U23825 (N_23825,N_17200,N_17026);
or U23826 (N_23826,N_17068,N_15096);
nor U23827 (N_23827,N_18383,N_14713);
or U23828 (N_23828,N_17901,N_15637);
nand U23829 (N_23829,N_16173,N_15412);
nor U23830 (N_23830,N_13692,N_15276);
nor U23831 (N_23831,N_16989,N_18609);
and U23832 (N_23832,N_17996,N_16193);
nand U23833 (N_23833,N_14933,N_14885);
and U23834 (N_23834,N_16194,N_18400);
nand U23835 (N_23835,N_18435,N_17161);
and U23836 (N_23836,N_15420,N_15746);
and U23837 (N_23837,N_13329,N_13931);
nand U23838 (N_23838,N_13749,N_18478);
and U23839 (N_23839,N_14090,N_16851);
and U23840 (N_23840,N_17596,N_17490);
nand U23841 (N_23841,N_16057,N_18629);
nand U23842 (N_23842,N_15952,N_15376);
xor U23843 (N_23843,N_17689,N_18026);
and U23844 (N_23844,N_15299,N_13447);
and U23845 (N_23845,N_18536,N_13974);
nand U23846 (N_23846,N_16453,N_16422);
nand U23847 (N_23847,N_14884,N_15257);
nor U23848 (N_23848,N_15610,N_17745);
or U23849 (N_23849,N_15850,N_18111);
and U23850 (N_23850,N_13865,N_17600);
and U23851 (N_23851,N_17506,N_17747);
nor U23852 (N_23852,N_14228,N_16825);
nor U23853 (N_23853,N_16269,N_13901);
or U23854 (N_23854,N_15684,N_13286);
nand U23855 (N_23855,N_12514,N_15902);
nor U23856 (N_23856,N_17074,N_13975);
nor U23857 (N_23857,N_17834,N_18013);
or U23858 (N_23858,N_17074,N_15387);
nand U23859 (N_23859,N_18425,N_17331);
nor U23860 (N_23860,N_13420,N_16474);
nand U23861 (N_23861,N_17175,N_17834);
or U23862 (N_23862,N_12678,N_15858);
nand U23863 (N_23863,N_13145,N_17572);
nand U23864 (N_23864,N_18465,N_17198);
nor U23865 (N_23865,N_17970,N_16262);
xor U23866 (N_23866,N_12733,N_13455);
or U23867 (N_23867,N_12833,N_14288);
or U23868 (N_23868,N_16927,N_15541);
or U23869 (N_23869,N_17627,N_14616);
nand U23870 (N_23870,N_16881,N_17858);
and U23871 (N_23871,N_13717,N_16402);
nand U23872 (N_23872,N_17735,N_17511);
and U23873 (N_23873,N_16769,N_13616);
or U23874 (N_23874,N_17399,N_14032);
and U23875 (N_23875,N_13154,N_13961);
and U23876 (N_23876,N_13762,N_13922);
nand U23877 (N_23877,N_13807,N_17956);
or U23878 (N_23878,N_16137,N_15258);
or U23879 (N_23879,N_14464,N_12869);
or U23880 (N_23880,N_14085,N_13436);
and U23881 (N_23881,N_18427,N_14316);
or U23882 (N_23882,N_16286,N_17327);
or U23883 (N_23883,N_13416,N_16920);
or U23884 (N_23884,N_17687,N_16628);
nor U23885 (N_23885,N_15009,N_13570);
and U23886 (N_23886,N_18641,N_16297);
and U23887 (N_23887,N_15376,N_17167);
nand U23888 (N_23888,N_16870,N_16011);
xnor U23889 (N_23889,N_14956,N_17127);
and U23890 (N_23890,N_16833,N_12821);
nand U23891 (N_23891,N_15000,N_12884);
and U23892 (N_23892,N_12946,N_13039);
or U23893 (N_23893,N_18641,N_17178);
and U23894 (N_23894,N_15908,N_14973);
nand U23895 (N_23895,N_18122,N_18488);
nand U23896 (N_23896,N_17119,N_18369);
and U23897 (N_23897,N_14772,N_18310);
nor U23898 (N_23898,N_16511,N_13480);
nor U23899 (N_23899,N_14818,N_16086);
or U23900 (N_23900,N_17464,N_13527);
nand U23901 (N_23901,N_14084,N_13998);
and U23902 (N_23902,N_18245,N_17644);
nor U23903 (N_23903,N_13790,N_18510);
nand U23904 (N_23904,N_17416,N_16988);
or U23905 (N_23905,N_17996,N_14350);
or U23906 (N_23906,N_18534,N_17151);
or U23907 (N_23907,N_14031,N_15637);
and U23908 (N_23908,N_14336,N_17290);
and U23909 (N_23909,N_13990,N_15694);
or U23910 (N_23910,N_13608,N_13995);
nor U23911 (N_23911,N_12731,N_13386);
or U23912 (N_23912,N_13809,N_16820);
and U23913 (N_23913,N_16653,N_16735);
nor U23914 (N_23914,N_14355,N_14186);
and U23915 (N_23915,N_17723,N_15005);
and U23916 (N_23916,N_13168,N_17439);
nor U23917 (N_23917,N_16341,N_13120);
nor U23918 (N_23918,N_12876,N_13395);
nor U23919 (N_23919,N_17503,N_12844);
or U23920 (N_23920,N_15509,N_16045);
nand U23921 (N_23921,N_18032,N_18303);
and U23922 (N_23922,N_13836,N_14051);
nand U23923 (N_23923,N_15416,N_13622);
or U23924 (N_23924,N_15975,N_12777);
nand U23925 (N_23925,N_16143,N_16030);
nor U23926 (N_23926,N_16210,N_17595);
nor U23927 (N_23927,N_18604,N_16211);
nor U23928 (N_23928,N_13220,N_15262);
or U23929 (N_23929,N_18596,N_15847);
nand U23930 (N_23930,N_16809,N_14799);
and U23931 (N_23931,N_16249,N_13078);
nor U23932 (N_23932,N_13083,N_13971);
or U23933 (N_23933,N_13417,N_16710);
nor U23934 (N_23934,N_12530,N_18533);
nand U23935 (N_23935,N_13607,N_14757);
nand U23936 (N_23936,N_16392,N_18257);
or U23937 (N_23937,N_15513,N_17794);
and U23938 (N_23938,N_17432,N_18399);
and U23939 (N_23939,N_18495,N_13084);
and U23940 (N_23940,N_13945,N_18621);
nand U23941 (N_23941,N_17262,N_17129);
and U23942 (N_23942,N_15424,N_12678);
and U23943 (N_23943,N_12549,N_17916);
nand U23944 (N_23944,N_18281,N_12697);
or U23945 (N_23945,N_14201,N_15323);
and U23946 (N_23946,N_16985,N_12876);
or U23947 (N_23947,N_16773,N_17736);
nand U23948 (N_23948,N_17172,N_17141);
nand U23949 (N_23949,N_18735,N_15714);
nor U23950 (N_23950,N_15703,N_14228);
nand U23951 (N_23951,N_13272,N_13088);
nand U23952 (N_23952,N_18722,N_13017);
and U23953 (N_23953,N_18393,N_15599);
or U23954 (N_23954,N_17245,N_14790);
and U23955 (N_23955,N_14875,N_14212);
or U23956 (N_23956,N_18683,N_17534);
and U23957 (N_23957,N_12925,N_15070);
and U23958 (N_23958,N_14847,N_13123);
nand U23959 (N_23959,N_18648,N_13879);
or U23960 (N_23960,N_14598,N_14059);
nand U23961 (N_23961,N_16773,N_15011);
or U23962 (N_23962,N_13334,N_13513);
nand U23963 (N_23963,N_13570,N_16325);
nand U23964 (N_23964,N_15737,N_13776);
nand U23965 (N_23965,N_12979,N_17771);
nand U23966 (N_23966,N_13179,N_13875);
nor U23967 (N_23967,N_16257,N_13739);
nand U23968 (N_23968,N_15744,N_13715);
nor U23969 (N_23969,N_12809,N_15321);
and U23970 (N_23970,N_14597,N_17183);
nand U23971 (N_23971,N_15022,N_16833);
nor U23972 (N_23972,N_14398,N_18529);
or U23973 (N_23973,N_14152,N_15796);
and U23974 (N_23974,N_17664,N_15544);
nand U23975 (N_23975,N_13981,N_15676);
nor U23976 (N_23976,N_15169,N_14635);
or U23977 (N_23977,N_13099,N_14341);
nand U23978 (N_23978,N_17768,N_15189);
or U23979 (N_23979,N_17597,N_15716);
nor U23980 (N_23980,N_15326,N_12607);
and U23981 (N_23981,N_17089,N_17695);
nand U23982 (N_23982,N_15000,N_13268);
nand U23983 (N_23983,N_12754,N_12769);
and U23984 (N_23984,N_16086,N_14189);
nand U23985 (N_23985,N_15541,N_13771);
nand U23986 (N_23986,N_16898,N_13688);
nor U23987 (N_23987,N_13963,N_16467);
nor U23988 (N_23988,N_16779,N_18470);
nor U23989 (N_23989,N_17548,N_14839);
or U23990 (N_23990,N_12807,N_16802);
nor U23991 (N_23991,N_13151,N_16461);
nand U23992 (N_23992,N_12733,N_16133);
xnor U23993 (N_23993,N_13071,N_14950);
nor U23994 (N_23994,N_16355,N_14835);
nor U23995 (N_23995,N_15090,N_17865);
nor U23996 (N_23996,N_14839,N_14628);
nor U23997 (N_23997,N_17880,N_14597);
nor U23998 (N_23998,N_13292,N_15005);
nor U23999 (N_23999,N_12631,N_16078);
or U24000 (N_24000,N_18433,N_16273);
or U24001 (N_24001,N_17541,N_14457);
or U24002 (N_24002,N_13360,N_14597);
nor U24003 (N_24003,N_15063,N_13370);
nor U24004 (N_24004,N_17041,N_13350);
or U24005 (N_24005,N_15789,N_17300);
and U24006 (N_24006,N_18338,N_15572);
and U24007 (N_24007,N_15540,N_13355);
or U24008 (N_24008,N_17198,N_14026);
nor U24009 (N_24009,N_13585,N_17657);
nor U24010 (N_24010,N_13071,N_14489);
nand U24011 (N_24011,N_17008,N_14904);
nand U24012 (N_24012,N_14580,N_17419);
nor U24013 (N_24013,N_13583,N_14039);
nand U24014 (N_24014,N_16901,N_15717);
or U24015 (N_24015,N_17024,N_16002);
and U24016 (N_24016,N_14609,N_16435);
or U24017 (N_24017,N_16498,N_15199);
and U24018 (N_24018,N_17803,N_13630);
nand U24019 (N_24019,N_15136,N_14537);
and U24020 (N_24020,N_15588,N_13565);
nand U24021 (N_24021,N_14771,N_14596);
nor U24022 (N_24022,N_17786,N_16199);
and U24023 (N_24023,N_16426,N_15131);
or U24024 (N_24024,N_14010,N_13522);
or U24025 (N_24025,N_15708,N_14337);
nand U24026 (N_24026,N_18548,N_17715);
or U24027 (N_24027,N_13825,N_17435);
and U24028 (N_24028,N_13501,N_13056);
nand U24029 (N_24029,N_15867,N_14469);
and U24030 (N_24030,N_15277,N_14887);
nor U24031 (N_24031,N_15999,N_16485);
and U24032 (N_24032,N_15390,N_13457);
and U24033 (N_24033,N_13689,N_17817);
nor U24034 (N_24034,N_13368,N_17592);
nor U24035 (N_24035,N_16728,N_18058);
or U24036 (N_24036,N_14694,N_14927);
nand U24037 (N_24037,N_17322,N_17366);
and U24038 (N_24038,N_17610,N_14352);
or U24039 (N_24039,N_12667,N_15092);
and U24040 (N_24040,N_16889,N_14528);
and U24041 (N_24041,N_15430,N_13080);
or U24042 (N_24042,N_12902,N_15972);
nor U24043 (N_24043,N_18470,N_17536);
or U24044 (N_24044,N_15124,N_12681);
and U24045 (N_24045,N_12776,N_18133);
and U24046 (N_24046,N_15942,N_16229);
or U24047 (N_24047,N_16077,N_15415);
and U24048 (N_24048,N_17264,N_14255);
and U24049 (N_24049,N_13037,N_12510);
or U24050 (N_24050,N_18469,N_16088);
nor U24051 (N_24051,N_13650,N_13756);
nor U24052 (N_24052,N_16960,N_13798);
nor U24053 (N_24053,N_18153,N_18460);
and U24054 (N_24054,N_16013,N_14860);
or U24055 (N_24055,N_13159,N_16126);
nor U24056 (N_24056,N_17237,N_14786);
nor U24057 (N_24057,N_13522,N_17965);
nor U24058 (N_24058,N_13493,N_16130);
nor U24059 (N_24059,N_15063,N_13590);
nand U24060 (N_24060,N_15770,N_16741);
and U24061 (N_24061,N_13985,N_16613);
nor U24062 (N_24062,N_16989,N_13608);
and U24063 (N_24063,N_16618,N_17746);
and U24064 (N_24064,N_18308,N_15785);
nor U24065 (N_24065,N_13343,N_16712);
or U24066 (N_24066,N_13023,N_15417);
nor U24067 (N_24067,N_17446,N_17154);
nand U24068 (N_24068,N_15017,N_18219);
and U24069 (N_24069,N_13953,N_16980);
nand U24070 (N_24070,N_15142,N_14761);
and U24071 (N_24071,N_16759,N_13889);
nor U24072 (N_24072,N_15601,N_16884);
nor U24073 (N_24073,N_15316,N_12605);
nor U24074 (N_24074,N_16924,N_16719);
and U24075 (N_24075,N_18171,N_17896);
or U24076 (N_24076,N_18049,N_13554);
and U24077 (N_24077,N_16096,N_18092);
nand U24078 (N_24078,N_17640,N_14436);
nor U24079 (N_24079,N_13982,N_14720);
and U24080 (N_24080,N_13670,N_13563);
or U24081 (N_24081,N_14212,N_16874);
nor U24082 (N_24082,N_15623,N_15465);
nor U24083 (N_24083,N_13537,N_15648);
or U24084 (N_24084,N_13892,N_16077);
and U24085 (N_24085,N_13264,N_13434);
nand U24086 (N_24086,N_16395,N_16753);
or U24087 (N_24087,N_15061,N_16788);
nor U24088 (N_24088,N_14518,N_17223);
or U24089 (N_24089,N_12541,N_13517);
nor U24090 (N_24090,N_12808,N_17128);
and U24091 (N_24091,N_14075,N_14327);
or U24092 (N_24092,N_15461,N_16546);
or U24093 (N_24093,N_15389,N_15681);
or U24094 (N_24094,N_14482,N_16241);
or U24095 (N_24095,N_17229,N_14864);
and U24096 (N_24096,N_14770,N_12590);
or U24097 (N_24097,N_14314,N_14564);
or U24098 (N_24098,N_16839,N_12800);
and U24099 (N_24099,N_15207,N_13876);
nand U24100 (N_24100,N_15262,N_13786);
nor U24101 (N_24101,N_17731,N_15919);
or U24102 (N_24102,N_14536,N_12863);
and U24103 (N_24103,N_13333,N_15838);
and U24104 (N_24104,N_18605,N_15546);
nor U24105 (N_24105,N_16521,N_15485);
and U24106 (N_24106,N_18199,N_17202);
nor U24107 (N_24107,N_12794,N_15413);
and U24108 (N_24108,N_15205,N_13351);
and U24109 (N_24109,N_18248,N_12994);
nor U24110 (N_24110,N_14342,N_17088);
or U24111 (N_24111,N_16957,N_15920);
nand U24112 (N_24112,N_17429,N_16201);
or U24113 (N_24113,N_17320,N_16276);
or U24114 (N_24114,N_14026,N_15746);
and U24115 (N_24115,N_17472,N_17514);
and U24116 (N_24116,N_17559,N_18136);
and U24117 (N_24117,N_15617,N_13900);
xor U24118 (N_24118,N_18310,N_14691);
xor U24119 (N_24119,N_12625,N_12851);
and U24120 (N_24120,N_16640,N_18426);
and U24121 (N_24121,N_18599,N_15448);
nand U24122 (N_24122,N_16978,N_14234);
or U24123 (N_24123,N_15570,N_16654);
nand U24124 (N_24124,N_15873,N_16436);
or U24125 (N_24125,N_17695,N_15104);
and U24126 (N_24126,N_17531,N_13601);
nor U24127 (N_24127,N_16829,N_13445);
nor U24128 (N_24128,N_13886,N_15197);
xor U24129 (N_24129,N_14033,N_18179);
xor U24130 (N_24130,N_15083,N_13232);
and U24131 (N_24131,N_12766,N_16940);
or U24132 (N_24132,N_16514,N_18435);
and U24133 (N_24133,N_17436,N_15891);
nand U24134 (N_24134,N_14757,N_16459);
nor U24135 (N_24135,N_17083,N_15690);
and U24136 (N_24136,N_15510,N_17687);
or U24137 (N_24137,N_15310,N_18352);
nand U24138 (N_24138,N_17187,N_17826);
nand U24139 (N_24139,N_16832,N_17283);
nand U24140 (N_24140,N_15942,N_14542);
nor U24141 (N_24141,N_14496,N_16126);
and U24142 (N_24142,N_18394,N_12723);
and U24143 (N_24143,N_17908,N_18420);
or U24144 (N_24144,N_18166,N_14817);
nand U24145 (N_24145,N_16058,N_16546);
nand U24146 (N_24146,N_17879,N_17405);
or U24147 (N_24147,N_14265,N_14748);
nand U24148 (N_24148,N_12982,N_13338);
nand U24149 (N_24149,N_16816,N_14175);
and U24150 (N_24150,N_17973,N_13576);
or U24151 (N_24151,N_15981,N_14416);
and U24152 (N_24152,N_15746,N_12782);
or U24153 (N_24153,N_17328,N_17223);
nand U24154 (N_24154,N_13850,N_14989);
or U24155 (N_24155,N_16862,N_16394);
nand U24156 (N_24156,N_13096,N_13750);
nand U24157 (N_24157,N_15533,N_13869);
or U24158 (N_24158,N_14125,N_12732);
and U24159 (N_24159,N_15068,N_15188);
or U24160 (N_24160,N_17887,N_14721);
and U24161 (N_24161,N_16948,N_16158);
or U24162 (N_24162,N_16494,N_13918);
or U24163 (N_24163,N_14982,N_17037);
nand U24164 (N_24164,N_12706,N_12754);
or U24165 (N_24165,N_18273,N_17366);
and U24166 (N_24166,N_15074,N_17382);
and U24167 (N_24167,N_13313,N_15286);
nand U24168 (N_24168,N_14880,N_14523);
or U24169 (N_24169,N_17871,N_16791);
nor U24170 (N_24170,N_17376,N_14070);
or U24171 (N_24171,N_13384,N_13777);
nor U24172 (N_24172,N_14063,N_12713);
xnor U24173 (N_24173,N_15816,N_17097);
or U24174 (N_24174,N_16925,N_13400);
and U24175 (N_24175,N_16405,N_17280);
and U24176 (N_24176,N_13035,N_12842);
and U24177 (N_24177,N_17694,N_17036);
and U24178 (N_24178,N_13997,N_15347);
nand U24179 (N_24179,N_13787,N_14230);
and U24180 (N_24180,N_16275,N_13155);
or U24181 (N_24181,N_14184,N_16938);
nor U24182 (N_24182,N_15337,N_18381);
and U24183 (N_24183,N_14573,N_14908);
nand U24184 (N_24184,N_12995,N_13575);
nand U24185 (N_24185,N_18577,N_15940);
nand U24186 (N_24186,N_12898,N_18389);
nand U24187 (N_24187,N_15393,N_14806);
or U24188 (N_24188,N_14106,N_18393);
nand U24189 (N_24189,N_15195,N_12579);
and U24190 (N_24190,N_12755,N_17467);
nor U24191 (N_24191,N_13534,N_16389);
or U24192 (N_24192,N_12915,N_13305);
or U24193 (N_24193,N_16166,N_15803);
and U24194 (N_24194,N_16518,N_16418);
or U24195 (N_24195,N_16979,N_14896);
and U24196 (N_24196,N_14919,N_14594);
nand U24197 (N_24197,N_12542,N_14453);
nand U24198 (N_24198,N_18318,N_14905);
nor U24199 (N_24199,N_12695,N_12891);
or U24200 (N_24200,N_18536,N_17258);
nor U24201 (N_24201,N_12546,N_14361);
nand U24202 (N_24202,N_17654,N_18168);
or U24203 (N_24203,N_14251,N_13626);
or U24204 (N_24204,N_13246,N_16802);
and U24205 (N_24205,N_15348,N_17505);
or U24206 (N_24206,N_14852,N_15310);
nand U24207 (N_24207,N_15517,N_14115);
nor U24208 (N_24208,N_17958,N_15048);
or U24209 (N_24209,N_16071,N_15732);
or U24210 (N_24210,N_15850,N_15025);
nor U24211 (N_24211,N_14640,N_18602);
or U24212 (N_24212,N_18035,N_17877);
nand U24213 (N_24213,N_14145,N_15164);
and U24214 (N_24214,N_16866,N_15416);
nor U24215 (N_24215,N_14469,N_16980);
nor U24216 (N_24216,N_16753,N_17838);
and U24217 (N_24217,N_17955,N_14722);
or U24218 (N_24218,N_13250,N_15799);
and U24219 (N_24219,N_18211,N_17060);
nor U24220 (N_24220,N_17195,N_14603);
nor U24221 (N_24221,N_15312,N_14525);
nor U24222 (N_24222,N_12966,N_15145);
nor U24223 (N_24223,N_16102,N_13517);
nor U24224 (N_24224,N_17093,N_13194);
or U24225 (N_24225,N_18555,N_17169);
and U24226 (N_24226,N_16656,N_15704);
and U24227 (N_24227,N_13470,N_14447);
nor U24228 (N_24228,N_13142,N_14395);
or U24229 (N_24229,N_17994,N_13192);
nor U24230 (N_24230,N_13483,N_18472);
nand U24231 (N_24231,N_17389,N_13366);
and U24232 (N_24232,N_16017,N_15795);
and U24233 (N_24233,N_14471,N_15767);
nor U24234 (N_24234,N_17817,N_13418);
nor U24235 (N_24235,N_13976,N_14452);
or U24236 (N_24236,N_16313,N_16767);
and U24237 (N_24237,N_18006,N_13533);
and U24238 (N_24238,N_13166,N_14896);
and U24239 (N_24239,N_18321,N_13467);
and U24240 (N_24240,N_14813,N_18324);
and U24241 (N_24241,N_17721,N_13549);
or U24242 (N_24242,N_16471,N_17077);
and U24243 (N_24243,N_15351,N_13478);
nand U24244 (N_24244,N_16424,N_17042);
or U24245 (N_24245,N_16813,N_18638);
or U24246 (N_24246,N_15335,N_15122);
nand U24247 (N_24247,N_15964,N_12874);
or U24248 (N_24248,N_15317,N_13307);
and U24249 (N_24249,N_16852,N_14374);
nor U24250 (N_24250,N_15522,N_14950);
and U24251 (N_24251,N_17719,N_17259);
nand U24252 (N_24252,N_16027,N_16494);
or U24253 (N_24253,N_14862,N_13306);
nor U24254 (N_24254,N_13715,N_16671);
or U24255 (N_24255,N_18180,N_14608);
nand U24256 (N_24256,N_12577,N_15755);
and U24257 (N_24257,N_13097,N_15437);
nor U24258 (N_24258,N_13159,N_16732);
nor U24259 (N_24259,N_15212,N_16973);
and U24260 (N_24260,N_16309,N_15380);
or U24261 (N_24261,N_17950,N_13857);
nor U24262 (N_24262,N_12605,N_15666);
and U24263 (N_24263,N_12702,N_16209);
and U24264 (N_24264,N_15121,N_17701);
nor U24265 (N_24265,N_12820,N_15579);
nand U24266 (N_24266,N_16218,N_14205);
and U24267 (N_24267,N_13036,N_14995);
and U24268 (N_24268,N_12624,N_17844);
and U24269 (N_24269,N_13829,N_16559);
nand U24270 (N_24270,N_14198,N_13569);
and U24271 (N_24271,N_17089,N_14509);
and U24272 (N_24272,N_13031,N_12701);
xnor U24273 (N_24273,N_13445,N_14006);
and U24274 (N_24274,N_13551,N_12813);
or U24275 (N_24275,N_14938,N_12849);
nor U24276 (N_24276,N_15567,N_14200);
and U24277 (N_24277,N_14176,N_14363);
and U24278 (N_24278,N_12662,N_14308);
and U24279 (N_24279,N_14078,N_14686);
and U24280 (N_24280,N_14615,N_16797);
nand U24281 (N_24281,N_16770,N_16976);
or U24282 (N_24282,N_13249,N_13097);
nor U24283 (N_24283,N_18209,N_17371);
and U24284 (N_24284,N_18309,N_18195);
nor U24285 (N_24285,N_14089,N_15526);
nor U24286 (N_24286,N_14498,N_12877);
or U24287 (N_24287,N_14648,N_15782);
or U24288 (N_24288,N_13291,N_15966);
nor U24289 (N_24289,N_18575,N_18365);
nand U24290 (N_24290,N_13068,N_14418);
or U24291 (N_24291,N_13525,N_14904);
xor U24292 (N_24292,N_15424,N_17159);
nor U24293 (N_24293,N_16734,N_13678);
or U24294 (N_24294,N_18000,N_16866);
nor U24295 (N_24295,N_12586,N_14361);
nand U24296 (N_24296,N_16546,N_16321);
xnor U24297 (N_24297,N_16294,N_14859);
nand U24298 (N_24298,N_14736,N_12907);
or U24299 (N_24299,N_18085,N_14689);
nand U24300 (N_24300,N_18039,N_16535);
nor U24301 (N_24301,N_16231,N_12920);
or U24302 (N_24302,N_12793,N_18568);
and U24303 (N_24303,N_13865,N_18378);
nor U24304 (N_24304,N_16634,N_12943);
or U24305 (N_24305,N_16200,N_12886);
nand U24306 (N_24306,N_17447,N_14417);
nor U24307 (N_24307,N_17806,N_15291);
and U24308 (N_24308,N_12899,N_16708);
nor U24309 (N_24309,N_17476,N_16298);
and U24310 (N_24310,N_15821,N_17242);
or U24311 (N_24311,N_14010,N_14734);
nand U24312 (N_24312,N_15597,N_17348);
or U24313 (N_24313,N_15650,N_16588);
nor U24314 (N_24314,N_15550,N_14861);
nor U24315 (N_24315,N_18091,N_15105);
nor U24316 (N_24316,N_16801,N_18053);
and U24317 (N_24317,N_14050,N_13486);
nand U24318 (N_24318,N_13531,N_18660);
and U24319 (N_24319,N_16719,N_17551);
nand U24320 (N_24320,N_13940,N_17779);
nand U24321 (N_24321,N_18615,N_17328);
nor U24322 (N_24322,N_17438,N_13657);
or U24323 (N_24323,N_18032,N_13531);
and U24324 (N_24324,N_12676,N_14257);
and U24325 (N_24325,N_17320,N_14887);
nand U24326 (N_24326,N_16644,N_13377);
or U24327 (N_24327,N_17950,N_15798);
nand U24328 (N_24328,N_14824,N_14925);
or U24329 (N_24329,N_14120,N_13331);
nand U24330 (N_24330,N_16015,N_16055);
or U24331 (N_24331,N_17352,N_16663);
and U24332 (N_24332,N_18603,N_17730);
or U24333 (N_24333,N_13325,N_14280);
nor U24334 (N_24334,N_18217,N_17282);
or U24335 (N_24335,N_13751,N_16928);
and U24336 (N_24336,N_14510,N_14171);
and U24337 (N_24337,N_18167,N_14227);
or U24338 (N_24338,N_14662,N_16880);
and U24339 (N_24339,N_13513,N_18632);
nor U24340 (N_24340,N_13173,N_13891);
or U24341 (N_24341,N_12514,N_15652);
and U24342 (N_24342,N_18737,N_17074);
xnor U24343 (N_24343,N_13233,N_16371);
nand U24344 (N_24344,N_17160,N_16289);
nor U24345 (N_24345,N_12547,N_15780);
and U24346 (N_24346,N_16082,N_13341);
and U24347 (N_24347,N_16052,N_15718);
nor U24348 (N_24348,N_18098,N_12798);
or U24349 (N_24349,N_13487,N_16725);
or U24350 (N_24350,N_14080,N_13649);
or U24351 (N_24351,N_14662,N_14314);
or U24352 (N_24352,N_16301,N_16467);
or U24353 (N_24353,N_17815,N_12861);
nor U24354 (N_24354,N_17631,N_18205);
or U24355 (N_24355,N_14824,N_18716);
and U24356 (N_24356,N_13503,N_18071);
and U24357 (N_24357,N_17026,N_17170);
nand U24358 (N_24358,N_12680,N_13096);
and U24359 (N_24359,N_15464,N_15606);
nand U24360 (N_24360,N_16463,N_13187);
and U24361 (N_24361,N_12647,N_13850);
or U24362 (N_24362,N_12983,N_14589);
and U24363 (N_24363,N_13306,N_17520);
or U24364 (N_24364,N_18624,N_13289);
and U24365 (N_24365,N_13634,N_14275);
nand U24366 (N_24366,N_15135,N_16777);
nor U24367 (N_24367,N_15160,N_15050);
nor U24368 (N_24368,N_18340,N_14393);
nor U24369 (N_24369,N_12736,N_16858);
or U24370 (N_24370,N_16838,N_12660);
nor U24371 (N_24371,N_17079,N_17332);
or U24372 (N_24372,N_14015,N_14525);
or U24373 (N_24373,N_13484,N_16862);
and U24374 (N_24374,N_13567,N_14300);
and U24375 (N_24375,N_12837,N_16341);
nor U24376 (N_24376,N_14942,N_15140);
and U24377 (N_24377,N_17290,N_13004);
and U24378 (N_24378,N_18217,N_16607);
nor U24379 (N_24379,N_18179,N_14818);
or U24380 (N_24380,N_16459,N_12910);
nand U24381 (N_24381,N_15202,N_16304);
or U24382 (N_24382,N_15361,N_15182);
and U24383 (N_24383,N_15509,N_17400);
xor U24384 (N_24384,N_13885,N_18218);
and U24385 (N_24385,N_16099,N_16444);
nor U24386 (N_24386,N_14213,N_16553);
nor U24387 (N_24387,N_16331,N_13297);
nand U24388 (N_24388,N_16766,N_14241);
or U24389 (N_24389,N_18244,N_15930);
nand U24390 (N_24390,N_17946,N_15924);
nand U24391 (N_24391,N_14597,N_16438);
nand U24392 (N_24392,N_18163,N_14015);
or U24393 (N_24393,N_13485,N_18047);
nand U24394 (N_24394,N_14664,N_17550);
nor U24395 (N_24395,N_16700,N_15715);
or U24396 (N_24396,N_12703,N_13712);
nor U24397 (N_24397,N_16591,N_13976);
nand U24398 (N_24398,N_18460,N_13177);
and U24399 (N_24399,N_15873,N_18121);
and U24400 (N_24400,N_13837,N_15264);
and U24401 (N_24401,N_13624,N_16516);
nand U24402 (N_24402,N_16700,N_15203);
nand U24403 (N_24403,N_17428,N_14489);
and U24404 (N_24404,N_12670,N_18225);
nor U24405 (N_24405,N_12704,N_16012);
and U24406 (N_24406,N_18149,N_12641);
nor U24407 (N_24407,N_15903,N_13516);
nor U24408 (N_24408,N_16933,N_14065);
nand U24409 (N_24409,N_13692,N_16842);
nor U24410 (N_24410,N_13209,N_17295);
nand U24411 (N_24411,N_16730,N_14205);
nor U24412 (N_24412,N_15133,N_14430);
nor U24413 (N_24413,N_18735,N_16203);
nand U24414 (N_24414,N_16880,N_18504);
nand U24415 (N_24415,N_18037,N_14785);
or U24416 (N_24416,N_15541,N_14714);
and U24417 (N_24417,N_18326,N_17769);
nand U24418 (N_24418,N_17543,N_13014);
or U24419 (N_24419,N_18114,N_14994);
nor U24420 (N_24420,N_15190,N_18028);
or U24421 (N_24421,N_14513,N_16552);
or U24422 (N_24422,N_16801,N_18317);
nor U24423 (N_24423,N_13618,N_17357);
nor U24424 (N_24424,N_13718,N_15086);
nand U24425 (N_24425,N_18174,N_13725);
nand U24426 (N_24426,N_17668,N_15559);
nor U24427 (N_24427,N_12923,N_13583);
or U24428 (N_24428,N_17134,N_15337);
nand U24429 (N_24429,N_18604,N_13137);
nor U24430 (N_24430,N_13030,N_13396);
and U24431 (N_24431,N_18558,N_13898);
and U24432 (N_24432,N_14065,N_14356);
nor U24433 (N_24433,N_16783,N_14665);
nor U24434 (N_24434,N_16900,N_16539);
or U24435 (N_24435,N_14301,N_15740);
or U24436 (N_24436,N_17303,N_18171);
or U24437 (N_24437,N_13092,N_16421);
and U24438 (N_24438,N_16468,N_17180);
nand U24439 (N_24439,N_14422,N_16787);
nand U24440 (N_24440,N_16978,N_13748);
nand U24441 (N_24441,N_12958,N_15500);
nand U24442 (N_24442,N_12718,N_12805);
and U24443 (N_24443,N_13144,N_16447);
or U24444 (N_24444,N_13479,N_18072);
nand U24445 (N_24445,N_15580,N_15433);
nand U24446 (N_24446,N_15665,N_13489);
and U24447 (N_24447,N_13347,N_17214);
or U24448 (N_24448,N_18018,N_15885);
and U24449 (N_24449,N_17828,N_16158);
nand U24450 (N_24450,N_17199,N_13960);
nor U24451 (N_24451,N_18322,N_17516);
or U24452 (N_24452,N_13730,N_13744);
or U24453 (N_24453,N_17876,N_16569);
and U24454 (N_24454,N_14695,N_18365);
nor U24455 (N_24455,N_18287,N_15681);
nand U24456 (N_24456,N_14321,N_18496);
or U24457 (N_24457,N_13759,N_14270);
or U24458 (N_24458,N_12998,N_16131);
nand U24459 (N_24459,N_18513,N_15248);
nand U24460 (N_24460,N_14170,N_16061);
or U24461 (N_24461,N_17311,N_15709);
nor U24462 (N_24462,N_18689,N_14275);
or U24463 (N_24463,N_15847,N_16294);
or U24464 (N_24464,N_17547,N_16085);
nor U24465 (N_24465,N_17591,N_14250);
or U24466 (N_24466,N_14244,N_14380);
nand U24467 (N_24467,N_14568,N_16283);
nand U24468 (N_24468,N_17359,N_12756);
nand U24469 (N_24469,N_17233,N_17676);
nor U24470 (N_24470,N_12860,N_14071);
nand U24471 (N_24471,N_15351,N_17455);
or U24472 (N_24472,N_14232,N_16457);
nand U24473 (N_24473,N_13321,N_15662);
nor U24474 (N_24474,N_14121,N_15010);
nor U24475 (N_24475,N_16274,N_17611);
nand U24476 (N_24476,N_18490,N_18154);
or U24477 (N_24477,N_14507,N_12575);
nor U24478 (N_24478,N_14750,N_16188);
and U24479 (N_24479,N_12781,N_18507);
and U24480 (N_24480,N_15443,N_13600);
nor U24481 (N_24481,N_17393,N_16181);
xor U24482 (N_24482,N_12834,N_15623);
nor U24483 (N_24483,N_14199,N_16268);
and U24484 (N_24484,N_15289,N_17262);
nand U24485 (N_24485,N_16821,N_12943);
nor U24486 (N_24486,N_16912,N_15486);
or U24487 (N_24487,N_13953,N_16890);
nand U24488 (N_24488,N_13223,N_15279);
or U24489 (N_24489,N_14865,N_17215);
nor U24490 (N_24490,N_13819,N_12653);
nand U24491 (N_24491,N_17262,N_17642);
nor U24492 (N_24492,N_16493,N_17300);
or U24493 (N_24493,N_14869,N_14902);
nand U24494 (N_24494,N_14589,N_12846);
nor U24495 (N_24495,N_18426,N_15884);
nand U24496 (N_24496,N_16759,N_15402);
and U24497 (N_24497,N_18628,N_16914);
and U24498 (N_24498,N_18087,N_13240);
and U24499 (N_24499,N_18274,N_13054);
nand U24500 (N_24500,N_14482,N_15537);
and U24501 (N_24501,N_15866,N_16810);
nand U24502 (N_24502,N_18714,N_15363);
and U24503 (N_24503,N_15957,N_15452);
or U24504 (N_24504,N_17561,N_13997);
or U24505 (N_24505,N_13565,N_17970);
and U24506 (N_24506,N_18697,N_16311);
and U24507 (N_24507,N_15215,N_16082);
and U24508 (N_24508,N_12893,N_13917);
nand U24509 (N_24509,N_12702,N_13756);
nand U24510 (N_24510,N_16997,N_12639);
or U24511 (N_24511,N_18085,N_16517);
nand U24512 (N_24512,N_15181,N_12771);
and U24513 (N_24513,N_15424,N_16022);
and U24514 (N_24514,N_18185,N_18336);
nand U24515 (N_24515,N_15616,N_17793);
nand U24516 (N_24516,N_17487,N_15017);
or U24517 (N_24517,N_15091,N_15298);
or U24518 (N_24518,N_13903,N_13382);
nand U24519 (N_24519,N_16602,N_18674);
or U24520 (N_24520,N_12689,N_12990);
or U24521 (N_24521,N_13269,N_13680);
nand U24522 (N_24522,N_12898,N_13100);
or U24523 (N_24523,N_17452,N_17100);
or U24524 (N_24524,N_12889,N_15839);
nand U24525 (N_24525,N_16527,N_15863);
or U24526 (N_24526,N_15698,N_15324);
nand U24527 (N_24527,N_14229,N_13006);
and U24528 (N_24528,N_13352,N_13094);
and U24529 (N_24529,N_15348,N_14738);
or U24530 (N_24530,N_18097,N_15369);
nor U24531 (N_24531,N_14559,N_17310);
or U24532 (N_24532,N_18654,N_14117);
nand U24533 (N_24533,N_13424,N_15242);
nor U24534 (N_24534,N_17112,N_14365);
nand U24535 (N_24535,N_13525,N_14731);
or U24536 (N_24536,N_16806,N_16247);
nand U24537 (N_24537,N_16022,N_17621);
and U24538 (N_24538,N_13239,N_18047);
and U24539 (N_24539,N_17234,N_17400);
and U24540 (N_24540,N_14803,N_17220);
nor U24541 (N_24541,N_15877,N_17256);
or U24542 (N_24542,N_17395,N_12545);
and U24543 (N_24543,N_17330,N_15072);
nor U24544 (N_24544,N_14494,N_13641);
or U24545 (N_24545,N_18158,N_17390);
or U24546 (N_24546,N_14087,N_12983);
nor U24547 (N_24547,N_17312,N_15831);
and U24548 (N_24548,N_13511,N_15311);
and U24549 (N_24549,N_18387,N_15738);
nor U24550 (N_24550,N_17202,N_18243);
nor U24551 (N_24551,N_12609,N_16294);
nor U24552 (N_24552,N_16060,N_16206);
nor U24553 (N_24553,N_17402,N_14716);
nand U24554 (N_24554,N_15791,N_18014);
nand U24555 (N_24555,N_18336,N_18309);
or U24556 (N_24556,N_14558,N_14362);
nand U24557 (N_24557,N_18488,N_14571);
nor U24558 (N_24558,N_16430,N_16182);
and U24559 (N_24559,N_14021,N_13080);
and U24560 (N_24560,N_16512,N_16842);
nor U24561 (N_24561,N_13678,N_14279);
nor U24562 (N_24562,N_17192,N_15807);
nor U24563 (N_24563,N_17736,N_12538);
or U24564 (N_24564,N_16176,N_13340);
or U24565 (N_24565,N_14275,N_12833);
and U24566 (N_24566,N_16711,N_13728);
nand U24567 (N_24567,N_12917,N_18047);
and U24568 (N_24568,N_15828,N_15107);
nor U24569 (N_24569,N_16012,N_14760);
nor U24570 (N_24570,N_17900,N_16925);
and U24571 (N_24571,N_13505,N_12709);
and U24572 (N_24572,N_17559,N_16867);
or U24573 (N_24573,N_15746,N_18607);
or U24574 (N_24574,N_14936,N_12804);
nand U24575 (N_24575,N_15834,N_12889);
nor U24576 (N_24576,N_14643,N_14025);
nand U24577 (N_24577,N_12901,N_15826);
or U24578 (N_24578,N_17594,N_17392);
or U24579 (N_24579,N_14214,N_18261);
and U24580 (N_24580,N_17311,N_17741);
and U24581 (N_24581,N_13125,N_12854);
nand U24582 (N_24582,N_15115,N_15014);
or U24583 (N_24583,N_16980,N_15678);
or U24584 (N_24584,N_14947,N_12789);
nor U24585 (N_24585,N_17991,N_15476);
nand U24586 (N_24586,N_17897,N_12898);
nor U24587 (N_24587,N_18705,N_17188);
or U24588 (N_24588,N_18705,N_17862);
and U24589 (N_24589,N_17259,N_12652);
and U24590 (N_24590,N_18644,N_16862);
or U24591 (N_24591,N_15105,N_16907);
and U24592 (N_24592,N_13943,N_15238);
or U24593 (N_24593,N_12862,N_18009);
or U24594 (N_24594,N_14212,N_17609);
nand U24595 (N_24595,N_13955,N_18604);
and U24596 (N_24596,N_12925,N_15367);
nor U24597 (N_24597,N_17134,N_18070);
and U24598 (N_24598,N_13195,N_17727);
nand U24599 (N_24599,N_15456,N_14383);
nand U24600 (N_24600,N_16116,N_18318);
nand U24601 (N_24601,N_14805,N_18412);
and U24602 (N_24602,N_14911,N_15737);
nand U24603 (N_24603,N_14707,N_14398);
and U24604 (N_24604,N_18446,N_13835);
nand U24605 (N_24605,N_17127,N_14866);
and U24606 (N_24606,N_15824,N_13346);
and U24607 (N_24607,N_12716,N_13447);
nor U24608 (N_24608,N_15332,N_16831);
or U24609 (N_24609,N_18552,N_12581);
or U24610 (N_24610,N_15956,N_15018);
or U24611 (N_24611,N_17352,N_17712);
nand U24612 (N_24612,N_13694,N_12772);
and U24613 (N_24613,N_15972,N_14285);
or U24614 (N_24614,N_18310,N_14333);
or U24615 (N_24615,N_16332,N_12724);
and U24616 (N_24616,N_15314,N_15354);
xor U24617 (N_24617,N_12843,N_14356);
nor U24618 (N_24618,N_16833,N_13778);
or U24619 (N_24619,N_12618,N_17752);
and U24620 (N_24620,N_16867,N_14281);
nand U24621 (N_24621,N_16485,N_15144);
and U24622 (N_24622,N_15004,N_17969);
and U24623 (N_24623,N_14220,N_12657);
nand U24624 (N_24624,N_14200,N_15860);
or U24625 (N_24625,N_16190,N_13741);
nor U24626 (N_24626,N_16998,N_17118);
or U24627 (N_24627,N_18327,N_15456);
and U24628 (N_24628,N_12878,N_15747);
and U24629 (N_24629,N_17960,N_16104);
nand U24630 (N_24630,N_14479,N_17260);
or U24631 (N_24631,N_12681,N_15839);
nor U24632 (N_24632,N_14120,N_16381);
nor U24633 (N_24633,N_14185,N_15264);
nor U24634 (N_24634,N_13702,N_16441);
nor U24635 (N_24635,N_13134,N_16840);
or U24636 (N_24636,N_12599,N_15992);
and U24637 (N_24637,N_15366,N_16052);
and U24638 (N_24638,N_12935,N_17797);
nand U24639 (N_24639,N_13468,N_16142);
nand U24640 (N_24640,N_18672,N_18492);
nand U24641 (N_24641,N_13441,N_13746);
xnor U24642 (N_24642,N_16460,N_17938);
or U24643 (N_24643,N_16618,N_18001);
or U24644 (N_24644,N_15606,N_16301);
or U24645 (N_24645,N_15505,N_12939);
or U24646 (N_24646,N_18289,N_15725);
nand U24647 (N_24647,N_13526,N_14223);
nor U24648 (N_24648,N_15730,N_14467);
or U24649 (N_24649,N_14260,N_12590);
and U24650 (N_24650,N_17848,N_14139);
and U24651 (N_24651,N_15273,N_17932);
nand U24652 (N_24652,N_15054,N_13058);
nand U24653 (N_24653,N_17386,N_13852);
nor U24654 (N_24654,N_17392,N_15737);
nand U24655 (N_24655,N_15503,N_14383);
nor U24656 (N_24656,N_14399,N_16256);
or U24657 (N_24657,N_13161,N_13326);
nor U24658 (N_24658,N_15422,N_18234);
and U24659 (N_24659,N_16336,N_18449);
or U24660 (N_24660,N_17559,N_16498);
or U24661 (N_24661,N_12839,N_15089);
and U24662 (N_24662,N_17213,N_16495);
xor U24663 (N_24663,N_16990,N_18124);
nor U24664 (N_24664,N_15523,N_14701);
or U24665 (N_24665,N_14025,N_13510);
nor U24666 (N_24666,N_14900,N_17781);
nand U24667 (N_24667,N_14296,N_14414);
nand U24668 (N_24668,N_14011,N_17083);
nor U24669 (N_24669,N_17421,N_13645);
and U24670 (N_24670,N_17094,N_15300);
nand U24671 (N_24671,N_14001,N_16245);
nor U24672 (N_24672,N_15840,N_17205);
or U24673 (N_24673,N_13557,N_15590);
nand U24674 (N_24674,N_17008,N_14038);
and U24675 (N_24675,N_13231,N_15602);
nor U24676 (N_24676,N_14670,N_15557);
and U24677 (N_24677,N_18658,N_16274);
or U24678 (N_24678,N_18642,N_17838);
and U24679 (N_24679,N_14885,N_16058);
and U24680 (N_24680,N_17141,N_15662);
nor U24681 (N_24681,N_15352,N_13245);
nor U24682 (N_24682,N_18312,N_13741);
and U24683 (N_24683,N_14612,N_15616);
or U24684 (N_24684,N_18686,N_15925);
and U24685 (N_24685,N_14987,N_16351);
and U24686 (N_24686,N_14468,N_16501);
nor U24687 (N_24687,N_16772,N_16188);
and U24688 (N_24688,N_16015,N_15257);
or U24689 (N_24689,N_17772,N_14677);
and U24690 (N_24690,N_15141,N_14315);
nand U24691 (N_24691,N_13875,N_14903);
and U24692 (N_24692,N_15879,N_13121);
and U24693 (N_24693,N_16227,N_13852);
nor U24694 (N_24694,N_17883,N_16508);
and U24695 (N_24695,N_12740,N_13945);
and U24696 (N_24696,N_14705,N_16590);
nor U24697 (N_24697,N_16827,N_16874);
and U24698 (N_24698,N_17241,N_15791);
xnor U24699 (N_24699,N_14811,N_14912);
and U24700 (N_24700,N_14235,N_12787);
nor U24701 (N_24701,N_18406,N_16212);
or U24702 (N_24702,N_16833,N_17123);
or U24703 (N_24703,N_13078,N_14003);
or U24704 (N_24704,N_14706,N_18676);
or U24705 (N_24705,N_14428,N_14577);
nand U24706 (N_24706,N_16940,N_18621);
nand U24707 (N_24707,N_17084,N_12529);
or U24708 (N_24708,N_13866,N_15012);
and U24709 (N_24709,N_13895,N_13243);
nand U24710 (N_24710,N_13831,N_17053);
and U24711 (N_24711,N_15906,N_16543);
or U24712 (N_24712,N_14038,N_18280);
or U24713 (N_24713,N_14554,N_16872);
or U24714 (N_24714,N_15246,N_17880);
and U24715 (N_24715,N_17811,N_15741);
or U24716 (N_24716,N_16158,N_17858);
nand U24717 (N_24717,N_15231,N_17977);
nor U24718 (N_24718,N_18536,N_17419);
nand U24719 (N_24719,N_18164,N_17550);
and U24720 (N_24720,N_13138,N_18439);
and U24721 (N_24721,N_16814,N_17752);
nand U24722 (N_24722,N_16471,N_18714);
and U24723 (N_24723,N_16524,N_15672);
nor U24724 (N_24724,N_13582,N_17242);
nor U24725 (N_24725,N_14714,N_17189);
nor U24726 (N_24726,N_15989,N_14707);
or U24727 (N_24727,N_14183,N_15516);
or U24728 (N_24728,N_14945,N_16758);
nor U24729 (N_24729,N_17669,N_16220);
or U24730 (N_24730,N_16233,N_13765);
nor U24731 (N_24731,N_14665,N_13239);
nor U24732 (N_24732,N_16187,N_13025);
and U24733 (N_24733,N_16496,N_18049);
and U24734 (N_24734,N_18612,N_15295);
or U24735 (N_24735,N_17317,N_16523);
and U24736 (N_24736,N_18289,N_16290);
or U24737 (N_24737,N_17715,N_14065);
nand U24738 (N_24738,N_18224,N_16530);
nand U24739 (N_24739,N_15668,N_13766);
or U24740 (N_24740,N_14962,N_15540);
nand U24741 (N_24741,N_16563,N_17395);
and U24742 (N_24742,N_15397,N_14785);
and U24743 (N_24743,N_17627,N_16094);
nor U24744 (N_24744,N_17802,N_14589);
nor U24745 (N_24745,N_13600,N_15840);
and U24746 (N_24746,N_12676,N_16609);
and U24747 (N_24747,N_17882,N_15041);
and U24748 (N_24748,N_15972,N_12808);
nor U24749 (N_24749,N_16758,N_14101);
or U24750 (N_24750,N_17501,N_16632);
and U24751 (N_24751,N_17683,N_15306);
and U24752 (N_24752,N_12940,N_14884);
nand U24753 (N_24753,N_13436,N_13265);
and U24754 (N_24754,N_15856,N_14518);
or U24755 (N_24755,N_13618,N_17588);
and U24756 (N_24756,N_14662,N_17059);
or U24757 (N_24757,N_12834,N_13054);
nand U24758 (N_24758,N_15154,N_15246);
and U24759 (N_24759,N_17163,N_13250);
and U24760 (N_24760,N_14939,N_18185);
or U24761 (N_24761,N_15609,N_14219);
nor U24762 (N_24762,N_14778,N_14399);
nor U24763 (N_24763,N_17312,N_16432);
xor U24764 (N_24764,N_14199,N_14464);
nor U24765 (N_24765,N_12767,N_17086);
or U24766 (N_24766,N_17979,N_13662);
nor U24767 (N_24767,N_15676,N_12740);
and U24768 (N_24768,N_12529,N_15035);
and U24769 (N_24769,N_14686,N_13026);
nand U24770 (N_24770,N_13543,N_15794);
nand U24771 (N_24771,N_13728,N_13223);
or U24772 (N_24772,N_16992,N_13379);
nor U24773 (N_24773,N_18480,N_12625);
or U24774 (N_24774,N_14606,N_15930);
nand U24775 (N_24775,N_17092,N_16187);
and U24776 (N_24776,N_18503,N_13418);
or U24777 (N_24777,N_15011,N_15896);
and U24778 (N_24778,N_17696,N_13524);
or U24779 (N_24779,N_15688,N_16329);
or U24780 (N_24780,N_17843,N_16810);
nand U24781 (N_24781,N_17085,N_17582);
nand U24782 (N_24782,N_17809,N_17867);
nand U24783 (N_24783,N_13219,N_13704);
nor U24784 (N_24784,N_15694,N_12908);
and U24785 (N_24785,N_18707,N_16061);
or U24786 (N_24786,N_15415,N_17029);
or U24787 (N_24787,N_16118,N_16069);
or U24788 (N_24788,N_16463,N_16323);
nor U24789 (N_24789,N_18599,N_12554);
nand U24790 (N_24790,N_17893,N_13685);
and U24791 (N_24791,N_17287,N_18227);
nor U24792 (N_24792,N_14224,N_17960);
and U24793 (N_24793,N_17511,N_17904);
or U24794 (N_24794,N_16261,N_13402);
nand U24795 (N_24795,N_14707,N_17411);
nor U24796 (N_24796,N_14501,N_13796);
nor U24797 (N_24797,N_15431,N_16874);
nand U24798 (N_24798,N_17507,N_14657);
nand U24799 (N_24799,N_17966,N_12915);
nand U24800 (N_24800,N_14737,N_15094);
and U24801 (N_24801,N_17266,N_17296);
and U24802 (N_24802,N_17954,N_15988);
or U24803 (N_24803,N_12505,N_15795);
nor U24804 (N_24804,N_13942,N_18316);
nand U24805 (N_24805,N_18172,N_16632);
and U24806 (N_24806,N_18618,N_16234);
nand U24807 (N_24807,N_16405,N_13204);
and U24808 (N_24808,N_17648,N_14286);
or U24809 (N_24809,N_15792,N_18450);
nor U24810 (N_24810,N_17495,N_17062);
nor U24811 (N_24811,N_13759,N_16358);
nor U24812 (N_24812,N_13744,N_15718);
nor U24813 (N_24813,N_14066,N_18593);
and U24814 (N_24814,N_14296,N_14738);
nand U24815 (N_24815,N_13915,N_16196);
nand U24816 (N_24816,N_18554,N_15800);
nor U24817 (N_24817,N_12999,N_16933);
or U24818 (N_24818,N_17371,N_16309);
and U24819 (N_24819,N_13907,N_18565);
and U24820 (N_24820,N_14377,N_16081);
xnor U24821 (N_24821,N_15566,N_17916);
nand U24822 (N_24822,N_15686,N_14072);
and U24823 (N_24823,N_18692,N_16069);
nand U24824 (N_24824,N_14262,N_15320);
or U24825 (N_24825,N_18214,N_17835);
nor U24826 (N_24826,N_16430,N_13522);
nand U24827 (N_24827,N_14065,N_17396);
nor U24828 (N_24828,N_15293,N_18658);
or U24829 (N_24829,N_14846,N_18297);
or U24830 (N_24830,N_17505,N_14564);
nand U24831 (N_24831,N_18745,N_14517);
or U24832 (N_24832,N_15084,N_18017);
nor U24833 (N_24833,N_17106,N_17750);
or U24834 (N_24834,N_12609,N_15343);
nand U24835 (N_24835,N_15826,N_16888);
and U24836 (N_24836,N_14480,N_14512);
or U24837 (N_24837,N_17747,N_14902);
or U24838 (N_24838,N_14704,N_17996);
nand U24839 (N_24839,N_16531,N_16804);
and U24840 (N_24840,N_12821,N_14530);
and U24841 (N_24841,N_14239,N_12696);
or U24842 (N_24842,N_14282,N_18019);
or U24843 (N_24843,N_14073,N_14293);
nor U24844 (N_24844,N_14641,N_12572);
or U24845 (N_24845,N_18165,N_13814);
nand U24846 (N_24846,N_13755,N_16787);
or U24847 (N_24847,N_13430,N_14447);
nand U24848 (N_24848,N_14911,N_13086);
or U24849 (N_24849,N_18357,N_15217);
or U24850 (N_24850,N_17065,N_17542);
and U24851 (N_24851,N_13881,N_16646);
nand U24852 (N_24852,N_14559,N_14415);
nor U24853 (N_24853,N_14657,N_15026);
and U24854 (N_24854,N_16472,N_18419);
nor U24855 (N_24855,N_14013,N_18679);
nor U24856 (N_24856,N_16077,N_16976);
or U24857 (N_24857,N_17430,N_15384);
and U24858 (N_24858,N_17211,N_17427);
nor U24859 (N_24859,N_15444,N_13672);
nor U24860 (N_24860,N_13399,N_15549);
and U24861 (N_24861,N_17188,N_12543);
or U24862 (N_24862,N_13279,N_13620);
nand U24863 (N_24863,N_15642,N_13853);
nand U24864 (N_24864,N_13301,N_14876);
nand U24865 (N_24865,N_14140,N_12546);
nand U24866 (N_24866,N_14998,N_16771);
nor U24867 (N_24867,N_13621,N_15689);
nand U24868 (N_24868,N_12791,N_17839);
nor U24869 (N_24869,N_18169,N_16100);
or U24870 (N_24870,N_16165,N_17045);
nor U24871 (N_24871,N_13344,N_13260);
nand U24872 (N_24872,N_16056,N_16974);
and U24873 (N_24873,N_17506,N_18169);
or U24874 (N_24874,N_13931,N_13809);
or U24875 (N_24875,N_15440,N_12938);
and U24876 (N_24876,N_15790,N_17746);
and U24877 (N_24877,N_15787,N_15978);
nand U24878 (N_24878,N_18319,N_15071);
nand U24879 (N_24879,N_13946,N_16579);
or U24880 (N_24880,N_14575,N_15252);
nor U24881 (N_24881,N_17197,N_13039);
or U24882 (N_24882,N_12826,N_15689);
and U24883 (N_24883,N_13376,N_17620);
nor U24884 (N_24884,N_15152,N_15016);
or U24885 (N_24885,N_15360,N_16574);
nor U24886 (N_24886,N_16383,N_16438);
or U24887 (N_24887,N_13706,N_12534);
and U24888 (N_24888,N_18312,N_15347);
or U24889 (N_24889,N_14299,N_13776);
nor U24890 (N_24890,N_14507,N_18445);
xor U24891 (N_24891,N_17954,N_16415);
nand U24892 (N_24892,N_14506,N_13754);
and U24893 (N_24893,N_13180,N_16270);
or U24894 (N_24894,N_14141,N_15668);
nand U24895 (N_24895,N_18739,N_16554);
or U24896 (N_24896,N_15060,N_12575);
nor U24897 (N_24897,N_13546,N_18606);
nand U24898 (N_24898,N_17939,N_13541);
or U24899 (N_24899,N_14040,N_14319);
nand U24900 (N_24900,N_16424,N_18394);
nor U24901 (N_24901,N_14313,N_12847);
or U24902 (N_24902,N_17348,N_16214);
nor U24903 (N_24903,N_18557,N_13453);
or U24904 (N_24904,N_17876,N_12932);
or U24905 (N_24905,N_17326,N_16600);
nor U24906 (N_24906,N_14741,N_15162);
and U24907 (N_24907,N_12599,N_12739);
and U24908 (N_24908,N_18414,N_16552);
or U24909 (N_24909,N_14945,N_17317);
and U24910 (N_24910,N_15285,N_15397);
or U24911 (N_24911,N_13056,N_12773);
nand U24912 (N_24912,N_17845,N_16380);
and U24913 (N_24913,N_15411,N_17083);
or U24914 (N_24914,N_17917,N_14429);
or U24915 (N_24915,N_12864,N_18112);
nor U24916 (N_24916,N_16077,N_17174);
and U24917 (N_24917,N_13782,N_16858);
or U24918 (N_24918,N_16009,N_14990);
or U24919 (N_24919,N_14212,N_16755);
nand U24920 (N_24920,N_13919,N_13475);
nand U24921 (N_24921,N_13497,N_14521);
nor U24922 (N_24922,N_14484,N_14147);
nor U24923 (N_24923,N_13680,N_16561);
or U24924 (N_24924,N_13397,N_17338);
nand U24925 (N_24925,N_16081,N_17894);
nand U24926 (N_24926,N_18744,N_17997);
and U24927 (N_24927,N_18251,N_12929);
nor U24928 (N_24928,N_18632,N_15866);
nand U24929 (N_24929,N_15455,N_14609);
and U24930 (N_24930,N_17468,N_14894);
or U24931 (N_24931,N_13347,N_16500);
nor U24932 (N_24932,N_15800,N_16637);
and U24933 (N_24933,N_16214,N_17174);
nand U24934 (N_24934,N_13459,N_18691);
or U24935 (N_24935,N_18518,N_13303);
nor U24936 (N_24936,N_16160,N_16742);
or U24937 (N_24937,N_13819,N_16572);
nor U24938 (N_24938,N_17056,N_12676);
nand U24939 (N_24939,N_15444,N_15809);
or U24940 (N_24940,N_14047,N_12972);
and U24941 (N_24941,N_17475,N_16873);
nand U24942 (N_24942,N_18039,N_12917);
or U24943 (N_24943,N_14163,N_14407);
or U24944 (N_24944,N_14430,N_17273);
nor U24945 (N_24945,N_16085,N_14537);
or U24946 (N_24946,N_17512,N_13338);
nand U24947 (N_24947,N_17648,N_12816);
or U24948 (N_24948,N_18731,N_13483);
nand U24949 (N_24949,N_14863,N_18347);
and U24950 (N_24950,N_14557,N_17719);
or U24951 (N_24951,N_17610,N_18208);
nand U24952 (N_24952,N_16973,N_15617);
nor U24953 (N_24953,N_12972,N_18602);
nor U24954 (N_24954,N_16959,N_14836);
or U24955 (N_24955,N_12820,N_14446);
nand U24956 (N_24956,N_14792,N_15269);
xnor U24957 (N_24957,N_17741,N_18098);
and U24958 (N_24958,N_14789,N_14691);
and U24959 (N_24959,N_13580,N_13600);
nor U24960 (N_24960,N_17652,N_18329);
and U24961 (N_24961,N_14298,N_14117);
or U24962 (N_24962,N_16915,N_15001);
nand U24963 (N_24963,N_15712,N_15592);
or U24964 (N_24964,N_14670,N_13067);
nor U24965 (N_24965,N_13177,N_16697);
nand U24966 (N_24966,N_18279,N_18625);
nor U24967 (N_24967,N_17363,N_13823);
nor U24968 (N_24968,N_12627,N_18706);
xor U24969 (N_24969,N_17462,N_14079);
or U24970 (N_24970,N_17628,N_15210);
nor U24971 (N_24971,N_14638,N_17602);
nor U24972 (N_24972,N_12609,N_16494);
nand U24973 (N_24973,N_18699,N_13266);
nand U24974 (N_24974,N_14093,N_16297);
or U24975 (N_24975,N_17745,N_13315);
and U24976 (N_24976,N_12708,N_16253);
and U24977 (N_24977,N_13123,N_16005);
or U24978 (N_24978,N_15191,N_17017);
or U24979 (N_24979,N_17504,N_17368);
nand U24980 (N_24980,N_17395,N_16862);
nor U24981 (N_24981,N_13224,N_18586);
nand U24982 (N_24982,N_13769,N_18019);
nand U24983 (N_24983,N_17432,N_13059);
nand U24984 (N_24984,N_13563,N_13333);
and U24985 (N_24985,N_14733,N_14171);
nand U24986 (N_24986,N_14492,N_17665);
nor U24987 (N_24987,N_17948,N_12794);
nor U24988 (N_24988,N_17914,N_14758);
or U24989 (N_24989,N_13581,N_12902);
xor U24990 (N_24990,N_12861,N_17432);
nor U24991 (N_24991,N_17516,N_16478);
or U24992 (N_24992,N_12780,N_12765);
nor U24993 (N_24993,N_15180,N_17727);
or U24994 (N_24994,N_13249,N_16686);
nor U24995 (N_24995,N_15511,N_18738);
and U24996 (N_24996,N_15838,N_16241);
and U24997 (N_24997,N_14045,N_15812);
nand U24998 (N_24998,N_18566,N_18465);
or U24999 (N_24999,N_18377,N_14117);
nand UO_0 (O_0,N_20765,N_24892);
nor UO_1 (O_1,N_23675,N_21760);
and UO_2 (O_2,N_22385,N_24491);
nor UO_3 (O_3,N_23674,N_20599);
or UO_4 (O_4,N_24806,N_24968);
or UO_5 (O_5,N_23089,N_18881);
nor UO_6 (O_6,N_23000,N_23645);
nor UO_7 (O_7,N_21101,N_21861);
or UO_8 (O_8,N_24399,N_19723);
nand UO_9 (O_9,N_24655,N_21252);
nor UO_10 (O_10,N_19074,N_19530);
and UO_11 (O_11,N_24186,N_24605);
or UO_12 (O_12,N_20221,N_23498);
or UO_13 (O_13,N_20457,N_21331);
nor UO_14 (O_14,N_24206,N_19985);
nand UO_15 (O_15,N_21068,N_22742);
and UO_16 (O_16,N_23928,N_19899);
nand UO_17 (O_17,N_20962,N_20402);
and UO_18 (O_18,N_23287,N_22351);
nand UO_19 (O_19,N_20636,N_22034);
nand UO_20 (O_20,N_18988,N_19451);
or UO_21 (O_21,N_22074,N_22063);
and UO_22 (O_22,N_21881,N_21471);
or UO_23 (O_23,N_21132,N_22284);
nor UO_24 (O_24,N_24606,N_21805);
nor UO_25 (O_25,N_19466,N_22401);
nor UO_26 (O_26,N_20133,N_19916);
and UO_27 (O_27,N_24950,N_21496);
nand UO_28 (O_28,N_22184,N_19027);
nand UO_29 (O_29,N_24500,N_21555);
nand UO_30 (O_30,N_21350,N_20925);
or UO_31 (O_31,N_24735,N_19687);
nand UO_32 (O_32,N_19460,N_21369);
nor UO_33 (O_33,N_22528,N_19111);
nor UO_34 (O_34,N_19239,N_23256);
nor UO_35 (O_35,N_24585,N_20981);
or UO_36 (O_36,N_23460,N_24634);
or UO_37 (O_37,N_24397,N_22199);
or UO_38 (O_38,N_20440,N_19492);
or UO_39 (O_39,N_23319,N_24444);
or UO_40 (O_40,N_20776,N_24420);
and UO_41 (O_41,N_24984,N_24907);
nor UO_42 (O_42,N_23960,N_19395);
nand UO_43 (O_43,N_21097,N_20818);
nand UO_44 (O_44,N_20578,N_21173);
nand UO_45 (O_45,N_23078,N_19811);
and UO_46 (O_46,N_20008,N_21701);
or UO_47 (O_47,N_22209,N_19784);
or UO_48 (O_48,N_20680,N_20842);
or UO_49 (O_49,N_24107,N_24717);
and UO_50 (O_50,N_21014,N_18899);
and UO_51 (O_51,N_22053,N_21988);
nand UO_52 (O_52,N_18941,N_18978);
or UO_53 (O_53,N_22890,N_23916);
nand UO_54 (O_54,N_19310,N_20459);
and UO_55 (O_55,N_21951,N_19612);
and UO_56 (O_56,N_18750,N_18879);
nand UO_57 (O_57,N_18951,N_23998);
nand UO_58 (O_58,N_21931,N_21077);
nor UO_59 (O_59,N_22461,N_22843);
nand UO_60 (O_60,N_19750,N_19386);
and UO_61 (O_61,N_24249,N_23457);
nand UO_62 (O_62,N_19232,N_23889);
nor UO_63 (O_63,N_21591,N_24245);
nor UO_64 (O_64,N_23496,N_22277);
nor UO_65 (O_65,N_22878,N_19988);
nand UO_66 (O_66,N_24689,N_19447);
or UO_67 (O_67,N_23828,N_23357);
and UO_68 (O_68,N_24244,N_24346);
or UO_69 (O_69,N_23131,N_19198);
nand UO_70 (O_70,N_21636,N_18914);
nand UO_71 (O_71,N_22166,N_23023);
or UO_72 (O_72,N_19497,N_24729);
or UO_73 (O_73,N_18940,N_19375);
nor UO_74 (O_74,N_21593,N_20983);
or UO_75 (O_75,N_22368,N_23571);
or UO_76 (O_76,N_22410,N_18907);
nand UO_77 (O_77,N_21012,N_19088);
or UO_78 (O_78,N_21122,N_19862);
or UO_79 (O_79,N_23350,N_20786);
or UO_80 (O_80,N_19818,N_24364);
nand UO_81 (O_81,N_21544,N_22856);
or UO_82 (O_82,N_22397,N_23033);
and UO_83 (O_83,N_20860,N_21606);
or UO_84 (O_84,N_21687,N_21113);
nand UO_85 (O_85,N_24487,N_22172);
and UO_86 (O_86,N_23903,N_22934);
nor UO_87 (O_87,N_19880,N_21570);
and UO_88 (O_88,N_21052,N_20834);
nand UO_89 (O_89,N_22723,N_24144);
nand UO_90 (O_90,N_22235,N_19775);
and UO_91 (O_91,N_24303,N_21065);
or UO_92 (O_92,N_22904,N_18765);
and UO_93 (O_93,N_20760,N_22243);
or UO_94 (O_94,N_23567,N_23810);
or UO_95 (O_95,N_21958,N_20618);
or UO_96 (O_96,N_19156,N_20428);
nor UO_97 (O_97,N_20613,N_21312);
or UO_98 (O_98,N_19150,N_22588);
nand UO_99 (O_99,N_20126,N_21270);
or UO_100 (O_100,N_20731,N_23205);
and UO_101 (O_101,N_23341,N_22148);
and UO_102 (O_102,N_24123,N_23364);
nand UO_103 (O_103,N_19578,N_23862);
and UO_104 (O_104,N_22840,N_22605);
nor UO_105 (O_105,N_19514,N_24767);
nor UO_106 (O_106,N_21159,N_21415);
or UO_107 (O_107,N_21104,N_24507);
nor UO_108 (O_108,N_20381,N_23587);
nor UO_109 (O_109,N_22041,N_19914);
and UO_110 (O_110,N_20972,N_23672);
nand UO_111 (O_111,N_21664,N_20898);
nor UO_112 (O_112,N_19738,N_19149);
or UO_113 (O_113,N_18771,N_22771);
nand UO_114 (O_114,N_23080,N_22822);
and UO_115 (O_115,N_21454,N_19356);
and UO_116 (O_116,N_19052,N_19132);
nor UO_117 (O_117,N_19755,N_19203);
nand UO_118 (O_118,N_24895,N_21236);
nand UO_119 (O_119,N_22473,N_23215);
and UO_120 (O_120,N_22331,N_24292);
nand UO_121 (O_121,N_23973,N_19828);
nor UO_122 (O_122,N_22377,N_22699);
nand UO_123 (O_123,N_23744,N_23549);
or UO_124 (O_124,N_23171,N_23783);
and UO_125 (O_125,N_19978,N_18864);
nand UO_126 (O_126,N_22868,N_20890);
nor UO_127 (O_127,N_23879,N_19399);
or UO_128 (O_128,N_23584,N_21314);
or UO_129 (O_129,N_21961,N_23302);
nor UO_130 (O_130,N_20878,N_23663);
nor UO_131 (O_131,N_19291,N_20416);
nor UO_132 (O_132,N_19090,N_22295);
nor UO_133 (O_133,N_18963,N_19167);
and UO_134 (O_134,N_23667,N_23137);
nand UO_135 (O_135,N_22222,N_22242);
nand UO_136 (O_136,N_22884,N_22135);
nand UO_137 (O_137,N_22874,N_19333);
nor UO_138 (O_138,N_19147,N_22719);
nand UO_139 (O_139,N_23905,N_21876);
nand UO_140 (O_140,N_19876,N_22931);
nor UO_141 (O_141,N_21645,N_24589);
and UO_142 (O_142,N_18909,N_19691);
nor UO_143 (O_143,N_23884,N_18930);
or UO_144 (O_144,N_20749,N_24406);
or UO_145 (O_145,N_24023,N_23228);
and UO_146 (O_146,N_22753,N_23925);
and UO_147 (O_147,N_20741,N_19917);
nor UO_148 (O_148,N_21436,N_21420);
nor UO_149 (O_149,N_19494,N_21180);
or UO_150 (O_150,N_20280,N_24565);
and UO_151 (O_151,N_21199,N_19306);
or UO_152 (O_152,N_22881,N_23451);
and UO_153 (O_153,N_19973,N_23176);
nor UO_154 (O_154,N_22518,N_22975);
nor UO_155 (O_155,N_20059,N_23401);
nor UO_156 (O_156,N_21061,N_24704);
nor UO_157 (O_157,N_22767,N_24104);
nand UO_158 (O_158,N_24009,N_19801);
or UO_159 (O_159,N_24029,N_21624);
nor UO_160 (O_160,N_20173,N_22550);
nor UO_161 (O_161,N_21105,N_20443);
nand UO_162 (O_162,N_20614,N_20671);
nand UO_163 (O_163,N_21188,N_24548);
nor UO_164 (O_164,N_21321,N_23692);
and UO_165 (O_165,N_21184,N_22661);
nor UO_166 (O_166,N_20335,N_24925);
and UO_167 (O_167,N_24527,N_24948);
or UO_168 (O_168,N_19431,N_21397);
nand UO_169 (O_169,N_21348,N_20035);
or UO_170 (O_170,N_18984,N_22134);
and UO_171 (O_171,N_19429,N_21856);
nor UO_172 (O_172,N_21776,N_24665);
nor UO_173 (O_173,N_21774,N_21527);
nor UO_174 (O_174,N_21909,N_24996);
and UO_175 (O_175,N_19675,N_22180);
and UO_176 (O_176,N_24854,N_24642);
nor UO_177 (O_177,N_19703,N_22865);
and UO_178 (O_178,N_24870,N_24998);
nand UO_179 (O_179,N_23258,N_20552);
nand UO_180 (O_180,N_20110,N_22052);
and UO_181 (O_181,N_21970,N_23948);
nor UO_182 (O_182,N_20598,N_24198);
nor UO_183 (O_183,N_21452,N_21937);
and UO_184 (O_184,N_21536,N_21901);
or UO_185 (O_185,N_20142,N_22342);
nand UO_186 (O_186,N_24656,N_21578);
or UO_187 (O_187,N_24618,N_19142);
or UO_188 (O_188,N_24674,N_22972);
and UO_189 (O_189,N_20564,N_20120);
nor UO_190 (O_190,N_24416,N_22477);
nand UO_191 (O_191,N_23754,N_24307);
and UO_192 (O_192,N_19152,N_23867);
nand UO_193 (O_193,N_22191,N_20712);
nor UO_194 (O_194,N_21275,N_23230);
and UO_195 (O_195,N_21764,N_21064);
nand UO_196 (O_196,N_23740,N_20820);
nand UO_197 (O_197,N_23226,N_23468);
or UO_198 (O_198,N_24248,N_23238);
nand UO_199 (O_199,N_22775,N_19015);
and UO_200 (O_200,N_19556,N_23222);
nor UO_201 (O_201,N_22799,N_20411);
nor UO_202 (O_202,N_19279,N_22125);
nor UO_203 (O_203,N_22549,N_24766);
nand UO_204 (O_204,N_23144,N_22422);
and UO_205 (O_205,N_24869,N_19596);
or UO_206 (O_206,N_19062,N_19083);
or UO_207 (O_207,N_19947,N_24289);
nand UO_208 (O_208,N_24881,N_22221);
or UO_209 (O_209,N_24865,N_24372);
and UO_210 (O_210,N_19186,N_20768);
nand UO_211 (O_211,N_23559,N_20991);
or UO_212 (O_212,N_20990,N_21094);
and UO_213 (O_213,N_19734,N_22995);
nand UO_214 (O_214,N_23432,N_23293);
and UO_215 (O_215,N_20913,N_24679);
nand UO_216 (O_216,N_18897,N_19297);
nor UO_217 (O_217,N_20242,N_20829);
nor UO_218 (O_218,N_20306,N_24228);
or UO_219 (O_219,N_22254,N_18846);
nand UO_220 (O_220,N_21772,N_19528);
and UO_221 (O_221,N_24727,N_20727);
nor UO_222 (O_222,N_23373,N_23677);
nand UO_223 (O_223,N_24152,N_19676);
xnor UO_224 (O_224,N_24122,N_23619);
or UO_225 (O_225,N_18974,N_20263);
xnor UO_226 (O_226,N_23014,N_24290);
and UO_227 (O_227,N_24554,N_18763);
nand UO_228 (O_228,N_24038,N_23852);
nor UO_229 (O_229,N_24782,N_20295);
or UO_230 (O_230,N_24193,N_23169);
or UO_231 (O_231,N_21716,N_19573);
and UO_232 (O_232,N_19402,N_24083);
nor UO_233 (O_233,N_21387,N_24298);
or UO_234 (O_234,N_22894,N_20424);
or UO_235 (O_235,N_21470,N_22071);
or UO_236 (O_236,N_24989,N_20927);
or UO_237 (O_237,N_20294,N_22914);
or UO_238 (O_238,N_23035,N_21254);
or UO_239 (O_239,N_23052,N_23513);
or UO_240 (O_240,N_20436,N_22023);
or UO_241 (O_241,N_22713,N_22694);
and UO_242 (O_242,N_24539,N_21377);
or UO_243 (O_243,N_22412,N_23883);
nand UO_244 (O_244,N_22864,N_18815);
nand UO_245 (O_245,N_21417,N_22309);
and UO_246 (O_246,N_19075,N_19348);
and UO_247 (O_247,N_22375,N_22568);
nor UO_248 (O_248,N_21295,N_24811);
nor UO_249 (O_249,N_19362,N_20384);
or UO_250 (O_250,N_20177,N_21922);
and UO_251 (O_251,N_24498,N_21010);
and UO_252 (O_252,N_21965,N_21507);
and UO_253 (O_253,N_22077,N_22746);
or UO_254 (O_254,N_24916,N_24924);
and UO_255 (O_255,N_22535,N_20903);
nand UO_256 (O_256,N_22983,N_23262);
nor UO_257 (O_257,N_19694,N_23086);
or UO_258 (O_258,N_20445,N_20698);
nor UO_259 (O_259,N_21734,N_24293);
and UO_260 (O_260,N_24374,N_19454);
nor UO_261 (O_261,N_23771,N_23400);
or UO_262 (O_262,N_24235,N_23651);
or UO_263 (O_263,N_23168,N_19996);
nand UO_264 (O_264,N_24367,N_22157);
and UO_265 (O_265,N_19699,N_21674);
and UO_266 (O_266,N_20856,N_22198);
and UO_267 (O_267,N_22098,N_24440);
and UO_268 (O_268,N_22163,N_23272);
nor UO_269 (O_269,N_20137,N_20654);
and UO_270 (O_270,N_20066,N_24306);
nand UO_271 (O_271,N_22067,N_19215);
and UO_272 (O_272,N_22059,N_21375);
or UO_273 (O_273,N_20415,N_23485);
nand UO_274 (O_274,N_22882,N_24599);
or UO_275 (O_275,N_22030,N_21950);
nor UO_276 (O_276,N_24324,N_24779);
nand UO_277 (O_277,N_24714,N_20905);
and UO_278 (O_278,N_21247,N_22784);
nand UO_279 (O_279,N_20350,N_20260);
or UO_280 (O_280,N_20579,N_21859);
and UO_281 (O_281,N_24770,N_20471);
nand UO_282 (O_282,N_22489,N_21819);
and UO_283 (O_283,N_23402,N_24652);
or UO_284 (O_284,N_19457,N_23066);
or UO_285 (O_285,N_22658,N_21911);
nor UO_286 (O_286,N_19435,N_19638);
or UO_287 (O_287,N_23770,N_22122);
or UO_288 (O_288,N_21157,N_19318);
or UO_289 (O_289,N_20858,N_18993);
and UO_290 (O_290,N_24930,N_19821);
nor UO_291 (O_291,N_19473,N_21343);
and UO_292 (O_292,N_22248,N_23094);
nor UO_293 (O_293,N_24496,N_19382);
nand UO_294 (O_294,N_23776,N_20434);
or UO_295 (O_295,N_24211,N_20096);
nor UO_296 (O_296,N_23199,N_22371);
or UO_297 (O_297,N_21363,N_22569);
and UO_298 (O_298,N_20147,N_22193);
or UO_299 (O_299,N_22003,N_23027);
nand UO_300 (O_300,N_20511,N_20315);
and UO_301 (O_301,N_20451,N_23077);
nor UO_302 (O_302,N_22926,N_21647);
nand UO_303 (O_303,N_23465,N_21288);
and UO_304 (O_304,N_24824,N_20105);
or UO_305 (O_305,N_19854,N_24316);
nand UO_306 (O_306,N_21038,N_21755);
nor UO_307 (O_307,N_20462,N_23767);
and UO_308 (O_308,N_24976,N_19108);
and UO_309 (O_309,N_21661,N_20502);
nand UO_310 (O_310,N_21231,N_22420);
nor UO_311 (O_311,N_22596,N_21627);
nand UO_312 (O_312,N_18976,N_23611);
nand UO_313 (O_313,N_18912,N_23897);
nor UO_314 (O_314,N_19439,N_23792);
nand UO_315 (O_315,N_19120,N_18962);
and UO_316 (O_316,N_19436,N_21494);
nor UO_317 (O_317,N_24810,N_20634);
nor UO_318 (O_318,N_23885,N_23734);
nor UO_319 (O_319,N_21696,N_23607);
or UO_320 (O_320,N_21673,N_24200);
nand UO_321 (O_321,N_19491,N_23486);
nor UO_322 (O_322,N_22659,N_20193);
nand UO_323 (O_323,N_21004,N_19553);
nand UO_324 (O_324,N_23683,N_19354);
nor UO_325 (O_325,N_22306,N_21528);
nand UO_326 (O_326,N_24985,N_22324);
and UO_327 (O_327,N_21552,N_21724);
or UO_328 (O_328,N_20036,N_20156);
or UO_329 (O_329,N_22940,N_24624);
and UO_330 (O_330,N_23294,N_24260);
nand UO_331 (O_331,N_19325,N_24006);
or UO_332 (O_332,N_21437,N_22231);
or UO_333 (O_333,N_23655,N_21893);
nand UO_334 (O_334,N_20098,N_21500);
or UO_335 (O_335,N_24684,N_19419);
or UO_336 (O_336,N_20797,N_24032);
nor UO_337 (O_337,N_22600,N_20841);
nor UO_338 (O_338,N_22345,N_20746);
and UO_339 (O_339,N_22217,N_24213);
and UO_340 (O_340,N_19894,N_24343);
and UO_341 (O_341,N_18795,N_19741);
nand UO_342 (O_342,N_23214,N_21090);
and UO_343 (O_343,N_24345,N_23914);
and UO_344 (O_344,N_19790,N_22687);
nor UO_345 (O_345,N_21336,N_18994);
nand UO_346 (O_346,N_20086,N_22548);
or UO_347 (O_347,N_24419,N_19406);
and UO_348 (O_348,N_22520,N_20321);
or UO_349 (O_349,N_21468,N_24120);
and UO_350 (O_350,N_23524,N_21813);
and UO_351 (O_351,N_20267,N_21341);
nand UO_352 (O_352,N_24489,N_22635);
nand UO_353 (O_353,N_24282,N_24541);
and UO_354 (O_354,N_19305,N_24163);
or UO_355 (O_355,N_21986,N_19848);
and UO_356 (O_356,N_18852,N_23836);
nor UO_357 (O_357,N_22611,N_23411);
and UO_358 (O_358,N_22019,N_18863);
nor UO_359 (O_359,N_23251,N_21934);
nand UO_360 (O_360,N_21971,N_18786);
nor UO_361 (O_361,N_22989,N_20136);
or UO_362 (O_362,N_21581,N_20607);
nand UO_363 (O_363,N_19885,N_23352);
or UO_364 (O_364,N_21839,N_23068);
nor UO_365 (O_365,N_20718,N_21932);
nand UO_366 (O_366,N_24961,N_21884);
and UO_367 (O_367,N_24871,N_24941);
nand UO_368 (O_368,N_19913,N_19507);
nand UO_369 (O_369,N_21845,N_20076);
and UO_370 (O_370,N_24012,N_22114);
nand UO_371 (O_371,N_22440,N_22104);
nor UO_372 (O_372,N_21587,N_24903);
nand UO_373 (O_373,N_24394,N_19041);
nor UO_374 (O_374,N_21968,N_21668);
or UO_375 (O_375,N_23437,N_18900);
nand UO_376 (O_376,N_22128,N_22445);
or UO_377 (O_377,N_24312,N_18992);
and UO_378 (O_378,N_24972,N_20380);
and UO_379 (O_379,N_21583,N_24271);
and UO_380 (O_380,N_21690,N_21510);
nor UO_381 (O_381,N_21823,N_22218);
nor UO_382 (O_382,N_19277,N_20220);
nand UO_383 (O_383,N_24567,N_24993);
nor UO_384 (O_384,N_22498,N_21498);
and UO_385 (O_385,N_24338,N_22824);
nor UO_386 (O_386,N_24061,N_22138);
nand UO_387 (O_387,N_19760,N_23083);
nor UO_388 (O_388,N_22112,N_22612);
and UO_389 (O_389,N_24995,N_20969);
nand UO_390 (O_390,N_22102,N_20734);
and UO_391 (O_391,N_24758,N_20201);
and UO_392 (O_392,N_22066,N_23387);
nand UO_393 (O_393,N_19896,N_24167);
nand UO_394 (O_394,N_20009,N_23664);
nand UO_395 (O_395,N_21781,N_20234);
or UO_396 (O_396,N_24273,N_23508);
nand UO_397 (O_397,N_20500,N_24469);
and UO_398 (O_398,N_19991,N_20893);
and UO_399 (O_399,N_21258,N_20849);
nand UO_400 (O_400,N_19846,N_24938);
and UO_401 (O_401,N_23616,N_23138);
nand UO_402 (O_402,N_21463,N_20674);
or UO_403 (O_403,N_19192,N_22585);
nand UO_404 (O_404,N_23946,N_21039);
nor UO_405 (O_405,N_23381,N_22298);
or UO_406 (O_406,N_19833,N_23864);
nor UO_407 (O_407,N_21358,N_19272);
nor UO_408 (O_408,N_19891,N_22078);
and UO_409 (O_409,N_21410,N_20493);
and UO_410 (O_410,N_22213,N_20010);
nand UO_411 (O_411,N_22757,N_23860);
and UO_412 (O_412,N_19806,N_23386);
nor UO_413 (O_413,N_23536,N_21187);
nor UO_414 (O_414,N_20997,N_21542);
or UO_415 (O_415,N_22762,N_21633);
nand UO_416 (O_416,N_20425,N_24400);
nand UO_417 (O_417,N_24463,N_24602);
and UO_418 (O_418,N_19179,N_23330);
nor UO_419 (O_419,N_21733,N_22072);
or UO_420 (O_420,N_20043,N_20284);
nand UO_421 (O_421,N_22603,N_20496);
or UO_422 (O_422,N_24021,N_19365);
or UO_423 (O_423,N_20720,N_23097);
and UO_424 (O_424,N_20401,N_20696);
nand UO_425 (O_425,N_21216,N_20633);
nor UO_426 (O_426,N_19523,N_23165);
nor UO_427 (O_427,N_21183,N_24650);
nor UO_428 (O_428,N_22815,N_22821);
or UO_429 (O_429,N_22976,N_19904);
or UO_430 (O_430,N_20737,N_22674);
nand UO_431 (O_431,N_19739,N_21704);
or UO_432 (O_432,N_24351,N_20024);
xor UO_433 (O_433,N_21582,N_19593);
or UO_434 (O_434,N_23842,N_20965);
nand UO_435 (O_435,N_21391,N_19166);
or UO_436 (O_436,N_24016,N_19314);
and UO_437 (O_437,N_21834,N_23535);
nand UO_438 (O_438,N_21866,N_18925);
nor UO_439 (O_439,N_21054,N_22921);
nand UO_440 (O_440,N_24888,N_24118);
or UO_441 (O_441,N_23344,N_19216);
nor UO_442 (O_442,N_19855,N_21917);
nand UO_443 (O_443,N_24035,N_22725);
nand UO_444 (O_444,N_24196,N_19069);
nand UO_445 (O_445,N_20183,N_19839);
and UO_446 (O_446,N_20788,N_21170);
and UO_447 (O_447,N_21305,N_20054);
and UO_448 (O_448,N_19600,N_23185);
or UO_449 (O_449,N_19674,N_22705);
and UO_450 (O_450,N_20164,N_22977);
nor UO_451 (O_451,N_18830,N_24558);
and UO_452 (O_452,N_24571,N_23115);
nand UO_453 (O_453,N_24090,N_24612);
or UO_454 (O_454,N_20419,N_20794);
nor UO_455 (O_455,N_22798,N_22094);
and UO_456 (O_456,N_19282,N_22374);
or UO_457 (O_457,N_19469,N_20146);
nand UO_458 (O_458,N_23718,N_19199);
nor UO_459 (O_459,N_18813,N_23067);
and UO_460 (O_460,N_22090,N_23993);
and UO_461 (O_461,N_20334,N_23275);
or UO_462 (O_462,N_24174,N_20119);
and UO_463 (O_463,N_23626,N_21034);
or UO_464 (O_464,N_21364,N_24771);
nand UO_465 (O_465,N_22282,N_20687);
nand UO_466 (O_466,N_22182,N_24636);
or UO_467 (O_467,N_24076,N_24043);
nor UO_468 (O_468,N_22407,N_21092);
nor UO_469 (O_469,N_23530,N_19563);
nor UO_470 (O_470,N_20787,N_22500);
and UO_471 (O_471,N_22836,N_24720);
nand UO_472 (O_472,N_23714,N_19815);
nand UO_473 (O_473,N_22637,N_24834);
and UO_474 (O_474,N_20057,N_24763);
nand UO_475 (O_475,N_22085,N_19471);
nand UO_476 (O_476,N_19420,N_19928);
nand UO_477 (O_477,N_23087,N_20288);
or UO_478 (O_478,N_22204,N_23659);
or UO_479 (O_479,N_21066,N_24979);
and UO_480 (O_480,N_22149,N_20979);
and UO_481 (O_481,N_21425,N_19048);
or UO_482 (O_482,N_22850,N_24693);
and UO_483 (O_483,N_19433,N_23609);
nor UO_484 (O_484,N_21440,N_23826);
nor UO_485 (O_485,N_20733,N_20084);
and UO_486 (O_486,N_21297,N_22153);
nand UO_487 (O_487,N_23184,N_22920);
and UO_488 (O_488,N_22599,N_24891);
nand UO_489 (O_489,N_23252,N_23753);
or UO_490 (O_490,N_23875,N_23976);
nor UO_491 (O_491,N_21462,N_24615);
or UO_492 (O_492,N_18980,N_21210);
nand UO_493 (O_493,N_24184,N_22404);
nor UO_494 (O_494,N_20246,N_20346);
nand UO_495 (O_495,N_18956,N_20199);
and UO_496 (O_496,N_23469,N_22393);
and UO_497 (O_497,N_19789,N_23996);
xor UO_498 (O_498,N_23190,N_20376);
nand UO_499 (O_499,N_24899,N_24927);
or UO_500 (O_500,N_23721,N_21164);
nand UO_501 (O_501,N_23612,N_22390);
nor UO_502 (O_502,N_20840,N_19577);
nor UO_503 (O_503,N_21726,N_21757);
and UO_504 (O_504,N_20883,N_20782);
nor UO_505 (O_505,N_21708,N_21790);
or UO_506 (O_506,N_24027,N_24268);
and UO_507 (O_507,N_22980,N_22991);
or UO_508 (O_508,N_19918,N_24874);
nand UO_509 (O_509,N_24819,N_21298);
nand UO_510 (O_510,N_21233,N_23371);
nand UO_511 (O_511,N_22755,N_23504);
or UO_512 (O_512,N_19072,N_23463);
nor UO_513 (O_513,N_22618,N_23523);
nor UO_514 (O_514,N_24868,N_20602);
nor UO_515 (O_515,N_19881,N_22591);
nor UO_516 (O_516,N_19057,N_22766);
or UO_517 (O_517,N_20964,N_23906);
nand UO_518 (O_518,N_21530,N_22304);
nor UO_519 (O_519,N_18756,N_20846);
nand UO_520 (O_520,N_24926,N_20854);
nor UO_521 (O_521,N_19458,N_24134);
nand UO_522 (O_522,N_23271,N_20819);
nand UO_523 (O_523,N_19540,N_24457);
nor UO_524 (O_524,N_22139,N_24386);
and UO_525 (O_525,N_19634,N_23269);
and UO_526 (O_526,N_21574,N_22210);
nor UO_527 (O_527,N_20413,N_20866);
or UO_528 (O_528,N_21206,N_19586);
or UO_529 (O_529,N_24033,N_19778);
and UO_530 (O_530,N_23552,N_19478);
nand UO_531 (O_531,N_20711,N_19550);
or UO_532 (O_532,N_21131,N_23586);
or UO_533 (O_533,N_21995,N_21519);
or UO_534 (O_534,N_18990,N_24433);
or UO_535 (O_535,N_19210,N_21136);
nand UO_536 (O_536,N_20118,N_21863);
nor UO_537 (O_537,N_23121,N_21936);
nand UO_538 (O_538,N_23312,N_24915);
nor UO_539 (O_539,N_24809,N_23594);
nand UO_540 (O_540,N_24230,N_22318);
nor UO_541 (O_541,N_21511,N_24019);
and UO_542 (O_542,N_20966,N_23551);
and UO_543 (O_543,N_22642,N_22579);
nor UO_544 (O_544,N_22251,N_21482);
and UO_545 (O_545,N_21407,N_22126);
or UO_546 (O_546,N_21629,N_18904);
nor UO_547 (O_547,N_22534,N_19668);
nor UO_548 (O_548,N_23041,N_20536);
nor UO_549 (O_549,N_20676,N_23034);
and UO_550 (O_550,N_21637,N_24800);
and UO_551 (O_551,N_21124,N_22325);
nand UO_552 (O_552,N_19560,N_24086);
xor UO_553 (O_553,N_24096,N_20989);
nand UO_554 (O_554,N_22580,N_24906);
and UO_555 (O_555,N_20215,N_22910);
nor UO_556 (O_556,N_21488,N_24366);
and UO_557 (O_557,N_24817,N_21260);
nand UO_558 (O_558,N_24370,N_24588);
nand UO_559 (O_559,N_22680,N_24000);
nand UO_560 (O_560,N_23661,N_22932);
or UO_561 (O_561,N_19515,N_19817);
nor UO_562 (O_562,N_24195,N_19317);
or UO_563 (O_563,N_24951,N_19287);
nor UO_564 (O_564,N_22359,N_22729);
nor UO_565 (O_565,N_20894,N_21143);
nand UO_566 (O_566,N_21771,N_21443);
xnor UO_567 (O_567,N_21837,N_23181);
and UO_568 (O_568,N_24581,N_23188);
nand UO_569 (O_569,N_22337,N_20523);
and UO_570 (O_570,N_19412,N_20753);
nand UO_571 (O_571,N_19391,N_22168);
or UO_572 (O_572,N_21096,N_21860);
nor UO_573 (O_573,N_23557,N_19626);
nor UO_574 (O_574,N_24520,N_23556);
and UO_575 (O_575,N_23116,N_24034);
or UO_576 (O_576,N_23966,N_22089);
xor UO_577 (O_577,N_22514,N_21589);
nor UO_578 (O_578,N_22647,N_21345);
and UO_579 (O_579,N_22866,N_21631);
nor UO_580 (O_580,N_20252,N_21230);
nand UO_581 (O_581,N_20662,N_24887);
and UO_582 (O_582,N_23924,N_24802);
nand UO_583 (O_583,N_18759,N_22281);
or UO_584 (O_584,N_20940,N_19990);
nand UO_585 (O_585,N_24455,N_20907);
nor UO_586 (O_586,N_22455,N_23930);
nor UO_587 (O_587,N_24936,N_23365);
nand UO_588 (O_588,N_24521,N_23656);
and UO_589 (O_589,N_24451,N_24238);
nor UO_590 (O_590,N_20777,N_22038);
or UO_591 (O_591,N_22981,N_24672);
nor UO_592 (O_592,N_18872,N_20576);
or UO_593 (O_593,N_22927,N_19155);
nand UO_594 (O_594,N_23982,N_19234);
and UO_595 (O_595,N_21836,N_20115);
nor UO_596 (O_596,N_19986,N_19557);
and UO_597 (O_597,N_21458,N_20683);
nand UO_598 (O_598,N_20393,N_22383);
and UO_599 (O_599,N_24205,N_19543);
and UO_600 (O_600,N_19262,N_21703);
nor UO_601 (O_601,N_19976,N_22115);
nor UO_602 (O_602,N_22257,N_23938);
and UO_603 (O_603,N_20895,N_22413);
or UO_604 (O_604,N_24465,N_23913);
nand UO_605 (O_605,N_20938,N_24363);
nand UO_606 (O_606,N_23853,N_19281);
and UO_607 (O_607,N_20216,N_24681);
or UO_608 (O_608,N_23355,N_19380);
or UO_609 (O_609,N_24830,N_18966);
and UO_610 (O_610,N_21824,N_23809);
nand UO_611 (O_611,N_19463,N_22923);
and UO_612 (O_612,N_21071,N_23084);
and UO_613 (O_613,N_24667,N_18917);
and UO_614 (O_614,N_19408,N_23636);
nand UO_615 (O_615,N_21818,N_19746);
nor UO_616 (O_616,N_19525,N_22091);
and UO_617 (O_617,N_21179,N_22169);
nor UO_618 (O_618,N_23697,N_21365);
or UO_619 (O_619,N_24795,N_24572);
and UO_620 (O_620,N_18973,N_20487);
and UO_621 (O_621,N_19953,N_22226);
nor UO_622 (O_622,N_24078,N_20495);
nor UO_623 (O_623,N_19025,N_22435);
nor UO_624 (O_624,N_19432,N_22544);
nor UO_625 (O_625,N_20808,N_21318);
or UO_626 (O_626,N_18995,N_21380);
nand UO_627 (O_627,N_23348,N_22967);
nand UO_628 (O_628,N_19587,N_23446);
nor UO_629 (O_629,N_21939,N_24328);
nor UO_630 (O_630,N_19009,N_20862);
nor UO_631 (O_631,N_24214,N_23336);
nor UO_632 (O_632,N_23992,N_23648);
and UO_633 (O_633,N_23781,N_20984);
and UO_634 (O_634,N_23849,N_23475);
nand UO_635 (O_635,N_20286,N_24917);
or UO_636 (O_636,N_24431,N_20960);
or UO_637 (O_637,N_23687,N_22696);
nor UO_638 (O_638,N_24039,N_21277);
nand UO_639 (O_639,N_20229,N_19427);
and UO_640 (O_640,N_21626,N_19168);
and UO_641 (O_641,N_23983,N_20655);
and UO_642 (O_642,N_24007,N_19319);
and UO_643 (O_643,N_23494,N_22205);
and UO_644 (O_644,N_20591,N_23830);
nand UO_645 (O_645,N_20557,N_20888);
or UO_646 (O_646,N_19517,N_21361);
nand UO_647 (O_647,N_20512,N_22652);
nand UO_648 (O_648,N_22315,N_23732);
nand UO_649 (O_649,N_22174,N_19893);
and UO_650 (O_650,N_22510,N_22414);
and UO_651 (O_651,N_19014,N_24897);
or UO_652 (O_652,N_19171,N_22382);
nand UO_653 (O_653,N_21219,N_23241);
and UO_654 (O_654,N_21993,N_23383);
nor UO_655 (O_655,N_22769,N_18843);
nor UO_656 (O_656,N_24053,N_20929);
nor UO_657 (O_657,N_21347,N_20278);
nor UO_658 (O_658,N_20735,N_21622);
nand UO_659 (O_659,N_22847,N_19663);
nor UO_660 (O_660,N_20410,N_24052);
or UO_661 (O_661,N_21897,N_23491);
or UO_662 (O_662,N_21145,N_23384);
nor UO_663 (O_663,N_23742,N_23904);
nand UO_664 (O_664,N_22253,N_24576);
nand UO_665 (O_665,N_21729,N_22188);
nand UO_666 (O_666,N_22679,N_23265);
and UO_667 (O_667,N_20473,N_23015);
nand UO_668 (O_668,N_20538,N_23461);
nor UO_669 (O_669,N_22565,N_20392);
or UO_670 (O_670,N_23391,N_23324);
nand UO_671 (O_671,N_23777,N_24492);
nand UO_672 (O_672,N_20917,N_24922);
or UO_673 (O_673,N_21329,N_22763);
or UO_674 (O_674,N_20170,N_20601);
or UO_675 (O_675,N_19542,N_24755);
or UO_676 (O_676,N_20593,N_21251);
nor UO_677 (O_677,N_23308,N_21503);
and UO_678 (O_678,N_21838,N_21870);
and UO_679 (O_679,N_22870,N_21568);
or UO_680 (O_680,N_21955,N_22262);
nand UO_681 (O_681,N_24402,N_19858);
nor UO_682 (O_682,N_24531,N_22717);
nor UO_683 (O_683,N_20677,N_22291);
nor UO_684 (O_684,N_18901,N_21609);
nand UO_685 (O_685,N_24511,N_20980);
and UO_686 (O_686,N_23686,N_24827);
and UO_687 (O_687,N_21080,N_21902);
or UO_688 (O_688,N_19835,N_20919);
nor UO_689 (O_689,N_23354,N_19303);
or UO_690 (O_690,N_19221,N_21682);
or UO_691 (O_691,N_20070,N_20742);
nor UO_692 (O_692,N_18935,N_20574);
nand UO_693 (O_693,N_24659,N_19226);
or UO_694 (O_694,N_19685,N_19360);
and UO_695 (O_695,N_24099,N_21411);
nor UO_696 (O_696,N_24317,N_24106);
nor UO_697 (O_697,N_22136,N_19335);
nand UO_698 (O_698,N_23440,N_21028);
and UO_699 (O_699,N_22178,N_22482);
nor UO_700 (O_700,N_21031,N_21656);
nor UO_701 (O_701,N_23788,N_22517);
or UO_702 (O_702,N_24327,N_19804);
nand UO_703 (O_703,N_22432,N_19308);
and UO_704 (O_704,N_24705,N_23789);
nor UO_705 (O_705,N_20791,N_23456);
nand UO_706 (O_706,N_21560,N_21050);
nor UO_707 (O_707,N_22802,N_24158);
or UO_708 (O_708,N_19561,N_20936);
nor UO_709 (O_709,N_19126,N_20505);
nand UO_710 (O_710,N_19650,N_19081);
xor UO_711 (O_711,N_18833,N_19982);
and UO_712 (O_712,N_21871,N_19707);
nand UO_713 (O_713,N_20967,N_21310);
or UO_714 (O_714,N_21709,N_24932);
and UO_715 (O_715,N_21573,N_23146);
or UO_716 (O_716,N_22527,N_22279);
nor UO_717 (O_717,N_24333,N_19964);
or UO_718 (O_718,N_20504,N_21161);
nor UO_719 (O_719,N_19337,N_21702);
or UO_720 (O_720,N_23422,N_24886);
or UO_721 (O_721,N_19558,N_23926);
nand UO_722 (O_722,N_23338,N_24820);
or UO_723 (O_723,N_23007,N_19309);
or UO_724 (O_724,N_21453,N_21195);
nor UO_725 (O_725,N_22389,N_23236);
nor UO_726 (O_726,N_19640,N_20046);
nor UO_727 (O_727,N_21473,N_19865);
and UO_728 (O_728,N_19665,N_19647);
or UO_729 (O_729,N_23246,N_19263);
and UO_730 (O_730,N_21205,N_20901);
or UO_731 (O_731,N_24449,N_21502);
nor UO_732 (O_732,N_24647,N_19901);
or UO_733 (O_733,N_21176,N_24743);
and UO_734 (O_734,N_19390,N_22502);
nand UO_735 (O_735,N_23538,N_19629);
and UO_736 (O_736,N_20111,N_20114);
xnor UO_737 (O_737,N_19264,N_20627);
and UO_738 (O_738,N_21652,N_22590);
or UO_739 (O_739,N_20207,N_22559);
nor UO_740 (O_740,N_24165,N_21960);
and UO_741 (O_741,N_21087,N_22054);
or UO_742 (O_742,N_20241,N_23970);
or UO_743 (O_743,N_19946,N_22488);
nand UO_744 (O_744,N_19030,N_22589);
nor UO_745 (O_745,N_19255,N_21135);
or UO_746 (O_746,N_20853,N_20514);
nor UO_747 (O_747,N_18919,N_18888);
nor UO_748 (O_748,N_23449,N_22715);
nand UO_749 (O_749,N_22439,N_21356);
nor UO_750 (O_750,N_22770,N_21337);
or UO_751 (O_751,N_24908,N_23517);
nand UO_752 (O_752,N_19595,N_20912);
and UO_753 (O_753,N_21431,N_20722);
nor UO_754 (O_754,N_23772,N_21478);
and UO_755 (O_755,N_19623,N_24805);
xor UO_756 (O_756,N_21785,N_20461);
nor UO_757 (O_757,N_24774,N_24975);
and UO_758 (O_758,N_19312,N_19227);
nand UO_759 (O_759,N_20986,N_23931);
nor UO_760 (O_760,N_20957,N_24586);
nand UO_761 (O_761,N_23418,N_23315);
or UO_762 (O_762,N_23179,N_24721);
or UO_763 (O_763,N_20752,N_23473);
nor UO_764 (O_764,N_22310,N_19231);
or UO_765 (O_765,N_21404,N_19829);
or UO_766 (O_766,N_22442,N_20045);
or UO_767 (O_767,N_19401,N_19237);
or UO_768 (O_768,N_24553,N_20153);
nand UO_769 (O_769,N_19984,N_22379);
or UO_770 (O_770,N_21432,N_22055);
nor UO_771 (O_771,N_23815,N_21238);
nor UO_772 (O_772,N_23910,N_22745);
nand UO_773 (O_773,N_20441,N_23602);
nand UO_774 (O_774,N_24592,N_20454);
nand UO_775 (O_775,N_20802,N_22244);
or UO_776 (O_776,N_20172,N_24724);
nand UO_777 (O_777,N_18855,N_20583);
nand UO_778 (O_778,N_23243,N_19275);
nor UO_779 (O_779,N_19934,N_22880);
nand UO_780 (O_780,N_19810,N_21241);
and UO_781 (O_781,N_21620,N_22552);
nand UO_782 (O_782,N_23150,N_24716);
and UO_783 (O_783,N_21450,N_20328);
and UO_784 (O_784,N_23896,N_19350);
nand UO_785 (O_785,N_19735,N_23444);
nor UO_786 (O_786,N_20621,N_23614);
nor UO_787 (O_787,N_23285,N_19748);
nor UO_788 (O_788,N_23075,N_24526);
nand UO_789 (O_789,N_21487,N_22893);
nor UO_790 (O_790,N_20001,N_24172);
and UO_791 (O_791,N_22595,N_19056);
or UO_792 (O_792,N_19219,N_23593);
nand UO_793 (O_793,N_20298,N_19849);
or UO_794 (O_794,N_20304,N_19797);
nand UO_795 (O_795,N_20659,N_21894);
and UO_796 (O_796,N_23588,N_24300);
nand UO_797 (O_797,N_22357,N_23142);
and UO_798 (O_798,N_20358,N_19658);
nor UO_799 (O_799,N_24192,N_22959);
or UO_800 (O_800,N_21767,N_19185);
nor UO_801 (O_801,N_19603,N_24013);
nor UO_802 (O_802,N_21915,N_22311);
or UO_803 (O_803,N_21049,N_23527);
and UO_804 (O_804,N_20789,N_24997);
nand UO_805 (O_805,N_22430,N_19278);
nor UO_806 (O_806,N_20682,N_21634);
nor UO_807 (O_807,N_22519,N_21381);
and UO_808 (O_808,N_20619,N_23309);
nor UO_809 (O_809,N_21197,N_21671);
nand UO_810 (O_810,N_23237,N_23711);
or UO_811 (O_811,N_23572,N_20437);
nand UO_812 (O_812,N_20269,N_23745);
or UO_813 (O_813,N_23466,N_21280);
nand UO_814 (O_814,N_22644,N_19823);
or UO_815 (O_815,N_22272,N_24269);
or UO_816 (O_816,N_21426,N_22280);
or UO_817 (O_817,N_19915,N_22734);
nand UO_818 (O_818,N_21806,N_20464);
or UO_819 (O_819,N_23868,N_22669);
or UO_820 (O_820,N_20844,N_20793);
or UO_821 (O_821,N_22999,N_20541);
nand UO_822 (O_822,N_23577,N_24462);
or UO_823 (O_823,N_22170,N_22070);
or UO_824 (O_824,N_23940,N_22956);
or UO_825 (O_825,N_21607,N_20049);
and UO_826 (O_826,N_22269,N_20418);
and UO_827 (O_827,N_22754,N_19396);
nand UO_828 (O_828,N_22787,N_24285);
nand UO_829 (O_829,N_21684,N_18876);
nor UO_830 (O_830,N_23701,N_24559);
or UO_831 (O_831,N_22451,N_22845);
and UO_832 (O_832,N_19265,N_23854);
or UO_833 (O_833,N_19922,N_23986);
or UO_834 (O_834,N_20700,N_21869);
or UO_835 (O_835,N_19258,N_19448);
or UO_836 (O_836,N_19747,N_23666);
nor UO_837 (O_837,N_23065,N_24815);
nor UO_838 (O_838,N_23671,N_23927);
nor UO_839 (O_839,N_24730,N_24879);
or UO_840 (O_840,N_19089,N_23113);
nand UO_841 (O_841,N_21543,N_20590);
xor UO_842 (O_842,N_23710,N_24383);
nor UO_843 (O_843,N_23347,N_22364);
and UO_844 (O_844,N_22245,N_22366);
and UO_845 (O_845,N_20719,N_22758);
and UO_846 (O_846,N_24227,N_20726);
nand UO_847 (O_847,N_20909,N_23773);
xnor UO_848 (O_848,N_24988,N_19224);
nand UO_849 (O_849,N_20432,N_21385);
and UO_850 (O_850,N_19611,N_19423);
nand UO_851 (O_851,N_19582,N_20078);
or UO_852 (O_852,N_24713,N_24785);
nor UO_853 (O_853,N_21118,N_19956);
and UO_854 (O_854,N_18875,N_20880);
nor UO_855 (O_855,N_21883,N_21567);
and UO_856 (O_856,N_21362,N_18961);
and UO_857 (O_857,N_22973,N_19462);
and UO_858 (O_858,N_19481,N_20869);
nand UO_859 (O_859,N_22930,N_20870);
nand UO_860 (O_860,N_19417,N_22530);
or UO_861 (O_861,N_19585,N_24942);
and UO_862 (O_862,N_20080,N_20332);
or UO_863 (O_863,N_23876,N_21207);
or UO_864 (O_864,N_23414,N_19134);
and UO_865 (O_865,N_23186,N_20446);
and UO_866 (O_866,N_22871,N_22685);
nor UO_867 (O_867,N_21725,N_21335);
nor UO_868 (O_868,N_21406,N_24410);
or UO_869 (O_869,N_21472,N_19389);
or UO_870 (O_870,N_21079,N_22604);
nand UO_871 (O_871,N_18831,N_24417);
nand UO_872 (O_872,N_24348,N_19957);
nand UO_873 (O_873,N_20283,N_22289);
or UO_874 (O_874,N_23154,N_23331);
or UO_875 (O_875,N_21151,N_22162);
and UO_876 (O_876,N_20305,N_24411);
nor UO_877 (O_877,N_22313,N_21203);
nand UO_878 (O_878,N_21693,N_19455);
nor UO_879 (O_879,N_23895,N_22782);
nor UO_880 (O_880,N_20482,N_22061);
nor UO_881 (O_881,N_20679,N_21250);
nor UO_882 (O_882,N_19965,N_21062);
nor UO_883 (O_883,N_19324,N_19017);
or UO_884 (O_884,N_20926,N_18754);
nand UO_885 (O_885,N_18867,N_21129);
and UO_886 (O_886,N_23439,N_20999);
nand UO_887 (O_887,N_21892,N_24421);
nand UO_888 (O_888,N_22419,N_23561);
or UO_889 (O_889,N_19633,N_22968);
and UO_890 (O_890,N_22141,N_24683);
and UO_891 (O_891,N_20522,N_19332);
nand UO_892 (O_892,N_23130,N_23975);
nor UO_893 (O_893,N_24628,N_24461);
nand UO_894 (O_894,N_20217,N_20852);
nand UO_895 (O_895,N_22877,N_23055);
nand UO_896 (O_896,N_23221,N_20996);
nor UO_897 (O_897,N_21189,N_19771);
nand UO_898 (O_898,N_22578,N_20341);
and UO_899 (O_899,N_19099,N_21679);
xor UO_900 (O_900,N_24794,N_20433);
nor UO_901 (O_901,N_20225,N_18957);
nor UO_902 (O_902,N_23580,N_20815);
nand UO_903 (O_903,N_19445,N_24133);
nand UO_904 (O_904,N_24506,N_24054);
nand UO_905 (O_905,N_21579,N_23025);
or UO_906 (O_906,N_22886,N_23208);
nor UO_907 (O_907,N_19843,N_22012);
and UO_908 (O_908,N_22859,N_21273);
nor UO_909 (O_909,N_21718,N_20656);
and UO_910 (O_910,N_23134,N_21735);
nand UO_911 (O_911,N_22320,N_23441);
nor UO_912 (O_912,N_19223,N_21885);
and UO_913 (O_913,N_23715,N_24127);
or UO_914 (O_914,N_22584,N_23886);
or UO_915 (O_915,N_22275,N_23694);
or UO_916 (O_916,N_23901,N_24084);
or UO_917 (O_917,N_18751,N_20339);
or UO_918 (O_918,N_18788,N_23640);
nand UO_919 (O_919,N_18819,N_19446);
nor UO_920 (O_920,N_23912,N_20822);
and UO_921 (O_921,N_23526,N_20756);
and UO_922 (O_922,N_22818,N_23048);
nor UO_923 (O_923,N_19902,N_21608);
nor UO_924 (O_924,N_19624,N_24332);
nand UO_925 (O_925,N_19501,N_24182);
or UO_926 (O_926,N_21501,N_21821);
or UO_927 (O_927,N_23500,N_19300);
or UO_928 (O_928,N_24640,N_24803);
or UO_929 (O_929,N_23964,N_18818);
nand UO_930 (O_930,N_20000,N_20721);
nand UO_931 (O_931,N_21505,N_19930);
or UO_932 (O_932,N_22928,N_21163);
or UO_933 (O_933,N_24991,N_23757);
nand UO_934 (O_934,N_24251,N_24164);
nor UO_935 (O_935,N_24858,N_24414);
or UO_936 (O_936,N_22150,N_19720);
or UO_937 (O_937,N_23794,N_21401);
or UO_938 (O_938,N_23969,N_23510);
nand UO_939 (O_939,N_22646,N_19019);
nand UO_940 (O_940,N_19477,N_24784);
or UO_941 (O_941,N_20900,N_22143);
nand UO_942 (O_942,N_20174,N_22862);
or UO_943 (O_943,N_19342,N_19535);
nand UO_944 (O_944,N_19125,N_21353);
and UO_945 (O_945,N_20403,N_23888);
and UO_946 (O_946,N_19713,N_22437);
nor UO_947 (O_947,N_21566,N_19882);
or UO_948 (O_948,N_23107,N_22471);
or UO_949 (O_949,N_19766,N_19207);
nor UO_950 (O_950,N_19467,N_24826);
nand UO_951 (O_951,N_20099,N_24751);
nand UO_952 (O_952,N_19710,N_21957);
xnor UO_953 (O_953,N_20396,N_23070);
or UO_954 (O_954,N_19374,N_24791);
or UO_955 (O_955,N_21830,N_21569);
nand UO_956 (O_956,N_21378,N_20617);
or UO_957 (O_957,N_23736,N_20472);
nand UO_958 (O_958,N_21360,N_21518);
nor UO_959 (O_959,N_22487,N_20902);
and UO_960 (O_960,N_20817,N_20365);
nor UO_961 (O_961,N_20356,N_24215);
nor UO_962 (O_962,N_23209,N_21166);
or UO_963 (O_963,N_24540,N_23657);
nor UO_964 (O_964,N_19673,N_24232);
nor UO_965 (O_965,N_24436,N_21677);
and UO_966 (O_966,N_19559,N_23578);
nand UO_967 (O_967,N_19409,N_22872);
and UO_968 (O_968,N_21602,N_22945);
nand UO_969 (O_969,N_19502,N_24011);
or UO_970 (O_970,N_24604,N_20264);
nor UO_971 (O_971,N_21516,N_22395);
or UO_972 (O_972,N_23274,N_23708);
nand UO_973 (O_973,N_20691,N_24187);
or UO_974 (O_974,N_18762,N_24093);
and UO_975 (O_975,N_21923,N_20087);
nor UO_976 (O_976,N_21978,N_18775);
or UO_977 (O_977,N_20647,N_24631);
nand UO_978 (O_978,N_23010,N_20747);
and UO_979 (O_979,N_23001,N_21059);
or UO_980 (O_980,N_19714,N_23300);
nand UO_981 (O_981,N_21994,N_20361);
and UO_982 (O_982,N_22774,N_20019);
or UO_983 (O_983,N_24745,N_22321);
and UO_984 (O_984,N_19376,N_19706);
or UO_985 (O_985,N_23629,N_23601);
nand UO_986 (O_986,N_20041,N_24673);
nor UO_987 (O_987,N_19442,N_19437);
and UO_988 (O_988,N_23442,N_22454);
nand UO_989 (O_989,N_22233,N_21742);
nand UO_990 (O_990,N_21935,N_24909);
nor UO_991 (O_991,N_19565,N_24790);
and UO_992 (O_992,N_23920,N_22841);
and UO_993 (O_993,N_23218,N_18861);
nor UO_994 (O_994,N_24534,N_22582);
and UO_995 (O_995,N_22467,N_22747);
nand UO_996 (O_996,N_23890,N_19245);
nand UO_997 (O_997,N_22545,N_22670);
or UO_998 (O_998,N_22147,N_20958);
nand UO_999 (O_999,N_21023,N_23119);
nor UO_1000 (O_1000,N_24059,N_19769);
and UO_1001 (O_1001,N_19851,N_21382);
nor UO_1002 (O_1002,N_21428,N_23952);
nor UO_1003 (O_1003,N_24046,N_21751);
or UO_1004 (O_1004,N_22974,N_22748);
nor UO_1005 (O_1005,N_21089,N_19567);
nand UO_1006 (O_1006,N_22381,N_21438);
and UO_1007 (O_1007,N_19002,N_24661);
or UO_1008 (O_1008,N_23128,N_23972);
nand UO_1009 (O_1009,N_22449,N_20478);
and UO_1010 (O_1010,N_20650,N_18996);
nand UO_1011 (O_1011,N_21374,N_24762);
nor UO_1012 (O_1012,N_24295,N_19434);
nor UO_1013 (O_1013,N_20448,N_20179);
or UO_1014 (O_1014,N_24898,N_21040);
nand UO_1015 (O_1015,N_22958,N_23295);
nor UO_1016 (O_1016,N_22614,N_22146);
nor UO_1017 (O_1017,N_23823,N_24657);
xnor UO_1018 (O_1018,N_22634,N_22287);
or UO_1019 (O_1019,N_19519,N_20744);
and UO_1020 (O_1020,N_19315,N_19133);
nand UO_1021 (O_1021,N_21888,N_23507);
and UO_1022 (O_1022,N_24468,N_24212);
or UO_1023 (O_1023,N_21814,N_24347);
nand UO_1024 (O_1024,N_23812,N_21256);
nand UO_1025 (O_1025,N_23741,N_22587);
or UO_1026 (O_1026,N_21854,N_21743);
nand UO_1027 (O_1027,N_19034,N_24336);
and UO_1028 (O_1028,N_24369,N_23547);
or UO_1029 (O_1029,N_19388,N_20134);
nand UO_1030 (O_1030,N_20668,N_20378);
or UO_1031 (O_1031,N_22511,N_23502);
nand UO_1032 (O_1032,N_23288,N_22516);
nor UO_1033 (O_1033,N_21396,N_20939);
or UO_1034 (O_1034,N_23314,N_23421);
nand UO_1035 (O_1035,N_20342,N_21712);
nand UO_1036 (O_1036,N_23790,N_24159);
nor UO_1037 (O_1037,N_22006,N_21201);
or UO_1038 (O_1038,N_21169,N_19809);
nand UO_1039 (O_1039,N_22058,N_24940);
and UO_1040 (O_1040,N_22607,N_23725);
and UO_1041 (O_1041,N_19989,N_22698);
nand UO_1042 (O_1042,N_21959,N_23737);
nand UO_1043 (O_1043,N_21149,N_22728);
or UO_1044 (O_1044,N_22338,N_19521);
and UO_1045 (O_1045,N_21429,N_19666);
or UO_1046 (O_1046,N_20175,N_21933);
or UO_1047 (O_1047,N_19532,N_24929);
nand UO_1048 (O_1048,N_23161,N_19043);
nor UO_1049 (O_1049,N_22808,N_23049);
and UO_1050 (O_1050,N_22509,N_24380);
or UO_1051 (O_1051,N_20836,N_19547);
nor UO_1052 (O_1052,N_19493,N_20157);
and UO_1053 (O_1053,N_24956,N_19980);
or UO_1054 (O_1054,N_24413,N_18837);
and UO_1055 (O_1055,N_23220,N_20743);
nor UO_1056 (O_1056,N_23847,N_21001);
nand UO_1057 (O_1057,N_19428,N_22227);
and UO_1058 (O_1058,N_22386,N_23892);
nor UO_1059 (O_1059,N_23676,N_20660);
nand UO_1060 (O_1060,N_20359,N_23022);
and UO_1061 (O_1061,N_18931,N_19449);
and UO_1062 (O_1062,N_23553,N_20366);
nor UO_1063 (O_1063,N_23627,N_24843);
or UO_1064 (O_1064,N_22951,N_20180);
nor UO_1065 (O_1065,N_20809,N_24799);
or UO_1066 (O_1066,N_23390,N_22394);
xnor UO_1067 (O_1067,N_19689,N_20703);
or UO_1068 (O_1068,N_19697,N_20587);
or UO_1069 (O_1069,N_19659,N_19726);
or UO_1070 (O_1070,N_23827,N_23795);
nand UO_1071 (O_1071,N_20005,N_21603);
and UO_1072 (O_1072,N_23484,N_22630);
nor UO_1073 (O_1073,N_24253,N_21435);
and UO_1074 (O_1074,N_19887,N_23764);
and UO_1075 (O_1075,N_23242,N_19060);
nand UO_1076 (O_1076,N_21338,N_23159);
nor UO_1077 (O_1077,N_21857,N_20723);
nand UO_1078 (O_1078,N_24831,N_20645);
nand UO_1079 (O_1079,N_23480,N_20558);
nand UO_1080 (O_1080,N_24801,N_24797);
and UO_1081 (O_1081,N_22483,N_20051);
and UO_1082 (O_1082,N_23785,N_22875);
or UO_1083 (O_1083,N_19012,N_23525);
nand UO_1084 (O_1084,N_23187,N_24116);
nor UO_1085 (O_1085,N_22617,N_19594);
nor UO_1086 (O_1086,N_20063,N_22613);
and UO_1087 (O_1087,N_19574,N_22801);
or UO_1088 (O_1088,N_19159,N_23207);
or UO_1089 (O_1089,N_23665,N_24079);
nor UO_1090 (O_1090,N_19398,N_20933);
or UO_1091 (O_1091,N_22867,N_23630);
and UO_1092 (O_1092,N_24472,N_24765);
nor UO_1093 (O_1093,N_20324,N_22228);
or UO_1094 (O_1094,N_19644,N_23392);
and UO_1095 (O_1095,N_19397,N_20083);
nand UO_1096 (O_1096,N_22131,N_18884);
nor UO_1097 (O_1097,N_23817,N_24970);
nor UO_1098 (O_1098,N_24741,N_21232);
nand UO_1099 (O_1099,N_22167,N_24177);
and UO_1100 (O_1100,N_20272,N_24600);
and UO_1101 (O_1101,N_22062,N_19511);
or UO_1102 (O_1102,N_20608,N_19538);
and UO_1103 (O_1103,N_22456,N_24203);
nand UO_1104 (O_1104,N_24884,N_23178);
and UO_1105 (O_1105,N_20644,N_21952);
nor UO_1106 (O_1106,N_18808,N_20253);
nor UO_1107 (O_1107,N_22812,N_21616);
and UO_1108 (O_1108,N_24931,N_23372);
xor UO_1109 (O_1109,N_21667,N_21737);
nor UO_1110 (O_1110,N_19966,N_24609);
and UO_1111 (O_1111,N_19782,N_22888);
and UO_1112 (O_1112,N_23499,N_23170);
nand UO_1113 (O_1113,N_21194,N_23542);
or UO_1114 (O_1114,N_23136,N_21921);
and UO_1115 (O_1115,N_23623,N_23098);
nand UO_1116 (O_1116,N_20148,N_20693);
and UO_1117 (O_1117,N_22293,N_22737);
or UO_1118 (O_1118,N_21752,N_19536);
nand UO_1119 (O_1119,N_23279,N_22964);
and UO_1120 (O_1120,N_20620,N_22918);
nand UO_1121 (O_1121,N_21017,N_24422);
nand UO_1122 (O_1122,N_20612,N_20145);
nor UO_1123 (O_1123,N_19472,N_21940);
or UO_1124 (O_1124,N_20707,N_21308);
or UO_1125 (O_1125,N_21303,N_19944);
nand UO_1126 (O_1126,N_23162,N_18752);
and UO_1127 (O_1127,N_20998,N_22691);
nand UO_1128 (O_1128,N_23404,N_24178);
and UO_1129 (O_1129,N_19688,N_22855);
nand UO_1130 (O_1130,N_22929,N_20549);
or UO_1131 (O_1131,N_23157,N_21590);
or UO_1132 (O_1132,N_22037,N_20839);
or UO_1133 (O_1133,N_22294,N_24946);
xor UO_1134 (O_1134,N_21102,N_23990);
nor UO_1135 (O_1135,N_18797,N_21697);
nor UO_1136 (O_1136,N_23047,N_23974);
nor UO_1137 (O_1137,N_22503,N_21676);
and UO_1138 (O_1138,N_24070,N_20023);
and UO_1139 (O_1139,N_21522,N_24538);
and UO_1140 (O_1140,N_21121,N_24570);
nand UO_1141 (O_1141,N_19932,N_19995);
nor UO_1142 (O_1142,N_21840,N_20071);
or UO_1143 (O_1143,N_20474,N_19130);
and UO_1144 (O_1144,N_21980,N_19725);
or UO_1145 (O_1145,N_20399,N_23759);
nand UO_1146 (O_1146,N_20928,N_21864);
nor UO_1147 (O_1147,N_23079,N_21833);
or UO_1148 (O_1148,N_19488,N_24669);
and UO_1149 (O_1149,N_20219,N_22212);
nor UO_1150 (O_1150,N_21808,N_22852);
or UO_1151 (O_1151,N_23965,N_21662);
nand UO_1152 (O_1152,N_24958,N_20992);
or UO_1153 (O_1153,N_19958,N_21198);
nor UO_1154 (O_1154,N_22402,N_19609);
and UO_1155 (O_1155,N_18766,N_22376);
nand UO_1156 (O_1156,N_19844,N_22982);
and UO_1157 (O_1157,N_20218,N_24889);
nor UO_1158 (O_1158,N_19840,N_19724);
or UO_1159 (O_1159,N_21359,N_20973);
or UO_1160 (O_1160,N_21658,N_24437);
and UO_1161 (O_1161,N_22505,N_23174);
and UO_1162 (O_1162,N_19566,N_23472);
or UO_1163 (O_1163,N_22329,N_19627);
nand UO_1164 (O_1164,N_24482,N_22008);
or UO_1165 (O_1165,N_19482,N_22361);
or UO_1166 (O_1166,N_22107,N_22779);
and UO_1167 (O_1167,N_23540,N_24732);
or UO_1168 (O_1168,N_19925,N_22796);
or UO_1169 (O_1169,N_24808,N_21846);
or UO_1170 (O_1170,N_18761,N_19018);
and UO_1171 (O_1171,N_19136,N_24773);
and UO_1172 (O_1172,N_24291,N_21974);
and UO_1173 (O_1173,N_21196,N_19021);
and UO_1174 (O_1174,N_24955,N_23668);
nand UO_1175 (O_1175,N_23204,N_22616);
nor UO_1176 (O_1176,N_22155,N_22948);
nor UO_1177 (O_1177,N_24041,N_18997);
and UO_1178 (O_1178,N_21540,N_23425);
nand UO_1179 (O_1179,N_19094,N_20184);
nor UO_1180 (O_1180,N_24512,N_23476);
nand UO_1181 (O_1181,N_21789,N_19864);
and UO_1182 (O_1182,N_22899,N_19575);
and UO_1183 (O_1183,N_24002,N_21490);
or UO_1184 (O_1184,N_19877,N_21384);
or UO_1185 (O_1185,N_22816,N_23303);
and UO_1186 (O_1186,N_21807,N_20692);
and UO_1187 (O_1187,N_23229,N_23999);
and UO_1188 (O_1188,N_20513,N_24302);
and UO_1189 (O_1189,N_21872,N_24190);
nand UO_1190 (O_1190,N_21067,N_19029);
nor UO_1191 (O_1191,N_24376,N_23006);
or UO_1192 (O_1192,N_19008,N_21486);
nand UO_1193 (O_1193,N_24485,N_23978);
nand UO_1194 (O_1194,N_23851,N_20771);
or UO_1195 (O_1195,N_21388,N_20189);
and UO_1196 (O_1196,N_18868,N_23152);
and UO_1197 (O_1197,N_24835,N_20697);
nor UO_1198 (O_1198,N_20383,N_20369);
and UO_1199 (O_1199,N_19054,N_21621);
or UO_1200 (O_1200,N_20439,N_23519);
nor UO_1201 (O_1201,N_24071,N_20847);
nand UO_1202 (O_1202,N_22547,N_20129);
nor UO_1203 (O_1203,N_19326,N_24037);
nand UO_1204 (O_1204,N_24629,N_21267);
nand UO_1205 (O_1205,N_22558,N_24686);
and UO_1206 (O_1206,N_23762,N_18971);
nor UO_1207 (O_1207,N_24513,N_23899);
nand UO_1208 (O_1208,N_19124,N_22660);
or UO_1209 (O_1209,N_22797,N_23393);
and UO_1210 (O_1210,N_24490,N_22283);
and UO_1211 (O_1211,N_24523,N_22017);
and UO_1212 (O_1212,N_22858,N_21403);
nand UO_1213 (O_1213,N_20649,N_24675);
nor UO_1214 (O_1214,N_20955,N_20003);
or UO_1215 (O_1215,N_22409,N_19169);
nor UO_1216 (O_1216,N_22900,N_19055);
nand UO_1217 (O_1217,N_22615,N_19832);
or UO_1218 (O_1218,N_20409,N_22978);
or UO_1219 (O_1219,N_23063,N_22593);
nand UO_1220 (O_1220,N_19678,N_23071);
and UO_1221 (O_1221,N_21053,N_20160);
or UO_1222 (O_1222,N_21600,N_23635);
and UO_1223 (O_1223,N_22905,N_22834);
nand UO_1224 (O_1224,N_22800,N_20658);
nor UO_1225 (O_1225,N_21650,N_22171);
nor UO_1226 (O_1226,N_20222,N_21117);
and UO_1227 (O_1227,N_22206,N_23739);
and UO_1228 (O_1228,N_20293,N_23193);
and UO_1229 (O_1229,N_18916,N_20355);
nand UO_1230 (O_1230,N_23305,N_23245);
nand UO_1231 (O_1231,N_23575,N_24170);
nand UO_1232 (O_1232,N_23706,N_21831);
and UO_1233 (O_1233,N_24453,N_19866);
nand UO_1234 (O_1234,N_19708,N_22436);
nand UO_1235 (O_1235,N_24443,N_19076);
nand UO_1236 (O_1236,N_21000,N_21956);
or UO_1237 (O_1237,N_20586,N_19347);
or UO_1238 (O_1238,N_20181,N_18753);
nand UO_1239 (O_1239,N_23670,N_21926);
nor UO_1240 (O_1240,N_20483,N_20489);
nor UO_1241 (O_1241,N_19727,N_19032);
and UO_1242 (O_1242,N_22076,N_19235);
or UO_1243 (O_1243,N_20127,N_24219);
or UO_1244 (O_1244,N_20832,N_21354);
and UO_1245 (O_1245,N_23802,N_22752);
nor UO_1246 (O_1246,N_21076,N_23297);
nor UO_1247 (O_1247,N_21272,N_23397);
and UO_1248 (O_1248,N_20918,N_23919);
nor UO_1249 (O_1249,N_21304,N_24426);
nand UO_1250 (O_1250,N_20835,N_20303);
and UO_1251 (O_1251,N_19475,N_24545);
nand UO_1252 (O_1252,N_24097,N_23088);
nor UO_1253 (O_1253,N_22879,N_19555);
nand UO_1254 (O_1254,N_24546,N_22504);
nor UO_1255 (O_1255,N_19998,N_21914);
nand UO_1256 (O_1256,N_20609,N_20017);
nand UO_1257 (O_1257,N_23962,N_23682);
or UO_1258 (O_1258,N_22316,N_23147);
and UO_1259 (O_1259,N_21562,N_21924);
or UO_1260 (O_1260,N_18986,N_18791);
and UO_1261 (O_1261,N_24708,N_20778);
nor UO_1262 (O_1262,N_23104,N_20945);
and UO_1263 (O_1263,N_22913,N_19077);
or UO_1264 (O_1264,N_22441,N_21811);
nor UO_1265 (O_1265,N_24362,N_22667);
nand UO_1266 (O_1266,N_21265,N_21393);
and UO_1267 (O_1267,N_21796,N_21835);
and UO_1268 (O_1268,N_19774,N_18922);
and UO_1269 (O_1269,N_22640,N_23735);
and UO_1270 (O_1270,N_19660,N_23505);
nor UO_1271 (O_1271,N_19943,N_24275);
or UO_1272 (O_1272,N_21047,N_22566);
xnor UO_1273 (O_1273,N_19597,N_24591);
or UO_1274 (O_1274,N_21744,N_22497);
or UO_1275 (O_1275,N_21144,N_21412);
nor UO_1276 (O_1276,N_24723,N_19144);
and UO_1277 (O_1277,N_23669,N_19487);
nand UO_1278 (O_1278,N_23843,N_21274);
or UO_1279 (O_1279,N_20466,N_20540);
and UO_1280 (O_1280,N_21451,N_24877);
nand UO_1281 (O_1281,N_23028,N_24151);
nor UO_1282 (O_1282,N_18817,N_24759);
or UO_1283 (O_1283,N_23233,N_21945);
or UO_1284 (O_1284,N_24959,N_22478);
and UO_1285 (O_1285,N_20764,N_24582);
nor UO_1286 (O_1286,N_23545,N_18814);
nor UO_1287 (O_1287,N_21722,N_24048);
nor UO_1288 (O_1288,N_20517,N_24949);
or UO_1289 (O_1289,N_19834,N_23407);
nor UO_1290 (O_1290,N_19213,N_21095);
or UO_1291 (O_1291,N_19102,N_19236);
nand UO_1292 (O_1292,N_24593,N_20404);
and UO_1293 (O_1293,N_23908,N_19615);
or UO_1294 (O_1294,N_23123,N_23634);
nor UO_1295 (O_1295,N_24319,N_19269);
nor UO_1296 (O_1296,N_23249,N_21119);
nand UO_1297 (O_1297,N_23483,N_20953);
nor UO_1298 (O_1298,N_19545,N_22811);
and UO_1299 (O_1299,N_21174,N_19172);
or UO_1300 (O_1300,N_23183,N_20908);
nand UO_1301 (O_1301,N_19639,N_22429);
nand UO_1302 (O_1302,N_20896,N_21509);
and UO_1303 (O_1303,N_22194,N_19570);
or UO_1304 (O_1304,N_21630,N_18924);
and UO_1305 (O_1305,N_23329,N_19814);
nor UO_1306 (O_1306,N_24100,N_23712);
and UO_1307 (O_1307,N_22444,N_23132);
and UO_1308 (O_1308,N_21043,N_22466);
or UO_1309 (O_1309,N_24355,N_21446);
or UO_1310 (O_1310,N_24459,N_19544);
or UO_1311 (O_1311,N_22513,N_19343);
nand UO_1312 (O_1312,N_23433,N_20572);
nor UO_1313 (O_1313,N_22574,N_20701);
or UO_1314 (O_1314,N_19217,N_20689);
nor UO_1315 (O_1315,N_18851,N_19951);
nand UO_1316 (O_1316,N_22005,N_20262);
or UO_1317 (O_1317,N_24893,N_20881);
and UO_1318 (O_1318,N_22088,N_23932);
or UO_1319 (O_1319,N_19939,N_23378);
and UO_1320 (O_1320,N_24065,N_24533);
nand UO_1321 (O_1321,N_23375,N_22686);
nand UO_1322 (O_1322,N_21448,N_22671);
nand UO_1323 (O_1323,N_20600,N_20565);
nor UO_1324 (O_1324,N_21060,N_22015);
nand UO_1325 (O_1325,N_22581,N_24937);
nand UO_1326 (O_1326,N_19372,N_24234);
and UO_1327 (O_1327,N_24365,N_21171);
nor UO_1328 (O_1328,N_22570,N_24660);
and UO_1329 (O_1329,N_23189,N_23122);
nand UO_1330 (O_1330,N_20632,N_21996);
and UO_1331 (O_1331,N_24876,N_24094);
nand UO_1332 (O_1332,N_24147,N_21103);
nor UO_1333 (O_1333,N_23477,N_19323);
and UO_1334 (O_1334,N_19960,N_24202);
nor UO_1335 (O_1335,N_20141,N_22426);
and UO_1336 (O_1336,N_23224,N_20060);
or UO_1337 (O_1337,N_21571,N_22817);
and UO_1338 (O_1338,N_24429,N_19393);
or UO_1339 (O_1339,N_18874,N_22029);
and UO_1340 (O_1340,N_22411,N_22837);
nor UO_1341 (O_1341,N_19898,N_24698);
nand UO_1342 (O_1342,N_22458,N_24573);
nor UO_1343 (O_1343,N_23717,N_18949);
or UO_1344 (O_1344,N_23092,N_20616);
nor UO_1345 (O_1345,N_20924,N_22116);
or UO_1346 (O_1346,N_21313,N_22490);
xnor UO_1347 (O_1347,N_22190,N_19751);
or UO_1348 (O_1348,N_20757,N_21366);
or UO_1349 (O_1349,N_19252,N_22399);
and UO_1350 (O_1350,N_23774,N_23613);
nand UO_1351 (O_1351,N_22047,N_18880);
nand UO_1352 (O_1352,N_20313,N_23434);
nor UO_1353 (O_1353,N_24101,N_23277);
or UO_1354 (O_1354,N_23470,N_19468);
nor UO_1355 (O_1355,N_22353,N_24074);
or UO_1356 (O_1356,N_24102,N_24015);
or UO_1357 (O_1357,N_24286,N_22722);
or UO_1358 (O_1358,N_20037,N_18910);
or UO_1359 (O_1359,N_24166,N_24726);
or UO_1360 (O_1360,N_19230,N_24505);
nor UO_1361 (O_1361,N_20429,N_22760);
nand UO_1362 (O_1362,N_22460,N_23213);
and UO_1363 (O_1363,N_22192,N_21419);
or UO_1364 (O_1364,N_23192,N_20309);
and UO_1365 (O_1365,N_23947,N_21727);
nand UO_1366 (O_1366,N_20803,N_20875);
and UO_1367 (O_1367,N_23095,N_23362);
and UO_1368 (O_1368,N_24504,N_21981);
nand UO_1369 (O_1369,N_20149,N_22009);
nand UO_1370 (O_1370,N_19921,N_21115);
nand UO_1371 (O_1371,N_18947,N_18929);
nand UO_1372 (O_1372,N_23323,N_23596);
and UO_1373 (O_1373,N_22572,N_22120);
or UO_1374 (O_1374,N_21078,N_22996);
nor UO_1375 (O_1375,N_23195,N_19244);
or UO_1376 (O_1376,N_24734,N_23865);
nor UO_1377 (O_1377,N_22942,N_22416);
nand UO_1378 (O_1378,N_19031,N_21929);
nand UO_1379 (O_1379,N_21083,N_22234);
or UO_1380 (O_1380,N_20308,N_21644);
nand UO_1381 (O_1381,N_19304,N_23898);
and UO_1382 (O_1382,N_24261,N_19116);
or UO_1383 (O_1383,N_21992,N_20061);
xnor UO_1384 (O_1384,N_22688,N_22632);
or UO_1385 (O_1385,N_21531,N_23038);
nor UO_1386 (O_1386,N_23699,N_23318);
or UO_1387 (O_1387,N_19552,N_23566);
and UO_1388 (O_1388,N_24753,N_21927);
nor UO_1389 (O_1389,N_21882,N_21269);
nand UO_1390 (O_1390,N_22979,N_24447);
or UO_1391 (O_1391,N_24045,N_22849);
or UO_1392 (O_1392,N_21614,N_22810);
nand UO_1393 (O_1393,N_20364,N_24804);
and UO_1394 (O_1394,N_21787,N_23644);
nand UO_1395 (O_1395,N_22586,N_20212);
nand UO_1396 (O_1396,N_20074,N_19757);
nand UO_1397 (O_1397,N_24438,N_19929);
nor UO_1398 (O_1398,N_19190,N_20316);
and UO_1399 (O_1399,N_20395,N_19320);
nand UO_1400 (O_1400,N_19712,N_23646);
and UO_1401 (O_1401,N_20162,N_22014);
or UO_1402 (O_1402,N_21850,N_19173);
or UO_1403 (O_1403,N_21046,N_22963);
and UO_1404 (O_1404,N_20202,N_22537);
nand UO_1405 (O_1405,N_21467,N_20805);
nand UO_1406 (O_1406,N_20628,N_21221);
and UO_1407 (O_1407,N_21286,N_19777);
nor UO_1408 (O_1408,N_23652,N_21640);
or UO_1409 (O_1409,N_24578,N_20363);
or UO_1410 (O_1410,N_20772,N_19961);
nand UO_1411 (O_1411,N_22480,N_23957);
and UO_1412 (O_1412,N_18945,N_23819);
and UO_1413 (O_1413,N_23278,N_18902);
or UO_1414 (O_1414,N_19271,N_20139);
nor UO_1415 (O_1415,N_24484,N_23448);
or UO_1416 (O_1416,N_19867,N_24711);
or UO_1417 (O_1417,N_20344,N_21211);
and UO_1418 (O_1418,N_19824,N_22663);
nand UO_1419 (O_1419,N_20301,N_22093);
and UO_1420 (O_1420,N_19807,N_19500);
nor UO_1421 (O_1421,N_23343,N_22406);
and UO_1422 (O_1422,N_22121,N_20006);
or UO_1423 (O_1423,N_24560,N_24590);
or UO_1424 (O_1424,N_22060,N_20904);
or UO_1425 (O_1425,N_22346,N_19299);
or UO_1426 (O_1426,N_21218,N_19584);
nor UO_1427 (O_1427,N_19349,N_21706);
and UO_1428 (O_1428,N_19608,N_23296);
nor UO_1429 (O_1429,N_23758,N_23340);
or UO_1430 (O_1430,N_19912,N_23281);
nor UO_1431 (O_1431,N_24377,N_21798);
and UO_1432 (O_1432,N_23863,N_24412);
nor UO_1433 (O_1433,N_23177,N_23239);
nand UO_1434 (O_1434,N_22653,N_24252);
and UO_1435 (O_1435,N_20769,N_22629);
and UO_1436 (O_1436,N_24786,N_24671);
or UO_1437 (O_1437,N_20476,N_20588);
nand UO_1438 (O_1438,N_20255,N_23564);
and UO_1439 (O_1439,N_23997,N_23012);
nand UO_1440 (O_1440,N_18862,N_23370);
nand UO_1441 (O_1441,N_24160,N_22463);
and UO_1442 (O_1442,N_19035,N_21324);
and UO_1443 (O_1443,N_24839,N_23462);
nand UO_1444 (O_1444,N_22403,N_22312);
nand UO_1445 (O_1445,N_20921,N_21106);
or UO_1446 (O_1446,N_19200,N_20532);
and UO_1447 (O_1447,N_23529,N_20209);
nand UO_1448 (O_1448,N_22418,N_24075);
or UO_1449 (O_1449,N_20494,N_23112);
or UO_1450 (O_1450,N_21158,N_24233);
nand UO_1451 (O_1451,N_23148,N_22986);
and UO_1452 (O_1452,N_24692,N_18777);
and UO_1453 (O_1453,N_24064,N_23073);
nand UO_1454 (O_1454,N_20150,N_22915);
or UO_1455 (O_1455,N_23415,N_19779);
or UO_1456 (O_1456,N_21459,N_19743);
nor UO_1457 (O_1457,N_22154,N_21005);
nor UO_1458 (O_1458,N_20652,N_24382);
nand UO_1459 (O_1459,N_19852,N_24494);
nor UO_1460 (O_1460,N_19331,N_24254);
and UO_1461 (O_1461,N_20104,N_20203);
and UO_1462 (O_1462,N_21016,N_23009);
nor UO_1463 (O_1463,N_19233,N_24340);
or UO_1464 (O_1464,N_21907,N_23907);
nand UO_1465 (O_1465,N_23037,N_18758);
nor UO_1466 (O_1466,N_22803,N_21474);
nor UO_1467 (O_1467,N_22703,N_19064);
and UO_1468 (O_1468,N_19722,N_19328);
or UO_1469 (O_1469,N_22726,N_22902);
and UO_1470 (O_1470,N_21003,N_22438);
nand UO_1471 (O_1471,N_20566,N_24601);
or UO_1472 (O_1472,N_24658,N_22476);
nand UO_1473 (O_1473,N_24191,N_23544);
nor UO_1474 (O_1474,N_20412,N_24073);
nand UO_1475 (O_1475,N_19461,N_20850);
nand UO_1476 (O_1476,N_24761,N_19170);
nand UO_1477 (O_1477,N_24003,N_23953);
or UO_1478 (O_1478,N_22987,N_24480);
or UO_1479 (O_1479,N_19900,N_19524);
and UO_1480 (O_1480,N_21928,N_21287);
or UO_1481 (O_1481,N_18873,N_22943);
or UO_1482 (O_1482,N_19670,N_21875);
or UO_1483 (O_1483,N_22828,N_23267);
nor UO_1484 (O_1484,N_21966,N_19534);
or UO_1485 (O_1485,N_18823,N_23716);
nor UO_1486 (O_1486,N_22339,N_21548);
nand UO_1487 (O_1487,N_22883,N_19330);
nand UO_1488 (O_1488,N_22417,N_21300);
nor UO_1489 (O_1489,N_21843,N_24329);
or UO_1490 (O_1490,N_21750,N_20783);
and UO_1491 (O_1491,N_18920,N_22103);
and UO_1492 (O_1492,N_23002,N_20977);
or UO_1493 (O_1493,N_24240,N_21797);
nor UO_1494 (O_1494,N_18792,N_23353);
nor UO_1495 (O_1495,N_23149,N_21612);
nor UO_1496 (O_1496,N_22011,N_21214);
nor UO_1497 (O_1497,N_24150,N_21120);
or UO_1498 (O_1498,N_24222,N_21565);
nor UO_1499 (O_1499,N_19911,N_21070);
xnor UO_1500 (O_1500,N_23787,N_23936);
nand UO_1501 (O_1501,N_22308,N_19355);
or UO_1502 (O_1502,N_23984,N_21495);
or UO_1503 (O_1503,N_20821,N_23647);
and UO_1504 (O_1504,N_24789,N_19533);
nand UO_1505 (O_1505,N_18967,N_20625);
and UO_1506 (O_1506,N_24395,N_22542);
or UO_1507 (O_1507,N_24701,N_22507);
nor UO_1508 (O_1508,N_19321,N_22751);
nor UO_1509 (O_1509,N_20265,N_20186);
nand UO_1510 (O_1510,N_21880,N_22051);
and UO_1511 (O_1511,N_24947,N_20091);
nand UO_1512 (O_1512,N_19622,N_21392);
nor UO_1513 (O_1513,N_24446,N_19938);
or UO_1514 (O_1514,N_24404,N_20798);
and UO_1515 (O_1515,N_24424,N_20672);
nand UO_1516 (O_1516,N_24360,N_21619);
nor UO_1517 (O_1517,N_22388,N_21355);
nand UO_1518 (O_1518,N_23950,N_24638);
xnor UO_1519 (O_1519,N_21592,N_23958);
nand UO_1520 (O_1520,N_19000,N_20430);
xnor UO_1521 (O_1521,N_23713,N_18886);
nand UO_1522 (O_1522,N_20528,N_19909);
or UO_1523 (O_1523,N_19842,N_21349);
nor UO_1524 (O_1524,N_24466,N_21657);
and UO_1525 (O_1525,N_22099,N_20646);
nor UO_1526 (O_1526,N_18838,N_21224);
nand UO_1527 (O_1527,N_18946,N_21237);
nand UO_1528 (O_1528,N_20827,N_21598);
and UO_1529 (O_1529,N_23798,N_20258);
and UO_1530 (O_1530,N_20611,N_23846);
and UO_1531 (O_1531,N_21421,N_20515);
nor UO_1532 (O_1532,N_24861,N_20695);
or UO_1533 (O_1533,N_23325,N_19630);
nor UO_1534 (O_1534,N_18903,N_24115);
nand UO_1535 (O_1535,N_23528,N_20876);
nor UO_1536 (O_1536,N_24334,N_20182);
xor UO_1537 (O_1537,N_23511,N_19803);
or UO_1538 (O_1538,N_24626,N_20874);
or UO_1539 (O_1539,N_24550,N_24089);
nand UO_1540 (O_1540,N_24274,N_21628);
and UO_1541 (O_1541,N_21985,N_23450);
nand UO_1542 (O_1542,N_22540,N_20296);
and UO_1543 (O_1543,N_18870,N_20571);
and UO_1544 (O_1544,N_21134,N_21242);
nand UO_1545 (O_1545,N_23702,N_23779);
and UO_1546 (O_1546,N_19669,N_22086);
or UO_1547 (O_1547,N_22700,N_24913);
nand UO_1548 (O_1548,N_21793,N_24350);
or UO_1549 (O_1549,N_18982,N_23662);
or UO_1550 (O_1550,N_19138,N_18850);
nand UO_1551 (O_1551,N_20028,N_22236);
nand UO_1552 (O_1552,N_19963,N_20709);
and UO_1553 (O_1553,N_21938,N_18987);
and UO_1554 (O_1554,N_23518,N_22425);
or UO_1555 (O_1555,N_22641,N_19158);
and UO_1556 (O_1556,N_19704,N_20048);
or UO_1557 (O_1557,N_22106,N_24902);
nand UO_1558 (O_1558,N_22966,N_22197);
nor UO_1559 (O_1559,N_20740,N_24829);
nor UO_1560 (O_1560,N_21694,N_22187);
and UO_1561 (O_1561,N_19997,N_24371);
nor UO_1562 (O_1562,N_22334,N_20519);
or UO_1563 (O_1563,N_19863,N_23382);
nor UO_1564 (O_1564,N_24320,N_19050);
or UO_1565 (O_1565,N_23167,N_20417);
and UO_1566 (O_1566,N_20640,N_24928);
and UO_1567 (O_1567,N_20993,N_22493);
and UO_1568 (O_1568,N_24277,N_21919);
or UO_1569 (O_1569,N_24358,N_21780);
nor UO_1570 (O_1570,N_22922,N_23752);
nand UO_1571 (O_1571,N_19730,N_18828);
or UO_1572 (O_1572,N_20724,N_21713);
nand UO_1573 (O_1573,N_23840,N_19403);
nand UO_1574 (O_1574,N_21262,N_21346);
and UO_1575 (O_1575,N_23482,N_21476);
nand UO_1576 (O_1576,N_21517,N_22273);
or UO_1577 (O_1577,N_23436,N_20131);
and UO_1578 (O_1578,N_19937,N_24189);
and UO_1579 (O_1579,N_22954,N_23579);
nor UO_1580 (O_1580,N_23497,N_24030);
and UO_1581 (O_1581,N_22369,N_24962);
nand UO_1582 (O_1582,N_22384,N_19672);
or UO_1583 (O_1583,N_22684,N_24243);
or UO_1584 (O_1584,N_21414,N_23695);
nor UO_1585 (O_1585,N_22764,N_21730);
or UO_1586 (O_1586,N_22889,N_21368);
and UO_1587 (O_1587,N_20077,N_19994);
or UO_1588 (O_1588,N_24373,N_21623);
nor UO_1589 (O_1589,N_19715,N_24031);
nor UO_1590 (O_1590,N_20879,N_24524);
and UO_1591 (O_1591,N_21867,N_20575);
nor UO_1592 (O_1592,N_20274,N_21800);
nand UO_1593 (O_1593,N_20020,N_23398);
nand UO_1594 (O_1594,N_22118,N_18958);
nand UO_1595 (O_1595,N_21799,N_24047);
and UO_1596 (O_1596,N_20453,N_20337);
or UO_1597 (O_1597,N_18890,N_21748);
nand UO_1598 (O_1598,N_23922,N_19601);
nor UO_1599 (O_1599,N_22898,N_23219);
and UO_1600 (O_1600,N_23013,N_23929);
nor UO_1601 (O_1601,N_24495,N_24536);
or UO_1602 (O_1602,N_19861,N_24836);
or UO_1603 (O_1603,N_20754,N_24954);
or UO_1604 (O_1604,N_22271,N_21100);
nor UO_1605 (O_1605,N_24969,N_23358);
nor UO_1606 (O_1606,N_21549,N_19098);
nor UO_1607 (O_1607,N_22161,N_24337);
nor UO_1608 (O_1608,N_19562,N_20635);
nand UO_1609 (O_1609,N_20730,N_24305);
nand UO_1610 (O_1610,N_23124,N_20710);
nand UO_1611 (O_1611,N_23591,N_24069);
or UO_1612 (O_1612,N_20750,N_21460);
and UO_1613 (O_1613,N_21801,N_19180);
and UO_1614 (O_1614,N_24544,N_24154);
or UO_1615 (O_1615,N_24646,N_22896);
nand UO_1616 (O_1616,N_22946,N_20914);
nand UO_1617 (O_1617,N_19182,N_24140);
and UO_1618 (O_1618,N_19529,N_19268);
or UO_1619 (O_1619,N_22081,N_22124);
and UO_1620 (O_1620,N_20813,N_21112);
nor UO_1621 (O_1621,N_23806,N_21455);
or UO_1622 (O_1622,N_22571,N_22731);
or UO_1623 (O_1623,N_23949,N_23459);
or UO_1624 (O_1624,N_24532,N_24418);
or UO_1625 (O_1625,N_20307,N_23981);
and UO_1626 (O_1626,N_20567,N_20013);
nor UO_1627 (O_1627,N_20770,N_21873);
or UO_1628 (O_1628,N_24199,N_20555);
nor UO_1629 (O_1629,N_19981,N_24407);
or UO_1630 (O_1630,N_21848,N_19010);
nor UO_1631 (O_1631,N_21257,N_21057);
nor UO_1632 (O_1632,N_21449,N_23396);
and UO_1633 (O_1633,N_22693,N_20774);
nand UO_1634 (O_1634,N_20047,N_21983);
and UO_1635 (O_1635,N_23814,N_20553);
nand UO_1636 (O_1636,N_19992,N_18764);
or UO_1637 (O_1637,N_18832,N_20067);
nor UO_1638 (O_1638,N_21390,N_21167);
nor UO_1639 (O_1639,N_22601,N_21946);
nor UO_1640 (O_1640,N_18896,N_20509);
nor UO_1641 (O_1641,N_19589,N_21009);
nand UO_1642 (O_1642,N_19968,N_19571);
nor UO_1643 (O_1643,N_23951,N_24768);
or UO_1644 (O_1644,N_23598,N_20343);
nor UO_1645 (O_1645,N_24832,N_18953);
and UO_1646 (O_1646,N_23696,N_21243);
nand UO_1647 (O_1647,N_21075,N_24475);
or UO_1648 (O_1648,N_20651,N_22113);
nor UO_1649 (O_1649,N_20062,N_22007);
or UO_1650 (O_1650,N_22095,N_23082);
nand UO_1651 (O_1651,N_22689,N_19195);
and UO_1652 (O_1652,N_19253,N_23313);
or UO_1653 (O_1653,N_23280,N_21513);
and UO_1654 (O_1654,N_23822,N_19927);
nand UO_1655 (O_1655,N_19588,N_19352);
or UO_1656 (O_1656,N_19086,N_20814);
nor UO_1657 (O_1657,N_22183,N_21477);
nand UO_1658 (O_1658,N_23801,N_19879);
nor UO_1659 (O_1659,N_18933,N_18937);
and UO_1660 (O_1660,N_24415,N_21154);
or UO_1661 (O_1661,N_21641,N_19082);
or UO_1662 (O_1662,N_24270,N_24114);
and UO_1663 (O_1663,N_19404,N_18885);
and UO_1664 (O_1664,N_24700,N_19758);
nor UO_1665 (O_1665,N_22173,N_19001);
nand UO_1666 (O_1666,N_19948,N_19869);
and UO_1667 (O_1667,N_23820,N_21383);
or UO_1668 (O_1668,N_21153,N_20055);
nand UO_1669 (O_1669,N_19744,N_21137);
and UO_1670 (O_1670,N_20004,N_23101);
or UO_1671 (O_1671,N_20971,N_21213);
xnor UO_1672 (O_1672,N_24921,N_21178);
or UO_1673 (O_1673,N_21855,N_22949);
and UO_1674 (O_1674,N_22792,N_18845);
nand UO_1675 (O_1675,N_24648,N_24691);
and UO_1676 (O_1676,N_19825,N_21779);
and UO_1677 (O_1677,N_20982,N_22319);
nand UO_1678 (O_1678,N_20125,N_20163);
or UO_1679 (O_1679,N_19479,N_21109);
or UO_1680 (O_1680,N_20922,N_20312);
or UO_1681 (O_1681,N_21172,N_22706);
nor UO_1682 (O_1682,N_23247,N_22010);
or UO_1683 (O_1683,N_18926,N_23824);
and UO_1684 (O_1684,N_21293,N_22185);
or UO_1685 (O_1685,N_23834,N_22887);
nand UO_1686 (O_1686,N_19539,N_21617);
nor UO_1687 (O_1687,N_22761,N_18829);
nand UO_1688 (O_1688,N_24125,N_22056);
and UO_1689 (O_1689,N_21423,N_19498);
nor UO_1690 (O_1690,N_19614,N_21018);
nand UO_1691 (O_1691,N_21024,N_20034);
and UO_1692 (O_1692,N_23156,N_23310);
and UO_1693 (O_1693,N_19378,N_19148);
xor UO_1694 (O_1694,N_19808,N_20188);
and UO_1695 (O_1695,N_23125,N_19373);
or UO_1696 (O_1696,N_21182,N_21091);
and UO_1697 (O_1697,N_22651,N_19022);
nand UO_1698 (O_1698,N_22064,N_20270);
nor UO_1699 (O_1699,N_24707,N_23298);
and UO_1700 (O_1700,N_23166,N_20843);
nor UO_1701 (O_1701,N_20642,N_23534);
xor UO_1702 (O_1702,N_21055,N_23050);
nand UO_1703 (O_1703,N_23316,N_20490);
nor UO_1704 (O_1704,N_22021,N_19871);
nand UO_1705 (O_1705,N_22853,N_24464);
or UO_1706 (O_1706,N_22790,N_22533);
nand UO_1707 (O_1707,N_18778,N_19646);
and UO_1708 (O_1708,N_19206,N_19716);
nand UO_1709 (O_1709,N_20694,N_21282);
or UO_1710 (O_1710,N_24952,N_21504);
nor UO_1711 (O_1711,N_20577,N_21977);
or UO_1712 (O_1712,N_22479,N_22619);
nand UO_1713 (O_1713,N_21309,N_22960);
nand UO_1714 (O_1714,N_24058,N_23240);
or UO_1715 (O_1715,N_20427,N_24709);
or UO_1716 (O_1716,N_22869,N_20192);
and UO_1717 (O_1717,N_22560,N_23805);
or UO_1718 (O_1718,N_20082,N_19641);
or UO_1719 (O_1719,N_22538,N_24085);
nor UO_1720 (O_1720,N_21759,N_19100);
nand UO_1721 (O_1721,N_18969,N_24957);
xor UO_1722 (O_1722,N_20570,N_24666);
nand UO_1723 (O_1723,N_24515,N_24173);
and UO_1724 (O_1724,N_22274,N_19820);
nand UO_1725 (O_1725,N_20390,N_19788);
nand UO_1726 (O_1726,N_19259,N_23420);
nand UO_1727 (O_1727,N_20056,N_20806);
nor UO_1728 (O_1728,N_20052,N_22165);
or UO_1729 (O_1729,N_22314,N_21408);
and UO_1730 (O_1730,N_24682,N_24635);
and UO_1731 (O_1731,N_19248,N_23120);
nand UO_1732 (O_1732,N_20816,N_19607);
or UO_1733 (O_1733,N_24257,N_19700);
or UO_1734 (O_1734,N_19122,N_24321);
nand UO_1735 (O_1735,N_21891,N_24643);
and UO_1736 (O_1736,N_22250,N_23959);
or UO_1737 (O_1737,N_22123,N_24737);
nand UO_1738 (O_1738,N_19020,N_20240);
nand UO_1739 (O_1739,N_23838,N_24391);
nor UO_1740 (O_1740,N_20516,N_24814);
nand UO_1741 (O_1741,N_22457,N_23719);
nor UO_1742 (O_1742,N_22529,N_19193);
or UO_1743 (O_1743,N_22594,N_22202);
nand UO_1744 (O_1744,N_20450,N_20845);
nand UO_1745 (O_1745,N_21002,N_23109);
nor UO_1746 (O_1746,N_23617,N_19590);
nand UO_1747 (O_1747,N_20254,N_23388);
nand UO_1748 (O_1748,N_24180,N_24853);
and UO_1749 (O_1749,N_23320,N_20911);
nor UO_1750 (O_1750,N_24139,N_20251);
or UO_1751 (O_1751,N_21580,N_23419);
nand UO_1752 (O_1752,N_18981,N_24168);
nand UO_1753 (O_1753,N_20347,N_21191);
and UO_1754 (O_1754,N_21784,N_21227);
and UO_1755 (O_1755,N_23349,N_21535);
nand UO_1756 (O_1756,N_21193,N_21665);
nor UO_1757 (O_1757,N_23290,N_18859);
nand UO_1758 (O_1758,N_19637,N_19453);
or UO_1759 (O_1759,N_19450,N_20889);
nand UO_1760 (O_1760,N_19643,N_24072);
nor UO_1761 (O_1761,N_23746,N_21910);
or UO_1762 (O_1762,N_22848,N_24776);
nand UO_1763 (O_1763,N_19290,N_22714);
or UO_1764 (O_1764,N_22672,N_21074);
nand UO_1765 (O_1765,N_23615,N_21761);
nor UO_1766 (O_1766,N_22000,N_24738);
and UO_1767 (O_1767,N_23099,N_19664);
or UO_1768 (O_1768,N_19499,N_23100);
nand UO_1769 (O_1769,N_19016,N_22825);
or UO_1770 (O_1770,N_21508,N_20594);
nor UO_1771 (O_1771,N_23681,N_22829);
and UO_1772 (O_1772,N_19289,N_23625);
nor UO_1773 (O_1773,N_19819,N_19506);
or UO_1774 (O_1774,N_20167,N_24439);
nor UO_1775 (O_1775,N_23558,N_23621);
xnor UO_1776 (O_1776,N_19605,N_19084);
or UO_1777 (O_1777,N_19931,N_21920);
or UO_1778 (O_1778,N_23004,N_23029);
nor UO_1779 (O_1779,N_23995,N_19813);
nand UO_1780 (O_1780,N_24375,N_19246);
nor UO_1781 (O_1781,N_19800,N_20781);
nand UO_1782 (O_1782,N_23085,N_21208);
nand UO_1783 (O_1783,N_24297,N_24722);
nand UO_1784 (O_1784,N_18905,N_20592);
or UO_1785 (O_1785,N_23282,N_22097);
nand UO_1786 (O_1786,N_21723,N_24068);
nand UO_1787 (O_1787,N_19046,N_22446);
nor UO_1788 (O_1788,N_24018,N_20584);
nand UO_1789 (O_1789,N_22372,N_19679);
or UO_1790 (O_1790,N_22622,N_22296);
nand UO_1791 (O_1791,N_23729,N_24280);
nor UO_1792 (O_1792,N_20375,N_23887);
or UO_1793 (O_1793,N_20521,N_22258);
and UO_1794 (O_1794,N_21973,N_22577);
nand UO_1795 (O_1795,N_19411,N_24994);
nand UO_1796 (O_1796,N_19160,N_19201);
nand UO_1797 (O_1797,N_24136,N_24639);
nor UO_1798 (O_1798,N_23289,N_22484);
or UO_1799 (O_1799,N_19178,N_24561);
nor UO_1800 (O_1800,N_23299,N_18812);
and UO_1801 (O_1801,N_22341,N_23512);
nor UO_1802 (O_1802,N_19363,N_22523);
nor UO_1803 (O_1803,N_18811,N_19225);
nor UO_1804 (O_1804,N_20368,N_20421);
and UO_1805 (O_1805,N_22891,N_24176);
and UO_1806 (O_1806,N_21905,N_21296);
nand UO_1807 (O_1807,N_23453,N_24175);
and UO_1808 (O_1808,N_20297,N_24860);
nand UO_1809 (O_1809,N_21610,N_24813);
nand UO_1810 (O_1810,N_19903,N_22682);
nand UO_1811 (O_1811,N_24664,N_23837);
nor UO_1812 (O_1812,N_22083,N_19202);
or UO_1813 (O_1813,N_23631,N_22344);
and UO_1814 (O_1814,N_20106,N_22749);
nand UO_1815 (O_1815,N_22133,N_23599);
nand UO_1816 (O_1816,N_24409,N_20259);
nor UO_1817 (O_1817,N_19551,N_22907);
nand UO_1818 (O_1818,N_22906,N_21266);
nand UO_1819 (O_1819,N_21756,N_20492);
nor UO_1820 (O_1820,N_20178,N_22839);
nand UO_1821 (O_1821,N_19344,N_20529);
or UO_1822 (O_1822,N_18776,N_19400);
nor UO_1823 (O_1823,N_19197,N_20140);
nand UO_1824 (O_1824,N_21558,N_22857);
and UO_1825 (O_1825,N_19063,N_20030);
nand UO_1826 (O_1826,N_23217,N_22421);
nand UO_1827 (O_1827,N_22620,N_22863);
or UO_1828 (O_1828,N_19085,N_19857);
nand UO_1829 (O_1829,N_21745,N_20582);
nand UO_1830 (O_1830,N_24263,N_22994);
and UO_1831 (O_1831,N_23987,N_24568);
or UO_1832 (O_1832,N_19926,N_23061);
and UO_1833 (O_1833,N_20029,N_21877);
and UO_1834 (O_1834,N_21212,N_22740);
nand UO_1835 (O_1835,N_21444,N_24313);
nor UO_1836 (O_1836,N_22984,N_19387);
nand UO_1837 (O_1837,N_20527,N_23231);
nand UO_1838 (O_1838,N_20715,N_21714);
nand UO_1839 (O_1839,N_23304,N_24026);
nand UO_1840 (O_1840,N_23431,N_19798);
or UO_1841 (O_1841,N_21044,N_19208);
nand UO_1842 (O_1842,N_22823,N_23417);
nand UO_1843 (O_1843,N_19642,N_24311);
and UO_1844 (O_1844,N_20330,N_23541);
nor UO_1845 (O_1845,N_19218,N_23322);
nor UO_1846 (O_1846,N_22501,N_24818);
and UO_1847 (O_1847,N_21290,N_19334);
nor UO_1848 (O_1848,N_23679,N_20331);
and UO_1849 (O_1849,N_23261,N_24408);
nor UO_1850 (O_1850,N_22592,N_24308);
and UO_1851 (O_1851,N_22326,N_23731);
and UO_1852 (O_1852,N_19040,N_23581);
nor UO_1853 (O_1853,N_20920,N_18804);
and UO_1854 (O_1854,N_21307,N_24008);
or UO_1855 (O_1855,N_22380,N_21520);
nor UO_1856 (O_1856,N_20377,N_22333);
and UO_1857 (O_1857,N_20824,N_24610);
nand UO_1858 (O_1858,N_23533,N_24535);
or UO_1859 (O_1859,N_23202,N_21809);
nand UO_1860 (O_1860,N_24678,N_24405);
nand UO_1861 (O_1861,N_20485,N_22695);
and UO_1862 (O_1862,N_24750,N_21586);
nand UO_1863 (O_1863,N_24798,N_19799);
nand UO_1864 (O_1864,N_23054,N_21022);
nand UO_1865 (O_1865,N_23791,N_19793);
or UO_1866 (O_1866,N_21344,N_21879);
and UO_1867 (O_1867,N_22772,N_23660);
or UO_1868 (O_1868,N_20681,N_20228);
and UO_1869 (O_1869,N_20573,N_19367);
and UO_1870 (O_1870,N_20548,N_19358);
nor UO_1871 (O_1871,N_21111,N_21906);
nor UO_1872 (O_1872,N_20985,N_19940);
or UO_1873 (O_1873,N_20021,N_23873);
nand UO_1874 (O_1874,N_20556,N_19006);
or UO_1875 (O_1875,N_21908,N_22117);
nand UO_1876 (O_1876,N_18780,N_20271);
and UO_1877 (O_1877,N_23180,N_24379);
or UO_1878 (O_1878,N_19247,N_22130);
nand UO_1879 (O_1879,N_24171,N_24982);
and UO_1880 (O_1880,N_22195,N_21705);
and UO_1881 (O_1881,N_20550,N_23191);
and UO_1882 (O_1882,N_19520,N_24702);
or UO_1883 (O_1883,N_24594,N_18883);
and UO_1884 (O_1884,N_24393,N_19033);
or UO_1885 (O_1885,N_20211,N_19394);
nor UO_1886 (O_1886,N_23977,N_18891);
and UO_1887 (O_1887,N_21029,N_21301);
nor UO_1888 (O_1888,N_19003,N_20185);
or UO_1889 (O_1889,N_22057,N_24825);
and UO_1890 (O_1890,N_20318,N_23797);
nand UO_1891 (O_1891,N_20916,N_19301);
nor UO_1892 (O_1892,N_24778,N_21584);
nor UO_1893 (O_1893,N_20408,N_18983);
nor UO_1894 (O_1894,N_20970,N_22208);
nor UO_1895 (O_1895,N_20317,N_23942);
nand UO_1896 (O_1896,N_20595,N_24914);
and UO_1897 (O_1897,N_24999,N_20475);
nor UO_1898 (O_1898,N_20423,N_22831);
or UO_1899 (O_1899,N_18787,N_20069);
or UO_1900 (O_1900,N_19654,N_23031);
nor UO_1901 (O_1901,N_23250,N_21975);
and UO_1902 (O_1902,N_21255,N_23618);
nor UO_1903 (O_1903,N_21371,N_21898);
or UO_1904 (O_1904,N_20103,N_19745);
and UO_1905 (O_1905,N_23546,N_22957);
nand UO_1906 (O_1906,N_20465,N_24359);
nand UO_1907 (O_1907,N_22806,N_24688);
and UO_1908 (O_1908,N_22415,N_23877);
xor UO_1909 (O_1909,N_23111,N_22539);
or UO_1910 (O_1910,N_20002,N_24473);
and UO_1911 (O_1911,N_21698,N_19384);
nor UO_1912 (O_1912,N_24728,N_22990);
nor UO_1913 (O_1913,N_20235,N_20224);
nand UO_1914 (O_1914,N_21604,N_20664);
and UO_1915 (O_1915,N_22704,N_23749);
or UO_1916 (O_1916,N_20643,N_24098);
and UO_1917 (O_1917,N_22068,N_23800);
nor UO_1918 (O_1918,N_23196,N_23554);
nand UO_1919 (O_1919,N_19702,N_21700);
nand UO_1920 (O_1920,N_20790,N_22997);
nor UO_1921 (O_1921,N_20370,N_23270);
and UO_1922 (O_1922,N_21056,N_24556);
and UO_1923 (O_1923,N_20154,N_24703);
and UO_1924 (O_1924,N_23175,N_21685);
and UO_1925 (O_1925,N_19831,N_19671);
nor UO_1926 (O_1926,N_21483,N_20191);
or UO_1927 (O_1927,N_23452,N_22323);
or UO_1928 (O_1928,N_23410,N_20861);
and UO_1929 (O_1929,N_22736,N_21788);
nor UO_1930 (O_1930,N_23727,N_21599);
and UO_1931 (O_1931,N_23481,N_21736);
nor UO_1932 (O_1932,N_22336,N_19868);
nor UO_1933 (O_1933,N_24522,N_20038);
and UO_1934 (O_1934,N_19781,N_24055);
nand UO_1935 (O_1935,N_22332,N_20885);
nand UO_1936 (O_1936,N_20230,N_24905);
and UO_1937 (O_1937,N_21042,N_22668);
or UO_1938 (O_1938,N_19205,N_23839);
and UO_1939 (O_1939,N_24971,N_19662);
and UO_1940 (O_1940,N_24963,N_23008);
nor UO_1941 (O_1941,N_23939,N_24145);
and UO_1942 (O_1942,N_22335,N_22108);
nor UO_1943 (O_1943,N_22355,N_24284);
nor UO_1944 (O_1944,N_23620,N_21322);
or UO_1945 (O_1945,N_20551,N_21152);
or UO_1946 (O_1946,N_23520,N_23114);
and UO_1947 (O_1947,N_24856,N_19631);
and UO_1948 (O_1948,N_22186,N_20941);
nand UO_1949 (O_1949,N_22255,N_22330);
nor UO_1950 (O_1950,N_20345,N_24185);
or UO_1951 (O_1951,N_21405,N_23861);
or UO_1952 (O_1952,N_19188,N_24852);
nor UO_1953 (O_1953,N_20581,N_23019);
and UO_1954 (O_1954,N_21538,N_24183);
and UO_1955 (O_1955,N_23638,N_19153);
nand UO_1956 (O_1956,N_21632,N_22428);
or UO_1957 (O_1957,N_24067,N_24236);
nand UO_1958 (O_1958,N_19661,N_23882);
nor UO_1959 (O_1959,N_24616,N_22780);
and UO_1960 (O_1960,N_23406,N_18796);
nand UO_1961 (O_1961,N_22639,N_22004);
nor UO_1962 (O_1962,N_24454,N_20637);
nand UO_1963 (O_1963,N_24281,N_19288);
and UO_1964 (O_1964,N_20479,N_24663);
nor UO_1965 (O_1965,N_24501,N_22370);
xnor UO_1966 (O_1966,N_20367,N_21235);
nand UO_1967 (O_1967,N_23968,N_21123);
or UO_1968 (O_1968,N_23750,N_22631);
nand UO_1969 (O_1969,N_20040,N_23194);
and UO_1970 (O_1970,N_21778,N_22576);
nand UO_1971 (O_1971,N_21030,N_19987);
or UO_1972 (O_1972,N_19999,N_22288);
nand UO_1973 (O_1973,N_24748,N_22765);
nand UO_1974 (O_1974,N_20638,N_23426);
nor UO_1975 (O_1975,N_20546,N_24042);
and UO_1976 (O_1976,N_24598,N_24024);
or UO_1977 (O_1977,N_19112,N_21827);
or UO_1978 (O_1978,N_23658,N_19636);
nand UO_1979 (O_1979,N_23521,N_24361);
and UO_1980 (O_1980,N_22947,N_20261);
nor UO_1981 (O_1981,N_24077,N_22328);
and UO_1982 (O_1982,N_22340,N_22773);
or UO_1983 (O_1983,N_24966,N_23989);
nand UO_1984 (O_1984,N_19296,N_19954);
xnor UO_1985 (O_1985,N_24028,N_23292);
nor UO_1986 (O_1986,N_22352,N_24105);
nor UO_1987 (O_1987,N_24694,N_23780);
nor UO_1988 (O_1988,N_20537,N_23722);
nand UO_1989 (O_1989,N_19853,N_20379);
and UO_1990 (O_1990,N_22903,N_23064);
nand UO_1991 (O_1991,N_24108,N_19346);
nand UO_1992 (O_1992,N_23608,N_24088);
and UO_1993 (O_1993,N_20606,N_24036);
or UO_1994 (O_1994,N_19189,N_19421);
xor UO_1995 (O_1995,N_19763,N_21689);
or UO_1996 (O_1996,N_24226,N_20812);
nor UO_1997 (O_1997,N_18809,N_24974);
and UO_1998 (O_1998,N_22813,N_24493);
and UO_1999 (O_1999,N_22759,N_23597);
or UO_2000 (O_2000,N_23766,N_22491);
and UO_2001 (O_2001,N_19440,N_19812);
nand UO_2002 (O_2002,N_20152,N_21890);
nor UO_2003 (O_2003,N_19260,N_22789);
xor UO_2004 (O_2004,N_18866,N_21229);
nor UO_2005 (O_2005,N_19942,N_20166);
nor UO_2006 (O_2006,N_20848,N_21289);
xnor UO_2007 (O_2007,N_23210,N_23408);
or UO_2008 (O_2008,N_19274,N_19756);
nand UO_2009 (O_2009,N_20266,N_24050);
nor UO_2010 (O_2010,N_22160,N_24980);
or UO_2011 (O_2011,N_20526,N_22036);
and UO_2012 (O_2012,N_19243,N_23405);
and UO_2013 (O_2013,N_23478,N_21672);
nand UO_2014 (O_2014,N_22241,N_20867);
nand UO_2015 (O_2015,N_19366,N_22785);
or UO_2016 (O_2016,N_19692,N_19174);
and UO_2017 (O_2017,N_21020,N_23747);
nand UO_2018 (O_2018,N_22827,N_22101);
or UO_2019 (O_2019,N_22795,N_22285);
nor UO_2020 (O_2020,N_24736,N_18860);
and UO_2021 (O_2021,N_22470,N_21947);
nand UO_2022 (O_2022,N_22665,N_23971);
or UO_2023 (O_2023,N_22405,N_20353);
and UO_2024 (O_2024,N_19079,N_20887);
or UO_2025 (O_2025,N_20187,N_21710);
nand UO_2026 (O_2026,N_19119,N_20873);
and UO_2027 (O_2027,N_22935,N_21782);
nand UO_2028 (O_2028,N_24896,N_24620);
or UO_2029 (O_2029,N_24258,N_21225);
nor UO_2030 (O_2030,N_24044,N_20484);
nand UO_2031 (O_2031,N_19145,N_23985);
or UO_2032 (O_2032,N_24356,N_22741);
and UO_2033 (O_2033,N_24597,N_21533);
nor UO_2034 (O_2034,N_23633,N_19183);
and UO_2035 (O_2035,N_24878,N_22625);
or UO_2036 (O_2036,N_24943,N_24919);
nor UO_2037 (O_2037,N_20449,N_20372);
nor UO_2038 (O_2038,N_24733,N_21765);
or UO_2039 (O_2039,N_19736,N_19496);
or UO_2040 (O_2040,N_22830,N_21045);
and UO_2041 (O_2041,N_23934,N_21984);
nor UO_2042 (O_2042,N_23569,N_24566);
and UO_2043 (O_2043,N_19476,N_23141);
or UO_2044 (O_2044,N_22526,N_23334);
nand UO_2045 (O_2045,N_19711,N_21524);
nor UO_2046 (O_2046,N_18895,N_21747);
nor UO_2047 (O_2047,N_21126,N_20204);
or UO_2048 (O_2048,N_23869,N_18871);
nor UO_2049 (O_2049,N_21521,N_20456);
or UO_2050 (O_2050,N_20801,N_22678);
or UO_2051 (O_2051,N_20273,N_20678);
xnor UO_2052 (O_2052,N_21485,N_23870);
nor UO_2053 (O_2053,N_20533,N_22084);
nand UO_2054 (O_2054,N_24384,N_21114);
or UO_2055 (O_2055,N_24633,N_24231);
nor UO_2056 (O_2056,N_23016,N_22447);
or UO_2057 (O_2057,N_22392,N_20100);
nor UO_2058 (O_2058,N_23653,N_20831);
and UO_2059 (O_2059,N_21557,N_23072);
nor UO_2060 (O_2060,N_22721,N_23212);
or UO_2061 (O_2061,N_21395,N_22400);
nand UO_2062 (O_2062,N_20670,N_20325);
nor UO_2063 (O_2063,N_19656,N_20420);
or UO_2064 (O_2064,N_20524,N_21422);
nand UO_2065 (O_2065,N_21138,N_24423);
nor UO_2066 (O_2066,N_22939,N_22016);
and UO_2067 (O_2067,N_18825,N_19883);
or UO_2068 (O_2068,N_24756,N_24978);
nand UO_2069 (O_2069,N_21204,N_22649);
nor UO_2070 (O_2070,N_24514,N_19592);
and UO_2071 (O_2071,N_19765,N_18911);
nor UO_2072 (O_2072,N_23738,N_22278);
nor UO_2073 (O_2073,N_24223,N_19211);
nand UO_2074 (O_2074,N_20210,N_23153);
nor UO_2075 (O_2075,N_22348,N_19920);
and UO_2076 (O_2076,N_22750,N_20302);
or UO_2077 (O_2077,N_20244,N_19157);
or UO_2078 (O_2078,N_21852,N_21749);
nor UO_2079 (O_2079,N_22901,N_20622);
nand UO_2080 (O_2080,N_21142,N_24617);
nand UO_2081 (O_2081,N_21643,N_24109);
and UO_2082 (O_2082,N_18783,N_19256);
nor UO_2083 (O_2083,N_19752,N_20143);
nor UO_2084 (O_2084,N_23537,N_21202);
or UO_2085 (O_2085,N_22735,N_24153);
nand UO_2086 (O_2086,N_22933,N_22002);
nand UO_2087 (O_2087,N_21969,N_24080);
and UO_2088 (O_2088,N_18770,N_18781);
nand UO_2089 (O_2089,N_22778,N_24542);
nand UO_2090 (O_2090,N_24587,N_24197);
xnor UO_2091 (O_2091,N_20499,N_19414);
nor UO_2092 (O_2092,N_19759,N_19721);
nand UO_2093 (O_2093,N_19889,N_20648);
and UO_2094 (O_2094,N_22300,N_20121);
or UO_2095 (O_2095,N_23135,N_23501);
or UO_2096 (O_2096,N_24022,N_24670);
nand UO_2097 (O_2097,N_19129,N_24066);
or UO_2098 (O_2098,N_23003,N_23755);
nor UO_2099 (O_2099,N_21155,N_23455);
nand UO_2100 (O_2100,N_22481,N_19895);
nand UO_2101 (O_2101,N_19950,N_23244);
nand UO_2102 (O_2102,N_22127,N_22556);
nand UO_2103 (O_2103,N_22892,N_19993);
nor UO_2104 (O_2104,N_21447,N_22860);
nor UO_2105 (O_2105,N_19826,N_20064);
and UO_2106 (O_2106,N_23307,N_24020);
and UO_2107 (O_2107,N_20422,N_18789);
or UO_2108 (O_2108,N_22936,N_20223);
and UO_2109 (O_2109,N_22885,N_20508);
and UO_2110 (O_2110,N_24965,N_24392);
nand UO_2111 (O_2111,N_19456,N_23751);
and UO_2112 (O_2112,N_20855,N_23637);
nand UO_2113 (O_2113,N_20320,N_23366);
nand UO_2114 (O_2114,N_20641,N_19113);
nand UO_2115 (O_2115,N_20773,N_22557);
and UO_2116 (O_2116,N_22621,N_24595);
and UO_2117 (O_2117,N_21865,N_22292);
and UO_2118 (O_2118,N_24934,N_21317);
or UO_2119 (O_2119,N_21886,N_22515);
xor UO_2120 (O_2120,N_24900,N_24676);
nand UO_2121 (O_2121,N_19770,N_20994);
and UO_2122 (O_2122,N_19742,N_22786);
nand UO_2123 (O_2123,N_21165,N_23160);
and UO_2124 (O_2124,N_20117,N_24266);
or UO_2125 (O_2125,N_24822,N_20333);
and UO_2126 (O_2126,N_21357,N_20732);
or UO_2127 (O_2127,N_24265,N_20987);
nor UO_2128 (O_2128,N_22650,N_23223);
and UO_2129 (O_2129,N_23891,N_23489);
nand UO_2130 (O_2130,N_21133,N_22643);
nand UO_2131 (O_2131,N_22224,N_23956);
nor UO_2132 (O_2132,N_20562,N_20884);
or UO_2133 (O_2133,N_22908,N_24103);
and UO_2134 (O_2134,N_21740,N_18985);
and UO_2135 (O_2135,N_20535,N_20011);
nor UO_2136 (O_2136,N_24569,N_20657);
or UO_2137 (O_2137,N_24378,N_20108);
nand UO_2138 (O_2138,N_19761,N_20400);
nor UO_2139 (O_2139,N_23030,N_23866);
and UO_2140 (O_2140,N_24503,N_24143);
and UO_2141 (O_2141,N_23684,N_20804);
and UO_2142 (O_2142,N_21008,N_19261);
or UO_2143 (O_2143,N_24126,N_20329);
nor UO_2144 (O_2144,N_18942,N_18932);
nand UO_2145 (O_2145,N_19270,N_22712);
and UO_2146 (O_2146,N_20256,N_22727);
nor UO_2147 (O_2147,N_19480,N_24848);
and UO_2148 (O_2148,N_19972,N_22532);
nor UO_2149 (O_2149,N_19364,N_23763);
and UO_2150 (O_2150,N_20792,N_22602);
nor UO_2151 (O_2151,N_24699,N_22508);
or UO_2152 (O_2152,N_19870,N_19822);
nand UO_2153 (O_2153,N_20530,N_19080);
nor UO_2154 (O_2154,N_23967,N_20360);
or UO_2155 (O_2155,N_23057,N_24204);
or UO_2156 (O_2156,N_20092,N_22809);
nand UO_2157 (O_2157,N_18944,N_19979);
nand UO_2158 (O_2158,N_22079,N_22512);
or UO_2159 (O_2159,N_21918,N_24428);
and UO_2160 (O_2160,N_20623,N_22025);
nand UO_2161 (O_2161,N_23380,N_22082);
and UO_2162 (O_2162,N_21642,N_22583);
nand UO_2163 (O_2163,N_21093,N_23858);
and UO_2164 (O_2164,N_21731,N_24885);
or UO_2165 (O_2165,N_24596,N_20702);
and UO_2166 (O_2166,N_20761,N_23311);
or UO_2167 (O_2167,N_20169,N_21851);
nand UO_2168 (O_2168,N_23273,N_23902);
or UO_2169 (O_2169,N_21352,N_24335);
and UO_2170 (O_2170,N_19884,N_24890);
nor UO_2171 (O_2171,N_22302,N_23979);
nand UO_2172 (O_2172,N_24680,N_23413);
and UO_2173 (O_2173,N_20407,N_19613);
nor UO_2174 (O_2174,N_19970,N_24194);
nand UO_2175 (O_2175,N_23163,N_24935);
nand UO_2176 (O_2176,N_23423,N_21019);
or UO_2177 (O_2177,N_24846,N_22832);
nor UO_2178 (O_2178,N_20245,N_21325);
nand UO_2179 (O_2179,N_19222,N_21186);
nand UO_2180 (O_2180,N_20455,N_22506);
or UO_2181 (O_2181,N_22805,N_23698);
nor UO_2182 (O_2182,N_19059,N_22073);
or UO_2183 (O_2183,N_20944,N_19847);
or UO_2184 (O_2184,N_22657,N_22196);
nor UO_2185 (O_2185,N_21775,N_18826);
nor UO_2186 (O_2186,N_22475,N_23337);
and UO_2187 (O_2187,N_23367,N_20825);
nor UO_2188 (O_2188,N_21442,N_23775);
and UO_2189 (O_2189,N_19194,N_23550);
nor UO_2190 (O_2190,N_23327,N_23724);
nor UO_2191 (O_2191,N_20124,N_21073);
and UO_2192 (O_2192,N_22238,N_20669);
and UO_2193 (O_2193,N_22358,N_24322);
or UO_2194 (O_2194,N_19292,N_20122);
nor UO_2195 (O_2195,N_21868,N_21841);
nand UO_2196 (O_2196,N_20506,N_23988);
nand UO_2197 (O_2197,N_23173,N_23574);
or UO_2198 (O_2198,N_22239,N_24967);
nand UO_2199 (O_2199,N_22176,N_21276);
xor UO_2200 (O_2200,N_21433,N_23360);
and UO_2201 (O_2201,N_22567,N_23871);
nor UO_2202 (O_2202,N_19667,N_20975);
nand UO_2203 (O_2203,N_21326,N_24110);
nor UO_2204 (O_2204,N_20872,N_18965);
nor UO_2205 (O_2205,N_23603,N_20751);
or UO_2206 (O_2206,N_22494,N_23096);
nor UO_2207 (O_2207,N_22223,N_22638);
and UO_2208 (O_2208,N_21678,N_20291);
or UO_2209 (O_2209,N_24483,N_23639);
nand UO_2210 (O_2210,N_19772,N_24833);
or UO_2211 (O_2211,N_21332,N_21330);
nand UO_2212 (O_2212,N_22347,N_21943);
or UO_2213 (O_2213,N_19787,N_24060);
or UO_2214 (O_2214,N_24519,N_24403);
nand UO_2215 (O_2215,N_20196,N_24452);
and UO_2216 (O_2216,N_23831,N_19293);
nand UO_2217 (O_2217,N_22819,N_20554);
nand UO_2218 (O_2218,N_20950,N_21795);
and UO_2219 (O_2219,N_24137,N_24715);
or UO_2220 (O_2220,N_24621,N_24181);
or UO_2221 (O_2221,N_21497,N_23118);
and UO_2222 (O_2222,N_24435,N_20276);
nand UO_2223 (O_2223,N_24218,N_20444);
nand UO_2224 (O_2224,N_23606,N_22941);
or UO_2225 (O_2225,N_22624,N_20543);
and UO_2226 (O_2226,N_19139,N_22181);
nand UO_2227 (O_2227,N_22018,N_19767);
or UO_2228 (O_2228,N_20068,N_20197);
nand UO_2229 (O_2229,N_22681,N_24653);
and UO_2230 (O_2230,N_23158,N_19549);
or UO_2231 (O_2231,N_19313,N_18790);
nand UO_2232 (O_2232,N_20725,N_19065);
nand UO_2233 (O_2233,N_22842,N_22229);
and UO_2234 (O_2234,N_22024,N_19681);
nand UO_2235 (O_2235,N_24237,N_21964);
or UO_2236 (O_2236,N_22111,N_19209);
and UO_2237 (O_2237,N_24611,N_21681);
nor UO_2238 (O_2238,N_19121,N_20171);
and UO_2239 (O_2239,N_20200,N_24637);
nor UO_2240 (O_2240,N_20631,N_23680);
and UO_2241 (O_2241,N_23129,N_21715);
nand UO_2242 (O_2242,N_24863,N_20319);
nor UO_2243 (O_2243,N_21889,N_24161);
nand UO_2244 (O_2244,N_20397,N_22027);
nor UO_2245 (O_2245,N_20667,N_22256);
nand UO_2246 (O_2246,N_24499,N_22365);
or UO_2247 (O_2247,N_21659,N_19096);
nor UO_2248 (O_2248,N_20559,N_21469);
nor UO_2249 (O_2249,N_24169,N_24001);
nor UO_2250 (O_2250,N_22237,N_19579);
nor UO_2251 (O_2251,N_19483,N_23026);
and UO_2252 (O_2252,N_24649,N_21399);
or UO_2253 (O_2253,N_22623,N_22854);
nand UO_2254 (O_2254,N_23133,N_20498);
or UO_2255 (O_2255,N_21997,N_21434);
nand UO_2256 (O_2256,N_19181,N_19486);
or UO_2257 (O_2257,N_19042,N_23039);
nor UO_2258 (O_2258,N_19370,N_23803);
nor UO_2259 (O_2259,N_24918,N_19625);
or UO_2260 (O_2260,N_22720,N_20932);
or UO_2261 (O_2261,N_23430,N_21537);
nand UO_2262 (O_2262,N_22396,N_24525);
or UO_2263 (O_2263,N_19377,N_21013);
or UO_2264 (O_2264,N_22268,N_18847);
nor UO_2265 (O_2265,N_23424,N_20285);
nand UO_2266 (O_2266,N_21386,N_22807);
or UO_2267 (O_2267,N_24155,N_22408);
and UO_2268 (O_2268,N_19302,N_21512);
and UO_2269 (O_2269,N_21618,N_19422);
nand UO_2270 (O_2270,N_21181,N_20673);
nand UO_2271 (O_2271,N_20510,N_21261);
and UO_2272 (O_2272,N_21815,N_19338);
nor UO_2273 (O_2273,N_22788,N_21223);
nand UO_2274 (O_2274,N_18975,N_20563);
or UO_2275 (O_2275,N_24239,N_21085);
and UO_2276 (O_2276,N_23043,N_21048);
nor UO_2277 (O_2277,N_18952,N_20351);
nand UO_2278 (O_2278,N_19886,N_19242);
nand UO_2279 (O_2279,N_23632,N_23857);
or UO_2280 (O_2280,N_19684,N_23103);
nand UO_2281 (O_2281,N_19764,N_20268);
or UO_2282 (O_2282,N_19773,N_23102);
or UO_2283 (O_2283,N_18802,N_20081);
and UO_2284 (O_2284,N_19251,N_24623);
nor UO_2285 (O_2285,N_20486,N_19307);
nor UO_2286 (O_2286,N_21732,N_24339);
nand UO_2287 (O_2287,N_21394,N_19191);
nand UO_2288 (O_2288,N_23203,N_22826);
nand UO_2289 (O_2289,N_21925,N_21327);
nor UO_2290 (O_2290,N_18807,N_24760);
nand UO_2291 (O_2291,N_21669,N_18839);
and UO_2292 (O_2292,N_24622,N_24796);
or UO_2293 (O_2293,N_21372,N_21930);
and UO_2294 (O_2294,N_24855,N_20931);
or UO_2295 (O_2295,N_22562,N_24842);
and UO_2296 (O_2296,N_18892,N_18767);
or UO_2297 (O_2297,N_18835,N_19011);
xnor UO_2298 (O_2298,N_19091,N_23069);
or UO_2299 (O_2299,N_18959,N_21595);
and UO_2300 (O_2300,N_24837,N_24557);
nand UO_2301 (O_2301,N_21670,N_19516);
or UO_2302 (O_2302,N_22851,N_22716);
nand UO_2303 (O_2303,N_22189,N_20373);
nor UO_2304 (O_2304,N_20388,N_19971);
and UO_2305 (O_2305,N_22561,N_18977);
or UO_2306 (O_2306,N_20603,N_23678);
and UO_2307 (O_2307,N_19838,N_19137);
nand UO_2308 (O_2308,N_20243,N_21794);
and UO_2309 (O_2309,N_20250,N_19068);
or UO_2310 (O_2310,N_18889,N_24224);
nor UO_2311 (O_2311,N_18921,N_20398);
nand UO_2312 (O_2312,N_21699,N_24279);
and UO_2313 (O_2313,N_19220,N_23227);
and UO_2314 (O_2314,N_21413,N_23488);
or UO_2315 (O_2315,N_21140,N_22317);
or UO_2316 (O_2316,N_24458,N_22045);
and UO_2317 (O_2317,N_20807,N_23335);
or UO_2318 (O_2318,N_24149,N_20327);
and UO_2319 (O_2319,N_23845,N_23880);
or UO_2320 (O_2320,N_19092,N_18821);
nor UO_2321 (O_2321,N_24752,N_23933);
nand UO_2322 (O_2322,N_22677,N_19161);
and UO_2323 (O_2323,N_20231,N_19336);
nand UO_2324 (O_2324,N_24862,N_20568);
nand UO_2325 (O_2325,N_20213,N_20811);
nor UO_2326 (O_2326,N_24812,N_23435);
or UO_2327 (O_2327,N_24754,N_20629);
and UO_2328 (O_2328,N_19531,N_22035);
and UO_2329 (O_2329,N_21550,N_21246);
nor UO_2330 (O_2330,N_23563,N_24517);
nor UO_2331 (O_2331,N_20090,N_22362);
nand UO_2332 (O_2332,N_21942,N_24990);
nand UO_2333 (O_2333,N_22838,N_24740);
nand UO_2334 (O_2334,N_22970,N_21340);
or UO_2335 (O_2335,N_19276,N_21461);
nand UO_2336 (O_2336,N_19572,N_20123);
or UO_2337 (O_2337,N_22499,N_18908);
nor UO_2338 (O_2338,N_21021,N_23874);
nand UO_2339 (O_2339,N_21139,N_24627);
and UO_2340 (O_2340,N_21389,N_21291);
xnor UO_2341 (O_2341,N_20374,N_22230);
or UO_2342 (O_2342,N_20569,N_19628);
or UO_2343 (O_2343,N_22276,N_23317);
nor UO_2344 (O_2344,N_19392,N_22225);
and UO_2345 (O_2345,N_20239,N_22215);
or UO_2346 (O_2346,N_21342,N_20075);
nand UO_2347 (O_2347,N_20311,N_24960);
or UO_2348 (O_2348,N_20469,N_22367);
nor UO_2349 (O_2349,N_19051,N_24502);
nor UO_2350 (O_2350,N_19101,N_23399);
or UO_2351 (O_2351,N_21299,N_24685);
or UO_2352 (O_2352,N_23108,N_24537);
nor UO_2353 (O_2353,N_22307,N_21895);
nand UO_2354 (O_2354,N_19698,N_23225);
nand UO_2355 (O_2355,N_18893,N_20684);
nand UO_2356 (O_2356,N_20716,N_22216);
and UO_2357 (O_2357,N_23726,N_21954);
nor UO_2358 (O_2358,N_20976,N_22031);
nor UO_2359 (O_2359,N_22201,N_24025);
nand UO_2360 (O_2360,N_22156,N_24749);
or UO_2361 (O_2361,N_21217,N_19569);
or UO_2362 (O_2362,N_19284,N_21594);
or UO_2363 (O_2363,N_19740,N_23020);
or UO_2364 (O_2364,N_23495,N_20503);
nand UO_2365 (O_2365,N_20015,N_24396);
nand UO_2366 (O_2366,N_19705,N_22794);
nor UO_2367 (O_2367,N_20589,N_18939);
nand UO_2368 (O_2368,N_24479,N_18857);
and UO_2369 (O_2369,N_21786,N_20042);
or UO_2370 (O_2370,N_20865,N_20915);
and UO_2371 (O_2371,N_19805,N_24551);
nor UO_2372 (O_2372,N_21007,N_21515);
or UO_2373 (O_2373,N_21491,N_24563);
and UO_2374 (O_2374,N_19097,N_20685);
or UO_2375 (O_2375,N_21585,N_19345);
xor UO_2376 (O_2376,N_21949,N_23376);
nor UO_2377 (O_2377,N_21036,N_23941);
or UO_2378 (O_2378,N_22013,N_21982);
nand UO_2379 (O_2379,N_21264,N_19361);
and UO_2380 (O_2380,N_19619,N_22378);
nand UO_2381 (O_2381,N_24687,N_21635);
nand UO_2382 (O_2382,N_23447,N_24247);
nand UO_2383 (O_2383,N_19339,N_23286);
nor UO_2384 (O_2384,N_24241,N_23900);
nand UO_2385 (O_2385,N_20362,N_21554);
and UO_2386 (O_2386,N_18836,N_18822);
or UO_2387 (O_2387,N_23622,N_22676);
nand UO_2388 (O_2388,N_19583,N_20387);
nand UO_2389 (O_2389,N_23994,N_19518);
and UO_2390 (O_2390,N_24017,N_20675);
nand UO_2391 (O_2391,N_24840,N_22783);
or UO_2392 (O_2392,N_20176,N_22777);
or UO_2393 (O_2393,N_19013,N_22756);
nand UO_2394 (O_2394,N_21912,N_20952);
and UO_2395 (O_2395,N_20025,N_22299);
and UO_2396 (O_2396,N_23106,N_20282);
nand UO_2397 (O_2397,N_22001,N_23200);
and UO_2398 (O_2398,N_18760,N_19505);
and UO_2399 (O_2399,N_20292,N_24945);
nand UO_2400 (O_2400,N_20767,N_24352);
nor UO_2401 (O_2401,N_22861,N_22427);
or UO_2402 (O_2402,N_19908,N_20336);
or UO_2403 (O_2403,N_21832,N_23894);
or UO_2404 (O_2404,N_21268,N_24883);
nor UO_2405 (O_2405,N_18794,N_23515);
or UO_2406 (O_2406,N_21783,N_20686);
nor UO_2407 (O_2407,N_22266,N_19340);
nor UO_2408 (O_2408,N_20300,N_22909);
nor UO_2409 (O_2409,N_20580,N_24481);
and UO_2410 (O_2410,N_22247,N_23881);
nor UO_2411 (O_2411,N_20963,N_21035);
and UO_2412 (O_2412,N_23503,N_24497);
and UO_2413 (O_2413,N_21990,N_19316);
or UO_2414 (O_2414,N_23260,N_19241);
nand UO_2415 (O_2415,N_23565,N_23799);
and UO_2416 (O_2416,N_23786,N_22110);
xor UO_2417 (O_2417,N_19067,N_19424);
nor UO_2418 (O_2418,N_18915,N_22267);
nand UO_2419 (O_2419,N_22833,N_21319);
nand UO_2420 (O_2420,N_24225,N_23673);
and UO_2421 (O_2421,N_18827,N_20605);
nor UO_2422 (O_2422,N_22955,N_19620);
nand UO_2423 (O_2423,N_21239,N_24179);
or UO_2424 (O_2424,N_24841,N_23259);
nand UO_2425 (O_2425,N_23377,N_19677);
and UO_2426 (O_2426,N_20097,N_19383);
and UO_2427 (O_2427,N_21762,N_18894);
nand UO_2428 (O_2428,N_23492,N_22662);
nand UO_2429 (O_2429,N_19266,N_20974);
nor UO_2430 (O_2430,N_21563,N_19240);
or UO_2431 (O_2431,N_21107,N_23127);
or UO_2432 (O_2432,N_23821,N_23126);
or UO_2433 (O_2433,N_20534,N_24849);
nand UO_2434 (O_2434,N_19786,N_21829);
nor UO_2435 (O_2435,N_24381,N_24477);
or UO_2436 (O_2436,N_19537,N_22050);
and UO_2437 (O_2437,N_22119,N_23833);
nand UO_2438 (O_2438,N_24549,N_23688);
xnor UO_2439 (O_2439,N_19444,N_23804);
nand UO_2440 (O_2440,N_22919,N_22080);
and UO_2441 (O_2441,N_24354,N_20155);
or UO_2442 (O_2442,N_21746,N_23216);
and UO_2443 (O_2443,N_21279,N_23428);
nand UO_2444 (O_2444,N_21006,N_24983);
or UO_2445 (O_2445,N_20470,N_21234);
nand UO_2446 (O_2446,N_21088,N_22744);
xnor UO_2447 (O_2447,N_22673,N_20072);
nand UO_2448 (O_2448,N_22961,N_21215);
and UO_2449 (O_2449,N_20830,N_21185);
nor UO_2450 (O_2450,N_18853,N_19591);
nor UO_2451 (O_2451,N_20859,N_22132);
and UO_2452 (O_2452,N_22259,N_20480);
nor UO_2453 (O_2453,N_22087,N_23532);
or UO_2454 (O_2454,N_19830,N_19510);
nand UO_2455 (O_2455,N_20058,N_23164);
and UO_2456 (O_2456,N_22969,N_19359);
nand UO_2457 (O_2457,N_20357,N_20033);
and UO_2458 (O_2458,N_19058,N_23531);
nand UO_2459 (O_2459,N_20232,N_21972);
or UO_2460 (O_2460,N_20094,N_21011);
nand UO_2461 (O_2461,N_23044,N_20690);
and UO_2462 (O_2462,N_20954,N_19049);
nand UO_2463 (O_2463,N_24010,N_19214);
nor UO_2464 (O_2464,N_19490,N_20248);
and UO_2465 (O_2465,N_23479,N_21828);
and UO_2466 (O_2466,N_23855,N_22022);
and UO_2467 (O_2467,N_24442,N_21200);
and UO_2468 (O_2468,N_23351,N_21802);
nor UO_2469 (O_2469,N_18877,N_23685);
nor UO_2470 (O_2470,N_18989,N_21773);
or UO_2471 (O_2471,N_24353,N_20910);
or UO_2472 (O_2472,N_19073,N_23796);
or UO_2473 (O_2473,N_20833,N_20352);
nor UO_2474 (O_2474,N_19105,N_19791);
and UO_2475 (O_2475,N_21162,N_24148);
and UO_2476 (O_2476,N_18865,N_21063);
and UO_2477 (O_2477,N_19093,N_23514);
nand UO_2478 (O_2478,N_24777,N_20864);
nand UO_2479 (O_2479,N_24508,N_20763);
or UO_2480 (O_2480,N_22645,N_20158);
nor UO_2481 (O_2481,N_21770,N_21916);
or UO_2482 (O_2482,N_21150,N_24739);
or UO_2483 (O_2483,N_23326,N_19526);
nor UO_2484 (O_2484,N_21409,N_18755);
and UO_2485 (O_2485,N_19728,N_24121);
nor UO_2486 (O_2486,N_22718,N_23918);
or UO_2487 (O_2487,N_21576,N_22020);
and UO_2488 (O_2488,N_22627,N_24510);
nand UO_2489 (O_2489,N_22993,N_22776);
nand UO_2490 (O_2490,N_23568,N_21989);
nand UO_2491 (O_2491,N_19104,N_24113);
and UO_2492 (O_2492,N_23076,N_20542);
nor UO_2493 (O_2493,N_24901,N_24910);
and UO_2494 (O_2494,N_23813,N_19794);
and UO_2495 (O_2495,N_20014,N_19701);
nand UO_2496 (O_2496,N_23374,N_22211);
nand UO_2497 (O_2497,N_24156,N_19935);
and UO_2498 (O_2498,N_22286,N_22597);
nor UO_2499 (O_2499,N_23074,N_19418);
and UO_2500 (O_2500,N_24547,N_20882);
nand UO_2501 (O_2501,N_24142,N_21226);
and UO_2502 (O_2502,N_23841,N_23691);
nor UO_2503 (O_2503,N_24516,N_23761);
and UO_2504 (O_2504,N_22232,N_23140);
or UO_2505 (O_2505,N_20214,N_19581);
and UO_2506 (O_2506,N_24344,N_21037);
nand UO_2507 (O_2507,N_23720,N_23923);
nor UO_2508 (O_2508,N_24478,N_20877);
nand UO_2509 (O_2509,N_22553,N_21546);
nor UO_2510 (O_2510,N_23264,N_19443);
or UO_2511 (O_2511,N_21086,N_20249);
nor UO_2512 (O_2512,N_23560,N_23266);
nor UO_2513 (O_2513,N_18841,N_20688);
nand UO_2514 (O_2514,N_21506,N_23961);
or UO_2515 (O_2515,N_21529,N_21545);
nand UO_2516 (O_2516,N_19107,N_19616);
xor UO_2517 (O_2517,N_20959,N_24267);
nor UO_2518 (O_2518,N_24864,N_22965);
nand UO_2519 (O_2519,N_20442,N_22048);
nand UO_2520 (O_2520,N_22988,N_21015);
and UO_2521 (O_2521,N_24625,N_21660);
nand UO_2522 (O_2522,N_19381,N_20168);
and UO_2523 (O_2523,N_20128,N_19836);
or UO_2524 (O_2524,N_22220,N_22459);
and UO_2525 (O_2525,N_19026,N_24425);
and UO_2526 (O_2526,N_24696,N_19410);
nor UO_2527 (O_2527,N_24188,N_24987);
or UO_2528 (O_2528,N_18991,N_21464);
or UO_2529 (O_2529,N_23493,N_19257);
or UO_2530 (O_2530,N_20431,N_22895);
nand UO_2531 (O_2531,N_22992,N_22781);
and UO_2532 (O_2532,N_24781,N_19036);
nand UO_2533 (O_2533,N_22462,N_23445);
or UO_2534 (O_2534,N_24857,N_19484);
and UO_2535 (O_2535,N_20665,N_23816);
nand UO_2536 (O_2536,N_24904,N_24651);
nand UO_2537 (O_2537,N_21480,N_22246);
and UO_2538 (O_2538,N_18834,N_20978);
nor UO_2539 (O_2539,N_18928,N_20338);
nor UO_2540 (O_2540,N_23201,N_24894);
nor UO_2541 (O_2541,N_23060,N_21192);
nand UO_2542 (O_2542,N_22521,N_24764);
or UO_2543 (O_2543,N_24229,N_20728);
or UO_2544 (O_2544,N_19754,N_21948);
and UO_2545 (O_2545,N_23412,N_24129);
nor UO_2546 (O_2546,N_21953,N_22327);
or UO_2547 (O_2547,N_24518,N_18887);
nor UO_2548 (O_2548,N_21547,N_24004);
and UO_2549 (O_2549,N_21904,N_20022);
or UO_2550 (O_2550,N_20799,N_19438);
and UO_2551 (O_2551,N_23056,N_23333);
nor UO_2552 (O_2552,N_19452,N_20699);
nor UO_2553 (O_2553,N_21402,N_20851);
xor UO_2554 (O_2554,N_24259,N_21666);
nor UO_2555 (O_2555,N_24341,N_23516);
nand UO_2556 (O_2556,N_20102,N_23395);
nand UO_2557 (O_2557,N_24579,N_21177);
nand UO_2558 (O_2558,N_20085,N_23429);
or UO_2559 (O_2559,N_21099,N_19140);
or UO_2560 (O_2560,N_22075,N_22835);
and UO_2561 (O_2561,N_21739,N_22655);
or UO_2562 (O_2562,N_23878,N_23911);
nor UO_2563 (O_2563,N_23641,N_19066);
and UO_2564 (O_2564,N_20460,N_21858);
xor UO_2565 (O_2565,N_24220,N_24543);
or UO_2566 (O_2566,N_22543,N_19967);
nor UO_2567 (O_2567,N_22912,N_24331);
and UO_2568 (O_2568,N_21853,N_24607);
nor UO_2569 (O_2569,N_20386,N_24095);
nor UO_2570 (O_2570,N_24262,N_19162);
nor UO_2571 (O_2571,N_21763,N_24706);
nand UO_2572 (O_2572,N_24845,N_24654);
nand UO_2573 (O_2573,N_19604,N_19785);
nor UO_2574 (O_2574,N_24283,N_20144);
nand UO_2575 (O_2575,N_22485,N_24807);
and UO_2576 (O_2576,N_21398,N_21639);
and UO_2577 (O_2577,N_24112,N_21611);
nor UO_2578 (O_2578,N_19087,N_20012);
or UO_2579 (O_2579,N_18768,N_23234);
nor UO_2580 (O_2580,N_24385,N_20481);
or UO_2581 (O_2581,N_24662,N_18858);
or UO_2582 (O_2582,N_24509,N_20988);
and UO_2583 (O_2583,N_21316,N_19682);
nand UO_2584 (O_2584,N_22450,N_24250);
or UO_2585 (O_2585,N_21175,N_20227);
nor UO_2586 (O_2586,N_22708,N_19859);
nand UO_2587 (O_2587,N_21456,N_21376);
and UO_2588 (O_2588,N_21944,N_24432);
nor UO_2589 (O_2589,N_22732,N_20518);
nor UO_2590 (O_2590,N_20525,N_20837);
nand UO_2591 (O_2591,N_19651,N_19117);
or UO_2592 (O_2592,N_20785,N_21228);
nor UO_2593 (O_2593,N_19039,N_24644);
nor UO_2594 (O_2594,N_22692,N_21041);
or UO_2595 (O_2595,N_24325,N_24138);
and UO_2596 (O_2596,N_19115,N_23690);
and UO_2597 (O_2597,N_23018,N_19285);
and UO_2598 (O_2598,N_23110,N_24040);
and UO_2599 (O_2599,N_21082,N_22303);
nor UO_2600 (O_2600,N_19273,N_23628);
and UO_2601 (O_2601,N_20405,N_24851);
or UO_2602 (O_2602,N_19485,N_20027);
nor UO_2603 (O_2603,N_22938,N_21649);
nor UO_2604 (O_2604,N_19649,N_23385);
and UO_2605 (O_2605,N_23848,N_21738);
or UO_2606 (O_2606,N_19341,N_22690);
nand UO_2607 (O_2607,N_19617,N_20299);
nor UO_2608 (O_2608,N_24315,N_22846);
nand UO_2609 (O_2609,N_19907,N_21683);
or UO_2610 (O_2610,N_19645,N_22469);
nand UO_2611 (O_2611,N_20784,N_24255);
nor UO_2612 (O_2612,N_21663,N_24788);
nor UO_2613 (O_2613,N_24574,N_21979);
or UO_2614 (O_2614,N_18898,N_22301);
nor UO_2615 (O_2615,N_19905,N_20624);
xor UO_2616 (O_2616,N_19146,N_21646);
nand UO_2617 (O_2617,N_20477,N_21962);
and UO_2618 (O_2618,N_19683,N_24583);
nand UO_2619 (O_2619,N_21526,N_19184);
and UO_2620 (O_2620,N_23342,N_23368);
nor UO_2621 (O_2621,N_19371,N_22711);
nand UO_2622 (O_2622,N_23943,N_23733);
and UO_2623 (O_2623,N_23689,N_19165);
nor UO_2624 (O_2624,N_20597,N_24488);
nor UO_2625 (O_2625,N_19610,N_20923);
or UO_2626 (O_2626,N_21148,N_21653);
nor UO_2627 (O_2627,N_23301,N_22129);
and UO_2628 (O_2628,N_19878,N_18806);
nor UO_2629 (O_2629,N_18784,N_19053);
nand UO_2630 (O_2630,N_23253,N_24389);
and UO_2631 (O_2631,N_19653,N_20452);
and UO_2632 (O_2632,N_19892,N_23832);
or UO_2633 (O_2633,N_20065,N_22724);
nand UO_2634 (O_2634,N_19941,N_22363);
nor UO_2635 (O_2635,N_24742,N_22628);
nor UO_2636 (O_2636,N_24608,N_24445);
or UO_2637 (O_2637,N_23649,N_19109);
nor UO_2638 (O_2638,N_23467,N_20615);
or UO_2639 (O_2639,N_22448,N_24873);
nand UO_2640 (O_2640,N_22633,N_19936);
and UO_2641 (O_2641,N_23454,N_19576);
or UO_2642 (O_2642,N_19776,N_20093);
nor UO_2643 (O_2643,N_24209,N_24529);
nand UO_2644 (O_2644,N_20899,N_22145);
nand UO_2645 (O_2645,N_21284,N_23359);
nor UO_2646 (O_2646,N_20113,N_21896);
or UO_2647 (O_2647,N_18848,N_20326);
nand UO_2648 (O_2648,N_22158,N_21033);
and UO_2649 (O_2649,N_19632,N_20762);
and UO_2650 (O_2650,N_19294,N_20758);
nand UO_2651 (O_2651,N_19768,N_19952);
and UO_2652 (O_2652,N_24986,N_23850);
nor UO_2653 (O_2653,N_23284,N_22350);
or UO_2654 (O_2654,N_22702,N_19873);
and UO_2655 (O_2655,N_21826,N_19322);
nand UO_2656 (O_2656,N_22214,N_24746);
nor UO_2657 (O_2657,N_21720,N_19955);
nand UO_2658 (O_2658,N_20151,N_24082);
nand UO_2659 (O_2659,N_19379,N_23143);
or UO_2660 (O_2660,N_24056,N_19731);
or UO_2661 (O_2661,N_22525,N_24368);
and UO_2662 (O_2662,N_18972,N_22069);
nor UO_2663 (O_2663,N_21717,N_18948);
and UO_2664 (O_2664,N_20458,N_19564);
and UO_2665 (O_2665,N_21245,N_20995);
and UO_2666 (O_2666,N_22710,N_21240);
or UO_2667 (O_2667,N_23765,N_18782);
and UO_2668 (O_2668,N_22039,N_21244);
nor UO_2669 (O_2669,N_22626,N_19512);
or UO_2670 (O_2670,N_24264,N_21654);
nand UO_2671 (O_2671,N_19164,N_20194);
nor UO_2672 (O_2672,N_24476,N_21128);
nand UO_2673 (O_2673,N_20354,N_22541);
and UO_2674 (O_2674,N_23464,N_19949);
and UO_2675 (O_2675,N_24613,N_20717);
and UO_2676 (O_2676,N_20892,N_20138);
or UO_2677 (O_2677,N_19464,N_18934);
nor UO_2678 (O_2678,N_19513,N_23042);
or UO_2679 (O_2679,N_24920,N_21058);
and UO_2680 (O_2680,N_19327,N_21108);
or UO_2681 (O_2681,N_23600,N_22925);
or UO_2682 (O_2682,N_20116,N_20539);
and UO_2683 (O_2683,N_23935,N_23306);
nand UO_2684 (O_2684,N_23276,N_19474);
nand UO_2685 (O_2685,N_23197,N_19695);
nand UO_2686 (O_2686,N_18918,N_22100);
nand UO_2687 (O_2687,N_22971,N_21127);
or UO_2688 (O_2688,N_20547,N_22453);
or UO_2689 (O_2689,N_24630,N_18960);
nand UO_2690 (O_2690,N_22636,N_21141);
nand UO_2691 (O_2691,N_21489,N_20279);
nor UO_2692 (O_2692,N_23051,N_24783);
nand UO_2693 (O_2693,N_22356,N_24130);
or UO_2694 (O_2694,N_24911,N_21532);
nand UO_2695 (O_2695,N_19280,N_21874);
nor UO_2696 (O_2696,N_23807,N_23909);
or UO_2697 (O_2697,N_23332,N_21315);
or UO_2698 (O_2698,N_20026,N_24314);
nor UO_2699 (O_2699,N_21400,N_19238);
nand UO_2700 (O_2700,N_22240,N_19212);
or UO_2701 (O_2701,N_21691,N_18772);
and UO_2702 (O_2702,N_23046,N_21844);
and UO_2703 (O_2703,N_22952,N_21976);
or UO_2704 (O_2704,N_19095,N_20775);
and UO_2705 (O_2705,N_22683,N_19495);
or UO_2706 (O_2706,N_22916,N_24309);
or UO_2707 (O_2707,N_19983,N_23605);
nand UO_2708 (O_2708,N_22152,N_23945);
or UO_2709 (O_2709,N_22096,N_20891);
xor UO_2710 (O_2710,N_20745,N_19103);
or UO_2711 (O_2711,N_20190,N_22563);
and UO_2712 (O_2712,N_20348,N_24349);
or UO_2713 (O_2713,N_23490,N_19845);
nor UO_2714 (O_2714,N_23818,N_22360);
or UO_2715 (O_2715,N_20310,N_24062);
or UO_2716 (O_2716,N_24757,N_19546);
nor UO_2717 (O_2717,N_18954,N_20828);
or UO_2718 (O_2718,N_21688,N_24398);
or UO_2719 (O_2719,N_24828,N_24564);
nand UO_2720 (O_2720,N_19733,N_19047);
and UO_2721 (O_2721,N_19933,N_24695);
or UO_2722 (O_2722,N_18849,N_21441);
and UO_2723 (O_2723,N_19004,N_21615);
nor UO_2724 (O_2724,N_21601,N_23643);
nand UO_2725 (O_2725,N_20748,N_19635);
and UO_2726 (O_2726,N_21271,N_23403);
nand UO_2727 (O_2727,N_23980,N_22648);
nor UO_2728 (O_2728,N_22524,N_24207);
nand UO_2729 (O_2729,N_22985,N_21648);
nand UO_2730 (O_2730,N_23040,N_20435);
or UO_2731 (O_2731,N_23917,N_23053);
nor UO_2732 (O_2732,N_21220,N_19351);
or UO_2733 (O_2733,N_19070,N_23409);
or UO_2734 (O_2734,N_20838,N_22814);
nor UO_2735 (O_2735,N_21525,N_19407);
nand UO_2736 (O_2736,N_22468,N_24973);
and UO_2737 (O_2737,N_20132,N_23835);
or UO_2738 (O_2738,N_22924,N_23963);
nor UO_2739 (O_2739,N_21987,N_24014);
nor UO_2740 (O_2740,N_19045,N_23257);
nand UO_2741 (O_2741,N_21373,N_23471);
nand UO_2742 (O_2742,N_23856,N_21320);
nand UO_2743 (O_2743,N_22666,N_24882);
or UO_2744 (O_2744,N_23784,N_21481);
or UO_2745 (O_2745,N_23703,N_19254);
nand UO_2746 (O_2746,N_22804,N_24216);
nand UO_2747 (O_2747,N_20779,N_20032);
nand UO_2748 (O_2748,N_20653,N_21493);
nor UO_2749 (O_2749,N_24460,N_20323);
nand UO_2750 (O_2750,N_22536,N_24718);
nor UO_2751 (O_2751,N_24390,N_23339);
and UO_2752 (O_2752,N_19078,N_22105);
nor UO_2753 (O_2753,N_21564,N_22897);
nand UO_2754 (O_2754,N_20759,N_21248);
nor UO_2755 (O_2755,N_21263,N_19368);
or UO_2756 (O_2756,N_24787,N_18810);
or UO_2757 (O_2757,N_23509,N_21514);
nor UO_2758 (O_2758,N_19024,N_21588);
nand UO_2759 (O_2759,N_20886,N_22387);
nor UO_2760 (O_2760,N_19151,N_20531);
xor UO_2761 (O_2761,N_24063,N_20414);
or UO_2762 (O_2762,N_23058,N_19696);
nor UO_2763 (O_2763,N_24850,N_21370);
nor UO_2764 (O_2764,N_22164,N_24357);
or UO_2765 (O_2765,N_18936,N_24880);
or UO_2766 (O_2766,N_21339,N_20039);
and UO_2767 (O_2767,N_21707,N_20016);
nor UO_2768 (O_2768,N_20281,N_21572);
nand UO_2769 (O_2769,N_21680,N_21539);
or UO_2770 (O_2770,N_21333,N_20780);
nor UO_2771 (O_2771,N_22349,N_19923);
nand UO_2772 (O_2772,N_21754,N_22598);
and UO_2773 (O_2773,N_24530,N_19749);
nand UO_2774 (O_2774,N_24135,N_24304);
nor UO_2775 (O_2775,N_20314,N_20406);
nor UO_2776 (O_2776,N_21625,N_19023);
xnor UO_2777 (O_2777,N_19127,N_24769);
nor UO_2778 (O_2778,N_21379,N_19780);
nand UO_2779 (O_2779,N_19762,N_22911);
or UO_2780 (O_2780,N_19128,N_20385);
and UO_2781 (O_2781,N_20247,N_20630);
nor UO_2782 (O_2782,N_24246,N_22738);
and UO_2783 (O_2783,N_20706,N_20795);
nand UO_2784 (O_2784,N_23232,N_24330);
or UO_2785 (O_2785,N_21825,N_24614);
nor UO_2786 (O_2786,N_24731,N_19680);
nand UO_2787 (O_2787,N_24294,N_20968);
or UO_2788 (O_2788,N_23944,N_22531);
and UO_2789 (O_2789,N_23650,N_23937);
or UO_2790 (O_2790,N_24201,N_21692);
nor UO_2791 (O_2791,N_23728,N_22144);
nor UO_2792 (O_2792,N_24276,N_22305);
and UO_2793 (O_2793,N_21027,N_19621);
and UO_2794 (O_2794,N_20349,N_20868);
or UO_2795 (O_2795,N_20101,N_24772);
nand UO_2796 (O_2796,N_23543,N_23829);
and UO_2797 (O_2797,N_24792,N_21328);
nor UO_2798 (O_2798,N_20233,N_21842);
or UO_2799 (O_2799,N_21812,N_20823);
nor UO_2800 (O_2800,N_23893,N_23756);
nand UO_2801 (O_2801,N_22028,N_21130);
nor UO_2802 (O_2802,N_20491,N_24603);
and UO_2803 (O_2803,N_21686,N_19541);
and UO_2804 (O_2804,N_19655,N_19856);
nor UO_2805 (O_2805,N_20800,N_19718);
nand UO_2806 (O_2806,N_20007,N_22820);
or UO_2807 (O_2807,N_18999,N_22495);
and UO_2808 (O_2808,N_23036,N_19465);
nand UO_2809 (O_2809,N_22701,N_18979);
or UO_2810 (O_2810,N_19580,N_24981);
and UO_2811 (O_2811,N_18923,N_23151);
and UO_2812 (O_2812,N_23021,N_23090);
and UO_2813 (O_2813,N_19850,N_20488);
nand UO_2814 (O_2814,N_19897,N_20507);
or UO_2815 (O_2815,N_21998,N_24141);
nor UO_2816 (O_2816,N_24528,N_20322);
or UO_2817 (O_2817,N_20604,N_22709);
nor UO_2818 (O_2818,N_22142,N_19888);
and UO_2819 (O_2819,N_20906,N_18793);
and UO_2820 (O_2820,N_19425,N_20708);
nor UO_2821 (O_2821,N_22697,N_24057);
nand UO_2822 (O_2822,N_20468,N_18950);
nand UO_2823 (O_2823,N_21792,N_21334);
or UO_2824 (O_2824,N_19709,N_18970);
nand UO_2825 (O_2825,N_20663,N_22109);
nor UO_2826 (O_2826,N_21424,N_24668);
nor UO_2827 (O_2827,N_24111,N_24859);
or UO_2828 (O_2828,N_21484,N_21900);
and UO_2829 (O_2829,N_20389,N_18801);
nand UO_2830 (O_2830,N_21804,N_21613);
and UO_2831 (O_2831,N_20135,N_20257);
and UO_2832 (O_2832,N_19038,N_19044);
or UO_2833 (O_2833,N_22675,N_19229);
nand UO_2834 (O_2834,N_20109,N_19405);
and UO_2835 (O_2835,N_19329,N_20560);
or UO_2836 (O_2836,N_19267,N_24005);
and UO_2837 (O_2837,N_22768,N_21156);
or UO_2838 (O_2838,N_22606,N_20714);
or UO_2839 (O_2839,N_24456,N_19975);
nor UO_2840 (O_2840,N_24434,N_21457);
nand UO_2841 (O_2841,N_22200,N_19509);
or UO_2842 (O_2842,N_23211,N_23730);
nand UO_2843 (O_2843,N_20195,N_24964);
nor UO_2844 (O_2844,N_24555,N_22546);
nor UO_2845 (O_2845,N_23915,N_21430);
nor UO_2846 (O_2846,N_23458,N_22876);
or UO_2847 (O_2847,N_22261,N_19286);
and UO_2848 (O_2848,N_20275,N_24747);
and UO_2849 (O_2849,N_21323,N_24128);
nor UO_2850 (O_2850,N_21903,N_24875);
and UO_2851 (O_2851,N_24467,N_19385);
nand UO_2852 (O_2852,N_18820,N_21146);
nor UO_2853 (O_2853,N_20713,N_18824);
nor UO_2854 (O_2854,N_22203,N_20165);
nor UO_2855 (O_2855,N_23859,N_19816);
or UO_2856 (O_2856,N_24242,N_21561);
nand UO_2857 (O_2857,N_19753,N_24272);
and UO_2858 (O_2858,N_23589,N_23811);
nand UO_2859 (O_2859,N_19977,N_24912);
nand UO_2860 (O_2860,N_22496,N_24092);
nor UO_2861 (O_2861,N_20897,N_19686);
nand UO_2862 (O_2862,N_23991,N_24310);
or UO_2863 (O_2863,N_20705,N_19441);
and UO_2864 (O_2864,N_19732,N_21675);
nor UO_2865 (O_2865,N_20729,N_23011);
nor UO_2866 (O_2866,N_23590,N_19037);
or UO_2867 (O_2867,N_21292,N_19802);
and UO_2868 (O_2868,N_21032,N_23654);
nand UO_2869 (O_2869,N_21899,N_19875);
or UO_2870 (O_2870,N_21816,N_20796);
and UO_2871 (O_2871,N_22609,N_21026);
nor UO_2872 (O_2872,N_22950,N_24256);
and UO_2873 (O_2873,N_22707,N_20206);
nand UO_2874 (O_2874,N_20371,N_18805);
nand UO_2875 (O_2875,N_23443,N_22793);
nand UO_2876 (O_2876,N_21081,N_19827);
nor UO_2877 (O_2877,N_23592,N_19554);
nand UO_2878 (O_2878,N_23427,N_24051);
and UO_2879 (O_2879,N_21719,N_22443);
and UO_2880 (O_2880,N_23346,N_20467);
nor UO_2881 (O_2881,N_24712,N_19969);
nor UO_2882 (O_2882,N_20289,N_24944);
or UO_2883 (O_2883,N_23793,N_24450);
nor UO_2884 (O_2884,N_21306,N_19719);
nand UO_2885 (O_2885,N_23778,N_19874);
and UO_2886 (O_2886,N_19311,N_23573);
nand UO_2887 (O_2887,N_23105,N_22472);
or UO_2888 (O_2888,N_23709,N_22743);
nor UO_2889 (O_2889,N_19729,N_19606);
nand UO_2890 (O_2890,N_19187,N_20238);
nand UO_2891 (O_2891,N_21249,N_19141);
nor UO_2892 (O_2892,N_22398,N_23921);
and UO_2893 (O_2893,N_18773,N_24939);
and UO_2894 (O_2894,N_24448,N_21311);
nor UO_2895 (O_2895,N_24470,N_20948);
or UO_2896 (O_2896,N_21479,N_19007);
nand UO_2897 (O_2897,N_21541,N_19415);
nand UO_2898 (O_2898,N_24430,N_24577);
or UO_2899 (O_2899,N_23642,N_22739);
or UO_2900 (O_2900,N_22937,N_21534);
nand UO_2901 (O_2901,N_19693,N_23198);
nor UO_2902 (O_2902,N_20426,N_20810);
nor UO_2903 (O_2903,N_19110,N_19962);
nor UO_2904 (O_2904,N_19114,N_20237);
or UO_2905 (O_2905,N_22424,N_19568);
nor UO_2906 (O_2906,N_20930,N_22140);
nand UO_2907 (O_2907,N_19618,N_22844);
nand UO_2908 (O_2908,N_21222,N_18844);
nor UO_2909 (O_2909,N_20205,N_20935);
nand UO_2910 (O_2910,N_20942,N_20596);
nor UO_2911 (O_2911,N_19204,N_21294);
nand UO_2912 (O_2912,N_20236,N_21810);
nand UO_2913 (O_2913,N_24844,N_24441);
nor UO_2914 (O_2914,N_19489,N_21556);
or UO_2915 (O_2915,N_22354,N_18878);
or UO_2916 (O_2916,N_20226,N_22486);
nor UO_2917 (O_2917,N_23539,N_18998);
nor UO_2918 (O_2918,N_24744,N_23769);
and UO_2919 (O_2919,N_21803,N_24816);
xor UO_2920 (O_2920,N_21822,N_19795);
or UO_2921 (O_2921,N_24326,N_23872);
and UO_2922 (O_2922,N_22554,N_24296);
or UO_2923 (O_2923,N_24427,N_22092);
nand UO_2924 (O_2924,N_20463,N_21941);
nor UO_2925 (O_2925,N_22046,N_20447);
or UO_2926 (O_2926,N_19005,N_22175);
nand UO_2927 (O_2927,N_21475,N_20382);
nor UO_2928 (O_2928,N_21638,N_20089);
nand UO_2929 (O_2929,N_19175,N_19504);
and UO_2930 (O_2930,N_23062,N_24867);
nand UO_2931 (O_2931,N_24866,N_18842);
nand UO_2932 (O_2932,N_20208,N_19919);
and UO_2933 (O_2933,N_22065,N_23093);
or UO_2934 (O_2934,N_22917,N_19430);
nand UO_2935 (O_2935,N_24838,N_24221);
or UO_2936 (O_2936,N_20107,N_24087);
nand UO_2937 (O_2937,N_19295,N_23438);
nand UO_2938 (O_2938,N_20112,N_23585);
nor UO_2939 (O_2939,N_23548,N_20018);
nand UO_2940 (O_2940,N_19792,N_20946);
or UO_2941 (O_2941,N_19459,N_21259);
nand UO_2942 (O_2942,N_22654,N_24132);
xnor UO_2943 (O_2943,N_19503,N_22608);
nor UO_2944 (O_2944,N_23955,N_18779);
nor UO_2945 (O_2945,N_24562,N_20739);
and UO_2946 (O_2946,N_24933,N_23474);
and UO_2947 (O_2947,N_24821,N_18774);
nand UO_2948 (O_2948,N_20290,N_21913);
and UO_2949 (O_2949,N_23624,N_20130);
or UO_2950 (O_2950,N_23487,N_22032);
or UO_2951 (O_2951,N_19737,N_18927);
and UO_2952 (O_2952,N_22391,N_19690);
nand UO_2953 (O_2953,N_19369,N_19890);
nand UO_2954 (O_2954,N_21596,N_22177);
or UO_2955 (O_2955,N_22343,N_21499);
nand UO_2956 (O_2956,N_21967,N_23562);
and UO_2957 (O_2957,N_19353,N_22260);
nand UO_2958 (O_2958,N_19717,N_21168);
and UO_2959 (O_2959,N_21721,N_21791);
and UO_2960 (O_2960,N_22265,N_21766);
nor UO_2961 (O_2961,N_20736,N_23283);
and UO_2962 (O_2962,N_23045,N_21991);
or UO_2963 (O_2963,N_19131,N_21445);
or UO_2964 (O_2964,N_24725,N_19527);
or UO_2965 (O_2965,N_18955,N_22264);
or UO_2966 (O_2966,N_22290,N_19657);
and UO_2967 (O_2967,N_22322,N_20857);
nand UO_2968 (O_2968,N_21116,N_22791);
nor UO_2969 (O_2969,N_22219,N_19416);
nor UO_2970 (O_2970,N_22730,N_20561);
nand UO_2971 (O_2971,N_22137,N_23091);
or UO_2972 (O_2972,N_21553,N_23700);
and UO_2973 (O_2973,N_20501,N_21367);
nor UO_2974 (O_2974,N_22953,N_20704);
nor UO_2975 (O_2975,N_19548,N_19910);
nor UO_2976 (O_2976,N_23155,N_19426);
or UO_2977 (O_2977,N_20394,N_23139);
nor UO_2978 (O_2978,N_24690,N_22998);
and UO_2979 (O_2979,N_22522,N_21559);
nand UO_2980 (O_2980,N_24162,N_24401);
and UO_2981 (O_2981,N_23263,N_19413);
nand UO_2982 (O_2982,N_24288,N_24923);
and UO_2983 (O_2983,N_20161,N_24387);
and UO_2984 (O_2984,N_23768,N_23235);
nand UO_2985 (O_2985,N_21849,N_23117);
nor UO_2986 (O_2986,N_23610,N_19648);
nor UO_2987 (O_2987,N_20937,N_20956);
nor UO_2988 (O_2988,N_21253,N_23595);
and UO_2989 (O_2989,N_21651,N_20497);
and UO_2990 (O_2990,N_23555,N_24552);
or UO_2991 (O_2991,N_19959,N_18854);
and UO_2992 (O_2992,N_24632,N_21465);
nand UO_2993 (O_2993,N_24091,N_20391);
nand UO_2994 (O_2994,N_21285,N_19163);
nand UO_2995 (O_2995,N_21655,N_22431);
or UO_2996 (O_2996,N_21492,N_19071);
and UO_2997 (O_2997,N_20050,N_23743);
nor UO_2998 (O_2998,N_21025,N_22040);
or UO_2999 (O_2999,N_22042,N_23583);
endmodule