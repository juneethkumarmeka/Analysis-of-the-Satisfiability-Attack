module basic_1000_10000_1500_4_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_302,In_670);
nand U1 (N_1,In_730,In_387);
nand U2 (N_2,In_309,In_767);
xnor U3 (N_3,In_757,In_173);
nand U4 (N_4,In_347,In_53);
nand U5 (N_5,In_36,In_571);
nor U6 (N_6,In_884,In_439);
nand U7 (N_7,In_429,In_837);
nand U8 (N_8,In_545,In_324);
nand U9 (N_9,In_154,In_821);
nor U10 (N_10,In_880,In_345);
and U11 (N_11,In_51,In_400);
xnor U12 (N_12,In_944,In_856);
and U13 (N_13,In_591,In_224);
nor U14 (N_14,In_13,In_815);
nor U15 (N_15,In_564,In_71);
nand U16 (N_16,In_306,In_391);
xor U17 (N_17,In_998,In_747);
and U18 (N_18,In_540,In_739);
nand U19 (N_19,In_983,In_311);
xor U20 (N_20,In_640,In_575);
nor U21 (N_21,In_548,In_431);
nor U22 (N_22,In_130,In_1);
nand U23 (N_23,In_898,In_796);
nand U24 (N_24,In_599,In_312);
nor U25 (N_25,In_82,In_723);
xnor U26 (N_26,In_337,In_778);
nor U27 (N_27,In_368,In_425);
nand U28 (N_28,In_350,In_847);
and U29 (N_29,In_577,In_83);
or U30 (N_30,In_166,In_681);
xnor U31 (N_31,In_634,In_612);
or U32 (N_32,In_893,In_822);
nor U33 (N_33,In_164,In_489);
and U34 (N_34,In_26,In_220);
nand U35 (N_35,In_786,In_121);
nand U36 (N_36,In_642,In_484);
nand U37 (N_37,In_505,In_385);
or U38 (N_38,In_946,In_92);
nor U39 (N_39,In_56,In_346);
or U40 (N_40,In_883,In_222);
xor U41 (N_41,In_19,In_60);
nor U42 (N_42,In_945,In_598);
or U43 (N_43,In_982,In_626);
or U44 (N_44,In_218,In_0);
and U45 (N_45,In_755,In_105);
nand U46 (N_46,In_442,In_31);
nor U47 (N_47,In_999,In_911);
nor U48 (N_48,In_234,In_852);
or U49 (N_49,In_838,In_625);
nand U50 (N_50,In_644,In_759);
nand U51 (N_51,In_78,In_86);
nand U52 (N_52,In_353,In_799);
nand U53 (N_53,In_965,In_968);
or U54 (N_54,In_809,In_994);
or U55 (N_55,In_95,In_433);
nand U56 (N_56,In_419,In_294);
or U57 (N_57,In_443,In_453);
or U58 (N_58,In_647,In_89);
nand U59 (N_59,In_33,In_275);
and U60 (N_60,In_136,In_572);
or U61 (N_61,In_280,In_584);
nor U62 (N_62,In_903,In_587);
and U63 (N_63,In_805,In_395);
xor U64 (N_64,In_282,In_909);
and U65 (N_65,In_293,In_219);
nor U66 (N_66,In_549,In_25);
nor U67 (N_67,In_621,In_300);
nand U68 (N_68,In_596,In_382);
nand U69 (N_69,In_356,In_555);
nor U70 (N_70,In_529,In_694);
or U71 (N_71,In_11,In_349);
nor U72 (N_72,In_891,In_508);
xor U73 (N_73,In_230,In_12);
nor U74 (N_74,In_863,In_886);
nand U75 (N_75,In_14,In_929);
nand U76 (N_76,In_476,In_848);
and U77 (N_77,In_660,In_969);
and U78 (N_78,In_704,In_99);
or U79 (N_79,In_738,In_879);
nor U80 (N_80,In_372,In_791);
or U81 (N_81,In_284,In_562);
nand U82 (N_82,In_779,In_298);
nand U83 (N_83,In_351,In_790);
or U84 (N_84,In_180,In_393);
nand U85 (N_85,In_134,In_265);
and U86 (N_86,In_978,In_645);
and U87 (N_87,In_405,In_766);
nor U88 (N_88,In_470,In_861);
nand U89 (N_89,In_373,In_97);
nor U90 (N_90,In_711,In_667);
xor U91 (N_91,In_643,In_620);
and U92 (N_92,In_594,In_524);
nor U93 (N_93,In_227,In_901);
nand U94 (N_94,In_194,In_836);
and U95 (N_95,In_788,In_183);
nor U96 (N_96,In_614,In_283);
and U97 (N_97,In_421,In_709);
or U98 (N_98,In_876,In_396);
and U99 (N_99,In_444,In_123);
nor U100 (N_100,In_938,In_897);
and U101 (N_101,In_922,In_192);
or U102 (N_102,In_966,In_942);
xor U103 (N_103,In_521,In_812);
nor U104 (N_104,In_633,In_910);
nor U105 (N_105,In_558,In_992);
or U106 (N_106,In_731,In_223);
and U107 (N_107,In_141,In_517);
nand U108 (N_108,In_606,In_961);
or U109 (N_109,In_912,In_195);
nor U110 (N_110,In_157,In_340);
and U111 (N_111,In_343,In_330);
and U112 (N_112,In_394,In_556);
nor U113 (N_113,In_972,In_253);
nand U114 (N_114,In_240,In_468);
nor U115 (N_115,In_652,In_427);
and U116 (N_116,In_725,In_657);
or U117 (N_117,In_760,In_986);
or U118 (N_118,In_658,In_635);
and U119 (N_119,In_701,In_55);
nor U120 (N_120,In_366,In_411);
and U121 (N_121,In_816,In_187);
nor U122 (N_122,In_299,In_472);
and U123 (N_123,In_827,In_46);
and U124 (N_124,In_979,In_456);
nor U125 (N_125,In_441,In_563);
nor U126 (N_126,In_930,In_65);
nand U127 (N_127,In_926,In_266);
and U128 (N_128,In_737,In_34);
or U129 (N_129,In_868,In_169);
xor U130 (N_130,In_313,In_526);
or U131 (N_131,In_402,In_301);
and U132 (N_132,In_954,In_384);
xor U133 (N_133,In_165,In_920);
and U134 (N_134,In_995,In_291);
nor U135 (N_135,In_10,In_480);
nor U136 (N_136,In_754,In_854);
and U137 (N_137,In_650,In_318);
xor U138 (N_138,In_941,In_120);
nand U139 (N_139,In_707,In_904);
nand U140 (N_140,In_244,In_708);
and U141 (N_141,In_215,In_566);
and U142 (N_142,In_264,In_878);
or U143 (N_143,In_487,In_964);
or U144 (N_144,In_465,In_7);
or U145 (N_145,In_363,In_700);
or U146 (N_146,In_722,In_321);
and U147 (N_147,In_664,In_889);
xnor U148 (N_148,In_984,In_124);
xnor U149 (N_149,In_580,In_370);
or U150 (N_150,In_261,In_870);
nor U151 (N_151,In_437,In_864);
nand U152 (N_152,In_432,In_699);
or U153 (N_153,In_826,In_902);
nor U154 (N_154,In_934,In_676);
or U155 (N_155,In_404,In_256);
and U156 (N_156,In_270,In_32);
and U157 (N_157,In_628,In_849);
and U158 (N_158,In_939,In_597);
nand U159 (N_159,In_706,In_618);
nand U160 (N_160,In_109,In_996);
nor U161 (N_161,In_734,In_793);
or U162 (N_162,In_937,In_501);
nand U163 (N_163,In_203,In_845);
nor U164 (N_164,In_415,In_406);
nor U165 (N_165,In_41,In_317);
nand U166 (N_166,In_463,In_91);
or U167 (N_167,In_414,In_874);
xor U168 (N_168,In_248,In_712);
nor U169 (N_169,In_50,In_450);
and U170 (N_170,In_703,In_710);
xnor U171 (N_171,In_981,In_561);
nand U172 (N_172,In_27,In_947);
or U173 (N_173,In_473,In_47);
and U174 (N_174,In_288,In_895);
or U175 (N_175,In_601,In_960);
xnor U176 (N_176,In_813,In_289);
nor U177 (N_177,In_532,In_331);
nor U178 (N_178,In_528,In_377);
or U179 (N_179,In_327,In_853);
nand U180 (N_180,In_833,In_546);
or U181 (N_181,In_617,In_527);
nand U182 (N_182,In_560,In_719);
nor U183 (N_183,In_509,In_673);
nor U184 (N_184,In_497,In_492);
nor U185 (N_185,In_503,In_653);
xor U186 (N_186,In_107,In_314);
and U187 (N_187,In_976,In_956);
xor U188 (N_188,In_76,In_892);
nand U189 (N_189,In_254,In_949);
nand U190 (N_190,In_943,In_133);
and U191 (N_191,In_398,In_684);
or U192 (N_192,In_842,In_125);
nand U193 (N_193,In_379,In_721);
or U194 (N_194,In_418,In_957);
or U195 (N_195,In_307,In_808);
nand U196 (N_196,In_221,In_325);
xor U197 (N_197,In_761,In_771);
nand U198 (N_198,In_170,In_735);
nand U199 (N_199,In_604,In_88);
nand U200 (N_200,In_666,In_654);
nand U201 (N_201,In_553,In_334);
or U202 (N_202,In_101,In_649);
or U203 (N_203,In_504,In_900);
and U204 (N_204,In_452,In_49);
nand U205 (N_205,In_629,In_206);
or U206 (N_206,In_818,In_322);
or U207 (N_207,In_514,In_257);
and U208 (N_208,In_551,In_229);
and U209 (N_209,In_365,In_190);
nand U210 (N_210,In_840,In_66);
or U211 (N_211,In_646,In_679);
nand U212 (N_212,In_171,In_455);
and U213 (N_213,In_44,In_205);
or U214 (N_214,In_179,In_932);
xnor U215 (N_215,In_690,In_691);
nor U216 (N_216,In_438,In_153);
nand U217 (N_217,In_919,In_603);
nand U218 (N_218,In_905,In_583);
or U219 (N_219,In_714,In_186);
and U220 (N_220,In_637,In_290);
nand U221 (N_221,In_554,In_209);
or U222 (N_222,In_595,In_374);
and U223 (N_223,In_537,In_485);
and U224 (N_224,In_212,In_682);
or U225 (N_225,In_616,In_252);
xnor U226 (N_226,In_775,In_515);
or U227 (N_227,In_882,In_364);
and U228 (N_228,In_339,In_63);
xor U229 (N_229,In_510,In_449);
nand U230 (N_230,In_871,In_37);
nor U231 (N_231,In_499,In_407);
xnor U232 (N_232,In_336,In_718);
and U233 (N_233,In_104,In_522);
or U234 (N_234,In_2,In_610);
nor U235 (N_235,In_217,In_776);
xnor U236 (N_236,In_144,In_830);
and U237 (N_237,In_990,In_733);
and U238 (N_238,In_651,In_924);
nand U239 (N_239,In_100,In_857);
nand U240 (N_240,In_401,In_588);
nand U241 (N_241,In_81,In_615);
and U242 (N_242,In_268,In_512);
or U243 (N_243,In_114,In_239);
nor U244 (N_244,In_272,In_305);
nor U245 (N_245,In_632,In_825);
nor U246 (N_246,In_115,In_17);
nand U247 (N_247,In_168,In_894);
xnor U248 (N_248,In_783,In_787);
nor U249 (N_249,In_989,In_316);
or U250 (N_250,In_116,In_211);
nor U251 (N_251,In_814,In_977);
xnor U252 (N_252,In_410,In_887);
or U253 (N_253,In_841,In_24);
and U254 (N_254,In_683,In_959);
and U255 (N_255,In_151,In_281);
nand U256 (N_256,In_279,In_623);
or U257 (N_257,In_536,In_225);
xnor U258 (N_258,In_355,In_152);
nor U259 (N_259,In_399,In_200);
and U260 (N_260,In_59,In_611);
xnor U261 (N_261,In_69,In_255);
xor U262 (N_262,In_263,In_810);
xor U263 (N_263,In_908,In_925);
nor U264 (N_264,In_35,In_175);
nor U265 (N_265,In_498,In_451);
or U266 (N_266,In_110,In_196);
nor U267 (N_267,In_742,In_412);
nand U268 (N_268,In_42,In_278);
nand U269 (N_269,In_927,In_477);
nand U270 (N_270,In_770,In_851);
and U271 (N_271,In_692,In_106);
or U272 (N_272,In_435,In_403);
nand U273 (N_273,In_541,In_570);
nand U274 (N_274,In_763,In_208);
nand U275 (N_275,In_161,In_112);
or U276 (N_276,In_496,In_693);
nor U277 (N_277,In_579,In_122);
xor U278 (N_278,In_697,In_585);
nand U279 (N_279,In_466,In_8);
or U280 (N_280,In_30,In_963);
nor U281 (N_281,In_216,In_5);
nand U282 (N_282,In_834,In_54);
nand U283 (N_283,In_147,In_543);
or U284 (N_284,In_875,In_860);
nor U285 (N_285,In_191,In_310);
nand U286 (N_286,In_544,In_469);
or U287 (N_287,In_138,In_328);
nor U288 (N_288,In_803,In_375);
or U289 (N_289,In_409,In_181);
and U290 (N_290,In_74,In_952);
nand U291 (N_291,In_352,In_802);
and U292 (N_292,In_746,In_460);
nor U293 (N_293,In_378,In_48);
nor U294 (N_294,In_865,In_478);
nor U295 (N_295,In_798,In_668);
and U296 (N_296,In_806,In_890);
and U297 (N_297,In_576,In_581);
and U298 (N_298,In_573,In_578);
and U299 (N_299,In_777,In_250);
nand U300 (N_300,In_592,In_705);
nand U301 (N_301,In_717,In_511);
xor U302 (N_302,In_974,In_332);
nand U303 (N_303,In_145,In_677);
or U304 (N_304,In_381,In_502);
and U305 (N_305,In_914,In_420);
or U306 (N_306,In_749,In_28);
or U307 (N_307,In_523,In_607);
nor U308 (N_308,In_988,In_648);
nor U309 (N_309,In_163,In_695);
or U310 (N_310,In_308,In_490);
nand U311 (N_311,In_156,In_780);
or U312 (N_312,In_459,In_199);
nand U313 (N_313,In_481,In_987);
and U314 (N_314,In_90,In_804);
nor U315 (N_315,In_96,In_129);
nand U316 (N_316,In_390,In_817);
nand U317 (N_317,In_341,In_127);
nand U318 (N_318,In_784,In_167);
or U319 (N_319,In_367,In_567);
nand U320 (N_320,In_881,In_338);
nand U321 (N_321,In_862,In_622);
nand U322 (N_322,In_831,In_792);
and U323 (N_323,In_687,In_689);
and U324 (N_324,In_126,In_462);
nand U325 (N_325,In_111,In_855);
nand U326 (N_326,In_743,In_619);
and U327 (N_327,In_58,In_609);
and U328 (N_328,In_29,In_258);
and U329 (N_329,In_608,In_907);
or U330 (N_330,In_534,In_574);
and U331 (N_331,In_500,In_568);
nor U332 (N_332,In_659,In_928);
xor U333 (N_333,In_386,In_146);
nor U334 (N_334,In_149,In_117);
and U335 (N_335,In_829,In_613);
nor U336 (N_336,In_57,In_531);
xor U337 (N_337,In_962,In_600);
nand U338 (N_338,In_461,In_906);
nand U339 (N_339,In_304,In_103);
and U340 (N_340,In_23,In_846);
nand U341 (N_341,In_177,In_62);
nor U342 (N_342,In_440,In_773);
and U343 (N_343,In_686,In_271);
or U344 (N_344,In_39,In_15);
or U345 (N_345,In_362,In_899);
and U346 (N_346,In_231,In_296);
nor U347 (N_347,In_232,In_507);
nand U348 (N_348,In_586,In_408);
nand U349 (N_349,In_955,In_745);
nand U350 (N_350,In_980,In_267);
nor U351 (N_351,In_233,In_67);
or U352 (N_352,In_843,In_729);
and U353 (N_353,In_589,In_688);
and U354 (N_354,In_744,In_765);
nand U355 (N_355,In_542,In_174);
or U356 (N_356,In_132,In_732);
and U357 (N_357,In_727,In_446);
nand U358 (N_358,In_159,In_495);
and U359 (N_359,In_416,In_975);
nor U360 (N_360,In_417,In_9);
or U361 (N_361,In_479,In_696);
nand U362 (N_362,In_389,In_716);
and U363 (N_363,In_913,In_728);
or U364 (N_364,In_75,In_935);
nand U365 (N_365,In_226,In_18);
xor U366 (N_366,In_552,In_228);
nor U367 (N_367,In_627,In_519);
or U368 (N_368,In_781,In_471);
and U369 (N_369,In_207,In_768);
nand U370 (N_370,In_663,In_276);
or U371 (N_371,In_486,In_859);
xor U372 (N_372,In_87,In_756);
and U373 (N_373,In_474,In_630);
and U374 (N_374,In_950,In_789);
and U375 (N_375,In_369,In_794);
xnor U376 (N_376,In_197,In_392);
xor U377 (N_377,In_98,In_188);
and U378 (N_378,In_292,In_538);
and U379 (N_379,In_158,In_342);
xnor U380 (N_380,In_413,In_713);
or U381 (N_381,In_454,In_702);
and U382 (N_382,In_774,In_850);
nor U383 (N_383,In_971,In_533);
and U384 (N_384,In_494,In_249);
nand U385 (N_385,In_820,In_624);
nand U386 (N_386,In_520,In_204);
nand U387 (N_387,In_866,In_491);
nand U388 (N_388,In_269,In_436);
nor U389 (N_389,In_344,In_973);
and U390 (N_390,In_602,In_287);
or U391 (N_391,In_237,In_93);
and U392 (N_392,In_726,In_434);
nor U393 (N_393,In_458,In_493);
nor U394 (N_394,In_286,In_172);
nand U395 (N_395,In_967,In_769);
nand U396 (N_396,In_750,In_662);
nand U397 (N_397,In_131,In_128);
nand U398 (N_398,In_764,In_641);
nor U399 (N_399,In_285,In_869);
and U400 (N_400,In_724,In_631);
nand U401 (N_401,In_669,In_210);
or U402 (N_402,In_819,In_84);
nand U403 (N_403,In_80,In_917);
and U404 (N_404,In_751,In_467);
nor U405 (N_405,In_247,In_506);
xor U406 (N_406,In_916,In_605);
nor U407 (N_407,In_569,In_64);
and U408 (N_408,In_828,In_656);
nor U409 (N_409,In_148,In_108);
nor U410 (N_410,In_260,In_685);
or U411 (N_411,In_674,In_915);
or U412 (N_412,In_397,In_273);
and U413 (N_413,In_251,In_4);
or U414 (N_414,In_135,In_297);
xor U415 (N_415,In_274,In_795);
and U416 (N_416,In_348,In_422);
nand U417 (N_417,In_22,In_16);
nand U418 (N_418,In_277,In_448);
or U419 (N_419,In_762,In_953);
xnor U420 (N_420,In_445,In_245);
nor U421 (N_421,In_991,In_753);
and U422 (N_422,In_680,In_741);
xor U423 (N_423,In_513,In_72);
nor U424 (N_424,In_931,In_383);
and U425 (N_425,In_464,In_748);
nor U426 (N_426,In_782,In_358);
xor U427 (N_427,In_636,In_740);
nand U428 (N_428,In_118,In_77);
xnor U429 (N_429,In_142,In_638);
nor U430 (N_430,In_807,In_426);
nor U431 (N_431,In_357,In_319);
and U432 (N_432,In_3,In_678);
nor U433 (N_433,In_736,In_525);
and U434 (N_434,In_715,In_326);
nand U435 (N_435,In_213,In_354);
or U436 (N_436,In_535,In_888);
nand U437 (N_437,In_593,In_102);
nand U438 (N_438,In_189,In_198);
or U439 (N_439,In_315,In_94);
or U440 (N_440,In_997,In_238);
xnor U441 (N_441,In_371,In_482);
nand U442 (N_442,In_185,In_178);
or U443 (N_443,In_359,In_52);
xor U444 (N_444,In_655,In_182);
nor U445 (N_445,In_201,In_639);
nor U446 (N_446,In_333,In_885);
and U447 (N_447,In_6,In_475);
nor U448 (N_448,In_993,In_867);
and U449 (N_449,In_423,In_119);
or U450 (N_450,In_45,In_162);
nand U451 (N_451,In_832,In_590);
nand U452 (N_452,In_150,In_143);
or U453 (N_453,In_457,In_539);
or U454 (N_454,In_70,In_202);
nand U455 (N_455,In_447,In_155);
xnor U456 (N_456,In_236,In_246);
or U457 (N_457,In_262,In_139);
nand U458 (N_458,In_193,In_320);
nand U459 (N_459,In_985,In_241);
and U460 (N_460,In_797,In_872);
and U461 (N_461,In_698,In_758);
nand U462 (N_462,In_38,In_675);
nand U463 (N_463,In_488,In_259);
or U464 (N_464,In_811,In_380);
and U465 (N_465,In_20,In_235);
or U466 (N_466,In_951,In_68);
nand U467 (N_467,In_918,In_823);
xor U468 (N_468,In_582,In_335);
and U469 (N_469,In_160,In_933);
and U470 (N_470,In_873,In_214);
nor U471 (N_471,In_958,In_295);
or U472 (N_472,In_559,In_360);
nand U473 (N_473,In_361,In_921);
nand U474 (N_474,In_79,In_176);
and U475 (N_475,In_323,In_40);
nand U476 (N_476,In_923,In_21);
xnor U477 (N_477,In_671,In_672);
or U478 (N_478,In_388,In_550);
nand U479 (N_479,In_428,In_530);
nor U480 (N_480,In_184,In_785);
nand U481 (N_481,In_43,In_303);
and U482 (N_482,In_329,In_970);
nand U483 (N_483,In_877,In_800);
nand U484 (N_484,In_565,In_85);
nor U485 (N_485,In_430,In_73);
or U486 (N_486,In_801,In_824);
and U487 (N_487,In_424,In_940);
nor U488 (N_488,In_720,In_140);
and U489 (N_489,In_665,In_844);
or U490 (N_490,In_936,In_483);
nor U491 (N_491,In_61,In_752);
nor U492 (N_492,In_518,In_113);
and U493 (N_493,In_557,In_858);
nor U494 (N_494,In_839,In_376);
nor U495 (N_495,In_948,In_243);
or U496 (N_496,In_547,In_516);
nand U497 (N_497,In_896,In_242);
and U498 (N_498,In_661,In_137);
or U499 (N_499,In_835,In_772);
nand U500 (N_500,In_887,In_281);
nor U501 (N_501,In_97,In_764);
and U502 (N_502,In_468,In_467);
or U503 (N_503,In_483,In_670);
nor U504 (N_504,In_199,In_802);
nand U505 (N_505,In_119,In_933);
nor U506 (N_506,In_243,In_337);
and U507 (N_507,In_250,In_377);
nor U508 (N_508,In_755,In_983);
or U509 (N_509,In_566,In_461);
nand U510 (N_510,In_359,In_146);
nand U511 (N_511,In_452,In_15);
nand U512 (N_512,In_528,In_850);
or U513 (N_513,In_345,In_264);
nor U514 (N_514,In_305,In_523);
nand U515 (N_515,In_607,In_744);
nand U516 (N_516,In_478,In_534);
or U517 (N_517,In_60,In_756);
xnor U518 (N_518,In_680,In_325);
and U519 (N_519,In_329,In_352);
or U520 (N_520,In_513,In_179);
and U521 (N_521,In_682,In_581);
or U522 (N_522,In_293,In_859);
nor U523 (N_523,In_13,In_912);
nand U524 (N_524,In_250,In_6);
nor U525 (N_525,In_703,In_514);
or U526 (N_526,In_873,In_255);
nor U527 (N_527,In_220,In_686);
or U528 (N_528,In_377,In_242);
nor U529 (N_529,In_607,In_761);
nor U530 (N_530,In_538,In_210);
or U531 (N_531,In_374,In_792);
nand U532 (N_532,In_308,In_357);
and U533 (N_533,In_452,In_524);
nand U534 (N_534,In_811,In_94);
or U535 (N_535,In_536,In_849);
xor U536 (N_536,In_181,In_815);
or U537 (N_537,In_698,In_379);
nor U538 (N_538,In_718,In_719);
nand U539 (N_539,In_288,In_943);
or U540 (N_540,In_685,In_813);
and U541 (N_541,In_541,In_360);
and U542 (N_542,In_583,In_401);
nor U543 (N_543,In_315,In_999);
nor U544 (N_544,In_758,In_993);
and U545 (N_545,In_861,In_9);
nand U546 (N_546,In_86,In_339);
and U547 (N_547,In_306,In_326);
or U548 (N_548,In_117,In_373);
or U549 (N_549,In_563,In_664);
or U550 (N_550,In_880,In_598);
and U551 (N_551,In_824,In_232);
or U552 (N_552,In_796,In_984);
and U553 (N_553,In_554,In_319);
nor U554 (N_554,In_54,In_303);
and U555 (N_555,In_569,In_76);
nand U556 (N_556,In_985,In_299);
xor U557 (N_557,In_706,In_829);
xnor U558 (N_558,In_400,In_702);
nor U559 (N_559,In_123,In_75);
and U560 (N_560,In_992,In_577);
or U561 (N_561,In_592,In_908);
nand U562 (N_562,In_73,In_150);
and U563 (N_563,In_478,In_916);
and U564 (N_564,In_804,In_114);
nor U565 (N_565,In_477,In_180);
or U566 (N_566,In_628,In_799);
and U567 (N_567,In_797,In_353);
nand U568 (N_568,In_770,In_897);
or U569 (N_569,In_746,In_133);
or U570 (N_570,In_901,In_35);
nor U571 (N_571,In_586,In_663);
or U572 (N_572,In_731,In_949);
nor U573 (N_573,In_669,In_508);
or U574 (N_574,In_965,In_564);
and U575 (N_575,In_115,In_448);
and U576 (N_576,In_839,In_938);
nand U577 (N_577,In_6,In_14);
and U578 (N_578,In_896,In_992);
xnor U579 (N_579,In_685,In_930);
xor U580 (N_580,In_223,In_968);
nor U581 (N_581,In_137,In_622);
nand U582 (N_582,In_360,In_480);
nor U583 (N_583,In_456,In_207);
nor U584 (N_584,In_50,In_771);
nor U585 (N_585,In_919,In_639);
and U586 (N_586,In_581,In_934);
and U587 (N_587,In_69,In_870);
nand U588 (N_588,In_772,In_78);
nand U589 (N_589,In_141,In_806);
and U590 (N_590,In_616,In_471);
or U591 (N_591,In_172,In_215);
or U592 (N_592,In_773,In_270);
or U593 (N_593,In_390,In_120);
or U594 (N_594,In_897,In_774);
and U595 (N_595,In_23,In_839);
nand U596 (N_596,In_902,In_74);
nor U597 (N_597,In_897,In_204);
and U598 (N_598,In_601,In_968);
xnor U599 (N_599,In_377,In_129);
xor U600 (N_600,In_124,In_559);
and U601 (N_601,In_209,In_488);
nand U602 (N_602,In_75,In_0);
or U603 (N_603,In_801,In_277);
and U604 (N_604,In_429,In_64);
nor U605 (N_605,In_112,In_666);
xnor U606 (N_606,In_398,In_193);
and U607 (N_607,In_219,In_566);
xor U608 (N_608,In_726,In_737);
nor U609 (N_609,In_603,In_834);
xor U610 (N_610,In_845,In_664);
nor U611 (N_611,In_622,In_393);
nand U612 (N_612,In_16,In_607);
nor U613 (N_613,In_611,In_803);
nor U614 (N_614,In_162,In_215);
nor U615 (N_615,In_232,In_944);
nand U616 (N_616,In_283,In_881);
nand U617 (N_617,In_161,In_587);
and U618 (N_618,In_303,In_632);
nand U619 (N_619,In_921,In_293);
or U620 (N_620,In_673,In_115);
or U621 (N_621,In_558,In_769);
or U622 (N_622,In_963,In_459);
and U623 (N_623,In_456,In_298);
nand U624 (N_624,In_959,In_807);
and U625 (N_625,In_506,In_543);
nor U626 (N_626,In_520,In_119);
and U627 (N_627,In_982,In_800);
and U628 (N_628,In_390,In_613);
and U629 (N_629,In_351,In_182);
or U630 (N_630,In_819,In_293);
nor U631 (N_631,In_309,In_549);
nand U632 (N_632,In_258,In_177);
nand U633 (N_633,In_794,In_901);
and U634 (N_634,In_495,In_639);
and U635 (N_635,In_100,In_388);
or U636 (N_636,In_447,In_173);
nand U637 (N_637,In_905,In_787);
xnor U638 (N_638,In_147,In_814);
xor U639 (N_639,In_614,In_324);
or U640 (N_640,In_852,In_257);
and U641 (N_641,In_195,In_909);
nand U642 (N_642,In_563,In_297);
or U643 (N_643,In_632,In_228);
nand U644 (N_644,In_757,In_17);
and U645 (N_645,In_166,In_153);
and U646 (N_646,In_400,In_374);
nor U647 (N_647,In_844,In_975);
or U648 (N_648,In_721,In_269);
xnor U649 (N_649,In_898,In_896);
or U650 (N_650,In_667,In_529);
xnor U651 (N_651,In_976,In_483);
xor U652 (N_652,In_678,In_624);
and U653 (N_653,In_443,In_835);
nor U654 (N_654,In_22,In_686);
nor U655 (N_655,In_764,In_402);
or U656 (N_656,In_459,In_394);
nand U657 (N_657,In_579,In_533);
or U658 (N_658,In_20,In_370);
xor U659 (N_659,In_804,In_346);
nor U660 (N_660,In_738,In_674);
nor U661 (N_661,In_323,In_554);
nand U662 (N_662,In_793,In_918);
nand U663 (N_663,In_618,In_222);
or U664 (N_664,In_993,In_289);
nor U665 (N_665,In_619,In_735);
or U666 (N_666,In_856,In_541);
nor U667 (N_667,In_756,In_921);
nor U668 (N_668,In_68,In_380);
nor U669 (N_669,In_123,In_700);
and U670 (N_670,In_691,In_553);
and U671 (N_671,In_611,In_889);
nor U672 (N_672,In_327,In_370);
xor U673 (N_673,In_361,In_901);
nand U674 (N_674,In_347,In_946);
nor U675 (N_675,In_902,In_265);
nor U676 (N_676,In_740,In_470);
nor U677 (N_677,In_10,In_533);
or U678 (N_678,In_215,In_774);
nand U679 (N_679,In_240,In_173);
nand U680 (N_680,In_517,In_870);
and U681 (N_681,In_461,In_544);
nand U682 (N_682,In_598,In_242);
nand U683 (N_683,In_103,In_837);
or U684 (N_684,In_666,In_378);
and U685 (N_685,In_218,In_690);
xor U686 (N_686,In_563,In_772);
or U687 (N_687,In_608,In_260);
nand U688 (N_688,In_726,In_952);
and U689 (N_689,In_493,In_911);
or U690 (N_690,In_691,In_359);
or U691 (N_691,In_758,In_345);
nor U692 (N_692,In_652,In_327);
xor U693 (N_693,In_907,In_485);
xor U694 (N_694,In_31,In_151);
or U695 (N_695,In_2,In_382);
nand U696 (N_696,In_76,In_419);
nor U697 (N_697,In_108,In_279);
nand U698 (N_698,In_675,In_817);
and U699 (N_699,In_428,In_743);
nor U700 (N_700,In_984,In_205);
nand U701 (N_701,In_652,In_971);
nand U702 (N_702,In_116,In_790);
or U703 (N_703,In_95,In_144);
nand U704 (N_704,In_181,In_913);
xor U705 (N_705,In_927,In_158);
nand U706 (N_706,In_466,In_548);
nand U707 (N_707,In_454,In_934);
nor U708 (N_708,In_123,In_789);
or U709 (N_709,In_415,In_150);
or U710 (N_710,In_219,In_386);
nor U711 (N_711,In_552,In_847);
nand U712 (N_712,In_252,In_349);
nand U713 (N_713,In_955,In_17);
nand U714 (N_714,In_892,In_731);
nand U715 (N_715,In_26,In_29);
or U716 (N_716,In_317,In_237);
nand U717 (N_717,In_357,In_957);
nor U718 (N_718,In_455,In_562);
and U719 (N_719,In_70,In_654);
or U720 (N_720,In_131,In_516);
xor U721 (N_721,In_375,In_141);
and U722 (N_722,In_438,In_770);
and U723 (N_723,In_913,In_733);
nand U724 (N_724,In_209,In_72);
and U725 (N_725,In_901,In_700);
or U726 (N_726,In_313,In_110);
nand U727 (N_727,In_949,In_921);
or U728 (N_728,In_251,In_705);
nand U729 (N_729,In_241,In_939);
nor U730 (N_730,In_95,In_913);
nand U731 (N_731,In_158,In_130);
xnor U732 (N_732,In_620,In_918);
or U733 (N_733,In_983,In_731);
xnor U734 (N_734,In_108,In_869);
or U735 (N_735,In_12,In_391);
and U736 (N_736,In_472,In_249);
nand U737 (N_737,In_832,In_189);
or U738 (N_738,In_883,In_476);
nand U739 (N_739,In_899,In_749);
nor U740 (N_740,In_91,In_328);
xnor U741 (N_741,In_630,In_350);
and U742 (N_742,In_946,In_643);
xor U743 (N_743,In_408,In_685);
nand U744 (N_744,In_45,In_375);
nand U745 (N_745,In_934,In_217);
nand U746 (N_746,In_238,In_585);
or U747 (N_747,In_892,In_836);
nand U748 (N_748,In_547,In_109);
and U749 (N_749,In_76,In_916);
nand U750 (N_750,In_866,In_684);
nand U751 (N_751,In_303,In_326);
nand U752 (N_752,In_71,In_345);
xor U753 (N_753,In_416,In_642);
or U754 (N_754,In_936,In_693);
and U755 (N_755,In_410,In_955);
nor U756 (N_756,In_391,In_258);
or U757 (N_757,In_526,In_648);
or U758 (N_758,In_569,In_237);
or U759 (N_759,In_465,In_938);
and U760 (N_760,In_971,In_474);
xor U761 (N_761,In_843,In_49);
nor U762 (N_762,In_719,In_170);
nor U763 (N_763,In_902,In_459);
or U764 (N_764,In_67,In_563);
nand U765 (N_765,In_493,In_867);
nand U766 (N_766,In_224,In_598);
xor U767 (N_767,In_680,In_701);
or U768 (N_768,In_109,In_437);
xnor U769 (N_769,In_327,In_500);
nor U770 (N_770,In_798,In_787);
nand U771 (N_771,In_830,In_994);
and U772 (N_772,In_437,In_972);
and U773 (N_773,In_794,In_921);
and U774 (N_774,In_690,In_881);
and U775 (N_775,In_466,In_47);
xnor U776 (N_776,In_381,In_670);
nor U777 (N_777,In_77,In_751);
or U778 (N_778,In_720,In_84);
and U779 (N_779,In_658,In_402);
and U780 (N_780,In_900,In_155);
and U781 (N_781,In_497,In_307);
nand U782 (N_782,In_550,In_179);
nand U783 (N_783,In_583,In_443);
or U784 (N_784,In_308,In_39);
nand U785 (N_785,In_175,In_530);
xor U786 (N_786,In_226,In_627);
and U787 (N_787,In_903,In_445);
and U788 (N_788,In_116,In_284);
and U789 (N_789,In_921,In_790);
and U790 (N_790,In_854,In_827);
nand U791 (N_791,In_646,In_733);
nor U792 (N_792,In_201,In_8);
or U793 (N_793,In_718,In_949);
and U794 (N_794,In_277,In_479);
nand U795 (N_795,In_182,In_742);
nand U796 (N_796,In_696,In_564);
nor U797 (N_797,In_664,In_923);
nor U798 (N_798,In_543,In_841);
or U799 (N_799,In_444,In_107);
or U800 (N_800,In_467,In_907);
nor U801 (N_801,In_183,In_904);
nand U802 (N_802,In_984,In_758);
nor U803 (N_803,In_999,In_949);
and U804 (N_804,In_660,In_418);
and U805 (N_805,In_256,In_917);
nand U806 (N_806,In_274,In_472);
or U807 (N_807,In_118,In_40);
nor U808 (N_808,In_541,In_527);
nand U809 (N_809,In_759,In_219);
and U810 (N_810,In_714,In_879);
nand U811 (N_811,In_415,In_167);
xor U812 (N_812,In_556,In_288);
nor U813 (N_813,In_648,In_571);
and U814 (N_814,In_82,In_387);
and U815 (N_815,In_438,In_103);
and U816 (N_816,In_263,In_251);
nand U817 (N_817,In_97,In_752);
nand U818 (N_818,In_72,In_600);
and U819 (N_819,In_565,In_343);
and U820 (N_820,In_569,In_345);
or U821 (N_821,In_154,In_751);
nand U822 (N_822,In_306,In_301);
nor U823 (N_823,In_393,In_588);
nor U824 (N_824,In_128,In_314);
nor U825 (N_825,In_688,In_649);
nor U826 (N_826,In_187,In_318);
or U827 (N_827,In_349,In_302);
xor U828 (N_828,In_190,In_200);
nor U829 (N_829,In_829,In_843);
nor U830 (N_830,In_834,In_84);
and U831 (N_831,In_617,In_464);
and U832 (N_832,In_979,In_81);
or U833 (N_833,In_300,In_976);
nand U834 (N_834,In_506,In_558);
and U835 (N_835,In_884,In_822);
or U836 (N_836,In_572,In_876);
nand U837 (N_837,In_445,In_298);
or U838 (N_838,In_523,In_672);
and U839 (N_839,In_181,In_840);
xnor U840 (N_840,In_701,In_53);
nor U841 (N_841,In_792,In_128);
xor U842 (N_842,In_474,In_594);
or U843 (N_843,In_681,In_151);
or U844 (N_844,In_752,In_365);
nand U845 (N_845,In_930,In_330);
nor U846 (N_846,In_356,In_678);
nand U847 (N_847,In_899,In_694);
nor U848 (N_848,In_25,In_290);
nor U849 (N_849,In_562,In_561);
and U850 (N_850,In_435,In_181);
or U851 (N_851,In_738,In_774);
or U852 (N_852,In_355,In_584);
nor U853 (N_853,In_64,In_484);
xor U854 (N_854,In_362,In_925);
or U855 (N_855,In_709,In_248);
nor U856 (N_856,In_32,In_372);
nand U857 (N_857,In_70,In_201);
nand U858 (N_858,In_66,In_136);
nand U859 (N_859,In_684,In_557);
and U860 (N_860,In_902,In_932);
nand U861 (N_861,In_775,In_39);
or U862 (N_862,In_967,In_850);
xnor U863 (N_863,In_514,In_827);
nand U864 (N_864,In_864,In_354);
and U865 (N_865,In_965,In_628);
or U866 (N_866,In_627,In_97);
nand U867 (N_867,In_989,In_437);
nor U868 (N_868,In_600,In_693);
nor U869 (N_869,In_552,In_514);
nor U870 (N_870,In_77,In_603);
or U871 (N_871,In_272,In_135);
or U872 (N_872,In_261,In_162);
nor U873 (N_873,In_853,In_905);
nand U874 (N_874,In_988,In_382);
nor U875 (N_875,In_178,In_341);
xor U876 (N_876,In_390,In_923);
nor U877 (N_877,In_854,In_196);
or U878 (N_878,In_890,In_814);
nand U879 (N_879,In_672,In_99);
nand U880 (N_880,In_794,In_117);
nand U881 (N_881,In_358,In_734);
nor U882 (N_882,In_989,In_532);
and U883 (N_883,In_927,In_425);
nand U884 (N_884,In_133,In_236);
and U885 (N_885,In_750,In_243);
or U886 (N_886,In_247,In_427);
nand U887 (N_887,In_715,In_705);
nor U888 (N_888,In_818,In_67);
nand U889 (N_889,In_45,In_589);
nand U890 (N_890,In_286,In_529);
xor U891 (N_891,In_54,In_783);
or U892 (N_892,In_404,In_269);
nand U893 (N_893,In_372,In_316);
nand U894 (N_894,In_879,In_14);
and U895 (N_895,In_12,In_162);
nor U896 (N_896,In_326,In_101);
xnor U897 (N_897,In_923,In_304);
and U898 (N_898,In_614,In_736);
nand U899 (N_899,In_777,In_869);
nand U900 (N_900,In_458,In_308);
and U901 (N_901,In_841,In_399);
and U902 (N_902,In_407,In_759);
or U903 (N_903,In_874,In_908);
or U904 (N_904,In_111,In_754);
nor U905 (N_905,In_625,In_943);
and U906 (N_906,In_493,In_616);
or U907 (N_907,In_477,In_320);
nand U908 (N_908,In_209,In_75);
nand U909 (N_909,In_150,In_220);
nor U910 (N_910,In_439,In_125);
nor U911 (N_911,In_810,In_596);
nand U912 (N_912,In_608,In_475);
nand U913 (N_913,In_312,In_128);
and U914 (N_914,In_296,In_770);
nor U915 (N_915,In_897,In_941);
nand U916 (N_916,In_852,In_461);
or U917 (N_917,In_982,In_883);
nor U918 (N_918,In_597,In_747);
and U919 (N_919,In_409,In_647);
and U920 (N_920,In_776,In_249);
xor U921 (N_921,In_751,In_659);
and U922 (N_922,In_731,In_91);
xor U923 (N_923,In_586,In_204);
or U924 (N_924,In_111,In_511);
and U925 (N_925,In_80,In_984);
nand U926 (N_926,In_89,In_562);
and U927 (N_927,In_791,In_240);
and U928 (N_928,In_493,In_886);
nor U929 (N_929,In_670,In_361);
nand U930 (N_930,In_658,In_568);
xor U931 (N_931,In_626,In_394);
nor U932 (N_932,In_896,In_191);
xnor U933 (N_933,In_676,In_608);
nor U934 (N_934,In_241,In_853);
nor U935 (N_935,In_840,In_653);
xor U936 (N_936,In_972,In_82);
nand U937 (N_937,In_882,In_885);
nand U938 (N_938,In_895,In_517);
and U939 (N_939,In_271,In_471);
nand U940 (N_940,In_389,In_736);
nand U941 (N_941,In_87,In_932);
nor U942 (N_942,In_962,In_75);
or U943 (N_943,In_366,In_813);
and U944 (N_944,In_488,In_366);
nand U945 (N_945,In_281,In_226);
or U946 (N_946,In_56,In_609);
and U947 (N_947,In_441,In_916);
xnor U948 (N_948,In_433,In_507);
or U949 (N_949,In_410,In_386);
nor U950 (N_950,In_85,In_50);
or U951 (N_951,In_195,In_46);
xor U952 (N_952,In_382,In_766);
and U953 (N_953,In_99,In_112);
nand U954 (N_954,In_131,In_692);
and U955 (N_955,In_587,In_421);
and U956 (N_956,In_105,In_952);
xnor U957 (N_957,In_313,In_427);
and U958 (N_958,In_105,In_4);
nand U959 (N_959,In_536,In_751);
nand U960 (N_960,In_249,In_252);
and U961 (N_961,In_763,In_880);
and U962 (N_962,In_949,In_768);
nand U963 (N_963,In_867,In_815);
nor U964 (N_964,In_764,In_184);
and U965 (N_965,In_73,In_493);
nand U966 (N_966,In_457,In_259);
and U967 (N_967,In_367,In_947);
nor U968 (N_968,In_634,In_4);
or U969 (N_969,In_257,In_206);
and U970 (N_970,In_983,In_94);
and U971 (N_971,In_525,In_270);
nor U972 (N_972,In_806,In_687);
xnor U973 (N_973,In_565,In_974);
nor U974 (N_974,In_814,In_804);
and U975 (N_975,In_993,In_35);
nand U976 (N_976,In_288,In_771);
nor U977 (N_977,In_819,In_851);
nand U978 (N_978,In_800,In_935);
nor U979 (N_979,In_989,In_911);
nor U980 (N_980,In_19,In_448);
nand U981 (N_981,In_438,In_710);
nor U982 (N_982,In_964,In_346);
and U983 (N_983,In_854,In_142);
or U984 (N_984,In_230,In_183);
and U985 (N_985,In_716,In_113);
nand U986 (N_986,In_622,In_799);
nor U987 (N_987,In_254,In_209);
xnor U988 (N_988,In_362,In_600);
and U989 (N_989,In_105,In_655);
nor U990 (N_990,In_707,In_199);
nor U991 (N_991,In_299,In_251);
and U992 (N_992,In_804,In_718);
nand U993 (N_993,In_326,In_829);
nand U994 (N_994,In_339,In_428);
or U995 (N_995,In_677,In_844);
and U996 (N_996,In_141,In_843);
or U997 (N_997,In_338,In_88);
and U998 (N_998,In_525,In_296);
or U999 (N_999,In_424,In_802);
or U1000 (N_1000,In_669,In_524);
nor U1001 (N_1001,In_223,In_633);
and U1002 (N_1002,In_191,In_642);
or U1003 (N_1003,In_796,In_356);
or U1004 (N_1004,In_789,In_531);
or U1005 (N_1005,In_963,In_81);
or U1006 (N_1006,In_492,In_46);
or U1007 (N_1007,In_383,In_893);
or U1008 (N_1008,In_878,In_290);
xor U1009 (N_1009,In_35,In_826);
nor U1010 (N_1010,In_600,In_819);
or U1011 (N_1011,In_432,In_158);
nand U1012 (N_1012,In_865,In_247);
or U1013 (N_1013,In_487,In_914);
or U1014 (N_1014,In_992,In_681);
and U1015 (N_1015,In_744,In_999);
and U1016 (N_1016,In_664,In_934);
or U1017 (N_1017,In_12,In_889);
nor U1018 (N_1018,In_116,In_372);
and U1019 (N_1019,In_211,In_761);
and U1020 (N_1020,In_947,In_306);
and U1021 (N_1021,In_925,In_528);
or U1022 (N_1022,In_721,In_258);
xnor U1023 (N_1023,In_65,In_675);
or U1024 (N_1024,In_2,In_955);
and U1025 (N_1025,In_621,In_71);
nor U1026 (N_1026,In_452,In_789);
nand U1027 (N_1027,In_91,In_660);
and U1028 (N_1028,In_437,In_658);
nor U1029 (N_1029,In_307,In_982);
nand U1030 (N_1030,In_48,In_521);
xnor U1031 (N_1031,In_72,In_454);
or U1032 (N_1032,In_694,In_936);
or U1033 (N_1033,In_887,In_976);
nand U1034 (N_1034,In_396,In_15);
and U1035 (N_1035,In_241,In_406);
or U1036 (N_1036,In_827,In_935);
nor U1037 (N_1037,In_436,In_740);
nand U1038 (N_1038,In_186,In_63);
nand U1039 (N_1039,In_134,In_367);
nand U1040 (N_1040,In_717,In_10);
xor U1041 (N_1041,In_26,In_862);
nor U1042 (N_1042,In_30,In_651);
nand U1043 (N_1043,In_6,In_885);
nand U1044 (N_1044,In_699,In_911);
or U1045 (N_1045,In_959,In_366);
nor U1046 (N_1046,In_232,In_657);
nor U1047 (N_1047,In_164,In_653);
or U1048 (N_1048,In_33,In_161);
nand U1049 (N_1049,In_425,In_159);
and U1050 (N_1050,In_226,In_540);
nor U1051 (N_1051,In_116,In_34);
nand U1052 (N_1052,In_873,In_332);
nor U1053 (N_1053,In_174,In_979);
nor U1054 (N_1054,In_329,In_935);
xor U1055 (N_1055,In_929,In_295);
nor U1056 (N_1056,In_416,In_6);
or U1057 (N_1057,In_202,In_8);
or U1058 (N_1058,In_720,In_352);
xnor U1059 (N_1059,In_525,In_934);
xor U1060 (N_1060,In_602,In_982);
and U1061 (N_1061,In_560,In_499);
or U1062 (N_1062,In_855,In_533);
nor U1063 (N_1063,In_305,In_464);
nor U1064 (N_1064,In_910,In_801);
nand U1065 (N_1065,In_919,In_298);
or U1066 (N_1066,In_785,In_164);
nor U1067 (N_1067,In_249,In_372);
nand U1068 (N_1068,In_970,In_79);
nor U1069 (N_1069,In_526,In_418);
nor U1070 (N_1070,In_894,In_661);
xor U1071 (N_1071,In_883,In_616);
nor U1072 (N_1072,In_915,In_810);
or U1073 (N_1073,In_432,In_632);
or U1074 (N_1074,In_587,In_81);
and U1075 (N_1075,In_312,In_750);
or U1076 (N_1076,In_480,In_558);
or U1077 (N_1077,In_859,In_223);
nand U1078 (N_1078,In_537,In_602);
nor U1079 (N_1079,In_88,In_328);
nand U1080 (N_1080,In_904,In_359);
nor U1081 (N_1081,In_937,In_73);
and U1082 (N_1082,In_170,In_301);
nand U1083 (N_1083,In_423,In_685);
nor U1084 (N_1084,In_188,In_40);
and U1085 (N_1085,In_437,In_331);
nand U1086 (N_1086,In_387,In_642);
nand U1087 (N_1087,In_25,In_123);
xnor U1088 (N_1088,In_357,In_182);
and U1089 (N_1089,In_620,In_192);
and U1090 (N_1090,In_999,In_125);
nand U1091 (N_1091,In_654,In_252);
nor U1092 (N_1092,In_87,In_869);
nand U1093 (N_1093,In_419,In_404);
nand U1094 (N_1094,In_185,In_602);
nor U1095 (N_1095,In_387,In_829);
nand U1096 (N_1096,In_699,In_380);
xor U1097 (N_1097,In_140,In_319);
and U1098 (N_1098,In_792,In_582);
xnor U1099 (N_1099,In_523,In_345);
nor U1100 (N_1100,In_829,In_688);
or U1101 (N_1101,In_40,In_144);
nand U1102 (N_1102,In_453,In_398);
xnor U1103 (N_1103,In_704,In_595);
nor U1104 (N_1104,In_925,In_856);
nand U1105 (N_1105,In_318,In_655);
nor U1106 (N_1106,In_657,In_715);
or U1107 (N_1107,In_50,In_974);
nor U1108 (N_1108,In_94,In_362);
nand U1109 (N_1109,In_981,In_551);
nand U1110 (N_1110,In_240,In_419);
nor U1111 (N_1111,In_613,In_223);
and U1112 (N_1112,In_88,In_839);
and U1113 (N_1113,In_736,In_832);
or U1114 (N_1114,In_900,In_973);
and U1115 (N_1115,In_337,In_946);
or U1116 (N_1116,In_933,In_193);
nand U1117 (N_1117,In_191,In_433);
nand U1118 (N_1118,In_293,In_415);
nor U1119 (N_1119,In_788,In_233);
and U1120 (N_1120,In_786,In_818);
nor U1121 (N_1121,In_601,In_817);
xor U1122 (N_1122,In_889,In_754);
xnor U1123 (N_1123,In_978,In_917);
and U1124 (N_1124,In_963,In_757);
and U1125 (N_1125,In_86,In_819);
nand U1126 (N_1126,In_202,In_113);
nor U1127 (N_1127,In_770,In_510);
nand U1128 (N_1128,In_851,In_195);
nand U1129 (N_1129,In_738,In_936);
nor U1130 (N_1130,In_196,In_861);
or U1131 (N_1131,In_732,In_460);
nand U1132 (N_1132,In_418,In_829);
nor U1133 (N_1133,In_348,In_478);
nand U1134 (N_1134,In_12,In_778);
and U1135 (N_1135,In_99,In_961);
or U1136 (N_1136,In_874,In_29);
nand U1137 (N_1137,In_898,In_21);
or U1138 (N_1138,In_285,In_966);
or U1139 (N_1139,In_280,In_47);
or U1140 (N_1140,In_449,In_796);
nor U1141 (N_1141,In_87,In_648);
or U1142 (N_1142,In_490,In_599);
or U1143 (N_1143,In_39,In_958);
or U1144 (N_1144,In_875,In_611);
or U1145 (N_1145,In_86,In_104);
or U1146 (N_1146,In_185,In_225);
and U1147 (N_1147,In_925,In_23);
xor U1148 (N_1148,In_334,In_885);
and U1149 (N_1149,In_391,In_711);
and U1150 (N_1150,In_23,In_318);
and U1151 (N_1151,In_521,In_71);
nor U1152 (N_1152,In_391,In_752);
nand U1153 (N_1153,In_621,In_360);
xor U1154 (N_1154,In_49,In_507);
nand U1155 (N_1155,In_872,In_652);
xnor U1156 (N_1156,In_250,In_709);
xor U1157 (N_1157,In_745,In_258);
and U1158 (N_1158,In_368,In_117);
or U1159 (N_1159,In_720,In_758);
nor U1160 (N_1160,In_533,In_378);
and U1161 (N_1161,In_434,In_703);
xor U1162 (N_1162,In_425,In_387);
nand U1163 (N_1163,In_974,In_324);
or U1164 (N_1164,In_553,In_607);
and U1165 (N_1165,In_989,In_47);
or U1166 (N_1166,In_281,In_852);
nand U1167 (N_1167,In_154,In_45);
and U1168 (N_1168,In_814,In_323);
or U1169 (N_1169,In_887,In_394);
and U1170 (N_1170,In_151,In_237);
xor U1171 (N_1171,In_900,In_272);
nor U1172 (N_1172,In_706,In_687);
and U1173 (N_1173,In_776,In_644);
nor U1174 (N_1174,In_127,In_776);
nand U1175 (N_1175,In_509,In_319);
nor U1176 (N_1176,In_593,In_732);
and U1177 (N_1177,In_161,In_811);
and U1178 (N_1178,In_415,In_189);
or U1179 (N_1179,In_924,In_647);
nand U1180 (N_1180,In_505,In_862);
nor U1181 (N_1181,In_674,In_679);
and U1182 (N_1182,In_890,In_766);
or U1183 (N_1183,In_833,In_75);
and U1184 (N_1184,In_13,In_486);
nand U1185 (N_1185,In_261,In_586);
or U1186 (N_1186,In_530,In_374);
nor U1187 (N_1187,In_843,In_16);
nand U1188 (N_1188,In_958,In_647);
or U1189 (N_1189,In_355,In_941);
nor U1190 (N_1190,In_436,In_90);
nand U1191 (N_1191,In_316,In_330);
nor U1192 (N_1192,In_17,In_540);
xnor U1193 (N_1193,In_443,In_904);
and U1194 (N_1194,In_167,In_62);
nand U1195 (N_1195,In_637,In_323);
nor U1196 (N_1196,In_873,In_83);
and U1197 (N_1197,In_412,In_522);
or U1198 (N_1198,In_5,In_772);
and U1199 (N_1199,In_691,In_71);
and U1200 (N_1200,In_915,In_218);
nor U1201 (N_1201,In_32,In_473);
and U1202 (N_1202,In_256,In_441);
and U1203 (N_1203,In_838,In_207);
nor U1204 (N_1204,In_476,In_863);
and U1205 (N_1205,In_79,In_195);
nor U1206 (N_1206,In_33,In_857);
nand U1207 (N_1207,In_133,In_255);
nor U1208 (N_1208,In_141,In_437);
nand U1209 (N_1209,In_945,In_972);
and U1210 (N_1210,In_266,In_611);
nand U1211 (N_1211,In_245,In_381);
nor U1212 (N_1212,In_796,In_210);
xnor U1213 (N_1213,In_632,In_87);
nor U1214 (N_1214,In_2,In_723);
and U1215 (N_1215,In_55,In_921);
nor U1216 (N_1216,In_477,In_155);
nand U1217 (N_1217,In_557,In_767);
nor U1218 (N_1218,In_756,In_214);
or U1219 (N_1219,In_562,In_884);
and U1220 (N_1220,In_519,In_128);
nor U1221 (N_1221,In_380,In_362);
or U1222 (N_1222,In_274,In_339);
nor U1223 (N_1223,In_907,In_376);
nor U1224 (N_1224,In_877,In_492);
or U1225 (N_1225,In_655,In_601);
nand U1226 (N_1226,In_368,In_223);
or U1227 (N_1227,In_999,In_733);
and U1228 (N_1228,In_616,In_969);
or U1229 (N_1229,In_684,In_293);
nand U1230 (N_1230,In_799,In_142);
and U1231 (N_1231,In_139,In_772);
xor U1232 (N_1232,In_998,In_31);
nand U1233 (N_1233,In_210,In_22);
xnor U1234 (N_1234,In_89,In_997);
nand U1235 (N_1235,In_779,In_735);
nor U1236 (N_1236,In_552,In_255);
nand U1237 (N_1237,In_633,In_579);
or U1238 (N_1238,In_406,In_828);
nand U1239 (N_1239,In_5,In_492);
or U1240 (N_1240,In_119,In_811);
or U1241 (N_1241,In_738,In_583);
nor U1242 (N_1242,In_728,In_907);
nor U1243 (N_1243,In_878,In_706);
nor U1244 (N_1244,In_533,In_852);
nand U1245 (N_1245,In_354,In_232);
nor U1246 (N_1246,In_524,In_264);
nand U1247 (N_1247,In_513,In_142);
or U1248 (N_1248,In_978,In_364);
and U1249 (N_1249,In_232,In_892);
or U1250 (N_1250,In_115,In_824);
and U1251 (N_1251,In_91,In_666);
nand U1252 (N_1252,In_945,In_526);
and U1253 (N_1253,In_682,In_298);
or U1254 (N_1254,In_666,In_787);
and U1255 (N_1255,In_87,In_983);
xor U1256 (N_1256,In_984,In_657);
nor U1257 (N_1257,In_109,In_377);
nor U1258 (N_1258,In_916,In_321);
or U1259 (N_1259,In_564,In_368);
xor U1260 (N_1260,In_943,In_3);
nand U1261 (N_1261,In_13,In_40);
and U1262 (N_1262,In_663,In_591);
and U1263 (N_1263,In_763,In_392);
or U1264 (N_1264,In_202,In_133);
nor U1265 (N_1265,In_145,In_952);
nand U1266 (N_1266,In_980,In_407);
xnor U1267 (N_1267,In_321,In_809);
nor U1268 (N_1268,In_577,In_25);
and U1269 (N_1269,In_956,In_607);
nand U1270 (N_1270,In_107,In_694);
nand U1271 (N_1271,In_334,In_460);
and U1272 (N_1272,In_206,In_549);
and U1273 (N_1273,In_621,In_872);
or U1274 (N_1274,In_114,In_388);
nor U1275 (N_1275,In_169,In_425);
and U1276 (N_1276,In_989,In_220);
nand U1277 (N_1277,In_595,In_495);
nand U1278 (N_1278,In_324,In_198);
xnor U1279 (N_1279,In_188,In_47);
nand U1280 (N_1280,In_515,In_167);
nand U1281 (N_1281,In_346,In_420);
nor U1282 (N_1282,In_67,In_197);
or U1283 (N_1283,In_250,In_941);
nand U1284 (N_1284,In_45,In_734);
nor U1285 (N_1285,In_804,In_670);
nand U1286 (N_1286,In_380,In_231);
nand U1287 (N_1287,In_488,In_563);
nand U1288 (N_1288,In_720,In_378);
nand U1289 (N_1289,In_555,In_381);
or U1290 (N_1290,In_877,In_785);
nor U1291 (N_1291,In_560,In_515);
and U1292 (N_1292,In_102,In_721);
nand U1293 (N_1293,In_654,In_80);
and U1294 (N_1294,In_324,In_322);
nor U1295 (N_1295,In_598,In_315);
or U1296 (N_1296,In_35,In_643);
and U1297 (N_1297,In_547,In_314);
and U1298 (N_1298,In_16,In_487);
nor U1299 (N_1299,In_789,In_759);
xnor U1300 (N_1300,In_517,In_242);
nor U1301 (N_1301,In_713,In_148);
xor U1302 (N_1302,In_641,In_462);
nor U1303 (N_1303,In_50,In_307);
xor U1304 (N_1304,In_848,In_356);
nor U1305 (N_1305,In_608,In_52);
or U1306 (N_1306,In_918,In_670);
nand U1307 (N_1307,In_300,In_813);
nand U1308 (N_1308,In_524,In_599);
or U1309 (N_1309,In_690,In_479);
or U1310 (N_1310,In_238,In_605);
nor U1311 (N_1311,In_390,In_477);
nand U1312 (N_1312,In_110,In_223);
xor U1313 (N_1313,In_695,In_801);
xor U1314 (N_1314,In_437,In_288);
and U1315 (N_1315,In_517,In_135);
nor U1316 (N_1316,In_889,In_771);
nor U1317 (N_1317,In_366,In_732);
and U1318 (N_1318,In_192,In_773);
or U1319 (N_1319,In_171,In_554);
or U1320 (N_1320,In_543,In_883);
or U1321 (N_1321,In_564,In_847);
nand U1322 (N_1322,In_417,In_544);
or U1323 (N_1323,In_819,In_312);
nand U1324 (N_1324,In_717,In_169);
nor U1325 (N_1325,In_566,In_256);
xnor U1326 (N_1326,In_154,In_414);
nor U1327 (N_1327,In_994,In_218);
or U1328 (N_1328,In_439,In_206);
nand U1329 (N_1329,In_244,In_95);
and U1330 (N_1330,In_213,In_161);
or U1331 (N_1331,In_904,In_686);
and U1332 (N_1332,In_247,In_899);
nand U1333 (N_1333,In_843,In_664);
nor U1334 (N_1334,In_23,In_445);
xor U1335 (N_1335,In_794,In_91);
or U1336 (N_1336,In_373,In_709);
nand U1337 (N_1337,In_295,In_76);
nor U1338 (N_1338,In_776,In_137);
xnor U1339 (N_1339,In_238,In_940);
and U1340 (N_1340,In_460,In_694);
nor U1341 (N_1341,In_653,In_634);
nor U1342 (N_1342,In_221,In_826);
nand U1343 (N_1343,In_297,In_121);
nand U1344 (N_1344,In_391,In_666);
nand U1345 (N_1345,In_63,In_272);
and U1346 (N_1346,In_172,In_254);
or U1347 (N_1347,In_276,In_749);
nand U1348 (N_1348,In_530,In_104);
nand U1349 (N_1349,In_717,In_868);
and U1350 (N_1350,In_760,In_733);
nor U1351 (N_1351,In_288,In_845);
or U1352 (N_1352,In_734,In_282);
or U1353 (N_1353,In_225,In_49);
and U1354 (N_1354,In_861,In_359);
nor U1355 (N_1355,In_926,In_561);
and U1356 (N_1356,In_401,In_536);
nor U1357 (N_1357,In_412,In_696);
nand U1358 (N_1358,In_604,In_422);
nand U1359 (N_1359,In_509,In_220);
or U1360 (N_1360,In_833,In_642);
or U1361 (N_1361,In_553,In_127);
nor U1362 (N_1362,In_258,In_815);
nor U1363 (N_1363,In_131,In_385);
xnor U1364 (N_1364,In_98,In_946);
or U1365 (N_1365,In_458,In_582);
nor U1366 (N_1366,In_312,In_314);
and U1367 (N_1367,In_783,In_294);
and U1368 (N_1368,In_666,In_714);
nor U1369 (N_1369,In_760,In_384);
nand U1370 (N_1370,In_734,In_699);
nor U1371 (N_1371,In_923,In_768);
nor U1372 (N_1372,In_431,In_981);
or U1373 (N_1373,In_962,In_681);
nand U1374 (N_1374,In_969,In_69);
or U1375 (N_1375,In_371,In_845);
xnor U1376 (N_1376,In_229,In_112);
nor U1377 (N_1377,In_12,In_364);
nor U1378 (N_1378,In_216,In_366);
and U1379 (N_1379,In_731,In_248);
nand U1380 (N_1380,In_748,In_322);
or U1381 (N_1381,In_241,In_538);
xor U1382 (N_1382,In_205,In_178);
nand U1383 (N_1383,In_220,In_30);
or U1384 (N_1384,In_429,In_609);
nor U1385 (N_1385,In_459,In_503);
xor U1386 (N_1386,In_16,In_816);
xor U1387 (N_1387,In_955,In_807);
xor U1388 (N_1388,In_80,In_151);
and U1389 (N_1389,In_196,In_90);
or U1390 (N_1390,In_931,In_429);
and U1391 (N_1391,In_906,In_630);
nand U1392 (N_1392,In_452,In_662);
and U1393 (N_1393,In_211,In_22);
and U1394 (N_1394,In_574,In_718);
nand U1395 (N_1395,In_344,In_811);
xnor U1396 (N_1396,In_396,In_203);
and U1397 (N_1397,In_116,In_672);
nand U1398 (N_1398,In_476,In_480);
or U1399 (N_1399,In_227,In_565);
and U1400 (N_1400,In_583,In_365);
nand U1401 (N_1401,In_128,In_558);
nor U1402 (N_1402,In_328,In_888);
nor U1403 (N_1403,In_62,In_781);
nand U1404 (N_1404,In_522,In_289);
nand U1405 (N_1405,In_734,In_474);
and U1406 (N_1406,In_673,In_457);
and U1407 (N_1407,In_134,In_718);
nor U1408 (N_1408,In_529,In_367);
and U1409 (N_1409,In_302,In_86);
and U1410 (N_1410,In_601,In_525);
nor U1411 (N_1411,In_606,In_512);
xnor U1412 (N_1412,In_79,In_439);
nor U1413 (N_1413,In_259,In_798);
nand U1414 (N_1414,In_15,In_218);
and U1415 (N_1415,In_753,In_917);
and U1416 (N_1416,In_653,In_650);
nand U1417 (N_1417,In_25,In_251);
nor U1418 (N_1418,In_825,In_791);
xor U1419 (N_1419,In_676,In_736);
nor U1420 (N_1420,In_442,In_738);
xor U1421 (N_1421,In_313,In_785);
and U1422 (N_1422,In_200,In_716);
nor U1423 (N_1423,In_579,In_811);
nand U1424 (N_1424,In_957,In_763);
xnor U1425 (N_1425,In_34,In_821);
or U1426 (N_1426,In_6,In_781);
or U1427 (N_1427,In_811,In_26);
xnor U1428 (N_1428,In_715,In_821);
nor U1429 (N_1429,In_218,In_341);
nand U1430 (N_1430,In_35,In_809);
and U1431 (N_1431,In_501,In_800);
xnor U1432 (N_1432,In_799,In_244);
nor U1433 (N_1433,In_422,In_978);
xor U1434 (N_1434,In_148,In_969);
or U1435 (N_1435,In_601,In_556);
nor U1436 (N_1436,In_273,In_52);
nand U1437 (N_1437,In_425,In_332);
nand U1438 (N_1438,In_892,In_488);
xnor U1439 (N_1439,In_610,In_934);
nand U1440 (N_1440,In_182,In_592);
nand U1441 (N_1441,In_968,In_317);
nor U1442 (N_1442,In_656,In_775);
nor U1443 (N_1443,In_120,In_709);
and U1444 (N_1444,In_859,In_385);
nand U1445 (N_1445,In_841,In_923);
and U1446 (N_1446,In_913,In_961);
nor U1447 (N_1447,In_338,In_915);
xnor U1448 (N_1448,In_729,In_155);
nor U1449 (N_1449,In_88,In_33);
or U1450 (N_1450,In_951,In_316);
and U1451 (N_1451,In_89,In_859);
nor U1452 (N_1452,In_560,In_259);
nand U1453 (N_1453,In_36,In_553);
nor U1454 (N_1454,In_827,In_705);
or U1455 (N_1455,In_68,In_968);
nor U1456 (N_1456,In_59,In_14);
nor U1457 (N_1457,In_869,In_904);
xor U1458 (N_1458,In_92,In_670);
and U1459 (N_1459,In_996,In_776);
and U1460 (N_1460,In_311,In_561);
or U1461 (N_1461,In_994,In_558);
or U1462 (N_1462,In_90,In_349);
nand U1463 (N_1463,In_310,In_988);
nor U1464 (N_1464,In_262,In_389);
and U1465 (N_1465,In_749,In_396);
nor U1466 (N_1466,In_389,In_679);
nand U1467 (N_1467,In_204,In_701);
nor U1468 (N_1468,In_442,In_726);
and U1469 (N_1469,In_667,In_246);
xnor U1470 (N_1470,In_492,In_764);
nand U1471 (N_1471,In_844,In_646);
or U1472 (N_1472,In_316,In_518);
or U1473 (N_1473,In_287,In_299);
nand U1474 (N_1474,In_916,In_398);
and U1475 (N_1475,In_237,In_478);
nor U1476 (N_1476,In_673,In_572);
nand U1477 (N_1477,In_899,In_267);
nand U1478 (N_1478,In_793,In_727);
nand U1479 (N_1479,In_310,In_868);
nand U1480 (N_1480,In_963,In_578);
nor U1481 (N_1481,In_423,In_350);
nand U1482 (N_1482,In_607,In_686);
nor U1483 (N_1483,In_561,In_563);
and U1484 (N_1484,In_293,In_128);
nor U1485 (N_1485,In_370,In_782);
nor U1486 (N_1486,In_246,In_90);
nor U1487 (N_1487,In_783,In_784);
and U1488 (N_1488,In_333,In_463);
or U1489 (N_1489,In_617,In_942);
or U1490 (N_1490,In_286,In_746);
and U1491 (N_1491,In_476,In_516);
and U1492 (N_1492,In_55,In_729);
nand U1493 (N_1493,In_297,In_615);
nand U1494 (N_1494,In_612,In_227);
nand U1495 (N_1495,In_124,In_912);
or U1496 (N_1496,In_246,In_397);
or U1497 (N_1497,In_729,In_32);
nor U1498 (N_1498,In_845,In_550);
nand U1499 (N_1499,In_713,In_390);
or U1500 (N_1500,In_629,In_918);
or U1501 (N_1501,In_909,In_369);
or U1502 (N_1502,In_870,In_676);
nand U1503 (N_1503,In_772,In_338);
nand U1504 (N_1504,In_983,In_321);
nand U1505 (N_1505,In_601,In_79);
and U1506 (N_1506,In_676,In_229);
xnor U1507 (N_1507,In_469,In_637);
or U1508 (N_1508,In_800,In_807);
nand U1509 (N_1509,In_696,In_243);
or U1510 (N_1510,In_538,In_406);
xor U1511 (N_1511,In_87,In_439);
nor U1512 (N_1512,In_798,In_466);
nand U1513 (N_1513,In_304,In_553);
and U1514 (N_1514,In_174,In_151);
and U1515 (N_1515,In_764,In_162);
and U1516 (N_1516,In_124,In_843);
and U1517 (N_1517,In_760,In_925);
nand U1518 (N_1518,In_455,In_308);
nor U1519 (N_1519,In_884,In_593);
xnor U1520 (N_1520,In_748,In_786);
xnor U1521 (N_1521,In_331,In_800);
or U1522 (N_1522,In_267,In_882);
and U1523 (N_1523,In_708,In_949);
nand U1524 (N_1524,In_647,In_879);
nand U1525 (N_1525,In_406,In_914);
and U1526 (N_1526,In_78,In_620);
xnor U1527 (N_1527,In_497,In_702);
and U1528 (N_1528,In_132,In_185);
nand U1529 (N_1529,In_497,In_379);
nand U1530 (N_1530,In_191,In_44);
nor U1531 (N_1531,In_452,In_19);
or U1532 (N_1532,In_904,In_765);
and U1533 (N_1533,In_442,In_589);
nor U1534 (N_1534,In_855,In_970);
or U1535 (N_1535,In_871,In_239);
nor U1536 (N_1536,In_427,In_910);
and U1537 (N_1537,In_945,In_641);
nor U1538 (N_1538,In_76,In_146);
nand U1539 (N_1539,In_838,In_712);
and U1540 (N_1540,In_842,In_355);
nand U1541 (N_1541,In_336,In_856);
or U1542 (N_1542,In_50,In_941);
or U1543 (N_1543,In_41,In_99);
and U1544 (N_1544,In_412,In_553);
nand U1545 (N_1545,In_366,In_406);
nor U1546 (N_1546,In_781,In_35);
nor U1547 (N_1547,In_340,In_44);
and U1548 (N_1548,In_226,In_739);
or U1549 (N_1549,In_2,In_6);
and U1550 (N_1550,In_337,In_275);
nand U1551 (N_1551,In_532,In_324);
and U1552 (N_1552,In_927,In_997);
nand U1553 (N_1553,In_188,In_261);
nor U1554 (N_1554,In_562,In_544);
nor U1555 (N_1555,In_226,In_922);
or U1556 (N_1556,In_59,In_190);
or U1557 (N_1557,In_651,In_35);
nand U1558 (N_1558,In_160,In_76);
nor U1559 (N_1559,In_562,In_393);
xnor U1560 (N_1560,In_62,In_40);
and U1561 (N_1561,In_506,In_171);
or U1562 (N_1562,In_136,In_373);
nor U1563 (N_1563,In_825,In_966);
and U1564 (N_1564,In_141,In_793);
nor U1565 (N_1565,In_766,In_786);
nand U1566 (N_1566,In_646,In_362);
nand U1567 (N_1567,In_13,In_173);
nor U1568 (N_1568,In_175,In_508);
and U1569 (N_1569,In_188,In_128);
and U1570 (N_1570,In_366,In_903);
and U1571 (N_1571,In_808,In_192);
nor U1572 (N_1572,In_417,In_36);
xor U1573 (N_1573,In_986,In_763);
or U1574 (N_1574,In_230,In_103);
nor U1575 (N_1575,In_634,In_964);
and U1576 (N_1576,In_570,In_12);
or U1577 (N_1577,In_199,In_33);
nor U1578 (N_1578,In_917,In_222);
nor U1579 (N_1579,In_95,In_450);
nand U1580 (N_1580,In_280,In_417);
nor U1581 (N_1581,In_640,In_427);
and U1582 (N_1582,In_4,In_789);
nor U1583 (N_1583,In_891,In_355);
nor U1584 (N_1584,In_555,In_323);
or U1585 (N_1585,In_36,In_131);
and U1586 (N_1586,In_413,In_699);
nor U1587 (N_1587,In_623,In_691);
or U1588 (N_1588,In_728,In_700);
and U1589 (N_1589,In_503,In_279);
nor U1590 (N_1590,In_277,In_127);
and U1591 (N_1591,In_224,In_798);
nand U1592 (N_1592,In_651,In_7);
and U1593 (N_1593,In_372,In_445);
and U1594 (N_1594,In_302,In_179);
nand U1595 (N_1595,In_390,In_740);
nand U1596 (N_1596,In_803,In_909);
and U1597 (N_1597,In_522,In_414);
and U1598 (N_1598,In_860,In_857);
nor U1599 (N_1599,In_59,In_24);
and U1600 (N_1600,In_839,In_883);
and U1601 (N_1601,In_433,In_263);
and U1602 (N_1602,In_126,In_139);
or U1603 (N_1603,In_405,In_939);
or U1604 (N_1604,In_351,In_321);
nor U1605 (N_1605,In_645,In_367);
and U1606 (N_1606,In_590,In_364);
nor U1607 (N_1607,In_809,In_626);
nand U1608 (N_1608,In_424,In_720);
nand U1609 (N_1609,In_792,In_738);
nand U1610 (N_1610,In_631,In_82);
nand U1611 (N_1611,In_710,In_27);
or U1612 (N_1612,In_729,In_561);
and U1613 (N_1613,In_523,In_909);
nand U1614 (N_1614,In_279,In_141);
nand U1615 (N_1615,In_259,In_60);
or U1616 (N_1616,In_777,In_301);
and U1617 (N_1617,In_576,In_80);
or U1618 (N_1618,In_629,In_142);
or U1619 (N_1619,In_64,In_989);
and U1620 (N_1620,In_435,In_135);
xor U1621 (N_1621,In_37,In_660);
and U1622 (N_1622,In_687,In_502);
xor U1623 (N_1623,In_829,In_409);
or U1624 (N_1624,In_463,In_519);
nor U1625 (N_1625,In_46,In_508);
xor U1626 (N_1626,In_628,In_194);
or U1627 (N_1627,In_88,In_548);
and U1628 (N_1628,In_179,In_31);
and U1629 (N_1629,In_783,In_289);
nor U1630 (N_1630,In_786,In_473);
and U1631 (N_1631,In_708,In_347);
or U1632 (N_1632,In_935,In_942);
xor U1633 (N_1633,In_749,In_500);
or U1634 (N_1634,In_55,In_840);
or U1635 (N_1635,In_244,In_658);
or U1636 (N_1636,In_153,In_141);
or U1637 (N_1637,In_324,In_528);
or U1638 (N_1638,In_332,In_103);
nor U1639 (N_1639,In_966,In_450);
and U1640 (N_1640,In_429,In_672);
or U1641 (N_1641,In_367,In_273);
nand U1642 (N_1642,In_527,In_671);
xnor U1643 (N_1643,In_966,In_427);
nor U1644 (N_1644,In_147,In_464);
and U1645 (N_1645,In_461,In_679);
or U1646 (N_1646,In_325,In_877);
or U1647 (N_1647,In_714,In_953);
xor U1648 (N_1648,In_631,In_109);
xor U1649 (N_1649,In_990,In_899);
xor U1650 (N_1650,In_839,In_916);
and U1651 (N_1651,In_220,In_805);
or U1652 (N_1652,In_90,In_91);
and U1653 (N_1653,In_745,In_888);
nand U1654 (N_1654,In_996,In_953);
or U1655 (N_1655,In_363,In_299);
nor U1656 (N_1656,In_0,In_835);
or U1657 (N_1657,In_702,In_567);
nor U1658 (N_1658,In_880,In_635);
nand U1659 (N_1659,In_937,In_266);
nor U1660 (N_1660,In_205,In_516);
nor U1661 (N_1661,In_151,In_668);
or U1662 (N_1662,In_839,In_92);
nor U1663 (N_1663,In_997,In_137);
nand U1664 (N_1664,In_260,In_791);
or U1665 (N_1665,In_409,In_530);
nor U1666 (N_1666,In_73,In_145);
or U1667 (N_1667,In_240,In_47);
or U1668 (N_1668,In_226,In_115);
or U1669 (N_1669,In_46,In_268);
nand U1670 (N_1670,In_384,In_236);
nand U1671 (N_1671,In_892,In_313);
and U1672 (N_1672,In_880,In_951);
nand U1673 (N_1673,In_153,In_807);
nand U1674 (N_1674,In_486,In_166);
and U1675 (N_1675,In_888,In_484);
and U1676 (N_1676,In_997,In_183);
and U1677 (N_1677,In_212,In_713);
nor U1678 (N_1678,In_374,In_259);
nand U1679 (N_1679,In_407,In_220);
and U1680 (N_1680,In_538,In_37);
or U1681 (N_1681,In_758,In_708);
and U1682 (N_1682,In_881,In_779);
nand U1683 (N_1683,In_174,In_394);
or U1684 (N_1684,In_646,In_209);
and U1685 (N_1685,In_948,In_23);
and U1686 (N_1686,In_697,In_361);
nor U1687 (N_1687,In_329,In_660);
xnor U1688 (N_1688,In_403,In_920);
and U1689 (N_1689,In_135,In_363);
nand U1690 (N_1690,In_935,In_674);
nand U1691 (N_1691,In_509,In_140);
nor U1692 (N_1692,In_574,In_200);
and U1693 (N_1693,In_378,In_20);
or U1694 (N_1694,In_192,In_660);
nor U1695 (N_1695,In_284,In_106);
xor U1696 (N_1696,In_445,In_70);
and U1697 (N_1697,In_758,In_177);
nor U1698 (N_1698,In_311,In_633);
nand U1699 (N_1699,In_848,In_678);
nor U1700 (N_1700,In_337,In_404);
and U1701 (N_1701,In_46,In_664);
nand U1702 (N_1702,In_467,In_914);
and U1703 (N_1703,In_185,In_195);
nor U1704 (N_1704,In_128,In_963);
nor U1705 (N_1705,In_744,In_140);
nor U1706 (N_1706,In_473,In_996);
and U1707 (N_1707,In_882,In_507);
nor U1708 (N_1708,In_298,In_795);
or U1709 (N_1709,In_400,In_259);
nand U1710 (N_1710,In_939,In_845);
or U1711 (N_1711,In_458,In_448);
or U1712 (N_1712,In_498,In_603);
nor U1713 (N_1713,In_393,In_83);
nor U1714 (N_1714,In_866,In_674);
xnor U1715 (N_1715,In_831,In_9);
xnor U1716 (N_1716,In_707,In_872);
nand U1717 (N_1717,In_276,In_696);
or U1718 (N_1718,In_610,In_990);
xor U1719 (N_1719,In_704,In_330);
or U1720 (N_1720,In_498,In_518);
and U1721 (N_1721,In_415,In_418);
and U1722 (N_1722,In_162,In_878);
and U1723 (N_1723,In_792,In_420);
nor U1724 (N_1724,In_682,In_477);
nand U1725 (N_1725,In_336,In_799);
and U1726 (N_1726,In_340,In_329);
nor U1727 (N_1727,In_780,In_332);
nand U1728 (N_1728,In_988,In_756);
nand U1729 (N_1729,In_509,In_963);
or U1730 (N_1730,In_776,In_486);
and U1731 (N_1731,In_492,In_113);
xnor U1732 (N_1732,In_149,In_244);
and U1733 (N_1733,In_302,In_110);
or U1734 (N_1734,In_96,In_829);
xnor U1735 (N_1735,In_333,In_642);
nor U1736 (N_1736,In_157,In_991);
or U1737 (N_1737,In_939,In_64);
nor U1738 (N_1738,In_93,In_686);
nand U1739 (N_1739,In_909,In_133);
or U1740 (N_1740,In_551,In_856);
or U1741 (N_1741,In_584,In_750);
nor U1742 (N_1742,In_362,In_321);
nand U1743 (N_1743,In_847,In_327);
nor U1744 (N_1744,In_807,In_997);
or U1745 (N_1745,In_199,In_905);
nor U1746 (N_1746,In_212,In_881);
or U1747 (N_1747,In_742,In_121);
nor U1748 (N_1748,In_681,In_240);
and U1749 (N_1749,In_37,In_208);
and U1750 (N_1750,In_724,In_120);
xor U1751 (N_1751,In_969,In_652);
nor U1752 (N_1752,In_949,In_591);
and U1753 (N_1753,In_178,In_957);
xor U1754 (N_1754,In_97,In_757);
or U1755 (N_1755,In_614,In_484);
nor U1756 (N_1756,In_699,In_250);
or U1757 (N_1757,In_598,In_918);
nor U1758 (N_1758,In_618,In_868);
nand U1759 (N_1759,In_872,In_164);
xnor U1760 (N_1760,In_265,In_959);
nor U1761 (N_1761,In_993,In_76);
and U1762 (N_1762,In_114,In_663);
nor U1763 (N_1763,In_431,In_726);
nand U1764 (N_1764,In_388,In_189);
nor U1765 (N_1765,In_868,In_693);
xnor U1766 (N_1766,In_259,In_187);
nor U1767 (N_1767,In_642,In_946);
xor U1768 (N_1768,In_756,In_567);
and U1769 (N_1769,In_572,In_932);
xor U1770 (N_1770,In_284,In_546);
xnor U1771 (N_1771,In_749,In_829);
nand U1772 (N_1772,In_461,In_645);
or U1773 (N_1773,In_468,In_482);
xor U1774 (N_1774,In_261,In_406);
nand U1775 (N_1775,In_720,In_705);
or U1776 (N_1776,In_739,In_685);
xnor U1777 (N_1777,In_585,In_480);
nand U1778 (N_1778,In_567,In_139);
nand U1779 (N_1779,In_477,In_440);
nand U1780 (N_1780,In_412,In_100);
or U1781 (N_1781,In_427,In_651);
or U1782 (N_1782,In_376,In_101);
nand U1783 (N_1783,In_366,In_924);
nand U1784 (N_1784,In_421,In_93);
and U1785 (N_1785,In_85,In_489);
or U1786 (N_1786,In_766,In_797);
nand U1787 (N_1787,In_928,In_178);
nand U1788 (N_1788,In_882,In_398);
nor U1789 (N_1789,In_486,In_439);
or U1790 (N_1790,In_993,In_157);
xnor U1791 (N_1791,In_74,In_496);
nor U1792 (N_1792,In_84,In_1);
and U1793 (N_1793,In_819,In_615);
nand U1794 (N_1794,In_547,In_228);
nand U1795 (N_1795,In_477,In_30);
nor U1796 (N_1796,In_351,In_224);
and U1797 (N_1797,In_710,In_632);
nor U1798 (N_1798,In_950,In_755);
nand U1799 (N_1799,In_743,In_775);
and U1800 (N_1800,In_222,In_712);
nand U1801 (N_1801,In_771,In_596);
nand U1802 (N_1802,In_854,In_21);
or U1803 (N_1803,In_282,In_789);
nand U1804 (N_1804,In_573,In_871);
and U1805 (N_1805,In_930,In_33);
nand U1806 (N_1806,In_127,In_402);
or U1807 (N_1807,In_573,In_976);
and U1808 (N_1808,In_31,In_59);
xnor U1809 (N_1809,In_421,In_499);
xor U1810 (N_1810,In_242,In_832);
nor U1811 (N_1811,In_104,In_493);
or U1812 (N_1812,In_584,In_480);
nor U1813 (N_1813,In_28,In_302);
and U1814 (N_1814,In_816,In_646);
and U1815 (N_1815,In_823,In_382);
or U1816 (N_1816,In_413,In_773);
and U1817 (N_1817,In_112,In_639);
and U1818 (N_1818,In_23,In_772);
or U1819 (N_1819,In_668,In_200);
nand U1820 (N_1820,In_336,In_591);
nand U1821 (N_1821,In_351,In_476);
and U1822 (N_1822,In_899,In_438);
nand U1823 (N_1823,In_409,In_625);
or U1824 (N_1824,In_616,In_623);
or U1825 (N_1825,In_72,In_845);
nand U1826 (N_1826,In_351,In_225);
xor U1827 (N_1827,In_650,In_132);
nor U1828 (N_1828,In_678,In_688);
and U1829 (N_1829,In_762,In_566);
nand U1830 (N_1830,In_948,In_54);
nand U1831 (N_1831,In_484,In_76);
nor U1832 (N_1832,In_649,In_363);
xnor U1833 (N_1833,In_820,In_287);
nor U1834 (N_1834,In_442,In_914);
or U1835 (N_1835,In_140,In_823);
nand U1836 (N_1836,In_720,In_406);
and U1837 (N_1837,In_822,In_596);
or U1838 (N_1838,In_752,In_222);
and U1839 (N_1839,In_865,In_515);
and U1840 (N_1840,In_165,In_509);
or U1841 (N_1841,In_233,In_349);
nor U1842 (N_1842,In_760,In_732);
nor U1843 (N_1843,In_362,In_377);
nand U1844 (N_1844,In_529,In_452);
and U1845 (N_1845,In_659,In_131);
nand U1846 (N_1846,In_382,In_522);
or U1847 (N_1847,In_483,In_526);
nand U1848 (N_1848,In_276,In_506);
or U1849 (N_1849,In_156,In_848);
nor U1850 (N_1850,In_54,In_932);
or U1851 (N_1851,In_584,In_764);
nand U1852 (N_1852,In_571,In_815);
nor U1853 (N_1853,In_313,In_187);
xnor U1854 (N_1854,In_693,In_451);
nand U1855 (N_1855,In_532,In_42);
nand U1856 (N_1856,In_905,In_727);
or U1857 (N_1857,In_444,In_374);
nand U1858 (N_1858,In_523,In_368);
or U1859 (N_1859,In_263,In_450);
and U1860 (N_1860,In_663,In_19);
xnor U1861 (N_1861,In_6,In_293);
nand U1862 (N_1862,In_261,In_14);
and U1863 (N_1863,In_640,In_861);
nor U1864 (N_1864,In_563,In_265);
xor U1865 (N_1865,In_961,In_253);
nand U1866 (N_1866,In_270,In_818);
and U1867 (N_1867,In_675,In_362);
or U1868 (N_1868,In_956,In_12);
nor U1869 (N_1869,In_360,In_499);
nand U1870 (N_1870,In_350,In_92);
nand U1871 (N_1871,In_486,In_191);
and U1872 (N_1872,In_742,In_571);
xor U1873 (N_1873,In_545,In_989);
and U1874 (N_1874,In_293,In_154);
xor U1875 (N_1875,In_56,In_530);
and U1876 (N_1876,In_946,In_853);
xor U1877 (N_1877,In_783,In_700);
nor U1878 (N_1878,In_414,In_974);
xnor U1879 (N_1879,In_152,In_581);
or U1880 (N_1880,In_503,In_143);
nor U1881 (N_1881,In_57,In_950);
nand U1882 (N_1882,In_676,In_271);
xor U1883 (N_1883,In_320,In_514);
or U1884 (N_1884,In_944,In_612);
nand U1885 (N_1885,In_935,In_816);
nand U1886 (N_1886,In_898,In_864);
nor U1887 (N_1887,In_215,In_581);
and U1888 (N_1888,In_583,In_22);
nor U1889 (N_1889,In_422,In_942);
or U1890 (N_1890,In_961,In_118);
or U1891 (N_1891,In_995,In_576);
nor U1892 (N_1892,In_665,In_782);
and U1893 (N_1893,In_487,In_342);
or U1894 (N_1894,In_963,In_6);
or U1895 (N_1895,In_6,In_20);
xnor U1896 (N_1896,In_929,In_282);
and U1897 (N_1897,In_282,In_72);
and U1898 (N_1898,In_765,In_957);
nor U1899 (N_1899,In_276,In_345);
nor U1900 (N_1900,In_595,In_957);
xnor U1901 (N_1901,In_515,In_367);
nor U1902 (N_1902,In_857,In_294);
xor U1903 (N_1903,In_126,In_453);
xor U1904 (N_1904,In_272,In_849);
or U1905 (N_1905,In_155,In_160);
or U1906 (N_1906,In_567,In_606);
nand U1907 (N_1907,In_670,In_99);
or U1908 (N_1908,In_643,In_84);
nand U1909 (N_1909,In_852,In_890);
xnor U1910 (N_1910,In_438,In_503);
nor U1911 (N_1911,In_191,In_536);
or U1912 (N_1912,In_8,In_745);
and U1913 (N_1913,In_241,In_836);
and U1914 (N_1914,In_355,In_716);
and U1915 (N_1915,In_104,In_909);
nor U1916 (N_1916,In_773,In_699);
nor U1917 (N_1917,In_265,In_723);
and U1918 (N_1918,In_133,In_1);
nand U1919 (N_1919,In_720,In_748);
or U1920 (N_1920,In_961,In_374);
and U1921 (N_1921,In_707,In_202);
or U1922 (N_1922,In_895,In_966);
xor U1923 (N_1923,In_223,In_488);
nor U1924 (N_1924,In_948,In_646);
nor U1925 (N_1925,In_555,In_29);
and U1926 (N_1926,In_228,In_944);
nor U1927 (N_1927,In_42,In_692);
and U1928 (N_1928,In_909,In_643);
nor U1929 (N_1929,In_0,In_3);
or U1930 (N_1930,In_253,In_845);
nor U1931 (N_1931,In_688,In_593);
xnor U1932 (N_1932,In_480,In_646);
or U1933 (N_1933,In_904,In_756);
nor U1934 (N_1934,In_916,In_911);
xnor U1935 (N_1935,In_242,In_462);
or U1936 (N_1936,In_855,In_801);
nand U1937 (N_1937,In_408,In_203);
xor U1938 (N_1938,In_105,In_692);
or U1939 (N_1939,In_28,In_69);
xor U1940 (N_1940,In_99,In_171);
nand U1941 (N_1941,In_193,In_466);
or U1942 (N_1942,In_209,In_272);
and U1943 (N_1943,In_318,In_195);
nand U1944 (N_1944,In_525,In_363);
xor U1945 (N_1945,In_41,In_294);
nor U1946 (N_1946,In_790,In_612);
nor U1947 (N_1947,In_721,In_870);
xnor U1948 (N_1948,In_155,In_4);
and U1949 (N_1949,In_836,In_978);
and U1950 (N_1950,In_42,In_806);
nand U1951 (N_1951,In_247,In_684);
nor U1952 (N_1952,In_161,In_508);
nor U1953 (N_1953,In_682,In_206);
and U1954 (N_1954,In_522,In_387);
and U1955 (N_1955,In_617,In_383);
and U1956 (N_1956,In_863,In_400);
nand U1957 (N_1957,In_177,In_333);
nor U1958 (N_1958,In_169,In_978);
and U1959 (N_1959,In_355,In_805);
nand U1960 (N_1960,In_514,In_941);
nand U1961 (N_1961,In_500,In_624);
nand U1962 (N_1962,In_945,In_363);
and U1963 (N_1963,In_698,In_871);
nor U1964 (N_1964,In_857,In_73);
or U1965 (N_1965,In_606,In_149);
nor U1966 (N_1966,In_803,In_61);
nor U1967 (N_1967,In_938,In_219);
xnor U1968 (N_1968,In_868,In_87);
and U1969 (N_1969,In_157,In_582);
nor U1970 (N_1970,In_407,In_890);
and U1971 (N_1971,In_907,In_716);
xor U1972 (N_1972,In_473,In_501);
nor U1973 (N_1973,In_425,In_928);
and U1974 (N_1974,In_756,In_196);
nand U1975 (N_1975,In_546,In_443);
nor U1976 (N_1976,In_958,In_84);
nor U1977 (N_1977,In_236,In_843);
and U1978 (N_1978,In_209,In_26);
nand U1979 (N_1979,In_36,In_550);
or U1980 (N_1980,In_125,In_540);
nand U1981 (N_1981,In_98,In_509);
and U1982 (N_1982,In_206,In_668);
xnor U1983 (N_1983,In_379,In_21);
nand U1984 (N_1984,In_356,In_634);
nand U1985 (N_1985,In_188,In_730);
nor U1986 (N_1986,In_296,In_388);
xnor U1987 (N_1987,In_632,In_180);
nor U1988 (N_1988,In_495,In_43);
and U1989 (N_1989,In_346,In_849);
nand U1990 (N_1990,In_883,In_811);
or U1991 (N_1991,In_661,In_86);
and U1992 (N_1992,In_257,In_521);
and U1993 (N_1993,In_610,In_634);
xor U1994 (N_1994,In_904,In_260);
nor U1995 (N_1995,In_931,In_867);
and U1996 (N_1996,In_77,In_663);
nor U1997 (N_1997,In_584,In_675);
nand U1998 (N_1998,In_53,In_697);
and U1999 (N_1999,In_852,In_56);
nand U2000 (N_2000,In_235,In_906);
nor U2001 (N_2001,In_855,In_46);
nor U2002 (N_2002,In_924,In_943);
and U2003 (N_2003,In_560,In_63);
xor U2004 (N_2004,In_153,In_604);
and U2005 (N_2005,In_695,In_825);
xor U2006 (N_2006,In_258,In_822);
nand U2007 (N_2007,In_471,In_224);
or U2008 (N_2008,In_707,In_274);
nor U2009 (N_2009,In_135,In_362);
nand U2010 (N_2010,In_72,In_868);
or U2011 (N_2011,In_690,In_792);
nor U2012 (N_2012,In_875,In_583);
and U2013 (N_2013,In_45,In_979);
and U2014 (N_2014,In_574,In_734);
nand U2015 (N_2015,In_716,In_282);
nand U2016 (N_2016,In_556,In_194);
or U2017 (N_2017,In_869,In_573);
nor U2018 (N_2018,In_112,In_137);
or U2019 (N_2019,In_836,In_618);
nand U2020 (N_2020,In_95,In_168);
nand U2021 (N_2021,In_829,In_360);
or U2022 (N_2022,In_810,In_213);
nor U2023 (N_2023,In_842,In_145);
and U2024 (N_2024,In_68,In_890);
nand U2025 (N_2025,In_994,In_762);
nor U2026 (N_2026,In_287,In_965);
or U2027 (N_2027,In_120,In_690);
or U2028 (N_2028,In_49,In_809);
and U2029 (N_2029,In_745,In_323);
or U2030 (N_2030,In_616,In_337);
nand U2031 (N_2031,In_161,In_69);
or U2032 (N_2032,In_91,In_362);
xor U2033 (N_2033,In_135,In_633);
xnor U2034 (N_2034,In_540,In_157);
nand U2035 (N_2035,In_637,In_888);
and U2036 (N_2036,In_467,In_543);
nor U2037 (N_2037,In_46,In_651);
nand U2038 (N_2038,In_864,In_257);
xnor U2039 (N_2039,In_430,In_713);
or U2040 (N_2040,In_750,In_647);
xor U2041 (N_2041,In_506,In_103);
xor U2042 (N_2042,In_942,In_482);
xnor U2043 (N_2043,In_320,In_143);
and U2044 (N_2044,In_411,In_88);
nand U2045 (N_2045,In_704,In_297);
and U2046 (N_2046,In_726,In_401);
nor U2047 (N_2047,In_913,In_795);
nor U2048 (N_2048,In_333,In_18);
or U2049 (N_2049,In_677,In_786);
nand U2050 (N_2050,In_221,In_373);
nand U2051 (N_2051,In_613,In_754);
xor U2052 (N_2052,In_226,In_550);
nand U2053 (N_2053,In_936,In_3);
nand U2054 (N_2054,In_333,In_845);
or U2055 (N_2055,In_282,In_357);
xor U2056 (N_2056,In_489,In_469);
or U2057 (N_2057,In_999,In_638);
and U2058 (N_2058,In_85,In_73);
and U2059 (N_2059,In_413,In_176);
and U2060 (N_2060,In_489,In_795);
nand U2061 (N_2061,In_296,In_533);
or U2062 (N_2062,In_346,In_365);
nor U2063 (N_2063,In_628,In_652);
and U2064 (N_2064,In_437,In_142);
and U2065 (N_2065,In_504,In_987);
and U2066 (N_2066,In_862,In_725);
nand U2067 (N_2067,In_308,In_782);
and U2068 (N_2068,In_800,In_951);
and U2069 (N_2069,In_290,In_372);
xnor U2070 (N_2070,In_764,In_92);
nor U2071 (N_2071,In_538,In_985);
or U2072 (N_2072,In_25,In_712);
nor U2073 (N_2073,In_712,In_847);
and U2074 (N_2074,In_895,In_749);
or U2075 (N_2075,In_435,In_675);
nor U2076 (N_2076,In_226,In_558);
nor U2077 (N_2077,In_286,In_249);
nor U2078 (N_2078,In_271,In_455);
or U2079 (N_2079,In_857,In_855);
nor U2080 (N_2080,In_680,In_136);
and U2081 (N_2081,In_406,In_248);
and U2082 (N_2082,In_418,In_608);
xor U2083 (N_2083,In_482,In_985);
nor U2084 (N_2084,In_922,In_462);
and U2085 (N_2085,In_322,In_62);
and U2086 (N_2086,In_176,In_330);
nor U2087 (N_2087,In_704,In_367);
and U2088 (N_2088,In_406,In_316);
and U2089 (N_2089,In_346,In_925);
nand U2090 (N_2090,In_438,In_699);
nor U2091 (N_2091,In_706,In_219);
nand U2092 (N_2092,In_499,In_354);
and U2093 (N_2093,In_892,In_50);
nand U2094 (N_2094,In_89,In_658);
nand U2095 (N_2095,In_964,In_226);
nand U2096 (N_2096,In_137,In_282);
nor U2097 (N_2097,In_776,In_99);
and U2098 (N_2098,In_834,In_666);
and U2099 (N_2099,In_479,In_122);
or U2100 (N_2100,In_140,In_462);
or U2101 (N_2101,In_985,In_731);
nand U2102 (N_2102,In_469,In_902);
nor U2103 (N_2103,In_351,In_8);
nor U2104 (N_2104,In_853,In_454);
nor U2105 (N_2105,In_394,In_981);
nor U2106 (N_2106,In_205,In_267);
or U2107 (N_2107,In_541,In_607);
and U2108 (N_2108,In_989,In_284);
nand U2109 (N_2109,In_40,In_859);
and U2110 (N_2110,In_815,In_650);
nand U2111 (N_2111,In_973,In_204);
nand U2112 (N_2112,In_568,In_20);
or U2113 (N_2113,In_103,In_827);
xnor U2114 (N_2114,In_509,In_903);
xnor U2115 (N_2115,In_303,In_660);
nor U2116 (N_2116,In_819,In_48);
and U2117 (N_2117,In_459,In_470);
nand U2118 (N_2118,In_509,In_919);
xor U2119 (N_2119,In_233,In_724);
nand U2120 (N_2120,In_526,In_116);
and U2121 (N_2121,In_959,In_257);
nor U2122 (N_2122,In_987,In_976);
or U2123 (N_2123,In_264,In_890);
xor U2124 (N_2124,In_625,In_659);
or U2125 (N_2125,In_841,In_884);
or U2126 (N_2126,In_532,In_829);
or U2127 (N_2127,In_759,In_929);
nand U2128 (N_2128,In_113,In_160);
or U2129 (N_2129,In_683,In_273);
nor U2130 (N_2130,In_494,In_623);
xnor U2131 (N_2131,In_313,In_695);
nor U2132 (N_2132,In_211,In_721);
and U2133 (N_2133,In_121,In_867);
nand U2134 (N_2134,In_958,In_420);
nand U2135 (N_2135,In_833,In_870);
nand U2136 (N_2136,In_678,In_105);
xor U2137 (N_2137,In_598,In_753);
nand U2138 (N_2138,In_45,In_712);
nand U2139 (N_2139,In_461,In_318);
nand U2140 (N_2140,In_623,In_839);
and U2141 (N_2141,In_922,In_437);
nand U2142 (N_2142,In_840,In_75);
nand U2143 (N_2143,In_456,In_452);
or U2144 (N_2144,In_591,In_599);
or U2145 (N_2145,In_704,In_194);
nand U2146 (N_2146,In_522,In_180);
and U2147 (N_2147,In_401,In_627);
xnor U2148 (N_2148,In_95,In_836);
and U2149 (N_2149,In_975,In_653);
nor U2150 (N_2150,In_712,In_691);
nand U2151 (N_2151,In_721,In_848);
nor U2152 (N_2152,In_384,In_385);
nand U2153 (N_2153,In_872,In_126);
xnor U2154 (N_2154,In_919,In_133);
and U2155 (N_2155,In_857,In_511);
nor U2156 (N_2156,In_634,In_596);
nand U2157 (N_2157,In_678,In_902);
or U2158 (N_2158,In_726,In_878);
and U2159 (N_2159,In_149,In_426);
nor U2160 (N_2160,In_492,In_480);
nor U2161 (N_2161,In_943,In_500);
or U2162 (N_2162,In_984,In_557);
nand U2163 (N_2163,In_140,In_652);
nand U2164 (N_2164,In_304,In_959);
xor U2165 (N_2165,In_456,In_350);
or U2166 (N_2166,In_834,In_28);
or U2167 (N_2167,In_509,In_143);
nand U2168 (N_2168,In_718,In_211);
or U2169 (N_2169,In_989,In_204);
nor U2170 (N_2170,In_879,In_615);
or U2171 (N_2171,In_177,In_578);
or U2172 (N_2172,In_426,In_898);
nand U2173 (N_2173,In_553,In_608);
nor U2174 (N_2174,In_265,In_37);
nor U2175 (N_2175,In_939,In_543);
xnor U2176 (N_2176,In_600,In_125);
or U2177 (N_2177,In_900,In_696);
nand U2178 (N_2178,In_754,In_351);
and U2179 (N_2179,In_281,In_49);
xnor U2180 (N_2180,In_948,In_160);
nand U2181 (N_2181,In_41,In_606);
nor U2182 (N_2182,In_892,In_988);
nor U2183 (N_2183,In_894,In_839);
or U2184 (N_2184,In_45,In_622);
nor U2185 (N_2185,In_398,In_772);
xor U2186 (N_2186,In_183,In_497);
and U2187 (N_2187,In_794,In_245);
and U2188 (N_2188,In_420,In_652);
or U2189 (N_2189,In_195,In_616);
or U2190 (N_2190,In_83,In_110);
nand U2191 (N_2191,In_926,In_414);
nor U2192 (N_2192,In_127,In_516);
nor U2193 (N_2193,In_981,In_961);
nand U2194 (N_2194,In_725,In_824);
nand U2195 (N_2195,In_739,In_300);
nor U2196 (N_2196,In_71,In_450);
nor U2197 (N_2197,In_806,In_263);
and U2198 (N_2198,In_8,In_735);
nor U2199 (N_2199,In_377,In_617);
xor U2200 (N_2200,In_632,In_998);
nand U2201 (N_2201,In_130,In_708);
nor U2202 (N_2202,In_678,In_239);
nand U2203 (N_2203,In_164,In_619);
xor U2204 (N_2204,In_82,In_761);
nor U2205 (N_2205,In_276,In_237);
nand U2206 (N_2206,In_610,In_532);
nand U2207 (N_2207,In_505,In_464);
or U2208 (N_2208,In_38,In_648);
nand U2209 (N_2209,In_600,In_213);
or U2210 (N_2210,In_165,In_221);
or U2211 (N_2211,In_767,In_92);
nor U2212 (N_2212,In_764,In_694);
and U2213 (N_2213,In_820,In_272);
and U2214 (N_2214,In_837,In_938);
or U2215 (N_2215,In_784,In_87);
nand U2216 (N_2216,In_264,In_743);
or U2217 (N_2217,In_597,In_759);
and U2218 (N_2218,In_627,In_546);
nor U2219 (N_2219,In_90,In_399);
nand U2220 (N_2220,In_731,In_8);
nand U2221 (N_2221,In_232,In_743);
nor U2222 (N_2222,In_308,In_875);
nand U2223 (N_2223,In_213,In_286);
and U2224 (N_2224,In_858,In_138);
nand U2225 (N_2225,In_275,In_638);
nand U2226 (N_2226,In_140,In_931);
xnor U2227 (N_2227,In_765,In_487);
or U2228 (N_2228,In_185,In_623);
or U2229 (N_2229,In_237,In_492);
or U2230 (N_2230,In_825,In_280);
or U2231 (N_2231,In_707,In_676);
nand U2232 (N_2232,In_377,In_601);
nand U2233 (N_2233,In_350,In_292);
nand U2234 (N_2234,In_619,In_687);
nand U2235 (N_2235,In_815,In_61);
nand U2236 (N_2236,In_938,In_574);
and U2237 (N_2237,In_667,In_46);
nor U2238 (N_2238,In_627,In_594);
nand U2239 (N_2239,In_319,In_79);
nand U2240 (N_2240,In_975,In_803);
or U2241 (N_2241,In_926,In_229);
nand U2242 (N_2242,In_582,In_84);
and U2243 (N_2243,In_43,In_839);
nor U2244 (N_2244,In_414,In_306);
nor U2245 (N_2245,In_510,In_56);
nor U2246 (N_2246,In_484,In_775);
nor U2247 (N_2247,In_296,In_765);
and U2248 (N_2248,In_986,In_442);
and U2249 (N_2249,In_480,In_506);
or U2250 (N_2250,In_742,In_315);
and U2251 (N_2251,In_76,In_705);
nand U2252 (N_2252,In_141,In_822);
nand U2253 (N_2253,In_828,In_52);
and U2254 (N_2254,In_474,In_413);
and U2255 (N_2255,In_768,In_206);
or U2256 (N_2256,In_511,In_618);
nand U2257 (N_2257,In_474,In_537);
nand U2258 (N_2258,In_790,In_197);
nand U2259 (N_2259,In_376,In_120);
and U2260 (N_2260,In_722,In_284);
or U2261 (N_2261,In_847,In_277);
and U2262 (N_2262,In_683,In_684);
or U2263 (N_2263,In_642,In_730);
and U2264 (N_2264,In_908,In_944);
nand U2265 (N_2265,In_579,In_128);
nor U2266 (N_2266,In_317,In_648);
nand U2267 (N_2267,In_210,In_670);
and U2268 (N_2268,In_171,In_114);
nor U2269 (N_2269,In_9,In_260);
nand U2270 (N_2270,In_745,In_218);
or U2271 (N_2271,In_79,In_899);
or U2272 (N_2272,In_871,In_263);
nor U2273 (N_2273,In_243,In_735);
nor U2274 (N_2274,In_857,In_475);
nor U2275 (N_2275,In_166,In_471);
nand U2276 (N_2276,In_774,In_755);
nor U2277 (N_2277,In_121,In_714);
or U2278 (N_2278,In_874,In_407);
nand U2279 (N_2279,In_917,In_654);
nand U2280 (N_2280,In_608,In_480);
xnor U2281 (N_2281,In_136,In_454);
xnor U2282 (N_2282,In_302,In_979);
and U2283 (N_2283,In_74,In_56);
and U2284 (N_2284,In_241,In_447);
and U2285 (N_2285,In_74,In_512);
nand U2286 (N_2286,In_196,In_448);
nor U2287 (N_2287,In_494,In_436);
xor U2288 (N_2288,In_752,In_552);
or U2289 (N_2289,In_831,In_896);
nor U2290 (N_2290,In_316,In_449);
xor U2291 (N_2291,In_462,In_593);
nand U2292 (N_2292,In_377,In_871);
and U2293 (N_2293,In_589,In_841);
xnor U2294 (N_2294,In_388,In_700);
and U2295 (N_2295,In_579,In_395);
or U2296 (N_2296,In_326,In_443);
or U2297 (N_2297,In_555,In_590);
or U2298 (N_2298,In_249,In_238);
nand U2299 (N_2299,In_937,In_99);
or U2300 (N_2300,In_680,In_404);
nand U2301 (N_2301,In_963,In_932);
nor U2302 (N_2302,In_31,In_690);
or U2303 (N_2303,In_979,In_887);
nor U2304 (N_2304,In_885,In_954);
nor U2305 (N_2305,In_700,In_482);
or U2306 (N_2306,In_807,In_953);
and U2307 (N_2307,In_650,In_944);
or U2308 (N_2308,In_318,In_241);
nand U2309 (N_2309,In_454,In_762);
nand U2310 (N_2310,In_633,In_661);
nand U2311 (N_2311,In_260,In_965);
and U2312 (N_2312,In_836,In_551);
nand U2313 (N_2313,In_392,In_250);
nand U2314 (N_2314,In_473,In_339);
and U2315 (N_2315,In_419,In_255);
nor U2316 (N_2316,In_553,In_755);
or U2317 (N_2317,In_961,In_280);
nand U2318 (N_2318,In_52,In_914);
and U2319 (N_2319,In_627,In_101);
or U2320 (N_2320,In_317,In_976);
xor U2321 (N_2321,In_931,In_398);
and U2322 (N_2322,In_54,In_462);
or U2323 (N_2323,In_877,In_225);
nor U2324 (N_2324,In_741,In_943);
nor U2325 (N_2325,In_294,In_593);
xor U2326 (N_2326,In_274,In_503);
xnor U2327 (N_2327,In_759,In_554);
nor U2328 (N_2328,In_704,In_874);
nor U2329 (N_2329,In_31,In_51);
and U2330 (N_2330,In_199,In_254);
nand U2331 (N_2331,In_493,In_678);
or U2332 (N_2332,In_816,In_557);
nand U2333 (N_2333,In_328,In_876);
nand U2334 (N_2334,In_370,In_787);
and U2335 (N_2335,In_511,In_448);
and U2336 (N_2336,In_168,In_476);
xor U2337 (N_2337,In_208,In_277);
nor U2338 (N_2338,In_924,In_538);
nand U2339 (N_2339,In_993,In_904);
nor U2340 (N_2340,In_128,In_306);
or U2341 (N_2341,In_695,In_305);
nor U2342 (N_2342,In_41,In_91);
nor U2343 (N_2343,In_978,In_190);
or U2344 (N_2344,In_11,In_294);
and U2345 (N_2345,In_505,In_921);
nand U2346 (N_2346,In_591,In_290);
nand U2347 (N_2347,In_996,In_755);
nor U2348 (N_2348,In_186,In_124);
xor U2349 (N_2349,In_36,In_647);
nor U2350 (N_2350,In_672,In_294);
nand U2351 (N_2351,In_85,In_929);
xor U2352 (N_2352,In_37,In_963);
nand U2353 (N_2353,In_605,In_619);
nand U2354 (N_2354,In_577,In_90);
nand U2355 (N_2355,In_115,In_201);
xor U2356 (N_2356,In_930,In_680);
nand U2357 (N_2357,In_638,In_170);
or U2358 (N_2358,In_102,In_350);
and U2359 (N_2359,In_148,In_441);
or U2360 (N_2360,In_882,In_224);
nor U2361 (N_2361,In_695,In_423);
nand U2362 (N_2362,In_769,In_944);
nand U2363 (N_2363,In_673,In_142);
and U2364 (N_2364,In_953,In_886);
nor U2365 (N_2365,In_539,In_780);
xnor U2366 (N_2366,In_769,In_728);
xnor U2367 (N_2367,In_554,In_567);
nor U2368 (N_2368,In_536,In_943);
nor U2369 (N_2369,In_787,In_815);
nand U2370 (N_2370,In_173,In_334);
or U2371 (N_2371,In_636,In_961);
nor U2372 (N_2372,In_189,In_79);
and U2373 (N_2373,In_787,In_509);
nor U2374 (N_2374,In_606,In_199);
and U2375 (N_2375,In_60,In_613);
nor U2376 (N_2376,In_929,In_793);
and U2377 (N_2377,In_22,In_650);
nor U2378 (N_2378,In_383,In_122);
or U2379 (N_2379,In_787,In_909);
or U2380 (N_2380,In_713,In_405);
and U2381 (N_2381,In_165,In_793);
nor U2382 (N_2382,In_224,In_465);
and U2383 (N_2383,In_385,In_275);
and U2384 (N_2384,In_66,In_124);
and U2385 (N_2385,In_979,In_752);
nor U2386 (N_2386,In_677,In_212);
nor U2387 (N_2387,In_539,In_142);
nor U2388 (N_2388,In_273,In_837);
nor U2389 (N_2389,In_919,In_40);
and U2390 (N_2390,In_667,In_172);
nor U2391 (N_2391,In_407,In_402);
nor U2392 (N_2392,In_521,In_628);
and U2393 (N_2393,In_619,In_182);
xnor U2394 (N_2394,In_197,In_607);
nor U2395 (N_2395,In_612,In_860);
or U2396 (N_2396,In_822,In_452);
nor U2397 (N_2397,In_667,In_476);
xor U2398 (N_2398,In_279,In_84);
xnor U2399 (N_2399,In_430,In_933);
nor U2400 (N_2400,In_974,In_222);
or U2401 (N_2401,In_326,In_984);
nand U2402 (N_2402,In_286,In_962);
nor U2403 (N_2403,In_651,In_467);
nand U2404 (N_2404,In_421,In_322);
or U2405 (N_2405,In_30,In_877);
and U2406 (N_2406,In_592,In_48);
xor U2407 (N_2407,In_3,In_715);
nor U2408 (N_2408,In_960,In_169);
and U2409 (N_2409,In_618,In_503);
or U2410 (N_2410,In_540,In_68);
or U2411 (N_2411,In_37,In_228);
nor U2412 (N_2412,In_396,In_54);
nand U2413 (N_2413,In_198,In_992);
nor U2414 (N_2414,In_640,In_931);
xnor U2415 (N_2415,In_128,In_710);
and U2416 (N_2416,In_747,In_543);
nor U2417 (N_2417,In_477,In_344);
or U2418 (N_2418,In_103,In_693);
nand U2419 (N_2419,In_274,In_387);
and U2420 (N_2420,In_356,In_819);
nand U2421 (N_2421,In_739,In_225);
nor U2422 (N_2422,In_351,In_677);
and U2423 (N_2423,In_375,In_775);
or U2424 (N_2424,In_637,In_720);
or U2425 (N_2425,In_498,In_850);
and U2426 (N_2426,In_381,In_418);
or U2427 (N_2427,In_381,In_994);
nand U2428 (N_2428,In_118,In_638);
and U2429 (N_2429,In_593,In_494);
or U2430 (N_2430,In_30,In_982);
nand U2431 (N_2431,In_611,In_463);
or U2432 (N_2432,In_428,In_716);
nand U2433 (N_2433,In_628,In_758);
nor U2434 (N_2434,In_951,In_673);
nor U2435 (N_2435,In_145,In_511);
xnor U2436 (N_2436,In_443,In_252);
nor U2437 (N_2437,In_588,In_392);
nor U2438 (N_2438,In_486,In_703);
nand U2439 (N_2439,In_104,In_481);
and U2440 (N_2440,In_891,In_330);
and U2441 (N_2441,In_105,In_191);
and U2442 (N_2442,In_508,In_614);
nand U2443 (N_2443,In_582,In_436);
nor U2444 (N_2444,In_49,In_560);
or U2445 (N_2445,In_619,In_39);
nand U2446 (N_2446,In_163,In_233);
nand U2447 (N_2447,In_44,In_665);
xnor U2448 (N_2448,In_952,In_77);
or U2449 (N_2449,In_19,In_623);
and U2450 (N_2450,In_126,In_424);
nor U2451 (N_2451,In_726,In_333);
nand U2452 (N_2452,In_425,In_897);
nand U2453 (N_2453,In_682,In_821);
xor U2454 (N_2454,In_879,In_891);
or U2455 (N_2455,In_479,In_718);
nand U2456 (N_2456,In_664,In_513);
or U2457 (N_2457,In_696,In_699);
or U2458 (N_2458,In_552,In_37);
nand U2459 (N_2459,In_837,In_781);
nor U2460 (N_2460,In_517,In_552);
nor U2461 (N_2461,In_86,In_242);
nor U2462 (N_2462,In_867,In_657);
nor U2463 (N_2463,In_799,In_634);
and U2464 (N_2464,In_195,In_892);
or U2465 (N_2465,In_593,In_585);
and U2466 (N_2466,In_831,In_527);
or U2467 (N_2467,In_730,In_488);
and U2468 (N_2468,In_716,In_1);
nor U2469 (N_2469,In_290,In_117);
and U2470 (N_2470,In_756,In_84);
and U2471 (N_2471,In_424,In_244);
or U2472 (N_2472,In_883,In_469);
nand U2473 (N_2473,In_335,In_857);
nand U2474 (N_2474,In_586,In_790);
and U2475 (N_2475,In_973,In_966);
or U2476 (N_2476,In_873,In_312);
or U2477 (N_2477,In_941,In_272);
xor U2478 (N_2478,In_479,In_533);
or U2479 (N_2479,In_43,In_163);
or U2480 (N_2480,In_814,In_463);
nor U2481 (N_2481,In_621,In_874);
nand U2482 (N_2482,In_792,In_0);
nand U2483 (N_2483,In_788,In_974);
xnor U2484 (N_2484,In_274,In_728);
nand U2485 (N_2485,In_464,In_823);
xor U2486 (N_2486,In_994,In_639);
nand U2487 (N_2487,In_826,In_581);
and U2488 (N_2488,In_960,In_423);
and U2489 (N_2489,In_63,In_454);
or U2490 (N_2490,In_904,In_791);
or U2491 (N_2491,In_34,In_518);
or U2492 (N_2492,In_868,In_249);
and U2493 (N_2493,In_168,In_929);
nand U2494 (N_2494,In_919,In_845);
nand U2495 (N_2495,In_52,In_642);
and U2496 (N_2496,In_773,In_281);
or U2497 (N_2497,In_233,In_88);
xnor U2498 (N_2498,In_681,In_565);
and U2499 (N_2499,In_47,In_288);
or U2500 (N_2500,N_170,N_1519);
xnor U2501 (N_2501,N_1171,N_1521);
or U2502 (N_2502,N_507,N_868);
nand U2503 (N_2503,N_608,N_1516);
nand U2504 (N_2504,N_602,N_518);
xnor U2505 (N_2505,N_1738,N_1283);
nand U2506 (N_2506,N_1024,N_846);
or U2507 (N_2507,N_543,N_1682);
or U2508 (N_2508,N_718,N_715);
nor U2509 (N_2509,N_259,N_678);
or U2510 (N_2510,N_1836,N_1623);
and U2511 (N_2511,N_137,N_1853);
nand U2512 (N_2512,N_370,N_2309);
nand U2513 (N_2513,N_169,N_2385);
or U2514 (N_2514,N_1637,N_2460);
or U2515 (N_2515,N_2069,N_977);
nand U2516 (N_2516,N_1008,N_510);
nand U2517 (N_2517,N_1823,N_311);
and U2518 (N_2518,N_1176,N_1857);
nor U2519 (N_2519,N_304,N_1935);
and U2520 (N_2520,N_2198,N_388);
xnor U2521 (N_2521,N_2290,N_859);
nand U2522 (N_2522,N_1760,N_605);
nor U2523 (N_2523,N_579,N_2495);
nor U2524 (N_2524,N_1724,N_1380);
and U2525 (N_2525,N_1622,N_1494);
xor U2526 (N_2526,N_1215,N_2033);
and U2527 (N_2527,N_922,N_251);
or U2528 (N_2528,N_1896,N_329);
nor U2529 (N_2529,N_905,N_1302);
or U2530 (N_2530,N_622,N_1107);
nor U2531 (N_2531,N_164,N_618);
or U2532 (N_2532,N_1360,N_2348);
nor U2533 (N_2533,N_469,N_955);
or U2534 (N_2534,N_932,N_1767);
or U2535 (N_2535,N_1467,N_2444);
nand U2536 (N_2536,N_731,N_382);
xnor U2537 (N_2537,N_2381,N_2097);
nor U2538 (N_2538,N_939,N_691);
nor U2539 (N_2539,N_1750,N_398);
and U2540 (N_2540,N_1872,N_1928);
or U2541 (N_2541,N_942,N_1814);
or U2542 (N_2542,N_941,N_1725);
nor U2543 (N_2543,N_504,N_1644);
nor U2544 (N_2544,N_1390,N_2325);
and U2545 (N_2545,N_1414,N_30);
nand U2546 (N_2546,N_574,N_663);
nor U2547 (N_2547,N_235,N_295);
or U2548 (N_2548,N_289,N_577);
or U2549 (N_2549,N_16,N_2240);
and U2550 (N_2550,N_1621,N_88);
nand U2551 (N_2551,N_1581,N_98);
and U2552 (N_2552,N_179,N_529);
or U2553 (N_2553,N_1227,N_1676);
xnor U2554 (N_2554,N_314,N_2032);
nand U2555 (N_2555,N_644,N_2117);
nand U2556 (N_2556,N_843,N_769);
nand U2557 (N_2557,N_476,N_1709);
nand U2558 (N_2558,N_2091,N_813);
nor U2559 (N_2559,N_1347,N_2286);
and U2560 (N_2560,N_1148,N_869);
or U2561 (N_2561,N_340,N_856);
and U2562 (N_2562,N_805,N_1728);
or U2563 (N_2563,N_2367,N_2114);
and U2564 (N_2564,N_944,N_1334);
or U2565 (N_2565,N_1358,N_2284);
and U2566 (N_2566,N_2236,N_836);
and U2567 (N_2567,N_426,N_162);
xor U2568 (N_2568,N_109,N_756);
and U2569 (N_2569,N_218,N_828);
nor U2570 (N_2570,N_584,N_1807);
nor U2571 (N_2571,N_1319,N_1815);
or U2572 (N_2572,N_1554,N_190);
and U2573 (N_2573,N_1982,N_2071);
nand U2574 (N_2574,N_2010,N_1971);
xor U2575 (N_2575,N_509,N_1580);
nand U2576 (N_2576,N_2149,N_1256);
nand U2577 (N_2577,N_1714,N_430);
nand U2578 (N_2578,N_196,N_435);
or U2579 (N_2579,N_403,N_397);
nand U2580 (N_2580,N_1752,N_297);
or U2581 (N_2581,N_1469,N_1432);
xnor U2582 (N_2582,N_822,N_1963);
or U2583 (N_2583,N_1854,N_659);
nand U2584 (N_2584,N_1568,N_1055);
nor U2585 (N_2585,N_1450,N_1100);
nor U2586 (N_2586,N_1680,N_904);
nand U2587 (N_2587,N_146,N_848);
nand U2588 (N_2588,N_776,N_159);
nand U2589 (N_2589,N_2353,N_188);
nor U2590 (N_2590,N_2441,N_273);
nand U2591 (N_2591,N_2219,N_2062);
and U2592 (N_2592,N_2055,N_1995);
nand U2593 (N_2593,N_2394,N_1754);
nor U2594 (N_2594,N_1921,N_1603);
or U2595 (N_2595,N_1789,N_734);
and U2596 (N_2596,N_1242,N_1972);
nand U2597 (N_2597,N_2247,N_2014);
nand U2598 (N_2598,N_1050,N_632);
nor U2599 (N_2599,N_645,N_1882);
nor U2600 (N_2600,N_724,N_399);
nor U2601 (N_2601,N_1371,N_409);
nor U2602 (N_2602,N_1488,N_864);
nor U2603 (N_2603,N_472,N_1284);
nand U2604 (N_2604,N_2250,N_1240);
nand U2605 (N_2605,N_199,N_626);
or U2606 (N_2606,N_1718,N_1298);
xnor U2607 (N_2607,N_566,N_432);
or U2608 (N_2608,N_407,N_2281);
nor U2609 (N_2609,N_1914,N_1939);
or U2610 (N_2610,N_1431,N_231);
nor U2611 (N_2611,N_604,N_1268);
nor U2612 (N_2612,N_606,N_406);
and U2613 (N_2613,N_1213,N_594);
nor U2614 (N_2614,N_1786,N_1065);
nand U2615 (N_2615,N_2100,N_1926);
or U2616 (N_2616,N_1003,N_2446);
nor U2617 (N_2617,N_132,N_1465);
and U2618 (N_2618,N_107,N_1799);
nor U2619 (N_2619,N_819,N_1341);
nor U2620 (N_2620,N_466,N_1688);
nor U2621 (N_2621,N_375,N_1920);
or U2622 (N_2622,N_893,N_160);
or U2623 (N_2623,N_286,N_1210);
or U2624 (N_2624,N_910,N_1613);
and U2625 (N_2625,N_569,N_2392);
nand U2626 (N_2626,N_2244,N_110);
nand U2627 (N_2627,N_1626,N_797);
xnor U2628 (N_2628,N_2484,N_1652);
and U2629 (N_2629,N_2169,N_1784);
nor U2630 (N_2630,N_1706,N_924);
and U2631 (N_2631,N_1229,N_177);
and U2632 (N_2632,N_1116,N_275);
nand U2633 (N_2633,N_1906,N_272);
or U2634 (N_2634,N_1086,N_2153);
or U2635 (N_2635,N_2344,N_654);
nor U2636 (N_2636,N_442,N_1424);
or U2637 (N_2637,N_559,N_371);
or U2638 (N_2638,N_60,N_1440);
xor U2639 (N_2639,N_1657,N_1707);
nand U2640 (N_2640,N_1635,N_1727);
or U2641 (N_2641,N_637,N_1983);
xor U2642 (N_2642,N_330,N_2180);
or U2643 (N_2643,N_1113,N_1878);
xor U2644 (N_2644,N_2186,N_281);
nor U2645 (N_2645,N_2369,N_2081);
or U2646 (N_2646,N_589,N_1606);
xor U2647 (N_2647,N_1902,N_908);
nand U2648 (N_2648,N_1550,N_1220);
nand U2649 (N_2649,N_1620,N_940);
or U2650 (N_2650,N_243,N_1000);
nor U2651 (N_2651,N_2245,N_37);
nor U2652 (N_2652,N_1993,N_1861);
nand U2653 (N_2653,N_2220,N_532);
and U2654 (N_2654,N_1761,N_2422);
nor U2655 (N_2655,N_439,N_1091);
and U2656 (N_2656,N_1595,N_981);
and U2657 (N_2657,N_542,N_1930);
or U2658 (N_2658,N_624,N_154);
xnor U2659 (N_2659,N_1910,N_1559);
or U2660 (N_2660,N_1455,N_555);
nor U2661 (N_2661,N_158,N_706);
or U2662 (N_2662,N_1933,N_392);
and U2663 (N_2663,N_413,N_593);
nor U2664 (N_2664,N_1967,N_1740);
nor U2665 (N_2665,N_1437,N_827);
nand U2666 (N_2666,N_1439,N_2261);
and U2667 (N_2667,N_1790,N_29);
and U2668 (N_2668,N_517,N_2167);
nor U2669 (N_2669,N_2351,N_2395);
nor U2670 (N_2670,N_1045,N_293);
or U2671 (N_2671,N_2104,N_809);
or U2672 (N_2672,N_1479,N_1736);
nor U2673 (N_2673,N_309,N_2194);
or U2674 (N_2674,N_866,N_2451);
nand U2675 (N_2675,N_2354,N_1246);
nor U2676 (N_2676,N_2205,N_2127);
nand U2677 (N_2677,N_50,N_2306);
or U2678 (N_2678,N_775,N_1075);
nor U2679 (N_2679,N_1571,N_1397);
and U2680 (N_2680,N_1490,N_1837);
nor U2681 (N_2681,N_1041,N_1865);
and U2682 (N_2682,N_919,N_1043);
and U2683 (N_2683,N_473,N_96);
and U2684 (N_2684,N_2314,N_2263);
nor U2685 (N_2685,N_1140,N_308);
xnor U2686 (N_2686,N_198,N_488);
or U2687 (N_2687,N_1452,N_1286);
nand U2688 (N_2688,N_2120,N_1591);
nor U2689 (N_2689,N_909,N_172);
nor U2690 (N_2690,N_2289,N_581);
or U2691 (N_2691,N_357,N_1124);
and U2692 (N_2692,N_523,N_355);
and U2693 (N_2693,N_2073,N_2461);
or U2694 (N_2694,N_1764,N_679);
and U2695 (N_2695,N_2349,N_524);
nor U2696 (N_2696,N_2296,N_512);
nand U2697 (N_2697,N_52,N_2378);
nand U2698 (N_2698,N_511,N_1868);
nand U2699 (N_2699,N_873,N_2402);
and U2700 (N_2700,N_45,N_1946);
or U2701 (N_2701,N_693,N_2278);
nor U2702 (N_2702,N_935,N_625);
xor U2703 (N_2703,N_1405,N_2195);
or U2704 (N_2704,N_571,N_300);
nor U2705 (N_2705,N_248,N_1998);
and U2706 (N_2706,N_182,N_1570);
nand U2707 (N_2707,N_2485,N_482);
nor U2708 (N_2708,N_2360,N_484);
and U2709 (N_2709,N_1968,N_2396);
xnor U2710 (N_2710,N_751,N_389);
nor U2711 (N_2711,N_1632,N_2438);
nand U2712 (N_2712,N_1014,N_1083);
nand U2713 (N_2713,N_168,N_2018);
or U2714 (N_2714,N_1458,N_1330);
or U2715 (N_2715,N_1012,N_149);
nor U2716 (N_2716,N_1354,N_214);
nor U2717 (N_2717,N_546,N_1106);
or U2718 (N_2718,N_669,N_1834);
or U2719 (N_2719,N_1819,N_43);
nor U2720 (N_2720,N_2144,N_268);
or U2721 (N_2721,N_665,N_2199);
or U2722 (N_2722,N_2406,N_140);
nand U2723 (N_2723,N_1959,N_1451);
nand U2724 (N_2724,N_1406,N_2355);
nor U2725 (N_2725,N_1460,N_1313);
and U2726 (N_2726,N_239,N_1957);
nand U2727 (N_2727,N_233,N_1700);
xor U2728 (N_2728,N_2039,N_287);
and U2729 (N_2729,N_264,N_642);
nand U2730 (N_2730,N_1690,N_1130);
or U2731 (N_2731,N_2159,N_368);
nand U2732 (N_2732,N_1534,N_1942);
and U2733 (N_2733,N_1847,N_242);
and U2734 (N_2734,N_1185,N_62);
xnor U2735 (N_2735,N_1687,N_2157);
or U2736 (N_2736,N_1053,N_2259);
or U2737 (N_2737,N_26,N_2356);
nor U2738 (N_2738,N_1333,N_70);
or U2739 (N_2739,N_1990,N_1303);
or U2740 (N_2740,N_232,N_2374);
xor U2741 (N_2741,N_2022,N_1427);
nor U2742 (N_2742,N_1395,N_1594);
nand U2743 (N_2743,N_2376,N_2477);
nor U2744 (N_2744,N_1773,N_1007);
and U2745 (N_2745,N_1785,N_1156);
nor U2746 (N_2746,N_2177,N_2212);
or U2747 (N_2747,N_2099,N_1264);
or U2748 (N_2748,N_1127,N_1295);
nand U2749 (N_2749,N_470,N_1708);
and U2750 (N_2750,N_1989,N_2276);
nand U2751 (N_2751,N_796,N_2175);
nor U2752 (N_2752,N_1111,N_1693);
xor U2753 (N_2753,N_1239,N_2472);
and U2754 (N_2754,N_993,N_334);
or U2755 (N_2755,N_24,N_420);
nand U2756 (N_2756,N_47,N_2308);
nor U2757 (N_2757,N_2371,N_163);
nand U2758 (N_2758,N_206,N_408);
and U2759 (N_2759,N_477,N_1563);
nor U2760 (N_2760,N_1511,N_1590);
or U2761 (N_2761,N_1310,N_486);
nor U2762 (N_2762,N_1378,N_987);
and U2763 (N_2763,N_1179,N_2137);
or U2764 (N_2764,N_479,N_2124);
and U2765 (N_2765,N_968,N_1308);
xor U2766 (N_2766,N_203,N_1673);
nor U2767 (N_2767,N_535,N_774);
nor U2768 (N_2768,N_1775,N_2035);
nand U2769 (N_2769,N_156,N_1477);
and U2770 (N_2770,N_2103,N_830);
or U2771 (N_2771,N_781,N_1842);
or U2772 (N_2772,N_305,N_1574);
xor U2773 (N_2773,N_570,N_1115);
nand U2774 (N_2774,N_551,N_94);
and U2775 (N_2775,N_36,N_241);
or U2776 (N_2776,N_2203,N_640);
nor U2777 (N_2777,N_789,N_2383);
nor U2778 (N_2778,N_1901,N_597);
nor U2779 (N_2779,N_2301,N_1869);
nand U2780 (N_2780,N_2453,N_1871);
nand U2781 (N_2781,N_2054,N_2478);
xor U2782 (N_2782,N_2012,N_966);
or U2783 (N_2783,N_750,N_1146);
and U2784 (N_2784,N_252,N_1355);
nor U2785 (N_2785,N_2115,N_684);
nand U2786 (N_2786,N_1028,N_347);
and U2787 (N_2787,N_1481,N_770);
and U2788 (N_2788,N_1648,N_82);
or U2789 (N_2789,N_1304,N_658);
nand U2790 (N_2790,N_262,N_880);
nand U2791 (N_2791,N_1938,N_1058);
xnor U2792 (N_2792,N_758,N_2304);
nand U2793 (N_2793,N_2227,N_267);
nand U2794 (N_2794,N_1833,N_1974);
xnor U2795 (N_2795,N_1634,N_1300);
nand U2796 (N_2796,N_204,N_1748);
xnor U2797 (N_2797,N_19,N_1779);
and U2798 (N_2798,N_1248,N_683);
nand U2799 (N_2799,N_2345,N_2454);
and U2800 (N_2800,N_2447,N_1154);
nor U2801 (N_2801,N_1658,N_1429);
or U2802 (N_2802,N_326,N_1562);
nand U2803 (N_2803,N_902,N_2106);
nor U2804 (N_2804,N_1801,N_1607);
or U2805 (N_2805,N_741,N_2098);
and U2806 (N_2806,N_2173,N_906);
nand U2807 (N_2807,N_849,N_1020);
nand U2808 (N_2808,N_590,N_1164);
or U2809 (N_2809,N_1653,N_483);
nand U2810 (N_2810,N_1218,N_1040);
and U2811 (N_2811,N_35,N_953);
nor U2812 (N_2812,N_1198,N_2464);
nand U2813 (N_2813,N_1977,N_1943);
or U2814 (N_2814,N_301,N_950);
or U2815 (N_2815,N_653,N_844);
nand U2816 (N_2816,N_898,N_1739);
nand U2817 (N_2817,N_1763,N_1699);
or U2818 (N_2818,N_2246,N_1484);
nand U2819 (N_2819,N_2067,N_2299);
nand U2820 (N_2820,N_1586,N_2235);
and U2821 (N_2821,N_2229,N_1120);
nand U2822 (N_2822,N_2206,N_97);
and U2823 (N_2823,N_1951,N_1415);
or U2824 (N_2824,N_1464,N_2211);
nand U2825 (N_2825,N_84,N_1636);
or U2826 (N_2826,N_2498,N_205);
or U2827 (N_2827,N_1755,N_2338);
nor U2828 (N_2828,N_1069,N_2074);
nand U2829 (N_2829,N_851,N_900);
and U2830 (N_2830,N_708,N_318);
and U2831 (N_2831,N_2357,N_1889);
and U2832 (N_2832,N_554,N_1093);
nand U2833 (N_2833,N_2092,N_564);
or U2834 (N_2834,N_1022,N_2189);
and U2835 (N_2835,N_807,N_1202);
and U2836 (N_2836,N_2280,N_1772);
nand U2837 (N_2837,N_285,N_219);
and U2838 (N_2838,N_2427,N_1403);
nand U2839 (N_2839,N_220,N_1436);
nor U2840 (N_2840,N_129,N_1733);
or U2841 (N_2841,N_2486,N_2366);
xor U2842 (N_2842,N_2285,N_1895);
or U2843 (N_2843,N_607,N_1238);
or U2844 (N_2844,N_531,N_2430);
xor U2845 (N_2845,N_991,N_565);
or U2846 (N_2846,N_1207,N_8);
xor U2847 (N_2847,N_387,N_1487);
or U2848 (N_2848,N_346,N_612);
nor U2849 (N_2849,N_2494,N_1247);
nand U2850 (N_2850,N_1862,N_1316);
or U2851 (N_2851,N_1698,N_1234);
and U2852 (N_2852,N_401,N_1717);
nor U2853 (N_2853,N_1810,N_1670);
nor U2854 (N_2854,N_1934,N_1720);
or U2855 (N_2855,N_694,N_1966);
nand U2856 (N_2856,N_316,N_2408);
or U2857 (N_2857,N_1241,N_2463);
or U2858 (N_2858,N_276,N_258);
or U2859 (N_2859,N_891,N_1922);
xor U2860 (N_2860,N_460,N_467);
or U2861 (N_2861,N_2416,N_1281);
and U2862 (N_2862,N_537,N_530);
xnor U2863 (N_2863,N_1030,N_2048);
xor U2864 (N_2864,N_506,N_761);
nor U2865 (N_2865,N_391,N_480);
nor U2866 (N_2866,N_970,N_2028);
xnor U2867 (N_2867,N_2087,N_1541);
and U2868 (N_2868,N_2056,N_1150);
nand U2869 (N_2869,N_767,N_277);
nor U2870 (N_2870,N_1749,N_2213);
nor U2871 (N_2871,N_2340,N_1409);
xnor U2872 (N_2872,N_328,N_38);
and U2873 (N_2873,N_1449,N_1924);
or U2874 (N_2874,N_651,N_911);
xor U2875 (N_2875,N_870,N_1734);
nand U2876 (N_2876,N_918,N_1816);
nor U2877 (N_2877,N_1004,N_1025);
or U2878 (N_2878,N_490,N_437);
and U2879 (N_2879,N_829,N_1167);
nor U2880 (N_2880,N_675,N_178);
nand U2881 (N_2881,N_1619,N_553);
and U2882 (N_2882,N_1592,N_1293);
xor U2883 (N_2883,N_1279,N_254);
nand U2884 (N_2884,N_87,N_2359);
and U2885 (N_2885,N_1155,N_1471);
or U2886 (N_2886,N_1413,N_863);
and U2887 (N_2887,N_1518,N_2027);
and U2888 (N_2888,N_1737,N_1783);
nand U2889 (N_2889,N_702,N_1766);
and U2890 (N_2890,N_2119,N_2493);
xnor U2891 (N_2891,N_485,N_1110);
nand U2892 (N_2892,N_886,N_945);
nor U2893 (N_2893,N_973,N_985);
or U2894 (N_2894,N_1422,N_996);
nand U2895 (N_2895,N_1265,N_1078);
nor U2896 (N_2896,N_974,N_1735);
or U2897 (N_2897,N_1407,N_106);
xnor U2898 (N_2898,N_1999,N_882);
and U2899 (N_2899,N_1660,N_1042);
nor U2900 (N_2900,N_2118,N_1224);
nor U2901 (N_2901,N_1369,N_1362);
and U2902 (N_2902,N_151,N_1618);
and U2903 (N_2903,N_760,N_1715);
nand U2904 (N_2904,N_112,N_324);
and U2905 (N_2905,N_1074,N_1668);
xnor U2906 (N_2906,N_447,N_1037);
xnor U2907 (N_2907,N_519,N_200);
or U2908 (N_2908,N_1143,N_1480);
nor U2909 (N_2909,N_253,N_575);
and U2910 (N_2910,N_855,N_1884);
nor U2911 (N_2911,N_1153,N_157);
nand U2912 (N_2912,N_1824,N_1525);
nor U2913 (N_2913,N_1252,N_343);
and U2914 (N_2914,N_1945,N_723);
or U2915 (N_2915,N_647,N_730);
xor U2916 (N_2916,N_2252,N_1894);
nand U2917 (N_2917,N_1776,N_1898);
nand U2918 (N_2918,N_260,N_302);
or U2919 (N_2919,N_2372,N_1142);
xor U2920 (N_2920,N_2302,N_325);
or U2921 (N_2921,N_2421,N_717);
nand U2922 (N_2922,N_1551,N_321);
xnor U2923 (N_2923,N_1170,N_838);
nand U2924 (N_2924,N_126,N_1498);
and U2925 (N_2925,N_1345,N_705);
nand U2926 (N_2926,N_2313,N_1235);
or U2927 (N_2927,N_458,N_1604);
and U2928 (N_2928,N_1643,N_1492);
or U2929 (N_2929,N_1031,N_1923);
and U2930 (N_2930,N_411,N_646);
nand U2931 (N_2931,N_2168,N_93);
or U2932 (N_2932,N_609,N_513);
nor U2933 (N_2933,N_1173,N_729);
nand U2934 (N_2934,N_1290,N_1875);
or U2935 (N_2935,N_634,N_1088);
and U2936 (N_2936,N_23,N_1965);
nor U2937 (N_2937,N_1629,N_2139);
and U2938 (N_2938,N_2011,N_2476);
xnor U2939 (N_2939,N_785,N_1277);
nand U2940 (N_2940,N_2434,N_1121);
and U2941 (N_2941,N_1332,N_2174);
xor U2942 (N_2942,N_374,N_1956);
and U2943 (N_2943,N_739,N_1909);
or U2944 (N_2944,N_1561,N_10);
nor U2945 (N_2945,N_2499,N_1805);
and U2946 (N_2946,N_587,N_410);
nand U2947 (N_2947,N_2185,N_2002);
nor U2948 (N_2948,N_2342,N_144);
nand U2949 (N_2949,N_448,N_2319);
nand U2950 (N_2950,N_2347,N_2231);
nand U2951 (N_2951,N_1062,N_1986);
or U2952 (N_2952,N_703,N_290);
nor U2953 (N_2953,N_320,N_2249);
and U2954 (N_2954,N_1245,N_1496);
nand U2955 (N_2955,N_766,N_103);
nor U2956 (N_2956,N_2310,N_496);
xor U2957 (N_2957,N_440,N_635);
or U2958 (N_2958,N_857,N_453);
xnor U2959 (N_2959,N_240,N_15);
nor U2960 (N_2960,N_424,N_53);
or U2961 (N_2961,N_712,N_1102);
nor U2962 (N_2962,N_892,N_319);
nor U2963 (N_2963,N_428,N_1681);
nor U2964 (N_2964,N_487,N_465);
or U2965 (N_2965,N_2420,N_788);
nor U2966 (N_2966,N_135,N_211);
and U2967 (N_2967,N_1122,N_1444);
xnor U2968 (N_2968,N_130,N_79);
nand U2969 (N_2969,N_527,N_1015);
nor U2970 (N_2970,N_595,N_1157);
nand U2971 (N_2971,N_1159,N_299);
and U2972 (N_2972,N_1840,N_377);
xor U2973 (N_2973,N_1915,N_643);
xor U2974 (N_2974,N_1510,N_2196);
and U2975 (N_2975,N_349,N_1070);
and U2976 (N_2976,N_2152,N_1001);
nand U2977 (N_2977,N_2192,N_1199);
xor U2978 (N_2978,N_984,N_284);
nand U2979 (N_2979,N_1255,N_2140);
or U2980 (N_2980,N_1839,N_429);
or U2981 (N_2981,N_433,N_1677);
or U2982 (N_2982,N_1539,N_2215);
or U2983 (N_2983,N_2233,N_2);
nand U2984 (N_2984,N_2232,N_274);
nand U2985 (N_2985,N_1389,N_64);
nor U2986 (N_2986,N_2172,N_786);
nand U2987 (N_2987,N_494,N_1294);
nand U2988 (N_2988,N_2007,N_457);
and U2989 (N_2989,N_1565,N_95);
nand U2990 (N_2990,N_2295,N_394);
or U2991 (N_2991,N_44,N_2228);
or U2992 (N_2992,N_1524,N_1285);
and U2993 (N_2993,N_733,N_1232);
nand U2994 (N_2994,N_655,N_216);
nand U2995 (N_2995,N_1503,N_1309);
or U2996 (N_2996,N_68,N_1529);
or U2997 (N_2997,N_1585,N_752);
or U2998 (N_2998,N_1970,N_247);
or U2999 (N_2999,N_2082,N_1152);
nand U3000 (N_3000,N_461,N_1278);
and U3001 (N_3001,N_127,N_719);
or U3002 (N_3002,N_1411,N_2428);
and U3003 (N_3003,N_361,N_2467);
nand U3004 (N_3004,N_1583,N_695);
or U3005 (N_3005,N_1843,N_948);
nand U3006 (N_3006,N_1271,N_1456);
nor U3007 (N_3007,N_315,N_115);
or U3008 (N_3008,N_2274,N_1689);
nand U3009 (N_3009,N_871,N_1434);
and U3010 (N_3010,N_1954,N_1892);
or U3011 (N_3011,N_1701,N_2487);
xor U3012 (N_3012,N_826,N_2272);
nor U3013 (N_3013,N_656,N_1447);
xnor U3014 (N_3014,N_337,N_1553);
and U3015 (N_3015,N_2390,N_1064);
nand U3016 (N_3016,N_1722,N_888);
nand U3017 (N_3017,N_2025,N_1705);
or U3018 (N_3018,N_1532,N_54);
or U3019 (N_3019,N_815,N_623);
or U3020 (N_3020,N_1537,N_1289);
nand U3021 (N_3021,N_66,N_2145);
and U3022 (N_3022,N_1557,N_1117);
or U3023 (N_3023,N_456,N_2459);
and U3024 (N_3024,N_1393,N_215);
nor U3025 (N_3025,N_1588,N_257);
nand U3026 (N_3026,N_2267,N_1335);
xor U3027 (N_3027,N_999,N_2490);
nand U3028 (N_3028,N_503,N_2497);
nand U3029 (N_3029,N_806,N_1034);
or U3030 (N_3030,N_1504,N_1713);
or U3031 (N_3031,N_1791,N_2411);
xnor U3032 (N_3032,N_2305,N_74);
nand U3033 (N_3033,N_1474,N_842);
nor U3034 (N_3034,N_1796,N_1082);
nor U3035 (N_3035,N_794,N_847);
xor U3036 (N_3036,N_936,N_183);
nand U3037 (N_3037,N_2243,N_954);
nand U3038 (N_3038,N_998,N_613);
nor U3039 (N_3039,N_2405,N_283);
xor U3040 (N_3040,N_920,N_2270);
and U3041 (N_3041,N_256,N_313);
and U3042 (N_3042,N_1134,N_2455);
nand U3043 (N_3043,N_1527,N_2101);
nand U3044 (N_3044,N_816,N_1408);
nand U3045 (N_3045,N_148,N_463);
and U3046 (N_3046,N_1359,N_883);
or U3047 (N_3047,N_526,N_1960);
or U3048 (N_3048,N_2064,N_1009);
nand U3049 (N_3049,N_1169,N_1318);
nor U3050 (N_3050,N_495,N_1297);
or U3051 (N_3051,N_185,N_1367);
and U3052 (N_3052,N_586,N_221);
nand U3053 (N_3053,N_744,N_2297);
nand U3054 (N_3054,N_475,N_1777);
and U3055 (N_3055,N_1747,N_765);
and U3056 (N_3056,N_1640,N_2063);
and U3057 (N_3057,N_2134,N_2316);
nand U3058 (N_3058,N_1052,N_657);
or U3059 (N_3059,N_61,N_1231);
nand U3060 (N_3060,N_995,N_2225);
nand U3061 (N_3061,N_1112,N_2343);
or U3062 (N_3062,N_1349,N_1443);
and U3063 (N_3063,N_331,N_896);
or U3064 (N_3064,N_2321,N_818);
or U3065 (N_3065,N_812,N_306);
and U3066 (N_3066,N_2387,N_1459);
nor U3067 (N_3067,N_1187,N_2045);
and U3068 (N_3068,N_1947,N_56);
xnor U3069 (N_3069,N_1927,N_99);
or U3070 (N_3070,N_1695,N_136);
or U3071 (N_3071,N_1655,N_2257);
nor U3072 (N_3072,N_1396,N_1765);
nand U3073 (N_3073,N_2448,N_294);
xnor U3074 (N_3074,N_1589,N_76);
nor U3075 (N_3075,N_2068,N_307);
and U3076 (N_3076,N_1958,N_17);
nand U3077 (N_3077,N_86,N_1282);
or U3078 (N_3078,N_1582,N_2210);
nand U3079 (N_3079,N_2088,N_1575);
nor U3080 (N_3080,N_1178,N_427);
or U3081 (N_3081,N_2005,N_1536);
and U3082 (N_3082,N_1806,N_497);
nor U3083 (N_3083,N_648,N_2468);
or U3084 (N_3084,N_1654,N_3);
nor U3085 (N_3085,N_1356,N_2176);
nand U3086 (N_3086,N_1782,N_1194);
and U3087 (N_3087,N_1685,N_1953);
and U3088 (N_3088,N_1531,N_2475);
and U3089 (N_3089,N_1005,N_2260);
nor U3090 (N_3090,N_1036,N_887);
nand U3091 (N_3091,N_743,N_1139);
nand U3092 (N_3092,N_1916,N_1890);
or U3093 (N_3093,N_1686,N_1105);
or U3094 (N_3094,N_1096,N_978);
and U3095 (N_3095,N_638,N_2125);
and U3096 (N_3096,N_1352,N_2143);
and U3097 (N_3097,N_1802,N_41);
and U3098 (N_3098,N_2489,N_2191);
nand U3099 (N_3099,N_1628,N_1244);
or U3100 (N_3100,N_2160,N_1952);
nor U3101 (N_3101,N_425,N_2377);
xnor U3102 (N_3102,N_2337,N_1988);
or U3103 (N_3103,N_2047,N_187);
or U3104 (N_3104,N_1420,N_2293);
or U3105 (N_3105,N_989,N_592);
and U3106 (N_3106,N_1128,N_867);
nor U3107 (N_3107,N_1072,N_2327);
nand U3108 (N_3108,N_732,N_1800);
and U3109 (N_3109,N_2161,N_124);
and U3110 (N_3110,N_489,N_755);
or U3111 (N_3111,N_345,N_2188);
nand U3112 (N_3112,N_1375,N_1021);
nor U3113 (N_3113,N_1267,N_2141);
or U3114 (N_3114,N_245,N_2436);
and U3115 (N_3115,N_949,N_1716);
nand U3116 (N_3116,N_1486,N_714);
and U3117 (N_3117,N_1425,N_1351);
nand U3118 (N_3118,N_1119,N_1320);
or U3119 (N_3119,N_1056,N_1991);
xnor U3120 (N_3120,N_1336,N_83);
or U3121 (N_3121,N_353,N_1841);
nor U3122 (N_3122,N_1160,N_1394);
or U3123 (N_3123,N_778,N_2057);
nor U3124 (N_3124,N_1593,N_2426);
or U3125 (N_3125,N_152,N_652);
and U3126 (N_3126,N_229,N_762);
nor U3127 (N_3127,N_464,N_1505);
xor U3128 (N_3128,N_1192,N_620);
and U3129 (N_3129,N_1327,N_350);
and U3130 (N_3130,N_808,N_699);
nor U3131 (N_3131,N_1388,N_116);
and U3132 (N_3132,N_1338,N_1826);
and U3133 (N_3133,N_840,N_1501);
nand U3134 (N_3134,N_1314,N_223);
and U3135 (N_3135,N_972,N_1201);
nor U3136 (N_3136,N_2020,N_1797);
xnor U3137 (N_3137,N_1305,N_1339);
nor U3138 (N_3138,N_1039,N_434);
or U3139 (N_3139,N_1675,N_1002);
and U3140 (N_3140,N_2331,N_884);
or U3141 (N_3141,N_1950,N_2109);
or U3142 (N_3142,N_2197,N_649);
or U3143 (N_3143,N_1175,N_2004);
or U3144 (N_3144,N_1666,N_1177);
and U3145 (N_3145,N_2275,N_81);
nor U3146 (N_3146,N_986,N_481);
and U3147 (N_3147,N_824,N_764);
nor U3148 (N_3148,N_598,N_1948);
nand U3149 (N_3149,N_1208,N_1742);
and U3150 (N_3150,N_1962,N_2183);
nand U3151 (N_3151,N_1900,N_525);
nand U3152 (N_3152,N_1381,N_141);
and U3153 (N_3153,N_516,N_1145);
nand U3154 (N_3154,N_498,N_1168);
and U3155 (N_3155,N_7,N_131);
nand U3156 (N_3156,N_263,N_2237);
or U3157 (N_3157,N_1528,N_100);
nor U3158 (N_3158,N_1697,N_1702);
nand U3159 (N_3159,N_119,N_1048);
nand U3160 (N_3160,N_195,N_1880);
nor U3161 (N_3161,N_212,N_1627);
nand U3162 (N_3162,N_134,N_249);
nor U3163 (N_3163,N_1641,N_1312);
and U3164 (N_3164,N_32,N_876);
nand U3165 (N_3165,N_1038,N_2061);
nand U3166 (N_3166,N_2207,N_1426);
and U3167 (N_3167,N_872,N_373);
or U3168 (N_3168,N_951,N_860);
nand U3169 (N_3169,N_934,N_378);
nand U3170 (N_3170,N_2365,N_1721);
and U3171 (N_3171,N_405,N_1225);
nor U3172 (N_3172,N_1821,N_1886);
nor U3173 (N_3173,N_1762,N_1756);
nor U3174 (N_3174,N_2065,N_2029);
nor U3175 (N_3175,N_451,N_75);
and U3176 (N_3176,N_1174,N_2031);
nor U3177 (N_3177,N_1092,N_933);
nand U3178 (N_3178,N_2178,N_1158);
and U3179 (N_3179,N_194,N_1493);
and U3180 (N_3180,N_2105,N_2059);
nor U3181 (N_3181,N_2364,N_383);
nor U3182 (N_3182,N_1412,N_2254);
and U3183 (N_3183,N_1694,N_422);
and U3184 (N_3184,N_1196,N_614);
nand U3185 (N_3185,N_250,N_2036);
nor U3186 (N_3186,N_2277,N_1126);
and U3187 (N_3187,N_2037,N_2303);
or U3188 (N_3188,N_664,N_1209);
and U3189 (N_3189,N_2096,N_390);
or U3190 (N_3190,N_416,N_1684);
xor U3191 (N_3191,N_333,N_114);
and U3192 (N_3192,N_1969,N_2413);
nor U3193 (N_3193,N_2329,N_1795);
or U3194 (N_3194,N_1377,N_417);
and U3195 (N_3195,N_367,N_1461);
xnor U3196 (N_3196,N_400,N_105);
nand U3197 (N_3197,N_2179,N_1323);
or U3198 (N_3198,N_875,N_2322);
xor U3199 (N_3199,N_795,N_1019);
and U3200 (N_3200,N_667,N_865);
nand U3201 (N_3201,N_2108,N_1584);
or U3202 (N_3202,N_722,N_358);
or U3203 (N_3203,N_1383,N_1770);
nor U3204 (N_3204,N_1071,N_983);
and U3205 (N_3205,N_562,N_748);
nor U3206 (N_3206,N_1470,N_2393);
nor U3207 (N_3207,N_698,N_2079);
or U3208 (N_3208,N_2042,N_2126);
or U3209 (N_3209,N_1273,N_552);
and U3210 (N_3210,N_351,N_1441);
and U3211 (N_3211,N_1350,N_943);
nor U3212 (N_3212,N_1221,N_2107);
nor U3213 (N_3213,N_2320,N_402);
or U3214 (N_3214,N_2222,N_339);
and U3215 (N_3215,N_1270,N_2480);
nand U3216 (N_3216,N_1611,N_1838);
xnor U3217 (N_3217,N_1184,N_2432);
or U3218 (N_3218,N_952,N_1817);
nor U3219 (N_3219,N_1975,N_2193);
xor U3220 (N_3220,N_1416,N_616);
nor U3221 (N_3221,N_568,N_1515);
or U3222 (N_3222,N_1032,N_1936);
nor U3223 (N_3223,N_2386,N_2256);
or U3224 (N_3224,N_1251,N_1276);
or U3225 (N_3225,N_2262,N_928);
nand U3226 (N_3226,N_2066,N_438);
or U3227 (N_3227,N_2085,N_2024);
or U3228 (N_3228,N_322,N_1822);
nand U3229 (N_3229,N_1642,N_207);
and U3230 (N_3230,N_1073,N_1731);
and U3231 (N_3231,N_1639,N_833);
nand U3232 (N_3232,N_1161,N_1080);
xor U3233 (N_3233,N_1798,N_1787);
or U3234 (N_3234,N_1633,N_1587);
or U3235 (N_3235,N_1147,N_1274);
nand U3236 (N_3236,N_1723,N_2015);
or U3237 (N_3237,N_967,N_1818);
and U3238 (N_3238,N_2379,N_521);
nand U3239 (N_3239,N_1261,N_1228);
and U3240 (N_3240,N_1077,N_1135);
nand U3241 (N_3241,N_404,N_1712);
nand U3242 (N_3242,N_557,N_852);
xor U3243 (N_3243,N_710,N_2184);
nor U3244 (N_3244,N_2016,N_1941);
or U3245 (N_3245,N_1195,N_2072);
or U3246 (N_3246,N_1605,N_854);
and U3247 (N_3247,N_1545,N_2216);
nor U3248 (N_3248,N_677,N_2221);
and U3249 (N_3249,N_336,N_55);
xor U3250 (N_3250,N_784,N_1744);
nand U3251 (N_3251,N_459,N_1512);
nand U3252 (N_3252,N_2391,N_436);
or U3253 (N_3253,N_1491,N_2241);
xor U3254 (N_3254,N_561,N_1730);
or U3255 (N_3255,N_421,N_1542);
and U3256 (N_3256,N_2496,N_150);
or U3257 (N_3257,N_20,N_1057);
nor U3258 (N_3258,N_1165,N_2401);
nor U3259 (N_3259,N_1059,N_668);
nor U3260 (N_3260,N_997,N_1366);
nand U3261 (N_3261,N_1912,N_77);
nor U3262 (N_3262,N_821,N_2491);
and U3263 (N_3263,N_926,N_800);
and U3264 (N_3264,N_798,N_1849);
or U3265 (N_3265,N_2449,N_1599);
nor U3266 (N_3266,N_1828,N_2412);
or U3267 (N_3267,N_1711,N_2008);
or U3268 (N_3268,N_222,N_927);
nor U3269 (N_3269,N_1769,N_58);
nor U3270 (N_3270,N_40,N_2429);
or U3271 (N_3271,N_963,N_740);
nor U3272 (N_3272,N_1526,N_671);
nor U3273 (N_3273,N_2419,N_2129);
nor U3274 (N_3274,N_631,N_2080);
or U3275 (N_3275,N_1908,N_201);
or U3276 (N_3276,N_964,N_27);
nand U3277 (N_3277,N_810,N_104);
nor U3278 (N_3278,N_171,N_1357);
or U3279 (N_3279,N_213,N_1976);
xnor U3280 (N_3280,N_468,N_672);
or U3281 (N_3281,N_1547,N_1287);
xnor U3282 (N_3282,N_2133,N_1249);
and U3283 (N_3283,N_5,N_538);
nand U3284 (N_3284,N_687,N_627);
and U3285 (N_3285,N_692,N_716);
nand U3286 (N_3286,N_1410,N_2264);
nor U3287 (N_3287,N_143,N_630);
and U3288 (N_3288,N_1011,N_2443);
and U3289 (N_3289,N_1507,N_2255);
nand U3290 (N_3290,N_230,N_728);
nor U3291 (N_3291,N_2445,N_960);
or U3292 (N_3292,N_1324,N_363);
and U3293 (N_3293,N_615,N_1035);
and U3294 (N_3294,N_957,N_688);
or U3295 (N_3295,N_1137,N_931);
nand U3296 (N_3296,N_1663,N_673);
nor U3297 (N_3297,N_22,N_1874);
and U3298 (N_3298,N_801,N_1253);
xor U3299 (N_3299,N_1579,N_2171);
nor U3300 (N_3300,N_814,N_721);
or U3301 (N_3301,N_1013,N_2242);
or U3302 (N_3302,N_1757,N_1981);
nor U3303 (N_3303,N_2218,N_2136);
nor U3304 (N_3304,N_246,N_1023);
nor U3305 (N_3305,N_92,N_2230);
and U3306 (N_3306,N_835,N_155);
and U3307 (N_3307,N_2093,N_754);
and U3308 (N_3308,N_2187,N_580);
and U3309 (N_3309,N_1538,N_2170);
nand U3310 (N_3310,N_916,N_332);
nor U3311 (N_3311,N_1468,N_444);
xor U3312 (N_3312,N_803,N_89);
nand U3313 (N_3313,N_1517,N_1417);
or U3314 (N_3314,N_128,N_1144);
nor U3315 (N_3315,N_759,N_1929);
nor U3316 (N_3316,N_1151,N_372);
nand U3317 (N_3317,N_2181,N_1596);
and U3318 (N_3318,N_528,N_1867);
xnor U3319 (N_3319,N_1743,N_2021);
xor U3320 (N_3320,N_2398,N_582);
and U3321 (N_3321,N_567,N_278);
and U3322 (N_3322,N_505,N_1321);
and U3323 (N_3323,N_2123,N_799);
and U3324 (N_3324,N_1651,N_946);
and U3325 (N_3325,N_817,N_2146);
or U3326 (N_3326,N_443,N_386);
and U3327 (N_3327,N_63,N_862);
nor U3328 (N_3328,N_2116,N_288);
or U3329 (N_3329,N_2458,N_1671);
nor U3330 (N_3330,N_2481,N_556);
or U3331 (N_3331,N_861,N_1669);
nor U3332 (N_3332,N_1223,N_1472);
nor U3333 (N_3333,N_1732,N_522);
nor U3334 (N_3334,N_209,N_1994);
nand U3335 (N_3335,N_1404,N_1311);
nor U3336 (N_3336,N_441,N_1476);
xor U3337 (N_3337,N_2238,N_1664);
nor U3338 (N_3338,N_921,N_877);
or U3339 (N_3339,N_2339,N_956);
or U3340 (N_3340,N_1212,N_720);
and U3341 (N_3341,N_186,N_903);
nor U3342 (N_3342,N_1418,N_1331);
or U3343 (N_3343,N_1095,N_167);
and U3344 (N_3344,N_1391,N_2113);
nand U3345 (N_3345,N_2307,N_549);
nand U3346 (N_3346,N_2182,N_2380);
or U3347 (N_3347,N_1197,N_2086);
and U3348 (N_3348,N_1329,N_2253);
or U3349 (N_3349,N_682,N_1576);
nor U3350 (N_3350,N_1704,N_515);
or U3351 (N_3351,N_1254,N_666);
nor U3352 (N_3352,N_2456,N_1919);
nor U3353 (N_3353,N_536,N_502);
nor U3354 (N_3354,N_1617,N_415);
and U3355 (N_3355,N_707,N_2332);
or U3356 (N_3356,N_1376,N_360);
or U3357 (N_3357,N_680,N_2282);
xor U3358 (N_3358,N_1384,N_462);
or U3359 (N_3359,N_689,N_1548);
nand U3360 (N_3360,N_1774,N_1662);
or U3361 (N_3361,N_1233,N_1961);
xor U3362 (N_3362,N_540,N_344);
or U3363 (N_3363,N_1870,N_2457);
xnor U3364 (N_3364,N_69,N_2158);
nand U3365 (N_3365,N_1386,N_1804);
or U3366 (N_3366,N_975,N_2318);
and U3367 (N_3367,N_979,N_117);
xor U3368 (N_3368,N_118,N_1692);
nand U3369 (N_3369,N_2424,N_1758);
or U3370 (N_3370,N_1189,N_191);
nand U3371 (N_3371,N_1672,N_414);
nor U3372 (N_3372,N_2095,N_1523);
or U3373 (N_3373,N_165,N_1094);
or U3374 (N_3374,N_773,N_2200);
or U3375 (N_3375,N_686,N_709);
nand U3376 (N_3376,N_1257,N_111);
and U3377 (N_3377,N_2102,N_2336);
nor U3378 (N_3378,N_1222,N_1535);
xnor U3379 (N_3379,N_853,N_13);
or U3380 (N_3380,N_2258,N_1949);
xnor U3381 (N_3381,N_2482,N_412);
and U3382 (N_3382,N_508,N_1090);
nor U3383 (N_3383,N_1616,N_2043);
xnor U3384 (N_3384,N_12,N_1136);
nor U3385 (N_3385,N_1552,N_208);
or U3386 (N_3386,N_591,N_2009);
or U3387 (N_3387,N_1500,N_1401);
and U3388 (N_3388,N_282,N_628);
nand U3389 (N_3389,N_1753,N_1741);
nor U3390 (N_3390,N_772,N_1027);
and U3391 (N_3391,N_1759,N_312);
or U3392 (N_3392,N_1944,N_1650);
and U3393 (N_3393,N_1141,N_2410);
nand U3394 (N_3394,N_1262,N_2417);
nand U3395 (N_3395,N_988,N_1863);
nand U3396 (N_3396,N_572,N_1746);
and U3397 (N_3397,N_2373,N_1567);
nor U3398 (N_3398,N_1462,N_1364);
or U3399 (N_3399,N_379,N_696);
xor U3400 (N_3400,N_1138,N_1216);
nor U3401 (N_3401,N_1646,N_2050);
or U3402 (N_3402,N_1703,N_491);
or U3403 (N_3403,N_31,N_2083);
and U3404 (N_3404,N_298,N_1230);
xor U3405 (N_3405,N_738,N_1133);
nand U3406 (N_3406,N_881,N_1659);
or U3407 (N_3407,N_478,N_2013);
and U3408 (N_3408,N_1315,N_629);
xor U3409 (N_3409,N_763,N_1017);
nand U3410 (N_3410,N_280,N_878);
nor U3411 (N_3411,N_685,N_2433);
nand U3412 (N_3412,N_1236,N_1382);
or U3413 (N_3413,N_1123,N_1845);
or U3414 (N_3414,N_2440,N_1630);
and U3415 (N_3415,N_1932,N_1864);
nor U3416 (N_3416,N_1556,N_914);
nand U3417 (N_3417,N_534,N_1076);
and U3418 (N_3418,N_700,N_1299);
or U3419 (N_3419,N_533,N_1602);
nor U3420 (N_3420,N_1219,N_1625);
nor U3421 (N_3421,N_342,N_1428);
or U3422 (N_3422,N_192,N_2112);
xor U3423 (N_3423,N_2294,N_1453);
nor U3424 (N_3424,N_1214,N_1181);
nand U3425 (N_3425,N_837,N_1322);
or U3426 (N_3426,N_255,N_711);
or U3427 (N_3427,N_1788,N_1615);
nand U3428 (N_3428,N_1466,N_228);
and U3429 (N_3429,N_1881,N_639);
nor U3430 (N_3430,N_385,N_1068);
or U3431 (N_3431,N_1387,N_2151);
or U3432 (N_3432,N_929,N_583);
and U3433 (N_3433,N_323,N_611);
nand U3434 (N_3434,N_1985,N_780);
or U3435 (N_3435,N_915,N_1645);
xnor U3436 (N_3436,N_2328,N_1899);
and U3437 (N_3437,N_2362,N_1280);
nor U3438 (N_3438,N_1291,N_1149);
or U3439 (N_3439,N_1768,N_1292);
nor U3440 (N_3440,N_1485,N_1044);
nand U3441 (N_3441,N_2147,N_514);
or U3442 (N_3442,N_558,N_1931);
nand U3443 (N_3443,N_1683,N_2334);
and U3444 (N_3444,N_2223,N_226);
and U3445 (N_3445,N_1558,N_2431);
and U3446 (N_3446,N_1609,N_1829);
or U3447 (N_3447,N_831,N_28);
or U3448 (N_3448,N_681,N_1087);
xnor U3449 (N_3449,N_176,N_1831);
nor U3450 (N_3450,N_782,N_184);
or U3451 (N_3451,N_792,N_1081);
or U3452 (N_3452,N_2471,N_1109);
or U3453 (N_3453,N_1457,N_548);
nand U3454 (N_3454,N_1997,N_2131);
nand U3455 (N_3455,N_21,N_2335);
xor U3456 (N_3456,N_1421,N_1661);
or U3457 (N_3457,N_113,N_674);
nor U3458 (N_3458,N_2311,N_2323);
and U3459 (N_3459,N_161,N_2162);
nand U3460 (N_3460,N_1973,N_166);
nand U3461 (N_3461,N_545,N_1751);
nor U3462 (N_3462,N_1079,N_450);
or U3463 (N_3463,N_2400,N_225);
xor U3464 (N_3464,N_1344,N_2418);
and U3465 (N_3465,N_725,N_335);
or U3466 (N_3466,N_57,N_6);
xor U3467 (N_3467,N_742,N_2266);
nor U3468 (N_3468,N_1016,N_1186);
nand U3469 (N_3469,N_14,N_1343);
xnor U3470 (N_3470,N_1827,N_2163);
nor U3471 (N_3471,N_2423,N_1060);
or U3472 (N_3472,N_376,N_747);
xnor U3473 (N_3473,N_990,N_1771);
nor U3474 (N_3474,N_2414,N_1848);
nor U3475 (N_3475,N_697,N_1873);
and U3476 (N_3476,N_1089,N_802);
nor U3477 (N_3477,N_2404,N_588);
xnor U3478 (N_3478,N_735,N_2469);
nor U3479 (N_3479,N_1903,N_1374);
and U3480 (N_3480,N_650,N_560);
and U3481 (N_3481,N_1846,N_2450);
nor U3482 (N_3482,N_108,N_961);
nor U3483 (N_3483,N_2370,N_1937);
or U3484 (N_3484,N_1372,N_1499);
nand U3485 (N_3485,N_2273,N_1328);
or U3486 (N_3486,N_520,N_1306);
nor U3487 (N_3487,N_917,N_266);
nor U3488 (N_3488,N_341,N_348);
or U3489 (N_3489,N_2053,N_271);
or U3490 (N_3490,N_1379,N_1275);
nor U3491 (N_3491,N_768,N_550);
nand U3492 (N_3492,N_123,N_2094);
nand U3493 (N_3493,N_2248,N_59);
nand U3494 (N_3494,N_2075,N_2312);
and U3495 (N_3495,N_1085,N_67);
and U3496 (N_3496,N_2268,N_418);
nor U3497 (N_3497,N_147,N_578);
or U3498 (N_3498,N_122,N_1996);
and U3499 (N_3499,N_2019,N_879);
xnor U3500 (N_3500,N_1463,N_1808);
and U3501 (N_3501,N_2326,N_1856);
xor U3502 (N_3502,N_2164,N_1363);
nand U3503 (N_3503,N_1851,N_834);
nand U3504 (N_3504,N_959,N_1084);
nor U3505 (N_3505,N_396,N_1337);
or U3506 (N_3506,N_1,N_1442);
or U3507 (N_3507,N_633,N_1614);
nand U3508 (N_3508,N_1911,N_2023);
nor U3509 (N_3509,N_1370,N_2350);
and U3510 (N_3510,N_1549,N_969);
xor U3511 (N_3511,N_820,N_34);
xor U3512 (N_3512,N_189,N_303);
nand U3513 (N_3513,N_901,N_1891);
nor U3514 (N_3514,N_2288,N_210);
nor U3515 (N_3515,N_2052,N_2315);
xnor U3516 (N_3516,N_2483,N_2415);
and U3517 (N_3517,N_238,N_1010);
and U3518 (N_3518,N_1392,N_1876);
or U3519 (N_3519,N_992,N_2403);
and U3520 (N_3520,N_958,N_874);
or U3521 (N_3521,N_1649,N_4);
or U3522 (N_3522,N_2283,N_1288);
xor U3523 (N_3523,N_895,N_994);
nor U3524 (N_3524,N_660,N_2142);
nand U3525 (N_3525,N_1781,N_1435);
nor U3526 (N_3526,N_1888,N_1696);
xor U3527 (N_3527,N_1978,N_173);
nor U3528 (N_3528,N_1260,N_1114);
nand U3529 (N_3529,N_1710,N_1250);
nand U3530 (N_3530,N_832,N_1263);
and U3531 (N_3531,N_2217,N_539);
or U3532 (N_3532,N_771,N_1897);
or U3533 (N_3533,N_1533,N_338);
xor U3534 (N_3534,N_619,N_1665);
or U3535 (N_3535,N_2041,N_352);
nand U3536 (N_3536,N_1745,N_1125);
and U3537 (N_3537,N_885,N_2006);
and U3538 (N_3538,N_133,N_600);
or U3539 (N_3539,N_2425,N_2165);
nor U3540 (N_3540,N_2279,N_563);
xor U3541 (N_3541,N_1830,N_541);
nor U3542 (N_3542,N_2224,N_1667);
and U3543 (N_3543,N_224,N_544);
or U3544 (N_3544,N_2470,N_1047);
xor U3545 (N_3545,N_1674,N_1729);
nor U3546 (N_3546,N_2058,N_1317);
nand U3547 (N_3547,N_823,N_380);
or U3548 (N_3548,N_48,N_2084);
and U3549 (N_3549,N_2089,N_1191);
nor U3550 (N_3550,N_982,N_2388);
or U3551 (N_3551,N_1206,N_1546);
or U3552 (N_3552,N_1482,N_1307);
and U3553 (N_3553,N_1508,N_1483);
nand U3554 (N_3554,N_980,N_804);
and U3555 (N_3555,N_125,N_1987);
or U3556 (N_3556,N_153,N_2000);
nand U3557 (N_3557,N_2389,N_1101);
nand U3558 (N_3558,N_610,N_1883);
and U3559 (N_3559,N_217,N_621);
nand U3560 (N_3560,N_2474,N_2399);
or U3561 (N_3561,N_180,N_2271);
nor U3562 (N_3562,N_193,N_690);
nor U3563 (N_3563,N_2287,N_1373);
and U3564 (N_3564,N_33,N_2208);
nand U3565 (N_3565,N_499,N_1506);
and U3566 (N_3566,N_1803,N_1877);
and U3567 (N_3567,N_1226,N_139);
or U3568 (N_3568,N_2361,N_1495);
nand U3569 (N_3569,N_1578,N_2204);
nand U3570 (N_3570,N_296,N_310);
nand U3571 (N_3571,N_1647,N_585);
and U3572 (N_3572,N_1678,N_2051);
or U3573 (N_3573,N_452,N_2479);
nand U3574 (N_3574,N_1211,N_1566);
or U3575 (N_3575,N_2078,N_1182);
nand U3576 (N_3576,N_449,N_1475);
or U3577 (N_3577,N_73,N_547);
xnor U3578 (N_3578,N_1513,N_1610);
nand U3579 (N_3579,N_573,N_1866);
xor U3580 (N_3580,N_1489,N_1980);
or U3581 (N_3581,N_1051,N_1832);
nand U3582 (N_3582,N_2044,N_393);
nand U3583 (N_3583,N_244,N_1368);
or U3584 (N_3584,N_1353,N_292);
nor U3585 (N_3585,N_1979,N_227);
or U3586 (N_3586,N_976,N_1726);
nand U3587 (N_3587,N_894,N_2121);
or U3588 (N_3588,N_175,N_1893);
or U3589 (N_3589,N_1543,N_701);
nand U3590 (N_3590,N_1205,N_2154);
or U3591 (N_3591,N_889,N_1850);
or U3592 (N_3592,N_1792,N_1419);
nand U3593 (N_3593,N_2465,N_2492);
and U3594 (N_3594,N_49,N_661);
nand U3595 (N_3595,N_493,N_937);
nor U3596 (N_3596,N_2214,N_1825);
nand U3597 (N_3597,N_2317,N_1243);
and U3598 (N_3598,N_2352,N_1029);
or U3599 (N_3599,N_39,N_500);
xor U3600 (N_3600,N_279,N_2358);
or U3601 (N_3601,N_1600,N_101);
nor U3602 (N_3602,N_1445,N_1183);
nor U3603 (N_3603,N_899,N_1385);
nand U3604 (N_3604,N_2437,N_1259);
nor U3605 (N_3605,N_841,N_1163);
nand U3606 (N_3606,N_1859,N_1794);
and U3607 (N_3607,N_1361,N_1063);
nor U3608 (N_3608,N_603,N_2090);
or U3609 (N_3609,N_1601,N_431);
nand U3610 (N_3610,N_1780,N_1166);
and U3611 (N_3611,N_2462,N_938);
nor U3612 (N_3612,N_1879,N_641);
nor U3613 (N_3613,N_745,N_793);
nor U3614 (N_3614,N_1180,N_1569);
nand U3615 (N_3615,N_2298,N_1448);
nor U3616 (N_3616,N_359,N_2409);
and U3617 (N_3617,N_1608,N_1204);
nand U3618 (N_3618,N_1400,N_2466);
nand U3619 (N_3619,N_1778,N_913);
nand U3620 (N_3620,N_1913,N_1473);
xnor U3621 (N_3621,N_1577,N_2166);
and U3622 (N_3622,N_1612,N_384);
or U3623 (N_3623,N_858,N_1638);
xnor U3624 (N_3624,N_1564,N_2130);
nand U3625 (N_3625,N_1066,N_85);
and U3626 (N_3626,N_1097,N_362);
and U3627 (N_3627,N_2003,N_965);
and U3628 (N_3628,N_18,N_1509);
or U3629 (N_3629,N_753,N_1544);
nor U3630 (N_3630,N_90,N_1520);
or U3631 (N_3631,N_1679,N_1497);
and U3632 (N_3632,N_1813,N_2076);
nor U3633 (N_3633,N_1522,N_381);
xnor U3634 (N_3634,N_42,N_1540);
nor U3635 (N_3635,N_1098,N_2017);
or U3636 (N_3636,N_1835,N_662);
and U3637 (N_3637,N_2435,N_783);
or U3638 (N_3638,N_2407,N_1402);
nor U3639 (N_3639,N_2049,N_1067);
xor U3640 (N_3640,N_1855,N_1033);
xnor U3641 (N_3641,N_1430,N_2292);
or U3642 (N_3642,N_234,N_1852);
or U3643 (N_3643,N_2150,N_1573);
or U3644 (N_3644,N_455,N_1217);
nor U3645 (N_3645,N_2077,N_2128);
nor U3646 (N_3646,N_270,N_1917);
nor U3647 (N_3647,N_0,N_369);
nor U3648 (N_3648,N_11,N_2201);
nor U3649 (N_3649,N_1904,N_1918);
nor U3650 (N_3650,N_202,N_356);
or U3651 (N_3651,N_811,N_2038);
or U3652 (N_3652,N_704,N_1162);
or U3653 (N_3653,N_907,N_1885);
or U3654 (N_3654,N_25,N_265);
nand U3655 (N_3655,N_1598,N_2138);
and U3656 (N_3656,N_261,N_423);
nor U3657 (N_3657,N_1190,N_1858);
and U3658 (N_3658,N_1046,N_446);
nor U3659 (N_3659,N_897,N_2110);
and U3660 (N_3660,N_1188,N_9);
or U3661 (N_3661,N_1200,N_749);
and U3662 (N_3662,N_713,N_947);
xor U3663 (N_3663,N_1820,N_2291);
nor U3664 (N_3664,N_121,N_80);
xor U3665 (N_3665,N_845,N_923);
and U3666 (N_3666,N_596,N_236);
nand U3667 (N_3667,N_2324,N_1984);
and U3668 (N_3668,N_474,N_2473);
and U3669 (N_3669,N_1809,N_779);
nand U3670 (N_3670,N_2155,N_746);
nand U3671 (N_3671,N_2251,N_1887);
or U3672 (N_3672,N_2439,N_1555);
and U3673 (N_3673,N_787,N_1907);
nand U3674 (N_3674,N_366,N_1118);
or U3675 (N_3675,N_72,N_1844);
nor U3676 (N_3676,N_1478,N_1193);
xnor U3677 (N_3677,N_1631,N_2226);
and U3678 (N_3678,N_2239,N_445);
nand U3679 (N_3679,N_1099,N_138);
or U3680 (N_3680,N_2488,N_930);
or U3681 (N_3681,N_1925,N_1104);
nor U3682 (N_3682,N_1301,N_142);
nor U3683 (N_3683,N_197,N_1811);
nor U3684 (N_3684,N_1269,N_354);
and U3685 (N_3685,N_1365,N_2269);
and U3686 (N_3686,N_145,N_1438);
and U3687 (N_3687,N_1018,N_790);
nor U3688 (N_3688,N_1940,N_2375);
nand U3689 (N_3689,N_1203,N_1348);
nor U3690 (N_3690,N_599,N_601);
nand U3691 (N_3691,N_1346,N_2333);
nor U3692 (N_3692,N_501,N_2135);
and U3693 (N_3693,N_576,N_839);
xnor U3694 (N_3694,N_2060,N_2330);
or U3695 (N_3695,N_1502,N_757);
or U3696 (N_3696,N_2346,N_2202);
nor U3697 (N_3697,N_1398,N_1572);
nand U3698 (N_3698,N_2132,N_1399);
nand U3699 (N_3699,N_2300,N_1530);
and U3700 (N_3700,N_777,N_962);
nand U3701 (N_3701,N_291,N_492);
nand U3702 (N_3702,N_2452,N_2001);
nand U3703 (N_3703,N_102,N_2442);
nor U3704 (N_3704,N_727,N_1026);
nor U3705 (N_3705,N_2234,N_2382);
nor U3706 (N_3706,N_890,N_676);
or U3707 (N_3707,N_1446,N_471);
nand U3708 (N_3708,N_364,N_1514);
xor U3709 (N_3709,N_2040,N_65);
or U3710 (N_3710,N_454,N_1108);
nor U3711 (N_3711,N_2026,N_1237);
nor U3712 (N_3712,N_1454,N_912);
nor U3713 (N_3713,N_2111,N_317);
nand U3714 (N_3714,N_617,N_1433);
or U3715 (N_3715,N_825,N_1129);
nor U3716 (N_3716,N_791,N_850);
or U3717 (N_3717,N_1793,N_327);
nand U3718 (N_3718,N_1964,N_2034);
nor U3719 (N_3719,N_174,N_1860);
nand U3720 (N_3720,N_71,N_1992);
and U3721 (N_3721,N_2030,N_2265);
nand U3722 (N_3722,N_2156,N_1656);
or U3723 (N_3723,N_46,N_2341);
nor U3724 (N_3724,N_1103,N_925);
nand U3725 (N_3725,N_1560,N_1624);
nand U3726 (N_3726,N_395,N_2384);
or U3727 (N_3727,N_365,N_1006);
nand U3728 (N_3728,N_91,N_1266);
nand U3729 (N_3729,N_1054,N_2368);
and U3730 (N_3730,N_670,N_2046);
and U3731 (N_3731,N_1719,N_1061);
or U3732 (N_3732,N_269,N_736);
or U3733 (N_3733,N_2209,N_2070);
nor U3734 (N_3734,N_1326,N_1340);
nand U3735 (N_3735,N_419,N_78);
or U3736 (N_3736,N_2190,N_737);
nor U3737 (N_3737,N_726,N_1955);
or U3738 (N_3738,N_1296,N_120);
xor U3739 (N_3739,N_1325,N_1131);
nor U3740 (N_3740,N_2148,N_971);
or U3741 (N_3741,N_51,N_1342);
or U3742 (N_3742,N_1132,N_181);
nor U3743 (N_3743,N_1812,N_636);
nor U3744 (N_3744,N_2363,N_1049);
nand U3745 (N_3745,N_1597,N_237);
nand U3746 (N_3746,N_1258,N_1272);
nand U3747 (N_3747,N_1905,N_1423);
nand U3748 (N_3748,N_1691,N_2397);
or U3749 (N_3749,N_1172,N_2122);
xnor U3750 (N_3750,N_474,N_329);
and U3751 (N_3751,N_183,N_543);
nor U3752 (N_3752,N_684,N_22);
nand U3753 (N_3753,N_1435,N_714);
nor U3754 (N_3754,N_819,N_902);
or U3755 (N_3755,N_334,N_1842);
nand U3756 (N_3756,N_1915,N_129);
nor U3757 (N_3757,N_1729,N_770);
and U3758 (N_3758,N_364,N_1397);
nand U3759 (N_3759,N_2023,N_482);
nor U3760 (N_3760,N_1125,N_1598);
nand U3761 (N_3761,N_372,N_2224);
and U3762 (N_3762,N_2205,N_633);
and U3763 (N_3763,N_771,N_904);
or U3764 (N_3764,N_399,N_349);
nand U3765 (N_3765,N_52,N_988);
and U3766 (N_3766,N_806,N_251);
nor U3767 (N_3767,N_1676,N_1973);
nand U3768 (N_3768,N_2085,N_2475);
nor U3769 (N_3769,N_926,N_733);
nor U3770 (N_3770,N_2246,N_1926);
and U3771 (N_3771,N_1145,N_830);
or U3772 (N_3772,N_2474,N_1946);
nor U3773 (N_3773,N_790,N_73);
and U3774 (N_3774,N_2015,N_1284);
and U3775 (N_3775,N_704,N_2377);
or U3776 (N_3776,N_1987,N_501);
and U3777 (N_3777,N_2140,N_760);
and U3778 (N_3778,N_755,N_205);
xor U3779 (N_3779,N_2418,N_2059);
nor U3780 (N_3780,N_2270,N_2344);
xor U3781 (N_3781,N_1936,N_1019);
xor U3782 (N_3782,N_1140,N_1053);
or U3783 (N_3783,N_144,N_889);
and U3784 (N_3784,N_1387,N_1095);
or U3785 (N_3785,N_696,N_482);
nand U3786 (N_3786,N_1459,N_1117);
nand U3787 (N_3787,N_1317,N_1943);
nand U3788 (N_3788,N_12,N_2219);
nor U3789 (N_3789,N_218,N_2477);
nor U3790 (N_3790,N_795,N_1218);
nand U3791 (N_3791,N_1657,N_2044);
and U3792 (N_3792,N_1041,N_259);
and U3793 (N_3793,N_1565,N_1709);
nor U3794 (N_3794,N_1958,N_179);
and U3795 (N_3795,N_767,N_231);
and U3796 (N_3796,N_1623,N_161);
and U3797 (N_3797,N_2313,N_898);
nand U3798 (N_3798,N_1885,N_131);
nand U3799 (N_3799,N_2427,N_209);
nor U3800 (N_3800,N_1712,N_1390);
nor U3801 (N_3801,N_2353,N_641);
and U3802 (N_3802,N_960,N_2148);
and U3803 (N_3803,N_545,N_346);
nor U3804 (N_3804,N_430,N_1928);
nor U3805 (N_3805,N_1668,N_1216);
or U3806 (N_3806,N_812,N_1959);
xnor U3807 (N_3807,N_1903,N_1124);
and U3808 (N_3808,N_1249,N_2459);
or U3809 (N_3809,N_230,N_2217);
and U3810 (N_3810,N_1511,N_892);
and U3811 (N_3811,N_1066,N_673);
nor U3812 (N_3812,N_1115,N_1331);
or U3813 (N_3813,N_720,N_1064);
and U3814 (N_3814,N_2069,N_1266);
xnor U3815 (N_3815,N_1861,N_1953);
and U3816 (N_3816,N_2142,N_1911);
nand U3817 (N_3817,N_2471,N_1835);
xor U3818 (N_3818,N_2179,N_394);
xor U3819 (N_3819,N_2446,N_1154);
xor U3820 (N_3820,N_1403,N_1226);
or U3821 (N_3821,N_2006,N_1619);
nor U3822 (N_3822,N_972,N_1763);
or U3823 (N_3823,N_7,N_1231);
or U3824 (N_3824,N_80,N_504);
and U3825 (N_3825,N_883,N_1145);
nor U3826 (N_3826,N_2253,N_1168);
and U3827 (N_3827,N_1214,N_1945);
nand U3828 (N_3828,N_127,N_296);
nor U3829 (N_3829,N_2251,N_1465);
nor U3830 (N_3830,N_519,N_2109);
nand U3831 (N_3831,N_2334,N_1844);
xnor U3832 (N_3832,N_601,N_1854);
xnor U3833 (N_3833,N_2237,N_1339);
nor U3834 (N_3834,N_442,N_380);
or U3835 (N_3835,N_663,N_1394);
xor U3836 (N_3836,N_2333,N_274);
nor U3837 (N_3837,N_717,N_1460);
nand U3838 (N_3838,N_610,N_991);
and U3839 (N_3839,N_1599,N_911);
or U3840 (N_3840,N_2413,N_1195);
nor U3841 (N_3841,N_983,N_1487);
and U3842 (N_3842,N_420,N_2453);
and U3843 (N_3843,N_969,N_1092);
or U3844 (N_3844,N_996,N_40);
xor U3845 (N_3845,N_1776,N_276);
nand U3846 (N_3846,N_279,N_801);
xor U3847 (N_3847,N_1192,N_2307);
nand U3848 (N_3848,N_1165,N_20);
nor U3849 (N_3849,N_1398,N_50);
nand U3850 (N_3850,N_11,N_210);
or U3851 (N_3851,N_378,N_1117);
nand U3852 (N_3852,N_840,N_1677);
nor U3853 (N_3853,N_991,N_1008);
xor U3854 (N_3854,N_1180,N_765);
or U3855 (N_3855,N_194,N_2349);
and U3856 (N_3856,N_2036,N_1628);
or U3857 (N_3857,N_1777,N_1913);
or U3858 (N_3858,N_1293,N_1040);
and U3859 (N_3859,N_514,N_1842);
nor U3860 (N_3860,N_1802,N_520);
or U3861 (N_3861,N_58,N_493);
and U3862 (N_3862,N_2457,N_1112);
nand U3863 (N_3863,N_1479,N_464);
and U3864 (N_3864,N_1213,N_1476);
nand U3865 (N_3865,N_54,N_95);
or U3866 (N_3866,N_401,N_592);
or U3867 (N_3867,N_677,N_972);
nor U3868 (N_3868,N_680,N_2385);
and U3869 (N_3869,N_1353,N_1594);
xor U3870 (N_3870,N_1015,N_49);
nor U3871 (N_3871,N_1110,N_944);
or U3872 (N_3872,N_1311,N_409);
nand U3873 (N_3873,N_2268,N_433);
or U3874 (N_3874,N_1081,N_1599);
and U3875 (N_3875,N_175,N_1328);
xor U3876 (N_3876,N_2447,N_1419);
or U3877 (N_3877,N_213,N_1180);
and U3878 (N_3878,N_208,N_986);
and U3879 (N_3879,N_2174,N_262);
nand U3880 (N_3880,N_1920,N_56);
and U3881 (N_3881,N_395,N_912);
nor U3882 (N_3882,N_257,N_1944);
nor U3883 (N_3883,N_1529,N_1749);
nor U3884 (N_3884,N_2157,N_2127);
xor U3885 (N_3885,N_1335,N_1537);
xor U3886 (N_3886,N_2092,N_604);
and U3887 (N_3887,N_230,N_130);
nand U3888 (N_3888,N_2077,N_702);
and U3889 (N_3889,N_801,N_1911);
nand U3890 (N_3890,N_173,N_1834);
nor U3891 (N_3891,N_1699,N_1758);
nand U3892 (N_3892,N_2215,N_1296);
and U3893 (N_3893,N_1128,N_2389);
and U3894 (N_3894,N_409,N_2424);
nor U3895 (N_3895,N_1255,N_133);
nor U3896 (N_3896,N_2200,N_1033);
or U3897 (N_3897,N_82,N_792);
nand U3898 (N_3898,N_307,N_1328);
or U3899 (N_3899,N_567,N_1869);
nor U3900 (N_3900,N_878,N_807);
and U3901 (N_3901,N_1790,N_2338);
or U3902 (N_3902,N_2081,N_988);
or U3903 (N_3903,N_789,N_393);
nor U3904 (N_3904,N_2072,N_2383);
nor U3905 (N_3905,N_1008,N_1707);
nor U3906 (N_3906,N_1660,N_786);
xnor U3907 (N_3907,N_2128,N_1466);
or U3908 (N_3908,N_812,N_1611);
nand U3909 (N_3909,N_1263,N_884);
or U3910 (N_3910,N_1966,N_1231);
nor U3911 (N_3911,N_1881,N_2045);
or U3912 (N_3912,N_1670,N_2369);
and U3913 (N_3913,N_2165,N_2256);
nor U3914 (N_3914,N_2495,N_440);
and U3915 (N_3915,N_2395,N_256);
nand U3916 (N_3916,N_2020,N_1556);
nor U3917 (N_3917,N_761,N_899);
nand U3918 (N_3918,N_2418,N_1006);
nor U3919 (N_3919,N_1345,N_1574);
xnor U3920 (N_3920,N_2285,N_1811);
nor U3921 (N_3921,N_687,N_1797);
nor U3922 (N_3922,N_551,N_1869);
or U3923 (N_3923,N_2376,N_2029);
xnor U3924 (N_3924,N_1012,N_534);
nor U3925 (N_3925,N_440,N_2361);
nand U3926 (N_3926,N_2176,N_830);
nand U3927 (N_3927,N_202,N_1416);
nor U3928 (N_3928,N_2326,N_1958);
nand U3929 (N_3929,N_862,N_1961);
nand U3930 (N_3930,N_84,N_257);
or U3931 (N_3931,N_1701,N_1898);
or U3932 (N_3932,N_114,N_1596);
and U3933 (N_3933,N_622,N_1091);
or U3934 (N_3934,N_847,N_939);
nand U3935 (N_3935,N_105,N_830);
and U3936 (N_3936,N_1823,N_2389);
nor U3937 (N_3937,N_1610,N_816);
and U3938 (N_3938,N_837,N_1280);
or U3939 (N_3939,N_2068,N_2137);
xnor U3940 (N_3940,N_731,N_19);
nand U3941 (N_3941,N_1158,N_2169);
and U3942 (N_3942,N_2041,N_879);
and U3943 (N_3943,N_1808,N_2282);
nand U3944 (N_3944,N_1790,N_2391);
nand U3945 (N_3945,N_130,N_706);
nor U3946 (N_3946,N_8,N_1487);
and U3947 (N_3947,N_2366,N_1962);
and U3948 (N_3948,N_1192,N_1805);
or U3949 (N_3949,N_2426,N_1742);
xnor U3950 (N_3950,N_926,N_997);
nor U3951 (N_3951,N_138,N_573);
nor U3952 (N_3952,N_1655,N_1427);
nor U3953 (N_3953,N_2428,N_2021);
nor U3954 (N_3954,N_1742,N_916);
or U3955 (N_3955,N_638,N_2223);
nand U3956 (N_3956,N_2429,N_2074);
nand U3957 (N_3957,N_252,N_1422);
or U3958 (N_3958,N_1047,N_2104);
or U3959 (N_3959,N_1795,N_555);
nor U3960 (N_3960,N_1700,N_1854);
nand U3961 (N_3961,N_167,N_2334);
nand U3962 (N_3962,N_2292,N_438);
nor U3963 (N_3963,N_239,N_1067);
nand U3964 (N_3964,N_2108,N_1397);
nand U3965 (N_3965,N_2179,N_1093);
or U3966 (N_3966,N_2023,N_909);
xnor U3967 (N_3967,N_1313,N_2075);
nor U3968 (N_3968,N_2258,N_495);
or U3969 (N_3969,N_2302,N_1139);
nand U3970 (N_3970,N_1037,N_2458);
and U3971 (N_3971,N_1405,N_20);
nand U3972 (N_3972,N_309,N_1509);
nand U3973 (N_3973,N_1502,N_1210);
or U3974 (N_3974,N_112,N_1051);
nand U3975 (N_3975,N_2320,N_1320);
xnor U3976 (N_3976,N_666,N_1296);
nor U3977 (N_3977,N_661,N_1072);
nor U3978 (N_3978,N_584,N_490);
xnor U3979 (N_3979,N_1142,N_2152);
or U3980 (N_3980,N_1208,N_1716);
or U3981 (N_3981,N_552,N_1654);
nand U3982 (N_3982,N_754,N_1939);
xnor U3983 (N_3983,N_2469,N_1569);
or U3984 (N_3984,N_2188,N_1869);
nand U3985 (N_3985,N_1013,N_431);
xnor U3986 (N_3986,N_2172,N_2039);
nor U3987 (N_3987,N_926,N_1193);
or U3988 (N_3988,N_2355,N_602);
nand U3989 (N_3989,N_2032,N_1968);
or U3990 (N_3990,N_1853,N_2414);
or U3991 (N_3991,N_1151,N_1761);
or U3992 (N_3992,N_1332,N_546);
or U3993 (N_3993,N_1850,N_1972);
nand U3994 (N_3994,N_364,N_1076);
nor U3995 (N_3995,N_2485,N_1801);
nand U3996 (N_3996,N_2217,N_155);
nand U3997 (N_3997,N_586,N_49);
or U3998 (N_3998,N_2159,N_1834);
and U3999 (N_3999,N_706,N_717);
nor U4000 (N_4000,N_794,N_1060);
nand U4001 (N_4001,N_2068,N_18);
or U4002 (N_4002,N_2105,N_386);
or U4003 (N_4003,N_682,N_320);
and U4004 (N_4004,N_966,N_47);
and U4005 (N_4005,N_315,N_268);
nor U4006 (N_4006,N_436,N_1377);
nor U4007 (N_4007,N_2093,N_80);
nand U4008 (N_4008,N_5,N_999);
nor U4009 (N_4009,N_1145,N_87);
or U4010 (N_4010,N_1719,N_1372);
nor U4011 (N_4011,N_1567,N_839);
nand U4012 (N_4012,N_1748,N_1781);
xor U4013 (N_4013,N_1312,N_6);
and U4014 (N_4014,N_1507,N_1415);
and U4015 (N_4015,N_1724,N_1546);
nand U4016 (N_4016,N_1788,N_1405);
and U4017 (N_4017,N_1424,N_1214);
nor U4018 (N_4018,N_2099,N_1635);
xor U4019 (N_4019,N_91,N_1274);
nor U4020 (N_4020,N_1753,N_1611);
nor U4021 (N_4021,N_2132,N_528);
nand U4022 (N_4022,N_845,N_1576);
nand U4023 (N_4023,N_2258,N_203);
or U4024 (N_4024,N_1555,N_2087);
nor U4025 (N_4025,N_2025,N_1095);
nor U4026 (N_4026,N_884,N_1044);
or U4027 (N_4027,N_1750,N_2111);
xnor U4028 (N_4028,N_757,N_1556);
nand U4029 (N_4029,N_1020,N_1109);
and U4030 (N_4030,N_826,N_1767);
nor U4031 (N_4031,N_778,N_1127);
and U4032 (N_4032,N_1727,N_608);
nand U4033 (N_4033,N_970,N_2307);
nand U4034 (N_4034,N_2396,N_1843);
and U4035 (N_4035,N_2293,N_1273);
nor U4036 (N_4036,N_628,N_1099);
xnor U4037 (N_4037,N_1433,N_283);
nor U4038 (N_4038,N_494,N_2445);
or U4039 (N_4039,N_2113,N_807);
nand U4040 (N_4040,N_2075,N_2047);
or U4041 (N_4041,N_1570,N_289);
or U4042 (N_4042,N_1670,N_342);
and U4043 (N_4043,N_1886,N_1669);
or U4044 (N_4044,N_1714,N_1973);
or U4045 (N_4045,N_254,N_338);
or U4046 (N_4046,N_1897,N_1664);
nor U4047 (N_4047,N_205,N_2087);
nand U4048 (N_4048,N_176,N_881);
nand U4049 (N_4049,N_2278,N_58);
nand U4050 (N_4050,N_1804,N_2280);
nand U4051 (N_4051,N_694,N_400);
nand U4052 (N_4052,N_2495,N_662);
nand U4053 (N_4053,N_1769,N_867);
nor U4054 (N_4054,N_789,N_2317);
nand U4055 (N_4055,N_1822,N_2457);
nor U4056 (N_4056,N_2242,N_1687);
and U4057 (N_4057,N_372,N_2361);
xor U4058 (N_4058,N_1749,N_1797);
and U4059 (N_4059,N_1692,N_40);
and U4060 (N_4060,N_2462,N_2474);
nor U4061 (N_4061,N_1551,N_2315);
nor U4062 (N_4062,N_101,N_878);
nor U4063 (N_4063,N_2210,N_1940);
and U4064 (N_4064,N_991,N_1194);
or U4065 (N_4065,N_1846,N_1743);
and U4066 (N_4066,N_235,N_2364);
or U4067 (N_4067,N_2465,N_2132);
and U4068 (N_4068,N_2043,N_221);
and U4069 (N_4069,N_634,N_2061);
nand U4070 (N_4070,N_1430,N_1188);
nor U4071 (N_4071,N_1539,N_2456);
nor U4072 (N_4072,N_1443,N_696);
and U4073 (N_4073,N_1054,N_2308);
nor U4074 (N_4074,N_2238,N_1617);
nand U4075 (N_4075,N_1997,N_50);
nand U4076 (N_4076,N_2497,N_1628);
nor U4077 (N_4077,N_1162,N_378);
xor U4078 (N_4078,N_2007,N_316);
and U4079 (N_4079,N_2366,N_1562);
and U4080 (N_4080,N_1284,N_1389);
or U4081 (N_4081,N_50,N_352);
xnor U4082 (N_4082,N_216,N_2389);
nor U4083 (N_4083,N_2261,N_562);
nor U4084 (N_4084,N_2185,N_999);
and U4085 (N_4085,N_51,N_1007);
xnor U4086 (N_4086,N_1088,N_973);
nor U4087 (N_4087,N_935,N_2228);
and U4088 (N_4088,N_465,N_716);
and U4089 (N_4089,N_1475,N_693);
nor U4090 (N_4090,N_1716,N_896);
nand U4091 (N_4091,N_1572,N_1583);
and U4092 (N_4092,N_836,N_651);
nor U4093 (N_4093,N_1564,N_1489);
nand U4094 (N_4094,N_406,N_282);
and U4095 (N_4095,N_2436,N_2018);
nor U4096 (N_4096,N_1123,N_457);
nand U4097 (N_4097,N_265,N_1153);
nor U4098 (N_4098,N_313,N_1935);
nand U4099 (N_4099,N_1817,N_2165);
nor U4100 (N_4100,N_893,N_2122);
and U4101 (N_4101,N_533,N_1833);
xnor U4102 (N_4102,N_1727,N_657);
nor U4103 (N_4103,N_1481,N_423);
and U4104 (N_4104,N_1561,N_1693);
nand U4105 (N_4105,N_2373,N_2370);
or U4106 (N_4106,N_2101,N_1943);
nor U4107 (N_4107,N_2318,N_1189);
or U4108 (N_4108,N_2054,N_45);
nor U4109 (N_4109,N_1320,N_1422);
or U4110 (N_4110,N_627,N_92);
or U4111 (N_4111,N_2268,N_277);
nor U4112 (N_4112,N_1153,N_355);
and U4113 (N_4113,N_1013,N_1573);
nand U4114 (N_4114,N_343,N_340);
or U4115 (N_4115,N_1610,N_1345);
or U4116 (N_4116,N_989,N_957);
and U4117 (N_4117,N_514,N_2033);
nor U4118 (N_4118,N_2241,N_2408);
nand U4119 (N_4119,N_1295,N_644);
or U4120 (N_4120,N_1819,N_1795);
nor U4121 (N_4121,N_712,N_551);
and U4122 (N_4122,N_1890,N_726);
nand U4123 (N_4123,N_1696,N_32);
and U4124 (N_4124,N_627,N_1304);
or U4125 (N_4125,N_596,N_1696);
nand U4126 (N_4126,N_885,N_54);
nor U4127 (N_4127,N_2348,N_512);
nor U4128 (N_4128,N_2222,N_643);
nand U4129 (N_4129,N_956,N_1869);
nor U4130 (N_4130,N_550,N_753);
xnor U4131 (N_4131,N_2113,N_2122);
and U4132 (N_4132,N_755,N_749);
xor U4133 (N_4133,N_2155,N_861);
or U4134 (N_4134,N_1206,N_1982);
xor U4135 (N_4135,N_1721,N_1557);
xor U4136 (N_4136,N_621,N_1872);
nor U4137 (N_4137,N_1624,N_40);
nor U4138 (N_4138,N_1045,N_1265);
nor U4139 (N_4139,N_1627,N_1512);
and U4140 (N_4140,N_1896,N_1299);
or U4141 (N_4141,N_823,N_841);
and U4142 (N_4142,N_1195,N_1781);
or U4143 (N_4143,N_24,N_107);
nand U4144 (N_4144,N_1989,N_1068);
nor U4145 (N_4145,N_1063,N_300);
nand U4146 (N_4146,N_1612,N_2174);
or U4147 (N_4147,N_592,N_1945);
and U4148 (N_4148,N_581,N_2377);
nor U4149 (N_4149,N_53,N_243);
or U4150 (N_4150,N_1550,N_2343);
or U4151 (N_4151,N_1163,N_1809);
nand U4152 (N_4152,N_2229,N_508);
and U4153 (N_4153,N_482,N_849);
and U4154 (N_4154,N_2120,N_2000);
nor U4155 (N_4155,N_780,N_87);
and U4156 (N_4156,N_1883,N_124);
or U4157 (N_4157,N_680,N_770);
nand U4158 (N_4158,N_450,N_645);
and U4159 (N_4159,N_1673,N_1806);
and U4160 (N_4160,N_854,N_527);
and U4161 (N_4161,N_1777,N_1859);
nor U4162 (N_4162,N_363,N_824);
nand U4163 (N_4163,N_1161,N_671);
or U4164 (N_4164,N_638,N_475);
and U4165 (N_4165,N_124,N_939);
or U4166 (N_4166,N_1834,N_2301);
or U4167 (N_4167,N_1108,N_2195);
xor U4168 (N_4168,N_662,N_2343);
and U4169 (N_4169,N_1575,N_2059);
nand U4170 (N_4170,N_1558,N_2159);
nor U4171 (N_4171,N_2272,N_2262);
nor U4172 (N_4172,N_1400,N_1958);
or U4173 (N_4173,N_69,N_165);
nor U4174 (N_4174,N_1269,N_882);
nor U4175 (N_4175,N_2159,N_2350);
nor U4176 (N_4176,N_727,N_2094);
nand U4177 (N_4177,N_2121,N_2328);
nand U4178 (N_4178,N_1778,N_351);
and U4179 (N_4179,N_269,N_98);
nand U4180 (N_4180,N_1210,N_606);
nor U4181 (N_4181,N_204,N_937);
and U4182 (N_4182,N_141,N_1667);
or U4183 (N_4183,N_395,N_372);
and U4184 (N_4184,N_1912,N_675);
or U4185 (N_4185,N_815,N_1866);
nand U4186 (N_4186,N_1831,N_2167);
and U4187 (N_4187,N_2437,N_484);
or U4188 (N_4188,N_222,N_1326);
and U4189 (N_4189,N_763,N_1055);
xor U4190 (N_4190,N_108,N_1011);
xor U4191 (N_4191,N_2011,N_1715);
nand U4192 (N_4192,N_570,N_306);
xor U4193 (N_4193,N_1984,N_2464);
or U4194 (N_4194,N_643,N_820);
nor U4195 (N_4195,N_397,N_1134);
nor U4196 (N_4196,N_2484,N_918);
xor U4197 (N_4197,N_839,N_630);
nand U4198 (N_4198,N_694,N_896);
nand U4199 (N_4199,N_522,N_440);
xnor U4200 (N_4200,N_1575,N_502);
xor U4201 (N_4201,N_1271,N_317);
or U4202 (N_4202,N_1309,N_872);
xnor U4203 (N_4203,N_1874,N_1130);
and U4204 (N_4204,N_967,N_1674);
xor U4205 (N_4205,N_618,N_544);
xnor U4206 (N_4206,N_1014,N_546);
and U4207 (N_4207,N_2,N_1955);
and U4208 (N_4208,N_1796,N_2048);
or U4209 (N_4209,N_1754,N_1880);
or U4210 (N_4210,N_1509,N_1493);
and U4211 (N_4211,N_928,N_1140);
xor U4212 (N_4212,N_669,N_64);
xnor U4213 (N_4213,N_2380,N_152);
nand U4214 (N_4214,N_1704,N_1201);
and U4215 (N_4215,N_2122,N_1650);
nor U4216 (N_4216,N_2026,N_660);
and U4217 (N_4217,N_1112,N_1401);
nor U4218 (N_4218,N_553,N_1096);
or U4219 (N_4219,N_1166,N_2377);
or U4220 (N_4220,N_306,N_1146);
nand U4221 (N_4221,N_81,N_1108);
nand U4222 (N_4222,N_796,N_2136);
or U4223 (N_4223,N_1231,N_1217);
nor U4224 (N_4224,N_1352,N_1121);
nand U4225 (N_4225,N_856,N_185);
nand U4226 (N_4226,N_1402,N_138);
and U4227 (N_4227,N_85,N_496);
nand U4228 (N_4228,N_764,N_669);
xnor U4229 (N_4229,N_453,N_142);
nor U4230 (N_4230,N_965,N_1227);
and U4231 (N_4231,N_611,N_144);
nand U4232 (N_4232,N_1499,N_2147);
xnor U4233 (N_4233,N_57,N_284);
and U4234 (N_4234,N_2379,N_1785);
or U4235 (N_4235,N_119,N_28);
and U4236 (N_4236,N_952,N_963);
or U4237 (N_4237,N_290,N_2060);
and U4238 (N_4238,N_1797,N_807);
and U4239 (N_4239,N_1172,N_2382);
nand U4240 (N_4240,N_720,N_865);
nand U4241 (N_4241,N_857,N_309);
and U4242 (N_4242,N_847,N_178);
or U4243 (N_4243,N_1170,N_325);
nand U4244 (N_4244,N_1985,N_331);
and U4245 (N_4245,N_2061,N_2469);
or U4246 (N_4246,N_1846,N_1210);
and U4247 (N_4247,N_48,N_2104);
and U4248 (N_4248,N_1441,N_40);
nand U4249 (N_4249,N_2022,N_2037);
and U4250 (N_4250,N_191,N_1684);
nand U4251 (N_4251,N_477,N_255);
and U4252 (N_4252,N_1656,N_627);
xnor U4253 (N_4253,N_1715,N_2350);
xor U4254 (N_4254,N_2174,N_1667);
and U4255 (N_4255,N_508,N_2158);
or U4256 (N_4256,N_1400,N_880);
nand U4257 (N_4257,N_1351,N_1165);
nor U4258 (N_4258,N_656,N_608);
nand U4259 (N_4259,N_1531,N_2286);
nor U4260 (N_4260,N_1210,N_475);
nand U4261 (N_4261,N_1403,N_440);
nand U4262 (N_4262,N_818,N_769);
and U4263 (N_4263,N_1884,N_1372);
nand U4264 (N_4264,N_2343,N_543);
and U4265 (N_4265,N_1749,N_2448);
and U4266 (N_4266,N_139,N_1091);
xnor U4267 (N_4267,N_1547,N_691);
nand U4268 (N_4268,N_1432,N_1431);
xor U4269 (N_4269,N_1028,N_2351);
nor U4270 (N_4270,N_863,N_843);
and U4271 (N_4271,N_1072,N_1464);
or U4272 (N_4272,N_284,N_2362);
and U4273 (N_4273,N_1746,N_1242);
and U4274 (N_4274,N_1727,N_260);
nor U4275 (N_4275,N_403,N_346);
nand U4276 (N_4276,N_1089,N_1997);
xor U4277 (N_4277,N_1005,N_737);
or U4278 (N_4278,N_2408,N_499);
nand U4279 (N_4279,N_911,N_2380);
nand U4280 (N_4280,N_1503,N_931);
and U4281 (N_4281,N_1808,N_105);
nand U4282 (N_4282,N_2250,N_2311);
nor U4283 (N_4283,N_1491,N_1053);
xor U4284 (N_4284,N_1202,N_1677);
nand U4285 (N_4285,N_124,N_860);
nand U4286 (N_4286,N_190,N_578);
nand U4287 (N_4287,N_1583,N_45);
and U4288 (N_4288,N_724,N_1465);
or U4289 (N_4289,N_1159,N_402);
nor U4290 (N_4290,N_1705,N_1166);
xor U4291 (N_4291,N_325,N_650);
and U4292 (N_4292,N_2058,N_1595);
or U4293 (N_4293,N_152,N_2478);
xor U4294 (N_4294,N_818,N_542);
or U4295 (N_4295,N_1748,N_2372);
or U4296 (N_4296,N_2263,N_2101);
and U4297 (N_4297,N_1704,N_1413);
and U4298 (N_4298,N_1437,N_1505);
nor U4299 (N_4299,N_1201,N_2049);
and U4300 (N_4300,N_1837,N_2124);
nor U4301 (N_4301,N_822,N_2415);
nand U4302 (N_4302,N_2057,N_1698);
and U4303 (N_4303,N_2099,N_2117);
nand U4304 (N_4304,N_2460,N_2262);
and U4305 (N_4305,N_365,N_2289);
nand U4306 (N_4306,N_1832,N_1475);
and U4307 (N_4307,N_1651,N_2127);
or U4308 (N_4308,N_1738,N_1811);
nand U4309 (N_4309,N_1763,N_1927);
nor U4310 (N_4310,N_1879,N_2424);
or U4311 (N_4311,N_483,N_2038);
or U4312 (N_4312,N_552,N_1746);
nor U4313 (N_4313,N_820,N_710);
and U4314 (N_4314,N_1099,N_166);
or U4315 (N_4315,N_1893,N_2277);
and U4316 (N_4316,N_1983,N_1675);
or U4317 (N_4317,N_286,N_2178);
or U4318 (N_4318,N_296,N_813);
nand U4319 (N_4319,N_1247,N_1105);
xnor U4320 (N_4320,N_1207,N_718);
nand U4321 (N_4321,N_230,N_66);
and U4322 (N_4322,N_1955,N_526);
and U4323 (N_4323,N_363,N_1415);
nor U4324 (N_4324,N_1266,N_1060);
and U4325 (N_4325,N_510,N_2127);
and U4326 (N_4326,N_996,N_30);
xnor U4327 (N_4327,N_411,N_499);
nand U4328 (N_4328,N_890,N_2234);
or U4329 (N_4329,N_242,N_2241);
nor U4330 (N_4330,N_1767,N_2125);
or U4331 (N_4331,N_2470,N_596);
or U4332 (N_4332,N_1229,N_1154);
and U4333 (N_4333,N_962,N_254);
nand U4334 (N_4334,N_1954,N_584);
nor U4335 (N_4335,N_270,N_782);
or U4336 (N_4336,N_2126,N_2020);
and U4337 (N_4337,N_1407,N_838);
nor U4338 (N_4338,N_2227,N_1993);
or U4339 (N_4339,N_359,N_863);
nand U4340 (N_4340,N_1132,N_1945);
or U4341 (N_4341,N_2056,N_775);
xnor U4342 (N_4342,N_953,N_50);
and U4343 (N_4343,N_495,N_1492);
nor U4344 (N_4344,N_2150,N_237);
or U4345 (N_4345,N_1962,N_1360);
and U4346 (N_4346,N_2497,N_1105);
nor U4347 (N_4347,N_999,N_3);
nor U4348 (N_4348,N_268,N_680);
and U4349 (N_4349,N_53,N_2262);
nand U4350 (N_4350,N_652,N_809);
and U4351 (N_4351,N_299,N_9);
nor U4352 (N_4352,N_700,N_2230);
and U4353 (N_4353,N_371,N_624);
and U4354 (N_4354,N_1960,N_1825);
nor U4355 (N_4355,N_1551,N_951);
and U4356 (N_4356,N_1431,N_2116);
or U4357 (N_4357,N_1472,N_400);
nand U4358 (N_4358,N_869,N_381);
nor U4359 (N_4359,N_1104,N_965);
or U4360 (N_4360,N_132,N_168);
nand U4361 (N_4361,N_2435,N_1649);
and U4362 (N_4362,N_2254,N_1067);
or U4363 (N_4363,N_620,N_1777);
nor U4364 (N_4364,N_489,N_1737);
nand U4365 (N_4365,N_805,N_1353);
nand U4366 (N_4366,N_257,N_1431);
and U4367 (N_4367,N_1125,N_773);
nand U4368 (N_4368,N_1783,N_105);
or U4369 (N_4369,N_943,N_1872);
nand U4370 (N_4370,N_741,N_1273);
or U4371 (N_4371,N_614,N_1884);
nand U4372 (N_4372,N_627,N_415);
or U4373 (N_4373,N_1298,N_2134);
nor U4374 (N_4374,N_2441,N_764);
nand U4375 (N_4375,N_622,N_822);
nand U4376 (N_4376,N_739,N_1237);
xnor U4377 (N_4377,N_114,N_211);
nor U4378 (N_4378,N_1940,N_38);
and U4379 (N_4379,N_384,N_2268);
or U4380 (N_4380,N_1863,N_19);
nand U4381 (N_4381,N_996,N_916);
xnor U4382 (N_4382,N_1491,N_2088);
or U4383 (N_4383,N_230,N_294);
and U4384 (N_4384,N_1081,N_2247);
nor U4385 (N_4385,N_2302,N_1626);
nor U4386 (N_4386,N_21,N_75);
nand U4387 (N_4387,N_2091,N_656);
nor U4388 (N_4388,N_357,N_1616);
nor U4389 (N_4389,N_951,N_1839);
nand U4390 (N_4390,N_1307,N_1954);
and U4391 (N_4391,N_2281,N_645);
xnor U4392 (N_4392,N_1176,N_1243);
nor U4393 (N_4393,N_2386,N_157);
nand U4394 (N_4394,N_976,N_226);
or U4395 (N_4395,N_1719,N_1746);
or U4396 (N_4396,N_1059,N_160);
nand U4397 (N_4397,N_1126,N_1976);
and U4398 (N_4398,N_2174,N_1196);
and U4399 (N_4399,N_550,N_1698);
or U4400 (N_4400,N_448,N_1934);
or U4401 (N_4401,N_1378,N_2016);
nand U4402 (N_4402,N_657,N_2206);
nor U4403 (N_4403,N_1605,N_230);
or U4404 (N_4404,N_2304,N_26);
or U4405 (N_4405,N_1235,N_31);
or U4406 (N_4406,N_2335,N_982);
or U4407 (N_4407,N_889,N_181);
nand U4408 (N_4408,N_689,N_1880);
nor U4409 (N_4409,N_1059,N_1322);
and U4410 (N_4410,N_1082,N_263);
nor U4411 (N_4411,N_498,N_194);
and U4412 (N_4412,N_1626,N_1375);
or U4413 (N_4413,N_1642,N_413);
or U4414 (N_4414,N_1296,N_526);
and U4415 (N_4415,N_2313,N_645);
xnor U4416 (N_4416,N_89,N_378);
and U4417 (N_4417,N_414,N_705);
nor U4418 (N_4418,N_967,N_2295);
or U4419 (N_4419,N_1812,N_1463);
nor U4420 (N_4420,N_1878,N_2102);
or U4421 (N_4421,N_1947,N_1455);
and U4422 (N_4422,N_1794,N_329);
nor U4423 (N_4423,N_2331,N_1054);
or U4424 (N_4424,N_910,N_1316);
xor U4425 (N_4425,N_1023,N_332);
and U4426 (N_4426,N_1807,N_2409);
nand U4427 (N_4427,N_622,N_1133);
nand U4428 (N_4428,N_435,N_738);
nand U4429 (N_4429,N_2225,N_2407);
xnor U4430 (N_4430,N_548,N_168);
or U4431 (N_4431,N_2327,N_1540);
nor U4432 (N_4432,N_2170,N_291);
or U4433 (N_4433,N_1552,N_108);
and U4434 (N_4434,N_2196,N_1424);
nor U4435 (N_4435,N_1029,N_2160);
and U4436 (N_4436,N_2218,N_1763);
and U4437 (N_4437,N_1057,N_1157);
or U4438 (N_4438,N_109,N_1513);
nor U4439 (N_4439,N_10,N_853);
or U4440 (N_4440,N_44,N_1814);
nor U4441 (N_4441,N_457,N_808);
nor U4442 (N_4442,N_2253,N_1011);
nand U4443 (N_4443,N_996,N_2045);
nand U4444 (N_4444,N_1024,N_1760);
nor U4445 (N_4445,N_793,N_1967);
nor U4446 (N_4446,N_1150,N_1110);
xor U4447 (N_4447,N_1935,N_1440);
nand U4448 (N_4448,N_1226,N_56);
and U4449 (N_4449,N_1972,N_1459);
and U4450 (N_4450,N_2139,N_26);
and U4451 (N_4451,N_836,N_394);
nand U4452 (N_4452,N_736,N_1129);
nand U4453 (N_4453,N_2181,N_192);
and U4454 (N_4454,N_2114,N_1497);
nand U4455 (N_4455,N_1891,N_987);
and U4456 (N_4456,N_25,N_742);
and U4457 (N_4457,N_869,N_456);
nand U4458 (N_4458,N_1841,N_48);
and U4459 (N_4459,N_771,N_1172);
or U4460 (N_4460,N_1746,N_1125);
or U4461 (N_4461,N_369,N_1417);
or U4462 (N_4462,N_281,N_2329);
xor U4463 (N_4463,N_1703,N_2452);
and U4464 (N_4464,N_985,N_886);
nor U4465 (N_4465,N_2417,N_659);
and U4466 (N_4466,N_1982,N_1292);
or U4467 (N_4467,N_376,N_1475);
and U4468 (N_4468,N_1151,N_2271);
nand U4469 (N_4469,N_258,N_183);
nor U4470 (N_4470,N_871,N_2345);
nand U4471 (N_4471,N_1256,N_1880);
nor U4472 (N_4472,N_2145,N_1785);
nor U4473 (N_4473,N_1666,N_1441);
and U4474 (N_4474,N_1555,N_1621);
nor U4475 (N_4475,N_404,N_2291);
nor U4476 (N_4476,N_2009,N_212);
nand U4477 (N_4477,N_1566,N_711);
nor U4478 (N_4478,N_1222,N_1245);
xor U4479 (N_4479,N_690,N_2339);
nand U4480 (N_4480,N_1859,N_905);
nor U4481 (N_4481,N_738,N_2451);
or U4482 (N_4482,N_1731,N_636);
nor U4483 (N_4483,N_1798,N_391);
or U4484 (N_4484,N_2174,N_1779);
or U4485 (N_4485,N_2251,N_588);
nand U4486 (N_4486,N_1607,N_285);
and U4487 (N_4487,N_1759,N_1549);
or U4488 (N_4488,N_720,N_514);
and U4489 (N_4489,N_1012,N_769);
or U4490 (N_4490,N_1929,N_1943);
nand U4491 (N_4491,N_465,N_1055);
nor U4492 (N_4492,N_1105,N_2107);
or U4493 (N_4493,N_1174,N_1747);
or U4494 (N_4494,N_390,N_298);
and U4495 (N_4495,N_486,N_935);
nor U4496 (N_4496,N_1655,N_1801);
nand U4497 (N_4497,N_834,N_223);
nand U4498 (N_4498,N_1631,N_34);
or U4499 (N_4499,N_1977,N_1661);
xnor U4500 (N_4500,N_1975,N_660);
nor U4501 (N_4501,N_188,N_1120);
and U4502 (N_4502,N_1331,N_2485);
nand U4503 (N_4503,N_500,N_1336);
and U4504 (N_4504,N_63,N_1489);
or U4505 (N_4505,N_162,N_396);
or U4506 (N_4506,N_1948,N_1824);
or U4507 (N_4507,N_1242,N_2119);
and U4508 (N_4508,N_2490,N_995);
nand U4509 (N_4509,N_1799,N_2211);
nor U4510 (N_4510,N_120,N_22);
xor U4511 (N_4511,N_32,N_1498);
and U4512 (N_4512,N_1360,N_247);
nor U4513 (N_4513,N_1749,N_632);
or U4514 (N_4514,N_2274,N_2488);
and U4515 (N_4515,N_290,N_1355);
or U4516 (N_4516,N_879,N_2381);
nand U4517 (N_4517,N_2230,N_452);
nand U4518 (N_4518,N_1321,N_2470);
or U4519 (N_4519,N_925,N_635);
and U4520 (N_4520,N_1282,N_132);
or U4521 (N_4521,N_466,N_360);
or U4522 (N_4522,N_703,N_2492);
nand U4523 (N_4523,N_2241,N_1574);
nand U4524 (N_4524,N_2335,N_1647);
nand U4525 (N_4525,N_1020,N_941);
nor U4526 (N_4526,N_378,N_2269);
and U4527 (N_4527,N_634,N_995);
or U4528 (N_4528,N_2006,N_961);
or U4529 (N_4529,N_1552,N_991);
nand U4530 (N_4530,N_1778,N_286);
nor U4531 (N_4531,N_1761,N_1275);
nand U4532 (N_4532,N_1748,N_1243);
nor U4533 (N_4533,N_2049,N_2416);
or U4534 (N_4534,N_1618,N_1048);
and U4535 (N_4535,N_694,N_1747);
or U4536 (N_4536,N_2048,N_1993);
nor U4537 (N_4537,N_1051,N_615);
xor U4538 (N_4538,N_1532,N_2314);
nand U4539 (N_4539,N_906,N_555);
nor U4540 (N_4540,N_1697,N_482);
nand U4541 (N_4541,N_665,N_661);
or U4542 (N_4542,N_2195,N_700);
nor U4543 (N_4543,N_1075,N_685);
xnor U4544 (N_4544,N_1474,N_2372);
xor U4545 (N_4545,N_2313,N_1963);
and U4546 (N_4546,N_2018,N_871);
and U4547 (N_4547,N_801,N_2327);
nand U4548 (N_4548,N_1016,N_1203);
or U4549 (N_4549,N_1026,N_578);
nand U4550 (N_4550,N_1448,N_2036);
xnor U4551 (N_4551,N_2052,N_1911);
and U4552 (N_4552,N_1240,N_672);
nand U4553 (N_4553,N_276,N_1197);
or U4554 (N_4554,N_784,N_750);
and U4555 (N_4555,N_336,N_1506);
nand U4556 (N_4556,N_731,N_1998);
nand U4557 (N_4557,N_2334,N_2289);
and U4558 (N_4558,N_1075,N_1634);
and U4559 (N_4559,N_1197,N_1230);
nand U4560 (N_4560,N_1551,N_2236);
nor U4561 (N_4561,N_1205,N_1947);
nor U4562 (N_4562,N_1356,N_502);
xnor U4563 (N_4563,N_297,N_1299);
nor U4564 (N_4564,N_2149,N_2475);
xor U4565 (N_4565,N_95,N_1606);
or U4566 (N_4566,N_1357,N_1055);
nand U4567 (N_4567,N_687,N_1463);
nor U4568 (N_4568,N_697,N_1921);
nand U4569 (N_4569,N_1124,N_899);
nor U4570 (N_4570,N_333,N_2294);
or U4571 (N_4571,N_2155,N_902);
or U4572 (N_4572,N_596,N_2327);
nand U4573 (N_4573,N_1479,N_2092);
or U4574 (N_4574,N_2374,N_632);
nand U4575 (N_4575,N_2366,N_1238);
nor U4576 (N_4576,N_483,N_363);
nand U4577 (N_4577,N_437,N_2237);
xor U4578 (N_4578,N_1835,N_1828);
nand U4579 (N_4579,N_1799,N_463);
or U4580 (N_4580,N_933,N_521);
xnor U4581 (N_4581,N_883,N_2043);
and U4582 (N_4582,N_1605,N_1169);
and U4583 (N_4583,N_521,N_578);
nor U4584 (N_4584,N_1031,N_1063);
nor U4585 (N_4585,N_2309,N_1134);
nand U4586 (N_4586,N_650,N_330);
xnor U4587 (N_4587,N_866,N_2308);
or U4588 (N_4588,N_839,N_1870);
nor U4589 (N_4589,N_969,N_826);
or U4590 (N_4590,N_1406,N_185);
nor U4591 (N_4591,N_1319,N_1520);
and U4592 (N_4592,N_120,N_2499);
nor U4593 (N_4593,N_1730,N_858);
and U4594 (N_4594,N_1844,N_1728);
and U4595 (N_4595,N_547,N_1637);
xor U4596 (N_4596,N_1990,N_656);
and U4597 (N_4597,N_671,N_935);
or U4598 (N_4598,N_2209,N_1253);
nand U4599 (N_4599,N_1065,N_2219);
nand U4600 (N_4600,N_147,N_641);
or U4601 (N_4601,N_386,N_157);
nor U4602 (N_4602,N_1905,N_1362);
nor U4603 (N_4603,N_749,N_831);
nor U4604 (N_4604,N_1258,N_334);
nor U4605 (N_4605,N_1403,N_732);
nand U4606 (N_4606,N_1607,N_900);
and U4607 (N_4607,N_380,N_2341);
nand U4608 (N_4608,N_2271,N_1621);
or U4609 (N_4609,N_1006,N_174);
nand U4610 (N_4610,N_551,N_2009);
nand U4611 (N_4611,N_1298,N_2463);
or U4612 (N_4612,N_1371,N_1140);
nand U4613 (N_4613,N_1626,N_1301);
and U4614 (N_4614,N_2169,N_1782);
nand U4615 (N_4615,N_109,N_2188);
or U4616 (N_4616,N_2032,N_1943);
nor U4617 (N_4617,N_216,N_972);
nor U4618 (N_4618,N_674,N_1483);
nor U4619 (N_4619,N_2077,N_624);
nand U4620 (N_4620,N_690,N_1299);
and U4621 (N_4621,N_2425,N_961);
and U4622 (N_4622,N_35,N_2270);
nor U4623 (N_4623,N_435,N_1224);
xor U4624 (N_4624,N_1480,N_777);
or U4625 (N_4625,N_2095,N_1375);
xor U4626 (N_4626,N_834,N_1201);
nor U4627 (N_4627,N_2498,N_571);
nand U4628 (N_4628,N_888,N_375);
xor U4629 (N_4629,N_1539,N_1706);
or U4630 (N_4630,N_1315,N_1098);
or U4631 (N_4631,N_911,N_1586);
nand U4632 (N_4632,N_867,N_1043);
or U4633 (N_4633,N_347,N_406);
nor U4634 (N_4634,N_151,N_1178);
nor U4635 (N_4635,N_833,N_461);
nor U4636 (N_4636,N_1742,N_1888);
nor U4637 (N_4637,N_585,N_1451);
and U4638 (N_4638,N_1789,N_1783);
nand U4639 (N_4639,N_2397,N_1753);
nor U4640 (N_4640,N_1086,N_1468);
or U4641 (N_4641,N_2420,N_1303);
nand U4642 (N_4642,N_922,N_181);
or U4643 (N_4643,N_2456,N_527);
nand U4644 (N_4644,N_488,N_1127);
or U4645 (N_4645,N_674,N_477);
nand U4646 (N_4646,N_1871,N_1952);
nor U4647 (N_4647,N_506,N_480);
or U4648 (N_4648,N_381,N_960);
nor U4649 (N_4649,N_2102,N_718);
nand U4650 (N_4650,N_458,N_986);
or U4651 (N_4651,N_39,N_758);
nor U4652 (N_4652,N_170,N_1679);
or U4653 (N_4653,N_2431,N_167);
nor U4654 (N_4654,N_1557,N_515);
and U4655 (N_4655,N_1262,N_2247);
nor U4656 (N_4656,N_1178,N_2252);
nor U4657 (N_4657,N_675,N_1549);
xnor U4658 (N_4658,N_755,N_469);
or U4659 (N_4659,N_1855,N_628);
xor U4660 (N_4660,N_148,N_1776);
nor U4661 (N_4661,N_187,N_656);
and U4662 (N_4662,N_251,N_1512);
or U4663 (N_4663,N_41,N_2406);
nand U4664 (N_4664,N_1834,N_589);
and U4665 (N_4665,N_2396,N_809);
nor U4666 (N_4666,N_1491,N_1004);
nand U4667 (N_4667,N_1062,N_2049);
and U4668 (N_4668,N_2406,N_1792);
or U4669 (N_4669,N_2282,N_1740);
or U4670 (N_4670,N_1184,N_32);
nand U4671 (N_4671,N_246,N_2210);
xnor U4672 (N_4672,N_1359,N_955);
or U4673 (N_4673,N_99,N_692);
or U4674 (N_4674,N_65,N_2390);
nor U4675 (N_4675,N_754,N_2239);
nor U4676 (N_4676,N_596,N_1319);
nand U4677 (N_4677,N_2363,N_744);
xor U4678 (N_4678,N_1076,N_793);
nor U4679 (N_4679,N_1938,N_1597);
and U4680 (N_4680,N_2236,N_1377);
nor U4681 (N_4681,N_603,N_2490);
xnor U4682 (N_4682,N_2444,N_1273);
nor U4683 (N_4683,N_465,N_1862);
nor U4684 (N_4684,N_852,N_491);
nand U4685 (N_4685,N_2062,N_1459);
and U4686 (N_4686,N_328,N_663);
nand U4687 (N_4687,N_492,N_701);
xor U4688 (N_4688,N_1133,N_1916);
nor U4689 (N_4689,N_252,N_397);
and U4690 (N_4690,N_1709,N_762);
and U4691 (N_4691,N_1547,N_1676);
nand U4692 (N_4692,N_1151,N_1414);
nor U4693 (N_4693,N_1216,N_1726);
and U4694 (N_4694,N_1075,N_848);
and U4695 (N_4695,N_808,N_988);
and U4696 (N_4696,N_1252,N_1555);
or U4697 (N_4697,N_2071,N_257);
nand U4698 (N_4698,N_1832,N_1146);
or U4699 (N_4699,N_1367,N_1502);
nor U4700 (N_4700,N_345,N_836);
or U4701 (N_4701,N_1015,N_1438);
or U4702 (N_4702,N_1214,N_2456);
nand U4703 (N_4703,N_1734,N_1561);
or U4704 (N_4704,N_1517,N_1804);
and U4705 (N_4705,N_1379,N_2267);
nand U4706 (N_4706,N_1663,N_377);
or U4707 (N_4707,N_2361,N_651);
and U4708 (N_4708,N_2330,N_506);
and U4709 (N_4709,N_648,N_618);
nor U4710 (N_4710,N_792,N_462);
and U4711 (N_4711,N_621,N_2487);
nand U4712 (N_4712,N_1328,N_1432);
nand U4713 (N_4713,N_2029,N_1258);
nand U4714 (N_4714,N_1736,N_926);
xnor U4715 (N_4715,N_1969,N_1989);
and U4716 (N_4716,N_1400,N_1858);
and U4717 (N_4717,N_2462,N_233);
nor U4718 (N_4718,N_859,N_258);
nand U4719 (N_4719,N_1335,N_1772);
and U4720 (N_4720,N_510,N_1133);
or U4721 (N_4721,N_1439,N_1746);
nor U4722 (N_4722,N_1579,N_187);
or U4723 (N_4723,N_2421,N_1569);
and U4724 (N_4724,N_536,N_944);
nand U4725 (N_4725,N_2403,N_453);
or U4726 (N_4726,N_22,N_1149);
nor U4727 (N_4727,N_1677,N_1670);
nor U4728 (N_4728,N_1721,N_4);
or U4729 (N_4729,N_878,N_2227);
or U4730 (N_4730,N_2083,N_1136);
nand U4731 (N_4731,N_1595,N_2338);
and U4732 (N_4732,N_1536,N_271);
nand U4733 (N_4733,N_1404,N_1726);
nor U4734 (N_4734,N_817,N_1474);
nor U4735 (N_4735,N_392,N_2310);
nor U4736 (N_4736,N_1645,N_1109);
nor U4737 (N_4737,N_103,N_552);
and U4738 (N_4738,N_1174,N_1856);
and U4739 (N_4739,N_1486,N_2442);
or U4740 (N_4740,N_2494,N_673);
nor U4741 (N_4741,N_1172,N_465);
and U4742 (N_4742,N_565,N_36);
nor U4743 (N_4743,N_154,N_956);
nand U4744 (N_4744,N_384,N_1929);
xnor U4745 (N_4745,N_1067,N_19);
and U4746 (N_4746,N_1879,N_222);
nor U4747 (N_4747,N_303,N_989);
and U4748 (N_4748,N_650,N_1133);
or U4749 (N_4749,N_785,N_1272);
nand U4750 (N_4750,N_1856,N_2150);
nand U4751 (N_4751,N_2293,N_396);
and U4752 (N_4752,N_1926,N_815);
nor U4753 (N_4753,N_1671,N_1231);
nor U4754 (N_4754,N_71,N_1525);
nand U4755 (N_4755,N_2184,N_1801);
nor U4756 (N_4756,N_1956,N_945);
and U4757 (N_4757,N_2178,N_2121);
and U4758 (N_4758,N_2448,N_2481);
and U4759 (N_4759,N_499,N_1135);
and U4760 (N_4760,N_2477,N_2307);
nor U4761 (N_4761,N_163,N_812);
nor U4762 (N_4762,N_1291,N_1420);
or U4763 (N_4763,N_1114,N_1737);
and U4764 (N_4764,N_613,N_1834);
nor U4765 (N_4765,N_280,N_97);
or U4766 (N_4766,N_2219,N_848);
or U4767 (N_4767,N_1747,N_2126);
nand U4768 (N_4768,N_1621,N_1821);
and U4769 (N_4769,N_424,N_846);
nand U4770 (N_4770,N_2138,N_1777);
and U4771 (N_4771,N_261,N_1170);
and U4772 (N_4772,N_1332,N_224);
or U4773 (N_4773,N_2264,N_34);
and U4774 (N_4774,N_2075,N_1230);
nor U4775 (N_4775,N_1745,N_142);
and U4776 (N_4776,N_2117,N_1310);
nor U4777 (N_4777,N_1255,N_254);
nor U4778 (N_4778,N_1534,N_1299);
nor U4779 (N_4779,N_516,N_1985);
xnor U4780 (N_4780,N_2445,N_1473);
xnor U4781 (N_4781,N_2295,N_2365);
or U4782 (N_4782,N_2475,N_2051);
xor U4783 (N_4783,N_1241,N_520);
nand U4784 (N_4784,N_2127,N_2352);
nor U4785 (N_4785,N_1043,N_364);
and U4786 (N_4786,N_491,N_2067);
nor U4787 (N_4787,N_1833,N_1124);
or U4788 (N_4788,N_120,N_2004);
nor U4789 (N_4789,N_2176,N_1924);
or U4790 (N_4790,N_1290,N_1942);
nor U4791 (N_4791,N_1477,N_568);
and U4792 (N_4792,N_2111,N_134);
or U4793 (N_4793,N_2340,N_614);
or U4794 (N_4794,N_2137,N_691);
and U4795 (N_4795,N_390,N_600);
or U4796 (N_4796,N_2222,N_1683);
xor U4797 (N_4797,N_1239,N_1776);
and U4798 (N_4798,N_984,N_31);
nand U4799 (N_4799,N_517,N_1803);
or U4800 (N_4800,N_576,N_1798);
nor U4801 (N_4801,N_2146,N_1332);
and U4802 (N_4802,N_414,N_76);
and U4803 (N_4803,N_1757,N_1759);
and U4804 (N_4804,N_1668,N_1164);
and U4805 (N_4805,N_2373,N_1769);
or U4806 (N_4806,N_813,N_1533);
or U4807 (N_4807,N_1878,N_2372);
nand U4808 (N_4808,N_747,N_1839);
nor U4809 (N_4809,N_210,N_589);
xor U4810 (N_4810,N_2481,N_570);
and U4811 (N_4811,N_976,N_566);
nand U4812 (N_4812,N_505,N_1912);
nand U4813 (N_4813,N_325,N_2128);
and U4814 (N_4814,N_1882,N_937);
nand U4815 (N_4815,N_1218,N_2144);
and U4816 (N_4816,N_1348,N_2345);
or U4817 (N_4817,N_2349,N_940);
and U4818 (N_4818,N_1119,N_618);
and U4819 (N_4819,N_172,N_1656);
or U4820 (N_4820,N_1283,N_1649);
and U4821 (N_4821,N_1580,N_1356);
nor U4822 (N_4822,N_1991,N_856);
and U4823 (N_4823,N_2257,N_1327);
and U4824 (N_4824,N_981,N_1655);
or U4825 (N_4825,N_976,N_1338);
and U4826 (N_4826,N_1756,N_501);
nor U4827 (N_4827,N_943,N_729);
and U4828 (N_4828,N_2345,N_536);
xnor U4829 (N_4829,N_808,N_1656);
or U4830 (N_4830,N_2391,N_2445);
nor U4831 (N_4831,N_672,N_74);
nand U4832 (N_4832,N_462,N_2166);
nand U4833 (N_4833,N_2369,N_1709);
nor U4834 (N_4834,N_506,N_1068);
nor U4835 (N_4835,N_1292,N_1282);
nor U4836 (N_4836,N_873,N_1974);
nor U4837 (N_4837,N_2170,N_287);
and U4838 (N_4838,N_1261,N_829);
and U4839 (N_4839,N_1179,N_1966);
or U4840 (N_4840,N_1164,N_538);
nor U4841 (N_4841,N_1549,N_2391);
or U4842 (N_4842,N_405,N_1800);
nor U4843 (N_4843,N_1527,N_1762);
nor U4844 (N_4844,N_1534,N_1017);
and U4845 (N_4845,N_157,N_980);
nor U4846 (N_4846,N_412,N_208);
nor U4847 (N_4847,N_1436,N_37);
xor U4848 (N_4848,N_1384,N_221);
nand U4849 (N_4849,N_1109,N_2281);
or U4850 (N_4850,N_1400,N_393);
nor U4851 (N_4851,N_1831,N_2130);
and U4852 (N_4852,N_1711,N_2345);
nor U4853 (N_4853,N_1553,N_2332);
nand U4854 (N_4854,N_1201,N_2206);
xnor U4855 (N_4855,N_846,N_1050);
and U4856 (N_4856,N_694,N_548);
and U4857 (N_4857,N_1149,N_1477);
nand U4858 (N_4858,N_1621,N_1481);
nand U4859 (N_4859,N_2458,N_1331);
or U4860 (N_4860,N_2435,N_1569);
xnor U4861 (N_4861,N_1707,N_114);
and U4862 (N_4862,N_2389,N_2497);
and U4863 (N_4863,N_1520,N_2199);
nor U4864 (N_4864,N_422,N_539);
nand U4865 (N_4865,N_1053,N_777);
and U4866 (N_4866,N_1099,N_2183);
nand U4867 (N_4867,N_436,N_1461);
xor U4868 (N_4868,N_633,N_1591);
nand U4869 (N_4869,N_1303,N_1769);
xor U4870 (N_4870,N_2067,N_857);
xnor U4871 (N_4871,N_1657,N_524);
or U4872 (N_4872,N_1209,N_671);
and U4873 (N_4873,N_1940,N_210);
xnor U4874 (N_4874,N_309,N_20);
or U4875 (N_4875,N_980,N_1390);
and U4876 (N_4876,N_589,N_411);
or U4877 (N_4877,N_2248,N_1503);
or U4878 (N_4878,N_1739,N_1528);
nor U4879 (N_4879,N_1272,N_2038);
or U4880 (N_4880,N_1905,N_860);
and U4881 (N_4881,N_30,N_331);
xnor U4882 (N_4882,N_2020,N_1140);
xor U4883 (N_4883,N_2481,N_696);
and U4884 (N_4884,N_1968,N_516);
or U4885 (N_4885,N_796,N_1582);
and U4886 (N_4886,N_2439,N_729);
nor U4887 (N_4887,N_83,N_2098);
and U4888 (N_4888,N_1827,N_1825);
and U4889 (N_4889,N_1351,N_821);
and U4890 (N_4890,N_1224,N_1531);
xor U4891 (N_4891,N_2219,N_834);
nor U4892 (N_4892,N_1277,N_616);
and U4893 (N_4893,N_1082,N_1450);
nor U4894 (N_4894,N_858,N_844);
nand U4895 (N_4895,N_1622,N_1637);
nor U4896 (N_4896,N_2240,N_1003);
and U4897 (N_4897,N_709,N_1259);
nand U4898 (N_4898,N_331,N_1858);
xnor U4899 (N_4899,N_1479,N_2210);
xor U4900 (N_4900,N_55,N_2270);
and U4901 (N_4901,N_606,N_2486);
or U4902 (N_4902,N_2275,N_1311);
xor U4903 (N_4903,N_2055,N_2013);
or U4904 (N_4904,N_676,N_2434);
or U4905 (N_4905,N_292,N_1879);
or U4906 (N_4906,N_2442,N_2386);
and U4907 (N_4907,N_907,N_1237);
or U4908 (N_4908,N_1623,N_1447);
nand U4909 (N_4909,N_101,N_1085);
nand U4910 (N_4910,N_569,N_2486);
nor U4911 (N_4911,N_78,N_2290);
and U4912 (N_4912,N_1033,N_2244);
and U4913 (N_4913,N_436,N_2474);
and U4914 (N_4914,N_1730,N_1397);
or U4915 (N_4915,N_1108,N_1377);
nand U4916 (N_4916,N_1215,N_1874);
and U4917 (N_4917,N_2130,N_694);
or U4918 (N_4918,N_848,N_2136);
xor U4919 (N_4919,N_937,N_2087);
xor U4920 (N_4920,N_71,N_518);
nand U4921 (N_4921,N_2035,N_2151);
and U4922 (N_4922,N_1514,N_862);
nand U4923 (N_4923,N_1443,N_862);
nand U4924 (N_4924,N_721,N_1868);
and U4925 (N_4925,N_719,N_2033);
nor U4926 (N_4926,N_1101,N_1471);
nand U4927 (N_4927,N_2294,N_1669);
nor U4928 (N_4928,N_636,N_1570);
xor U4929 (N_4929,N_1162,N_498);
nand U4930 (N_4930,N_1876,N_1554);
or U4931 (N_4931,N_323,N_134);
nor U4932 (N_4932,N_895,N_725);
nor U4933 (N_4933,N_1329,N_300);
nor U4934 (N_4934,N_2424,N_2370);
and U4935 (N_4935,N_2486,N_1158);
nor U4936 (N_4936,N_1163,N_843);
and U4937 (N_4937,N_1432,N_53);
nor U4938 (N_4938,N_715,N_1468);
nor U4939 (N_4939,N_1477,N_820);
and U4940 (N_4940,N_1292,N_932);
and U4941 (N_4941,N_2412,N_274);
and U4942 (N_4942,N_1349,N_161);
and U4943 (N_4943,N_1096,N_94);
or U4944 (N_4944,N_1847,N_1197);
nand U4945 (N_4945,N_2107,N_1874);
xor U4946 (N_4946,N_1465,N_423);
nand U4947 (N_4947,N_2293,N_1871);
nor U4948 (N_4948,N_1204,N_1164);
xor U4949 (N_4949,N_663,N_1513);
nor U4950 (N_4950,N_218,N_1552);
or U4951 (N_4951,N_795,N_2253);
nand U4952 (N_4952,N_1637,N_1630);
xnor U4953 (N_4953,N_929,N_2162);
or U4954 (N_4954,N_292,N_549);
nand U4955 (N_4955,N_1490,N_1010);
or U4956 (N_4956,N_1571,N_834);
and U4957 (N_4957,N_2283,N_2196);
nand U4958 (N_4958,N_2105,N_839);
nor U4959 (N_4959,N_1053,N_527);
and U4960 (N_4960,N_280,N_762);
nand U4961 (N_4961,N_2298,N_775);
or U4962 (N_4962,N_2134,N_1164);
nor U4963 (N_4963,N_886,N_1363);
and U4964 (N_4964,N_59,N_2444);
or U4965 (N_4965,N_161,N_1747);
and U4966 (N_4966,N_2282,N_388);
nand U4967 (N_4967,N_2226,N_2001);
xnor U4968 (N_4968,N_1342,N_1880);
nor U4969 (N_4969,N_1656,N_2239);
and U4970 (N_4970,N_2024,N_337);
and U4971 (N_4971,N_1584,N_1148);
nand U4972 (N_4972,N_935,N_100);
xnor U4973 (N_4973,N_2110,N_1677);
and U4974 (N_4974,N_2433,N_1866);
nand U4975 (N_4975,N_2489,N_1169);
nand U4976 (N_4976,N_1234,N_818);
xnor U4977 (N_4977,N_1154,N_537);
xor U4978 (N_4978,N_2408,N_413);
or U4979 (N_4979,N_1784,N_1857);
or U4980 (N_4980,N_96,N_72);
nand U4981 (N_4981,N_63,N_458);
nor U4982 (N_4982,N_666,N_1502);
nor U4983 (N_4983,N_867,N_2395);
and U4984 (N_4984,N_1641,N_1277);
or U4985 (N_4985,N_287,N_636);
or U4986 (N_4986,N_1515,N_2205);
or U4987 (N_4987,N_1407,N_2127);
or U4988 (N_4988,N_1296,N_531);
nand U4989 (N_4989,N_928,N_454);
and U4990 (N_4990,N_2092,N_2107);
nor U4991 (N_4991,N_218,N_1259);
xnor U4992 (N_4992,N_654,N_468);
nand U4993 (N_4993,N_1007,N_1905);
nor U4994 (N_4994,N_726,N_744);
nand U4995 (N_4995,N_323,N_1971);
nor U4996 (N_4996,N_2231,N_609);
nor U4997 (N_4997,N_1330,N_628);
and U4998 (N_4998,N_1993,N_1724);
nand U4999 (N_4999,N_2316,N_1289);
and U5000 (N_5000,N_3943,N_3314);
and U5001 (N_5001,N_2946,N_4893);
nand U5002 (N_5002,N_3996,N_4704);
nor U5003 (N_5003,N_4149,N_3437);
nand U5004 (N_5004,N_4346,N_2826);
nand U5005 (N_5005,N_4265,N_4304);
nand U5006 (N_5006,N_2845,N_4342);
or U5007 (N_5007,N_2839,N_3654);
nor U5008 (N_5008,N_4120,N_3723);
or U5009 (N_5009,N_4091,N_3827);
nand U5010 (N_5010,N_4288,N_4388);
nor U5011 (N_5011,N_3300,N_3375);
nand U5012 (N_5012,N_2999,N_3525);
and U5013 (N_5013,N_4336,N_4912);
or U5014 (N_5014,N_4038,N_2696);
or U5015 (N_5015,N_4549,N_3497);
nor U5016 (N_5016,N_3038,N_4041);
nand U5017 (N_5017,N_2564,N_3502);
nor U5018 (N_5018,N_3086,N_4080);
or U5019 (N_5019,N_4405,N_2661);
or U5020 (N_5020,N_2735,N_4755);
nand U5021 (N_5021,N_3863,N_2534);
xor U5022 (N_5022,N_4918,N_2979);
and U5023 (N_5023,N_2586,N_3735);
nor U5024 (N_5024,N_3492,N_3719);
xor U5025 (N_5025,N_3999,N_3264);
nand U5026 (N_5026,N_2719,N_3706);
nand U5027 (N_5027,N_4409,N_2940);
nand U5028 (N_5028,N_3130,N_3261);
or U5029 (N_5029,N_2553,N_2784);
or U5030 (N_5030,N_4477,N_2760);
and U5031 (N_5031,N_3642,N_3012);
xnor U5032 (N_5032,N_2765,N_3018);
xnor U5033 (N_5033,N_4017,N_3950);
xor U5034 (N_5034,N_3400,N_3600);
and U5035 (N_5035,N_2578,N_3188);
nand U5036 (N_5036,N_3243,N_3193);
and U5037 (N_5037,N_3043,N_3003);
nand U5038 (N_5038,N_4198,N_3818);
nor U5039 (N_5039,N_3832,N_3329);
nand U5040 (N_5040,N_4894,N_4228);
nand U5041 (N_5041,N_4908,N_4571);
nand U5042 (N_5042,N_4447,N_2959);
nand U5043 (N_5043,N_4535,N_3117);
and U5044 (N_5044,N_4012,N_4644);
nor U5045 (N_5045,N_4903,N_4117);
or U5046 (N_5046,N_2676,N_3305);
nor U5047 (N_5047,N_2909,N_3241);
nand U5048 (N_5048,N_3679,N_3078);
or U5049 (N_5049,N_3285,N_3147);
nand U5050 (N_5050,N_2939,N_3429);
or U5051 (N_5051,N_3280,N_3662);
nand U5052 (N_5052,N_3644,N_3697);
or U5053 (N_5053,N_3606,N_4179);
nand U5054 (N_5054,N_4946,N_3568);
or U5055 (N_5055,N_3196,N_4958);
or U5056 (N_5056,N_4039,N_4642);
nor U5057 (N_5057,N_3795,N_4694);
nor U5058 (N_5058,N_2509,N_4508);
nor U5059 (N_5059,N_4431,N_2832);
or U5060 (N_5060,N_3798,N_3883);
nand U5061 (N_5061,N_3744,N_3543);
nor U5062 (N_5062,N_3237,N_2781);
nor U5063 (N_5063,N_3528,N_4247);
nor U5064 (N_5064,N_3537,N_4978);
or U5065 (N_5065,N_4788,N_3076);
or U5066 (N_5066,N_3232,N_2823);
and U5067 (N_5067,N_3918,N_2730);
nand U5068 (N_5068,N_4709,N_3875);
and U5069 (N_5069,N_4167,N_4718);
or U5070 (N_5070,N_3660,N_3365);
or U5071 (N_5071,N_3794,N_4211);
nor U5072 (N_5072,N_3467,N_3974);
and U5073 (N_5073,N_4583,N_4671);
xor U5074 (N_5074,N_4769,N_4424);
nand U5075 (N_5075,N_4793,N_4900);
nor U5076 (N_5076,N_4492,N_3562);
nand U5077 (N_5077,N_4181,N_4019);
nand U5078 (N_5078,N_4837,N_3409);
and U5079 (N_5079,N_3404,N_4350);
nor U5080 (N_5080,N_4525,N_3396);
nor U5081 (N_5081,N_4130,N_4590);
nand U5082 (N_5082,N_2513,N_4372);
or U5083 (N_5083,N_4112,N_4058);
or U5084 (N_5084,N_3511,N_4851);
or U5085 (N_5085,N_4584,N_4257);
or U5086 (N_5086,N_2713,N_4282);
nand U5087 (N_5087,N_4259,N_4371);
nand U5088 (N_5088,N_3820,N_3657);
nand U5089 (N_5089,N_2917,N_3982);
and U5090 (N_5090,N_3036,N_3951);
nor U5091 (N_5091,N_3872,N_4480);
nand U5092 (N_5092,N_3821,N_2532);
nor U5093 (N_5093,N_3262,N_2809);
nor U5094 (N_5094,N_2922,N_4155);
nand U5095 (N_5095,N_2603,N_2745);
and U5096 (N_5096,N_3547,N_4801);
nand U5097 (N_5097,N_4143,N_2813);
and U5098 (N_5098,N_4542,N_4945);
nand U5099 (N_5099,N_4778,N_3037);
nand U5100 (N_5100,N_3961,N_4347);
or U5101 (N_5101,N_3700,N_2754);
or U5102 (N_5102,N_4471,N_2926);
nand U5103 (N_5103,N_4654,N_4066);
and U5104 (N_5104,N_2841,N_2698);
or U5105 (N_5105,N_3273,N_4623);
nor U5106 (N_5106,N_4427,N_3218);
nand U5107 (N_5107,N_3419,N_2865);
nand U5108 (N_5108,N_3810,N_3876);
or U5109 (N_5109,N_4938,N_3604);
and U5110 (N_5110,N_4736,N_4705);
or U5111 (N_5111,N_4649,N_2842);
nand U5112 (N_5112,N_4963,N_4454);
nand U5113 (N_5113,N_3512,N_3206);
or U5114 (N_5114,N_3407,N_3257);
nor U5115 (N_5115,N_4062,N_4760);
nand U5116 (N_5116,N_4854,N_2650);
and U5117 (N_5117,N_4308,N_3755);
nand U5118 (N_5118,N_3632,N_4981);
nand U5119 (N_5119,N_4049,N_3561);
nand U5120 (N_5120,N_4865,N_2533);
nor U5121 (N_5121,N_2976,N_3215);
or U5122 (N_5122,N_4597,N_3682);
or U5123 (N_5123,N_3139,N_4862);
nand U5124 (N_5124,N_4831,N_3111);
and U5125 (N_5125,N_4532,N_4082);
and U5126 (N_5126,N_4666,N_4917);
and U5127 (N_5127,N_4223,N_2975);
and U5128 (N_5128,N_3125,N_4678);
nor U5129 (N_5129,N_3855,N_2715);
nand U5130 (N_5130,N_4916,N_4042);
or U5131 (N_5131,N_2780,N_4108);
or U5132 (N_5132,N_3980,N_4768);
and U5133 (N_5133,N_3824,N_4383);
and U5134 (N_5134,N_2584,N_3886);
xnor U5135 (N_5135,N_3637,N_3819);
nand U5136 (N_5136,N_4224,N_4020);
xnor U5137 (N_5137,N_2554,N_3291);
nand U5138 (N_5138,N_3486,N_3090);
nor U5139 (N_5139,N_4183,N_4533);
xor U5140 (N_5140,N_2751,N_3267);
and U5141 (N_5141,N_3893,N_4048);
nand U5142 (N_5142,N_4613,N_3307);
nor U5143 (N_5143,N_2687,N_3705);
nor U5144 (N_5144,N_2794,N_3712);
nand U5145 (N_5145,N_4708,N_2512);
nand U5146 (N_5146,N_4685,N_3030);
and U5147 (N_5147,N_4081,N_3325);
xnor U5148 (N_5148,N_4460,N_4185);
nor U5149 (N_5149,N_2954,N_4615);
xor U5150 (N_5150,N_2852,N_4973);
nand U5151 (N_5151,N_3717,N_3734);
nand U5152 (N_5152,N_3754,N_4131);
and U5153 (N_5153,N_2771,N_4286);
and U5154 (N_5154,N_3524,N_4258);
nor U5155 (N_5155,N_2673,N_4182);
nand U5156 (N_5156,N_2675,N_4134);
and U5157 (N_5157,N_2507,N_4780);
nor U5158 (N_5158,N_4724,N_3411);
nand U5159 (N_5159,N_3665,N_3355);
and U5160 (N_5160,N_4920,N_4569);
nor U5161 (N_5161,N_3628,N_4115);
and U5162 (N_5162,N_4359,N_3924);
nand U5163 (N_5163,N_2536,N_3689);
or U5164 (N_5164,N_2669,N_3212);
or U5165 (N_5165,N_4832,N_4266);
nand U5166 (N_5166,N_2654,N_2848);
xnor U5167 (N_5167,N_3476,N_3531);
and U5168 (N_5168,N_3358,N_3320);
nor U5169 (N_5169,N_4728,N_3067);
xor U5170 (N_5170,N_4136,N_4199);
and U5171 (N_5171,N_3641,N_4753);
or U5172 (N_5172,N_4180,N_3327);
nor U5173 (N_5173,N_4972,N_4595);
or U5174 (N_5174,N_2645,N_2986);
and U5175 (N_5175,N_3839,N_3049);
nor U5176 (N_5176,N_3666,N_4161);
or U5177 (N_5177,N_4884,N_3146);
nand U5178 (N_5178,N_2680,N_2819);
nor U5179 (N_5179,N_3311,N_2824);
nand U5180 (N_5180,N_4098,N_3097);
nor U5181 (N_5181,N_4071,N_3994);
nor U5182 (N_5182,N_3173,N_4594);
nor U5183 (N_5183,N_2664,N_4621);
nor U5184 (N_5184,N_2652,N_4518);
and U5185 (N_5185,N_3334,N_3447);
nor U5186 (N_5186,N_2821,N_2911);
or U5187 (N_5187,N_4794,N_2605);
nand U5188 (N_5188,N_3091,N_3805);
and U5189 (N_5189,N_3519,N_3945);
nor U5190 (N_5190,N_4074,N_4469);
or U5191 (N_5191,N_3074,N_2526);
and U5192 (N_5192,N_4745,N_3073);
xnor U5193 (N_5193,N_2994,N_3461);
xnor U5194 (N_5194,N_3731,N_3969);
and U5195 (N_5195,N_4164,N_4821);
nor U5196 (N_5196,N_4393,N_4269);
nand U5197 (N_5197,N_2772,N_4194);
nand U5198 (N_5198,N_4501,N_3862);
and U5199 (N_5199,N_2670,N_4838);
nor U5200 (N_5200,N_4146,N_3573);
nand U5201 (N_5201,N_4540,N_2778);
or U5202 (N_5202,N_4422,N_4969);
nand U5203 (N_5203,N_3934,N_3826);
nand U5204 (N_5204,N_3572,N_3769);
and U5205 (N_5205,N_4682,N_4828);
or U5206 (N_5206,N_3465,N_3472);
and U5207 (N_5207,N_3837,N_2629);
xor U5208 (N_5208,N_4841,N_3549);
nand U5209 (N_5209,N_4355,N_3169);
or U5210 (N_5210,N_4614,N_3456);
or U5211 (N_5211,N_4345,N_4045);
nor U5212 (N_5212,N_3113,N_4640);
xor U5213 (N_5213,N_4648,N_2875);
and U5214 (N_5214,N_4683,N_2710);
and U5215 (N_5215,N_2623,N_2905);
or U5216 (N_5216,N_4586,N_4256);
nand U5217 (N_5217,N_2974,N_3101);
nor U5218 (N_5218,N_2796,N_4977);
nor U5219 (N_5219,N_2981,N_4738);
nor U5220 (N_5220,N_3425,N_4311);
or U5221 (N_5221,N_3834,N_4086);
or U5222 (N_5222,N_3052,N_4950);
xor U5223 (N_5223,N_3940,N_4213);
nand U5224 (N_5224,N_2686,N_2827);
nor U5225 (N_5225,N_2712,N_3768);
or U5226 (N_5226,N_4925,N_3217);
or U5227 (N_5227,N_4866,N_4309);
xnor U5228 (N_5228,N_3412,N_3841);
or U5229 (N_5229,N_2759,N_3381);
xor U5230 (N_5230,N_3624,N_2860);
xnor U5231 (N_5231,N_2508,N_3895);
or U5232 (N_5232,N_3114,N_4784);
and U5233 (N_5233,N_3301,N_4385);
or U5234 (N_5234,N_3439,N_2952);
nor U5235 (N_5235,N_3975,N_3014);
or U5236 (N_5236,N_4690,N_3061);
nor U5237 (N_5237,N_3812,N_4214);
nor U5238 (N_5238,N_4633,N_3621);
nor U5239 (N_5239,N_2583,N_2619);
and U5240 (N_5240,N_4065,N_2725);
nor U5241 (N_5241,N_3478,N_3565);
nand U5242 (N_5242,N_4706,N_2977);
or U5243 (N_5243,N_4193,N_3390);
nor U5244 (N_5244,N_3952,N_3133);
nor U5245 (N_5245,N_4739,N_3025);
nand U5246 (N_5246,N_2737,N_2683);
and U5247 (N_5247,N_2540,N_4545);
or U5248 (N_5248,N_4475,N_3395);
and U5249 (N_5249,N_3442,N_3462);
and U5250 (N_5250,N_4175,N_2896);
or U5251 (N_5251,N_3063,N_4524);
nand U5252 (N_5252,N_4717,N_3128);
or U5253 (N_5253,N_2748,N_2902);
nand U5254 (N_5254,N_3627,N_4552);
and U5255 (N_5255,N_4382,N_2704);
nand U5256 (N_5256,N_4757,N_4101);
and U5257 (N_5257,N_2838,N_4616);
nor U5258 (N_5258,N_2983,N_2665);
xor U5259 (N_5259,N_4300,N_4028);
and U5260 (N_5260,N_2872,N_3116);
nand U5261 (N_5261,N_3701,N_3578);
nor U5262 (N_5262,N_3482,N_4770);
or U5263 (N_5263,N_2828,N_2915);
nor U5264 (N_5264,N_3986,N_3319);
nand U5265 (N_5265,N_3770,N_3823);
or U5266 (N_5266,N_4001,N_3538);
and U5267 (N_5267,N_2520,N_4237);
and U5268 (N_5268,N_4902,N_3672);
nor U5269 (N_5269,N_4653,N_3900);
and U5270 (N_5270,N_4911,N_3613);
or U5271 (N_5271,N_4985,N_2613);
nand U5272 (N_5272,N_2503,N_2649);
nor U5273 (N_5273,N_2539,N_3213);
nand U5274 (N_5274,N_3773,N_4680);
nand U5275 (N_5275,N_4088,N_3633);
and U5276 (N_5276,N_2962,N_4468);
and U5277 (N_5277,N_3897,N_3098);
nand U5278 (N_5278,N_3057,N_3984);
nand U5279 (N_5279,N_3221,N_4401);
or U5280 (N_5280,N_3451,N_3027);
nand U5281 (N_5281,N_4940,N_4244);
and U5282 (N_5282,N_2970,N_4875);
or U5283 (N_5283,N_4909,N_4407);
or U5284 (N_5284,N_4796,N_2928);
nor U5285 (N_5285,N_4238,N_3313);
nand U5286 (N_5286,N_3751,N_2862);
or U5287 (N_5287,N_4126,N_4270);
or U5288 (N_5288,N_3048,N_4060);
or U5289 (N_5289,N_3151,N_4697);
xor U5290 (N_5290,N_4812,N_4096);
or U5291 (N_5291,N_3779,N_3726);
nand U5292 (N_5292,N_4581,N_3433);
nor U5293 (N_5293,N_3032,N_4069);
xnor U5294 (N_5294,N_3310,N_4712);
nand U5295 (N_5295,N_3214,N_3123);
and U5296 (N_5296,N_2559,N_4589);
and U5297 (N_5297,N_3523,N_4044);
nand U5298 (N_5298,N_3056,N_2885);
nand U5299 (N_5299,N_2808,N_4813);
nand U5300 (N_5300,N_3776,N_4947);
or U5301 (N_5301,N_3019,N_4668);
nor U5302 (N_5302,N_4929,N_4792);
or U5303 (N_5303,N_4710,N_4151);
nand U5304 (N_5304,N_4384,N_3000);
nor U5305 (N_5305,N_3535,N_2682);
or U5306 (N_5306,N_2866,N_3298);
nor U5307 (N_5307,N_3903,N_4976);
and U5308 (N_5308,N_2550,N_4937);
nor U5309 (N_5309,N_3747,N_4144);
nor U5310 (N_5310,N_3687,N_3248);
nand U5311 (N_5311,N_3740,N_4450);
nor U5312 (N_5312,N_3597,N_3473);
nor U5313 (N_5313,N_4530,N_2829);
nand U5314 (N_5314,N_2617,N_3575);
and U5315 (N_5315,N_4758,N_3234);
nand U5316 (N_5316,N_4290,N_3899);
or U5317 (N_5317,N_3949,N_3145);
xor U5318 (N_5318,N_3318,N_3361);
xor U5319 (N_5319,N_2987,N_4989);
nand U5320 (N_5320,N_4816,N_2768);
and U5321 (N_5321,N_4034,N_2563);
and U5322 (N_5322,N_3948,N_3675);
and U5323 (N_5323,N_4003,N_4833);
nand U5324 (N_5324,N_3496,N_4307);
nor U5325 (N_5325,N_2931,N_4085);
or U5326 (N_5326,N_4727,N_4898);
and U5327 (N_5327,N_2596,N_3605);
or U5328 (N_5328,N_3303,N_4629);
or U5329 (N_5329,N_3844,N_2883);
and U5330 (N_5330,N_3521,N_4320);
nor U5331 (N_5331,N_4729,N_3388);
nand U5332 (N_5332,N_3271,N_3607);
and U5333 (N_5333,N_4627,N_3667);
nor U5334 (N_5334,N_2543,N_2523);
nand U5335 (N_5335,N_4437,N_3083);
nand U5336 (N_5336,N_4996,N_4075);
and U5337 (N_5337,N_3539,N_3699);
nand U5338 (N_5338,N_2971,N_4510);
or U5339 (N_5339,N_4781,N_4624);
or U5340 (N_5340,N_4730,N_3269);
nand U5341 (N_5341,N_3432,N_4655);
and U5342 (N_5342,N_3788,N_4645);
nand U5343 (N_5343,N_3106,N_4883);
nor U5344 (N_5344,N_3552,N_2724);
xnor U5345 (N_5345,N_4141,N_4809);
nor U5346 (N_5346,N_3577,N_2919);
nand U5347 (N_5347,N_3711,N_3656);
xor U5348 (N_5348,N_2614,N_4817);
nand U5349 (N_5349,N_3275,N_2934);
nor U5350 (N_5350,N_4877,N_3131);
nand U5351 (N_5351,N_4895,N_4800);
nand U5352 (N_5352,N_4099,N_4373);
or U5353 (N_5353,N_3674,N_4111);
and U5354 (N_5354,N_3838,N_4491);
and U5355 (N_5355,N_4539,N_3742);
and U5356 (N_5356,N_4810,N_4274);
and U5357 (N_5357,N_4846,N_4466);
nand U5358 (N_5358,N_4849,N_4170);
nor U5359 (N_5359,N_3136,N_3080);
or U5360 (N_5360,N_2957,N_4752);
and U5361 (N_5361,N_4830,N_3871);
nor U5362 (N_5362,N_4497,N_2639);
nand U5363 (N_5363,N_2925,N_2727);
nand U5364 (N_5364,N_3828,N_3930);
nor U5365 (N_5365,N_4997,N_3176);
and U5366 (N_5366,N_4639,N_4625);
and U5367 (N_5367,N_4132,N_2871);
xnor U5368 (N_5368,N_2602,N_2929);
nor U5369 (N_5369,N_2666,N_4271);
xnor U5370 (N_5370,N_4232,N_3541);
nand U5371 (N_5371,N_3825,N_2773);
or U5372 (N_5372,N_2560,N_4029);
and U5373 (N_5373,N_4352,N_3878);
or U5374 (N_5374,N_2552,N_4139);
or U5375 (N_5375,N_3750,N_3759);
nor U5376 (N_5376,N_4476,N_2876);
and U5377 (N_5377,N_4462,N_4714);
nor U5378 (N_5378,N_4631,N_4516);
nand U5379 (N_5379,N_3323,N_3688);
nor U5380 (N_5380,N_4481,N_3845);
and U5381 (N_5381,N_3308,N_4439);
nand U5382 (N_5382,N_3907,N_4982);
and U5383 (N_5383,N_3926,N_4184);
nor U5384 (N_5384,N_4150,N_4285);
or U5385 (N_5385,N_4236,N_3695);
nand U5386 (N_5386,N_3421,N_4762);
nor U5387 (N_5387,N_2736,N_4692);
or U5388 (N_5388,N_4635,N_3588);
nand U5389 (N_5389,N_3691,N_4040);
or U5390 (N_5390,N_3517,N_2966);
or U5391 (N_5391,N_4924,N_3210);
or U5392 (N_5392,N_2622,N_4646);
xor U5393 (N_5393,N_2516,N_3702);
nor U5394 (N_5394,N_3718,N_4293);
and U5395 (N_5395,N_4482,N_4785);
xor U5396 (N_5396,N_3991,N_4297);
nor U5397 (N_5397,N_4856,N_3239);
nor U5398 (N_5398,N_2511,N_3162);
nor U5399 (N_5399,N_3126,N_3910);
nor U5400 (N_5400,N_4962,N_2893);
nand U5401 (N_5401,N_3460,N_3321);
or U5402 (N_5402,N_4328,N_3377);
and U5403 (N_5403,N_3348,N_4110);
and U5404 (N_5404,N_3504,N_3732);
nand U5405 (N_5405,N_4018,N_4484);
and U5406 (N_5406,N_2595,N_2636);
or U5407 (N_5407,N_2518,N_3513);
and U5408 (N_5408,N_4025,N_4394);
or U5409 (N_5409,N_2755,N_3865);
nand U5410 (N_5410,N_4208,N_3534);
or U5411 (N_5411,N_3047,N_3105);
and U5412 (N_5412,N_3911,N_2822);
nand U5413 (N_5413,N_3102,N_2610);
nand U5414 (N_5414,N_4528,N_2705);
or U5415 (N_5415,N_4414,N_3064);
and U5416 (N_5416,N_3645,N_3971);
nand U5417 (N_5417,N_3677,N_4226);
or U5418 (N_5418,N_4316,N_2956);
nand U5419 (N_5419,N_2963,N_2820);
nor U5420 (N_5420,N_4606,N_2898);
nor U5421 (N_5421,N_4036,N_3380);
or U5422 (N_5422,N_4312,N_4897);
nor U5423 (N_5423,N_3983,N_4957);
xnor U5424 (N_5424,N_4314,N_2731);
nand U5425 (N_5425,N_3491,N_2967);
nand U5426 (N_5426,N_4227,N_2935);
nand U5427 (N_5427,N_4177,N_3376);
nor U5428 (N_5428,N_4402,N_3743);
and U5429 (N_5429,N_3119,N_4489);
nand U5430 (N_5430,N_4622,N_4534);
and U5431 (N_5431,N_3207,N_2624);
or U5432 (N_5432,N_4863,N_4842);
nor U5433 (N_5433,N_2843,N_3919);
and U5434 (N_5434,N_2993,N_4751);
nor U5435 (N_5435,N_3704,N_2799);
xor U5436 (N_5436,N_2973,N_3516);
nand U5437 (N_5437,N_2817,N_2659);
xnor U5438 (N_5438,N_3345,N_3707);
or U5439 (N_5439,N_3874,N_4262);
or U5440 (N_5440,N_3661,N_3599);
nor U5441 (N_5441,N_3197,N_4790);
nand U5442 (N_5442,N_3935,N_2840);
xor U5443 (N_5443,N_3938,N_4910);
nand U5444 (N_5444,N_3941,N_2648);
and U5445 (N_5445,N_4289,N_4562);
nor U5446 (N_5446,N_4826,N_4901);
or U5447 (N_5447,N_3586,N_2515);
xor U5448 (N_5448,N_4847,N_3033);
nor U5449 (N_5449,N_3651,N_4876);
nor U5450 (N_5450,N_3725,N_3371);
xor U5451 (N_5451,N_2978,N_3564);
nor U5452 (N_5452,N_3585,N_4362);
xnor U5453 (N_5453,N_4171,N_3507);
nand U5454 (N_5454,N_3135,N_3916);
nor U5455 (N_5455,N_3004,N_4611);
or U5456 (N_5456,N_3163,N_4713);
nor U5457 (N_5457,N_2726,N_3490);
or U5458 (N_5458,N_3398,N_4163);
xnor U5459 (N_5459,N_4221,N_2743);
or U5460 (N_5460,N_3065,N_3322);
nand U5461 (N_5461,N_4196,N_3962);
and U5462 (N_5462,N_3850,N_3499);
or U5463 (N_5463,N_3787,N_4064);
or U5464 (N_5464,N_4953,N_3847);
nand U5465 (N_5465,N_3959,N_3339);
xnor U5466 (N_5466,N_4936,N_2572);
nand U5467 (N_5467,N_4746,N_3617);
nand U5468 (N_5468,N_4601,N_3194);
or U5469 (N_5469,N_3266,N_2776);
or U5470 (N_5470,N_4861,N_4191);
xor U5471 (N_5471,N_3710,N_3684);
nand U5472 (N_5472,N_2815,N_4425);
xnor U5473 (N_5473,N_2570,N_4890);
nor U5474 (N_5474,N_3591,N_3094);
nor U5475 (N_5475,N_3045,N_4827);
xnor U5476 (N_5476,N_3831,N_3998);
nor U5477 (N_5477,N_3625,N_4416);
nor U5478 (N_5478,N_3069,N_3686);
nand U5479 (N_5479,N_4965,N_3494);
and U5480 (N_5480,N_4000,N_3892);
nor U5481 (N_5481,N_3664,N_2812);
nand U5482 (N_5482,N_3190,N_4368);
or U5483 (N_5483,N_2601,N_4913);
nand U5484 (N_5484,N_4375,N_3579);
nor U5485 (N_5485,N_3115,N_4443);
or U5486 (N_5486,N_3973,N_4051);
and U5487 (N_5487,N_4664,N_3921);
nor U5488 (N_5488,N_4522,N_4766);
nand U5489 (N_5489,N_2877,N_3441);
nand U5490 (N_5490,N_3141,N_4448);
and U5491 (N_5491,N_4979,N_4716);
nor U5492 (N_5492,N_3009,N_4386);
xor U5493 (N_5493,N_3366,N_3925);
xnor U5494 (N_5494,N_2746,N_4203);
nand U5495 (N_5495,N_3160,N_4544);
and U5496 (N_5496,N_3121,N_3283);
nand U5497 (N_5497,N_3563,N_3995);
or U5498 (N_5498,N_3344,N_4617);
and U5499 (N_5499,N_3498,N_3035);
nor U5500 (N_5500,N_4774,N_4991);
and U5501 (N_5501,N_4551,N_4840);
nor U5502 (N_5502,N_3923,N_4546);
nor U5503 (N_5503,N_3955,N_4046);
nand U5504 (N_5504,N_3474,N_2500);
nor U5505 (N_5505,N_3284,N_3138);
nand U5506 (N_5506,N_4494,N_3374);
nor U5507 (N_5507,N_2647,N_4174);
nand U5508 (N_5508,N_4310,N_2567);
nand U5509 (N_5509,N_3008,N_4725);
or U5510 (N_5510,N_4162,N_4391);
and U5511 (N_5511,N_3898,N_4848);
nor U5512 (N_5512,N_4187,N_3333);
or U5513 (N_5513,N_4776,N_4914);
nand U5514 (N_5514,N_4899,N_3852);
or U5515 (N_5515,N_2936,N_2519);
and U5516 (N_5516,N_4123,N_4637);
xor U5517 (N_5517,N_3860,N_2545);
and U5518 (N_5518,N_3137,N_4090);
nor U5519 (N_5519,N_4092,N_3849);
nand U5520 (N_5520,N_4870,N_3520);
or U5521 (N_5521,N_4839,N_4951);
or U5522 (N_5522,N_3463,N_4740);
and U5523 (N_5523,N_2789,N_3683);
nand U5524 (N_5524,N_3763,N_4764);
or U5525 (N_5525,N_4296,N_3224);
nand U5526 (N_5526,N_4808,N_3576);
nor U5527 (N_5527,N_4882,N_3612);
or U5528 (N_5528,N_4076,N_4365);
xor U5529 (N_5529,N_3786,N_4173);
nor U5530 (N_5530,N_4575,N_4743);
or U5531 (N_5531,N_2625,N_4734);
or U5532 (N_5532,N_3861,N_3653);
nor U5533 (N_5533,N_4241,N_2895);
xnor U5534 (N_5534,N_4906,N_3784);
nand U5535 (N_5535,N_4487,N_3108);
xnor U5536 (N_5536,N_3954,N_4814);
nand U5537 (N_5537,N_4417,N_3185);
nor U5538 (N_5538,N_3889,N_4855);
nor U5539 (N_5539,N_3383,N_4675);
and U5540 (N_5540,N_3434,N_4698);
nand U5541 (N_5541,N_3175,N_2950);
and U5542 (N_5542,N_4031,N_3809);
and U5543 (N_5543,N_3988,N_4474);
nand U5544 (N_5544,N_3846,N_4054);
or U5545 (N_5545,N_4618,N_3487);
nor U5546 (N_5546,N_4234,N_3343);
nor U5547 (N_5547,N_4103,N_2612);
nor U5548 (N_5548,N_4463,N_4473);
and U5549 (N_5549,N_4521,N_3509);
and U5550 (N_5550,N_4915,N_3560);
nand U5551 (N_5551,N_4107,N_4943);
nand U5552 (N_5552,N_2927,N_3501);
or U5553 (N_5553,N_3529,N_4638);
nand U5554 (N_5554,N_2752,N_3391);
and U5555 (N_5555,N_4797,N_4189);
or U5556 (N_5556,N_2579,N_3570);
or U5557 (N_5557,N_3696,N_4672);
nand U5558 (N_5558,N_3405,N_3694);
xor U5559 (N_5559,N_4926,N_4845);
nand U5560 (N_5560,N_2568,N_3255);
or U5561 (N_5561,N_4952,N_4264);
nor U5562 (N_5562,N_4858,N_3580);
nand U5563 (N_5563,N_3894,N_4403);
and U5564 (N_5564,N_2879,N_2878);
nor U5565 (N_5565,N_4457,N_3615);
nand U5566 (N_5566,N_4479,N_3304);
nand U5567 (N_5567,N_3713,N_4824);
and U5568 (N_5568,N_3663,N_4853);
nand U5569 (N_5569,N_2801,N_4027);
or U5570 (N_5570,N_2679,N_2653);
nor U5571 (N_5571,N_3382,N_4283);
and U5572 (N_5572,N_4465,N_2800);
or U5573 (N_5573,N_3164,N_2923);
nand U5574 (N_5574,N_2677,N_3413);
nor U5575 (N_5575,N_4277,N_4119);
nand U5576 (N_5576,N_4333,N_4878);
nor U5577 (N_5577,N_4922,N_3294);
nor U5578 (N_5578,N_3222,N_3804);
nand U5579 (N_5579,N_3716,N_2904);
nand U5580 (N_5580,N_4599,N_2538);
nor U5581 (N_5581,N_4421,N_3085);
nor U5582 (N_5582,N_2767,N_2903);
nand U5583 (N_5583,N_4609,N_2678);
nor U5584 (N_5584,N_2996,N_4750);
xor U5585 (N_5585,N_4330,N_2945);
or U5586 (N_5586,N_3182,N_4249);
xor U5587 (N_5587,N_2591,N_3475);
xnor U5588 (N_5588,N_4412,N_2853);
or U5589 (N_5589,N_4657,N_3843);
xor U5590 (N_5590,N_2836,N_3031);
nand U5591 (N_5591,N_4341,N_3177);
xor U5592 (N_5592,N_2958,N_4426);
or U5593 (N_5593,N_3155,N_4693);
nand U5594 (N_5594,N_4243,N_4954);
nor U5595 (N_5595,N_3970,N_3670);
nand U5596 (N_5596,N_2604,N_2702);
or U5597 (N_5597,N_3592,N_4127);
nand U5598 (N_5598,N_4674,N_2889);
or U5599 (N_5599,N_2620,N_4715);
nand U5600 (N_5600,N_4026,N_4975);
nor U5601 (N_5601,N_3781,N_4104);
and U5602 (N_5602,N_4089,N_3316);
and U5603 (N_5603,N_4512,N_3783);
or U5604 (N_5604,N_2857,N_4660);
and U5605 (N_5605,N_2998,N_3917);
nand U5606 (N_5606,N_3546,N_4002);
nand U5607 (N_5607,N_3120,N_2920);
or U5608 (N_5608,N_4536,N_2632);
and U5609 (N_5609,N_4744,N_4869);
or U5610 (N_5610,N_2646,N_3937);
nand U5611 (N_5611,N_2858,N_4502);
nand U5612 (N_5612,N_4125,N_4050);
nand U5613 (N_5613,N_4634,N_4364);
and U5614 (N_5614,N_4923,N_3363);
or U5615 (N_5615,N_4490,N_2937);
and U5616 (N_5616,N_4287,N_3324);
and U5617 (N_5617,N_4579,N_4904);
or U5618 (N_5618,N_3830,N_3774);
nor U5619 (N_5619,N_4255,N_2944);
nand U5620 (N_5620,N_2616,N_2750);
and U5621 (N_5621,N_3144,N_4376);
or U5622 (N_5622,N_4907,N_4043);
and U5623 (N_5623,N_2891,N_3772);
nand U5624 (N_5624,N_4348,N_4547);
nand U5625 (N_5625,N_4138,N_4580);
nand U5626 (N_5626,N_4888,N_4588);
nand U5627 (N_5627,N_2779,N_4941);
nor U5628 (N_5628,N_4596,N_2761);
and U5629 (N_5629,N_4275,N_3720);
or U5630 (N_5630,N_4279,N_4114);
and U5631 (N_5631,N_3293,N_4379);
or U5632 (N_5632,N_3428,N_4073);
nand U5633 (N_5633,N_3811,N_2997);
and U5634 (N_5634,N_3542,N_3384);
nand U5635 (N_5635,N_4610,N_4102);
nor U5636 (N_5636,N_3851,N_3946);
nor U5637 (N_5637,N_3668,N_4887);
nor U5638 (N_5638,N_2656,N_3495);
nand U5639 (N_5639,N_4723,N_3459);
or U5640 (N_5640,N_2995,N_4077);
and U5641 (N_5641,N_3835,N_3676);
and U5642 (N_5642,N_2600,N_3530);
nor U5643 (N_5643,N_3142,N_4771);
or U5644 (N_5644,N_3931,N_3236);
and U5645 (N_5645,N_4932,N_3658);
and U5646 (N_5646,N_4056,N_3010);
and U5647 (N_5647,N_3039,N_2707);
nor U5648 (N_5648,N_4278,N_4295);
xor U5649 (N_5649,N_4548,N_2504);
nand U5650 (N_5650,N_2803,N_3802);
and U5651 (N_5651,N_2689,N_4231);
or U5652 (N_5652,N_3084,N_3964);
nor U5653 (N_5653,N_4229,N_4799);
and U5654 (N_5654,N_3330,N_4356);
xnor U5655 (N_5655,N_3558,N_2701);
nand U5656 (N_5656,N_3346,N_4928);
nor U5657 (N_5657,N_3159,N_3189);
or U5658 (N_5658,N_3006,N_2932);
nand U5659 (N_5659,N_3368,N_2753);
or U5660 (N_5660,N_2825,N_3545);
nand U5661 (N_5661,N_4325,N_3470);
or U5662 (N_5662,N_2522,N_4204);
and U5663 (N_5663,N_2658,N_4974);
and U5664 (N_5664,N_2790,N_4294);
nor U5665 (N_5665,N_4334,N_2798);
or U5666 (N_5666,N_4844,N_3928);
xor U5667 (N_5667,N_4689,N_4587);
nand U5668 (N_5668,N_3401,N_4529);
or U5669 (N_5669,N_4118,N_3180);
nor U5670 (N_5670,N_3598,N_3302);
and U5671 (N_5671,N_4677,N_4210);
nand U5672 (N_5672,N_4868,N_3208);
xor U5673 (N_5673,N_2739,N_4992);
and U5674 (N_5674,N_4772,N_4687);
or U5675 (N_5675,N_4434,N_3104);
nor U5676 (N_5676,N_4891,N_3226);
xor U5677 (N_5677,N_4470,N_2609);
and U5678 (N_5678,N_3295,N_4315);
nor U5679 (N_5679,N_2880,N_3258);
or U5680 (N_5680,N_4971,N_3864);
nand U5681 (N_5681,N_3797,N_3966);
nor U5682 (N_5682,N_4673,N_2668);
xnor U5683 (N_5683,N_3075,N_4935);
nor U5684 (N_5684,N_4215,N_4068);
or U5685 (N_5685,N_4240,N_3077);
xor U5686 (N_5686,N_3727,N_4822);
nand U5687 (N_5687,N_4216,N_2575);
xor U5688 (N_5688,N_4748,N_4128);
nand U5689 (N_5689,N_3639,N_4166);
and U5690 (N_5690,N_2949,N_2948);
or U5691 (N_5691,N_3369,N_3762);
and U5692 (N_5692,N_4133,N_2716);
or U5693 (N_5693,N_2606,N_3249);
and U5694 (N_5694,N_4819,N_3526);
xnor U5695 (N_5695,N_4327,N_3842);
nor U5696 (N_5696,N_3178,N_4021);
nor U5697 (N_5697,N_3251,N_4207);
nand U5698 (N_5698,N_3987,N_4742);
or U5699 (N_5699,N_4222,N_4700);
or U5700 (N_5700,N_4956,N_3168);
nand U5701 (N_5701,N_2742,N_2984);
nand U5702 (N_5702,N_3274,N_2867);
or U5703 (N_5703,N_3386,N_3796);
xnor U5704 (N_5704,N_3882,N_2571);
nor U5705 (N_5705,N_3896,N_4009);
nor U5706 (N_5706,N_2741,N_4097);
nand U5707 (N_5707,N_3238,N_4436);
or U5708 (N_5708,N_4573,N_4093);
or U5709 (N_5709,N_3247,N_3993);
nor U5710 (N_5710,N_3714,N_3479);
nand U5711 (N_5711,N_4659,N_4292);
or U5712 (N_5712,N_3960,N_3112);
xnor U5713 (N_5713,N_3873,N_2607);
or U5714 (N_5714,N_4349,N_3567);
nor U5715 (N_5715,N_2587,N_4686);
xnor U5716 (N_5716,N_4432,N_2881);
or U5717 (N_5717,N_4964,N_3480);
nand U5718 (N_5718,N_3452,N_3079);
nand U5719 (N_5719,N_4281,N_4321);
and U5720 (N_5720,N_3868,N_3756);
nor U5721 (N_5721,N_4340,N_3272);
xnor U5722 (N_5722,N_3416,N_3205);
or U5723 (N_5723,N_4366,N_4254);
xnor U5724 (N_5724,N_3183,N_2955);
nand U5725 (N_5725,N_3775,N_3245);
xnor U5726 (N_5726,N_4094,N_4619);
nor U5727 (N_5727,N_3011,N_2947);
or U5728 (N_5728,N_4100,N_2744);
or U5729 (N_5729,N_3767,N_3070);
or U5730 (N_5730,N_4949,N_2529);
nand U5731 (N_5731,N_2806,N_3187);
nor U5732 (N_5732,N_3989,N_4178);
nand U5733 (N_5733,N_2793,N_3179);
nand U5734 (N_5734,N_3054,N_2722);
nor U5735 (N_5735,N_2535,N_4410);
nand U5736 (N_5736,N_4335,N_3601);
nand U5737 (N_5737,N_4867,N_3227);
nand U5738 (N_5738,N_3997,N_3270);
xnor U5739 (N_5739,N_3614,N_3915);
nand U5740 (N_5740,N_3746,N_3813);
and U5741 (N_5741,N_3081,N_4600);
nand U5742 (N_5742,N_3933,N_3464);
nand U5743 (N_5743,N_3148,N_4968);
nor U5744 (N_5744,N_3282,N_3466);
xnor U5745 (N_5745,N_3044,N_4129);
nand U5746 (N_5746,N_4984,N_2907);
and U5747 (N_5747,N_2548,N_4015);
xnor U5748 (N_5748,N_3109,N_3853);
nor U5749 (N_5749,N_3392,N_2811);
xor U5750 (N_5750,N_3408,N_4142);
or U5751 (N_5751,N_3041,N_3922);
xnor U5752 (N_5752,N_2901,N_4721);
or U5753 (N_5753,N_4889,N_3216);
nor U5754 (N_5754,N_3440,N_3635);
xnor U5755 (N_5755,N_4011,N_4555);
xnor U5756 (N_5756,N_2630,N_4429);
xor U5757 (N_5757,N_2795,N_2684);
xnor U5758 (N_5758,N_3422,N_3780);
nand U5759 (N_5759,N_3082,N_3854);
nand U5760 (N_5760,N_2527,N_3231);
or U5761 (N_5761,N_4520,N_3254);
nand U5762 (N_5762,N_2662,N_4495);
nand U5763 (N_5763,N_2611,N_3058);
nand U5764 (N_5764,N_4319,N_3410);
nor U5765 (N_5765,N_3170,N_4156);
nand U5766 (N_5766,N_2758,N_3927);
or U5767 (N_5767,N_3315,N_4030);
and U5768 (N_5768,N_4543,N_3150);
or U5769 (N_5769,N_2830,N_4055);
xor U5770 (N_5770,N_2887,N_2850);
or U5771 (N_5771,N_3693,N_2638);
and U5772 (N_5772,N_3445,N_2943);
nor U5773 (N_5773,N_3869,N_4986);
nand U5774 (N_5774,N_2834,N_4843);
and U5775 (N_5775,N_2762,N_3556);
nand U5776 (N_5776,N_4557,N_4008);
and U5777 (N_5777,N_4933,N_4148);
or U5778 (N_5778,N_3739,N_3060);
nand U5779 (N_5779,N_3799,N_3681);
and U5780 (N_5780,N_4896,N_3939);
nor U5781 (N_5781,N_4688,N_4787);
or U5782 (N_5782,N_4313,N_3544);
xor U5783 (N_5783,N_2835,N_3088);
nor U5784 (N_5784,N_2599,N_4299);
or U5785 (N_5785,N_3692,N_2873);
and U5786 (N_5786,N_3709,N_3431);
xnor U5787 (N_5787,N_3471,N_2697);
nand U5788 (N_5788,N_3909,N_4807);
nor U5789 (N_5789,N_2694,N_3761);
and U5790 (N_5790,N_4284,N_4168);
nor U5791 (N_5791,N_4852,N_4070);
and U5792 (N_5792,N_4140,N_3867);
or U5793 (N_5793,N_4472,N_2549);
and U5794 (N_5794,N_4554,N_2708);
and U5795 (N_5795,N_4172,N_3200);
nor U5796 (N_5796,N_4419,N_4820);
nor U5797 (N_5797,N_3790,N_2734);
or U5798 (N_5798,N_3042,N_3584);
or U5799 (N_5799,N_3737,N_3378);
nand U5800 (N_5800,N_4433,N_3914);
nor U5801 (N_5801,N_2831,N_4550);
and U5802 (N_5802,N_3650,N_4572);
or U5803 (N_5803,N_2660,N_3087);
nor U5804 (N_5804,N_2908,N_4881);
and U5805 (N_5805,N_3963,N_4273);
or U5806 (N_5806,N_3335,N_4291);
or U5807 (N_5807,N_3240,N_4815);
or U5808 (N_5808,N_3611,N_4201);
nand U5809 (N_5809,N_4338,N_3631);
nor U5810 (N_5810,N_4113,N_4415);
nand U5811 (N_5811,N_4767,N_3808);
nor U5812 (N_5812,N_4367,N_3789);
nor U5813 (N_5813,N_3807,N_2818);
and U5814 (N_5814,N_3652,N_2810);
xor U5815 (N_5815,N_4779,N_3888);
or U5816 (N_5816,N_2807,N_3389);
nand U5817 (N_5817,N_3800,N_4301);
or U5818 (N_5818,N_3296,N_4298);
xnor U5819 (N_5819,N_4563,N_4998);
nand U5820 (N_5820,N_4420,N_4083);
nand U5821 (N_5821,N_3859,N_4825);
nor U5822 (N_5822,N_4514,N_2869);
nand U5823 (N_5823,N_4351,N_4124);
and U5824 (N_5824,N_3062,N_3469);
nor U5825 (N_5825,N_3936,N_2849);
or U5826 (N_5826,N_4067,N_4061);
or U5827 (N_5827,N_4592,N_3095);
and U5828 (N_5828,N_2969,N_4263);
nand U5829 (N_5829,N_4461,N_4652);
xor U5830 (N_5830,N_4245,N_3978);
or U5831 (N_5831,N_4095,N_2786);
or U5832 (N_5832,N_4084,N_3001);
nor U5833 (N_5833,N_3673,N_4445);
and U5834 (N_5834,N_2585,N_4306);
or U5835 (N_5835,N_3902,N_3253);
nor U5836 (N_5836,N_3942,N_3582);
nand U5837 (N_5837,N_2562,N_3757);
or U5838 (N_5838,N_3446,N_3454);
or U5839 (N_5839,N_3690,N_3174);
nand U5840 (N_5840,N_4880,N_4626);
nand U5841 (N_5841,N_2593,N_2941);
nor U5842 (N_5842,N_4802,N_2510);
nor U5843 (N_5843,N_3181,N_3708);
or U5844 (N_5844,N_2685,N_3265);
nand U5845 (N_5845,N_4159,N_4948);
nor U5846 (N_5846,N_3309,N_3051);
or U5847 (N_5847,N_3866,N_3581);
xnor U5848 (N_5848,N_3648,N_2863);
nand U5849 (N_5849,N_4722,N_3228);
nand U5850 (N_5850,N_3736,N_4190);
or U5851 (N_5851,N_4458,N_2557);
nand U5852 (N_5852,N_4116,N_4200);
or U5853 (N_5853,N_3152,N_3458);
nand U5854 (N_5854,N_4057,N_2621);
or U5855 (N_5855,N_4380,N_4679);
nor U5856 (N_5856,N_3029,N_3007);
xnor U5857 (N_5857,N_2938,N_3730);
and U5858 (N_5858,N_3777,N_3290);
or U5859 (N_5859,N_3124,N_4641);
and U5860 (N_5860,N_4523,N_4823);
nor U5861 (N_5861,N_2864,N_4775);
and U5862 (N_5862,N_2521,N_4398);
and U5863 (N_5863,N_3426,N_4662);
or U5864 (N_5864,N_4620,N_4591);
nand U5865 (N_5865,N_3848,N_3153);
nor U5866 (N_5866,N_3771,N_4343);
nand U5867 (N_5867,N_4370,N_4105);
or U5868 (N_5868,N_4578,N_2672);
and U5869 (N_5869,N_3527,N_3312);
nand U5870 (N_5870,N_3024,N_2699);
and U5871 (N_5871,N_3603,N_4658);
or U5872 (N_5872,N_2667,N_4276);
and U5873 (N_5873,N_4326,N_4691);
or U5874 (N_5874,N_2894,N_2899);
nand U5875 (N_5875,N_4553,N_4930);
nand U5876 (N_5876,N_4004,N_4235);
or U5877 (N_5877,N_4656,N_2546);
nor U5878 (N_5878,N_2637,N_2844);
nor U5879 (N_5879,N_2777,N_3020);
or U5880 (N_5880,N_4650,N_3906);
or U5881 (N_5881,N_3609,N_2942);
nor U5882 (N_5882,N_4360,N_3622);
and U5883 (N_5883,N_4905,N_4970);
nand U5884 (N_5884,N_4836,N_4186);
and U5885 (N_5885,N_3066,N_2537);
nor U5886 (N_5886,N_3092,N_4252);
nand U5887 (N_5887,N_4967,N_4078);
or U5888 (N_5888,N_2805,N_2633);
or U5889 (N_5889,N_4478,N_3418);
nand U5890 (N_5890,N_4137,N_4268);
nand U5891 (N_5891,N_2785,N_4438);
or U5892 (N_5892,N_3977,N_3566);
nor U5893 (N_5893,N_3729,N_3659);
or U5894 (N_5894,N_3250,N_3158);
nand U5895 (N_5895,N_4630,N_4442);
nor U5896 (N_5896,N_3957,N_3636);
nand U5897 (N_5897,N_4791,N_4504);
or U5898 (N_5898,N_3724,N_3268);
or U5899 (N_5899,N_4483,N_3161);
nand U5900 (N_5900,N_2663,N_3583);
xnor U5901 (N_5901,N_2693,N_2814);
and U5902 (N_5902,N_4732,N_4574);
and U5903 (N_5903,N_3619,N_4987);
nand U5904 (N_5904,N_3198,N_4990);
or U5905 (N_5905,N_4440,N_4741);
xor U5906 (N_5906,N_4667,N_4106);
or U5907 (N_5907,N_3016,N_3806);
and U5908 (N_5908,N_3026,N_4527);
nor U5909 (N_5909,N_2717,N_2589);
or U5910 (N_5910,N_3186,N_2965);
nor U5911 (N_5911,N_4805,N_2524);
nor U5912 (N_5912,N_2992,N_3292);
xnor U5913 (N_5913,N_4331,N_3219);
nand U5914 (N_5914,N_4961,N_3276);
and U5915 (N_5915,N_2897,N_4413);
and U5916 (N_5916,N_2816,N_4176);
nand U5917 (N_5917,N_4559,N_3394);
nand U5918 (N_5918,N_4651,N_2930);
nor U5919 (N_5919,N_2688,N_3351);
nand U5920 (N_5920,N_4121,N_3990);
nand U5921 (N_5921,N_3002,N_3457);
nor U5922 (N_5922,N_4576,N_4147);
nand U5923 (N_5923,N_3760,N_4993);
nor U5924 (N_5924,N_3602,N_3059);
or U5925 (N_5925,N_4765,N_3508);
or U5926 (N_5926,N_4063,N_4455);
nand U5927 (N_5927,N_3728,N_4339);
nor U5928 (N_5928,N_4195,N_4944);
nand U5929 (N_5929,N_3518,N_3968);
nand U5930 (N_5930,N_4665,N_4014);
or U5931 (N_5931,N_3072,N_4165);
nand U5932 (N_5932,N_4280,N_2854);
nor U5933 (N_5933,N_4406,N_4225);
and U5934 (N_5934,N_3510,N_3947);
or U5935 (N_5935,N_3402,N_3638);
and U5936 (N_5936,N_3484,N_2906);
or U5937 (N_5937,N_3191,N_2555);
nor U5938 (N_5938,N_3256,N_4703);
or U5939 (N_5939,N_4135,N_4242);
or U5940 (N_5940,N_2506,N_3540);
or U5941 (N_5941,N_3778,N_4496);
nor U5942 (N_5942,N_2783,N_2868);
or U5943 (N_5943,N_3979,N_3550);
nand U5944 (N_5944,N_3406,N_3655);
or U5945 (N_5945,N_4251,N_4253);
nor U5946 (N_5946,N_3733,N_3500);
nor U5947 (N_5947,N_4122,N_2914);
nor U5948 (N_5948,N_4160,N_2874);
nand U5949 (N_5949,N_3958,N_4711);
nor U5950 (N_5950,N_4873,N_2846);
and U5951 (N_5951,N_4577,N_2706);
nor U5952 (N_5952,N_4087,N_2530);
nor U5953 (N_5953,N_2655,N_3341);
or U5954 (N_5954,N_3110,N_2703);
nor U5955 (N_5955,N_2890,N_2590);
nand U5956 (N_5956,N_3204,N_4157);
nor U5957 (N_5957,N_3857,N_2770);
or U5958 (N_5958,N_4390,N_3887);
nand U5959 (N_5959,N_4485,N_3362);
and U5960 (N_5960,N_2588,N_2769);
nand U5961 (N_5961,N_4503,N_2573);
or U5962 (N_5962,N_4513,N_2980);
xnor U5963 (N_5963,N_2542,N_4506);
xnor U5964 (N_5964,N_3554,N_2691);
nand U5965 (N_5965,N_4500,N_4942);
nand U5966 (N_5966,N_2766,N_4464);
nor U5967 (N_5967,N_3533,N_3259);
or U5968 (N_5968,N_3920,N_3017);
and U5969 (N_5969,N_4267,N_3932);
nor U5970 (N_5970,N_4773,N_2561);
or U5971 (N_5971,N_3220,N_3068);
xnor U5972 (N_5972,N_3801,N_4980);
and U5973 (N_5973,N_3647,N_3448);
nor U5974 (N_5974,N_2985,N_2855);
nor U5975 (N_5975,N_3053,N_3833);
and U5976 (N_5976,N_3195,N_4022);
nor U5977 (N_5977,N_3822,N_2802);
or U5978 (N_5978,N_3040,N_4541);
nand U5979 (N_5979,N_3013,N_4035);
and U5980 (N_5980,N_3328,N_2912);
nand U5981 (N_5981,N_4250,N_4670);
nand U5982 (N_5982,N_2709,N_3559);
and U5983 (N_5983,N_3785,N_4582);
nor U5984 (N_5984,N_4006,N_4777);
and U5985 (N_5985,N_4804,N_4451);
nor U5986 (N_5986,N_3536,N_4919);
or U5987 (N_5987,N_4449,N_2528);
and U5988 (N_5988,N_3297,N_2900);
xnor U5989 (N_5989,N_4983,N_4885);
nand U5990 (N_5990,N_3229,N_4363);
or U5991 (N_5991,N_3129,N_3055);
nand U5992 (N_5992,N_3616,N_2690);
nor U5993 (N_5993,N_4834,N_4430);
and U5994 (N_5994,N_4921,N_2961);
nor U5995 (N_5995,N_2695,N_4441);
or U5996 (N_5996,N_4570,N_4032);
and U5997 (N_5997,N_2721,N_2626);
nor U5998 (N_5998,N_3127,N_3814);
nand U5999 (N_5999,N_4871,N_4378);
or U6000 (N_6000,N_2782,N_4197);
and U6001 (N_6001,N_3680,N_3233);
and U6002 (N_6002,N_2720,N_4811);
or U6003 (N_6003,N_4361,N_4218);
or U6004 (N_6004,N_2640,N_3373);
and U6005 (N_6005,N_3202,N_2989);
xor U6006 (N_6006,N_4829,N_3156);
nand U6007 (N_6007,N_2547,N_3354);
and U6008 (N_6008,N_3630,N_4158);
and U6009 (N_6009,N_4505,N_4305);
nand U6010 (N_6010,N_2791,N_4399);
nand U6011 (N_6011,N_3443,N_4747);
nor U6012 (N_6012,N_3100,N_3803);
nand U6013 (N_6013,N_2674,N_3571);
and U6014 (N_6014,N_2837,N_4789);
nor U6015 (N_6015,N_4818,N_3134);
or U6016 (N_6016,N_3551,N_3881);
or U6017 (N_6017,N_3488,N_3557);
or U6018 (N_6018,N_3235,N_4960);
xor U6019 (N_6019,N_3858,N_3669);
nor U6020 (N_6020,N_4966,N_4701);
xor U6021 (N_6021,N_2870,N_2608);
nand U6022 (N_6022,N_2892,N_3367);
or U6023 (N_6023,N_4302,N_4260);
nand U6024 (N_6024,N_2723,N_4835);
or U6025 (N_6025,N_4202,N_4053);
or U6026 (N_6026,N_4538,N_3792);
nand U6027 (N_6027,N_2718,N_3880);
nor U6028 (N_6028,N_3415,N_3555);
and U6029 (N_6029,N_3286,N_4632);
nor U6030 (N_6030,N_3481,N_3912);
nand U6031 (N_6031,N_3287,N_4684);
and U6032 (N_6032,N_3244,N_2833);
or U6033 (N_6033,N_3634,N_2913);
xnor U6034 (N_6034,N_3764,N_3364);
nand U6035 (N_6035,N_3223,N_4459);
nor U6036 (N_6036,N_2886,N_4988);
or U6037 (N_6037,N_2671,N_3569);
or U6038 (N_6038,N_4007,N_3929);
and U6039 (N_6039,N_3263,N_3417);
and U6040 (N_6040,N_4154,N_4795);
xor U6041 (N_6041,N_2775,N_4145);
or U6042 (N_6042,N_3506,N_3722);
nand U6043 (N_6043,N_3349,N_4358);
or U6044 (N_6044,N_2910,N_3172);
nand U6045 (N_6045,N_3748,N_4024);
nor U6046 (N_6046,N_3166,N_3944);
nor U6047 (N_6047,N_3610,N_3721);
nor U6048 (N_6048,N_2804,N_3165);
nor U6049 (N_6049,N_4239,N_3595);
nand U6050 (N_6050,N_4567,N_3698);
and U6051 (N_6051,N_2792,N_3438);
and U6052 (N_6052,N_4212,N_4737);
nor U6053 (N_6053,N_4509,N_3981);
or U6054 (N_6054,N_4568,N_4643);
nor U6055 (N_6055,N_3278,N_2577);
or U6056 (N_6056,N_3143,N_4999);
nor U6057 (N_6057,N_3884,N_4261);
and U6058 (N_6058,N_3252,N_2847);
nor U6059 (N_6059,N_4381,N_3908);
nor U6060 (N_6060,N_3972,N_3840);
nor U6061 (N_6061,N_2990,N_4759);
xor U6062 (N_6062,N_3356,N_4803);
nor U6063 (N_6063,N_4453,N_4531);
and U6064 (N_6064,N_2918,N_3034);
and U6065 (N_6065,N_2592,N_3856);
nand U6066 (N_6066,N_4435,N_4602);
or U6067 (N_6067,N_3485,N_3281);
xnor U6068 (N_6068,N_3154,N_3203);
nor U6069 (N_6069,N_3347,N_3477);
nor U6070 (N_6070,N_4109,N_3357);
and U6071 (N_6071,N_2569,N_2884);
and U6072 (N_6072,N_4047,N_3427);
and U6073 (N_6073,N_3745,N_2856);
nand U6074 (N_6074,N_4719,N_3379);
or U6075 (N_6075,N_4005,N_3643);
and U6076 (N_6076,N_2763,N_3230);
and U6077 (N_6077,N_4037,N_2628);
or U6078 (N_6078,N_2921,N_3953);
or U6079 (N_6079,N_4608,N_3199);
nor U6080 (N_6080,N_3099,N_4079);
nand U6081 (N_6081,N_3350,N_4152);
nor U6082 (N_6082,N_3791,N_3877);
or U6083 (N_6083,N_3468,N_4318);
nand U6084 (N_6084,N_4324,N_4344);
and U6085 (N_6085,N_3277,N_3435);
and U6086 (N_6086,N_3904,N_3766);
nor U6087 (N_6087,N_4389,N_4864);
nand U6088 (N_6088,N_3503,N_4209);
nor U6089 (N_6089,N_4377,N_3620);
or U6090 (N_6090,N_3532,N_4754);
nor U6091 (N_6091,N_2657,N_3765);
and U6092 (N_6092,N_4317,N_3370);
nand U6093 (N_6093,N_4593,N_4955);
xnor U6094 (N_6094,N_2924,N_2514);
nand U6095 (N_6095,N_3340,N_4763);
nand U6096 (N_6096,N_4357,N_3279);
nor U6097 (N_6097,N_4400,N_2972);
and U6098 (N_6098,N_3817,N_3260);
or U6099 (N_6099,N_4016,N_3167);
or U6100 (N_6100,N_4353,N_3629);
or U6101 (N_6101,N_4585,N_2581);
or U6102 (N_6102,N_4707,N_2517);
nor U6103 (N_6103,N_4493,N_2502);
nor U6104 (N_6104,N_4565,N_3171);
xnor U6105 (N_6105,N_2580,N_2642);
nor U6106 (N_6106,N_3184,N_4604);
or U6107 (N_6107,N_4444,N_4498);
or U6108 (N_6108,N_4994,N_3122);
or U6109 (N_6109,N_2635,N_3752);
or U6110 (N_6110,N_4558,N_3449);
and U6111 (N_6111,N_3140,N_3359);
or U6112 (N_6112,N_2594,N_4397);
or U6113 (N_6113,N_3885,N_4511);
nand U6114 (N_6114,N_4059,N_3424);
xor U6115 (N_6115,N_4647,N_2597);
nand U6116 (N_6116,N_3336,N_3905);
and U6117 (N_6117,N_4931,N_4013);
nor U6118 (N_6118,N_3965,N_2525);
and U6119 (N_6119,N_3306,N_2643);
nand U6120 (N_6120,N_4699,N_4857);
nand U6121 (N_6121,N_3589,N_4337);
xnor U6122 (N_6122,N_2574,N_4939);
nor U6123 (N_6123,N_3618,N_3015);
or U6124 (N_6124,N_4612,N_4598);
nor U6125 (N_6125,N_4233,N_3246);
or U6126 (N_6126,N_4696,N_4517);
and U6127 (N_6127,N_4272,N_2733);
nand U6128 (N_6128,N_4192,N_3956);
nor U6129 (N_6129,N_4702,N_4537);
and U6130 (N_6130,N_3192,N_3453);
and U6131 (N_6131,N_4749,N_2627);
or U6132 (N_6132,N_3608,N_3326);
and U6133 (N_6133,N_3005,N_2788);
nor U6134 (N_6134,N_3209,N_2501);
or U6135 (N_6135,N_3836,N_4859);
xnor U6136 (N_6136,N_4374,N_4782);
nor U6137 (N_6137,N_3420,N_3023);
nand U6138 (N_6138,N_2598,N_4153);
nand U6139 (N_6139,N_2531,N_4354);
nor U6140 (N_6140,N_3430,N_4879);
xor U6141 (N_6141,N_3646,N_4396);
and U6142 (N_6142,N_3132,N_4206);
nor U6143 (N_6143,N_4934,N_4248);
xnor U6144 (N_6144,N_2641,N_3590);
nor U6145 (N_6145,N_3385,N_2749);
nand U6146 (N_6146,N_3444,N_3050);
or U6147 (N_6147,N_2576,N_4217);
nor U6148 (N_6148,N_2631,N_2644);
or U6149 (N_6149,N_3626,N_3870);
nand U6150 (N_6150,N_3225,N_3337);
nand U6151 (N_6151,N_4663,N_3913);
nor U6152 (N_6152,N_4423,N_2968);
and U6153 (N_6153,N_4786,N_4408);
or U6154 (N_6154,N_3211,N_3574);
and U6155 (N_6155,N_4332,N_3793);
or U6156 (N_6156,N_3753,N_3403);
nor U6157 (N_6157,N_3976,N_4486);
or U6158 (N_6158,N_3089,N_4404);
nand U6159 (N_6159,N_4169,N_2651);
and U6160 (N_6160,N_3967,N_4726);
nand U6161 (N_6161,N_2565,N_4418);
nor U6162 (N_6162,N_3741,N_3816);
and U6163 (N_6163,N_4411,N_2988);
nor U6164 (N_6164,N_2711,N_4720);
nor U6165 (N_6165,N_4783,N_2964);
or U6166 (N_6166,N_2615,N_2582);
nor U6167 (N_6167,N_2991,N_3890);
and U6168 (N_6168,N_4456,N_3393);
or U6169 (N_6169,N_3317,N_2960);
or U6170 (N_6170,N_3514,N_3594);
nor U6171 (N_6171,N_4560,N_2551);
and U6172 (N_6172,N_4010,N_4488);
nand U6173 (N_6173,N_2505,N_2882);
nor U6174 (N_6174,N_2851,N_3738);
and U6175 (N_6175,N_3489,N_4323);
nand U6176 (N_6176,N_3107,N_4230);
or U6177 (N_6177,N_2757,N_4072);
nand U6178 (N_6178,N_2541,N_3553);
nor U6179 (N_6179,N_4219,N_2634);
nand U6180 (N_6180,N_4636,N_3046);
and U6181 (N_6181,N_2681,N_4387);
nand U6182 (N_6182,N_4392,N_4188);
nor U6183 (N_6183,N_2740,N_4246);
nand U6184 (N_6184,N_3749,N_4561);
and U6185 (N_6185,N_4806,N_4886);
or U6186 (N_6186,N_3640,N_3596);
nand U6187 (N_6187,N_4603,N_2933);
and U6188 (N_6188,N_3071,N_4605);
nand U6189 (N_6189,N_3331,N_2787);
and U6190 (N_6190,N_3399,N_3288);
and U6191 (N_6191,N_4850,N_3593);
nor U6192 (N_6192,N_2729,N_4628);
or U6193 (N_6193,N_3387,N_3372);
nand U6194 (N_6194,N_3703,N_3352);
and U6195 (N_6195,N_4731,N_3242);
or U6196 (N_6196,N_2714,N_2738);
and U6197 (N_6197,N_3548,N_4874);
nor U6198 (N_6198,N_2797,N_4892);
or U6199 (N_6199,N_4798,N_4515);
and U6200 (N_6200,N_3022,N_4761);
or U6201 (N_6201,N_4695,N_3450);
or U6202 (N_6202,N_3671,N_3623);
nand U6203 (N_6203,N_2982,N_4860);
nor U6204 (N_6204,N_3397,N_4499);
xnor U6205 (N_6205,N_2728,N_3985);
and U6206 (N_6206,N_4220,N_3342);
or U6207 (N_6207,N_2756,N_3028);
nor U6208 (N_6208,N_3829,N_4676);
nor U6209 (N_6209,N_4556,N_3891);
or U6210 (N_6210,N_4735,N_4205);
nor U6211 (N_6211,N_3103,N_3332);
and U6212 (N_6212,N_3522,N_2764);
and U6213 (N_6213,N_2747,N_3157);
or U6214 (N_6214,N_2566,N_4733);
and U6215 (N_6215,N_4681,N_2618);
or U6216 (N_6216,N_4995,N_2861);
or U6217 (N_6217,N_3758,N_2953);
nor U6218 (N_6218,N_4303,N_3096);
xnor U6219 (N_6219,N_3353,N_4446);
or U6220 (N_6220,N_2859,N_4428);
nor U6221 (N_6221,N_3649,N_2774);
and U6222 (N_6222,N_4872,N_2692);
nand U6223 (N_6223,N_3360,N_3021);
nor U6224 (N_6224,N_2732,N_3505);
or U6225 (N_6225,N_4322,N_3201);
nand U6226 (N_6226,N_4607,N_4369);
or U6227 (N_6227,N_4395,N_4566);
nor U6228 (N_6228,N_3423,N_3455);
and U6229 (N_6229,N_4467,N_4329);
xnor U6230 (N_6230,N_4927,N_2916);
and U6231 (N_6231,N_3782,N_3414);
and U6232 (N_6232,N_3678,N_3338);
or U6233 (N_6233,N_4669,N_3493);
nand U6234 (N_6234,N_3483,N_3118);
nand U6235 (N_6235,N_3992,N_3879);
or U6236 (N_6236,N_2888,N_4661);
or U6237 (N_6237,N_3299,N_3685);
nor U6238 (N_6238,N_2544,N_2558);
or U6239 (N_6239,N_3815,N_4023);
nor U6240 (N_6240,N_4452,N_3715);
and U6241 (N_6241,N_3901,N_3515);
or U6242 (N_6242,N_3093,N_3149);
nand U6243 (N_6243,N_2556,N_4052);
and U6244 (N_6244,N_4564,N_4519);
nor U6245 (N_6245,N_4959,N_3289);
and U6246 (N_6246,N_4033,N_4756);
or U6247 (N_6247,N_2700,N_3436);
nor U6248 (N_6248,N_3587,N_4507);
xnor U6249 (N_6249,N_2951,N_4526);
and U6250 (N_6250,N_3269,N_4934);
nand U6251 (N_6251,N_4308,N_4730);
nor U6252 (N_6252,N_3752,N_2609);
or U6253 (N_6253,N_3520,N_3684);
nor U6254 (N_6254,N_3028,N_3021);
xnor U6255 (N_6255,N_4117,N_2708);
and U6256 (N_6256,N_4356,N_2762);
nand U6257 (N_6257,N_3077,N_2637);
or U6258 (N_6258,N_4070,N_4858);
xnor U6259 (N_6259,N_4940,N_3640);
nand U6260 (N_6260,N_4594,N_4563);
and U6261 (N_6261,N_4788,N_3062);
nor U6262 (N_6262,N_3933,N_3979);
xor U6263 (N_6263,N_2973,N_4140);
or U6264 (N_6264,N_3976,N_4104);
or U6265 (N_6265,N_4572,N_3471);
nand U6266 (N_6266,N_2583,N_3495);
and U6267 (N_6267,N_3610,N_3480);
nor U6268 (N_6268,N_2650,N_3286);
or U6269 (N_6269,N_3022,N_4073);
and U6270 (N_6270,N_4208,N_2960);
nand U6271 (N_6271,N_3006,N_2977);
and U6272 (N_6272,N_4615,N_2685);
nand U6273 (N_6273,N_3539,N_4857);
or U6274 (N_6274,N_4318,N_4449);
nor U6275 (N_6275,N_2884,N_3940);
nand U6276 (N_6276,N_3021,N_4837);
and U6277 (N_6277,N_4376,N_2914);
and U6278 (N_6278,N_4809,N_2999);
nor U6279 (N_6279,N_3710,N_4803);
or U6280 (N_6280,N_2570,N_4059);
and U6281 (N_6281,N_3079,N_4635);
or U6282 (N_6282,N_4957,N_4593);
nor U6283 (N_6283,N_2771,N_4455);
and U6284 (N_6284,N_2942,N_3428);
xor U6285 (N_6285,N_3115,N_4554);
nand U6286 (N_6286,N_4344,N_3841);
or U6287 (N_6287,N_3503,N_2537);
nor U6288 (N_6288,N_2559,N_4211);
and U6289 (N_6289,N_3826,N_3960);
nand U6290 (N_6290,N_3461,N_4274);
nand U6291 (N_6291,N_3844,N_4485);
or U6292 (N_6292,N_3739,N_2694);
or U6293 (N_6293,N_4790,N_4464);
and U6294 (N_6294,N_3384,N_2553);
xnor U6295 (N_6295,N_2546,N_2655);
or U6296 (N_6296,N_3403,N_4852);
xor U6297 (N_6297,N_3974,N_4641);
nor U6298 (N_6298,N_3443,N_2598);
and U6299 (N_6299,N_4680,N_3355);
nand U6300 (N_6300,N_4407,N_3715);
and U6301 (N_6301,N_4344,N_3017);
or U6302 (N_6302,N_2622,N_2525);
nand U6303 (N_6303,N_4284,N_3050);
nor U6304 (N_6304,N_4015,N_4472);
xnor U6305 (N_6305,N_4941,N_4437);
xnor U6306 (N_6306,N_3738,N_3964);
and U6307 (N_6307,N_4903,N_4548);
or U6308 (N_6308,N_3263,N_3086);
nor U6309 (N_6309,N_3712,N_3832);
and U6310 (N_6310,N_4546,N_4926);
or U6311 (N_6311,N_4799,N_3561);
and U6312 (N_6312,N_4522,N_3002);
nor U6313 (N_6313,N_4145,N_3747);
and U6314 (N_6314,N_3411,N_4876);
nand U6315 (N_6315,N_4599,N_2695);
and U6316 (N_6316,N_3046,N_2994);
xnor U6317 (N_6317,N_4732,N_4722);
nand U6318 (N_6318,N_3765,N_2877);
or U6319 (N_6319,N_3176,N_3850);
nor U6320 (N_6320,N_4171,N_3529);
nor U6321 (N_6321,N_2511,N_3525);
and U6322 (N_6322,N_4545,N_4007);
nand U6323 (N_6323,N_4271,N_3439);
or U6324 (N_6324,N_4035,N_3807);
nor U6325 (N_6325,N_4563,N_4934);
and U6326 (N_6326,N_4503,N_2963);
nor U6327 (N_6327,N_4032,N_4425);
nand U6328 (N_6328,N_4003,N_3566);
nor U6329 (N_6329,N_4896,N_3543);
and U6330 (N_6330,N_3773,N_4455);
nand U6331 (N_6331,N_4771,N_3097);
nand U6332 (N_6332,N_3460,N_2685);
nand U6333 (N_6333,N_3567,N_3458);
xor U6334 (N_6334,N_2554,N_2533);
nor U6335 (N_6335,N_4397,N_3453);
or U6336 (N_6336,N_3064,N_2541);
and U6337 (N_6337,N_2955,N_3897);
nor U6338 (N_6338,N_3111,N_3817);
and U6339 (N_6339,N_2523,N_4939);
and U6340 (N_6340,N_3226,N_3686);
or U6341 (N_6341,N_3923,N_4660);
and U6342 (N_6342,N_4315,N_3659);
nand U6343 (N_6343,N_2871,N_4066);
and U6344 (N_6344,N_4944,N_2879);
nand U6345 (N_6345,N_2794,N_4721);
nand U6346 (N_6346,N_3821,N_4117);
nor U6347 (N_6347,N_3965,N_3924);
or U6348 (N_6348,N_4194,N_4477);
or U6349 (N_6349,N_3815,N_2640);
nor U6350 (N_6350,N_3324,N_4567);
or U6351 (N_6351,N_4798,N_4642);
nor U6352 (N_6352,N_2564,N_4148);
nor U6353 (N_6353,N_2641,N_4346);
and U6354 (N_6354,N_4022,N_4446);
and U6355 (N_6355,N_3238,N_4321);
and U6356 (N_6356,N_4899,N_3544);
xor U6357 (N_6357,N_3709,N_4130);
xor U6358 (N_6358,N_4623,N_3647);
and U6359 (N_6359,N_4795,N_4676);
xor U6360 (N_6360,N_4838,N_3920);
and U6361 (N_6361,N_4922,N_3741);
or U6362 (N_6362,N_4174,N_3224);
or U6363 (N_6363,N_3927,N_4401);
nor U6364 (N_6364,N_3874,N_3031);
nand U6365 (N_6365,N_4391,N_2545);
or U6366 (N_6366,N_4731,N_4765);
nand U6367 (N_6367,N_4594,N_3692);
nor U6368 (N_6368,N_3185,N_2747);
nand U6369 (N_6369,N_4531,N_4106);
or U6370 (N_6370,N_4149,N_3459);
and U6371 (N_6371,N_3550,N_4428);
and U6372 (N_6372,N_2808,N_3464);
nand U6373 (N_6373,N_3455,N_2767);
or U6374 (N_6374,N_3019,N_3819);
nand U6375 (N_6375,N_3806,N_4462);
or U6376 (N_6376,N_3207,N_4402);
nand U6377 (N_6377,N_4062,N_3905);
and U6378 (N_6378,N_3418,N_3792);
nand U6379 (N_6379,N_4093,N_3774);
nor U6380 (N_6380,N_4537,N_4962);
nor U6381 (N_6381,N_3373,N_4367);
nor U6382 (N_6382,N_4744,N_2815);
and U6383 (N_6383,N_2720,N_4737);
or U6384 (N_6384,N_3770,N_4224);
nor U6385 (N_6385,N_3016,N_3609);
and U6386 (N_6386,N_3112,N_4127);
xnor U6387 (N_6387,N_3661,N_3612);
or U6388 (N_6388,N_3636,N_2865);
nor U6389 (N_6389,N_3628,N_4704);
and U6390 (N_6390,N_3479,N_4559);
or U6391 (N_6391,N_2551,N_3773);
xor U6392 (N_6392,N_4637,N_3792);
or U6393 (N_6393,N_4929,N_4225);
and U6394 (N_6394,N_2870,N_4248);
nor U6395 (N_6395,N_3142,N_2725);
or U6396 (N_6396,N_4831,N_3454);
xor U6397 (N_6397,N_2987,N_2769);
and U6398 (N_6398,N_3348,N_4006);
nand U6399 (N_6399,N_3803,N_3382);
nand U6400 (N_6400,N_4327,N_4781);
or U6401 (N_6401,N_3090,N_3897);
and U6402 (N_6402,N_3798,N_3394);
xnor U6403 (N_6403,N_3266,N_3502);
and U6404 (N_6404,N_3004,N_4139);
or U6405 (N_6405,N_3779,N_2513);
or U6406 (N_6406,N_3861,N_4506);
nand U6407 (N_6407,N_3193,N_2631);
or U6408 (N_6408,N_2873,N_2946);
nand U6409 (N_6409,N_2511,N_4631);
nand U6410 (N_6410,N_4348,N_4101);
nor U6411 (N_6411,N_4421,N_4933);
or U6412 (N_6412,N_3713,N_3818);
nor U6413 (N_6413,N_3057,N_4880);
or U6414 (N_6414,N_4024,N_3303);
nor U6415 (N_6415,N_2731,N_4543);
nand U6416 (N_6416,N_3654,N_3303);
nor U6417 (N_6417,N_4130,N_4922);
or U6418 (N_6418,N_3207,N_4376);
or U6419 (N_6419,N_3410,N_4149);
xnor U6420 (N_6420,N_2840,N_3812);
or U6421 (N_6421,N_3518,N_3933);
nor U6422 (N_6422,N_3649,N_3413);
and U6423 (N_6423,N_4233,N_3954);
and U6424 (N_6424,N_3477,N_3525);
and U6425 (N_6425,N_2939,N_4211);
nand U6426 (N_6426,N_4935,N_2550);
nor U6427 (N_6427,N_4150,N_2606);
and U6428 (N_6428,N_2520,N_2999);
nor U6429 (N_6429,N_2958,N_4135);
nor U6430 (N_6430,N_4562,N_3123);
or U6431 (N_6431,N_4881,N_3998);
and U6432 (N_6432,N_3873,N_4958);
and U6433 (N_6433,N_3905,N_4649);
and U6434 (N_6434,N_2707,N_3426);
or U6435 (N_6435,N_3967,N_4240);
and U6436 (N_6436,N_3921,N_4864);
or U6437 (N_6437,N_3166,N_4206);
xor U6438 (N_6438,N_2717,N_3942);
or U6439 (N_6439,N_3465,N_4169);
nor U6440 (N_6440,N_4050,N_4215);
or U6441 (N_6441,N_4604,N_4548);
xor U6442 (N_6442,N_4314,N_3310);
and U6443 (N_6443,N_4397,N_4970);
nand U6444 (N_6444,N_3188,N_4495);
and U6445 (N_6445,N_4691,N_3931);
xor U6446 (N_6446,N_2592,N_4113);
nand U6447 (N_6447,N_3149,N_3378);
or U6448 (N_6448,N_4591,N_3154);
nor U6449 (N_6449,N_2906,N_3637);
and U6450 (N_6450,N_4116,N_3855);
nor U6451 (N_6451,N_3031,N_3750);
or U6452 (N_6452,N_3061,N_4327);
xor U6453 (N_6453,N_2717,N_3744);
or U6454 (N_6454,N_4214,N_4069);
and U6455 (N_6455,N_4600,N_2795);
nor U6456 (N_6456,N_4801,N_4787);
xor U6457 (N_6457,N_4488,N_3735);
nor U6458 (N_6458,N_4840,N_3130);
xnor U6459 (N_6459,N_3101,N_3477);
nor U6460 (N_6460,N_2649,N_2838);
nor U6461 (N_6461,N_3550,N_3585);
nand U6462 (N_6462,N_3438,N_3743);
and U6463 (N_6463,N_3115,N_2760);
nor U6464 (N_6464,N_4011,N_4568);
nand U6465 (N_6465,N_2735,N_3909);
xnor U6466 (N_6466,N_3662,N_3337);
nor U6467 (N_6467,N_4816,N_3277);
nor U6468 (N_6468,N_4330,N_4038);
or U6469 (N_6469,N_3708,N_4120);
nor U6470 (N_6470,N_4982,N_4434);
nand U6471 (N_6471,N_3839,N_2983);
xnor U6472 (N_6472,N_3638,N_2825);
and U6473 (N_6473,N_4044,N_3754);
nor U6474 (N_6474,N_4232,N_3511);
nand U6475 (N_6475,N_4758,N_4522);
and U6476 (N_6476,N_2807,N_3485);
xor U6477 (N_6477,N_4761,N_4069);
nand U6478 (N_6478,N_3335,N_3994);
nor U6479 (N_6479,N_3509,N_3676);
and U6480 (N_6480,N_4724,N_3697);
and U6481 (N_6481,N_3562,N_4450);
and U6482 (N_6482,N_3124,N_2506);
nor U6483 (N_6483,N_3631,N_4498);
xnor U6484 (N_6484,N_4368,N_2654);
nor U6485 (N_6485,N_2568,N_4958);
nor U6486 (N_6486,N_4008,N_4974);
nor U6487 (N_6487,N_3962,N_3951);
nand U6488 (N_6488,N_3134,N_3777);
and U6489 (N_6489,N_3881,N_3312);
and U6490 (N_6490,N_2706,N_2662);
nand U6491 (N_6491,N_4105,N_3906);
nor U6492 (N_6492,N_3497,N_4031);
or U6493 (N_6493,N_3050,N_3520);
or U6494 (N_6494,N_4879,N_3603);
nor U6495 (N_6495,N_3965,N_2997);
and U6496 (N_6496,N_3627,N_3933);
xnor U6497 (N_6497,N_4747,N_3379);
or U6498 (N_6498,N_4726,N_4236);
xnor U6499 (N_6499,N_4024,N_4323);
and U6500 (N_6500,N_2640,N_4685);
and U6501 (N_6501,N_3624,N_2623);
nand U6502 (N_6502,N_2963,N_2827);
or U6503 (N_6503,N_3258,N_2659);
and U6504 (N_6504,N_3439,N_3757);
or U6505 (N_6505,N_3825,N_4247);
and U6506 (N_6506,N_3120,N_4935);
nor U6507 (N_6507,N_2628,N_3509);
nand U6508 (N_6508,N_3555,N_4044);
or U6509 (N_6509,N_3704,N_4739);
nand U6510 (N_6510,N_3642,N_2986);
nand U6511 (N_6511,N_2650,N_4648);
nor U6512 (N_6512,N_3660,N_4035);
xnor U6513 (N_6513,N_2978,N_4325);
nand U6514 (N_6514,N_3186,N_3957);
or U6515 (N_6515,N_2624,N_4591);
xor U6516 (N_6516,N_4655,N_4043);
and U6517 (N_6517,N_2771,N_3527);
and U6518 (N_6518,N_4815,N_4951);
nand U6519 (N_6519,N_3834,N_3125);
and U6520 (N_6520,N_4851,N_2689);
nand U6521 (N_6521,N_4597,N_4234);
nor U6522 (N_6522,N_3735,N_3151);
and U6523 (N_6523,N_3634,N_4010);
nand U6524 (N_6524,N_2960,N_3855);
or U6525 (N_6525,N_3492,N_2880);
nand U6526 (N_6526,N_4209,N_4497);
or U6527 (N_6527,N_2843,N_2783);
nand U6528 (N_6528,N_3962,N_3695);
nand U6529 (N_6529,N_4716,N_4728);
or U6530 (N_6530,N_4207,N_3361);
or U6531 (N_6531,N_2879,N_4817);
or U6532 (N_6532,N_3014,N_4046);
or U6533 (N_6533,N_3183,N_4043);
nor U6534 (N_6534,N_3769,N_2733);
and U6535 (N_6535,N_3525,N_4344);
nor U6536 (N_6536,N_4516,N_2643);
xor U6537 (N_6537,N_3385,N_3084);
or U6538 (N_6538,N_3361,N_4540);
and U6539 (N_6539,N_4156,N_4158);
nand U6540 (N_6540,N_3405,N_3337);
nor U6541 (N_6541,N_4234,N_3834);
nor U6542 (N_6542,N_4961,N_3448);
and U6543 (N_6543,N_2721,N_4679);
nor U6544 (N_6544,N_4537,N_2970);
and U6545 (N_6545,N_3973,N_2805);
nor U6546 (N_6546,N_3546,N_4503);
xor U6547 (N_6547,N_2607,N_4813);
nor U6548 (N_6548,N_4408,N_4756);
nand U6549 (N_6549,N_4270,N_2657);
xnor U6550 (N_6550,N_3488,N_4925);
nand U6551 (N_6551,N_4687,N_4412);
or U6552 (N_6552,N_4723,N_4256);
nor U6553 (N_6553,N_3254,N_4820);
nand U6554 (N_6554,N_3836,N_3674);
and U6555 (N_6555,N_3864,N_4905);
nor U6556 (N_6556,N_2902,N_4836);
and U6557 (N_6557,N_3756,N_4308);
and U6558 (N_6558,N_4137,N_2639);
nand U6559 (N_6559,N_3422,N_2725);
and U6560 (N_6560,N_4476,N_4638);
or U6561 (N_6561,N_3473,N_4968);
and U6562 (N_6562,N_4996,N_2694);
nand U6563 (N_6563,N_2751,N_4182);
and U6564 (N_6564,N_3650,N_4384);
nor U6565 (N_6565,N_2698,N_4254);
nor U6566 (N_6566,N_3333,N_3886);
and U6567 (N_6567,N_2806,N_4276);
or U6568 (N_6568,N_3164,N_4134);
nand U6569 (N_6569,N_3323,N_4226);
and U6570 (N_6570,N_3287,N_2608);
and U6571 (N_6571,N_4764,N_4033);
nor U6572 (N_6572,N_3826,N_3828);
nor U6573 (N_6573,N_4282,N_3376);
or U6574 (N_6574,N_3400,N_2663);
or U6575 (N_6575,N_3917,N_4820);
nand U6576 (N_6576,N_4155,N_3236);
and U6577 (N_6577,N_4078,N_3167);
or U6578 (N_6578,N_2528,N_4315);
or U6579 (N_6579,N_4614,N_4628);
nand U6580 (N_6580,N_4402,N_3708);
and U6581 (N_6581,N_3434,N_3054);
nor U6582 (N_6582,N_4106,N_3023);
nor U6583 (N_6583,N_3354,N_3078);
or U6584 (N_6584,N_3464,N_2842);
nor U6585 (N_6585,N_3242,N_3911);
nand U6586 (N_6586,N_2767,N_2859);
and U6587 (N_6587,N_2665,N_4434);
nor U6588 (N_6588,N_4296,N_4546);
and U6589 (N_6589,N_3475,N_2723);
or U6590 (N_6590,N_3241,N_4375);
or U6591 (N_6591,N_4232,N_3509);
nor U6592 (N_6592,N_4773,N_4752);
or U6593 (N_6593,N_4317,N_3700);
or U6594 (N_6594,N_3512,N_4905);
or U6595 (N_6595,N_3373,N_2861);
and U6596 (N_6596,N_2507,N_3575);
nand U6597 (N_6597,N_3884,N_4810);
nor U6598 (N_6598,N_2594,N_2747);
nand U6599 (N_6599,N_4766,N_3242);
nand U6600 (N_6600,N_4279,N_4943);
nand U6601 (N_6601,N_4782,N_4144);
nand U6602 (N_6602,N_3516,N_3160);
and U6603 (N_6603,N_4652,N_3612);
or U6604 (N_6604,N_2525,N_4061);
or U6605 (N_6605,N_3284,N_3605);
and U6606 (N_6606,N_3659,N_3195);
nor U6607 (N_6607,N_2970,N_3764);
nand U6608 (N_6608,N_3423,N_3749);
and U6609 (N_6609,N_2605,N_3243);
nor U6610 (N_6610,N_2666,N_3328);
nor U6611 (N_6611,N_2605,N_3918);
and U6612 (N_6612,N_3604,N_3535);
or U6613 (N_6613,N_4926,N_3293);
or U6614 (N_6614,N_4330,N_3907);
nor U6615 (N_6615,N_3154,N_3817);
or U6616 (N_6616,N_4181,N_2909);
and U6617 (N_6617,N_3008,N_3612);
nor U6618 (N_6618,N_3128,N_4018);
and U6619 (N_6619,N_4167,N_3314);
nand U6620 (N_6620,N_4458,N_2501);
nand U6621 (N_6621,N_2907,N_4583);
or U6622 (N_6622,N_4057,N_2767);
xor U6623 (N_6623,N_3373,N_3457);
nor U6624 (N_6624,N_2791,N_3112);
or U6625 (N_6625,N_3323,N_4165);
nor U6626 (N_6626,N_3338,N_2512);
nor U6627 (N_6627,N_3190,N_3179);
or U6628 (N_6628,N_2669,N_4381);
or U6629 (N_6629,N_4834,N_3938);
or U6630 (N_6630,N_2995,N_4140);
nand U6631 (N_6631,N_3488,N_2798);
or U6632 (N_6632,N_3322,N_2745);
and U6633 (N_6633,N_4631,N_3064);
nand U6634 (N_6634,N_4542,N_4740);
or U6635 (N_6635,N_3176,N_3864);
nor U6636 (N_6636,N_4384,N_3736);
nor U6637 (N_6637,N_2936,N_2783);
nor U6638 (N_6638,N_3868,N_2599);
and U6639 (N_6639,N_4533,N_4308);
or U6640 (N_6640,N_2539,N_3155);
nand U6641 (N_6641,N_3268,N_4980);
or U6642 (N_6642,N_4469,N_3320);
nand U6643 (N_6643,N_4798,N_4887);
and U6644 (N_6644,N_4175,N_3516);
and U6645 (N_6645,N_2699,N_2672);
and U6646 (N_6646,N_2724,N_2616);
and U6647 (N_6647,N_3649,N_3801);
nand U6648 (N_6648,N_3624,N_4153);
or U6649 (N_6649,N_4699,N_3674);
nor U6650 (N_6650,N_4796,N_3201);
nand U6651 (N_6651,N_4386,N_4912);
and U6652 (N_6652,N_4880,N_4752);
nor U6653 (N_6653,N_3749,N_2766);
xnor U6654 (N_6654,N_4863,N_2998);
or U6655 (N_6655,N_3745,N_4777);
and U6656 (N_6656,N_2545,N_3804);
or U6657 (N_6657,N_4937,N_2749);
and U6658 (N_6658,N_4619,N_4020);
xnor U6659 (N_6659,N_2531,N_4823);
nand U6660 (N_6660,N_3006,N_4929);
or U6661 (N_6661,N_2921,N_4493);
and U6662 (N_6662,N_3632,N_2753);
and U6663 (N_6663,N_3590,N_3351);
nor U6664 (N_6664,N_4708,N_3205);
nor U6665 (N_6665,N_4445,N_2884);
or U6666 (N_6666,N_3884,N_3474);
nor U6667 (N_6667,N_3355,N_3170);
nor U6668 (N_6668,N_3727,N_2592);
and U6669 (N_6669,N_4562,N_4028);
xnor U6670 (N_6670,N_3957,N_2589);
and U6671 (N_6671,N_3431,N_3599);
or U6672 (N_6672,N_3514,N_3717);
xor U6673 (N_6673,N_3248,N_2763);
and U6674 (N_6674,N_3349,N_3180);
or U6675 (N_6675,N_4898,N_4269);
and U6676 (N_6676,N_4477,N_2912);
or U6677 (N_6677,N_4527,N_2829);
xor U6678 (N_6678,N_2856,N_4352);
and U6679 (N_6679,N_3709,N_4634);
or U6680 (N_6680,N_3084,N_3327);
and U6681 (N_6681,N_4838,N_3602);
or U6682 (N_6682,N_3639,N_4675);
nand U6683 (N_6683,N_4916,N_4155);
and U6684 (N_6684,N_4974,N_4668);
xor U6685 (N_6685,N_3906,N_3827);
xnor U6686 (N_6686,N_4768,N_3597);
or U6687 (N_6687,N_3163,N_4124);
and U6688 (N_6688,N_4786,N_3348);
or U6689 (N_6689,N_4334,N_3326);
xor U6690 (N_6690,N_4934,N_4385);
nand U6691 (N_6691,N_4995,N_4642);
nor U6692 (N_6692,N_4598,N_3263);
and U6693 (N_6693,N_3466,N_4657);
and U6694 (N_6694,N_2609,N_3260);
nor U6695 (N_6695,N_3879,N_3438);
or U6696 (N_6696,N_4908,N_3892);
and U6697 (N_6697,N_4694,N_4980);
and U6698 (N_6698,N_2866,N_4351);
and U6699 (N_6699,N_3847,N_4226);
xnor U6700 (N_6700,N_3449,N_4241);
and U6701 (N_6701,N_2994,N_4714);
or U6702 (N_6702,N_3662,N_3565);
or U6703 (N_6703,N_3502,N_3664);
and U6704 (N_6704,N_2645,N_4523);
or U6705 (N_6705,N_3700,N_3712);
nand U6706 (N_6706,N_4513,N_4997);
and U6707 (N_6707,N_3901,N_2933);
or U6708 (N_6708,N_2577,N_4688);
xor U6709 (N_6709,N_3209,N_3702);
nand U6710 (N_6710,N_3351,N_4083);
nor U6711 (N_6711,N_3006,N_3296);
xnor U6712 (N_6712,N_2510,N_4787);
nand U6713 (N_6713,N_3236,N_4174);
and U6714 (N_6714,N_4363,N_3832);
nor U6715 (N_6715,N_3461,N_2975);
or U6716 (N_6716,N_3018,N_4440);
xor U6717 (N_6717,N_3650,N_3742);
or U6718 (N_6718,N_3223,N_3080);
xor U6719 (N_6719,N_4709,N_4638);
or U6720 (N_6720,N_2571,N_4334);
or U6721 (N_6721,N_2639,N_2993);
and U6722 (N_6722,N_4589,N_4650);
and U6723 (N_6723,N_4470,N_4162);
nand U6724 (N_6724,N_2623,N_2862);
nor U6725 (N_6725,N_3211,N_2772);
and U6726 (N_6726,N_3710,N_3192);
or U6727 (N_6727,N_4704,N_4473);
nand U6728 (N_6728,N_3801,N_4026);
nor U6729 (N_6729,N_4815,N_4088);
nor U6730 (N_6730,N_4751,N_3226);
or U6731 (N_6731,N_4357,N_4445);
nand U6732 (N_6732,N_3475,N_2546);
xor U6733 (N_6733,N_2918,N_3189);
nand U6734 (N_6734,N_3227,N_4185);
nand U6735 (N_6735,N_4326,N_3501);
xor U6736 (N_6736,N_4932,N_3848);
or U6737 (N_6737,N_4228,N_3512);
and U6738 (N_6738,N_3694,N_2787);
nor U6739 (N_6739,N_3823,N_4153);
nor U6740 (N_6740,N_4133,N_2986);
or U6741 (N_6741,N_4600,N_4706);
nor U6742 (N_6742,N_4028,N_4623);
and U6743 (N_6743,N_4944,N_3787);
nand U6744 (N_6744,N_3585,N_3208);
nand U6745 (N_6745,N_2903,N_3203);
or U6746 (N_6746,N_4628,N_3400);
xnor U6747 (N_6747,N_4289,N_2590);
and U6748 (N_6748,N_3634,N_3928);
xnor U6749 (N_6749,N_3242,N_3531);
nand U6750 (N_6750,N_4826,N_3876);
and U6751 (N_6751,N_4284,N_4079);
nor U6752 (N_6752,N_4345,N_2774);
or U6753 (N_6753,N_4274,N_3596);
nor U6754 (N_6754,N_4484,N_2756);
and U6755 (N_6755,N_4622,N_3160);
nand U6756 (N_6756,N_2832,N_3857);
nand U6757 (N_6757,N_3567,N_2643);
nor U6758 (N_6758,N_2894,N_3648);
or U6759 (N_6759,N_4771,N_3061);
xnor U6760 (N_6760,N_3311,N_4196);
nand U6761 (N_6761,N_3176,N_3277);
and U6762 (N_6762,N_2828,N_2628);
or U6763 (N_6763,N_4891,N_3594);
and U6764 (N_6764,N_3205,N_4222);
or U6765 (N_6765,N_2587,N_2922);
and U6766 (N_6766,N_4173,N_4013);
or U6767 (N_6767,N_3909,N_3543);
or U6768 (N_6768,N_2502,N_4501);
nand U6769 (N_6769,N_4053,N_3573);
xor U6770 (N_6770,N_4687,N_4423);
and U6771 (N_6771,N_4903,N_3438);
xor U6772 (N_6772,N_3853,N_3146);
and U6773 (N_6773,N_3667,N_3513);
and U6774 (N_6774,N_2997,N_3033);
nand U6775 (N_6775,N_4878,N_4630);
and U6776 (N_6776,N_3654,N_4129);
or U6777 (N_6777,N_4063,N_3537);
and U6778 (N_6778,N_4716,N_3322);
and U6779 (N_6779,N_2839,N_2534);
or U6780 (N_6780,N_3744,N_4958);
xor U6781 (N_6781,N_3044,N_4007);
or U6782 (N_6782,N_2734,N_2766);
and U6783 (N_6783,N_3750,N_4341);
and U6784 (N_6784,N_3871,N_3597);
nor U6785 (N_6785,N_3799,N_3485);
nand U6786 (N_6786,N_4260,N_4426);
nand U6787 (N_6787,N_4294,N_3470);
or U6788 (N_6788,N_3955,N_4474);
nor U6789 (N_6789,N_3636,N_4686);
nor U6790 (N_6790,N_3640,N_4720);
xnor U6791 (N_6791,N_3936,N_3369);
and U6792 (N_6792,N_4584,N_3856);
nand U6793 (N_6793,N_4425,N_3954);
nor U6794 (N_6794,N_3776,N_3449);
and U6795 (N_6795,N_2623,N_3906);
nand U6796 (N_6796,N_3043,N_3632);
nand U6797 (N_6797,N_4290,N_4284);
nor U6798 (N_6798,N_2660,N_3905);
or U6799 (N_6799,N_4349,N_3478);
xnor U6800 (N_6800,N_4941,N_3078);
or U6801 (N_6801,N_3637,N_4910);
nand U6802 (N_6802,N_2961,N_4361);
and U6803 (N_6803,N_3848,N_4783);
and U6804 (N_6804,N_4848,N_4801);
or U6805 (N_6805,N_4650,N_2985);
nor U6806 (N_6806,N_3672,N_3053);
xor U6807 (N_6807,N_2554,N_3893);
xnor U6808 (N_6808,N_3826,N_3293);
nor U6809 (N_6809,N_3619,N_4379);
nand U6810 (N_6810,N_3218,N_3714);
or U6811 (N_6811,N_4548,N_4592);
or U6812 (N_6812,N_3746,N_3700);
nand U6813 (N_6813,N_3613,N_4872);
nand U6814 (N_6814,N_3858,N_3223);
nor U6815 (N_6815,N_4596,N_4764);
and U6816 (N_6816,N_2873,N_3094);
nor U6817 (N_6817,N_2851,N_3314);
nand U6818 (N_6818,N_4513,N_4479);
nand U6819 (N_6819,N_3635,N_4048);
and U6820 (N_6820,N_4109,N_2722);
nand U6821 (N_6821,N_3338,N_3293);
xor U6822 (N_6822,N_3453,N_3436);
or U6823 (N_6823,N_4785,N_3273);
nand U6824 (N_6824,N_4533,N_3811);
nand U6825 (N_6825,N_2907,N_3529);
or U6826 (N_6826,N_3743,N_3708);
or U6827 (N_6827,N_3522,N_4491);
nor U6828 (N_6828,N_3774,N_3478);
nor U6829 (N_6829,N_3473,N_4685);
or U6830 (N_6830,N_3349,N_3405);
nand U6831 (N_6831,N_2586,N_3636);
and U6832 (N_6832,N_4931,N_3392);
nand U6833 (N_6833,N_4997,N_4814);
and U6834 (N_6834,N_4138,N_3973);
nor U6835 (N_6835,N_3298,N_2766);
or U6836 (N_6836,N_4076,N_3352);
or U6837 (N_6837,N_4029,N_4659);
and U6838 (N_6838,N_4918,N_3540);
and U6839 (N_6839,N_3933,N_3014);
and U6840 (N_6840,N_4717,N_2940);
xnor U6841 (N_6841,N_3078,N_2843);
xnor U6842 (N_6842,N_3336,N_3665);
nand U6843 (N_6843,N_2724,N_4887);
nand U6844 (N_6844,N_4709,N_3073);
nor U6845 (N_6845,N_4707,N_4159);
and U6846 (N_6846,N_3389,N_4686);
nor U6847 (N_6847,N_2818,N_2566);
nand U6848 (N_6848,N_4942,N_3189);
xnor U6849 (N_6849,N_4922,N_3953);
and U6850 (N_6850,N_4585,N_4449);
or U6851 (N_6851,N_3284,N_3436);
nand U6852 (N_6852,N_2887,N_4388);
and U6853 (N_6853,N_2504,N_3132);
nor U6854 (N_6854,N_3542,N_2923);
xnor U6855 (N_6855,N_4670,N_4140);
and U6856 (N_6856,N_3436,N_4731);
or U6857 (N_6857,N_3958,N_2788);
nand U6858 (N_6858,N_4283,N_3998);
or U6859 (N_6859,N_2506,N_3429);
and U6860 (N_6860,N_2638,N_2746);
xor U6861 (N_6861,N_3688,N_2926);
or U6862 (N_6862,N_4440,N_4356);
or U6863 (N_6863,N_3269,N_4553);
nand U6864 (N_6864,N_4086,N_3477);
xor U6865 (N_6865,N_4043,N_4695);
xnor U6866 (N_6866,N_3123,N_4191);
nor U6867 (N_6867,N_3752,N_4653);
or U6868 (N_6868,N_2536,N_3034);
and U6869 (N_6869,N_3325,N_3280);
nand U6870 (N_6870,N_4274,N_4808);
or U6871 (N_6871,N_3078,N_2675);
nor U6872 (N_6872,N_4980,N_3585);
nor U6873 (N_6873,N_4472,N_3866);
xnor U6874 (N_6874,N_4967,N_3741);
nor U6875 (N_6875,N_3228,N_4783);
or U6876 (N_6876,N_2946,N_3657);
and U6877 (N_6877,N_3745,N_4549);
and U6878 (N_6878,N_3766,N_2542);
nand U6879 (N_6879,N_4599,N_4495);
or U6880 (N_6880,N_3249,N_4960);
and U6881 (N_6881,N_4511,N_3597);
or U6882 (N_6882,N_4286,N_2563);
xor U6883 (N_6883,N_4657,N_4941);
nor U6884 (N_6884,N_3270,N_2681);
nor U6885 (N_6885,N_4047,N_4486);
nand U6886 (N_6886,N_3417,N_3257);
or U6887 (N_6887,N_4471,N_3407);
and U6888 (N_6888,N_3274,N_2771);
nor U6889 (N_6889,N_2665,N_3403);
and U6890 (N_6890,N_3690,N_3573);
nand U6891 (N_6891,N_3628,N_4762);
nor U6892 (N_6892,N_4060,N_2995);
or U6893 (N_6893,N_4449,N_2617);
xnor U6894 (N_6894,N_2828,N_4239);
or U6895 (N_6895,N_3485,N_3842);
nand U6896 (N_6896,N_4512,N_3555);
nor U6897 (N_6897,N_4539,N_3960);
nor U6898 (N_6898,N_3161,N_4197);
or U6899 (N_6899,N_2939,N_3199);
nand U6900 (N_6900,N_4547,N_3865);
and U6901 (N_6901,N_4473,N_3430);
nand U6902 (N_6902,N_4896,N_4878);
nor U6903 (N_6903,N_4051,N_3412);
nor U6904 (N_6904,N_4735,N_2547);
and U6905 (N_6905,N_3605,N_2616);
nand U6906 (N_6906,N_2850,N_4056);
xor U6907 (N_6907,N_4999,N_3397);
nor U6908 (N_6908,N_4913,N_4211);
nand U6909 (N_6909,N_4722,N_3954);
nor U6910 (N_6910,N_2740,N_3655);
and U6911 (N_6911,N_4321,N_3757);
xor U6912 (N_6912,N_4424,N_2932);
or U6913 (N_6913,N_2899,N_3052);
nand U6914 (N_6914,N_4976,N_3523);
or U6915 (N_6915,N_3424,N_3449);
or U6916 (N_6916,N_3866,N_2545);
or U6917 (N_6917,N_2651,N_2592);
and U6918 (N_6918,N_4130,N_4366);
or U6919 (N_6919,N_4065,N_3710);
nor U6920 (N_6920,N_3604,N_3858);
nor U6921 (N_6921,N_3545,N_4050);
or U6922 (N_6922,N_2756,N_3987);
nor U6923 (N_6923,N_2962,N_3582);
or U6924 (N_6924,N_4825,N_4225);
nor U6925 (N_6925,N_4796,N_4999);
or U6926 (N_6926,N_4650,N_4477);
or U6927 (N_6927,N_2634,N_4104);
or U6928 (N_6928,N_4082,N_4445);
and U6929 (N_6929,N_3456,N_3305);
nand U6930 (N_6930,N_2778,N_3841);
nor U6931 (N_6931,N_4103,N_2608);
and U6932 (N_6932,N_4752,N_4810);
nand U6933 (N_6933,N_4712,N_4160);
nor U6934 (N_6934,N_2542,N_3097);
nand U6935 (N_6935,N_4775,N_4807);
or U6936 (N_6936,N_4953,N_2655);
and U6937 (N_6937,N_2652,N_3890);
and U6938 (N_6938,N_4833,N_4983);
nor U6939 (N_6939,N_4830,N_4665);
nor U6940 (N_6940,N_3097,N_4331);
nand U6941 (N_6941,N_4701,N_3617);
nand U6942 (N_6942,N_3899,N_3387);
nor U6943 (N_6943,N_2780,N_4879);
or U6944 (N_6944,N_3467,N_3704);
and U6945 (N_6945,N_4341,N_3341);
nor U6946 (N_6946,N_4842,N_4986);
and U6947 (N_6947,N_3459,N_4933);
or U6948 (N_6948,N_2501,N_4948);
nand U6949 (N_6949,N_2869,N_3545);
and U6950 (N_6950,N_3941,N_3897);
and U6951 (N_6951,N_2766,N_3729);
or U6952 (N_6952,N_2630,N_4057);
or U6953 (N_6953,N_3817,N_3652);
or U6954 (N_6954,N_4587,N_3680);
or U6955 (N_6955,N_2535,N_4724);
and U6956 (N_6956,N_4437,N_4444);
or U6957 (N_6957,N_4166,N_3337);
xnor U6958 (N_6958,N_4563,N_3487);
nor U6959 (N_6959,N_4260,N_2696);
xor U6960 (N_6960,N_3388,N_4977);
nand U6961 (N_6961,N_3460,N_3077);
nand U6962 (N_6962,N_3394,N_3368);
nand U6963 (N_6963,N_2513,N_4069);
and U6964 (N_6964,N_3929,N_4954);
or U6965 (N_6965,N_3674,N_4165);
and U6966 (N_6966,N_2642,N_4895);
and U6967 (N_6967,N_2630,N_3541);
and U6968 (N_6968,N_4397,N_4141);
or U6969 (N_6969,N_4843,N_2673);
and U6970 (N_6970,N_4966,N_2526);
nand U6971 (N_6971,N_2557,N_4183);
nor U6972 (N_6972,N_3254,N_4905);
xnor U6973 (N_6973,N_4030,N_3698);
nand U6974 (N_6974,N_3442,N_2647);
nor U6975 (N_6975,N_4434,N_3318);
and U6976 (N_6976,N_3309,N_2519);
nor U6977 (N_6977,N_2835,N_3243);
and U6978 (N_6978,N_3278,N_4475);
nand U6979 (N_6979,N_3451,N_2757);
and U6980 (N_6980,N_3799,N_4075);
nand U6981 (N_6981,N_2534,N_2985);
nand U6982 (N_6982,N_4951,N_3344);
nand U6983 (N_6983,N_3623,N_4030);
nand U6984 (N_6984,N_2707,N_3603);
nand U6985 (N_6985,N_4624,N_3587);
nand U6986 (N_6986,N_4196,N_4749);
nand U6987 (N_6987,N_4371,N_4157);
or U6988 (N_6988,N_2808,N_4357);
nand U6989 (N_6989,N_4483,N_3575);
nand U6990 (N_6990,N_2867,N_3241);
nor U6991 (N_6991,N_4695,N_4611);
nor U6992 (N_6992,N_4010,N_4378);
or U6993 (N_6993,N_3154,N_2752);
and U6994 (N_6994,N_4029,N_3003);
or U6995 (N_6995,N_3420,N_4925);
nand U6996 (N_6996,N_3359,N_2796);
nand U6997 (N_6997,N_2685,N_2830);
nand U6998 (N_6998,N_2664,N_4580);
nand U6999 (N_6999,N_2748,N_3966);
and U7000 (N_7000,N_4890,N_4459);
xnor U7001 (N_7001,N_2804,N_3028);
or U7002 (N_7002,N_4897,N_3779);
nor U7003 (N_7003,N_4478,N_3018);
nand U7004 (N_7004,N_3668,N_3282);
or U7005 (N_7005,N_3449,N_4109);
nor U7006 (N_7006,N_2942,N_3499);
nand U7007 (N_7007,N_3175,N_2989);
or U7008 (N_7008,N_3022,N_4595);
and U7009 (N_7009,N_3830,N_3889);
nand U7010 (N_7010,N_4608,N_4477);
xor U7011 (N_7011,N_4249,N_4224);
nand U7012 (N_7012,N_4280,N_4527);
nor U7013 (N_7013,N_3848,N_2636);
nand U7014 (N_7014,N_3922,N_4142);
nand U7015 (N_7015,N_4139,N_4082);
nand U7016 (N_7016,N_4091,N_2994);
nor U7017 (N_7017,N_3334,N_4410);
and U7018 (N_7018,N_4496,N_3098);
nand U7019 (N_7019,N_2903,N_2849);
or U7020 (N_7020,N_3168,N_2569);
nand U7021 (N_7021,N_4957,N_3890);
nand U7022 (N_7022,N_3766,N_3207);
and U7023 (N_7023,N_3988,N_4755);
nand U7024 (N_7024,N_3606,N_3727);
and U7025 (N_7025,N_2845,N_3878);
or U7026 (N_7026,N_4296,N_3185);
or U7027 (N_7027,N_4361,N_2945);
xnor U7028 (N_7028,N_4590,N_4905);
and U7029 (N_7029,N_3898,N_2660);
nor U7030 (N_7030,N_4238,N_3883);
nand U7031 (N_7031,N_3658,N_3136);
nor U7032 (N_7032,N_3272,N_3394);
nand U7033 (N_7033,N_2775,N_3938);
or U7034 (N_7034,N_4350,N_4638);
nand U7035 (N_7035,N_2815,N_2864);
and U7036 (N_7036,N_3763,N_3301);
nor U7037 (N_7037,N_4860,N_4337);
xnor U7038 (N_7038,N_3677,N_4052);
nor U7039 (N_7039,N_4431,N_2624);
nand U7040 (N_7040,N_4557,N_2858);
nand U7041 (N_7041,N_3840,N_4221);
or U7042 (N_7042,N_2740,N_3408);
and U7043 (N_7043,N_4147,N_3376);
nand U7044 (N_7044,N_4179,N_3025);
nor U7045 (N_7045,N_4099,N_4379);
nor U7046 (N_7046,N_3543,N_2583);
nor U7047 (N_7047,N_4061,N_3813);
nand U7048 (N_7048,N_4692,N_3370);
and U7049 (N_7049,N_4933,N_3151);
nor U7050 (N_7050,N_4169,N_2662);
and U7051 (N_7051,N_4071,N_4233);
nand U7052 (N_7052,N_4447,N_2528);
nand U7053 (N_7053,N_3946,N_4660);
nor U7054 (N_7054,N_2815,N_2836);
xnor U7055 (N_7055,N_4547,N_4768);
nor U7056 (N_7056,N_3481,N_3714);
or U7057 (N_7057,N_4125,N_4503);
and U7058 (N_7058,N_3960,N_4172);
nor U7059 (N_7059,N_4617,N_3003);
or U7060 (N_7060,N_4755,N_4688);
and U7061 (N_7061,N_4750,N_3583);
or U7062 (N_7062,N_3674,N_4742);
or U7063 (N_7063,N_4538,N_3528);
nor U7064 (N_7064,N_3203,N_2950);
or U7065 (N_7065,N_3124,N_3695);
or U7066 (N_7066,N_3720,N_2947);
or U7067 (N_7067,N_2989,N_2562);
nor U7068 (N_7068,N_2587,N_4573);
xor U7069 (N_7069,N_2765,N_3405);
nand U7070 (N_7070,N_3657,N_3301);
nand U7071 (N_7071,N_3622,N_3770);
nor U7072 (N_7072,N_4367,N_4897);
nand U7073 (N_7073,N_3962,N_4593);
or U7074 (N_7074,N_2750,N_3342);
nand U7075 (N_7075,N_3329,N_3595);
or U7076 (N_7076,N_2561,N_4240);
nor U7077 (N_7077,N_2695,N_3698);
xor U7078 (N_7078,N_3532,N_2657);
nor U7079 (N_7079,N_4167,N_4873);
xor U7080 (N_7080,N_3547,N_3493);
or U7081 (N_7081,N_3974,N_4056);
nor U7082 (N_7082,N_3005,N_4511);
and U7083 (N_7083,N_3167,N_3534);
xnor U7084 (N_7084,N_3059,N_2855);
or U7085 (N_7085,N_4564,N_4144);
nor U7086 (N_7086,N_4097,N_4258);
and U7087 (N_7087,N_2630,N_4670);
and U7088 (N_7088,N_3641,N_2730);
and U7089 (N_7089,N_3204,N_2771);
nand U7090 (N_7090,N_4120,N_4140);
nand U7091 (N_7091,N_4495,N_3151);
nand U7092 (N_7092,N_3917,N_3913);
nor U7093 (N_7093,N_4061,N_4226);
nor U7094 (N_7094,N_2918,N_4830);
xor U7095 (N_7095,N_4440,N_2703);
or U7096 (N_7096,N_4683,N_3475);
nand U7097 (N_7097,N_2824,N_2646);
nand U7098 (N_7098,N_4253,N_3485);
nand U7099 (N_7099,N_4662,N_4706);
or U7100 (N_7100,N_3836,N_4786);
or U7101 (N_7101,N_2893,N_3435);
xnor U7102 (N_7102,N_4243,N_4014);
and U7103 (N_7103,N_3628,N_3667);
and U7104 (N_7104,N_4460,N_4542);
nor U7105 (N_7105,N_3449,N_4633);
nand U7106 (N_7106,N_4738,N_3829);
nand U7107 (N_7107,N_4715,N_3130);
nor U7108 (N_7108,N_2519,N_3218);
or U7109 (N_7109,N_3653,N_2784);
nand U7110 (N_7110,N_3648,N_3007);
and U7111 (N_7111,N_2832,N_3919);
nand U7112 (N_7112,N_3004,N_4646);
xnor U7113 (N_7113,N_3924,N_2665);
nand U7114 (N_7114,N_4673,N_3663);
nor U7115 (N_7115,N_3049,N_4556);
nand U7116 (N_7116,N_2977,N_3187);
xnor U7117 (N_7117,N_3653,N_4376);
and U7118 (N_7118,N_4870,N_4070);
nor U7119 (N_7119,N_2687,N_4028);
and U7120 (N_7120,N_3077,N_4861);
xnor U7121 (N_7121,N_4939,N_3009);
or U7122 (N_7122,N_3498,N_2938);
or U7123 (N_7123,N_4171,N_3092);
nor U7124 (N_7124,N_4186,N_3780);
or U7125 (N_7125,N_3128,N_2691);
nor U7126 (N_7126,N_2635,N_4850);
xor U7127 (N_7127,N_4659,N_4196);
nand U7128 (N_7128,N_3477,N_2669);
nand U7129 (N_7129,N_3521,N_3307);
and U7130 (N_7130,N_3125,N_2767);
nor U7131 (N_7131,N_3119,N_4357);
nand U7132 (N_7132,N_2603,N_3497);
or U7133 (N_7133,N_3340,N_3760);
xnor U7134 (N_7134,N_3616,N_2985);
and U7135 (N_7135,N_2913,N_3313);
nand U7136 (N_7136,N_3893,N_3550);
nand U7137 (N_7137,N_4364,N_3057);
nor U7138 (N_7138,N_2889,N_3221);
or U7139 (N_7139,N_2565,N_4427);
and U7140 (N_7140,N_4644,N_4914);
nand U7141 (N_7141,N_4889,N_4657);
xor U7142 (N_7142,N_4954,N_4586);
nand U7143 (N_7143,N_4126,N_3808);
and U7144 (N_7144,N_2678,N_2596);
nand U7145 (N_7145,N_2935,N_4297);
nand U7146 (N_7146,N_4327,N_3147);
nand U7147 (N_7147,N_3284,N_3784);
and U7148 (N_7148,N_4257,N_3518);
nand U7149 (N_7149,N_4493,N_3941);
nand U7150 (N_7150,N_3564,N_4112);
and U7151 (N_7151,N_2523,N_3070);
and U7152 (N_7152,N_4818,N_3955);
nor U7153 (N_7153,N_4751,N_4049);
nand U7154 (N_7154,N_2528,N_3369);
and U7155 (N_7155,N_2624,N_3654);
nand U7156 (N_7156,N_3458,N_3648);
nor U7157 (N_7157,N_4509,N_3564);
nand U7158 (N_7158,N_2583,N_4941);
nor U7159 (N_7159,N_3675,N_3997);
or U7160 (N_7160,N_3638,N_4023);
or U7161 (N_7161,N_2722,N_3009);
and U7162 (N_7162,N_3838,N_2538);
and U7163 (N_7163,N_2949,N_3465);
nand U7164 (N_7164,N_3038,N_4102);
and U7165 (N_7165,N_4289,N_4079);
nand U7166 (N_7166,N_4789,N_2612);
xnor U7167 (N_7167,N_3991,N_3356);
xnor U7168 (N_7168,N_4534,N_3563);
or U7169 (N_7169,N_3352,N_4808);
and U7170 (N_7170,N_3322,N_2763);
nand U7171 (N_7171,N_3146,N_4551);
nor U7172 (N_7172,N_3429,N_4526);
nand U7173 (N_7173,N_3279,N_2749);
or U7174 (N_7174,N_4318,N_4600);
or U7175 (N_7175,N_2553,N_2508);
or U7176 (N_7176,N_4254,N_4804);
or U7177 (N_7177,N_4291,N_2658);
and U7178 (N_7178,N_4204,N_4523);
or U7179 (N_7179,N_2558,N_3898);
nor U7180 (N_7180,N_4141,N_3918);
nand U7181 (N_7181,N_3267,N_3205);
and U7182 (N_7182,N_3562,N_3508);
and U7183 (N_7183,N_2715,N_3537);
or U7184 (N_7184,N_2896,N_3992);
nor U7185 (N_7185,N_4289,N_2860);
or U7186 (N_7186,N_3582,N_2504);
nand U7187 (N_7187,N_3995,N_3822);
nor U7188 (N_7188,N_3600,N_2868);
xor U7189 (N_7189,N_3744,N_4513);
or U7190 (N_7190,N_4514,N_2829);
or U7191 (N_7191,N_3259,N_3358);
and U7192 (N_7192,N_4702,N_3966);
or U7193 (N_7193,N_3523,N_4895);
and U7194 (N_7194,N_4791,N_3210);
or U7195 (N_7195,N_4337,N_4971);
or U7196 (N_7196,N_3643,N_4868);
and U7197 (N_7197,N_2775,N_4271);
nor U7198 (N_7198,N_4047,N_3562);
nand U7199 (N_7199,N_3987,N_2668);
nand U7200 (N_7200,N_2951,N_2663);
or U7201 (N_7201,N_2974,N_4456);
or U7202 (N_7202,N_4938,N_4676);
nor U7203 (N_7203,N_3284,N_3118);
or U7204 (N_7204,N_4100,N_3850);
and U7205 (N_7205,N_4875,N_3288);
nand U7206 (N_7206,N_2902,N_3469);
nand U7207 (N_7207,N_4469,N_2549);
nor U7208 (N_7208,N_3724,N_3924);
xnor U7209 (N_7209,N_4082,N_4195);
or U7210 (N_7210,N_3917,N_3933);
nand U7211 (N_7211,N_4329,N_3522);
xor U7212 (N_7212,N_4453,N_3073);
nand U7213 (N_7213,N_2731,N_3985);
nor U7214 (N_7214,N_4571,N_2739);
nand U7215 (N_7215,N_2975,N_4056);
or U7216 (N_7216,N_3740,N_2857);
and U7217 (N_7217,N_2652,N_4430);
and U7218 (N_7218,N_4903,N_4243);
or U7219 (N_7219,N_2581,N_3406);
nor U7220 (N_7220,N_3536,N_2504);
xnor U7221 (N_7221,N_4780,N_3688);
and U7222 (N_7222,N_4926,N_2567);
and U7223 (N_7223,N_2533,N_3280);
or U7224 (N_7224,N_4511,N_3731);
xnor U7225 (N_7225,N_2728,N_3549);
and U7226 (N_7226,N_4038,N_4867);
and U7227 (N_7227,N_3652,N_4616);
or U7228 (N_7228,N_4513,N_4346);
and U7229 (N_7229,N_4173,N_3700);
or U7230 (N_7230,N_3493,N_3827);
and U7231 (N_7231,N_3231,N_4945);
and U7232 (N_7232,N_4409,N_4431);
or U7233 (N_7233,N_3552,N_4838);
nand U7234 (N_7234,N_4273,N_3061);
and U7235 (N_7235,N_4988,N_4109);
nand U7236 (N_7236,N_2722,N_4970);
nand U7237 (N_7237,N_4489,N_3102);
and U7238 (N_7238,N_4846,N_2592);
and U7239 (N_7239,N_2846,N_4971);
or U7240 (N_7240,N_3221,N_3534);
and U7241 (N_7241,N_4087,N_4001);
or U7242 (N_7242,N_2892,N_4114);
nand U7243 (N_7243,N_4867,N_3699);
nand U7244 (N_7244,N_3896,N_4419);
or U7245 (N_7245,N_3915,N_3673);
nand U7246 (N_7246,N_4534,N_3797);
or U7247 (N_7247,N_4441,N_3008);
or U7248 (N_7248,N_2978,N_4373);
or U7249 (N_7249,N_2948,N_3526);
nor U7250 (N_7250,N_2868,N_3719);
nand U7251 (N_7251,N_3360,N_3324);
nor U7252 (N_7252,N_3826,N_4830);
xnor U7253 (N_7253,N_4086,N_4809);
nand U7254 (N_7254,N_3433,N_4970);
nor U7255 (N_7255,N_4677,N_4336);
or U7256 (N_7256,N_4739,N_4312);
and U7257 (N_7257,N_4130,N_2776);
and U7258 (N_7258,N_3973,N_4709);
xnor U7259 (N_7259,N_2587,N_4632);
nand U7260 (N_7260,N_4189,N_4035);
and U7261 (N_7261,N_2826,N_3457);
or U7262 (N_7262,N_4637,N_4905);
or U7263 (N_7263,N_4943,N_2966);
nor U7264 (N_7264,N_2688,N_4922);
xnor U7265 (N_7265,N_4509,N_4895);
nor U7266 (N_7266,N_3040,N_4744);
nor U7267 (N_7267,N_4481,N_4855);
nand U7268 (N_7268,N_4387,N_4983);
xor U7269 (N_7269,N_3664,N_4664);
or U7270 (N_7270,N_2828,N_4576);
or U7271 (N_7271,N_4360,N_4962);
nor U7272 (N_7272,N_4525,N_3397);
and U7273 (N_7273,N_3842,N_4207);
and U7274 (N_7274,N_2596,N_2854);
xor U7275 (N_7275,N_3627,N_3473);
and U7276 (N_7276,N_4554,N_4615);
or U7277 (N_7277,N_3219,N_3220);
or U7278 (N_7278,N_3058,N_3674);
or U7279 (N_7279,N_4367,N_4839);
and U7280 (N_7280,N_4624,N_3479);
nand U7281 (N_7281,N_3044,N_3508);
nor U7282 (N_7282,N_2592,N_3606);
nor U7283 (N_7283,N_4175,N_3546);
nor U7284 (N_7284,N_2973,N_4918);
nand U7285 (N_7285,N_2914,N_4655);
or U7286 (N_7286,N_2696,N_4623);
and U7287 (N_7287,N_2500,N_4722);
nand U7288 (N_7288,N_4977,N_3736);
nand U7289 (N_7289,N_4370,N_3359);
xor U7290 (N_7290,N_2634,N_4534);
or U7291 (N_7291,N_2971,N_2871);
xor U7292 (N_7292,N_4251,N_3362);
nand U7293 (N_7293,N_4723,N_2777);
xor U7294 (N_7294,N_3916,N_3904);
and U7295 (N_7295,N_2874,N_3712);
nor U7296 (N_7296,N_2675,N_4063);
nor U7297 (N_7297,N_4050,N_3868);
or U7298 (N_7298,N_3502,N_2957);
nor U7299 (N_7299,N_3638,N_4564);
xnor U7300 (N_7300,N_4332,N_2967);
and U7301 (N_7301,N_2999,N_3956);
nor U7302 (N_7302,N_4646,N_3422);
and U7303 (N_7303,N_2669,N_3432);
and U7304 (N_7304,N_4131,N_3638);
and U7305 (N_7305,N_4920,N_3517);
and U7306 (N_7306,N_3835,N_4813);
and U7307 (N_7307,N_4700,N_3999);
and U7308 (N_7308,N_3864,N_4732);
nor U7309 (N_7309,N_3805,N_3894);
nand U7310 (N_7310,N_3136,N_4151);
and U7311 (N_7311,N_4359,N_3659);
nor U7312 (N_7312,N_3905,N_4195);
nor U7313 (N_7313,N_4705,N_3794);
nor U7314 (N_7314,N_4531,N_3660);
nor U7315 (N_7315,N_4318,N_4434);
nand U7316 (N_7316,N_4251,N_3300);
nand U7317 (N_7317,N_4195,N_4793);
xor U7318 (N_7318,N_4525,N_4244);
xnor U7319 (N_7319,N_3947,N_3922);
nor U7320 (N_7320,N_4688,N_2531);
and U7321 (N_7321,N_3150,N_4020);
nand U7322 (N_7322,N_2610,N_2521);
and U7323 (N_7323,N_3897,N_4601);
or U7324 (N_7324,N_4395,N_2717);
nand U7325 (N_7325,N_3702,N_2859);
xnor U7326 (N_7326,N_4286,N_2969);
nand U7327 (N_7327,N_3233,N_4054);
nand U7328 (N_7328,N_4880,N_3162);
and U7329 (N_7329,N_2513,N_3514);
and U7330 (N_7330,N_3670,N_2950);
nand U7331 (N_7331,N_3931,N_3975);
and U7332 (N_7332,N_4285,N_3032);
or U7333 (N_7333,N_4142,N_4201);
and U7334 (N_7334,N_4293,N_3253);
or U7335 (N_7335,N_4153,N_2801);
and U7336 (N_7336,N_4359,N_3270);
or U7337 (N_7337,N_3722,N_4936);
nand U7338 (N_7338,N_4044,N_3042);
and U7339 (N_7339,N_4732,N_4684);
nor U7340 (N_7340,N_3115,N_3612);
nor U7341 (N_7341,N_4480,N_3716);
and U7342 (N_7342,N_3373,N_3973);
nor U7343 (N_7343,N_4328,N_4937);
nor U7344 (N_7344,N_3222,N_2916);
nand U7345 (N_7345,N_3894,N_4414);
nor U7346 (N_7346,N_4417,N_4775);
nor U7347 (N_7347,N_3176,N_3038);
and U7348 (N_7348,N_3434,N_4512);
or U7349 (N_7349,N_2941,N_2663);
nor U7350 (N_7350,N_4521,N_4895);
or U7351 (N_7351,N_3400,N_3827);
and U7352 (N_7352,N_3161,N_4242);
and U7353 (N_7353,N_3207,N_2763);
and U7354 (N_7354,N_3087,N_3001);
nand U7355 (N_7355,N_4790,N_2670);
nand U7356 (N_7356,N_3716,N_2801);
xnor U7357 (N_7357,N_4106,N_3977);
nand U7358 (N_7358,N_4276,N_3463);
nand U7359 (N_7359,N_4577,N_3464);
and U7360 (N_7360,N_4529,N_2556);
or U7361 (N_7361,N_4906,N_2983);
and U7362 (N_7362,N_2742,N_3594);
nor U7363 (N_7363,N_3470,N_4218);
nor U7364 (N_7364,N_3555,N_4452);
nor U7365 (N_7365,N_3381,N_3183);
or U7366 (N_7366,N_4719,N_4077);
and U7367 (N_7367,N_2748,N_3767);
nor U7368 (N_7368,N_3955,N_3268);
and U7369 (N_7369,N_4200,N_4223);
or U7370 (N_7370,N_4392,N_4367);
or U7371 (N_7371,N_4735,N_3330);
xnor U7372 (N_7372,N_2923,N_3090);
nor U7373 (N_7373,N_3521,N_3825);
and U7374 (N_7374,N_3926,N_2854);
nor U7375 (N_7375,N_4401,N_3184);
nand U7376 (N_7376,N_4886,N_2754);
or U7377 (N_7377,N_4916,N_3323);
nor U7378 (N_7378,N_3327,N_3263);
nand U7379 (N_7379,N_4086,N_4322);
and U7380 (N_7380,N_3067,N_2575);
nor U7381 (N_7381,N_2980,N_3854);
nor U7382 (N_7382,N_3487,N_3697);
and U7383 (N_7383,N_4814,N_3775);
and U7384 (N_7384,N_4306,N_4961);
nand U7385 (N_7385,N_4251,N_3686);
nor U7386 (N_7386,N_3057,N_3237);
nor U7387 (N_7387,N_3836,N_3623);
nand U7388 (N_7388,N_3093,N_3969);
and U7389 (N_7389,N_2586,N_2921);
nand U7390 (N_7390,N_2718,N_2546);
or U7391 (N_7391,N_3821,N_2684);
xnor U7392 (N_7392,N_3318,N_2511);
nor U7393 (N_7393,N_3444,N_3654);
nor U7394 (N_7394,N_3785,N_3209);
xor U7395 (N_7395,N_3170,N_3880);
and U7396 (N_7396,N_4091,N_4593);
nand U7397 (N_7397,N_3122,N_2807);
nand U7398 (N_7398,N_2823,N_3819);
and U7399 (N_7399,N_3511,N_3831);
nor U7400 (N_7400,N_3891,N_3512);
or U7401 (N_7401,N_4703,N_3222);
nor U7402 (N_7402,N_3750,N_3311);
and U7403 (N_7403,N_2652,N_3015);
and U7404 (N_7404,N_3046,N_3988);
nor U7405 (N_7405,N_3042,N_3582);
or U7406 (N_7406,N_4011,N_3589);
or U7407 (N_7407,N_3950,N_3770);
and U7408 (N_7408,N_2535,N_4014);
nor U7409 (N_7409,N_2642,N_4543);
xor U7410 (N_7410,N_2770,N_4332);
and U7411 (N_7411,N_4542,N_4045);
or U7412 (N_7412,N_3267,N_3390);
or U7413 (N_7413,N_4677,N_3599);
and U7414 (N_7414,N_4597,N_4685);
nand U7415 (N_7415,N_4253,N_3066);
xor U7416 (N_7416,N_4884,N_4107);
nand U7417 (N_7417,N_2564,N_3858);
nand U7418 (N_7418,N_3213,N_4627);
xor U7419 (N_7419,N_4894,N_3201);
nand U7420 (N_7420,N_2588,N_4116);
nor U7421 (N_7421,N_2750,N_4186);
and U7422 (N_7422,N_4965,N_4454);
nor U7423 (N_7423,N_4794,N_4826);
and U7424 (N_7424,N_3778,N_4210);
nand U7425 (N_7425,N_4076,N_2667);
nor U7426 (N_7426,N_4294,N_3490);
nor U7427 (N_7427,N_2636,N_3751);
or U7428 (N_7428,N_4474,N_4395);
and U7429 (N_7429,N_2547,N_2929);
and U7430 (N_7430,N_4986,N_3816);
and U7431 (N_7431,N_2570,N_3988);
xor U7432 (N_7432,N_4746,N_4031);
or U7433 (N_7433,N_3770,N_4767);
or U7434 (N_7434,N_2818,N_3533);
and U7435 (N_7435,N_4127,N_4421);
or U7436 (N_7436,N_4529,N_4823);
xnor U7437 (N_7437,N_3415,N_3253);
and U7438 (N_7438,N_4157,N_3400);
xnor U7439 (N_7439,N_2742,N_4998);
and U7440 (N_7440,N_4633,N_3259);
or U7441 (N_7441,N_3834,N_2719);
and U7442 (N_7442,N_3878,N_3094);
and U7443 (N_7443,N_4738,N_3081);
or U7444 (N_7444,N_4935,N_3495);
or U7445 (N_7445,N_4016,N_4491);
and U7446 (N_7446,N_3831,N_2732);
nand U7447 (N_7447,N_3201,N_4585);
or U7448 (N_7448,N_3130,N_4770);
and U7449 (N_7449,N_3329,N_3341);
and U7450 (N_7450,N_4273,N_4899);
and U7451 (N_7451,N_3970,N_4331);
xnor U7452 (N_7452,N_4664,N_3875);
or U7453 (N_7453,N_3357,N_4865);
nor U7454 (N_7454,N_4768,N_3256);
or U7455 (N_7455,N_3614,N_3003);
nand U7456 (N_7456,N_4587,N_2822);
or U7457 (N_7457,N_3314,N_2728);
and U7458 (N_7458,N_2673,N_2512);
or U7459 (N_7459,N_3896,N_4975);
nand U7460 (N_7460,N_4628,N_4076);
nor U7461 (N_7461,N_3290,N_4697);
or U7462 (N_7462,N_2761,N_4466);
or U7463 (N_7463,N_4014,N_3746);
or U7464 (N_7464,N_4385,N_2779);
nand U7465 (N_7465,N_4134,N_3573);
nor U7466 (N_7466,N_2816,N_4384);
or U7467 (N_7467,N_3880,N_2605);
nand U7468 (N_7468,N_4240,N_3938);
and U7469 (N_7469,N_4849,N_3837);
nand U7470 (N_7470,N_4416,N_3734);
xor U7471 (N_7471,N_4575,N_3504);
or U7472 (N_7472,N_4873,N_4957);
or U7473 (N_7473,N_3487,N_4261);
and U7474 (N_7474,N_4808,N_4104);
or U7475 (N_7475,N_4507,N_2531);
nand U7476 (N_7476,N_4769,N_3048);
nand U7477 (N_7477,N_4292,N_4571);
xnor U7478 (N_7478,N_4849,N_3002);
or U7479 (N_7479,N_3436,N_3652);
or U7480 (N_7480,N_3573,N_2573);
and U7481 (N_7481,N_2746,N_3545);
and U7482 (N_7482,N_3374,N_3175);
nand U7483 (N_7483,N_3065,N_2928);
and U7484 (N_7484,N_3826,N_2982);
nor U7485 (N_7485,N_3165,N_2608);
or U7486 (N_7486,N_3482,N_4124);
and U7487 (N_7487,N_3942,N_4910);
and U7488 (N_7488,N_4116,N_3901);
nor U7489 (N_7489,N_4918,N_4168);
nand U7490 (N_7490,N_3037,N_2742);
nand U7491 (N_7491,N_4227,N_2751);
and U7492 (N_7492,N_4049,N_3218);
and U7493 (N_7493,N_2767,N_3986);
and U7494 (N_7494,N_4060,N_2733);
xor U7495 (N_7495,N_3264,N_4723);
nand U7496 (N_7496,N_3951,N_4565);
nand U7497 (N_7497,N_3962,N_4531);
nand U7498 (N_7498,N_4839,N_3587);
nor U7499 (N_7499,N_3830,N_4293);
and U7500 (N_7500,N_6150,N_7261);
xor U7501 (N_7501,N_7178,N_7065);
nor U7502 (N_7502,N_5307,N_5193);
nor U7503 (N_7503,N_5287,N_6666);
nand U7504 (N_7504,N_6165,N_5468);
nor U7505 (N_7505,N_7429,N_6289);
and U7506 (N_7506,N_6352,N_7066);
and U7507 (N_7507,N_6169,N_6513);
xnor U7508 (N_7508,N_5688,N_5346);
nor U7509 (N_7509,N_6815,N_6397);
nand U7510 (N_7510,N_5113,N_5571);
and U7511 (N_7511,N_5063,N_5845);
and U7512 (N_7512,N_6212,N_5835);
nand U7513 (N_7513,N_5487,N_6453);
or U7514 (N_7514,N_6442,N_6180);
nor U7515 (N_7515,N_7370,N_6953);
nor U7516 (N_7516,N_5486,N_6426);
and U7517 (N_7517,N_5036,N_6570);
nand U7518 (N_7518,N_7302,N_5413);
and U7519 (N_7519,N_5707,N_7124);
nand U7520 (N_7520,N_6187,N_5252);
nand U7521 (N_7521,N_6646,N_5878);
and U7522 (N_7522,N_6300,N_6901);
or U7523 (N_7523,N_5492,N_5118);
and U7524 (N_7524,N_6038,N_5148);
or U7525 (N_7525,N_6438,N_6896);
nor U7526 (N_7526,N_6299,N_5671);
nor U7527 (N_7527,N_6132,N_6813);
nand U7528 (N_7528,N_5777,N_7329);
nand U7529 (N_7529,N_7256,N_6204);
nand U7530 (N_7530,N_7001,N_7484);
nor U7531 (N_7531,N_6285,N_6358);
nand U7532 (N_7532,N_6366,N_5430);
or U7533 (N_7533,N_6819,N_7478);
nor U7534 (N_7534,N_5691,N_5060);
or U7535 (N_7535,N_7352,N_6529);
nor U7536 (N_7536,N_7462,N_6086);
nand U7537 (N_7537,N_6364,N_6807);
or U7538 (N_7538,N_5187,N_7092);
nand U7539 (N_7539,N_6345,N_5555);
or U7540 (N_7540,N_7162,N_6635);
nor U7541 (N_7541,N_6452,N_6462);
or U7542 (N_7542,N_5419,N_6724);
or U7543 (N_7543,N_6488,N_6975);
nand U7544 (N_7544,N_6247,N_5224);
and U7545 (N_7545,N_6855,N_5617);
nor U7546 (N_7546,N_6429,N_5935);
nor U7547 (N_7547,N_7368,N_5447);
or U7548 (N_7548,N_7167,N_5397);
or U7549 (N_7549,N_6142,N_6337);
nor U7550 (N_7550,N_7123,N_6129);
xnor U7551 (N_7551,N_7490,N_7436);
and U7552 (N_7552,N_6005,N_5647);
or U7553 (N_7553,N_5998,N_6049);
and U7554 (N_7554,N_6868,N_6259);
and U7555 (N_7555,N_5827,N_5303);
nor U7556 (N_7556,N_7037,N_7276);
or U7557 (N_7557,N_6680,N_5169);
nand U7558 (N_7558,N_6408,N_6054);
nor U7559 (N_7559,N_6088,N_7259);
nor U7560 (N_7560,N_6295,N_6475);
and U7561 (N_7561,N_6441,N_5210);
or U7562 (N_7562,N_6746,N_5417);
and U7563 (N_7563,N_5191,N_7392);
nand U7564 (N_7564,N_6261,N_6422);
nor U7565 (N_7565,N_7232,N_5585);
nor U7566 (N_7566,N_7204,N_7053);
or U7567 (N_7567,N_5847,N_5257);
and U7568 (N_7568,N_6158,N_6319);
nor U7569 (N_7569,N_5400,N_7113);
and U7570 (N_7570,N_6937,N_7190);
and U7571 (N_7571,N_6179,N_6772);
or U7572 (N_7572,N_6531,N_5043);
nor U7573 (N_7573,N_6239,N_7450);
or U7574 (N_7574,N_5735,N_6713);
nor U7575 (N_7575,N_5007,N_7476);
nor U7576 (N_7576,N_7347,N_5031);
or U7577 (N_7577,N_5629,N_5828);
or U7578 (N_7578,N_6178,N_6788);
nor U7579 (N_7579,N_7128,N_5919);
nand U7580 (N_7580,N_5609,N_6560);
nand U7581 (N_7581,N_5112,N_5124);
nand U7582 (N_7582,N_6501,N_7181);
xnor U7583 (N_7583,N_5258,N_5453);
or U7584 (N_7584,N_7293,N_5683);
or U7585 (N_7585,N_6894,N_6351);
or U7586 (N_7586,N_5752,N_6465);
nand U7587 (N_7587,N_6828,N_5766);
xor U7588 (N_7588,N_7015,N_5416);
and U7589 (N_7589,N_7254,N_5597);
nand U7590 (N_7590,N_5668,N_6495);
and U7591 (N_7591,N_6638,N_6837);
or U7592 (N_7592,N_5697,N_5563);
xor U7593 (N_7593,N_6954,N_5032);
nor U7594 (N_7594,N_7189,N_6175);
nor U7595 (N_7595,N_7220,N_6682);
nand U7596 (N_7596,N_6549,N_7471);
or U7597 (N_7597,N_6060,N_5738);
nor U7598 (N_7598,N_6105,N_5464);
and U7599 (N_7599,N_5232,N_5842);
nand U7600 (N_7600,N_6955,N_5675);
or U7601 (N_7601,N_5839,N_6334);
and U7602 (N_7602,N_5189,N_7454);
and U7603 (N_7603,N_6434,N_5913);
and U7604 (N_7604,N_6022,N_7393);
nand U7605 (N_7605,N_6691,N_6630);
nor U7606 (N_7606,N_5729,N_5127);
or U7607 (N_7607,N_6192,N_6144);
xnor U7608 (N_7608,N_5764,N_5944);
nand U7609 (N_7609,N_5182,N_5472);
or U7610 (N_7610,N_5573,N_6835);
or U7611 (N_7611,N_5361,N_6190);
and U7612 (N_7612,N_6493,N_5214);
and U7613 (N_7613,N_5639,N_5657);
nor U7614 (N_7614,N_5851,N_6653);
and U7615 (N_7615,N_6322,N_5605);
nor U7616 (N_7616,N_6803,N_6554);
nor U7617 (N_7617,N_6654,N_6193);
nand U7618 (N_7618,N_7428,N_6454);
or U7619 (N_7619,N_7332,N_5634);
nor U7620 (N_7620,N_7023,N_5785);
or U7621 (N_7621,N_5104,N_5306);
nor U7622 (N_7622,N_5779,N_5446);
xor U7623 (N_7623,N_7260,N_6237);
xnor U7624 (N_7624,N_7299,N_6384);
and U7625 (N_7625,N_5199,N_6128);
nor U7626 (N_7626,N_5864,N_5583);
xnor U7627 (N_7627,N_5511,N_7375);
or U7628 (N_7628,N_5497,N_6738);
and U7629 (N_7629,N_6057,N_5964);
or U7630 (N_7630,N_6458,N_6795);
nand U7631 (N_7631,N_5575,N_6845);
nand U7632 (N_7632,N_7283,N_7225);
nand U7633 (N_7633,N_6032,N_5577);
or U7634 (N_7634,N_6025,N_5283);
nor U7635 (N_7635,N_6498,N_6971);
or U7636 (N_7636,N_5372,N_5427);
nor U7637 (N_7637,N_5068,N_5170);
and U7638 (N_7638,N_5758,N_7487);
or U7639 (N_7639,N_5392,N_7343);
nand U7640 (N_7640,N_6238,N_6652);
nand U7641 (N_7641,N_6028,N_6817);
and U7642 (N_7642,N_5906,N_6913);
nand U7643 (N_7643,N_5667,N_6396);
xor U7644 (N_7644,N_6466,N_6866);
nor U7645 (N_7645,N_5314,N_5491);
and U7646 (N_7646,N_5876,N_5892);
nor U7647 (N_7647,N_6936,N_6849);
or U7648 (N_7648,N_6348,N_5882);
nand U7649 (N_7649,N_7154,N_5207);
nor U7650 (N_7650,N_7117,N_5601);
and U7651 (N_7651,N_5374,N_7390);
nand U7652 (N_7652,N_5734,N_7467);
or U7653 (N_7653,N_6555,N_6917);
nand U7654 (N_7654,N_6127,N_5884);
nand U7655 (N_7655,N_6891,N_5620);
nor U7656 (N_7656,N_5793,N_7337);
xor U7657 (N_7657,N_6869,N_5753);
and U7658 (N_7658,N_6617,N_6412);
or U7659 (N_7659,N_6651,N_6997);
and U7660 (N_7660,N_7074,N_5260);
nand U7661 (N_7661,N_6573,N_5650);
and U7662 (N_7662,N_5805,N_5269);
and U7663 (N_7663,N_5690,N_7272);
nand U7664 (N_7664,N_6659,N_5602);
or U7665 (N_7665,N_5975,N_6504);
nor U7666 (N_7666,N_6497,N_7342);
and U7667 (N_7667,N_5968,N_6760);
nor U7668 (N_7668,N_6419,N_6935);
and U7669 (N_7669,N_6643,N_5005);
or U7670 (N_7670,N_6339,N_5014);
or U7671 (N_7671,N_6544,N_5165);
nor U7672 (N_7672,N_5740,N_5941);
nor U7673 (N_7673,N_6590,N_5593);
nand U7674 (N_7674,N_5698,N_7325);
and U7675 (N_7675,N_6398,N_7383);
or U7676 (N_7676,N_7222,N_6741);
nand U7677 (N_7677,N_6965,N_7151);
and U7678 (N_7678,N_6061,N_6562);
and U7679 (N_7679,N_6494,N_5881);
nand U7680 (N_7680,N_6904,N_7381);
or U7681 (N_7681,N_6000,N_6679);
xnor U7682 (N_7682,N_5143,N_5772);
nand U7683 (N_7683,N_5385,N_6723);
nor U7684 (N_7684,N_7287,N_5613);
nand U7685 (N_7685,N_5358,N_5188);
nor U7686 (N_7686,N_7046,N_5808);
nand U7687 (N_7687,N_6140,N_7061);
or U7688 (N_7688,N_6897,N_6628);
or U7689 (N_7689,N_7042,N_6787);
nand U7690 (N_7690,N_7069,N_6314);
nand U7691 (N_7691,N_5404,N_6704);
or U7692 (N_7692,N_6424,N_7281);
nor U7693 (N_7693,N_5840,N_7071);
and U7694 (N_7694,N_5412,N_5539);
nand U7695 (N_7695,N_7171,N_6533);
xnor U7696 (N_7696,N_5322,N_6588);
nor U7697 (N_7697,N_7278,N_6149);
and U7698 (N_7698,N_6410,N_6737);
nand U7699 (N_7699,N_5332,N_6539);
and U7700 (N_7700,N_5423,N_6026);
and U7701 (N_7701,N_6446,N_6568);
and U7702 (N_7702,N_5426,N_6722);
nor U7703 (N_7703,N_5706,N_7206);
or U7704 (N_7704,N_5529,N_6739);
xor U7705 (N_7705,N_5353,N_6382);
nand U7706 (N_7706,N_5560,N_6431);
or U7707 (N_7707,N_7142,N_6847);
nand U7708 (N_7708,N_7280,N_7406);
nor U7709 (N_7709,N_6051,N_5564);
or U7710 (N_7710,N_6618,N_6268);
nand U7711 (N_7711,N_6296,N_5717);
or U7712 (N_7712,N_5556,N_6078);
nand U7713 (N_7713,N_7303,N_7183);
and U7714 (N_7714,N_5774,N_7161);
or U7715 (N_7715,N_6377,N_5645);
xor U7716 (N_7716,N_5438,N_6963);
nor U7717 (N_7717,N_5147,N_5598);
xnor U7718 (N_7718,N_6610,N_6068);
and U7719 (N_7719,N_5745,N_5914);
and U7720 (N_7720,N_5172,N_5183);
nand U7721 (N_7721,N_7486,N_5538);
xnor U7722 (N_7722,N_6075,N_5646);
nand U7723 (N_7723,N_6794,N_6425);
nor U7724 (N_7724,N_7099,N_5970);
nand U7725 (N_7725,N_7266,N_5027);
nor U7726 (N_7726,N_7039,N_5259);
nor U7727 (N_7727,N_5225,N_7473);
and U7728 (N_7728,N_7300,N_5162);
and U7729 (N_7729,N_6716,N_7141);
nand U7730 (N_7730,N_5315,N_6225);
nor U7731 (N_7731,N_7470,N_7430);
xnor U7732 (N_7732,N_5496,N_6706);
or U7733 (N_7733,N_5439,N_6899);
and U7734 (N_7734,N_5139,N_7267);
nor U7735 (N_7735,N_6589,N_5972);
nand U7736 (N_7736,N_6265,N_6644);
nor U7737 (N_7737,N_5985,N_7401);
or U7738 (N_7738,N_5362,N_5507);
and U7739 (N_7739,N_5720,N_5503);
nand U7740 (N_7740,N_7115,N_6229);
nor U7741 (N_7741,N_7415,N_6934);
nor U7742 (N_7742,N_5452,N_6689);
nand U7743 (N_7743,N_5903,N_5481);
and U7744 (N_7744,N_7120,N_5278);
or U7745 (N_7745,N_6566,N_6055);
nand U7746 (N_7746,N_6640,N_6528);
nor U7747 (N_7747,N_5859,N_6740);
xor U7748 (N_7748,N_5853,N_7262);
and U7749 (N_7749,N_7158,N_6962);
nand U7750 (N_7750,N_5298,N_5898);
and U7751 (N_7751,N_5489,N_7072);
nand U7752 (N_7752,N_7213,N_6515);
and U7753 (N_7753,N_6978,N_5467);
xnor U7754 (N_7754,N_7463,N_7121);
nor U7755 (N_7755,N_6782,N_5386);
or U7756 (N_7756,N_6464,N_5789);
nor U7757 (N_7757,N_5202,N_7294);
or U7758 (N_7758,N_6700,N_5059);
nor U7759 (N_7759,N_6893,N_7297);
xor U7760 (N_7760,N_6633,N_5345);
and U7761 (N_7761,N_6230,N_7147);
and U7762 (N_7762,N_6444,N_5180);
nor U7763 (N_7763,N_6607,N_7432);
nor U7764 (N_7764,N_6275,N_5705);
nand U7765 (N_7765,N_6305,N_5096);
and U7766 (N_7766,N_5863,N_6665);
xor U7767 (N_7767,N_5823,N_6625);
nand U7768 (N_7768,N_5787,N_6974);
and U7769 (N_7769,N_5451,N_7005);
and U7770 (N_7770,N_7047,N_5331);
nor U7771 (N_7771,N_5114,N_5606);
nand U7772 (N_7772,N_5149,N_5272);
and U7773 (N_7773,N_6764,N_5612);
and U7774 (N_7774,N_6487,N_6569);
or U7775 (N_7775,N_6509,N_6252);
nand U7776 (N_7776,N_5291,N_5756);
nand U7777 (N_7777,N_5541,N_5592);
nand U7778 (N_7778,N_6505,N_7067);
or U7779 (N_7779,N_5038,N_6156);
nor U7780 (N_7780,N_6201,N_5670);
xnor U7781 (N_7781,N_7041,N_6189);
nor U7782 (N_7782,N_5834,N_5900);
and U7783 (N_7783,N_7356,N_5536);
or U7784 (N_7784,N_6102,N_5531);
nor U7785 (N_7785,N_7057,N_7079);
nand U7786 (N_7786,N_7174,N_6362);
nor U7787 (N_7787,N_6460,N_7419);
xor U7788 (N_7788,N_5936,N_6214);
or U7789 (N_7789,N_5432,N_5865);
and U7790 (N_7790,N_5977,N_5672);
nor U7791 (N_7791,N_6530,N_5799);
or U7792 (N_7792,N_7150,N_5037);
or U7793 (N_7793,N_6063,N_5363);
or U7794 (N_7794,N_6882,N_6389);
nand U7795 (N_7795,N_5335,N_6099);
nor U7796 (N_7796,N_5796,N_6100);
and U7797 (N_7797,N_6262,N_6558);
or U7798 (N_7798,N_6004,N_5380);
nand U7799 (N_7799,N_6957,N_5953);
xor U7800 (N_7800,N_6084,N_6393);
or U7801 (N_7801,N_6368,N_5079);
nand U7802 (N_7802,N_5957,N_5039);
nand U7803 (N_7803,N_7211,N_7340);
nor U7804 (N_7804,N_6029,N_7423);
nand U7805 (N_7805,N_6964,N_5282);
and U7806 (N_7806,N_5070,N_6906);
and U7807 (N_7807,N_5221,N_6043);
nand U7808 (N_7808,N_7083,N_5482);
or U7809 (N_7809,N_7288,N_5965);
and U7810 (N_7810,N_5158,N_5950);
nand U7811 (N_7811,N_6952,N_6721);
nand U7812 (N_7812,N_5299,N_5390);
and U7813 (N_7813,N_6926,N_7184);
xnor U7814 (N_7814,N_6802,N_7170);
and U7815 (N_7815,N_5741,N_7103);
nor U7816 (N_7816,N_6522,N_7465);
nand U7817 (N_7817,N_6841,N_5547);
and U7818 (N_7818,N_6728,N_6293);
nand U7819 (N_7819,N_6650,N_6399);
nand U7820 (N_7820,N_5523,N_5157);
nand U7821 (N_7821,N_6670,N_6236);
and U7822 (N_7822,N_5230,N_5813);
nand U7823 (N_7823,N_7127,N_6346);
nor U7824 (N_7824,N_6830,N_7286);
nand U7825 (N_7825,N_5348,N_5356);
or U7826 (N_7826,N_6525,N_6220);
and U7827 (N_7827,N_7175,N_6082);
nand U7828 (N_7828,N_5553,N_5018);
xor U7829 (N_7829,N_5665,N_6669);
nand U7830 (N_7830,N_6940,N_5469);
nor U7831 (N_7831,N_7236,N_6394);
nor U7832 (N_7832,N_6980,N_5117);
or U7833 (N_7833,N_6681,N_5248);
nand U7834 (N_7834,N_6232,N_7197);
nand U7835 (N_7835,N_6079,N_6887);
or U7836 (N_7836,N_5044,N_6320);
and U7837 (N_7837,N_6853,N_6463);
or U7838 (N_7838,N_5323,N_6860);
and U7839 (N_7839,N_6073,N_6663);
nand U7840 (N_7840,N_6575,N_6930);
and U7841 (N_7841,N_7241,N_5341);
nand U7842 (N_7842,N_6542,N_6058);
or U7843 (N_7843,N_6120,N_5894);
or U7844 (N_7844,N_5213,N_5695);
and U7845 (N_7845,N_5991,N_6924);
and U7846 (N_7846,N_5686,N_6046);
xor U7847 (N_7847,N_6645,N_5234);
and U7848 (N_7848,N_5058,N_7081);
nand U7849 (N_7849,N_5076,N_5811);
nor U7850 (N_7850,N_6735,N_7126);
or U7851 (N_7851,N_6908,N_7144);
or U7852 (N_7852,N_6117,N_6593);
or U7853 (N_7853,N_5336,N_5373);
nand U7854 (N_7854,N_5266,N_6186);
nor U7855 (N_7855,N_5109,N_6626);
and U7856 (N_7856,N_6693,N_7425);
or U7857 (N_7857,N_5684,N_5663);
nor U7858 (N_7858,N_5728,N_5203);
nand U7859 (N_7859,N_5344,N_7418);
nand U7860 (N_7860,N_5398,N_5669);
and U7861 (N_7861,N_7243,N_5253);
and U7862 (N_7862,N_7024,N_5951);
or U7863 (N_7863,N_5444,N_5654);
xnor U7864 (N_7864,N_5211,N_6648);
or U7865 (N_7865,N_7255,N_6182);
or U7866 (N_7866,N_6263,N_6808);
nor U7867 (N_7867,N_6538,N_6851);
nand U7868 (N_7868,N_6245,N_7112);
nor U7869 (N_7869,N_5388,N_7051);
and U7870 (N_7870,N_5637,N_7318);
nor U7871 (N_7871,N_6479,N_6941);
or U7872 (N_7872,N_5186,N_5218);
or U7873 (N_7873,N_6499,N_6240);
xnor U7874 (N_7874,N_7304,N_5880);
and U7875 (N_7875,N_5576,N_5946);
and U7876 (N_7876,N_6091,N_5718);
nor U7877 (N_7877,N_5145,N_5247);
or U7878 (N_7878,N_7468,N_6571);
or U7879 (N_7879,N_6567,N_5736);
nand U7880 (N_7880,N_6563,N_5150);
nor U7881 (N_7881,N_5516,N_6483);
nand U7882 (N_7882,N_5514,N_5493);
nand U7883 (N_7883,N_5861,N_7087);
xnor U7884 (N_7884,N_6672,N_5791);
nand U7885 (N_7885,N_6077,N_6459);
or U7886 (N_7886,N_7224,N_5024);
nand U7887 (N_7887,N_5983,N_6730);
or U7888 (N_7888,N_7040,N_5460);
nor U7889 (N_7889,N_5558,N_7203);
nor U7890 (N_7890,N_6244,N_6662);
nor U7891 (N_7891,N_6769,N_7323);
nor U7892 (N_7892,N_6771,N_6565);
or U7893 (N_7893,N_6095,N_6200);
and U7894 (N_7894,N_6801,N_5784);
nand U7895 (N_7895,N_5624,N_7022);
and U7896 (N_7896,N_5582,N_6496);
or U7897 (N_7897,N_6223,N_7173);
nand U7898 (N_7898,N_6018,N_6705);
nor U7899 (N_7899,N_5241,N_5485);
or U7900 (N_7900,N_6030,N_6160);
nor U7901 (N_7901,N_5902,N_5956);
and U7902 (N_7902,N_6532,N_6406);
nor U7903 (N_7903,N_5229,N_6400);
or U7904 (N_7904,N_5517,N_7367);
or U7905 (N_7905,N_7054,N_5754);
and U7906 (N_7906,N_7165,N_6578);
nor U7907 (N_7907,N_5581,N_5151);
and U7908 (N_7908,N_6707,N_6253);
and U7909 (N_7909,N_6468,N_5548);
or U7910 (N_7910,N_6191,N_6123);
or U7911 (N_7911,N_5873,N_5085);
or U7912 (N_7912,N_7095,N_7427);
and U7913 (N_7913,N_7410,N_6800);
xor U7914 (N_7914,N_5860,N_6457);
or U7915 (N_7915,N_6195,N_5584);
and U7916 (N_7916,N_6793,N_7442);
nor U7917 (N_7917,N_5103,N_6692);
nor U7918 (N_7918,N_5175,N_6909);
xnor U7919 (N_7919,N_7159,N_6914);
or U7920 (N_7920,N_6832,N_6242);
nor U7921 (N_7921,N_5786,N_6042);
and U7922 (N_7922,N_6145,N_7078);
or U7923 (N_7923,N_6198,N_5131);
and U7924 (N_7924,N_5462,N_6547);
or U7925 (N_7925,N_5715,N_5969);
nor U7926 (N_7926,N_5871,N_6478);
nand U7927 (N_7927,N_5989,N_7312);
xor U7928 (N_7928,N_6729,N_7388);
xnor U7929 (N_7929,N_5001,N_6572);
and U7930 (N_7930,N_6090,N_6115);
nand U7931 (N_7931,N_7456,N_6347);
xor U7932 (N_7932,N_7135,N_5979);
and U7933 (N_7933,N_5848,N_5325);
nor U7934 (N_7934,N_6759,N_5411);
nand U7935 (N_7935,N_6264,N_7480);
or U7936 (N_7936,N_6816,N_6387);
nor U7937 (N_7937,N_5375,N_6846);
nand U7938 (N_7938,N_6217,N_5570);
nand U7939 (N_7939,N_5135,N_5856);
or U7940 (N_7940,N_7097,N_5960);
and U7941 (N_7941,N_7252,N_5226);
nand U7942 (N_7942,N_7437,N_7296);
or U7943 (N_7943,N_6686,N_7244);
and U7944 (N_7944,N_7034,N_5094);
and U7945 (N_7945,N_6137,N_6491);
nand U7946 (N_7946,N_6276,N_6318);
xnor U7947 (N_7947,N_6657,N_6744);
nand U7948 (N_7948,N_6605,N_5463);
xor U7949 (N_7949,N_5961,N_6629);
or U7950 (N_7950,N_5337,N_6768);
or U7951 (N_7951,N_7138,N_5703);
or U7952 (N_7952,N_6641,N_5589);
or U7953 (N_7953,N_6557,N_6708);
and U7954 (N_7954,N_7328,N_6642);
nor U7955 (N_7955,N_6649,N_5342);
xnor U7956 (N_7956,N_6623,N_6574);
or U7957 (N_7957,N_5071,N_5437);
nand U7958 (N_7958,N_6162,N_5759);
or U7959 (N_7959,N_6282,N_6792);
and U7960 (N_7960,N_6112,N_5123);
and U7961 (N_7961,N_7245,N_6451);
and U7962 (N_7962,N_7063,N_7435);
nor U7963 (N_7963,N_5751,N_6702);
and U7964 (N_7964,N_5664,N_5723);
and U7965 (N_7965,N_7314,N_6856);
nor U7966 (N_7966,N_5958,N_5982);
or U7967 (N_7967,N_6448,N_6982);
and U7968 (N_7968,N_5724,N_5783);
nand U7969 (N_7969,N_7143,N_5433);
and U7970 (N_7970,N_5270,N_6848);
and U7971 (N_7971,N_7003,N_6098);
nand U7972 (N_7972,N_6550,N_7050);
nor U7973 (N_7973,N_6443,N_6210);
or U7974 (N_7974,N_6674,N_5692);
nor U7975 (N_7975,N_5938,N_6014);
and U7976 (N_7976,N_6196,N_6278);
and U7977 (N_7977,N_6903,N_5674);
nand U7978 (N_7978,N_6251,N_5532);
xnor U7979 (N_7979,N_5274,N_5505);
nand U7980 (N_7980,N_6752,N_6173);
nand U7981 (N_7981,N_7009,N_7382);
nor U7982 (N_7982,N_5761,N_5767);
nor U7983 (N_7983,N_5512,N_5625);
or U7984 (N_7984,N_5990,N_6606);
nor U7985 (N_7985,N_5330,N_5488);
nand U7986 (N_7986,N_7132,N_5618);
nand U7987 (N_7987,N_6986,N_6271);
nand U7988 (N_7988,N_5614,N_5693);
and U7989 (N_7989,N_7271,N_6933);
nand U7990 (N_7990,N_5002,N_5069);
or U7991 (N_7991,N_6402,N_6361);
nor U7992 (N_7992,N_6037,N_7441);
or U7993 (N_7993,N_7140,N_6993);
or U7994 (N_7994,N_7493,N_7330);
or U7995 (N_7995,N_6889,N_7086);
and U7996 (N_7996,N_6227,N_7494);
and U7997 (N_7997,N_6482,N_5877);
or U7998 (N_7998,N_7335,N_5792);
xor U7999 (N_7999,N_5243,N_7229);
nand U8000 (N_8000,N_5909,N_6603);
or U8001 (N_8001,N_6035,N_7353);
nand U8002 (N_8002,N_5825,N_7373);
nor U8003 (N_8003,N_5713,N_6776);
or U8004 (N_8004,N_6857,N_7091);
nand U8005 (N_8005,N_5034,N_5474);
nand U8006 (N_8006,N_6166,N_6925);
or U8007 (N_8007,N_5632,N_6631);
or U8008 (N_8008,N_6333,N_5190);
and U8009 (N_8009,N_5681,N_5238);
or U8010 (N_8010,N_7200,N_6143);
nor U8011 (N_8011,N_5095,N_7369);
nor U8012 (N_8012,N_5450,N_7210);
nand U8013 (N_8013,N_5017,N_6354);
and U8014 (N_8014,N_6103,N_5458);
nand U8015 (N_8015,N_5804,N_5984);
xnor U8016 (N_8016,N_5948,N_7026);
or U8017 (N_8017,N_6066,N_6534);
nor U8018 (N_8018,N_6111,N_5644);
nor U8019 (N_8019,N_7350,N_6668);
or U8020 (N_8020,N_7131,N_7333);
and U8021 (N_8021,N_5384,N_6009);
xnor U8022 (N_8022,N_7461,N_7077);
nor U8023 (N_8023,N_6806,N_7451);
or U8024 (N_8024,N_6019,N_5534);
nor U8025 (N_8025,N_5292,N_7055);
nand U8026 (N_8026,N_6507,N_5177);
nor U8027 (N_8027,N_6797,N_5003);
or U8028 (N_8028,N_5009,N_6418);
nand U8029 (N_8029,N_5568,N_5311);
xor U8030 (N_8030,N_5347,N_5594);
nand U8031 (N_8031,N_5524,N_7191);
nand U8032 (N_8032,N_7075,N_7386);
nor U8033 (N_8033,N_6791,N_5097);
or U8034 (N_8034,N_6291,N_5142);
or U8035 (N_8035,N_5515,N_6420);
nor U8036 (N_8036,N_5120,N_7364);
and U8037 (N_8037,N_6131,N_7088);
nand U8038 (N_8038,N_6359,N_6745);
nand U8039 (N_8039,N_6308,N_6873);
and U8040 (N_8040,N_7137,N_6081);
nor U8041 (N_8041,N_5016,N_7230);
nand U8042 (N_8042,N_5803,N_6374);
or U8043 (N_8043,N_6254,N_7292);
and U8044 (N_8044,N_7365,N_7017);
nor U8045 (N_8045,N_5418,N_6224);
nor U8046 (N_8046,N_5651,N_6326);
and U8047 (N_8047,N_6249,N_6694);
and U8048 (N_8048,N_5604,N_5235);
nor U8049 (N_8049,N_5326,N_6017);
nand U8050 (N_8050,N_6136,N_5197);
or U8051 (N_8051,N_7007,N_6330);
and U8052 (N_8052,N_6332,N_7338);
nor U8053 (N_8053,N_6519,N_5810);
xor U8054 (N_8054,N_6089,N_6126);
nand U8055 (N_8055,N_6949,N_6428);
and U8056 (N_8056,N_7157,N_7434);
nor U8057 (N_8057,N_6241,N_5395);
or U8058 (N_8058,N_5184,N_6340);
or U8059 (N_8059,N_6774,N_5974);
nor U8060 (N_8060,N_5376,N_7176);
and U8061 (N_8061,N_5305,N_6763);
or U8062 (N_8062,N_6379,N_5242);
or U8063 (N_8063,N_7139,N_5535);
or U8064 (N_8064,N_5591,N_6439);
and U8065 (N_8065,N_6785,N_5893);
or U8066 (N_8066,N_7422,N_6407);
nand U8067 (N_8067,N_6071,N_5312);
nor U8068 (N_8068,N_6283,N_5300);
and U8069 (N_8069,N_6977,N_7013);
nor U8070 (N_8070,N_5630,N_7336);
xnor U8071 (N_8071,N_5047,N_7227);
and U8072 (N_8072,N_7030,N_5304);
xnor U8073 (N_8073,N_5995,N_7119);
and U8074 (N_8074,N_5261,N_5588);
and U8075 (N_8075,N_6258,N_7357);
nand U8076 (N_8076,N_5448,N_5920);
nor U8077 (N_8077,N_6878,N_5025);
nor U8078 (N_8078,N_5178,N_5833);
nor U8079 (N_8079,N_6118,N_6840);
and U8080 (N_8080,N_5233,N_5441);
or U8081 (N_8081,N_5732,N_7421);
and U8082 (N_8082,N_5750,N_5749);
and U8083 (N_8083,N_5506,N_5052);
nor U8084 (N_8084,N_5354,N_7483);
and U8085 (N_8085,N_7202,N_5159);
and U8086 (N_8086,N_7080,N_6898);
nor U8087 (N_8087,N_6500,N_6433);
nand U8088 (N_8088,N_5425,N_6135);
and U8089 (N_8089,N_6167,N_7105);
or U8090 (N_8090,N_5209,N_7032);
or U8091 (N_8091,N_5768,N_6155);
nor U8092 (N_8092,N_6002,N_5704);
or U8093 (N_8093,N_6536,N_6959);
and U8094 (N_8094,N_6709,N_5181);
nor U8095 (N_8095,N_5262,N_5442);
and U8096 (N_8096,N_5381,N_7045);
and U8097 (N_8097,N_6762,N_6315);
nand U8098 (N_8098,N_5627,N_6553);
nor U8099 (N_8099,N_6829,N_6233);
xnor U8100 (N_8100,N_6711,N_6045);
or U8101 (N_8101,N_5607,N_6932);
nor U8102 (N_8102,N_6409,N_5636);
and U8103 (N_8103,N_7407,N_6116);
xor U8104 (N_8104,N_6331,N_6492);
nor U8105 (N_8105,N_5371,N_5317);
nand U8106 (N_8106,N_7374,N_5527);
xnor U8107 (N_8107,N_5954,N_5256);
and U8108 (N_8108,N_6988,N_6033);
nand U8109 (N_8109,N_5940,N_5701);
nand U8110 (N_8110,N_5760,N_7366);
nor U8111 (N_8111,N_6222,N_6734);
or U8112 (N_8112,N_5185,N_6273);
nor U8113 (N_8113,N_7104,N_6474);
and U8114 (N_8114,N_5540,N_5473);
nor U8115 (N_8115,N_7320,N_5350);
and U8116 (N_8116,N_6344,N_5198);
or U8117 (N_8117,N_7491,N_7098);
and U8118 (N_8118,N_7306,N_7311);
or U8119 (N_8119,N_7495,N_5296);
nor U8120 (N_8120,N_6312,N_5267);
and U8121 (N_8121,N_6834,N_5140);
or U8122 (N_8122,N_6267,N_5421);
and U8123 (N_8123,N_5562,N_6228);
nand U8124 (N_8124,N_6867,N_7413);
and U8125 (N_8125,N_5478,N_6715);
and U8126 (N_8126,N_6376,N_5250);
and U8127 (N_8127,N_6750,N_5911);
nand U8128 (N_8128,N_6864,N_5340);
or U8129 (N_8129,N_5522,N_5134);
nor U8130 (N_8130,N_6798,N_5042);
nor U8131 (N_8131,N_5981,N_6307);
and U8132 (N_8132,N_6582,N_6311);
nor U8133 (N_8133,N_7403,N_5945);
and U8134 (N_8134,N_5319,N_5508);
nand U8135 (N_8135,N_5800,N_6328);
nor U8136 (N_8136,N_5775,N_5967);
nand U8137 (N_8137,N_6027,N_5023);
or U8138 (N_8138,N_5641,N_7146);
or U8139 (N_8139,N_7129,N_6056);
nand U8140 (N_8140,N_7497,N_5831);
or U8141 (N_8141,N_7209,N_6591);
nor U8142 (N_8142,N_6013,N_5895);
nand U8143 (N_8143,N_6287,N_6329);
or U8144 (N_8144,N_7059,N_6783);
or U8145 (N_8145,N_6209,N_6599);
or U8146 (N_8146,N_7064,N_6527);
xor U8147 (N_8147,N_6134,N_5966);
or U8148 (N_8148,N_7372,N_7351);
xnor U8149 (N_8149,N_6176,N_5494);
and U8150 (N_8150,N_5928,N_5952);
or U8151 (N_8151,N_6905,N_6881);
or U8152 (N_8152,N_5276,N_5685);
nand U8153 (N_8153,N_5843,N_7109);
nor U8154 (N_8154,N_6861,N_6298);
xnor U8155 (N_8155,N_6388,N_7417);
nor U8156 (N_8156,N_7094,N_5525);
nand U8157 (N_8157,N_6288,N_7474);
or U8158 (N_8158,N_6367,N_6620);
and U8159 (N_8159,N_5587,N_7315);
or U8160 (N_8160,N_6297,N_5841);
nand U8161 (N_8161,N_5389,N_5986);
xnor U8162 (N_8162,N_5616,N_6199);
or U8163 (N_8163,N_5318,N_5526);
and U8164 (N_8164,N_5237,N_7308);
or U8165 (N_8165,N_5888,N_5600);
nor U8166 (N_8166,N_7044,N_5678);
nand U8167 (N_8167,N_7316,N_5931);
nand U8168 (N_8168,N_7385,N_6727);
xor U8169 (N_8169,N_6773,N_5817);
nor U8170 (N_8170,N_6699,N_6206);
and U8171 (N_8171,N_6758,N_6811);
nor U8172 (N_8172,N_5082,N_5826);
or U8173 (N_8173,N_6580,N_7089);
xor U8174 (N_8174,N_6843,N_5498);
and U8175 (N_8175,N_6461,N_6995);
nor U8176 (N_8176,N_6435,N_6655);
nor U8177 (N_8177,N_5490,N_5921);
nand U8178 (N_8178,N_6614,N_6380);
nor U8179 (N_8179,N_5402,N_5466);
nor U8180 (N_8180,N_7362,N_7000);
nand U8181 (N_8181,N_6050,N_5012);
and U8182 (N_8182,N_6895,N_7391);
nor U8183 (N_8183,N_6021,N_6392);
nand U8184 (N_8184,N_6208,N_6613);
nor U8185 (N_8185,N_5056,N_5146);
xnor U8186 (N_8186,N_5136,N_5797);
nand U8187 (N_8187,N_6833,N_5574);
xnor U8188 (N_8188,N_5286,N_6943);
xor U8189 (N_8189,N_6520,N_7025);
xor U8190 (N_8190,N_5821,N_6877);
nand U8191 (N_8191,N_6024,N_5436);
nand U8192 (N_8192,N_5088,N_6579);
or U8193 (N_8193,N_7148,N_6621);
nor U8194 (N_8194,N_7279,N_6085);
or U8195 (N_8195,N_7027,N_7290);
or U8196 (N_8196,N_5901,N_6677);
and U8197 (N_8197,N_7379,N_6415);
nand U8198 (N_8198,N_6916,N_7208);
xor U8199 (N_8199,N_7195,N_6503);
or U8200 (N_8200,N_6324,N_6325);
nand U8201 (N_8201,N_7193,N_7475);
nor U8202 (N_8202,N_7008,N_6907);
nand U8203 (N_8203,N_6290,N_5887);
nor U8204 (N_8204,N_7444,N_5549);
and U8205 (N_8205,N_5696,N_5934);
xnor U8206 (N_8206,N_5816,N_6598);
xor U8207 (N_8207,N_5908,N_7111);
nor U8208 (N_8208,N_6432,N_6552);
xnor U8209 (N_8209,N_5382,N_6484);
nor U8210 (N_8210,N_7226,N_6097);
nand U8211 (N_8211,N_6257,N_7020);
and U8212 (N_8212,N_5457,N_5249);
nand U8213 (N_8213,N_6888,N_5566);
nand U8214 (N_8214,N_5798,N_6405);
nand U8215 (N_8215,N_6979,N_7363);
nor U8216 (N_8216,N_5742,N_7160);
nand U8217 (N_8217,N_6619,N_7334);
xor U8218 (N_8218,N_5141,N_6944);
nor U8219 (N_8219,N_5782,N_5443);
nor U8220 (N_8220,N_6586,N_5329);
and U8221 (N_8221,N_6360,N_7358);
or U8222 (N_8222,N_5366,N_6171);
and U8223 (N_8223,N_5167,N_5730);
or U8224 (N_8224,N_5781,N_6927);
nand U8225 (N_8225,N_6996,N_7360);
nand U8226 (N_8226,N_6577,N_5518);
or U8227 (N_8227,N_7149,N_5208);
nand U8228 (N_8228,N_5414,N_6011);
and U8229 (N_8229,N_6576,N_5275);
nor U8230 (N_8230,N_6234,N_5520);
nor U8231 (N_8231,N_6842,N_7246);
nor U8232 (N_8232,N_5778,N_5501);
and U8233 (N_8233,N_6733,N_6343);
xor U8234 (N_8234,N_6755,N_5890);
or U8235 (N_8235,N_6966,N_6044);
and U8236 (N_8236,N_5912,N_6248);
and U8237 (N_8237,N_5802,N_6754);
nand U8238 (N_8238,N_5010,N_6076);
or U8239 (N_8239,N_6277,N_5619);
and U8240 (N_8240,N_5780,N_5533);
nor U8241 (N_8241,N_5420,N_7499);
and U8242 (N_8242,N_6920,N_6756);
nor U8243 (N_8243,N_5976,N_7389);
nand U8244 (N_8244,N_7242,N_6153);
nand U8245 (N_8245,N_5923,N_6584);
nand U8246 (N_8246,N_5544,N_6070);
xor U8247 (N_8247,N_7082,N_5925);
and U8248 (N_8248,N_6034,N_7354);
or U8249 (N_8249,N_6911,N_5297);
nor U8250 (N_8250,N_6876,N_7116);
nand U8251 (N_8251,N_7397,N_5019);
nor U8252 (N_8252,N_5788,N_7496);
nand U8253 (N_8253,N_6656,N_5091);
nor U8254 (N_8254,N_6880,N_5580);
nand U8255 (N_8255,N_5309,N_7212);
and U8256 (N_8256,N_6615,N_5424);
or U8257 (N_8257,N_5343,N_6637);
and U8258 (N_8258,N_5471,N_5065);
or U8259 (N_8259,N_6818,N_5640);
nand U8260 (N_8260,N_6991,N_5687);
nand U8261 (N_8261,N_7093,N_5631);
nor U8262 (N_8262,N_5406,N_7180);
nand U8263 (N_8263,N_7305,N_6447);
and U8264 (N_8264,N_7458,N_5321);
or U8265 (N_8265,N_5708,N_5086);
nor U8266 (N_8266,N_5537,N_5456);
or U8267 (N_8267,N_6879,N_7118);
nand U8268 (N_8268,N_5359,N_5737);
nand U8269 (N_8269,N_7455,N_7447);
and U8270 (N_8270,N_5680,N_7043);
and U8271 (N_8271,N_6506,N_5073);
nand U8272 (N_8272,N_6161,N_5244);
and U8273 (N_8273,N_6976,N_6508);
or U8274 (N_8274,N_6765,N_6921);
or U8275 (N_8275,N_5116,N_7457);
xor U8276 (N_8276,N_5405,N_5215);
nand U8277 (N_8277,N_5057,N_6784);
and U8278 (N_8278,N_5351,N_5567);
and U8279 (N_8279,N_5850,N_6455);
or U8280 (N_8280,N_5658,N_6177);
nor U8281 (N_8281,N_5223,N_5092);
nor U8282 (N_8282,N_5115,N_6353);
nor U8283 (N_8283,N_6770,N_7182);
and U8284 (N_8284,N_6671,N_6356);
nor U8285 (N_8285,N_6202,N_5937);
nand U8286 (N_8286,N_5004,N_5926);
or U8287 (N_8287,N_5365,N_5176);
or U8288 (N_8288,N_7277,N_5929);
or U8289 (N_8289,N_6450,N_5870);
nor U8290 (N_8290,N_5874,N_5408);
nand U8291 (N_8291,N_6514,N_6912);
nand U8292 (N_8292,N_6062,N_5623);
or U8293 (N_8293,N_6872,N_5722);
xor U8294 (N_8294,N_6989,N_5013);
and U8295 (N_8295,N_7253,N_6931);
and U8296 (N_8296,N_5475,N_5858);
nand U8297 (N_8297,N_6647,N_6188);
and U8298 (N_8298,N_7107,N_7409);
nand U8299 (N_8299,N_5212,N_6583);
nand U8300 (N_8300,N_7201,N_6309);
or U8301 (N_8301,N_6545,N_5846);
nand U8302 (N_8302,N_7313,N_6313);
nor U8303 (N_8303,N_7298,N_5435);
nor U8304 (N_8304,N_5121,N_6609);
nor U8305 (N_8305,N_7301,N_5383);
and U8306 (N_8306,N_5391,N_6929);
nor U8307 (N_8307,N_6436,N_6736);
and U8308 (N_8308,N_5530,N_5824);
nor U8309 (N_8309,N_7469,N_6900);
nor U8310 (N_8310,N_5280,N_5962);
xnor U8311 (N_8311,N_6742,N_6718);
nor U8312 (N_8312,N_5899,N_6336);
and U8313 (N_8313,N_5978,N_5653);
and U8314 (N_8314,N_6973,N_5806);
or U8315 (N_8315,N_6007,N_7378);
nand U8316 (N_8316,N_5108,N_7076);
nor U8317 (N_8317,N_5812,N_6595);
nand U8318 (N_8318,N_6383,N_6250);
nor U8319 (N_8319,N_7048,N_6395);
nand U8320 (N_8320,N_7317,N_6859);
xor U8321 (N_8321,N_5727,N_7408);
or U8322 (N_8322,N_7033,N_5449);
nand U8323 (N_8323,N_5284,N_6083);
nand U8324 (N_8324,N_5080,N_6883);
or U8325 (N_8325,N_5205,N_6696);
nor U8326 (N_8326,N_7004,N_7221);
nor U8327 (N_8327,N_6948,N_6799);
and U8328 (N_8328,N_5125,N_7194);
nand U8329 (N_8329,N_6052,N_6181);
or U8330 (N_8330,N_6138,N_7394);
nand U8331 (N_8331,N_5028,N_5122);
nor U8332 (N_8332,N_5106,N_6417);
xnor U8333 (N_8333,N_5294,N_7341);
and U8334 (N_8334,N_6023,N_5910);
nor U8335 (N_8335,N_5048,N_7196);
nor U8336 (N_8336,N_5401,N_5277);
and U8337 (N_8337,N_5661,N_5020);
or U8338 (N_8338,N_5179,N_6826);
or U8339 (N_8339,N_5196,N_7185);
nand U8340 (N_8340,N_5652,N_6928);
or U8341 (N_8341,N_7399,N_6335);
or U8342 (N_8342,N_6805,N_7134);
nand U8343 (N_8343,N_7240,N_6923);
or U8344 (N_8344,N_5521,N_6703);
and U8345 (N_8345,N_5699,N_7062);
xor U8346 (N_8346,N_6942,N_6471);
nor U8347 (N_8347,N_5500,N_5716);
and U8348 (N_8348,N_5081,N_6106);
nor U8349 (N_8349,N_6981,N_6890);
or U8350 (N_8350,N_5886,N_5676);
and U8351 (N_8351,N_5822,N_6884);
or U8352 (N_8352,N_5219,N_5074);
or U8353 (N_8353,N_6281,N_6437);
or U8354 (N_8354,N_7346,N_5295);
and U8355 (N_8355,N_5355,N_5251);
and U8356 (N_8356,N_7400,N_6561);
or U8357 (N_8357,N_5217,N_5885);
nor U8358 (N_8358,N_7084,N_7345);
nand U8359 (N_8359,N_7449,N_5917);
nand U8360 (N_8360,N_7169,N_7416);
nor U8361 (N_8361,N_5132,N_7460);
or U8362 (N_8362,N_7404,N_6684);
nand U8363 (N_8363,N_5513,N_6119);
nand U8364 (N_8364,N_5545,N_6403);
xor U8365 (N_8365,N_6611,N_7361);
and U8366 (N_8366,N_6197,N_6753);
nor U8367 (N_8367,N_5726,N_7188);
and U8368 (N_8368,N_5656,N_5763);
nor U8369 (N_8369,N_5711,N_5153);
and U8370 (N_8370,N_5815,N_5862);
and U8371 (N_8371,N_7058,N_6092);
and U8372 (N_8372,N_5611,N_6292);
or U8373 (N_8373,N_7110,N_6404);
nand U8374 (N_8374,N_6279,N_5431);
xor U8375 (N_8375,N_7443,N_7238);
nor U8376 (N_8376,N_7035,N_6559);
nor U8377 (N_8377,N_6587,N_5477);
or U8378 (N_8378,N_6726,N_7215);
and U8379 (N_8379,N_7284,N_6109);
and U8380 (N_8380,N_5930,N_6870);
nor U8381 (N_8381,N_5565,N_5595);
or U8382 (N_8382,N_7348,N_6255);
xnor U8383 (N_8383,N_6316,N_5128);
or U8384 (N_8384,N_5195,N_6523);
or U8385 (N_8385,N_6168,N_5089);
and U8386 (N_8386,N_5554,N_5000);
xnor U8387 (N_8387,N_6968,N_6673);
or U8388 (N_8388,N_6036,N_6804);
and U8389 (N_8389,N_7327,N_7016);
and U8390 (N_8390,N_6147,N_5173);
xor U8391 (N_8391,N_5992,N_5164);
nand U8392 (N_8392,N_5483,N_5051);
or U8393 (N_8393,N_6581,N_6301);
nor U8394 (N_8394,N_6010,N_6537);
nand U8395 (N_8395,N_6001,N_6632);
and U8396 (N_8396,N_5891,N_5700);
xnor U8397 (N_8397,N_5083,N_6624);
or U8398 (N_8398,N_6967,N_7433);
nor U8399 (N_8399,N_6810,N_6902);
and U8400 (N_8400,N_5608,N_6341);
xnor U8401 (N_8401,N_6757,N_6006);
and U8402 (N_8402,N_6185,N_5399);
or U8403 (N_8403,N_5026,N_5171);
and U8404 (N_8404,N_5776,N_5702);
and U8405 (N_8405,N_5794,N_6113);
nand U8406 (N_8406,N_6939,N_6413);
and U8407 (N_8407,N_6517,N_6373);
and U8408 (N_8408,N_5897,N_5470);
or U8409 (N_8409,N_6477,N_5204);
or U8410 (N_8410,N_6731,N_6634);
nor U8411 (N_8411,N_6886,N_6521);
or U8412 (N_8412,N_6714,N_6749);
and U8413 (N_8413,N_6067,N_6094);
or U8414 (N_8414,N_6125,N_7163);
and U8415 (N_8415,N_6827,N_7339);
or U8416 (N_8416,N_5959,N_7466);
xor U8417 (N_8417,N_6636,N_6938);
or U8418 (N_8418,N_5293,N_5933);
nor U8419 (N_8419,N_7309,N_7038);
or U8420 (N_8420,N_6862,N_5743);
nand U8421 (N_8421,N_5947,N_5849);
nand U8422 (N_8422,N_7414,N_5055);
and U8423 (N_8423,N_6401,N_6486);
or U8424 (N_8424,N_6999,N_5216);
or U8425 (N_8425,N_7264,N_7018);
and U8426 (N_8426,N_7070,N_5852);
and U8427 (N_8427,N_6812,N_7155);
nand U8428 (N_8428,N_6751,N_5022);
nor U8429 (N_8429,N_5006,N_6365);
nor U8430 (N_8430,N_7331,N_6717);
or U8431 (N_8431,N_5324,N_6170);
and U8432 (N_8432,N_5387,N_5916);
nor U8433 (N_8433,N_5519,N_6675);
and U8434 (N_8434,N_6243,N_6124);
or U8435 (N_8435,N_7482,N_7028);
or U8436 (N_8436,N_5867,N_7060);
and U8437 (N_8437,N_5239,N_7488);
or U8438 (N_8438,N_6080,N_5642);
nor U8439 (N_8439,N_7219,N_7448);
and U8440 (N_8440,N_7387,N_6956);
nand U8441 (N_8441,N_5263,N_6059);
nor U8442 (N_8442,N_5502,N_6039);
or U8443 (N_8443,N_7235,N_7344);
and U8444 (N_8444,N_7177,N_6678);
nand U8445 (N_8445,N_5160,N_7411);
xnor U8446 (N_8446,N_5795,N_5206);
xor U8447 (N_8447,N_5528,N_6087);
nor U8448 (N_8448,N_6781,N_5271);
nand U8449 (N_8449,N_6676,N_5621);
or U8450 (N_8450,N_5285,N_5550);
nor U8451 (N_8451,N_6445,N_5932);
nor U8452 (N_8452,N_6616,N_5939);
or U8453 (N_8453,N_7090,N_7228);
or U8454 (N_8454,N_6701,N_7477);
nand U8455 (N_8455,N_5154,N_5993);
and U8456 (N_8456,N_7106,N_6594);
or U8457 (N_8457,N_5049,N_5710);
or U8458 (N_8458,N_5110,N_6272);
or U8459 (N_8459,N_5161,N_6789);
nor U8460 (N_8460,N_5360,N_5133);
or U8461 (N_8461,N_5635,N_7234);
nor U8462 (N_8462,N_5377,N_6743);
and U8463 (N_8463,N_5682,N_6414);
or U8464 (N_8464,N_6016,N_7479);
and U8465 (N_8465,N_7010,N_5721);
xor U8466 (N_8466,N_5035,N_5904);
nor U8467 (N_8467,N_5200,N_6600);
nand U8468 (N_8468,N_5552,N_7172);
xnor U8469 (N_8469,N_6003,N_6885);
or U8470 (N_8470,N_6040,N_5379);
and U8471 (N_8471,N_5084,N_5762);
nor U8472 (N_8472,N_5166,N_5454);
xnor U8473 (N_8473,N_6918,N_5062);
xnor U8474 (N_8474,N_5771,N_6020);
nor U8475 (N_8475,N_6342,N_6480);
xor U8476 (N_8476,N_7049,N_6719);
or U8477 (N_8477,N_6622,N_5268);
nand U8478 (N_8478,N_5790,N_6294);
nor U8479 (N_8479,N_6053,N_5349);
nand U8480 (N_8480,N_5105,N_5455);
nand U8481 (N_8481,N_5265,N_6838);
nor U8482 (N_8482,N_7326,N_7453);
nand U8483 (N_8483,N_7405,N_5543);
and U8484 (N_8484,N_7218,N_6183);
and U8485 (N_8485,N_5429,N_7198);
or U8486 (N_8486,N_7307,N_6154);
nor U8487 (N_8487,N_6712,N_6850);
nor U8488 (N_8488,N_6302,N_7164);
nand U8489 (N_8489,N_6690,N_5428);
nand U8490 (N_8490,N_6779,N_6355);
nor U8491 (N_8491,N_6858,N_5731);
xnor U8492 (N_8492,N_5679,N_6874);
or U8493 (N_8493,N_6683,N_6660);
xnor U8494 (N_8494,N_6852,N_7481);
nand U8495 (N_8495,N_6416,N_5367);
or U8496 (N_8496,N_7321,N_6524);
nor U8497 (N_8497,N_7489,N_7359);
or U8498 (N_8498,N_6221,N_5066);
nor U8499 (N_8499,N_6306,N_5029);
nand U8500 (N_8500,N_6865,N_7179);
or U8501 (N_8501,N_5561,N_5999);
or U8502 (N_8502,N_5633,N_6969);
nor U8503 (N_8503,N_6958,N_7452);
nor U8504 (N_8504,N_7056,N_5915);
nand U8505 (N_8505,N_6421,N_6121);
nor U8506 (N_8506,N_6323,N_5072);
nor U8507 (N_8507,N_5733,N_5615);
or U8508 (N_8508,N_7319,N_7355);
nand U8509 (N_8509,N_5100,N_6945);
nand U8510 (N_8510,N_5144,N_5155);
and U8511 (N_8511,N_5739,N_5814);
and U8512 (N_8512,N_6215,N_6518);
and U8513 (N_8513,N_6133,N_6725);
xnor U8514 (N_8514,N_7384,N_5045);
nor U8515 (N_8515,N_5119,N_5459);
nand U8516 (N_8516,N_7396,N_5245);
nand U8517 (N_8517,N_6350,N_5102);
and U8518 (N_8518,N_7295,N_6476);
and U8519 (N_8519,N_5077,N_6381);
nor U8520 (N_8520,N_7207,N_5394);
nor U8521 (N_8521,N_7133,N_7122);
and U8522 (N_8522,N_6602,N_5227);
xnor U8523 (N_8523,N_6766,N_5896);
nand U8524 (N_8524,N_6814,N_6216);
and U8525 (N_8525,N_6809,N_6639);
nor U8526 (N_8526,N_5854,N_5830);
or U8527 (N_8527,N_5996,N_6984);
xnor U8528 (N_8528,N_5662,N_5101);
xor U8529 (N_8529,N_5578,N_6449);
nand U8530 (N_8530,N_6685,N_6349);
and U8531 (N_8531,N_6777,N_6107);
and U8532 (N_8532,N_5130,N_5422);
nand U8533 (N_8533,N_5660,N_6951);
and U8534 (N_8534,N_5403,N_5228);
xor U8535 (N_8535,N_5137,N_6748);
and U8536 (N_8536,N_5465,N_7324);
or U8537 (N_8537,N_7310,N_7101);
or U8538 (N_8538,N_6317,N_5479);
and U8539 (N_8539,N_6556,N_6790);
or U8540 (N_8540,N_5273,N_5855);
or U8541 (N_8541,N_6831,N_7402);
and U8542 (N_8542,N_7258,N_6048);
or U8543 (N_8543,N_6110,N_5288);
nand U8544 (N_8544,N_6915,N_6564);
nor U8545 (N_8545,N_7145,N_7166);
or U8546 (N_8546,N_5744,N_6747);
nor U8547 (N_8547,N_5551,N_6440);
and U8548 (N_8548,N_6194,N_6998);
nor U8549 (N_8549,N_7250,N_7249);
nand U8550 (N_8550,N_5610,N_5495);
nor U8551 (N_8551,N_6159,N_7152);
xor U8552 (N_8552,N_7269,N_5078);
nand U8553 (N_8553,N_5765,N_6141);
nand U8554 (N_8554,N_5194,N_6987);
nor U8555 (N_8555,N_6548,N_5838);
and U8556 (N_8556,N_6512,N_6015);
nor U8557 (N_8557,N_7156,N_6151);
and U8558 (N_8558,N_7445,N_5579);
or U8559 (N_8559,N_6375,N_5883);
and U8560 (N_8560,N_7021,N_5364);
nor U8561 (N_8561,N_7168,N_5809);
and U8562 (N_8562,N_7012,N_5542);
or U8563 (N_8563,N_6472,N_7289);
nand U8564 (N_8564,N_5067,N_6761);
and U8565 (N_8565,N_5689,N_6065);
or U8566 (N_8566,N_6821,N_7153);
and U8567 (N_8567,N_5569,N_5075);
or U8568 (N_8568,N_6430,N_5370);
or U8569 (N_8569,N_6470,N_6994);
nand U8570 (N_8570,N_5709,N_6164);
xnor U8571 (N_8571,N_5053,N_6778);
or U8572 (N_8572,N_5628,N_6122);
xnor U8573 (N_8573,N_6825,N_5829);
and U8574 (N_8574,N_7412,N_6467);
xor U8575 (N_8575,N_5246,N_5879);
and U8576 (N_8576,N_6822,N_7247);
and U8577 (N_8577,N_6423,N_6469);
xor U8578 (N_8578,N_5254,N_5510);
or U8579 (N_8579,N_5922,N_6983);
and U8580 (N_8580,N_5168,N_6543);
or U8581 (N_8581,N_7380,N_7096);
and U8582 (N_8582,N_6163,N_5126);
nor U8583 (N_8583,N_7014,N_5087);
and U8584 (N_8584,N_6667,N_5869);
nor U8585 (N_8585,N_5769,N_5572);
nor U8586 (N_8586,N_5054,N_5484);
or U8587 (N_8587,N_6427,N_7068);
and U8588 (N_8588,N_5163,N_6338);
and U8589 (N_8589,N_6780,N_5339);
or U8590 (N_8590,N_6732,N_6390);
nor U8591 (N_8591,N_5807,N_7130);
nor U8592 (N_8592,N_6489,N_5770);
xnor U8593 (N_8593,N_6246,N_6108);
nor U8594 (N_8594,N_7231,N_7199);
nor U8595 (N_8595,N_6511,N_6152);
nor U8596 (N_8596,N_7011,N_5030);
nand U8597 (N_8597,N_5819,N_6697);
xnor U8598 (N_8598,N_7031,N_7239);
or U8599 (N_8599,N_6146,N_6130);
xnor U8600 (N_8600,N_6871,N_5963);
or U8601 (N_8601,N_6502,N_6456);
and U8602 (N_8602,N_5622,N_6370);
xnor U8603 (N_8603,N_6481,N_6386);
nor U8604 (N_8604,N_6950,N_5955);
or U8605 (N_8605,N_6008,N_6266);
or U8606 (N_8606,N_5222,N_5673);
or U8607 (N_8607,N_6786,N_7376);
or U8608 (N_8608,N_5313,N_5099);
nand U8609 (N_8609,N_5832,N_6836);
nand U8610 (N_8610,N_5719,N_6069);
nor U8611 (N_8611,N_6824,N_6256);
and U8612 (N_8612,N_5638,N_7237);
nand U8613 (N_8613,N_5308,N_5316);
xor U8614 (N_8614,N_5599,N_6985);
nand U8615 (N_8615,N_5889,N_5111);
nand U8616 (N_8616,N_7420,N_5844);
nand U8617 (N_8617,N_6101,N_5129);
nor U8618 (N_8618,N_7029,N_7125);
or U8619 (N_8619,N_5357,N_6235);
nand U8620 (N_8620,N_7248,N_6327);
or U8621 (N_8621,N_6226,N_5980);
nand U8622 (N_8622,N_7446,N_5393);
nor U8623 (N_8623,N_6627,N_7424);
or U8624 (N_8624,N_6012,N_7036);
or U8625 (N_8625,N_6139,N_5837);
nand U8626 (N_8626,N_5021,N_6854);
nor U8627 (N_8627,N_6207,N_5279);
xnor U8628 (N_8628,N_7270,N_6947);
or U8629 (N_8629,N_5666,N_7426);
nand U8630 (N_8630,N_6369,N_6148);
and U8631 (N_8631,N_6960,N_7223);
nor U8632 (N_8632,N_6844,N_5747);
nor U8633 (N_8633,N_5231,N_5649);
and U8634 (N_8634,N_6601,N_7136);
and U8635 (N_8635,N_7205,N_6990);
nand U8636 (N_8636,N_6270,N_6839);
and U8637 (N_8637,N_6597,N_7377);
nand U8638 (N_8638,N_6473,N_6796);
and U8639 (N_8639,N_6363,N_5648);
or U8640 (N_8640,N_6592,N_5725);
nand U8641 (N_8641,N_6516,N_6411);
nand U8642 (N_8642,N_5041,N_6688);
xor U8643 (N_8643,N_6231,N_6658);
nand U8644 (N_8644,N_6371,N_5918);
nor U8645 (N_8645,N_5655,N_5801);
nor U8646 (N_8646,N_7265,N_6820);
and U8647 (N_8647,N_6541,N_5694);
nor U8648 (N_8648,N_6664,N_6922);
nor U8649 (N_8649,N_5328,N_6661);
nand U8650 (N_8650,N_5927,N_6875);
and U8651 (N_8651,N_5677,N_7439);
nand U8652 (N_8652,N_5302,N_5773);
nor U8653 (N_8653,N_5461,N_5820);
nand U8654 (N_8654,N_5050,N_5192);
or U8655 (N_8655,N_6551,N_7440);
or U8656 (N_8656,N_5434,N_6174);
xnor U8657 (N_8657,N_6286,N_7349);
or U8658 (N_8658,N_6104,N_6970);
and U8659 (N_8659,N_6378,N_5264);
nor U8660 (N_8660,N_5603,N_5396);
and U8661 (N_8661,N_7263,N_6205);
nand U8662 (N_8662,N_6321,N_5352);
nor U8663 (N_8663,N_5174,N_6372);
nand U8664 (N_8664,N_5997,N_6695);
nand U8665 (N_8665,N_6710,N_6687);
xor U8666 (N_8666,N_7438,N_5714);
nor U8667 (N_8667,N_5064,N_6114);
nand U8668 (N_8668,N_5504,N_7186);
or U8669 (N_8669,N_5440,N_5201);
nor U8670 (N_8670,N_5327,N_7192);
nor U8671 (N_8671,N_5011,N_5480);
nand U8672 (N_8672,N_5590,N_5596);
nand U8673 (N_8673,N_6213,N_5301);
xnor U8674 (N_8674,N_5152,N_5090);
nand U8675 (N_8675,N_7282,N_7073);
nand U8676 (N_8676,N_6485,N_6698);
nand U8677 (N_8677,N_5836,N_5755);
nor U8678 (N_8678,N_6031,N_6585);
xor U8679 (N_8679,N_6608,N_5971);
nand U8680 (N_8680,N_7102,N_5866);
and U8681 (N_8681,N_7371,N_5290);
or U8682 (N_8682,N_6304,N_7291);
or U8683 (N_8683,N_7114,N_6767);
nor U8684 (N_8684,N_6310,N_5098);
nor U8685 (N_8685,N_7398,N_6526);
or U8686 (N_8686,N_6391,N_6269);
xor U8687 (N_8687,N_6972,N_5334);
nand U8688 (N_8688,N_6604,N_6910);
xor U8689 (N_8689,N_7257,N_7275);
and U8690 (N_8690,N_7485,N_5378);
or U8691 (N_8691,N_7464,N_5559);
nand U8692 (N_8692,N_5994,N_5872);
or U8693 (N_8693,N_7492,N_5643);
or U8694 (N_8694,N_7268,N_5868);
or U8695 (N_8695,N_6946,N_6992);
xnor U8696 (N_8696,N_6961,N_7395);
and U8697 (N_8697,N_7273,N_5746);
nor U8698 (N_8698,N_5499,N_5040);
nor U8699 (N_8699,N_5659,N_5156);
nand U8700 (N_8700,N_6775,N_5369);
or U8701 (N_8701,N_5942,N_6093);
and U8702 (N_8702,N_5509,N_5015);
or U8703 (N_8703,N_5320,N_5220);
or U8704 (N_8704,N_5033,N_6219);
nor U8705 (N_8705,N_5907,N_6490);
xnor U8706 (N_8706,N_7052,N_6064);
xor U8707 (N_8707,N_7233,N_6540);
and U8708 (N_8708,N_6892,N_5138);
or U8709 (N_8709,N_6919,N_6047);
nand U8710 (N_8710,N_6385,N_5445);
nand U8711 (N_8711,N_5557,N_6303);
nand U8712 (N_8712,N_5757,N_5236);
and U8713 (N_8713,N_5476,N_5281);
nand U8714 (N_8714,N_7217,N_6074);
nor U8715 (N_8715,N_7498,N_7216);
and U8716 (N_8716,N_5987,N_6596);
and U8717 (N_8717,N_7251,N_7108);
and U8718 (N_8718,N_5093,N_6211);
xor U8719 (N_8719,N_5046,N_6535);
nand U8720 (N_8720,N_6157,N_5818);
and U8721 (N_8721,N_7431,N_5988);
or U8722 (N_8722,N_5586,N_7187);
nand U8723 (N_8723,N_5943,N_5546);
or U8724 (N_8724,N_6612,N_6260);
xor U8725 (N_8725,N_7322,N_5240);
nor U8726 (N_8726,N_6863,N_5289);
nor U8727 (N_8727,N_5338,N_5333);
nand U8728 (N_8728,N_5407,N_5748);
nand U8729 (N_8729,N_5368,N_7285);
and U8730 (N_8730,N_7006,N_7214);
nand U8731 (N_8731,N_6072,N_7100);
xor U8732 (N_8732,N_7459,N_6184);
and U8733 (N_8733,N_6096,N_7472);
nand U8734 (N_8734,N_5857,N_5107);
and U8735 (N_8735,N_5875,N_5061);
nor U8736 (N_8736,N_6510,N_6284);
and U8737 (N_8737,N_5415,N_5973);
nor U8738 (N_8738,N_6274,N_7274);
or U8739 (N_8739,N_6546,N_7085);
nor U8740 (N_8740,N_7019,N_5712);
nor U8741 (N_8741,N_7002,N_5409);
xor U8742 (N_8742,N_6357,N_6041);
nor U8743 (N_8743,N_5626,N_5310);
nand U8744 (N_8744,N_5255,N_6280);
and U8745 (N_8745,N_5410,N_5905);
and U8746 (N_8746,N_5949,N_6203);
nor U8747 (N_8747,N_5008,N_6172);
nor U8748 (N_8748,N_6720,N_6823);
nand U8749 (N_8749,N_5924,N_6218);
and U8750 (N_8750,N_7154,N_5785);
nor U8751 (N_8751,N_6103,N_7311);
nand U8752 (N_8752,N_5776,N_5751);
or U8753 (N_8753,N_7327,N_7289);
or U8754 (N_8754,N_6707,N_7145);
nor U8755 (N_8755,N_5387,N_5337);
nor U8756 (N_8756,N_6514,N_6192);
nor U8757 (N_8757,N_5494,N_6553);
nor U8758 (N_8758,N_5819,N_5983);
nor U8759 (N_8759,N_7475,N_6646);
nor U8760 (N_8760,N_5318,N_6863);
or U8761 (N_8761,N_6060,N_5179);
xnor U8762 (N_8762,N_5349,N_5229);
and U8763 (N_8763,N_7243,N_6868);
or U8764 (N_8764,N_6403,N_6339);
nor U8765 (N_8765,N_5694,N_6764);
or U8766 (N_8766,N_5921,N_6337);
and U8767 (N_8767,N_7153,N_5439);
and U8768 (N_8768,N_5669,N_5130);
or U8769 (N_8769,N_7202,N_6554);
nor U8770 (N_8770,N_5702,N_6610);
or U8771 (N_8771,N_6782,N_6519);
or U8772 (N_8772,N_6848,N_5984);
and U8773 (N_8773,N_6822,N_5319);
and U8774 (N_8774,N_6004,N_6885);
nor U8775 (N_8775,N_7221,N_6511);
and U8776 (N_8776,N_6458,N_6405);
or U8777 (N_8777,N_6345,N_6461);
nand U8778 (N_8778,N_6933,N_6187);
or U8779 (N_8779,N_5307,N_5832);
xnor U8780 (N_8780,N_5918,N_6817);
and U8781 (N_8781,N_5217,N_7006);
nor U8782 (N_8782,N_5569,N_6385);
xor U8783 (N_8783,N_6028,N_6985);
and U8784 (N_8784,N_5334,N_5832);
nor U8785 (N_8785,N_5401,N_6675);
nor U8786 (N_8786,N_5759,N_5052);
and U8787 (N_8787,N_5313,N_5820);
nor U8788 (N_8788,N_5663,N_5551);
and U8789 (N_8789,N_5415,N_5439);
and U8790 (N_8790,N_5821,N_5252);
and U8791 (N_8791,N_5353,N_5380);
xor U8792 (N_8792,N_6221,N_6794);
and U8793 (N_8793,N_7420,N_7490);
or U8794 (N_8794,N_5414,N_5086);
and U8795 (N_8795,N_5332,N_5314);
nor U8796 (N_8796,N_5987,N_7027);
or U8797 (N_8797,N_5889,N_6747);
nand U8798 (N_8798,N_5911,N_7236);
nor U8799 (N_8799,N_5487,N_6975);
and U8800 (N_8800,N_5424,N_6011);
xor U8801 (N_8801,N_6606,N_6822);
nand U8802 (N_8802,N_6079,N_6019);
and U8803 (N_8803,N_6575,N_6881);
nand U8804 (N_8804,N_5909,N_7018);
nor U8805 (N_8805,N_6220,N_5454);
and U8806 (N_8806,N_7147,N_5228);
and U8807 (N_8807,N_7130,N_6226);
or U8808 (N_8808,N_7311,N_5683);
nor U8809 (N_8809,N_6248,N_5792);
nand U8810 (N_8810,N_6217,N_6918);
nor U8811 (N_8811,N_6932,N_7099);
nor U8812 (N_8812,N_5350,N_6623);
nand U8813 (N_8813,N_5708,N_6250);
xnor U8814 (N_8814,N_5778,N_6501);
or U8815 (N_8815,N_7075,N_6285);
and U8816 (N_8816,N_6026,N_6853);
nand U8817 (N_8817,N_5548,N_5901);
nor U8818 (N_8818,N_6119,N_6539);
and U8819 (N_8819,N_7344,N_7410);
and U8820 (N_8820,N_6489,N_5263);
xor U8821 (N_8821,N_5916,N_5606);
nand U8822 (N_8822,N_5638,N_6526);
or U8823 (N_8823,N_5456,N_6586);
nor U8824 (N_8824,N_6965,N_6643);
and U8825 (N_8825,N_5886,N_6118);
or U8826 (N_8826,N_7118,N_6304);
and U8827 (N_8827,N_7204,N_5230);
and U8828 (N_8828,N_5789,N_5731);
xnor U8829 (N_8829,N_5532,N_7304);
xor U8830 (N_8830,N_5994,N_7329);
nand U8831 (N_8831,N_5996,N_5159);
and U8832 (N_8832,N_5719,N_5281);
or U8833 (N_8833,N_6756,N_5269);
nand U8834 (N_8834,N_7298,N_6885);
and U8835 (N_8835,N_5701,N_7116);
nand U8836 (N_8836,N_7177,N_7429);
nand U8837 (N_8837,N_5817,N_6562);
and U8838 (N_8838,N_5787,N_7022);
nand U8839 (N_8839,N_6767,N_6845);
or U8840 (N_8840,N_6652,N_6209);
and U8841 (N_8841,N_6458,N_7470);
and U8842 (N_8842,N_5238,N_5270);
nor U8843 (N_8843,N_5509,N_5091);
nand U8844 (N_8844,N_6775,N_5125);
nand U8845 (N_8845,N_5472,N_5074);
xnor U8846 (N_8846,N_5890,N_6743);
or U8847 (N_8847,N_6810,N_5625);
or U8848 (N_8848,N_6477,N_5212);
and U8849 (N_8849,N_6972,N_5041);
nor U8850 (N_8850,N_5614,N_6241);
nor U8851 (N_8851,N_5839,N_5302);
nor U8852 (N_8852,N_5870,N_6127);
and U8853 (N_8853,N_6816,N_6697);
or U8854 (N_8854,N_5141,N_7450);
and U8855 (N_8855,N_5787,N_6514);
xor U8856 (N_8856,N_7428,N_6426);
and U8857 (N_8857,N_7460,N_6555);
or U8858 (N_8858,N_6324,N_5895);
xor U8859 (N_8859,N_6561,N_5102);
xor U8860 (N_8860,N_5687,N_6828);
or U8861 (N_8861,N_5116,N_7421);
nand U8862 (N_8862,N_5265,N_6729);
xnor U8863 (N_8863,N_5355,N_5037);
nor U8864 (N_8864,N_5854,N_5104);
nand U8865 (N_8865,N_6852,N_6058);
or U8866 (N_8866,N_6052,N_7438);
xnor U8867 (N_8867,N_6343,N_7081);
or U8868 (N_8868,N_6112,N_6304);
xor U8869 (N_8869,N_6292,N_5656);
nand U8870 (N_8870,N_6668,N_6086);
and U8871 (N_8871,N_5751,N_5229);
nand U8872 (N_8872,N_7470,N_5552);
or U8873 (N_8873,N_6248,N_5437);
nand U8874 (N_8874,N_5208,N_6149);
and U8875 (N_8875,N_6183,N_6118);
and U8876 (N_8876,N_6326,N_5927);
nand U8877 (N_8877,N_5300,N_7463);
nor U8878 (N_8878,N_6407,N_6994);
and U8879 (N_8879,N_5041,N_5303);
nor U8880 (N_8880,N_6131,N_7489);
nand U8881 (N_8881,N_6534,N_6193);
nand U8882 (N_8882,N_7103,N_5280);
nand U8883 (N_8883,N_7181,N_7356);
or U8884 (N_8884,N_7334,N_6398);
nand U8885 (N_8885,N_5335,N_6130);
nand U8886 (N_8886,N_5267,N_5940);
and U8887 (N_8887,N_7282,N_6985);
nor U8888 (N_8888,N_7409,N_5381);
or U8889 (N_8889,N_5622,N_5214);
and U8890 (N_8890,N_7197,N_7315);
and U8891 (N_8891,N_6128,N_6411);
nand U8892 (N_8892,N_6850,N_6223);
and U8893 (N_8893,N_6347,N_5973);
nor U8894 (N_8894,N_5463,N_5600);
and U8895 (N_8895,N_5611,N_6066);
nor U8896 (N_8896,N_6873,N_6438);
nor U8897 (N_8897,N_5886,N_6213);
or U8898 (N_8898,N_5778,N_6558);
and U8899 (N_8899,N_5093,N_5459);
or U8900 (N_8900,N_6965,N_6471);
nor U8901 (N_8901,N_7092,N_6689);
and U8902 (N_8902,N_7067,N_6188);
or U8903 (N_8903,N_7352,N_6382);
and U8904 (N_8904,N_5938,N_6381);
or U8905 (N_8905,N_5336,N_6902);
and U8906 (N_8906,N_7166,N_6764);
nor U8907 (N_8907,N_6632,N_6159);
and U8908 (N_8908,N_7492,N_6056);
nand U8909 (N_8909,N_5094,N_6206);
nor U8910 (N_8910,N_6826,N_6731);
xnor U8911 (N_8911,N_5620,N_7431);
and U8912 (N_8912,N_6202,N_5688);
nor U8913 (N_8913,N_5776,N_5595);
nand U8914 (N_8914,N_6040,N_6697);
and U8915 (N_8915,N_5286,N_5834);
nand U8916 (N_8916,N_7354,N_5055);
and U8917 (N_8917,N_6530,N_5377);
nor U8918 (N_8918,N_6305,N_6763);
or U8919 (N_8919,N_7097,N_5650);
nand U8920 (N_8920,N_7490,N_5336);
nand U8921 (N_8921,N_7103,N_6282);
and U8922 (N_8922,N_6752,N_6838);
xor U8923 (N_8923,N_6144,N_6378);
or U8924 (N_8924,N_5284,N_5572);
nand U8925 (N_8925,N_6335,N_5996);
nand U8926 (N_8926,N_6421,N_6985);
and U8927 (N_8927,N_7119,N_7115);
nor U8928 (N_8928,N_6207,N_6117);
and U8929 (N_8929,N_6129,N_7458);
nor U8930 (N_8930,N_5758,N_5605);
nand U8931 (N_8931,N_5247,N_5949);
nor U8932 (N_8932,N_5429,N_5991);
nor U8933 (N_8933,N_7129,N_7074);
and U8934 (N_8934,N_5535,N_7170);
and U8935 (N_8935,N_7043,N_6341);
nand U8936 (N_8936,N_6956,N_5657);
nand U8937 (N_8937,N_6463,N_6341);
and U8938 (N_8938,N_6580,N_6417);
nand U8939 (N_8939,N_5131,N_5012);
and U8940 (N_8940,N_6652,N_6595);
nand U8941 (N_8941,N_6233,N_5948);
nand U8942 (N_8942,N_7106,N_5526);
and U8943 (N_8943,N_5086,N_7040);
nand U8944 (N_8944,N_7071,N_5918);
nor U8945 (N_8945,N_5077,N_7133);
nor U8946 (N_8946,N_6352,N_7245);
or U8947 (N_8947,N_6912,N_5104);
nand U8948 (N_8948,N_6808,N_7301);
and U8949 (N_8949,N_5549,N_6287);
or U8950 (N_8950,N_6418,N_7460);
nand U8951 (N_8951,N_7355,N_6809);
and U8952 (N_8952,N_5363,N_6398);
nand U8953 (N_8953,N_7275,N_5882);
nor U8954 (N_8954,N_5585,N_6703);
or U8955 (N_8955,N_5364,N_6904);
xnor U8956 (N_8956,N_6527,N_5685);
or U8957 (N_8957,N_6895,N_5768);
nand U8958 (N_8958,N_6642,N_7332);
and U8959 (N_8959,N_5918,N_5228);
and U8960 (N_8960,N_5370,N_5881);
xor U8961 (N_8961,N_5891,N_6573);
nor U8962 (N_8962,N_6117,N_6801);
nand U8963 (N_8963,N_5536,N_5252);
or U8964 (N_8964,N_6950,N_7248);
nor U8965 (N_8965,N_5181,N_7332);
and U8966 (N_8966,N_6676,N_5966);
nor U8967 (N_8967,N_5803,N_7030);
and U8968 (N_8968,N_7125,N_5287);
and U8969 (N_8969,N_5853,N_5540);
nand U8970 (N_8970,N_5498,N_5861);
nand U8971 (N_8971,N_5663,N_5290);
nor U8972 (N_8972,N_6071,N_6765);
and U8973 (N_8973,N_7280,N_7034);
nand U8974 (N_8974,N_5970,N_6968);
and U8975 (N_8975,N_5801,N_5758);
and U8976 (N_8976,N_5973,N_7007);
xnor U8977 (N_8977,N_7083,N_6142);
nor U8978 (N_8978,N_6825,N_5939);
xnor U8979 (N_8979,N_6370,N_5562);
nor U8980 (N_8980,N_5520,N_6525);
and U8981 (N_8981,N_6257,N_6939);
nor U8982 (N_8982,N_6580,N_7494);
nor U8983 (N_8983,N_6611,N_5546);
nand U8984 (N_8984,N_5567,N_5928);
and U8985 (N_8985,N_5554,N_5749);
and U8986 (N_8986,N_5919,N_5964);
or U8987 (N_8987,N_6830,N_5890);
nand U8988 (N_8988,N_5514,N_7110);
nand U8989 (N_8989,N_7470,N_5034);
or U8990 (N_8990,N_6021,N_5772);
nand U8991 (N_8991,N_6461,N_5732);
nand U8992 (N_8992,N_6343,N_6015);
and U8993 (N_8993,N_5321,N_5654);
nand U8994 (N_8994,N_5417,N_6762);
or U8995 (N_8995,N_7063,N_6943);
or U8996 (N_8996,N_7360,N_6680);
nand U8997 (N_8997,N_5382,N_6124);
or U8998 (N_8998,N_5563,N_6108);
and U8999 (N_8999,N_7015,N_5983);
nand U9000 (N_9000,N_5442,N_6724);
and U9001 (N_9001,N_7387,N_5236);
nand U9002 (N_9002,N_7473,N_5582);
nor U9003 (N_9003,N_6351,N_6874);
nor U9004 (N_9004,N_6281,N_6270);
and U9005 (N_9005,N_7132,N_5718);
and U9006 (N_9006,N_7479,N_6672);
or U9007 (N_9007,N_6108,N_6642);
nand U9008 (N_9008,N_6182,N_6019);
nor U9009 (N_9009,N_7460,N_5364);
nor U9010 (N_9010,N_7438,N_7227);
xnor U9011 (N_9011,N_6089,N_6248);
and U9012 (N_9012,N_6242,N_6676);
or U9013 (N_9013,N_6572,N_6942);
nand U9014 (N_9014,N_6048,N_5501);
nand U9015 (N_9015,N_6438,N_5537);
or U9016 (N_9016,N_6136,N_5806);
xnor U9017 (N_9017,N_7144,N_5679);
or U9018 (N_9018,N_5419,N_5395);
and U9019 (N_9019,N_5686,N_7019);
nor U9020 (N_9020,N_5127,N_6376);
nand U9021 (N_9021,N_7111,N_5126);
nand U9022 (N_9022,N_6046,N_5700);
or U9023 (N_9023,N_5779,N_6545);
and U9024 (N_9024,N_5137,N_7231);
nor U9025 (N_9025,N_6684,N_5243);
or U9026 (N_9026,N_5622,N_5466);
or U9027 (N_9027,N_7039,N_5427);
and U9028 (N_9028,N_5692,N_5789);
xnor U9029 (N_9029,N_5359,N_5397);
nor U9030 (N_9030,N_5744,N_5448);
and U9031 (N_9031,N_6847,N_7013);
or U9032 (N_9032,N_5611,N_7404);
nor U9033 (N_9033,N_5029,N_5979);
and U9034 (N_9034,N_5790,N_5353);
xor U9035 (N_9035,N_5082,N_6527);
and U9036 (N_9036,N_5906,N_5379);
nand U9037 (N_9037,N_5885,N_5971);
nor U9038 (N_9038,N_7016,N_5664);
or U9039 (N_9039,N_7328,N_6216);
or U9040 (N_9040,N_6480,N_5971);
xnor U9041 (N_9041,N_5447,N_5552);
nor U9042 (N_9042,N_5617,N_6343);
nand U9043 (N_9043,N_7250,N_5745);
or U9044 (N_9044,N_6489,N_7335);
or U9045 (N_9045,N_5738,N_7167);
or U9046 (N_9046,N_6126,N_5421);
nor U9047 (N_9047,N_6694,N_6220);
and U9048 (N_9048,N_5024,N_7097);
and U9049 (N_9049,N_5386,N_5586);
xor U9050 (N_9050,N_5723,N_5347);
and U9051 (N_9051,N_5362,N_6957);
or U9052 (N_9052,N_6595,N_7033);
nor U9053 (N_9053,N_5266,N_6169);
nand U9054 (N_9054,N_6570,N_5810);
xor U9055 (N_9055,N_6230,N_5699);
nand U9056 (N_9056,N_5770,N_6310);
and U9057 (N_9057,N_5385,N_5153);
and U9058 (N_9058,N_5606,N_7222);
or U9059 (N_9059,N_5440,N_5820);
nand U9060 (N_9060,N_5902,N_5715);
nor U9061 (N_9061,N_6707,N_6522);
and U9062 (N_9062,N_5627,N_7051);
xor U9063 (N_9063,N_6295,N_5408);
nand U9064 (N_9064,N_6245,N_6685);
nand U9065 (N_9065,N_5309,N_6152);
or U9066 (N_9066,N_5185,N_5974);
or U9067 (N_9067,N_7110,N_6387);
or U9068 (N_9068,N_6238,N_7037);
xnor U9069 (N_9069,N_7110,N_7029);
xnor U9070 (N_9070,N_7298,N_6696);
and U9071 (N_9071,N_6727,N_5639);
and U9072 (N_9072,N_6324,N_5887);
or U9073 (N_9073,N_5114,N_6439);
nor U9074 (N_9074,N_7328,N_6878);
xnor U9075 (N_9075,N_5964,N_5785);
nand U9076 (N_9076,N_6132,N_5490);
nand U9077 (N_9077,N_6420,N_5981);
nor U9078 (N_9078,N_5557,N_7334);
nor U9079 (N_9079,N_6814,N_6597);
nor U9080 (N_9080,N_5369,N_5810);
or U9081 (N_9081,N_6184,N_5447);
and U9082 (N_9082,N_6430,N_5559);
and U9083 (N_9083,N_5583,N_6924);
nand U9084 (N_9084,N_6589,N_6429);
nor U9085 (N_9085,N_5149,N_7107);
or U9086 (N_9086,N_5719,N_6103);
xnor U9087 (N_9087,N_5009,N_5419);
nand U9088 (N_9088,N_6771,N_5588);
nand U9089 (N_9089,N_7449,N_6803);
and U9090 (N_9090,N_5191,N_5396);
nor U9091 (N_9091,N_5232,N_5857);
or U9092 (N_9092,N_5462,N_7129);
or U9093 (N_9093,N_7022,N_6471);
nor U9094 (N_9094,N_5801,N_6821);
nand U9095 (N_9095,N_6134,N_6063);
xor U9096 (N_9096,N_6229,N_5088);
and U9097 (N_9097,N_6841,N_5179);
xor U9098 (N_9098,N_5370,N_7478);
and U9099 (N_9099,N_5817,N_5951);
nand U9100 (N_9100,N_6487,N_6342);
nor U9101 (N_9101,N_6927,N_7156);
or U9102 (N_9102,N_6352,N_5786);
nand U9103 (N_9103,N_6254,N_6541);
or U9104 (N_9104,N_5197,N_7371);
and U9105 (N_9105,N_6064,N_6059);
or U9106 (N_9106,N_5610,N_5858);
and U9107 (N_9107,N_5144,N_5428);
or U9108 (N_9108,N_6418,N_5048);
or U9109 (N_9109,N_6464,N_5168);
and U9110 (N_9110,N_5918,N_5382);
nor U9111 (N_9111,N_7378,N_5018);
or U9112 (N_9112,N_5037,N_6304);
xor U9113 (N_9113,N_7232,N_6380);
nand U9114 (N_9114,N_7442,N_6853);
or U9115 (N_9115,N_6752,N_5561);
nand U9116 (N_9116,N_5169,N_6455);
and U9117 (N_9117,N_7290,N_5393);
and U9118 (N_9118,N_6397,N_5170);
and U9119 (N_9119,N_6738,N_5812);
nor U9120 (N_9120,N_5696,N_6912);
and U9121 (N_9121,N_6657,N_5057);
or U9122 (N_9122,N_5803,N_5374);
nor U9123 (N_9123,N_5165,N_6312);
or U9124 (N_9124,N_6518,N_5531);
and U9125 (N_9125,N_6822,N_5662);
or U9126 (N_9126,N_5525,N_6816);
nor U9127 (N_9127,N_5544,N_6878);
and U9128 (N_9128,N_6511,N_5511);
nor U9129 (N_9129,N_7291,N_7249);
or U9130 (N_9130,N_5225,N_7135);
nand U9131 (N_9131,N_7348,N_6285);
or U9132 (N_9132,N_7393,N_6194);
or U9133 (N_9133,N_6301,N_7434);
and U9134 (N_9134,N_6631,N_5875);
xnor U9135 (N_9135,N_5684,N_5855);
xor U9136 (N_9136,N_5804,N_6305);
nor U9137 (N_9137,N_7438,N_5645);
nand U9138 (N_9138,N_5315,N_7445);
and U9139 (N_9139,N_7011,N_6736);
and U9140 (N_9140,N_7100,N_5902);
nand U9141 (N_9141,N_6476,N_7422);
nand U9142 (N_9142,N_5266,N_6812);
nor U9143 (N_9143,N_5209,N_6663);
nor U9144 (N_9144,N_7180,N_5681);
xor U9145 (N_9145,N_5886,N_5005);
xor U9146 (N_9146,N_7435,N_6535);
nand U9147 (N_9147,N_6600,N_7166);
or U9148 (N_9148,N_5278,N_7329);
nor U9149 (N_9149,N_6211,N_6009);
and U9150 (N_9150,N_7408,N_6764);
nor U9151 (N_9151,N_5047,N_5050);
nor U9152 (N_9152,N_6094,N_5987);
nand U9153 (N_9153,N_5071,N_5141);
or U9154 (N_9154,N_7483,N_6180);
and U9155 (N_9155,N_5609,N_5967);
nor U9156 (N_9156,N_6296,N_5715);
nor U9157 (N_9157,N_5393,N_6704);
nor U9158 (N_9158,N_6175,N_5337);
or U9159 (N_9159,N_5858,N_5435);
xnor U9160 (N_9160,N_6632,N_6410);
and U9161 (N_9161,N_5234,N_7252);
xor U9162 (N_9162,N_5016,N_5146);
nor U9163 (N_9163,N_6951,N_6131);
nor U9164 (N_9164,N_6146,N_7209);
and U9165 (N_9165,N_6257,N_6389);
or U9166 (N_9166,N_6220,N_5281);
or U9167 (N_9167,N_6612,N_5939);
and U9168 (N_9168,N_5934,N_7497);
or U9169 (N_9169,N_5665,N_6757);
and U9170 (N_9170,N_5079,N_5855);
and U9171 (N_9171,N_5007,N_5418);
nor U9172 (N_9172,N_5460,N_7131);
or U9173 (N_9173,N_5190,N_5429);
xnor U9174 (N_9174,N_5468,N_6804);
xnor U9175 (N_9175,N_7245,N_5861);
nor U9176 (N_9176,N_6790,N_7037);
and U9177 (N_9177,N_5249,N_6160);
nand U9178 (N_9178,N_7320,N_5907);
and U9179 (N_9179,N_6873,N_5880);
or U9180 (N_9180,N_7371,N_5239);
nor U9181 (N_9181,N_5577,N_7095);
or U9182 (N_9182,N_6742,N_5129);
nand U9183 (N_9183,N_5873,N_6426);
xor U9184 (N_9184,N_6227,N_7036);
nor U9185 (N_9185,N_6555,N_5297);
or U9186 (N_9186,N_5439,N_5665);
nor U9187 (N_9187,N_7434,N_6946);
or U9188 (N_9188,N_5623,N_5390);
and U9189 (N_9189,N_5792,N_6291);
and U9190 (N_9190,N_7020,N_7428);
or U9191 (N_9191,N_5922,N_6369);
or U9192 (N_9192,N_6193,N_7105);
nand U9193 (N_9193,N_5312,N_5291);
and U9194 (N_9194,N_6849,N_5242);
or U9195 (N_9195,N_7069,N_6662);
nor U9196 (N_9196,N_5247,N_5466);
and U9197 (N_9197,N_7396,N_7393);
nand U9198 (N_9198,N_5795,N_7196);
nand U9199 (N_9199,N_5317,N_5755);
nor U9200 (N_9200,N_5039,N_5266);
nor U9201 (N_9201,N_6993,N_6295);
nand U9202 (N_9202,N_5838,N_7164);
nand U9203 (N_9203,N_7085,N_7470);
nor U9204 (N_9204,N_5745,N_6135);
or U9205 (N_9205,N_6355,N_5968);
and U9206 (N_9206,N_5103,N_6719);
nand U9207 (N_9207,N_6354,N_6394);
nor U9208 (N_9208,N_5125,N_6028);
and U9209 (N_9209,N_5685,N_7147);
nand U9210 (N_9210,N_7366,N_5275);
nand U9211 (N_9211,N_6800,N_6419);
and U9212 (N_9212,N_5949,N_5381);
and U9213 (N_9213,N_5106,N_7298);
or U9214 (N_9214,N_7204,N_7240);
and U9215 (N_9215,N_5857,N_7342);
nor U9216 (N_9216,N_6908,N_6411);
nor U9217 (N_9217,N_5280,N_6245);
and U9218 (N_9218,N_5981,N_7258);
nor U9219 (N_9219,N_5254,N_6417);
or U9220 (N_9220,N_5087,N_7250);
and U9221 (N_9221,N_7423,N_6582);
or U9222 (N_9222,N_6364,N_7335);
or U9223 (N_9223,N_6859,N_7363);
or U9224 (N_9224,N_5688,N_6848);
and U9225 (N_9225,N_5034,N_7109);
xor U9226 (N_9226,N_5937,N_7454);
and U9227 (N_9227,N_5963,N_5294);
or U9228 (N_9228,N_6391,N_5717);
and U9229 (N_9229,N_7078,N_6132);
and U9230 (N_9230,N_6838,N_5562);
nor U9231 (N_9231,N_6609,N_5579);
nor U9232 (N_9232,N_5097,N_6264);
or U9233 (N_9233,N_5381,N_7358);
xor U9234 (N_9234,N_7169,N_7310);
or U9235 (N_9235,N_7481,N_5001);
and U9236 (N_9236,N_5314,N_6887);
xor U9237 (N_9237,N_6429,N_7220);
xor U9238 (N_9238,N_5065,N_6475);
and U9239 (N_9239,N_7289,N_5323);
and U9240 (N_9240,N_5301,N_5940);
or U9241 (N_9241,N_6296,N_6091);
or U9242 (N_9242,N_6110,N_6093);
nand U9243 (N_9243,N_6572,N_6176);
nor U9244 (N_9244,N_5684,N_5313);
and U9245 (N_9245,N_6938,N_5827);
nand U9246 (N_9246,N_5282,N_7080);
and U9247 (N_9247,N_6050,N_5778);
nor U9248 (N_9248,N_6768,N_5908);
xnor U9249 (N_9249,N_7448,N_6767);
and U9250 (N_9250,N_7221,N_7050);
or U9251 (N_9251,N_5080,N_5564);
nand U9252 (N_9252,N_5355,N_5624);
xor U9253 (N_9253,N_6430,N_5360);
nand U9254 (N_9254,N_6433,N_5839);
nand U9255 (N_9255,N_7457,N_5950);
nand U9256 (N_9256,N_5159,N_7172);
xnor U9257 (N_9257,N_6978,N_7117);
nand U9258 (N_9258,N_6219,N_6522);
nand U9259 (N_9259,N_5838,N_5490);
nor U9260 (N_9260,N_5962,N_6000);
nor U9261 (N_9261,N_6380,N_5589);
nand U9262 (N_9262,N_6662,N_7141);
or U9263 (N_9263,N_5790,N_6590);
nor U9264 (N_9264,N_6419,N_6309);
and U9265 (N_9265,N_6460,N_6700);
nand U9266 (N_9266,N_6103,N_6591);
nand U9267 (N_9267,N_6527,N_5888);
nand U9268 (N_9268,N_7213,N_6681);
nand U9269 (N_9269,N_5797,N_6226);
nand U9270 (N_9270,N_7054,N_5458);
and U9271 (N_9271,N_6401,N_5042);
nor U9272 (N_9272,N_7185,N_5312);
xor U9273 (N_9273,N_5305,N_5568);
nand U9274 (N_9274,N_6365,N_5445);
or U9275 (N_9275,N_6051,N_7029);
nor U9276 (N_9276,N_6333,N_6227);
and U9277 (N_9277,N_5690,N_6860);
xnor U9278 (N_9278,N_5645,N_7011);
or U9279 (N_9279,N_7059,N_7026);
nor U9280 (N_9280,N_5180,N_5846);
xnor U9281 (N_9281,N_5250,N_5494);
and U9282 (N_9282,N_5919,N_6203);
xnor U9283 (N_9283,N_7005,N_5283);
nor U9284 (N_9284,N_5252,N_5630);
nor U9285 (N_9285,N_6536,N_6978);
nor U9286 (N_9286,N_5133,N_6069);
and U9287 (N_9287,N_6814,N_6062);
or U9288 (N_9288,N_7415,N_5375);
and U9289 (N_9289,N_5990,N_7224);
nor U9290 (N_9290,N_6121,N_6858);
nor U9291 (N_9291,N_5243,N_5240);
nor U9292 (N_9292,N_5166,N_5819);
nand U9293 (N_9293,N_5534,N_5875);
nor U9294 (N_9294,N_5369,N_5111);
nand U9295 (N_9295,N_5534,N_5710);
nand U9296 (N_9296,N_5917,N_5429);
nand U9297 (N_9297,N_7253,N_7367);
and U9298 (N_9298,N_5840,N_5585);
and U9299 (N_9299,N_5020,N_7490);
and U9300 (N_9300,N_7023,N_6661);
nand U9301 (N_9301,N_6113,N_5434);
nand U9302 (N_9302,N_5636,N_5625);
or U9303 (N_9303,N_7282,N_6372);
and U9304 (N_9304,N_7023,N_6774);
nand U9305 (N_9305,N_6615,N_5426);
nand U9306 (N_9306,N_7057,N_6883);
nand U9307 (N_9307,N_5026,N_7275);
nand U9308 (N_9308,N_6013,N_5697);
nor U9309 (N_9309,N_5704,N_5922);
nor U9310 (N_9310,N_6105,N_5098);
nor U9311 (N_9311,N_5589,N_7008);
or U9312 (N_9312,N_5818,N_6851);
xnor U9313 (N_9313,N_7421,N_6326);
nor U9314 (N_9314,N_7422,N_7293);
nand U9315 (N_9315,N_6103,N_6035);
nor U9316 (N_9316,N_5963,N_6897);
nand U9317 (N_9317,N_6429,N_6927);
nor U9318 (N_9318,N_6066,N_7071);
and U9319 (N_9319,N_5285,N_6540);
and U9320 (N_9320,N_5860,N_5331);
nand U9321 (N_9321,N_5794,N_6406);
or U9322 (N_9322,N_5530,N_5678);
nor U9323 (N_9323,N_7373,N_5614);
xnor U9324 (N_9324,N_6989,N_5801);
nand U9325 (N_9325,N_6985,N_6129);
nor U9326 (N_9326,N_6765,N_6068);
or U9327 (N_9327,N_6881,N_5015);
and U9328 (N_9328,N_5328,N_6822);
and U9329 (N_9329,N_7285,N_6631);
and U9330 (N_9330,N_6410,N_6734);
xor U9331 (N_9331,N_5528,N_7230);
nor U9332 (N_9332,N_6839,N_6056);
nand U9333 (N_9333,N_6939,N_6084);
or U9334 (N_9334,N_7470,N_5453);
nor U9335 (N_9335,N_5040,N_5368);
or U9336 (N_9336,N_6241,N_6406);
or U9337 (N_9337,N_7262,N_5096);
xor U9338 (N_9338,N_6562,N_5659);
nand U9339 (N_9339,N_7346,N_5199);
and U9340 (N_9340,N_5376,N_6126);
nor U9341 (N_9341,N_6026,N_5142);
nand U9342 (N_9342,N_6319,N_6393);
nor U9343 (N_9343,N_5037,N_6009);
xnor U9344 (N_9344,N_6668,N_6671);
xnor U9345 (N_9345,N_5122,N_5510);
nor U9346 (N_9346,N_6183,N_6792);
nand U9347 (N_9347,N_7189,N_6594);
and U9348 (N_9348,N_5594,N_6385);
nor U9349 (N_9349,N_5068,N_5752);
or U9350 (N_9350,N_6954,N_5622);
or U9351 (N_9351,N_5964,N_5723);
nor U9352 (N_9352,N_7094,N_5592);
xor U9353 (N_9353,N_6476,N_6143);
nand U9354 (N_9354,N_5389,N_7170);
nand U9355 (N_9355,N_6364,N_5683);
and U9356 (N_9356,N_7387,N_7245);
nor U9357 (N_9357,N_6232,N_7012);
or U9358 (N_9358,N_5832,N_5827);
nor U9359 (N_9359,N_6798,N_5510);
xnor U9360 (N_9360,N_7485,N_7460);
nand U9361 (N_9361,N_6252,N_5843);
or U9362 (N_9362,N_7498,N_5903);
and U9363 (N_9363,N_5528,N_5503);
nand U9364 (N_9364,N_5005,N_5037);
or U9365 (N_9365,N_6268,N_5310);
and U9366 (N_9366,N_5558,N_6097);
nand U9367 (N_9367,N_6333,N_6697);
or U9368 (N_9368,N_6715,N_6072);
xnor U9369 (N_9369,N_6994,N_6432);
or U9370 (N_9370,N_5831,N_6945);
nor U9371 (N_9371,N_6636,N_5582);
nor U9372 (N_9372,N_5969,N_5146);
nand U9373 (N_9373,N_6424,N_7186);
nand U9374 (N_9374,N_6934,N_5311);
nor U9375 (N_9375,N_6315,N_6442);
and U9376 (N_9376,N_6134,N_7206);
and U9377 (N_9377,N_7377,N_6827);
nor U9378 (N_9378,N_7440,N_6498);
or U9379 (N_9379,N_7437,N_6275);
nand U9380 (N_9380,N_6832,N_6254);
xor U9381 (N_9381,N_6899,N_5971);
or U9382 (N_9382,N_5097,N_7257);
and U9383 (N_9383,N_7331,N_6324);
nor U9384 (N_9384,N_6697,N_6384);
nor U9385 (N_9385,N_6552,N_6303);
nand U9386 (N_9386,N_7081,N_5273);
nand U9387 (N_9387,N_6925,N_5991);
and U9388 (N_9388,N_6026,N_5476);
nor U9389 (N_9389,N_5640,N_6415);
nor U9390 (N_9390,N_5430,N_6278);
or U9391 (N_9391,N_6789,N_5178);
and U9392 (N_9392,N_6577,N_7381);
or U9393 (N_9393,N_5433,N_6613);
or U9394 (N_9394,N_6010,N_6475);
and U9395 (N_9395,N_7177,N_7160);
or U9396 (N_9396,N_5512,N_6651);
nand U9397 (N_9397,N_5795,N_6292);
and U9398 (N_9398,N_6855,N_5090);
or U9399 (N_9399,N_5667,N_6475);
nand U9400 (N_9400,N_6402,N_7122);
nor U9401 (N_9401,N_7154,N_5893);
xor U9402 (N_9402,N_7063,N_5847);
nor U9403 (N_9403,N_5063,N_6023);
and U9404 (N_9404,N_6218,N_5700);
nand U9405 (N_9405,N_5464,N_6897);
or U9406 (N_9406,N_6009,N_5529);
and U9407 (N_9407,N_6142,N_5336);
or U9408 (N_9408,N_6671,N_6757);
or U9409 (N_9409,N_7411,N_5475);
xor U9410 (N_9410,N_6791,N_5388);
or U9411 (N_9411,N_5687,N_5598);
xnor U9412 (N_9412,N_6218,N_6513);
nor U9413 (N_9413,N_6118,N_7005);
xnor U9414 (N_9414,N_7353,N_6876);
or U9415 (N_9415,N_6170,N_7314);
and U9416 (N_9416,N_5386,N_6444);
or U9417 (N_9417,N_7113,N_6233);
nor U9418 (N_9418,N_6620,N_6208);
xnor U9419 (N_9419,N_5445,N_7107);
nor U9420 (N_9420,N_6388,N_5057);
nor U9421 (N_9421,N_6878,N_7466);
nand U9422 (N_9422,N_5796,N_7181);
xnor U9423 (N_9423,N_7104,N_6300);
nor U9424 (N_9424,N_5505,N_6724);
nand U9425 (N_9425,N_6133,N_6631);
nor U9426 (N_9426,N_6936,N_6980);
nor U9427 (N_9427,N_6190,N_7396);
nor U9428 (N_9428,N_7361,N_5104);
and U9429 (N_9429,N_7069,N_6117);
or U9430 (N_9430,N_5674,N_7045);
and U9431 (N_9431,N_5356,N_7402);
xnor U9432 (N_9432,N_5267,N_5063);
nand U9433 (N_9433,N_6967,N_7154);
nor U9434 (N_9434,N_5867,N_7436);
or U9435 (N_9435,N_5152,N_6686);
and U9436 (N_9436,N_5839,N_5644);
nor U9437 (N_9437,N_5272,N_6310);
and U9438 (N_9438,N_6962,N_5982);
nor U9439 (N_9439,N_7417,N_6908);
nand U9440 (N_9440,N_6994,N_6499);
or U9441 (N_9441,N_6160,N_5129);
or U9442 (N_9442,N_5506,N_6949);
or U9443 (N_9443,N_7493,N_5864);
and U9444 (N_9444,N_5815,N_5726);
or U9445 (N_9445,N_5242,N_6673);
nor U9446 (N_9446,N_7059,N_5800);
and U9447 (N_9447,N_6359,N_7005);
nor U9448 (N_9448,N_6721,N_6117);
xnor U9449 (N_9449,N_5844,N_5690);
nor U9450 (N_9450,N_6893,N_5764);
or U9451 (N_9451,N_5225,N_5487);
nand U9452 (N_9452,N_5582,N_5621);
nand U9453 (N_9453,N_5993,N_7415);
and U9454 (N_9454,N_5568,N_6983);
and U9455 (N_9455,N_6521,N_5331);
and U9456 (N_9456,N_7398,N_5619);
nand U9457 (N_9457,N_7235,N_6612);
or U9458 (N_9458,N_6060,N_5267);
and U9459 (N_9459,N_5335,N_5247);
xor U9460 (N_9460,N_7406,N_6315);
nand U9461 (N_9461,N_5167,N_6307);
nand U9462 (N_9462,N_7005,N_6756);
and U9463 (N_9463,N_7248,N_7458);
nand U9464 (N_9464,N_6517,N_6708);
xnor U9465 (N_9465,N_7046,N_5894);
or U9466 (N_9466,N_6352,N_6656);
nor U9467 (N_9467,N_6626,N_7088);
or U9468 (N_9468,N_5701,N_5804);
nand U9469 (N_9469,N_6974,N_6090);
and U9470 (N_9470,N_7432,N_6817);
or U9471 (N_9471,N_5859,N_6110);
and U9472 (N_9472,N_5305,N_6142);
or U9473 (N_9473,N_7218,N_6819);
or U9474 (N_9474,N_7338,N_6206);
nand U9475 (N_9475,N_7383,N_5383);
nor U9476 (N_9476,N_5264,N_5689);
nor U9477 (N_9477,N_6359,N_5037);
or U9478 (N_9478,N_6893,N_7411);
nand U9479 (N_9479,N_5769,N_7280);
nor U9480 (N_9480,N_5926,N_6137);
or U9481 (N_9481,N_6977,N_5827);
nand U9482 (N_9482,N_5292,N_7116);
and U9483 (N_9483,N_5492,N_6340);
and U9484 (N_9484,N_6313,N_7356);
nand U9485 (N_9485,N_5264,N_5076);
nor U9486 (N_9486,N_5403,N_6538);
or U9487 (N_9487,N_7271,N_5941);
nor U9488 (N_9488,N_6107,N_6480);
or U9489 (N_9489,N_5996,N_6424);
or U9490 (N_9490,N_5292,N_5105);
or U9491 (N_9491,N_6006,N_5821);
or U9492 (N_9492,N_6326,N_6488);
and U9493 (N_9493,N_6741,N_6286);
or U9494 (N_9494,N_6265,N_6403);
and U9495 (N_9495,N_7451,N_5366);
and U9496 (N_9496,N_5017,N_5746);
or U9497 (N_9497,N_5095,N_7451);
or U9498 (N_9498,N_7099,N_6435);
nor U9499 (N_9499,N_5886,N_6452);
nand U9500 (N_9500,N_6633,N_7136);
nor U9501 (N_9501,N_5879,N_5122);
nor U9502 (N_9502,N_7152,N_6962);
or U9503 (N_9503,N_6389,N_6371);
nor U9504 (N_9504,N_5519,N_6400);
nor U9505 (N_9505,N_6422,N_5237);
nor U9506 (N_9506,N_7072,N_5370);
nand U9507 (N_9507,N_7483,N_6889);
or U9508 (N_9508,N_5217,N_5431);
nor U9509 (N_9509,N_7149,N_7300);
and U9510 (N_9510,N_7227,N_6944);
nand U9511 (N_9511,N_6511,N_6928);
and U9512 (N_9512,N_5636,N_5299);
nor U9513 (N_9513,N_6541,N_6381);
and U9514 (N_9514,N_6378,N_6337);
nor U9515 (N_9515,N_7380,N_7141);
nor U9516 (N_9516,N_5931,N_7020);
or U9517 (N_9517,N_7223,N_5747);
and U9518 (N_9518,N_5461,N_7238);
or U9519 (N_9519,N_6006,N_5940);
nand U9520 (N_9520,N_5929,N_5312);
or U9521 (N_9521,N_5538,N_7394);
nor U9522 (N_9522,N_5278,N_5799);
nand U9523 (N_9523,N_6109,N_5174);
nand U9524 (N_9524,N_7187,N_5951);
nor U9525 (N_9525,N_5498,N_6870);
nor U9526 (N_9526,N_6671,N_7436);
nand U9527 (N_9527,N_5105,N_5829);
nand U9528 (N_9528,N_5916,N_5269);
or U9529 (N_9529,N_6186,N_6903);
nand U9530 (N_9530,N_7117,N_5846);
nor U9531 (N_9531,N_6601,N_6350);
or U9532 (N_9532,N_5902,N_5965);
nand U9533 (N_9533,N_6667,N_6316);
nor U9534 (N_9534,N_6721,N_5231);
and U9535 (N_9535,N_6888,N_5662);
nand U9536 (N_9536,N_7195,N_6419);
or U9537 (N_9537,N_5635,N_5725);
or U9538 (N_9538,N_5665,N_5899);
and U9539 (N_9539,N_5439,N_6825);
or U9540 (N_9540,N_7088,N_7383);
nor U9541 (N_9541,N_5433,N_7284);
xor U9542 (N_9542,N_6480,N_6811);
nand U9543 (N_9543,N_5043,N_5472);
nand U9544 (N_9544,N_7050,N_6066);
and U9545 (N_9545,N_6897,N_6416);
nand U9546 (N_9546,N_6388,N_6760);
nor U9547 (N_9547,N_6557,N_6519);
xnor U9548 (N_9548,N_5431,N_5724);
xor U9549 (N_9549,N_5616,N_6548);
nand U9550 (N_9550,N_5973,N_5073);
or U9551 (N_9551,N_5374,N_5908);
nor U9552 (N_9552,N_7354,N_5193);
or U9553 (N_9553,N_7044,N_5510);
or U9554 (N_9554,N_6475,N_6454);
nand U9555 (N_9555,N_5210,N_5870);
nor U9556 (N_9556,N_5878,N_5802);
xor U9557 (N_9557,N_7061,N_5063);
and U9558 (N_9558,N_7416,N_5630);
or U9559 (N_9559,N_5536,N_5316);
or U9560 (N_9560,N_5583,N_6141);
xnor U9561 (N_9561,N_5925,N_5204);
or U9562 (N_9562,N_6231,N_5361);
and U9563 (N_9563,N_5068,N_5322);
nor U9564 (N_9564,N_5370,N_6141);
or U9565 (N_9565,N_5276,N_5076);
nand U9566 (N_9566,N_7039,N_5021);
and U9567 (N_9567,N_6227,N_7165);
and U9568 (N_9568,N_6439,N_5465);
nor U9569 (N_9569,N_5942,N_6616);
or U9570 (N_9570,N_7424,N_6350);
xnor U9571 (N_9571,N_7175,N_5293);
and U9572 (N_9572,N_6245,N_7024);
nand U9573 (N_9573,N_6772,N_6512);
nor U9574 (N_9574,N_6388,N_6546);
or U9575 (N_9575,N_5485,N_5094);
or U9576 (N_9576,N_6964,N_5308);
and U9577 (N_9577,N_6133,N_6319);
nor U9578 (N_9578,N_7333,N_7287);
nand U9579 (N_9579,N_5440,N_7352);
or U9580 (N_9580,N_5586,N_5389);
and U9581 (N_9581,N_6090,N_6296);
and U9582 (N_9582,N_5658,N_7114);
xnor U9583 (N_9583,N_5475,N_5155);
nand U9584 (N_9584,N_7327,N_5627);
nand U9585 (N_9585,N_5697,N_5848);
and U9586 (N_9586,N_5733,N_7427);
xor U9587 (N_9587,N_5166,N_6647);
and U9588 (N_9588,N_7480,N_6528);
xnor U9589 (N_9589,N_5742,N_7389);
nand U9590 (N_9590,N_6874,N_7185);
nor U9591 (N_9591,N_5424,N_5916);
and U9592 (N_9592,N_5072,N_5116);
and U9593 (N_9593,N_6490,N_6569);
and U9594 (N_9594,N_7145,N_5247);
and U9595 (N_9595,N_7249,N_5415);
nand U9596 (N_9596,N_6976,N_7056);
or U9597 (N_9597,N_5361,N_5225);
nor U9598 (N_9598,N_5464,N_5989);
or U9599 (N_9599,N_5820,N_6398);
nand U9600 (N_9600,N_5941,N_7422);
xnor U9601 (N_9601,N_7306,N_6936);
and U9602 (N_9602,N_6639,N_7183);
nor U9603 (N_9603,N_5358,N_7187);
and U9604 (N_9604,N_5804,N_7435);
nor U9605 (N_9605,N_6004,N_6711);
or U9606 (N_9606,N_5525,N_6427);
nor U9607 (N_9607,N_5664,N_5068);
and U9608 (N_9608,N_5711,N_6332);
nand U9609 (N_9609,N_6658,N_6783);
nand U9610 (N_9610,N_6301,N_5538);
and U9611 (N_9611,N_7343,N_5331);
nor U9612 (N_9612,N_7460,N_6512);
and U9613 (N_9613,N_6210,N_6356);
nor U9614 (N_9614,N_6301,N_5350);
and U9615 (N_9615,N_5607,N_6298);
nand U9616 (N_9616,N_6960,N_5846);
nor U9617 (N_9617,N_5172,N_6759);
nand U9618 (N_9618,N_6489,N_6193);
nand U9619 (N_9619,N_6651,N_5514);
nor U9620 (N_9620,N_6902,N_6030);
or U9621 (N_9621,N_5465,N_7370);
nor U9622 (N_9622,N_5623,N_6728);
or U9623 (N_9623,N_5531,N_6963);
or U9624 (N_9624,N_6449,N_7439);
or U9625 (N_9625,N_5638,N_5101);
nor U9626 (N_9626,N_7139,N_5893);
xor U9627 (N_9627,N_5662,N_5804);
or U9628 (N_9628,N_7104,N_5699);
nor U9629 (N_9629,N_7347,N_6666);
xnor U9630 (N_9630,N_6122,N_7278);
xnor U9631 (N_9631,N_6553,N_5279);
nand U9632 (N_9632,N_7336,N_6358);
nor U9633 (N_9633,N_6178,N_6337);
nor U9634 (N_9634,N_5692,N_7180);
and U9635 (N_9635,N_5730,N_6682);
and U9636 (N_9636,N_6983,N_5481);
and U9637 (N_9637,N_6767,N_6757);
nor U9638 (N_9638,N_5366,N_5915);
nor U9639 (N_9639,N_5795,N_6801);
nand U9640 (N_9640,N_7205,N_5324);
and U9641 (N_9641,N_7166,N_6906);
nor U9642 (N_9642,N_5853,N_6847);
xor U9643 (N_9643,N_7340,N_6494);
nand U9644 (N_9644,N_5921,N_6997);
nor U9645 (N_9645,N_6304,N_6678);
or U9646 (N_9646,N_6568,N_5443);
and U9647 (N_9647,N_7076,N_5575);
and U9648 (N_9648,N_6098,N_6850);
nand U9649 (N_9649,N_6630,N_6124);
nor U9650 (N_9650,N_6158,N_5673);
nor U9651 (N_9651,N_6879,N_7486);
and U9652 (N_9652,N_5213,N_5828);
nor U9653 (N_9653,N_6806,N_6539);
or U9654 (N_9654,N_5812,N_5927);
or U9655 (N_9655,N_6738,N_5471);
nor U9656 (N_9656,N_5525,N_5126);
xor U9657 (N_9657,N_7373,N_5618);
xnor U9658 (N_9658,N_6859,N_7043);
or U9659 (N_9659,N_6512,N_6855);
or U9660 (N_9660,N_5228,N_7181);
nand U9661 (N_9661,N_6224,N_7148);
or U9662 (N_9662,N_6740,N_5338);
and U9663 (N_9663,N_6786,N_6849);
nand U9664 (N_9664,N_6410,N_5329);
or U9665 (N_9665,N_7393,N_6135);
or U9666 (N_9666,N_6771,N_6462);
or U9667 (N_9667,N_5315,N_5477);
nand U9668 (N_9668,N_6252,N_5687);
or U9669 (N_9669,N_7371,N_6314);
or U9670 (N_9670,N_6926,N_6227);
nor U9671 (N_9671,N_7259,N_7010);
nand U9672 (N_9672,N_6222,N_6748);
or U9673 (N_9673,N_5095,N_7154);
nand U9674 (N_9674,N_5325,N_7132);
nor U9675 (N_9675,N_7193,N_6539);
or U9676 (N_9676,N_5042,N_6252);
and U9677 (N_9677,N_6309,N_6109);
or U9678 (N_9678,N_7467,N_6569);
nand U9679 (N_9679,N_6053,N_6306);
nand U9680 (N_9680,N_5638,N_7279);
and U9681 (N_9681,N_6498,N_6096);
nor U9682 (N_9682,N_5195,N_6911);
or U9683 (N_9683,N_5652,N_6812);
nand U9684 (N_9684,N_6485,N_6566);
nand U9685 (N_9685,N_5326,N_6413);
and U9686 (N_9686,N_5868,N_5845);
and U9687 (N_9687,N_6496,N_5404);
nor U9688 (N_9688,N_6587,N_7366);
nand U9689 (N_9689,N_5336,N_7223);
or U9690 (N_9690,N_6018,N_7468);
and U9691 (N_9691,N_5614,N_6601);
and U9692 (N_9692,N_6140,N_5097);
nor U9693 (N_9693,N_6801,N_7131);
nor U9694 (N_9694,N_6931,N_6102);
nand U9695 (N_9695,N_6567,N_6845);
nand U9696 (N_9696,N_5143,N_6873);
nor U9697 (N_9697,N_6843,N_7217);
nor U9698 (N_9698,N_5984,N_7349);
nand U9699 (N_9699,N_6180,N_7300);
xnor U9700 (N_9700,N_7414,N_6684);
or U9701 (N_9701,N_7328,N_6584);
or U9702 (N_9702,N_6414,N_6371);
nand U9703 (N_9703,N_6282,N_6682);
nand U9704 (N_9704,N_5429,N_7287);
and U9705 (N_9705,N_6038,N_5033);
nor U9706 (N_9706,N_5801,N_5509);
nor U9707 (N_9707,N_5377,N_5496);
or U9708 (N_9708,N_6505,N_6806);
nor U9709 (N_9709,N_6922,N_5312);
nand U9710 (N_9710,N_5816,N_7320);
and U9711 (N_9711,N_6704,N_6428);
nand U9712 (N_9712,N_5447,N_6941);
nand U9713 (N_9713,N_5099,N_6166);
xor U9714 (N_9714,N_5610,N_5845);
xor U9715 (N_9715,N_6545,N_5483);
nor U9716 (N_9716,N_5789,N_6925);
or U9717 (N_9717,N_6609,N_6627);
nand U9718 (N_9718,N_5973,N_6769);
and U9719 (N_9719,N_7492,N_5870);
nor U9720 (N_9720,N_6431,N_7375);
nand U9721 (N_9721,N_6786,N_6335);
or U9722 (N_9722,N_7252,N_6652);
nor U9723 (N_9723,N_5464,N_6267);
xnor U9724 (N_9724,N_6224,N_6506);
or U9725 (N_9725,N_5620,N_5651);
nand U9726 (N_9726,N_6479,N_5864);
or U9727 (N_9727,N_7087,N_6363);
nand U9728 (N_9728,N_6494,N_5577);
or U9729 (N_9729,N_6136,N_6021);
nor U9730 (N_9730,N_5697,N_6399);
nor U9731 (N_9731,N_5294,N_6345);
and U9732 (N_9732,N_5726,N_6104);
or U9733 (N_9733,N_5803,N_7375);
nand U9734 (N_9734,N_5319,N_6678);
and U9735 (N_9735,N_5325,N_6519);
nand U9736 (N_9736,N_5645,N_6768);
or U9737 (N_9737,N_6669,N_7230);
nand U9738 (N_9738,N_7227,N_5768);
and U9739 (N_9739,N_7232,N_6423);
and U9740 (N_9740,N_5657,N_7029);
nor U9741 (N_9741,N_7346,N_5030);
nor U9742 (N_9742,N_5232,N_5880);
and U9743 (N_9743,N_7218,N_5014);
nor U9744 (N_9744,N_6314,N_7055);
nand U9745 (N_9745,N_5305,N_6192);
and U9746 (N_9746,N_5876,N_5463);
or U9747 (N_9747,N_7029,N_5284);
or U9748 (N_9748,N_5280,N_6422);
and U9749 (N_9749,N_5999,N_6734);
and U9750 (N_9750,N_5762,N_5442);
or U9751 (N_9751,N_5368,N_6950);
xnor U9752 (N_9752,N_7041,N_7004);
nor U9753 (N_9753,N_5852,N_6031);
and U9754 (N_9754,N_5924,N_5373);
nor U9755 (N_9755,N_6036,N_6887);
or U9756 (N_9756,N_5338,N_5616);
or U9757 (N_9757,N_5262,N_6184);
and U9758 (N_9758,N_5321,N_7452);
or U9759 (N_9759,N_5360,N_6168);
or U9760 (N_9760,N_6043,N_7400);
xnor U9761 (N_9761,N_5957,N_6328);
or U9762 (N_9762,N_7069,N_7143);
nand U9763 (N_9763,N_6102,N_7190);
xor U9764 (N_9764,N_7165,N_7160);
nor U9765 (N_9765,N_5247,N_5849);
and U9766 (N_9766,N_7201,N_5296);
or U9767 (N_9767,N_7119,N_7193);
nor U9768 (N_9768,N_6974,N_7185);
nand U9769 (N_9769,N_7333,N_6532);
xor U9770 (N_9770,N_5738,N_6633);
nand U9771 (N_9771,N_6334,N_5642);
nor U9772 (N_9772,N_5757,N_6099);
nor U9773 (N_9773,N_6129,N_7112);
and U9774 (N_9774,N_7387,N_5726);
and U9775 (N_9775,N_6624,N_5133);
or U9776 (N_9776,N_5941,N_6815);
or U9777 (N_9777,N_6522,N_7470);
nor U9778 (N_9778,N_6029,N_6569);
or U9779 (N_9779,N_6180,N_6272);
xor U9780 (N_9780,N_6132,N_6394);
and U9781 (N_9781,N_6129,N_6112);
nand U9782 (N_9782,N_7447,N_6314);
xnor U9783 (N_9783,N_6870,N_5073);
nand U9784 (N_9784,N_5850,N_5123);
nand U9785 (N_9785,N_5229,N_6379);
nand U9786 (N_9786,N_5233,N_5083);
nor U9787 (N_9787,N_6932,N_5034);
or U9788 (N_9788,N_6281,N_6825);
or U9789 (N_9789,N_5348,N_6201);
nand U9790 (N_9790,N_7324,N_5434);
nand U9791 (N_9791,N_5674,N_6328);
xnor U9792 (N_9792,N_5621,N_6139);
nand U9793 (N_9793,N_6219,N_6089);
and U9794 (N_9794,N_6146,N_7040);
xnor U9795 (N_9795,N_5440,N_5739);
nor U9796 (N_9796,N_5577,N_6157);
and U9797 (N_9797,N_6441,N_5157);
nand U9798 (N_9798,N_6008,N_6242);
nor U9799 (N_9799,N_5041,N_5611);
or U9800 (N_9800,N_5589,N_7242);
and U9801 (N_9801,N_6707,N_6227);
and U9802 (N_9802,N_5182,N_7121);
nand U9803 (N_9803,N_5455,N_7256);
nand U9804 (N_9804,N_7423,N_6947);
or U9805 (N_9805,N_5016,N_5271);
or U9806 (N_9806,N_7462,N_6495);
nand U9807 (N_9807,N_7345,N_7385);
or U9808 (N_9808,N_5448,N_6120);
or U9809 (N_9809,N_6077,N_5168);
or U9810 (N_9810,N_5143,N_6026);
nor U9811 (N_9811,N_5759,N_6669);
nor U9812 (N_9812,N_6658,N_5722);
xor U9813 (N_9813,N_6651,N_5162);
or U9814 (N_9814,N_5043,N_5206);
nor U9815 (N_9815,N_6194,N_5368);
xnor U9816 (N_9816,N_6730,N_7055);
nand U9817 (N_9817,N_5893,N_6568);
or U9818 (N_9818,N_5553,N_7016);
nor U9819 (N_9819,N_6834,N_5599);
nor U9820 (N_9820,N_6168,N_6320);
and U9821 (N_9821,N_5232,N_7314);
nor U9822 (N_9822,N_5689,N_6865);
nor U9823 (N_9823,N_5924,N_6285);
or U9824 (N_9824,N_6612,N_6160);
and U9825 (N_9825,N_5044,N_6990);
or U9826 (N_9826,N_7433,N_5589);
nand U9827 (N_9827,N_5393,N_6178);
xor U9828 (N_9828,N_5940,N_5296);
nand U9829 (N_9829,N_7445,N_6061);
or U9830 (N_9830,N_5100,N_6799);
or U9831 (N_9831,N_5492,N_6855);
or U9832 (N_9832,N_6923,N_7070);
nand U9833 (N_9833,N_6369,N_5180);
and U9834 (N_9834,N_6687,N_5167);
nand U9835 (N_9835,N_6645,N_6537);
or U9836 (N_9836,N_6134,N_7335);
nand U9837 (N_9837,N_6632,N_6601);
or U9838 (N_9838,N_6275,N_6028);
nand U9839 (N_9839,N_5481,N_6399);
and U9840 (N_9840,N_6706,N_6439);
nand U9841 (N_9841,N_5182,N_5361);
and U9842 (N_9842,N_5571,N_6543);
and U9843 (N_9843,N_7498,N_6262);
nor U9844 (N_9844,N_6099,N_5594);
or U9845 (N_9845,N_6506,N_6505);
nand U9846 (N_9846,N_5561,N_5919);
nand U9847 (N_9847,N_6805,N_7069);
nand U9848 (N_9848,N_5197,N_7433);
and U9849 (N_9849,N_5432,N_5062);
xor U9850 (N_9850,N_6987,N_6348);
and U9851 (N_9851,N_5933,N_6642);
nand U9852 (N_9852,N_6936,N_7262);
or U9853 (N_9853,N_7372,N_7162);
nor U9854 (N_9854,N_7003,N_6286);
xor U9855 (N_9855,N_6212,N_6757);
nand U9856 (N_9856,N_5434,N_6962);
and U9857 (N_9857,N_7066,N_5498);
nor U9858 (N_9858,N_5342,N_5186);
or U9859 (N_9859,N_7148,N_5133);
or U9860 (N_9860,N_6649,N_7303);
nor U9861 (N_9861,N_7305,N_6763);
and U9862 (N_9862,N_6983,N_5715);
nor U9863 (N_9863,N_5588,N_5807);
or U9864 (N_9864,N_6668,N_7223);
or U9865 (N_9865,N_7250,N_5775);
xor U9866 (N_9866,N_6495,N_6405);
and U9867 (N_9867,N_7113,N_6443);
nand U9868 (N_9868,N_5431,N_6315);
and U9869 (N_9869,N_6490,N_7402);
and U9870 (N_9870,N_6830,N_5227);
or U9871 (N_9871,N_7139,N_6337);
nor U9872 (N_9872,N_6025,N_5974);
nand U9873 (N_9873,N_5721,N_5333);
or U9874 (N_9874,N_6546,N_6659);
or U9875 (N_9875,N_5720,N_5777);
nor U9876 (N_9876,N_6801,N_7077);
and U9877 (N_9877,N_6361,N_7015);
and U9878 (N_9878,N_5876,N_6772);
nand U9879 (N_9879,N_6142,N_7349);
and U9880 (N_9880,N_6357,N_5868);
nor U9881 (N_9881,N_5448,N_7395);
nor U9882 (N_9882,N_7087,N_5341);
xnor U9883 (N_9883,N_5081,N_5387);
or U9884 (N_9884,N_6865,N_5618);
or U9885 (N_9885,N_5177,N_6018);
or U9886 (N_9886,N_5718,N_6429);
or U9887 (N_9887,N_7175,N_5216);
or U9888 (N_9888,N_5128,N_5836);
nand U9889 (N_9889,N_6395,N_5784);
nand U9890 (N_9890,N_6424,N_5948);
nand U9891 (N_9891,N_5377,N_5064);
nor U9892 (N_9892,N_6857,N_6324);
nand U9893 (N_9893,N_5466,N_5522);
xor U9894 (N_9894,N_7337,N_5139);
nand U9895 (N_9895,N_6344,N_7116);
and U9896 (N_9896,N_5340,N_5126);
and U9897 (N_9897,N_6243,N_7300);
nor U9898 (N_9898,N_5299,N_5917);
nand U9899 (N_9899,N_6207,N_6279);
xnor U9900 (N_9900,N_7360,N_5946);
nor U9901 (N_9901,N_6840,N_7034);
nand U9902 (N_9902,N_6081,N_5941);
nor U9903 (N_9903,N_6685,N_7442);
or U9904 (N_9904,N_6712,N_6375);
and U9905 (N_9905,N_6611,N_6431);
or U9906 (N_9906,N_5955,N_5807);
nor U9907 (N_9907,N_5513,N_6013);
nand U9908 (N_9908,N_5598,N_5542);
nor U9909 (N_9909,N_5633,N_7042);
and U9910 (N_9910,N_5653,N_6323);
nand U9911 (N_9911,N_7424,N_6630);
nor U9912 (N_9912,N_6522,N_5184);
or U9913 (N_9913,N_5010,N_6385);
nand U9914 (N_9914,N_7102,N_5776);
or U9915 (N_9915,N_5137,N_5680);
nand U9916 (N_9916,N_5199,N_6237);
nand U9917 (N_9917,N_5490,N_5764);
or U9918 (N_9918,N_7238,N_5868);
or U9919 (N_9919,N_6145,N_6537);
or U9920 (N_9920,N_5864,N_5506);
or U9921 (N_9921,N_6775,N_6679);
nor U9922 (N_9922,N_6231,N_6494);
nor U9923 (N_9923,N_6224,N_6248);
nor U9924 (N_9924,N_6568,N_6481);
and U9925 (N_9925,N_5644,N_7019);
nor U9926 (N_9926,N_5748,N_6381);
or U9927 (N_9927,N_7345,N_6225);
and U9928 (N_9928,N_5302,N_5907);
xor U9929 (N_9929,N_5286,N_5461);
nor U9930 (N_9930,N_6759,N_7153);
and U9931 (N_9931,N_7334,N_5562);
nor U9932 (N_9932,N_5795,N_7137);
nor U9933 (N_9933,N_6915,N_5874);
nor U9934 (N_9934,N_6330,N_5025);
and U9935 (N_9935,N_5835,N_5594);
or U9936 (N_9936,N_5860,N_5085);
nand U9937 (N_9937,N_5055,N_6644);
and U9938 (N_9938,N_6902,N_5786);
nand U9939 (N_9939,N_6218,N_7146);
xor U9940 (N_9940,N_5088,N_5363);
nor U9941 (N_9941,N_5938,N_6727);
nand U9942 (N_9942,N_6949,N_5984);
nor U9943 (N_9943,N_6454,N_6359);
nand U9944 (N_9944,N_5764,N_6712);
xor U9945 (N_9945,N_6084,N_6413);
nand U9946 (N_9946,N_5627,N_6314);
xor U9947 (N_9947,N_5737,N_5112);
nand U9948 (N_9948,N_6680,N_5876);
nor U9949 (N_9949,N_7027,N_6422);
nand U9950 (N_9950,N_6505,N_5209);
and U9951 (N_9951,N_5411,N_5867);
and U9952 (N_9952,N_5300,N_7317);
nand U9953 (N_9953,N_5984,N_5641);
and U9954 (N_9954,N_7403,N_5698);
and U9955 (N_9955,N_6541,N_5983);
and U9956 (N_9956,N_6320,N_5638);
xor U9957 (N_9957,N_6450,N_7108);
xor U9958 (N_9958,N_6104,N_6184);
and U9959 (N_9959,N_6889,N_5058);
nor U9960 (N_9960,N_6861,N_5047);
xor U9961 (N_9961,N_6254,N_6112);
or U9962 (N_9962,N_5336,N_5477);
xor U9963 (N_9963,N_6486,N_6382);
xnor U9964 (N_9964,N_6354,N_5960);
nand U9965 (N_9965,N_6035,N_5334);
nand U9966 (N_9966,N_5744,N_5591);
or U9967 (N_9967,N_6349,N_5171);
xor U9968 (N_9968,N_7465,N_5144);
or U9969 (N_9969,N_6047,N_5482);
and U9970 (N_9970,N_6250,N_6466);
or U9971 (N_9971,N_7045,N_6491);
or U9972 (N_9972,N_6395,N_6139);
or U9973 (N_9973,N_7294,N_5728);
and U9974 (N_9974,N_7133,N_7102);
or U9975 (N_9975,N_6091,N_5198);
and U9976 (N_9976,N_7002,N_5413);
and U9977 (N_9977,N_6519,N_6696);
nor U9978 (N_9978,N_5383,N_5429);
or U9979 (N_9979,N_6874,N_5722);
nand U9980 (N_9980,N_6475,N_6104);
nand U9981 (N_9981,N_5369,N_7185);
or U9982 (N_9982,N_6386,N_5827);
nor U9983 (N_9983,N_5779,N_6516);
and U9984 (N_9984,N_6923,N_6859);
or U9985 (N_9985,N_5850,N_7169);
and U9986 (N_9986,N_5827,N_6048);
and U9987 (N_9987,N_5692,N_7277);
xor U9988 (N_9988,N_6481,N_6754);
nand U9989 (N_9989,N_5862,N_5802);
or U9990 (N_9990,N_5212,N_6084);
nand U9991 (N_9991,N_5203,N_5954);
nor U9992 (N_9992,N_7154,N_6241);
nand U9993 (N_9993,N_7327,N_7228);
nor U9994 (N_9994,N_5507,N_6891);
and U9995 (N_9995,N_7118,N_6850);
nand U9996 (N_9996,N_6093,N_7127);
nor U9997 (N_9997,N_5237,N_5955);
or U9998 (N_9998,N_6072,N_5014);
nand U9999 (N_9999,N_6111,N_5091);
or UO_0 (O_0,N_8892,N_9007);
nand UO_1 (O_1,N_7650,N_9306);
and UO_2 (O_2,N_9985,N_9705);
or UO_3 (O_3,N_9297,N_7609);
nor UO_4 (O_4,N_8242,N_8549);
nand UO_5 (O_5,N_8719,N_9065);
and UO_6 (O_6,N_8486,N_9248);
nand UO_7 (O_7,N_8378,N_7613);
nor UO_8 (O_8,N_8603,N_9477);
nand UO_9 (O_9,N_8703,N_9743);
nor UO_10 (O_10,N_8034,N_8291);
nor UO_11 (O_11,N_7800,N_8890);
xor UO_12 (O_12,N_9046,N_7965);
nor UO_13 (O_13,N_8962,N_9425);
nor UO_14 (O_14,N_8701,N_7707);
nor UO_15 (O_15,N_8080,N_9259);
nand UO_16 (O_16,N_8094,N_9176);
or UO_17 (O_17,N_7601,N_8302);
nor UO_18 (O_18,N_9202,N_9878);
or UO_19 (O_19,N_9844,N_9055);
nand UO_20 (O_20,N_9278,N_7566);
nand UO_21 (O_21,N_8572,N_9390);
and UO_22 (O_22,N_7698,N_7579);
and UO_23 (O_23,N_9876,N_7668);
nor UO_24 (O_24,N_8609,N_8154);
or UO_25 (O_25,N_9106,N_7558);
or UO_26 (O_26,N_7894,N_9081);
or UO_27 (O_27,N_7665,N_9851);
and UO_28 (O_28,N_9508,N_7563);
nand UO_29 (O_29,N_9076,N_8573);
or UO_30 (O_30,N_8619,N_8313);
nand UO_31 (O_31,N_9734,N_7737);
or UO_32 (O_32,N_8553,N_9920);
nor UO_33 (O_33,N_7789,N_8853);
or UO_34 (O_34,N_9972,N_8206);
or UO_35 (O_35,N_8384,N_7733);
nor UO_36 (O_36,N_9562,N_8991);
nor UO_37 (O_37,N_8002,N_9690);
nor UO_38 (O_38,N_7876,N_9197);
nand UO_39 (O_39,N_9152,N_7856);
nand UO_40 (O_40,N_8941,N_7525);
nor UO_41 (O_41,N_9386,N_9184);
xor UO_42 (O_42,N_9245,N_9513);
and UO_43 (O_43,N_8851,N_8629);
xnor UO_44 (O_44,N_8237,N_8491);
nor UO_45 (O_45,N_9312,N_7997);
nand UO_46 (O_46,N_9244,N_9540);
nor UO_47 (O_47,N_8811,N_8031);
or UO_48 (O_48,N_7532,N_7598);
and UO_49 (O_49,N_7785,N_8540);
and UO_50 (O_50,N_9607,N_9216);
or UO_51 (O_51,N_8663,N_8321);
xnor UO_52 (O_52,N_8833,N_7996);
nor UO_53 (O_53,N_9915,N_9588);
and UO_54 (O_54,N_8781,N_8454);
nor UO_55 (O_55,N_7752,N_9012);
and UO_56 (O_56,N_7618,N_9883);
nor UO_57 (O_57,N_9196,N_7500);
or UO_58 (O_58,N_7725,N_7683);
and UO_59 (O_59,N_9582,N_9002);
nand UO_60 (O_60,N_8303,N_8896);
or UO_61 (O_61,N_9603,N_8182);
or UO_62 (O_62,N_8219,N_9472);
nand UO_63 (O_63,N_7773,N_8787);
nand UO_64 (O_64,N_8382,N_9810);
and UO_65 (O_65,N_8116,N_9892);
nand UO_66 (O_66,N_9195,N_9147);
and UO_67 (O_67,N_7635,N_8596);
nor UO_68 (O_68,N_7984,N_8944);
nand UO_69 (O_69,N_9489,N_8907);
or UO_70 (O_70,N_9396,N_7775);
nand UO_71 (O_71,N_8457,N_7592);
or UO_72 (O_72,N_9635,N_8058);
or UO_73 (O_73,N_9251,N_8394);
and UO_74 (O_74,N_9865,N_7763);
and UO_75 (O_75,N_9073,N_9090);
and UO_76 (O_76,N_7616,N_8104);
or UO_77 (O_77,N_8235,N_8396);
or UO_78 (O_78,N_8096,N_9449);
or UO_79 (O_79,N_8153,N_9101);
or UO_80 (O_80,N_9515,N_7565);
nand UO_81 (O_81,N_7739,N_7845);
xnor UO_82 (O_82,N_9178,N_7864);
nor UO_83 (O_83,N_7872,N_8584);
or UO_84 (O_84,N_7854,N_9177);
and UO_85 (O_85,N_8969,N_7813);
and UO_86 (O_86,N_9601,N_9187);
nor UO_87 (O_87,N_9256,N_9381);
or UO_88 (O_88,N_7895,N_9406);
nand UO_89 (O_89,N_8174,N_9080);
nand UO_90 (O_90,N_9547,N_8471);
or UO_91 (O_91,N_9591,N_7559);
nor UO_92 (O_92,N_9655,N_7780);
or UO_93 (O_93,N_9552,N_9824);
or UO_94 (O_94,N_7553,N_7719);
nand UO_95 (O_95,N_8751,N_8839);
and UO_96 (O_96,N_8708,N_8156);
nor UO_97 (O_97,N_8904,N_7806);
nand UO_98 (O_98,N_8957,N_8685);
and UO_99 (O_99,N_7961,N_7726);
and UO_100 (O_100,N_7514,N_7667);
nand UO_101 (O_101,N_9088,N_7906);
nor UO_102 (O_102,N_7839,N_9193);
and UO_103 (O_103,N_9203,N_9232);
nand UO_104 (O_104,N_8292,N_8450);
and UO_105 (O_105,N_8790,N_9079);
or UO_106 (O_106,N_7796,N_9509);
nor UO_107 (O_107,N_9965,N_9338);
nor UO_108 (O_108,N_7974,N_9186);
or UO_109 (O_109,N_8294,N_9541);
and UO_110 (O_110,N_8501,N_8379);
or UO_111 (O_111,N_8634,N_9872);
nor UO_112 (O_112,N_7907,N_8232);
nand UO_113 (O_113,N_8591,N_9052);
nor UO_114 (O_114,N_9426,N_9558);
or UO_115 (O_115,N_7717,N_9856);
nand UO_116 (O_116,N_8920,N_9314);
xnor UO_117 (O_117,N_7935,N_9355);
and UO_118 (O_118,N_9628,N_8534);
xor UO_119 (O_119,N_7824,N_9093);
nand UO_120 (O_120,N_8823,N_8914);
or UO_121 (O_121,N_8694,N_9014);
nor UO_122 (O_122,N_9040,N_8846);
nand UO_123 (O_123,N_8271,N_9163);
nor UO_124 (O_124,N_9910,N_8871);
nand UO_125 (O_125,N_8638,N_7669);
nand UO_126 (O_126,N_7643,N_8628);
and UO_127 (O_127,N_9740,N_8352);
and UO_128 (O_128,N_9776,N_9391);
nor UO_129 (O_129,N_9484,N_8929);
or UO_130 (O_130,N_8583,N_8247);
nor UO_131 (O_131,N_9836,N_7594);
and UO_132 (O_132,N_9980,N_9373);
and UO_133 (O_133,N_8420,N_8705);
and UO_134 (O_134,N_9399,N_9284);
and UO_135 (O_135,N_8903,N_9434);
nand UO_136 (O_136,N_9181,N_8806);
nand UO_137 (O_137,N_9099,N_8395);
or UO_138 (O_138,N_9718,N_7969);
xor UO_139 (O_139,N_8563,N_8084);
or UO_140 (O_140,N_9480,N_8802);
or UO_141 (O_141,N_9246,N_9201);
or UO_142 (O_142,N_9672,N_7639);
or UO_143 (O_143,N_9866,N_9868);
nor UO_144 (O_144,N_8455,N_8124);
or UO_145 (O_145,N_8590,N_8180);
and UO_146 (O_146,N_9648,N_9621);
and UO_147 (O_147,N_8356,N_7747);
nand UO_148 (O_148,N_7851,N_9975);
or UO_149 (O_149,N_8986,N_8643);
nand UO_150 (O_150,N_7917,N_8622);
or UO_151 (O_151,N_8776,N_8618);
and UO_152 (O_152,N_8073,N_7925);
nor UO_153 (O_153,N_9986,N_8223);
nand UO_154 (O_154,N_8524,N_9213);
nor UO_155 (O_155,N_9017,N_9961);
nand UO_156 (O_156,N_9930,N_8481);
nand UO_157 (O_157,N_9801,N_7597);
and UO_158 (O_158,N_8438,N_8865);
nor UO_159 (O_159,N_8998,N_8426);
nor UO_160 (O_160,N_7945,N_8308);
xnor UO_161 (O_161,N_8318,N_8211);
nor UO_162 (O_162,N_7896,N_8574);
and UO_163 (O_163,N_7831,N_7638);
nor UO_164 (O_164,N_8393,N_7644);
and UO_165 (O_165,N_9009,N_9673);
or UO_166 (O_166,N_8607,N_7509);
and UO_167 (O_167,N_7664,N_7911);
and UO_168 (O_168,N_8359,N_8770);
or UO_169 (O_169,N_8389,N_8692);
nor UO_170 (O_170,N_9899,N_7732);
nand UO_171 (O_171,N_7569,N_8550);
and UO_172 (O_172,N_8240,N_9759);
and UO_173 (O_173,N_8143,N_9574);
nor UO_174 (O_174,N_8829,N_8430);
nand UO_175 (O_175,N_9650,N_8671);
nand UO_176 (O_176,N_9544,N_9559);
or UO_177 (O_177,N_7611,N_8878);
nand UO_178 (O_178,N_9971,N_8078);
and UO_179 (O_179,N_8448,N_8456);
nand UO_180 (O_180,N_9863,N_8774);
xor UO_181 (O_181,N_7678,N_8431);
and UO_182 (O_182,N_9424,N_9159);
nand UO_183 (O_183,N_8905,N_7867);
xor UO_184 (O_184,N_9882,N_8830);
and UO_185 (O_185,N_7825,N_8676);
nand UO_186 (O_186,N_8891,N_9483);
nand UO_187 (O_187,N_8979,N_8244);
nor UO_188 (O_188,N_8465,N_8411);
nand UO_189 (O_189,N_9659,N_8256);
or UO_190 (O_190,N_9634,N_7966);
xor UO_191 (O_191,N_8314,N_8615);
nand UO_192 (O_192,N_8970,N_7718);
and UO_193 (O_193,N_8726,N_8516);
or UO_194 (O_194,N_8275,N_9991);
nor UO_195 (O_195,N_8898,N_8707);
nand UO_196 (O_196,N_9632,N_8295);
nor UO_197 (O_197,N_8548,N_7521);
and UO_198 (O_198,N_8300,N_8882);
or UO_199 (O_199,N_8383,N_8675);
nor UO_200 (O_200,N_9611,N_7786);
nor UO_201 (O_201,N_8526,N_9857);
and UO_202 (O_202,N_8155,N_8681);
and UO_203 (O_203,N_9457,N_9565);
nand UO_204 (O_204,N_7788,N_9885);
xnor UO_205 (O_205,N_7771,N_9416);
nand UO_206 (O_206,N_8644,N_9606);
xnor UO_207 (O_207,N_9904,N_9821);
nand UO_208 (O_208,N_9639,N_9614);
nand UO_209 (O_209,N_8228,N_8742);
and UO_210 (O_210,N_9198,N_9267);
nand UO_211 (O_211,N_7970,N_9658);
xnor UO_212 (O_212,N_9510,N_9078);
and UO_213 (O_213,N_8068,N_9696);
nand UO_214 (O_214,N_9160,N_8400);
xor UO_215 (O_215,N_8391,N_8207);
xor UO_216 (O_216,N_9794,N_7507);
xnor UO_217 (O_217,N_7673,N_8253);
nor UO_218 (O_218,N_8640,N_8786);
or UO_219 (O_219,N_8873,N_9733);
and UO_220 (O_220,N_9837,N_8995);
nand UO_221 (O_221,N_8737,N_9624);
or UO_222 (O_222,N_8799,N_8807);
or UO_223 (O_223,N_7899,N_8771);
or UO_224 (O_224,N_7715,N_8899);
or UO_225 (O_225,N_9567,N_8445);
and UO_226 (O_226,N_7921,N_9895);
nand UO_227 (O_227,N_9226,N_7955);
nand UO_228 (O_228,N_8693,N_8305);
and UO_229 (O_229,N_8441,N_8716);
nand UO_230 (O_230,N_9001,N_9324);
and UO_231 (O_231,N_8033,N_7994);
or UO_232 (O_232,N_8337,N_7617);
nor UO_233 (O_233,N_8290,N_8010);
and UO_234 (O_234,N_8557,N_8673);
nor UO_235 (O_235,N_7814,N_9485);
and UO_236 (O_236,N_9263,N_9296);
nor UO_237 (O_237,N_7977,N_9738);
or UO_238 (O_238,N_9933,N_9727);
nand UO_239 (O_239,N_8924,N_8349);
or UO_240 (O_240,N_9229,N_8564);
xor UO_241 (O_241,N_7608,N_9576);
and UO_242 (O_242,N_7588,N_9493);
and UO_243 (O_243,N_9927,N_9819);
and UO_244 (O_244,N_9891,N_9744);
nor UO_245 (O_245,N_7539,N_9110);
nand UO_246 (O_246,N_7656,N_8879);
nand UO_247 (O_247,N_9630,N_9735);
nor UO_248 (O_248,N_9652,N_8911);
nand UO_249 (O_249,N_8926,N_9905);
and UO_250 (O_250,N_8588,N_9726);
or UO_251 (O_251,N_8171,N_9115);
and UO_252 (O_252,N_7956,N_9664);
or UO_253 (O_253,N_7541,N_9311);
and UO_254 (O_254,N_7585,N_9988);
or UO_255 (O_255,N_9506,N_8505);
or UO_256 (O_256,N_9901,N_8993);
xor UO_257 (O_257,N_8141,N_7892);
and UO_258 (O_258,N_7741,N_9403);
and UO_259 (O_259,N_9966,N_8086);
and UO_260 (O_260,N_8630,N_7940);
or UO_261 (O_261,N_9709,N_9539);
nand UO_262 (O_262,N_9959,N_7950);
and UO_263 (O_263,N_9765,N_8076);
nor UO_264 (O_264,N_7686,N_8436);
nor UO_265 (O_265,N_8016,N_7783);
and UO_266 (O_266,N_9722,N_8815);
and UO_267 (O_267,N_9250,N_7684);
and UO_268 (O_268,N_8561,N_9584);
nor UO_269 (O_269,N_9520,N_8131);
nor UO_270 (O_270,N_8079,N_8385);
nand UO_271 (O_271,N_9505,N_7551);
or UO_272 (O_272,N_8442,N_9271);
and UO_273 (O_273,N_7760,N_7702);
nor UO_274 (O_274,N_8398,N_8810);
or UO_275 (O_275,N_8361,N_9304);
nor UO_276 (O_276,N_9784,N_7846);
or UO_277 (O_277,N_9981,N_9431);
xnor UO_278 (O_278,N_9122,N_7697);
nor UO_279 (O_279,N_9269,N_8040);
xnor UO_280 (O_280,N_9850,N_8115);
nand UO_281 (O_281,N_8416,N_9413);
and UO_282 (O_282,N_7999,N_9602);
xor UO_283 (O_283,N_9907,N_8162);
xor UO_284 (O_284,N_7808,N_8315);
and UO_285 (O_285,N_8281,N_7882);
nor UO_286 (O_286,N_9318,N_9841);
nor UO_287 (O_287,N_9149,N_9706);
nand UO_288 (O_288,N_7666,N_8888);
and UO_289 (O_289,N_7602,N_9037);
nor UO_290 (O_290,N_9770,N_8801);
xor UO_291 (O_291,N_9827,N_8097);
nor UO_292 (O_292,N_8554,N_8578);
and UO_293 (O_293,N_7502,N_8645);
or UO_294 (O_294,N_7904,N_7651);
nand UO_295 (O_295,N_7556,N_8813);
nor UO_296 (O_296,N_9687,N_8056);
nand UO_297 (O_297,N_9678,N_8380);
nor UO_298 (O_298,N_9380,N_7740);
or UO_299 (O_299,N_9649,N_8921);
and UO_300 (O_300,N_8089,N_9400);
and UO_301 (O_301,N_8325,N_8472);
nor UO_302 (O_302,N_7949,N_9613);
nand UO_303 (O_303,N_9916,N_8095);
or UO_304 (O_304,N_7934,N_9204);
nand UO_305 (O_305,N_9979,N_9501);
and UO_306 (O_306,N_9697,N_7570);
nand UO_307 (O_307,N_8772,N_8241);
nand UO_308 (O_308,N_9288,N_8566);
nor UO_309 (O_309,N_9473,N_8345);
nor UO_310 (O_310,N_9071,N_9121);
xor UO_311 (O_311,N_7908,N_9124);
nor UO_312 (O_312,N_7975,N_9041);
nand UO_313 (O_313,N_9045,N_8412);
or UO_314 (O_314,N_7630,N_8714);
nand UO_315 (O_315,N_8433,N_7843);
or UO_316 (O_316,N_8371,N_8715);
and UO_317 (O_317,N_9732,N_7875);
nor UO_318 (O_318,N_9710,N_9585);
nor UO_319 (O_319,N_8005,N_8468);
nand UO_320 (O_320,N_8976,N_7822);
and UO_321 (O_321,N_9166,N_7755);
xor UO_322 (O_322,N_8024,N_8977);
nor UO_323 (O_323,N_8082,N_8343);
or UO_324 (O_324,N_8243,N_8215);
nand UO_325 (O_325,N_9517,N_8949);
nor UO_326 (O_326,N_9035,N_8713);
and UO_327 (O_327,N_8023,N_9242);
and UO_328 (O_328,N_9643,N_7811);
and UO_329 (O_329,N_8170,N_7654);
and UO_330 (O_330,N_9623,N_9091);
nor UO_331 (O_331,N_9283,N_9771);
and UO_332 (O_332,N_8586,N_9908);
nor UO_333 (O_333,N_7535,N_8307);
and UO_334 (O_334,N_8667,N_9367);
or UO_335 (O_335,N_8906,N_7764);
nand UO_336 (O_336,N_8651,N_9977);
nor UO_337 (O_337,N_7998,N_9736);
nand UO_338 (O_338,N_9884,N_8221);
or UO_339 (O_339,N_7931,N_8199);
and UO_340 (O_340,N_7593,N_9793);
or UO_341 (O_341,N_9835,N_9702);
or UO_342 (O_342,N_8458,N_9873);
and UO_343 (O_343,N_9340,N_8494);
nor UO_344 (O_344,N_8852,N_9828);
xnor UO_345 (O_345,N_9536,N_9179);
nand UO_346 (O_346,N_8624,N_9225);
nand UO_347 (O_347,N_7634,N_9138);
nor UO_348 (O_348,N_8778,N_9523);
nand UO_349 (O_349,N_8710,N_7869);
nor UO_350 (O_350,N_8805,N_8504);
and UO_351 (O_351,N_9970,N_7818);
nand UO_352 (O_352,N_9504,N_8868);
and UO_353 (O_353,N_8869,N_8809);
nor UO_354 (O_354,N_8985,N_8777);
or UO_355 (O_355,N_8376,N_8533);
or UO_356 (O_356,N_7847,N_9731);
nor UO_357 (O_357,N_8014,N_8492);
and UO_358 (O_358,N_7736,N_9875);
nor UO_359 (O_359,N_8915,N_9212);
or UO_360 (O_360,N_9796,N_9174);
nand UO_361 (O_361,N_8405,N_9600);
nor UO_362 (O_362,N_7751,N_9345);
or UO_363 (O_363,N_8415,N_8796);
and UO_364 (O_364,N_9441,N_8425);
or UO_365 (O_365,N_9753,N_9125);
nand UO_366 (O_366,N_8886,N_8672);
nand UO_367 (O_367,N_8101,N_8184);
nor UO_368 (O_368,N_9350,N_8212);
and UO_369 (O_369,N_8114,N_9171);
nand UO_370 (O_370,N_9439,N_9569);
or UO_371 (O_371,N_8964,N_9502);
or UO_372 (O_372,N_7633,N_7768);
xnor UO_373 (O_373,N_8138,N_9689);
nor UO_374 (O_374,N_8453,N_7915);
nand UO_375 (O_375,N_9962,N_8439);
and UO_376 (O_376,N_9888,N_8353);
xnor UO_377 (O_377,N_8848,N_9165);
and UO_378 (O_378,N_8475,N_8547);
nor UO_379 (O_379,N_9303,N_8717);
nand UO_380 (O_380,N_9853,N_7920);
and UO_381 (O_381,N_8070,N_8085);
and UO_382 (O_382,N_8733,N_7642);
nand UO_383 (O_383,N_9437,N_9694);
nand UO_384 (O_384,N_8545,N_9307);
nor UO_385 (O_385,N_8265,N_9129);
or UO_386 (O_386,N_8019,N_8743);
and UO_387 (O_387,N_8397,N_8179);
or UO_388 (O_388,N_9754,N_8552);
nand UO_389 (O_389,N_9490,N_9742);
nor UO_390 (O_390,N_9192,N_7855);
or UO_391 (O_391,N_7770,N_8646);
nand UO_392 (O_392,N_8943,N_9221);
nand UO_393 (O_393,N_7816,N_7988);
nand UO_394 (O_394,N_9027,N_9825);
or UO_395 (O_395,N_9282,N_9462);
xnor UO_396 (O_396,N_9716,N_7624);
nand UO_397 (O_397,N_8178,N_9707);
xnor UO_398 (O_398,N_8377,N_7849);
nand UO_399 (O_399,N_9417,N_8580);
and UO_400 (O_400,N_9677,N_7636);
nand UO_401 (O_401,N_7508,N_8035);
and UO_402 (O_402,N_8766,N_7626);
xor UO_403 (O_403,N_9460,N_7672);
or UO_404 (O_404,N_8261,N_8664);
nand UO_405 (O_405,N_7972,N_9161);
and UO_406 (O_406,N_8351,N_9533);
nor UO_407 (O_407,N_8274,N_9812);
xor UO_408 (O_408,N_9932,N_9356);
xnor UO_409 (O_409,N_7914,N_9188);
nand UO_410 (O_410,N_7879,N_9089);
xor UO_411 (O_411,N_8090,N_9755);
nor UO_412 (O_412,N_8625,N_9261);
or UO_413 (O_413,N_9902,N_8158);
nand UO_414 (O_414,N_7659,N_8518);
nand UO_415 (O_415,N_7982,N_8474);
or UO_416 (O_416,N_9443,N_9459);
nand UO_417 (O_417,N_8370,N_8164);
or UO_418 (O_418,N_9749,N_7692);
and UO_419 (O_419,N_8043,N_7960);
and UO_420 (O_420,N_8169,N_9524);
nor UO_421 (O_421,N_8177,N_9336);
xor UO_422 (O_422,N_9537,N_9143);
and UO_423 (O_423,N_9398,N_7897);
nand UO_424 (O_424,N_8724,N_8473);
or UO_425 (O_425,N_7510,N_8250);
nand UO_426 (O_426,N_9056,N_9294);
and UO_427 (O_427,N_8832,N_8269);
and UO_428 (O_428,N_9456,N_9849);
or UO_429 (O_429,N_8927,N_7827);
nand UO_430 (O_430,N_9353,N_9943);
and UO_431 (O_431,N_7590,N_8061);
nor UO_432 (O_432,N_8015,N_9335);
xnor UO_433 (O_433,N_8935,N_9405);
nand UO_434 (O_434,N_8544,N_7989);
nor UO_435 (O_435,N_8060,N_7860);
or UO_436 (O_436,N_9082,N_8151);
and UO_437 (O_437,N_7710,N_9867);
and UO_438 (O_438,N_8510,N_8984);
or UO_439 (O_439,N_8133,N_9378);
or UO_440 (O_440,N_9167,N_8779);
or UO_441 (O_441,N_8857,N_8942);
and UO_442 (O_442,N_8200,N_8687);
and UO_443 (O_443,N_7620,N_8193);
and UO_444 (O_444,N_9262,N_8689);
and UO_445 (O_445,N_8668,N_8381);
xor UO_446 (O_446,N_9879,N_8827);
nor UO_447 (O_447,N_9713,N_7599);
and UO_448 (O_448,N_9931,N_8409);
or UO_449 (O_449,N_7951,N_8627);
and UO_450 (O_450,N_9741,N_8690);
and UO_451 (O_451,N_9407,N_9763);
nor UO_452 (O_452,N_8721,N_9917);
and UO_453 (O_453,N_8709,N_8637);
xnor UO_454 (O_454,N_9843,N_7689);
nand UO_455 (O_455,N_8582,N_8157);
and UO_456 (O_456,N_8662,N_8881);
nor UO_457 (O_457,N_8036,N_9098);
nand UO_458 (O_458,N_9522,N_8322);
or UO_459 (O_459,N_8604,N_8797);
xnor UO_460 (O_460,N_8083,N_8390);
nor UO_461 (O_461,N_8901,N_8804);
nand UO_462 (O_462,N_8679,N_8925);
nand UO_463 (O_463,N_9006,N_8319);
nor UO_464 (O_464,N_9656,N_8123);
nor UO_465 (O_465,N_8301,N_9155);
nor UO_466 (O_466,N_7954,N_7533);
and UO_467 (O_467,N_9570,N_9787);
and UO_468 (O_468,N_9802,N_9100);
nor UO_469 (O_469,N_7766,N_9890);
nor UO_470 (O_470,N_9450,N_8168);
nor UO_471 (O_471,N_8933,N_8183);
nand UO_472 (O_472,N_9036,N_9043);
nor UO_473 (O_473,N_8569,N_7889);
and UO_474 (O_474,N_8227,N_9935);
or UO_475 (O_475,N_9068,N_8052);
xor UO_476 (O_476,N_9973,N_9721);
and UO_477 (O_477,N_8258,N_7787);
nor UO_478 (O_478,N_7729,N_9886);
nand UO_479 (O_479,N_9496,N_9205);
nor UO_480 (O_480,N_8875,N_8022);
nor UO_481 (O_481,N_9848,N_8765);
nand UO_482 (O_482,N_8940,N_7591);
nor UO_483 (O_483,N_7587,N_8057);
or UO_484 (O_484,N_9325,N_7652);
and UO_485 (O_485,N_7835,N_8446);
nor UO_486 (O_486,N_8669,N_9379);
nand UO_487 (O_487,N_9060,N_9331);
nor UO_488 (O_488,N_9092,N_9468);
or UO_489 (O_489,N_7804,N_8417);
or UO_490 (O_490,N_9757,N_9339);
nor UO_491 (O_491,N_8568,N_8355);
and UO_492 (O_492,N_8152,N_9978);
or UO_493 (O_493,N_9466,N_9061);
and UO_494 (O_494,N_9804,N_9206);
nor UO_495 (O_495,N_7993,N_9219);
nand UO_496 (O_496,N_9969,N_8855);
nand UO_497 (O_497,N_9030,N_8289);
nor UO_498 (O_498,N_8858,N_8260);
nor UO_499 (O_499,N_9546,N_8191);
xor UO_500 (O_500,N_7571,N_9444);
nand UO_501 (O_501,N_8188,N_9921);
nor UO_502 (O_502,N_8113,N_9194);
nor UO_503 (O_503,N_9446,N_9788);
and UO_504 (O_504,N_9051,N_9136);
and UO_505 (O_505,N_7578,N_9640);
xnor UO_506 (O_506,N_9224,N_8632);
and UO_507 (O_507,N_9764,N_7730);
and UO_508 (O_508,N_8217,N_8102);
and UO_509 (O_509,N_8368,N_8042);
xor UO_510 (O_510,N_7797,N_8538);
and UO_511 (O_511,N_8283,N_7829);
xnor UO_512 (O_512,N_9730,N_8994);
and UO_513 (O_513,N_9668,N_8142);
nand UO_514 (O_514,N_9368,N_8650);
nand UO_515 (O_515,N_9990,N_8311);
or UO_516 (O_516,N_8838,N_8329);
nor UO_517 (O_517,N_7515,N_7589);
or UO_518 (O_518,N_8091,N_8821);
nor UO_519 (O_519,N_9308,N_9897);
nand UO_520 (O_520,N_9428,N_8203);
xnor UO_521 (O_521,N_7826,N_8530);
or UO_522 (O_522,N_7542,N_8362);
and UO_523 (O_523,N_9292,N_9947);
or UO_524 (O_524,N_8749,N_8758);
and UO_525 (O_525,N_8511,N_9922);
nor UO_526 (O_526,N_9815,N_8973);
or UO_527 (O_527,N_9527,N_8620);
and UO_528 (O_528,N_8469,N_9349);
and UO_529 (O_529,N_9135,N_8734);
nand UO_530 (O_530,N_7612,N_8648);
or UO_531 (O_531,N_9542,N_9107);
or UO_532 (O_532,N_8987,N_9097);
nor UO_533 (O_533,N_7820,N_8098);
or UO_534 (O_534,N_8388,N_9120);
nor UO_535 (O_535,N_7871,N_7980);
nand UO_536 (O_536,N_9382,N_8750);
nand UO_537 (O_537,N_9860,N_7695);
or UO_538 (O_538,N_9651,N_8722);
or UO_539 (O_539,N_9025,N_8556);
and UO_540 (O_540,N_8975,N_7898);
or UO_541 (O_541,N_8520,N_8285);
xor UO_542 (O_542,N_9786,N_9974);
nand UO_543 (O_543,N_9769,N_8497);
and UO_544 (O_544,N_9433,N_8950);
nand UO_545 (O_545,N_9346,N_8968);
or UO_546 (O_546,N_8559,N_9711);
nand UO_547 (O_547,N_9803,N_9560);
and UO_548 (O_548,N_8960,N_8507);
or UO_549 (O_549,N_8484,N_9033);
and UO_550 (O_550,N_7615,N_9085);
and UO_551 (O_551,N_9117,N_8895);
and UO_552 (O_552,N_8834,N_8862);
nor UO_553 (O_553,N_9792,N_8794);
and UO_554 (O_554,N_7720,N_8478);
or UO_555 (O_555,N_7544,N_9997);
and UO_556 (O_556,N_8812,N_8125);
nor UO_557 (O_557,N_7891,N_7704);
nand UO_558 (O_558,N_8589,N_8972);
nand UO_559 (O_559,N_7653,N_9881);
and UO_560 (O_560,N_8919,N_8616);
and UO_561 (O_561,N_7819,N_8529);
xnor UO_562 (O_562,N_7844,N_8118);
or UO_563 (O_563,N_9404,N_8826);
nor UO_564 (O_564,N_8233,N_9957);
xor UO_565 (O_565,N_8276,N_8006);
or UO_566 (O_566,N_8503,N_8932);
or UO_567 (O_567,N_8966,N_8761);
nand UO_568 (O_568,N_8246,N_9223);
nor UO_569 (O_569,N_9553,N_7504);
and UO_570 (O_570,N_8266,N_7756);
or UO_571 (O_571,N_9272,N_9724);
xor UO_572 (O_572,N_9684,N_8600);
and UO_573 (O_573,N_9592,N_8030);
nor UO_574 (O_574,N_7584,N_8198);
or UO_575 (O_575,N_7501,N_7953);
nand UO_576 (O_576,N_7782,N_8712);
nor UO_577 (O_577,N_8146,N_8166);
and UO_578 (O_578,N_9430,N_7530);
or UO_579 (O_579,N_7582,N_7762);
xnor UO_580 (O_580,N_8841,N_8009);
xor UO_581 (O_581,N_8769,N_7691);
xnor UO_582 (O_582,N_7681,N_9806);
or UO_583 (O_583,N_8176,N_9750);
xor UO_584 (O_584,N_9631,N_8818);
nor UO_585 (O_585,N_9185,N_7909);
or UO_586 (O_586,N_7546,N_8720);
or UO_587 (O_587,N_9680,N_7815);
nor UO_588 (O_588,N_9500,N_9387);
and UO_589 (O_589,N_8427,N_9666);
xnor UO_590 (O_590,N_8298,N_8360);
and UO_591 (O_591,N_9514,N_8999);
or UO_592 (O_592,N_7621,N_9029);
xnor UO_593 (O_593,N_8900,N_8467);
or UO_594 (O_594,N_9234,N_8462);
or UO_595 (O_595,N_9478,N_8894);
nor UO_596 (O_596,N_8817,N_7706);
nor UO_597 (O_597,N_9556,N_7675);
nand UO_598 (O_598,N_9157,N_9140);
or UO_599 (O_599,N_8512,N_8003);
or UO_600 (O_600,N_8730,N_8961);
or UO_601 (O_601,N_8930,N_9020);
nor UO_602 (O_602,N_9095,N_9671);
nor UO_603 (O_603,N_9062,N_8525);
nor UO_604 (O_604,N_7777,N_7640);
nor UO_605 (O_605,N_9454,N_8424);
nor UO_606 (O_606,N_9315,N_9550);
or UO_607 (O_607,N_8167,N_7884);
or UO_608 (O_608,N_7812,N_7523);
and UO_609 (O_609,N_9586,N_8686);
xor UO_610 (O_610,N_8195,N_9084);
nand UO_611 (O_611,N_9384,N_7807);
or UO_612 (O_612,N_8746,N_9479);
nor UO_613 (O_613,N_8161,N_9199);
or UO_614 (O_614,N_9751,N_8683);
nand UO_615 (O_615,N_9057,N_7610);
or UO_616 (O_616,N_8577,N_8051);
and UO_617 (O_617,N_8653,N_8137);
nor UO_618 (O_618,N_8341,N_9817);
or UO_619 (O_619,N_9829,N_8074);
nand UO_620 (O_620,N_7677,N_7878);
nand UO_621 (O_621,N_9005,N_8204);
nand UO_622 (O_622,N_9067,N_9328);
or UO_623 (O_623,N_8081,N_8414);
nand UO_624 (O_624,N_9992,N_9723);
or UO_625 (O_625,N_9305,N_7753);
and UO_626 (O_626,N_8947,N_8136);
nand UO_627 (O_627,N_8054,N_8286);
or UO_628 (O_628,N_7703,N_9545);
nand UO_629 (O_629,N_8087,N_8230);
nand UO_630 (O_630,N_8270,N_8952);
or UO_631 (O_631,N_9320,N_7723);
nor UO_632 (O_632,N_8028,N_8007);
xnor UO_633 (O_633,N_7838,N_9780);
nor UO_634 (O_634,N_7987,N_7671);
nand UO_635 (O_635,N_9243,N_8231);
or UO_636 (O_636,N_9000,N_9028);
and UO_637 (O_637,N_8513,N_9258);
xor UO_638 (O_638,N_9797,N_8602);
and UO_639 (O_639,N_9180,N_9064);
nor UO_640 (O_640,N_9604,N_7900);
nor UO_641 (O_641,N_8257,N_7924);
nand UO_642 (O_642,N_8037,N_9153);
nand UO_643 (O_643,N_7538,N_8088);
and UO_644 (O_644,N_8339,N_7606);
or UO_645 (O_645,N_7632,N_9032);
xnor UO_646 (O_646,N_9772,N_9590);
nor UO_647 (O_647,N_8522,N_9276);
or UO_648 (O_648,N_8419,N_9235);
nor UO_649 (O_649,N_7922,N_9429);
xnor UO_650 (O_650,N_9255,N_9436);
or UO_651 (O_651,N_9333,N_8762);
nand UO_652 (O_652,N_9401,N_9365);
nor UO_653 (O_653,N_9783,N_8612);
and UO_654 (O_654,N_8763,N_9495);
or UO_655 (O_655,N_9946,N_8075);
nand UO_656 (O_656,N_8366,N_8252);
or UO_657 (O_657,N_9692,N_9148);
or UO_658 (O_658,N_9170,N_7964);
nand UO_659 (O_659,N_8819,N_8536);
nor UO_660 (O_660,N_7959,N_7529);
and UO_661 (O_661,N_7991,N_8027);
nor UO_662 (O_662,N_8039,N_8249);
or UO_663 (O_663,N_8332,N_7688);
and UO_664 (O_664,N_8931,N_9548);
and UO_665 (O_665,N_8062,N_9214);
nand UO_666 (O_666,N_7870,N_7823);
and UO_667 (O_667,N_8887,N_8608);
or UO_668 (O_668,N_9217,N_9610);
or UO_669 (O_669,N_7676,N_7696);
and UO_670 (O_670,N_7901,N_7518);
or UO_671 (O_671,N_7792,N_7631);
and UO_672 (O_672,N_7645,N_9948);
or UO_673 (O_673,N_8132,N_8745);
or UO_674 (O_674,N_8691,N_9013);
nor UO_675 (O_675,N_7943,N_9452);
nor UO_676 (O_676,N_9112,N_9511);
xor UO_677 (O_677,N_9589,N_8435);
xnor UO_678 (O_678,N_8479,N_9383);
nand UO_679 (O_679,N_9074,N_8149);
nand UO_680 (O_680,N_7798,N_7694);
and UO_681 (O_681,N_8248,N_7776);
nor UO_682 (O_682,N_9240,N_8990);
and UO_683 (O_683,N_8657,N_9820);
and UO_684 (O_684,N_7809,N_8902);
nor UO_685 (O_685,N_8542,N_8238);
nor UO_686 (O_686,N_8917,N_8666);
and UO_687 (O_687,N_7603,N_9766);
nand UO_688 (O_688,N_9939,N_7754);
nand UO_689 (O_689,N_8309,N_7540);
or UO_690 (O_690,N_8674,N_9254);
nor UO_691 (O_691,N_8128,N_9289);
and UO_692 (O_692,N_7534,N_8443);
xnor UO_693 (O_693,N_9597,N_7767);
and UO_694 (O_694,N_8226,N_9938);
nor UO_695 (O_695,N_7958,N_9054);
and UO_696 (O_696,N_9549,N_8129);
or UO_697 (O_697,N_8842,N_9280);
nor UO_698 (O_698,N_9785,N_9964);
xnor UO_699 (O_699,N_8330,N_8463);
or UO_700 (O_700,N_9465,N_9911);
or UO_701 (O_701,N_8444,N_8122);
or UO_702 (O_702,N_8189,N_8912);
nor UO_703 (O_703,N_8992,N_8543);
and UO_704 (O_704,N_9693,N_9210);
xor UO_705 (O_705,N_7548,N_9344);
nand UO_706 (O_706,N_9323,N_7791);
or UO_707 (O_707,N_9715,N_8515);
and UO_708 (O_708,N_7577,N_7936);
or UO_709 (O_709,N_7942,N_8175);
or UO_710 (O_710,N_9087,N_9047);
nor UO_711 (O_711,N_8214,N_7790);
nor UO_712 (O_712,N_7928,N_9253);
xor UO_713 (O_713,N_8140,N_9528);
or UO_714 (O_714,N_8652,N_8585);
nand UO_715 (O_715,N_9994,N_8148);
nor UO_716 (O_716,N_9388,N_9354);
or UO_717 (O_717,N_9337,N_9467);
nor UO_718 (O_718,N_7604,N_9015);
nor UO_719 (O_719,N_7580,N_8725);
and UO_720 (O_720,N_8997,N_9626);
and UO_721 (O_721,N_9874,N_8423);
nand UO_722 (O_722,N_9535,N_8406);
and UO_723 (O_723,N_9960,N_8982);
and UO_724 (O_724,N_7622,N_7660);
xor UO_725 (O_725,N_8859,N_9720);
nor UO_726 (O_726,N_9116,N_9474);
nor UO_727 (O_727,N_7614,N_8793);
nand UO_728 (O_728,N_8660,N_7572);
or UO_729 (O_729,N_8392,N_7658);
or UO_730 (O_730,N_9637,N_9183);
nand UO_731 (O_731,N_7834,N_7619);
nor UO_732 (O_732,N_8410,N_9758);
nand UO_733 (O_733,N_7505,N_8099);
nor UO_734 (O_734,N_8364,N_7930);
nor UO_735 (O_735,N_9854,N_9364);
nor UO_736 (O_736,N_7657,N_7886);
nor UO_737 (O_737,N_9719,N_8342);
and UO_738 (O_738,N_7794,N_9956);
and UO_739 (O_739,N_8649,N_7522);
nand UO_740 (O_740,N_8754,N_8500);
nand UO_741 (O_741,N_8387,N_8631);
or UO_742 (O_742,N_8239,N_9215);
xnor UO_743 (O_743,N_7699,N_9858);
and UO_744 (O_744,N_9998,N_8567);
nor UO_745 (O_745,N_7765,N_9274);
and UO_746 (O_746,N_8934,N_7574);
or UO_747 (O_747,N_9945,N_8541);
and UO_748 (O_748,N_8610,N_7641);
nor UO_749 (O_749,N_9442,N_9127);
or UO_750 (O_750,N_9870,N_8092);
nor UO_751 (O_751,N_9929,N_9164);
or UO_752 (O_752,N_9332,N_8499);
xor UO_753 (O_753,N_9109,N_8334);
nand UO_754 (O_754,N_9317,N_7687);
or UO_755 (O_755,N_8704,N_8046);
nor UO_756 (O_756,N_7757,N_8320);
and UO_757 (O_757,N_7600,N_8049);
and UO_758 (O_758,N_9566,N_8048);
nand UO_759 (O_759,N_9982,N_9739);
or UO_760 (O_760,N_7913,N_8843);
or UO_761 (O_761,N_8803,N_9435);
nor UO_762 (O_762,N_8069,N_8555);
nand UO_763 (O_763,N_9775,N_9389);
nand UO_764 (O_764,N_7840,N_7848);
nor UO_765 (O_765,N_9334,N_9445);
or UO_766 (O_766,N_9189,N_7647);
nand UO_767 (O_767,N_9756,N_8403);
nand UO_768 (O_768,N_7865,N_9782);
nand UO_769 (O_769,N_7883,N_8658);
or UO_770 (O_770,N_9887,N_9923);
or UO_771 (O_771,N_8951,N_9228);
or UO_772 (O_772,N_7910,N_9855);
and UO_773 (O_773,N_8916,N_7561);
and UO_774 (O_774,N_9521,N_9293);
and UO_775 (O_775,N_8018,N_7583);
or UO_776 (O_776,N_9963,N_9778);
or UO_777 (O_777,N_9132,N_8288);
or UO_778 (O_778,N_9830,N_9674);
or UO_779 (O_779,N_9453,N_7511);
nor UO_780 (O_780,N_9319,N_9236);
or UO_781 (O_781,N_7554,N_9145);
xor UO_782 (O_782,N_8874,N_8654);
nor UO_783 (O_783,N_9557,N_7746);
nand UO_784 (O_784,N_9050,N_9665);
and UO_785 (O_785,N_9869,N_7957);
or UO_786 (O_786,N_9638,N_8127);
nand UO_787 (O_787,N_9846,N_8464);
nand UO_788 (O_788,N_7828,N_9989);
nor UO_789 (O_789,N_8741,N_9683);
nor UO_790 (O_790,N_8259,N_8702);
nand UO_791 (O_791,N_8185,N_9925);
xnor UO_792 (O_792,N_8918,N_8592);
and UO_793 (O_793,N_7575,N_9241);
xor UO_794 (O_794,N_8064,N_8344);
nand UO_795 (O_795,N_9661,N_9762);
and UO_796 (O_796,N_7774,N_9781);
nand UO_797 (O_797,N_7596,N_7701);
xor UO_798 (O_798,N_9555,N_8488);
nor UO_799 (O_799,N_9813,N_9377);
and UO_800 (O_800,N_8946,N_9952);
nor UO_801 (O_801,N_8621,N_8877);
nor UO_802 (O_802,N_8824,N_7758);
nor UO_803 (O_803,N_7948,N_9686);
nor UO_804 (O_804,N_9397,N_7662);
nor UO_805 (O_805,N_9412,N_8780);
nand UO_806 (O_806,N_9958,N_8866);
and UO_807 (O_807,N_9172,N_9499);
and UO_808 (O_808,N_7637,N_9936);
and UO_809 (O_809,N_8428,N_9207);
or UO_810 (O_810,N_7693,N_7890);
or UO_811 (O_811,N_8983,N_9023);
nand UO_812 (O_812,N_9369,N_8029);
nand UO_813 (O_813,N_8665,N_8593);
and UO_814 (O_814,N_8736,N_8144);
or UO_815 (O_815,N_9924,N_7560);
and UO_816 (O_816,N_8055,N_8537);
xnor UO_817 (O_817,N_9790,N_8363);
and UO_818 (O_818,N_9530,N_8883);
and UO_819 (O_819,N_9708,N_7506);
and UO_820 (O_820,N_9374,N_9955);
or UO_821 (O_821,N_7836,N_9746);
nand UO_822 (O_822,N_8974,N_9761);
xor UO_823 (O_823,N_7524,N_9414);
nor UO_824 (O_824,N_8328,N_9816);
or UO_825 (O_825,N_7781,N_8784);
nor UO_826 (O_826,N_9128,N_7576);
xor UO_827 (O_827,N_8756,N_9880);
and UO_828 (O_828,N_9996,N_9118);
nor UO_829 (O_829,N_8759,N_9004);
nor UO_830 (O_830,N_9463,N_7863);
and UO_831 (O_831,N_9075,N_8477);
nand UO_832 (O_832,N_8017,N_8375);
or UO_833 (O_833,N_8820,N_8788);
xor UO_834 (O_834,N_8539,N_8483);
xnor UO_835 (O_835,N_7923,N_8579);
nand UO_836 (O_836,N_9077,N_9395);
or UO_837 (O_837,N_8576,N_8044);
or UO_838 (O_838,N_9617,N_8192);
nand UO_839 (O_839,N_8789,N_9114);
or UO_840 (O_840,N_9421,N_7858);
or UO_841 (O_841,N_8626,N_7832);
or UO_842 (O_842,N_8978,N_8038);
and UO_843 (O_843,N_8312,N_9488);
and UO_844 (O_844,N_9838,N_8597);
and UO_845 (O_845,N_8502,N_9669);
nor UO_846 (O_846,N_8562,N_7866);
and UO_847 (O_847,N_9894,N_8767);
xor UO_848 (O_848,N_9275,N_9126);
nand UO_849 (O_849,N_7682,N_8963);
nor UO_850 (O_850,N_7526,N_9260);
nand UO_851 (O_851,N_9302,N_8245);
nor UO_852 (O_852,N_7680,N_8614);
nand UO_853 (O_853,N_9653,N_7679);
nand UO_854 (O_854,N_8041,N_8280);
nand UO_855 (O_855,N_8605,N_8773);
and UO_856 (O_856,N_8981,N_9371);
nand UO_857 (O_857,N_9491,N_9976);
and UO_858 (O_858,N_7712,N_9104);
or UO_859 (O_859,N_9968,N_7850);
nor UO_860 (O_860,N_8065,N_9455);
nand UO_861 (O_861,N_7841,N_8581);
and UO_862 (O_862,N_8365,N_9512);
nand UO_863 (O_863,N_8348,N_7852);
and UO_864 (O_864,N_9083,N_8025);
nand UO_865 (O_865,N_9605,N_9676);
xor UO_866 (O_866,N_9408,N_9264);
or UO_867 (O_867,N_9909,N_8587);
nand UO_868 (O_868,N_8013,N_9663);
and UO_869 (O_869,N_8971,N_9906);
and UO_870 (O_870,N_8760,N_9322);
xnor UO_871 (O_871,N_9279,N_8053);
nand UO_872 (O_872,N_8326,N_9779);
and UO_873 (O_873,N_7971,N_8867);
xnor UO_874 (O_874,N_7661,N_7905);
nand UO_875 (O_875,N_8922,N_9392);
nand UO_876 (O_876,N_8965,N_8523);
or UO_877 (O_877,N_7947,N_8711);
and UO_878 (O_878,N_9691,N_9898);
nor UO_879 (O_879,N_7670,N_8145);
nand UO_880 (O_880,N_8535,N_8159);
nand UO_881 (O_881,N_8263,N_9031);
nand UO_882 (O_882,N_7722,N_8367);
xor UO_883 (O_883,N_9728,N_9580);
or UO_884 (O_884,N_9247,N_9919);
xor UO_885 (O_885,N_7927,N_8954);
and UO_886 (O_886,N_8297,N_8354);
nand UO_887 (O_887,N_8066,N_9914);
nand UO_888 (O_888,N_9142,N_9394);
or UO_889 (O_889,N_8700,N_8835);
xnor UO_890 (O_890,N_8740,N_9102);
nand UO_891 (O_891,N_9249,N_9144);
and UO_892 (O_892,N_8884,N_8107);
nor UO_893 (O_893,N_8490,N_7552);
nand UO_894 (O_894,N_8437,N_9362);
or UO_895 (O_895,N_8744,N_9774);
xor UO_896 (O_896,N_8647,N_8636);
nor UO_897 (O_897,N_9290,N_9633);
nor UO_898 (O_898,N_8575,N_8310);
or UO_899 (O_899,N_9313,N_8277);
or UO_900 (O_900,N_9287,N_7516);
and UO_901 (O_901,N_8988,N_8755);
and UO_902 (O_902,N_9670,N_7537);
or UO_903 (O_903,N_8958,N_9644);
xor UO_904 (O_904,N_9069,N_8656);
nand UO_905 (O_905,N_9748,N_9807);
nor UO_906 (O_906,N_9657,N_8407);
nor UO_907 (O_907,N_9799,N_7918);
and UO_908 (O_908,N_9475,N_8357);
or UO_909 (O_909,N_8565,N_9049);
or UO_910 (O_910,N_7926,N_9158);
nor UO_911 (O_911,N_9551,N_9451);
or UO_912 (O_912,N_9507,N_9438);
or UO_913 (O_913,N_7893,N_8938);
or UO_914 (O_914,N_9823,N_7714);
nor UO_915 (O_915,N_9647,N_7881);
nor UO_916 (O_916,N_7952,N_8798);
nor UO_917 (O_917,N_9003,N_8739);
nor UO_918 (O_918,N_9608,N_8324);
nand UO_919 (O_919,N_8496,N_8861);
nor UO_920 (O_920,N_7607,N_7992);
or UO_921 (O_921,N_8727,N_8639);
and UO_922 (O_922,N_8126,N_8936);
and UO_923 (O_923,N_9498,N_7555);
and UO_924 (O_924,N_8278,N_9800);
and UO_925 (O_925,N_9326,N_9018);
and UO_926 (O_926,N_8482,N_7761);
or UO_927 (O_927,N_9190,N_8893);
or UO_928 (O_928,N_9791,N_9859);
nor UO_929 (O_929,N_9321,N_9675);
nand UO_930 (O_930,N_7685,N_8347);
nand UO_931 (O_931,N_8514,N_8718);
nand UO_932 (O_932,N_9285,N_8854);
nor UO_933 (O_933,N_7968,N_8531);
or UO_934 (O_934,N_9725,N_8659);
and UO_935 (O_935,N_8996,N_9777);
and UO_936 (O_936,N_7985,N_8856);
nand UO_937 (O_937,N_9329,N_8287);
xor UO_938 (O_938,N_9951,N_8209);
xor UO_939 (O_939,N_7527,N_7734);
xnor UO_940 (O_940,N_8208,N_7933);
and UO_941 (O_941,N_9795,N_9679);
and UO_942 (O_942,N_7779,N_7742);
nand UO_943 (O_943,N_9137,N_9151);
and UO_944 (O_944,N_8908,N_9309);
and UO_945 (O_945,N_9538,N_8521);
nand UO_946 (O_946,N_9348,N_9375);
nand UO_947 (O_947,N_9572,N_8201);
or UO_948 (O_948,N_9024,N_8595);
nor UO_949 (O_949,N_9347,N_9805);
and UO_950 (O_950,N_8165,N_9343);
nand UO_951 (O_951,N_8299,N_8190);
nor UO_952 (O_952,N_9481,N_8808);
nor UO_953 (O_953,N_8306,N_8460);
and UO_954 (O_954,N_9411,N_8785);
and UO_955 (O_955,N_8840,N_8955);
or UO_956 (O_956,N_7648,N_8753);
nor UO_957 (O_957,N_7885,N_8956);
nand UO_958 (O_958,N_7941,N_8909);
xnor UO_959 (O_959,N_8268,N_7595);
nand UO_960 (O_960,N_7903,N_8119);
and UO_961 (O_961,N_9230,N_8160);
or UO_962 (O_962,N_9529,N_9310);
xnor UO_963 (O_963,N_9105,N_9372);
nor UO_964 (O_964,N_7793,N_9847);
or UO_965 (O_965,N_9942,N_9086);
nand UO_966 (O_966,N_8452,N_7805);
or UO_967 (O_967,N_9363,N_7545);
and UO_968 (O_968,N_8661,N_8350);
or UO_969 (O_969,N_9615,N_9470);
nand UO_970 (O_970,N_9903,N_7859);
nor UO_971 (O_971,N_9461,N_8369);
nand UO_972 (O_972,N_9612,N_7674);
and UO_973 (O_973,N_9729,N_9912);
xor UO_974 (O_974,N_8723,N_8120);
and UO_975 (O_975,N_8135,N_8571);
and UO_976 (O_976,N_9222,N_7802);
and UO_977 (O_977,N_9182,N_9385);
and UO_978 (O_978,N_8836,N_7986);
nand UO_979 (O_979,N_9704,N_9094);
xnor UO_980 (O_980,N_8047,N_7627);
and UO_981 (O_981,N_8764,N_8599);
nor UO_982 (O_982,N_8897,N_9681);
nand UO_983 (O_983,N_8449,N_8953);
and UO_984 (O_984,N_9268,N_8373);
nor UO_985 (O_985,N_8850,N_8688);
nor UO_986 (O_986,N_9448,N_9423);
and UO_987 (O_987,N_7625,N_8284);
or UO_988 (O_988,N_9983,N_8021);
or UO_989 (O_989,N_9299,N_8606);
nand UO_990 (O_990,N_9237,N_8816);
and UO_991 (O_991,N_8333,N_8617);
xor UO_992 (O_992,N_7976,N_9871);
or UO_993 (O_993,N_8822,N_9351);
nor UO_994 (O_994,N_9596,N_8613);
and UO_995 (O_995,N_8980,N_8677);
and UO_996 (O_996,N_8293,N_9133);
nor UO_997 (O_997,N_8480,N_9516);
xnor UO_998 (O_998,N_9422,N_8358);
nor UO_999 (O_999,N_8495,N_8109);
and UO_1000 (O_1000,N_7724,N_8937);
nand UO_1001 (O_1001,N_9682,N_7711);
or UO_1002 (O_1002,N_8849,N_7520);
nor UO_1003 (O_1003,N_7573,N_8948);
xnor UO_1004 (O_1004,N_8000,N_7778);
xnor UO_1005 (O_1005,N_9044,N_8570);
nand UO_1006 (O_1006,N_9877,N_8121);
or UO_1007 (O_1007,N_9701,N_7531);
xnor UO_1008 (O_1008,N_8020,N_9048);
nor UO_1009 (O_1009,N_8747,N_9352);
nor UO_1010 (O_1010,N_7995,N_8234);
and UO_1011 (O_1011,N_9645,N_9066);
nor UO_1012 (O_1012,N_7944,N_8323);
or UO_1013 (O_1013,N_9581,N_9636);
nor UO_1014 (O_1014,N_9316,N_9941);
nand UO_1015 (O_1015,N_9359,N_9752);
and UO_1016 (O_1016,N_7745,N_9497);
xor UO_1017 (O_1017,N_9471,N_8775);
xor UO_1018 (O_1018,N_9928,N_9432);
and UO_1019 (O_1019,N_9503,N_9175);
nand UO_1020 (O_1020,N_9918,N_7512);
nand UO_1021 (O_1021,N_8267,N_9695);
nand UO_1022 (O_1022,N_9768,N_8111);
nand UO_1023 (O_1023,N_9156,N_8695);
nor UO_1024 (O_1024,N_8546,N_8989);
nor UO_1025 (O_1025,N_9818,N_7663);
nor UO_1026 (O_1026,N_8594,N_9300);
nor UO_1027 (O_1027,N_7716,N_8272);
nor UO_1028 (O_1028,N_8470,N_7517);
nor UO_1029 (O_1029,N_9984,N_7769);
or UO_1030 (O_1030,N_9376,N_9900);
and UO_1031 (O_1031,N_8317,N_9361);
or UO_1032 (O_1032,N_7902,N_8163);
nand UO_1033 (O_1033,N_9191,N_8611);
nor UO_1034 (O_1034,N_8845,N_8633);
nand UO_1035 (O_1035,N_7735,N_8560);
or UO_1036 (O_1036,N_8493,N_8814);
and UO_1037 (O_1037,N_9252,N_9231);
nor UO_1038 (O_1038,N_9896,N_8558);
xnor UO_1039 (O_1039,N_9599,N_7784);
nor UO_1040 (O_1040,N_7973,N_9808);
nor UO_1041 (O_1041,N_9218,N_7801);
and UO_1042 (O_1042,N_7880,N_9598);
nor UO_1043 (O_1043,N_8372,N_9146);
nor UO_1044 (O_1044,N_7629,N_9298);
or UO_1045 (O_1045,N_8117,N_8077);
xor UO_1046 (O_1046,N_9168,N_8872);
nand UO_1047 (O_1047,N_7727,N_9809);
or UO_1048 (O_1048,N_7568,N_9420);
or UO_1049 (O_1049,N_9660,N_9940);
nand UO_1050 (O_1050,N_9893,N_9967);
and UO_1051 (O_1051,N_8262,N_9458);
nand UO_1052 (O_1052,N_8225,N_9277);
or UO_1053 (O_1053,N_8509,N_9273);
and UO_1054 (O_1054,N_7938,N_7543);
and UO_1055 (O_1055,N_8528,N_8670);
nor UO_1056 (O_1056,N_8800,N_9554);
nor UO_1057 (O_1057,N_7581,N_8728);
or UO_1058 (O_1058,N_7919,N_9571);
and UO_1059 (O_1059,N_9627,N_8825);
and UO_1060 (O_1060,N_8335,N_9486);
and UO_1061 (O_1061,N_9415,N_8421);
nand UO_1062 (O_1062,N_9937,N_8642);
nor UO_1063 (O_1063,N_7649,N_9039);
and UO_1064 (O_1064,N_9950,N_7721);
and UO_1065 (O_1065,N_8205,N_8279);
nor UO_1066 (O_1066,N_8110,N_9531);
or UO_1067 (O_1067,N_8489,N_7744);
nor UO_1068 (O_1068,N_8844,N_9543);
or UO_1069 (O_1069,N_9281,N_9169);
and UO_1070 (O_1070,N_9227,N_9393);
xor UO_1071 (O_1071,N_8782,N_9712);
nor UO_1072 (O_1072,N_8434,N_9563);
or UO_1073 (O_1073,N_8828,N_8551);
or UO_1074 (O_1074,N_9096,N_8837);
and UO_1075 (O_1075,N_9341,N_9265);
or UO_1076 (O_1076,N_8706,N_8768);
nor UO_1077 (O_1077,N_8601,N_7916);
or UO_1078 (O_1078,N_9238,N_8459);
and UO_1079 (O_1079,N_8338,N_7547);
or UO_1080 (O_1080,N_9822,N_8680);
or UO_1081 (O_1081,N_8264,N_9573);
nor UO_1082 (O_1082,N_9594,N_8374);
nor UO_1083 (O_1083,N_9409,N_9593);
and UO_1084 (O_1084,N_7750,N_8186);
xnor UO_1085 (O_1085,N_9327,N_8729);
nand UO_1086 (O_1086,N_7862,N_7708);
nand UO_1087 (O_1087,N_8139,N_7623);
nand UO_1088 (O_1088,N_7743,N_9200);
or UO_1089 (O_1089,N_8792,N_8910);
xnor UO_1090 (O_1090,N_9266,N_7929);
xnor UO_1091 (O_1091,N_8923,N_8296);
nand UO_1092 (O_1092,N_9134,N_9833);
or UO_1093 (O_1093,N_9108,N_9688);
or UO_1094 (O_1094,N_9026,N_7861);
nand UO_1095 (O_1095,N_9440,N_9995);
nor UO_1096 (O_1096,N_8404,N_9402);
nor UO_1097 (O_1097,N_9123,N_7810);
nand UO_1098 (O_1098,N_8401,N_7567);
nor UO_1099 (O_1099,N_9568,N_8093);
nor UO_1100 (O_1100,N_7837,N_7990);
xnor UO_1101 (O_1101,N_9798,N_7868);
nand UO_1102 (O_1102,N_8451,N_9525);
xor UO_1103 (O_1103,N_9239,N_9717);
nand UO_1104 (O_1104,N_9038,N_8194);
and UO_1105 (O_1105,N_8508,N_8413);
nand UO_1106 (O_1106,N_9814,N_8063);
and UO_1107 (O_1107,N_8181,N_9131);
or UO_1108 (O_1108,N_8100,N_7519);
nor UO_1109 (O_1109,N_9685,N_9534);
nor UO_1110 (O_1110,N_9464,N_8880);
nor UO_1111 (O_1111,N_9587,N_9070);
nand UO_1112 (O_1112,N_9662,N_8130);
or UO_1113 (O_1113,N_9642,N_9913);
or UO_1114 (O_1114,N_9700,N_9953);
xor UO_1115 (O_1115,N_9141,N_9834);
nor UO_1116 (O_1116,N_9826,N_8218);
nand UO_1117 (O_1117,N_7939,N_8795);
nand UO_1118 (O_1118,N_9811,N_7513);
and UO_1119 (O_1119,N_8220,N_9747);
nand UO_1120 (O_1120,N_8732,N_9641);
and UO_1121 (O_1121,N_9053,N_8108);
xnor UO_1122 (O_1122,N_9773,N_9357);
nor UO_1123 (O_1123,N_8487,N_9058);
nor UO_1124 (O_1124,N_8008,N_9993);
or UO_1125 (O_1125,N_9010,N_9926);
nand UO_1126 (O_1126,N_9579,N_7586);
nand UO_1127 (O_1127,N_9301,N_7713);
nand UO_1128 (O_1128,N_7536,N_8752);
or UO_1129 (O_1129,N_9447,N_9209);
or UO_1130 (O_1130,N_8864,N_8429);
nand UO_1131 (O_1131,N_9831,N_8224);
and UO_1132 (O_1132,N_9620,N_7821);
nand UO_1133 (O_1133,N_9021,N_8134);
or UO_1134 (O_1134,N_8196,N_9366);
nand UO_1135 (O_1135,N_9703,N_9492);
nand UO_1136 (O_1136,N_8112,N_9270);
nor UO_1137 (O_1137,N_7557,N_8461);
nor UO_1138 (O_1138,N_9934,N_8304);
nand UO_1139 (O_1139,N_9954,N_7842);
and UO_1140 (O_1140,N_8173,N_8072);
and UO_1141 (O_1141,N_7550,N_8863);
nor UO_1142 (O_1142,N_9629,N_9119);
xnor UO_1143 (O_1143,N_8026,N_9113);
or UO_1144 (O_1144,N_9476,N_9482);
or UO_1145 (O_1145,N_9578,N_8641);
and UO_1146 (O_1146,N_8635,N_8001);
nand UO_1147 (O_1147,N_7549,N_8210);
nor UO_1148 (O_1148,N_9646,N_9034);
nand UO_1149 (O_1149,N_8506,N_8748);
nor UO_1150 (O_1150,N_9667,N_9575);
nand UO_1151 (O_1151,N_9842,N_7605);
nand UO_1152 (O_1152,N_8316,N_8699);
or UO_1153 (O_1153,N_8498,N_8071);
xnor UO_1154 (O_1154,N_7705,N_7946);
and UO_1155 (O_1155,N_7795,N_8422);
nand UO_1156 (O_1156,N_8527,N_9949);
nor UO_1157 (O_1157,N_8255,N_8251);
and UO_1158 (O_1158,N_8876,N_7803);
nor UO_1159 (O_1159,N_8150,N_9342);
and UO_1160 (O_1160,N_8885,N_8517);
nand UO_1161 (O_1161,N_8466,N_8831);
nand UO_1162 (O_1162,N_9518,N_7853);
nand UO_1163 (O_1163,N_7833,N_8032);
or UO_1164 (O_1164,N_7655,N_7646);
nand UO_1165 (O_1165,N_8336,N_9564);
nand UO_1166 (O_1166,N_9622,N_9840);
nand UO_1167 (O_1167,N_9519,N_8791);
nand UO_1168 (O_1168,N_8386,N_9861);
and UO_1169 (O_1169,N_7749,N_9360);
and UO_1170 (O_1170,N_9487,N_8216);
nand UO_1171 (O_1171,N_7700,N_8004);
or UO_1172 (O_1172,N_9654,N_9011);
and UO_1173 (O_1173,N_8889,N_9139);
or UO_1174 (O_1174,N_8939,N_8011);
or UO_1175 (O_1175,N_8783,N_8870);
nor UO_1176 (O_1176,N_8059,N_9370);
or UO_1177 (O_1177,N_9864,N_9944);
nand UO_1178 (O_1178,N_9211,N_8432);
or UO_1179 (O_1179,N_9162,N_8913);
nand UO_1180 (O_1180,N_8655,N_9619);
xor UO_1181 (O_1181,N_8229,N_8103);
and UO_1182 (O_1182,N_9233,N_9111);
or UO_1183 (O_1183,N_7932,N_7983);
and UO_1184 (O_1184,N_8860,N_7564);
nor UO_1185 (O_1185,N_7738,N_9019);
nor UO_1186 (O_1186,N_9595,N_8197);
nor UO_1187 (O_1187,N_9494,N_8045);
nor UO_1188 (O_1188,N_8187,N_7528);
and UO_1189 (O_1189,N_8598,N_8331);
nor UO_1190 (O_1190,N_9532,N_8447);
xor UO_1191 (O_1191,N_9286,N_7979);
nor UO_1192 (O_1192,N_8967,N_9583);
and UO_1193 (O_1193,N_9469,N_7690);
xnor UO_1194 (O_1194,N_9609,N_9059);
xor UO_1195 (O_1195,N_7981,N_7888);
and UO_1196 (O_1196,N_8327,N_9291);
and UO_1197 (O_1197,N_7978,N_9063);
and UO_1198 (O_1198,N_9618,N_8202);
and UO_1199 (O_1199,N_9714,N_9173);
and UO_1200 (O_1200,N_9208,N_7857);
nor UO_1201 (O_1201,N_8735,N_9130);
xor UO_1202 (O_1202,N_7912,N_9767);
nor UO_1203 (O_1203,N_8172,N_9999);
xnor UO_1204 (O_1204,N_8623,N_8067);
and UO_1205 (O_1205,N_7709,N_9295);
nand UO_1206 (O_1206,N_7628,N_8731);
nor UO_1207 (O_1207,N_9220,N_9154);
or UO_1208 (O_1208,N_8254,N_7963);
or UO_1209 (O_1209,N_9699,N_9008);
nor UO_1210 (O_1210,N_7817,N_8697);
xnor UO_1211 (O_1211,N_7962,N_9577);
nor UO_1212 (O_1212,N_8959,N_8399);
nand UO_1213 (O_1213,N_8696,N_9745);
nand UO_1214 (O_1214,N_9103,N_8678);
or UO_1215 (O_1215,N_8012,N_9737);
nor UO_1216 (O_1216,N_7874,N_8698);
nor UO_1217 (O_1217,N_7877,N_9072);
nor UO_1218 (O_1218,N_8757,N_9889);
and UO_1219 (O_1219,N_7799,N_8050);
and UO_1220 (O_1220,N_8273,N_8236);
or UO_1221 (O_1221,N_9042,N_7759);
xor UO_1222 (O_1222,N_9022,N_9418);
nand UO_1223 (O_1223,N_8213,N_9789);
nand UO_1224 (O_1224,N_7562,N_8682);
xnor UO_1225 (O_1225,N_9852,N_7728);
and UO_1226 (O_1226,N_9832,N_9862);
or UO_1227 (O_1227,N_9410,N_7731);
nand UO_1228 (O_1228,N_8408,N_9526);
nor UO_1229 (O_1229,N_9016,N_8519);
nor UO_1230 (O_1230,N_7873,N_9987);
and UO_1231 (O_1231,N_7937,N_8440);
nand UO_1232 (O_1232,N_9845,N_8106);
xnor UO_1233 (O_1233,N_7967,N_9561);
and UO_1234 (O_1234,N_8222,N_7887);
xor UO_1235 (O_1235,N_8147,N_9419);
and UO_1236 (O_1236,N_8684,N_9358);
nand UO_1237 (O_1237,N_8738,N_9616);
and UO_1238 (O_1238,N_8847,N_8945);
nand UO_1239 (O_1239,N_9257,N_8340);
and UO_1240 (O_1240,N_8928,N_9625);
nor UO_1241 (O_1241,N_8532,N_9330);
nand UO_1242 (O_1242,N_8418,N_9698);
xnor UO_1243 (O_1243,N_7503,N_8346);
nor UO_1244 (O_1244,N_9427,N_7830);
or UO_1245 (O_1245,N_8402,N_8485);
nor UO_1246 (O_1246,N_9760,N_7772);
nand UO_1247 (O_1247,N_9150,N_8476);
or UO_1248 (O_1248,N_9839,N_7748);
and UO_1249 (O_1249,N_8105,N_8282);
nand UO_1250 (O_1250,N_9626,N_8562);
nand UO_1251 (O_1251,N_9703,N_7676);
nor UO_1252 (O_1252,N_8698,N_8479);
nor UO_1253 (O_1253,N_7621,N_9188);
and UO_1254 (O_1254,N_8794,N_8411);
nor UO_1255 (O_1255,N_9262,N_7523);
or UO_1256 (O_1256,N_8349,N_8794);
nand UO_1257 (O_1257,N_9153,N_9799);
nor UO_1258 (O_1258,N_8419,N_8047);
or UO_1259 (O_1259,N_9335,N_8602);
nand UO_1260 (O_1260,N_9647,N_9604);
xnor UO_1261 (O_1261,N_9113,N_8262);
and UO_1262 (O_1262,N_9635,N_7705);
or UO_1263 (O_1263,N_8512,N_7766);
xor UO_1264 (O_1264,N_8434,N_9896);
nand UO_1265 (O_1265,N_8963,N_8776);
or UO_1266 (O_1266,N_8538,N_9380);
nor UO_1267 (O_1267,N_7996,N_8439);
nor UO_1268 (O_1268,N_8732,N_8784);
and UO_1269 (O_1269,N_8379,N_8777);
and UO_1270 (O_1270,N_7806,N_7998);
nand UO_1271 (O_1271,N_7994,N_8270);
or UO_1272 (O_1272,N_8483,N_9937);
and UO_1273 (O_1273,N_8882,N_8633);
nor UO_1274 (O_1274,N_8963,N_8855);
nand UO_1275 (O_1275,N_9965,N_8402);
and UO_1276 (O_1276,N_9455,N_8069);
and UO_1277 (O_1277,N_7795,N_8040);
or UO_1278 (O_1278,N_9981,N_8368);
nor UO_1279 (O_1279,N_8759,N_8875);
xnor UO_1280 (O_1280,N_8377,N_8790);
nand UO_1281 (O_1281,N_8363,N_8385);
or UO_1282 (O_1282,N_8774,N_8415);
xnor UO_1283 (O_1283,N_9168,N_7920);
nor UO_1284 (O_1284,N_9785,N_7907);
or UO_1285 (O_1285,N_7838,N_9171);
or UO_1286 (O_1286,N_8130,N_8733);
or UO_1287 (O_1287,N_7859,N_9569);
and UO_1288 (O_1288,N_7693,N_9674);
xnor UO_1289 (O_1289,N_8213,N_9100);
xnor UO_1290 (O_1290,N_7753,N_8186);
and UO_1291 (O_1291,N_9721,N_9256);
or UO_1292 (O_1292,N_8446,N_9370);
or UO_1293 (O_1293,N_9520,N_7568);
or UO_1294 (O_1294,N_7670,N_9385);
nor UO_1295 (O_1295,N_9313,N_8660);
or UO_1296 (O_1296,N_9172,N_8928);
or UO_1297 (O_1297,N_9086,N_8268);
nand UO_1298 (O_1298,N_9698,N_8570);
nand UO_1299 (O_1299,N_8296,N_8784);
nand UO_1300 (O_1300,N_8521,N_9204);
or UO_1301 (O_1301,N_8473,N_9937);
and UO_1302 (O_1302,N_8226,N_8062);
nor UO_1303 (O_1303,N_7588,N_8833);
or UO_1304 (O_1304,N_9143,N_7506);
and UO_1305 (O_1305,N_8517,N_9157);
or UO_1306 (O_1306,N_7799,N_7733);
nor UO_1307 (O_1307,N_8985,N_9419);
xnor UO_1308 (O_1308,N_8479,N_8055);
or UO_1309 (O_1309,N_9255,N_8214);
or UO_1310 (O_1310,N_9614,N_9684);
xnor UO_1311 (O_1311,N_9226,N_8022);
and UO_1312 (O_1312,N_8904,N_7729);
nand UO_1313 (O_1313,N_9218,N_9256);
or UO_1314 (O_1314,N_8151,N_7898);
nand UO_1315 (O_1315,N_8083,N_8697);
or UO_1316 (O_1316,N_7855,N_7860);
or UO_1317 (O_1317,N_9190,N_9768);
xnor UO_1318 (O_1318,N_9980,N_9951);
and UO_1319 (O_1319,N_8516,N_8049);
and UO_1320 (O_1320,N_7849,N_9457);
or UO_1321 (O_1321,N_9662,N_7917);
or UO_1322 (O_1322,N_9268,N_8990);
nor UO_1323 (O_1323,N_9139,N_9208);
nand UO_1324 (O_1324,N_8535,N_9653);
or UO_1325 (O_1325,N_9661,N_8784);
nand UO_1326 (O_1326,N_9919,N_8560);
or UO_1327 (O_1327,N_9050,N_8166);
and UO_1328 (O_1328,N_8408,N_8061);
or UO_1329 (O_1329,N_8167,N_8082);
or UO_1330 (O_1330,N_7868,N_7698);
and UO_1331 (O_1331,N_7953,N_9212);
xor UO_1332 (O_1332,N_9277,N_8161);
and UO_1333 (O_1333,N_8436,N_8431);
xnor UO_1334 (O_1334,N_8135,N_8640);
nand UO_1335 (O_1335,N_8986,N_9272);
and UO_1336 (O_1336,N_8827,N_8214);
and UO_1337 (O_1337,N_9080,N_8869);
nor UO_1338 (O_1338,N_8692,N_8481);
and UO_1339 (O_1339,N_8119,N_9301);
nand UO_1340 (O_1340,N_8281,N_8361);
and UO_1341 (O_1341,N_8950,N_9020);
and UO_1342 (O_1342,N_8047,N_9358);
and UO_1343 (O_1343,N_9933,N_9193);
or UO_1344 (O_1344,N_7977,N_9755);
and UO_1345 (O_1345,N_8753,N_8441);
nand UO_1346 (O_1346,N_8805,N_8579);
nand UO_1347 (O_1347,N_8224,N_7695);
and UO_1348 (O_1348,N_8661,N_9390);
and UO_1349 (O_1349,N_8315,N_8456);
nand UO_1350 (O_1350,N_8976,N_8571);
and UO_1351 (O_1351,N_8683,N_7673);
xnor UO_1352 (O_1352,N_8535,N_8636);
nand UO_1353 (O_1353,N_8290,N_8604);
nand UO_1354 (O_1354,N_7757,N_8694);
nand UO_1355 (O_1355,N_9777,N_9800);
or UO_1356 (O_1356,N_7872,N_9221);
nor UO_1357 (O_1357,N_9623,N_8359);
or UO_1358 (O_1358,N_7644,N_8720);
and UO_1359 (O_1359,N_9897,N_9301);
and UO_1360 (O_1360,N_9609,N_9221);
nor UO_1361 (O_1361,N_9954,N_8700);
nand UO_1362 (O_1362,N_9512,N_8631);
nor UO_1363 (O_1363,N_8188,N_9852);
nand UO_1364 (O_1364,N_8910,N_9517);
and UO_1365 (O_1365,N_8954,N_8397);
and UO_1366 (O_1366,N_8838,N_8064);
nand UO_1367 (O_1367,N_8613,N_7709);
xor UO_1368 (O_1368,N_8904,N_9997);
nand UO_1369 (O_1369,N_9485,N_7622);
xor UO_1370 (O_1370,N_7667,N_8640);
nand UO_1371 (O_1371,N_8862,N_7848);
or UO_1372 (O_1372,N_8141,N_9477);
nand UO_1373 (O_1373,N_9562,N_8377);
nor UO_1374 (O_1374,N_7971,N_8171);
nor UO_1375 (O_1375,N_8787,N_9466);
nand UO_1376 (O_1376,N_7696,N_8362);
xnor UO_1377 (O_1377,N_7937,N_8567);
nor UO_1378 (O_1378,N_8653,N_9168);
nor UO_1379 (O_1379,N_9045,N_7525);
and UO_1380 (O_1380,N_9175,N_9594);
nand UO_1381 (O_1381,N_9382,N_7672);
or UO_1382 (O_1382,N_9797,N_9236);
xor UO_1383 (O_1383,N_8218,N_8000);
nor UO_1384 (O_1384,N_8379,N_9443);
nand UO_1385 (O_1385,N_8672,N_8352);
nor UO_1386 (O_1386,N_9067,N_8920);
or UO_1387 (O_1387,N_9720,N_9651);
nor UO_1388 (O_1388,N_9287,N_9189);
nor UO_1389 (O_1389,N_8175,N_9801);
or UO_1390 (O_1390,N_8111,N_8460);
or UO_1391 (O_1391,N_9423,N_8092);
nor UO_1392 (O_1392,N_8734,N_8604);
nor UO_1393 (O_1393,N_9568,N_9311);
and UO_1394 (O_1394,N_8940,N_8377);
xor UO_1395 (O_1395,N_8199,N_8979);
nand UO_1396 (O_1396,N_9954,N_9686);
or UO_1397 (O_1397,N_8852,N_8138);
nand UO_1398 (O_1398,N_9566,N_7682);
nand UO_1399 (O_1399,N_9669,N_9953);
or UO_1400 (O_1400,N_8221,N_8365);
nor UO_1401 (O_1401,N_9198,N_7730);
nand UO_1402 (O_1402,N_9234,N_7816);
nor UO_1403 (O_1403,N_8203,N_9865);
or UO_1404 (O_1404,N_8238,N_9914);
xnor UO_1405 (O_1405,N_8650,N_9435);
nor UO_1406 (O_1406,N_7894,N_7741);
or UO_1407 (O_1407,N_9690,N_7881);
and UO_1408 (O_1408,N_9790,N_7984);
or UO_1409 (O_1409,N_9762,N_9894);
and UO_1410 (O_1410,N_8662,N_8242);
or UO_1411 (O_1411,N_8435,N_8578);
xnor UO_1412 (O_1412,N_8468,N_8475);
xnor UO_1413 (O_1413,N_9622,N_7631);
or UO_1414 (O_1414,N_8344,N_8945);
or UO_1415 (O_1415,N_9016,N_8212);
nor UO_1416 (O_1416,N_8523,N_9935);
and UO_1417 (O_1417,N_8287,N_9398);
nand UO_1418 (O_1418,N_9122,N_9497);
and UO_1419 (O_1419,N_8625,N_9021);
or UO_1420 (O_1420,N_9865,N_9028);
xor UO_1421 (O_1421,N_8352,N_9644);
xor UO_1422 (O_1422,N_9973,N_9788);
and UO_1423 (O_1423,N_7967,N_9537);
or UO_1424 (O_1424,N_7696,N_7595);
nand UO_1425 (O_1425,N_9783,N_7689);
or UO_1426 (O_1426,N_7918,N_8782);
nor UO_1427 (O_1427,N_8452,N_9105);
or UO_1428 (O_1428,N_9850,N_9952);
nand UO_1429 (O_1429,N_8483,N_9517);
nor UO_1430 (O_1430,N_9599,N_9786);
nand UO_1431 (O_1431,N_8382,N_7607);
or UO_1432 (O_1432,N_9579,N_7997);
nor UO_1433 (O_1433,N_7942,N_9817);
nand UO_1434 (O_1434,N_9117,N_8082);
xnor UO_1435 (O_1435,N_8207,N_8189);
and UO_1436 (O_1436,N_9232,N_8159);
nor UO_1437 (O_1437,N_9670,N_8851);
and UO_1438 (O_1438,N_7967,N_8169);
xor UO_1439 (O_1439,N_8686,N_8585);
or UO_1440 (O_1440,N_9521,N_8831);
nand UO_1441 (O_1441,N_8893,N_8797);
xnor UO_1442 (O_1442,N_9135,N_9392);
nand UO_1443 (O_1443,N_8312,N_9970);
nand UO_1444 (O_1444,N_9799,N_9069);
xnor UO_1445 (O_1445,N_9723,N_9442);
nand UO_1446 (O_1446,N_8527,N_8090);
and UO_1447 (O_1447,N_9246,N_9381);
nand UO_1448 (O_1448,N_8306,N_8020);
and UO_1449 (O_1449,N_9252,N_9261);
nor UO_1450 (O_1450,N_8737,N_9244);
nor UO_1451 (O_1451,N_9596,N_9238);
nor UO_1452 (O_1452,N_9521,N_9944);
nand UO_1453 (O_1453,N_9764,N_9419);
nor UO_1454 (O_1454,N_8490,N_8419);
nand UO_1455 (O_1455,N_8956,N_9514);
nor UO_1456 (O_1456,N_9763,N_9310);
or UO_1457 (O_1457,N_7864,N_8330);
nor UO_1458 (O_1458,N_7646,N_8531);
and UO_1459 (O_1459,N_8478,N_8834);
nand UO_1460 (O_1460,N_9297,N_8950);
nor UO_1461 (O_1461,N_9570,N_9745);
and UO_1462 (O_1462,N_7655,N_8259);
or UO_1463 (O_1463,N_8441,N_9068);
nand UO_1464 (O_1464,N_7516,N_9722);
nand UO_1465 (O_1465,N_8882,N_9782);
nor UO_1466 (O_1466,N_9652,N_7923);
and UO_1467 (O_1467,N_9896,N_9477);
xor UO_1468 (O_1468,N_9468,N_8593);
xor UO_1469 (O_1469,N_8653,N_7663);
or UO_1470 (O_1470,N_8012,N_9300);
or UO_1471 (O_1471,N_8171,N_9571);
and UO_1472 (O_1472,N_9706,N_9231);
and UO_1473 (O_1473,N_8256,N_8524);
nor UO_1474 (O_1474,N_8375,N_8850);
and UO_1475 (O_1475,N_9702,N_8049);
nand UO_1476 (O_1476,N_7793,N_7814);
nand UO_1477 (O_1477,N_9416,N_8745);
nand UO_1478 (O_1478,N_8643,N_9444);
nand UO_1479 (O_1479,N_7673,N_7983);
nor UO_1480 (O_1480,N_7839,N_8647);
and UO_1481 (O_1481,N_8532,N_7659);
and UO_1482 (O_1482,N_9049,N_8920);
and UO_1483 (O_1483,N_8505,N_7954);
or UO_1484 (O_1484,N_7971,N_8596);
nor UO_1485 (O_1485,N_8854,N_9196);
xnor UO_1486 (O_1486,N_9715,N_7614);
nor UO_1487 (O_1487,N_8853,N_8730);
or UO_1488 (O_1488,N_8436,N_9158);
nor UO_1489 (O_1489,N_9309,N_8915);
and UO_1490 (O_1490,N_9392,N_8015);
and UO_1491 (O_1491,N_8129,N_9574);
nor UO_1492 (O_1492,N_7940,N_8829);
and UO_1493 (O_1493,N_9412,N_8464);
nor UO_1494 (O_1494,N_8500,N_8540);
and UO_1495 (O_1495,N_8069,N_8771);
xnor UO_1496 (O_1496,N_9957,N_7852);
or UO_1497 (O_1497,N_9039,N_7979);
xnor UO_1498 (O_1498,N_9239,N_9675);
nand UO_1499 (O_1499,N_9827,N_8064);
endmodule