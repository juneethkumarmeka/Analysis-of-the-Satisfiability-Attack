module basic_1000_10000_1500_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_328,In_710);
and U1 (N_1,In_331,In_768);
and U2 (N_2,In_152,In_442);
nand U3 (N_3,In_717,In_953);
or U4 (N_4,In_956,In_410);
nand U5 (N_5,In_870,In_0);
and U6 (N_6,In_705,In_25);
nor U7 (N_7,In_608,In_995);
nand U8 (N_8,In_336,In_718);
nand U9 (N_9,In_851,In_888);
nor U10 (N_10,In_637,In_862);
nor U11 (N_11,In_639,In_631);
or U12 (N_12,In_855,In_940);
or U13 (N_13,In_651,In_313);
nor U14 (N_14,In_93,In_353);
and U15 (N_15,In_865,In_699);
nand U16 (N_16,In_561,In_920);
nor U17 (N_17,In_443,In_278);
and U18 (N_18,In_601,In_648);
nand U19 (N_19,In_885,In_293);
nand U20 (N_20,In_74,In_149);
xnor U21 (N_21,In_505,In_416);
and U22 (N_22,In_986,In_875);
nand U23 (N_23,In_943,In_967);
and U24 (N_24,In_607,In_213);
and U25 (N_25,In_635,In_736);
nor U26 (N_26,In_473,In_581);
nor U27 (N_27,In_341,In_950);
xnor U28 (N_28,In_951,In_26);
and U29 (N_29,In_909,In_167);
nor U30 (N_30,In_32,In_810);
nor U31 (N_31,In_729,In_179);
xor U32 (N_32,In_738,In_51);
nand U33 (N_33,In_873,In_627);
nand U34 (N_34,In_241,In_735);
xnor U35 (N_35,In_886,In_869);
nor U36 (N_36,In_252,In_982);
or U37 (N_37,In_515,In_551);
or U38 (N_38,In_359,In_333);
or U39 (N_39,In_948,In_508);
or U40 (N_40,In_526,In_579);
xor U41 (N_41,In_570,In_260);
or U42 (N_42,In_843,In_759);
nand U43 (N_43,In_461,In_67);
and U44 (N_44,In_853,In_249);
and U45 (N_45,In_709,In_617);
nor U46 (N_46,In_357,In_619);
nor U47 (N_47,In_449,In_225);
or U48 (N_48,In_676,In_457);
nand U49 (N_49,In_644,In_527);
nand U50 (N_50,In_118,In_86);
and U51 (N_51,In_406,In_592);
nand U52 (N_52,In_949,In_266);
xor U53 (N_53,In_150,In_606);
or U54 (N_54,In_616,In_75);
xnor U55 (N_55,In_689,In_966);
nand U56 (N_56,In_731,In_395);
nor U57 (N_57,In_444,In_196);
and U58 (N_58,In_254,In_866);
nand U59 (N_59,In_403,In_40);
and U60 (N_60,In_976,In_311);
and U61 (N_61,In_732,In_351);
or U62 (N_62,In_224,In_884);
nor U63 (N_63,In_271,In_358);
and U64 (N_64,In_912,In_952);
nand U65 (N_65,In_115,In_761);
and U66 (N_66,In_987,In_455);
xnor U67 (N_67,In_911,In_737);
xnor U68 (N_68,In_845,In_256);
nor U69 (N_69,In_429,In_823);
and U70 (N_70,In_286,In_90);
xnor U71 (N_71,In_273,In_100);
and U72 (N_72,In_202,In_335);
and U73 (N_73,In_261,In_70);
and U74 (N_74,In_301,In_168);
nor U75 (N_75,In_84,In_435);
and U76 (N_76,In_785,In_136);
or U77 (N_77,In_874,In_274);
nor U78 (N_78,In_483,In_18);
xor U79 (N_79,In_926,In_962);
and U80 (N_80,In_813,In_691);
xor U81 (N_81,In_33,In_656);
nand U82 (N_82,In_897,In_695);
xnor U83 (N_83,In_312,In_275);
and U84 (N_84,In_277,In_575);
xnor U85 (N_85,In_503,In_568);
xor U86 (N_86,In_177,In_172);
xnor U87 (N_87,In_753,In_822);
nand U88 (N_88,In_125,In_409);
nand U89 (N_89,In_217,In_445);
xnor U90 (N_90,In_584,In_158);
nand U91 (N_91,In_187,In_582);
and U92 (N_92,In_838,In_829);
or U93 (N_93,In_757,In_789);
xor U94 (N_94,In_56,In_560);
and U95 (N_95,In_433,In_268);
nand U96 (N_96,In_660,In_11);
and U97 (N_97,In_999,In_478);
nor U98 (N_98,In_858,In_216);
nand U99 (N_99,In_803,In_818);
xor U100 (N_100,In_151,In_265);
nor U101 (N_101,In_657,In_441);
and U102 (N_102,In_519,In_776);
or U103 (N_103,In_38,In_348);
nand U104 (N_104,In_628,In_383);
nor U105 (N_105,In_22,In_552);
nand U106 (N_106,In_233,In_758);
nand U107 (N_107,In_369,In_272);
xnor U108 (N_108,In_330,In_332);
and U109 (N_109,In_234,In_477);
or U110 (N_110,In_91,In_377);
xor U111 (N_111,In_209,In_345);
or U112 (N_112,In_462,In_605);
and U113 (N_113,In_509,In_498);
xor U114 (N_114,In_747,In_493);
or U115 (N_115,In_47,In_390);
and U116 (N_116,In_960,In_513);
and U117 (N_117,In_825,In_176);
xnor U118 (N_118,In_546,In_918);
xnor U119 (N_119,In_629,In_89);
nand U120 (N_120,In_915,In_380);
xnor U121 (N_121,In_171,In_255);
and U122 (N_122,In_205,In_147);
and U123 (N_123,In_430,In_37);
nor U124 (N_124,In_304,In_859);
nand U125 (N_125,In_517,In_440);
or U126 (N_126,In_368,In_935);
and U127 (N_127,In_895,In_454);
or U128 (N_128,In_308,In_901);
and U129 (N_129,In_913,In_385);
xnor U130 (N_130,In_835,In_655);
or U131 (N_131,In_796,In_63);
and U132 (N_132,In_238,In_214);
nand U133 (N_133,In_733,In_883);
nand U134 (N_134,In_700,In_334);
xnor U135 (N_135,In_134,In_578);
nand U136 (N_136,In_887,In_159);
xnor U137 (N_137,In_270,In_931);
nand U138 (N_138,In_1,In_276);
xnor U139 (N_139,In_927,In_95);
and U140 (N_140,In_237,In_46);
or U141 (N_141,In_882,In_683);
or U142 (N_142,In_425,In_791);
nand U143 (N_143,In_751,In_370);
and U144 (N_144,In_231,In_564);
or U145 (N_145,In_872,In_479);
and U146 (N_146,In_364,In_77);
and U147 (N_147,In_300,In_566);
nand U148 (N_148,In_191,In_8);
and U149 (N_149,In_988,In_557);
and U150 (N_150,In_499,In_230);
nand U151 (N_151,In_156,In_76);
and U152 (N_152,In_878,In_393);
xor U153 (N_153,In_431,In_958);
and U154 (N_154,In_981,In_208);
nor U155 (N_155,In_730,In_48);
nor U156 (N_156,In_204,In_421);
and U157 (N_157,In_316,In_830);
xnor U158 (N_158,In_668,In_924);
and U159 (N_159,In_685,In_131);
nor U160 (N_160,In_399,In_120);
nand U161 (N_161,In_108,In_130);
xnor U162 (N_162,In_674,In_57);
nand U163 (N_163,In_554,In_763);
nand U164 (N_164,In_98,In_414);
nor U165 (N_165,In_137,In_725);
nand U166 (N_166,In_540,In_665);
and U167 (N_167,In_2,In_30);
or U168 (N_168,In_867,In_921);
xnor U169 (N_169,In_583,In_60);
nor U170 (N_170,In_715,In_68);
or U171 (N_171,In_959,In_232);
and U172 (N_172,In_6,In_752);
nor U173 (N_173,In_460,In_365);
or U174 (N_174,In_597,In_437);
or U175 (N_175,In_24,In_847);
xnor U176 (N_176,In_910,In_684);
xor U177 (N_177,In_539,In_529);
and U178 (N_178,In_476,In_572);
xor U179 (N_179,In_113,In_81);
and U180 (N_180,In_842,In_550);
nor U181 (N_181,In_7,In_170);
or U182 (N_182,In_969,In_941);
and U183 (N_183,In_754,In_971);
nand U184 (N_184,In_946,In_615);
nor U185 (N_185,In_143,In_979);
nor U186 (N_186,In_94,In_604);
nor U187 (N_187,In_183,In_23);
or U188 (N_188,In_994,In_991);
nor U189 (N_189,In_44,In_259);
and U190 (N_190,In_97,In_315);
xnor U191 (N_191,In_997,In_190);
and U192 (N_192,In_317,In_871);
and U193 (N_193,In_640,In_139);
nor U194 (N_194,In_739,In_340);
nand U195 (N_195,In_844,In_481);
xor U196 (N_196,In_59,In_547);
nor U197 (N_197,In_598,In_447);
xor U198 (N_198,In_193,In_610);
or U199 (N_199,In_724,In_109);
or U200 (N_200,In_326,In_487);
xor U201 (N_201,In_291,In_543);
and U202 (N_202,In_974,In_128);
or U203 (N_203,In_675,In_577);
or U204 (N_204,In_993,In_397);
and U205 (N_205,In_45,In_376);
or U206 (N_206,In_964,In_211);
nand U207 (N_207,In_161,In_954);
or U208 (N_208,In_210,In_567);
and U209 (N_209,In_452,In_117);
or U210 (N_210,In_975,In_180);
xnor U211 (N_211,In_194,In_35);
nand U212 (N_212,In_215,In_73);
nor U213 (N_213,In_474,In_495);
or U214 (N_214,In_157,In_937);
and U215 (N_215,In_198,In_528);
nor U216 (N_216,In_595,In_630);
nor U217 (N_217,In_101,In_939);
xor U218 (N_218,In_625,In_189);
nand U219 (N_219,In_104,In_240);
or U220 (N_220,In_562,In_963);
xor U221 (N_221,In_203,In_185);
nor U222 (N_222,In_929,In_672);
nand U223 (N_223,In_679,In_839);
and U224 (N_224,In_992,In_782);
xor U225 (N_225,In_394,In_836);
nor U226 (N_226,In_13,In_78);
nand U227 (N_227,In_324,In_863);
and U228 (N_228,In_243,In_797);
nand U229 (N_229,In_388,In_165);
xor U230 (N_230,In_49,In_972);
and U231 (N_231,In_327,In_852);
and U232 (N_232,In_769,In_247);
xnor U233 (N_233,In_424,In_643);
or U234 (N_234,In_378,In_846);
nor U235 (N_235,In_296,In_961);
or U236 (N_236,In_690,In_632);
nand U237 (N_237,In_199,In_361);
or U238 (N_238,In_620,In_54);
nor U239 (N_239,In_893,In_880);
or U240 (N_240,In_347,In_749);
nand U241 (N_241,In_793,In_407);
and U242 (N_242,In_251,In_569);
xor U243 (N_243,In_4,In_633);
and U244 (N_244,In_670,In_760);
nor U245 (N_245,In_955,In_537);
nor U246 (N_246,In_827,In_52);
xnor U247 (N_247,In_110,In_538);
or U248 (N_248,In_850,In_322);
and U249 (N_249,In_523,In_779);
nand U250 (N_250,In_87,In_396);
nand U251 (N_251,In_646,In_669);
or U252 (N_252,In_290,In_50);
nor U253 (N_253,In_905,In_548);
or U254 (N_254,In_53,In_892);
nand U255 (N_255,In_908,In_775);
or U256 (N_256,In_762,In_766);
or U257 (N_257,In_363,In_80);
nor U258 (N_258,In_262,In_590);
nand U259 (N_259,In_857,In_141);
and U260 (N_260,In_898,In_711);
xnor U261 (N_261,In_244,In_352);
nand U262 (N_262,In_925,In_914);
xnor U263 (N_263,In_996,In_658);
or U264 (N_264,In_807,In_405);
or U265 (N_265,In_42,In_756);
and U266 (N_266,In_511,In_687);
nand U267 (N_267,In_748,In_422);
and U268 (N_268,In_549,In_745);
nand U269 (N_269,In_103,In_524);
and U270 (N_270,In_876,In_292);
xor U271 (N_271,In_587,In_781);
or U272 (N_272,In_153,In_666);
nor U273 (N_273,In_520,In_413);
or U274 (N_274,In_804,In_267);
and U275 (N_275,In_541,In_195);
nand U276 (N_276,In_34,In_408);
xor U277 (N_277,In_28,In_694);
nor U278 (N_278,In_916,In_212);
and U279 (N_279,In_486,In_226);
nand U280 (N_280,In_401,In_594);
nor U281 (N_281,In_612,In_106);
nand U282 (N_282,In_490,In_708);
xnor U283 (N_283,In_989,In_64);
and U284 (N_284,In_881,In_591);
nor U285 (N_285,In_382,In_384);
nor U286 (N_286,In_755,In_692);
nand U287 (N_287,In_400,In_121);
xor U288 (N_288,In_325,In_681);
nand U289 (N_289,In_418,In_228);
and U290 (N_290,In_320,In_798);
or U291 (N_291,In_491,In_889);
nor U292 (N_292,In_242,In_799);
or U293 (N_293,In_894,In_805);
and U294 (N_294,In_576,In_533);
and U295 (N_295,In_127,In_10);
nand U296 (N_296,In_178,In_907);
or U297 (N_297,In_9,In_821);
nand U298 (N_298,In_500,In_900);
or U299 (N_299,In_132,In_693);
nor U300 (N_300,In_603,In_864);
and U301 (N_301,In_174,In_415);
nor U302 (N_302,In_219,In_197);
and U303 (N_303,In_831,In_71);
nor U304 (N_304,In_419,In_970);
nor U305 (N_305,In_653,In_412);
nand U306 (N_306,In_636,In_555);
nor U307 (N_307,In_574,In_980);
nand U308 (N_308,In_772,In_932);
or U309 (N_309,In_140,In_107);
or U310 (N_310,In_79,In_471);
and U311 (N_311,In_114,In_281);
or U312 (N_312,In_246,In_744);
and U313 (N_313,In_426,In_323);
and U314 (N_314,In_227,In_62);
xor U315 (N_315,In_465,In_661);
xor U316 (N_316,In_82,In_743);
nand U317 (N_317,In_381,In_501);
nor U318 (N_318,In_391,In_722);
and U319 (N_319,In_464,In_404);
nor U320 (N_320,In_983,In_904);
or U321 (N_321,In_588,In_346);
and U322 (N_322,In_417,In_512);
and U323 (N_323,In_809,In_250);
and U324 (N_324,In_654,In_841);
xnor U325 (N_325,In_258,In_302);
and U326 (N_326,In_707,In_72);
nand U327 (N_327,In_860,In_245);
and U328 (N_328,In_902,In_531);
nor U329 (N_329,In_206,In_434);
or U330 (N_330,In_774,In_696);
xor U331 (N_331,In_706,In_641);
and U332 (N_332,In_16,In_423);
or U333 (N_333,In_239,In_734);
xor U334 (N_334,In_688,In_85);
nand U335 (N_335,In_530,In_39);
or U336 (N_336,In_126,In_832);
and U337 (N_337,In_626,In_535);
nor U338 (N_338,In_166,In_285);
nor U339 (N_339,In_697,In_297);
or U340 (N_340,In_146,In_321);
or U341 (N_341,In_236,In_990);
nand U342 (N_342,In_507,In_686);
and U343 (N_343,In_984,In_820);
nand U344 (N_344,In_788,In_542);
and U345 (N_345,In_815,In_624);
nand U346 (N_346,In_834,In_678);
nand U347 (N_347,In_398,In_310);
or U348 (N_348,In_379,In_145);
nand U349 (N_349,In_726,In_235);
xnor U350 (N_350,In_727,In_682);
nand U351 (N_351,In_155,In_504);
nand U352 (N_352,In_514,In_985);
xnor U353 (N_353,In_764,In_777);
and U354 (N_354,In_525,In_787);
xor U355 (N_355,In_484,In_448);
nor U356 (N_356,In_299,In_650);
nand U357 (N_357,In_922,In_497);
and U358 (N_358,In_536,In_329);
xor U359 (N_359,In_771,In_436);
nand U360 (N_360,In_502,In_428);
nor U361 (N_361,In_482,In_522);
or U362 (N_362,In_15,In_188);
xor U363 (N_363,In_468,In_184);
nand U364 (N_364,In_492,In_105);
xor U365 (N_365,In_309,In_634);
or U366 (N_366,In_220,In_494);
and U367 (N_367,In_21,In_667);
nand U368 (N_368,In_350,In_386);
xnor U369 (N_369,In_65,In_36);
nand U370 (N_370,In_456,In_14);
nor U371 (N_371,In_923,In_783);
nand U372 (N_372,In_896,In_942);
nand U373 (N_373,In_614,In_817);
nand U374 (N_374,In_207,In_600);
nor U375 (N_375,In_713,In_792);
and U376 (N_376,In_814,In_720);
or U377 (N_377,In_649,In_338);
nand U378 (N_378,In_780,In_192);
and U379 (N_379,In_928,In_319);
nor U380 (N_380,In_784,In_446);
nor U381 (N_381,In_945,In_826);
nand U382 (N_382,In_29,In_458);
or U383 (N_383,In_339,In_367);
or U384 (N_384,In_890,In_702);
and U385 (N_385,In_373,In_58);
nor U386 (N_386,In_162,In_119);
or U387 (N_387,In_420,In_613);
nand U388 (N_388,In_673,In_253);
or U389 (N_389,In_366,In_83);
xor U390 (N_390,In_934,In_102);
xnor U391 (N_391,In_573,In_279);
nand U392 (N_392,In_489,In_786);
xor U393 (N_393,In_99,In_111);
and U394 (N_394,In_998,In_343);
nand U395 (N_395,In_112,In_222);
nor U396 (N_396,In_585,In_116);
nand U397 (N_397,In_698,In_973);
or U398 (N_398,In_662,In_833);
nor U399 (N_399,In_741,In_765);
xnor U400 (N_400,In_510,In_704);
and U401 (N_401,In_919,In_257);
or U402 (N_402,In_534,In_387);
or U403 (N_403,In_621,In_719);
nor U404 (N_404,In_163,In_314);
and U405 (N_405,In_899,In_618);
and U406 (N_406,In_31,In_586);
nor U407 (N_407,In_712,In_728);
nor U408 (N_408,In_622,In_965);
and U409 (N_409,In_671,In_828);
and U410 (N_410,In_770,In_638);
and U411 (N_411,In_861,In_360);
nor U412 (N_412,In_27,In_506);
and U413 (N_413,In_453,In_794);
and U414 (N_414,In_559,In_544);
xnor U415 (N_415,In_740,In_41);
and U416 (N_416,In_186,In_611);
nor U417 (N_417,In_61,In_936);
or U418 (N_418,In_812,In_124);
xnor U419 (N_419,In_467,In_480);
and U420 (N_420,In_837,In_677);
xor U421 (N_421,In_288,In_659);
xnor U422 (N_422,In_17,In_282);
nand U423 (N_423,In_470,In_516);
and U424 (N_424,In_3,In_123);
and U425 (N_425,In_305,In_589);
or U426 (N_426,In_545,In_475);
nor U427 (N_427,In_596,In_303);
xnor U428 (N_428,In_466,In_801);
xnor U429 (N_429,In_808,In_294);
or U430 (N_430,In_280,In_978);
or U431 (N_431,In_680,In_652);
nor U432 (N_432,In_816,In_957);
and U433 (N_433,In_944,In_450);
nor U434 (N_434,In_55,In_571);
xnor U435 (N_435,In_349,In_451);
and U436 (N_436,In_938,In_647);
nand U437 (N_437,In_488,In_849);
xnor U438 (N_438,In_701,In_532);
nor U439 (N_439,In_355,In_848);
or U440 (N_440,In_565,In_703);
nand U441 (N_441,In_337,In_295);
nand U442 (N_442,In_795,In_664);
and U443 (N_443,In_773,In_558);
nor U444 (N_444,In_800,In_229);
or U445 (N_445,In_175,In_307);
nor U446 (N_446,In_200,In_891);
or U447 (N_447,In_133,In_371);
nand U448 (N_448,In_43,In_947);
xor U449 (N_449,In_356,In_411);
or U450 (N_450,In_742,In_223);
and U451 (N_451,In_372,In_389);
nand U452 (N_452,In_374,In_930);
xor U453 (N_453,In_767,In_802);
nand U454 (N_454,In_463,In_135);
and U455 (N_455,In_518,In_933);
or U456 (N_456,In_284,In_521);
xor U457 (N_457,In_906,In_609);
nand U458 (N_458,In_12,In_5);
xnor U459 (N_459,In_263,In_289);
nand U460 (N_460,In_623,In_593);
nor U461 (N_461,In_778,In_181);
or U462 (N_462,In_138,In_856);
nor U463 (N_463,In_221,In_714);
nand U464 (N_464,In_160,In_287);
or U465 (N_465,In_148,In_645);
nand U466 (N_466,In_459,In_269);
nor U467 (N_467,In_750,In_20);
and U468 (N_468,In_977,In_811);
or U469 (N_469,In_362,In_553);
or U470 (N_470,In_790,In_298);
and U471 (N_471,In_663,In_968);
nor U472 (N_472,In_580,In_840);
and U473 (N_473,In_642,In_164);
xor U474 (N_474,In_122,In_248);
xor U475 (N_475,In_88,In_169);
and U476 (N_476,In_19,In_92);
xnor U477 (N_477,In_917,In_264);
and U478 (N_478,In_69,In_496);
nand U479 (N_479,In_563,In_129);
nand U480 (N_480,In_599,In_868);
xnor U481 (N_481,In_879,In_154);
and U482 (N_482,In_556,In_439);
xor U483 (N_483,In_438,In_182);
nand U484 (N_484,In_283,In_218);
or U485 (N_485,In_819,In_485);
xor U486 (N_486,In_723,In_432);
nor U487 (N_487,In_318,In_402);
xnor U488 (N_488,In_472,In_903);
and U489 (N_489,In_716,In_354);
nand U490 (N_490,In_877,In_854);
and U491 (N_491,In_173,In_96);
or U492 (N_492,In_427,In_806);
or U493 (N_493,In_392,In_746);
xor U494 (N_494,In_142,In_469);
or U495 (N_495,In_602,In_342);
nand U496 (N_496,In_375,In_306);
and U497 (N_497,In_66,In_721);
and U498 (N_498,In_144,In_344);
nor U499 (N_499,In_824,In_201);
or U500 (N_500,In_782,In_339);
nor U501 (N_501,In_203,In_744);
nor U502 (N_502,In_875,In_189);
and U503 (N_503,In_154,In_96);
xnor U504 (N_504,In_836,In_237);
or U505 (N_505,In_24,In_3);
nor U506 (N_506,In_977,In_704);
and U507 (N_507,In_235,In_89);
or U508 (N_508,In_587,In_856);
xnor U509 (N_509,In_540,In_876);
nor U510 (N_510,In_657,In_417);
or U511 (N_511,In_504,In_515);
xor U512 (N_512,In_550,In_233);
nand U513 (N_513,In_529,In_292);
and U514 (N_514,In_358,In_769);
xnor U515 (N_515,In_909,In_417);
nor U516 (N_516,In_587,In_85);
and U517 (N_517,In_932,In_330);
nor U518 (N_518,In_110,In_962);
nor U519 (N_519,In_947,In_933);
nor U520 (N_520,In_45,In_43);
nor U521 (N_521,In_859,In_597);
and U522 (N_522,In_20,In_756);
xnor U523 (N_523,In_286,In_473);
nand U524 (N_524,In_743,In_145);
nand U525 (N_525,In_926,In_155);
nand U526 (N_526,In_907,In_341);
and U527 (N_527,In_849,In_601);
nand U528 (N_528,In_770,In_727);
or U529 (N_529,In_752,In_339);
xnor U530 (N_530,In_113,In_233);
xor U531 (N_531,In_98,In_541);
and U532 (N_532,In_756,In_108);
nand U533 (N_533,In_59,In_919);
xnor U534 (N_534,In_69,In_626);
xor U535 (N_535,In_453,In_44);
or U536 (N_536,In_1,In_56);
and U537 (N_537,In_177,In_226);
nand U538 (N_538,In_154,In_92);
nand U539 (N_539,In_870,In_937);
xor U540 (N_540,In_195,In_631);
and U541 (N_541,In_263,In_562);
nand U542 (N_542,In_27,In_863);
or U543 (N_543,In_143,In_698);
or U544 (N_544,In_770,In_135);
and U545 (N_545,In_530,In_801);
or U546 (N_546,In_944,In_128);
and U547 (N_547,In_302,In_329);
nor U548 (N_548,In_520,In_636);
nand U549 (N_549,In_77,In_550);
or U550 (N_550,In_961,In_468);
and U551 (N_551,In_858,In_221);
and U552 (N_552,In_308,In_231);
or U553 (N_553,In_862,In_453);
xor U554 (N_554,In_614,In_611);
xnor U555 (N_555,In_194,In_379);
nand U556 (N_556,In_514,In_833);
xnor U557 (N_557,In_68,In_176);
xnor U558 (N_558,In_109,In_983);
nor U559 (N_559,In_725,In_378);
nand U560 (N_560,In_520,In_358);
nand U561 (N_561,In_258,In_947);
and U562 (N_562,In_538,In_586);
nor U563 (N_563,In_198,In_925);
nor U564 (N_564,In_916,In_287);
or U565 (N_565,In_350,In_601);
xor U566 (N_566,In_305,In_241);
nor U567 (N_567,In_90,In_101);
nand U568 (N_568,In_328,In_804);
and U569 (N_569,In_19,In_146);
and U570 (N_570,In_726,In_443);
and U571 (N_571,In_466,In_944);
nand U572 (N_572,In_43,In_237);
and U573 (N_573,In_474,In_414);
xor U574 (N_574,In_113,In_784);
and U575 (N_575,In_903,In_690);
xnor U576 (N_576,In_945,In_277);
nor U577 (N_577,In_386,In_978);
nor U578 (N_578,In_324,In_658);
and U579 (N_579,In_499,In_442);
and U580 (N_580,In_193,In_465);
xnor U581 (N_581,In_462,In_602);
nor U582 (N_582,In_689,In_189);
and U583 (N_583,In_593,In_654);
nor U584 (N_584,In_429,In_715);
and U585 (N_585,In_275,In_172);
xnor U586 (N_586,In_566,In_245);
nor U587 (N_587,In_180,In_282);
and U588 (N_588,In_60,In_93);
or U589 (N_589,In_17,In_552);
and U590 (N_590,In_162,In_153);
and U591 (N_591,In_618,In_110);
and U592 (N_592,In_548,In_998);
nor U593 (N_593,In_372,In_367);
or U594 (N_594,In_115,In_16);
or U595 (N_595,In_524,In_215);
or U596 (N_596,In_311,In_923);
xnor U597 (N_597,In_61,In_270);
and U598 (N_598,In_746,In_241);
xor U599 (N_599,In_209,In_920);
nor U600 (N_600,In_278,In_619);
xnor U601 (N_601,In_398,In_685);
xnor U602 (N_602,In_769,In_185);
nor U603 (N_603,In_473,In_530);
and U604 (N_604,In_517,In_17);
and U605 (N_605,In_248,In_814);
and U606 (N_606,In_344,In_235);
xor U607 (N_607,In_401,In_752);
nand U608 (N_608,In_294,In_163);
or U609 (N_609,In_3,In_280);
nor U610 (N_610,In_254,In_174);
or U611 (N_611,In_921,In_538);
nand U612 (N_612,In_331,In_657);
or U613 (N_613,In_743,In_971);
xnor U614 (N_614,In_72,In_102);
nor U615 (N_615,In_669,In_105);
nor U616 (N_616,In_708,In_323);
or U617 (N_617,In_3,In_946);
nand U618 (N_618,In_695,In_578);
and U619 (N_619,In_453,In_6);
xnor U620 (N_620,In_34,In_51);
or U621 (N_621,In_13,In_902);
nor U622 (N_622,In_198,In_822);
or U623 (N_623,In_299,In_467);
and U624 (N_624,In_387,In_201);
nor U625 (N_625,In_8,In_271);
nor U626 (N_626,In_767,In_317);
nand U627 (N_627,In_861,In_88);
or U628 (N_628,In_166,In_293);
xnor U629 (N_629,In_872,In_384);
or U630 (N_630,In_788,In_151);
or U631 (N_631,In_6,In_497);
and U632 (N_632,In_147,In_543);
xnor U633 (N_633,In_747,In_262);
and U634 (N_634,In_787,In_412);
nor U635 (N_635,In_221,In_688);
or U636 (N_636,In_142,In_236);
xnor U637 (N_637,In_554,In_667);
xor U638 (N_638,In_548,In_666);
nor U639 (N_639,In_725,In_89);
nor U640 (N_640,In_69,In_958);
xor U641 (N_641,In_997,In_217);
nand U642 (N_642,In_368,In_763);
and U643 (N_643,In_571,In_712);
and U644 (N_644,In_97,In_848);
xnor U645 (N_645,In_354,In_932);
nor U646 (N_646,In_68,In_154);
or U647 (N_647,In_286,In_906);
or U648 (N_648,In_509,In_754);
nand U649 (N_649,In_180,In_657);
and U650 (N_650,In_47,In_882);
and U651 (N_651,In_998,In_556);
xor U652 (N_652,In_494,In_639);
nor U653 (N_653,In_192,In_648);
nor U654 (N_654,In_584,In_752);
nor U655 (N_655,In_444,In_273);
or U656 (N_656,In_162,In_824);
and U657 (N_657,In_536,In_481);
or U658 (N_658,In_400,In_53);
nand U659 (N_659,In_321,In_680);
xor U660 (N_660,In_533,In_177);
or U661 (N_661,In_586,In_579);
nand U662 (N_662,In_246,In_106);
nand U663 (N_663,In_155,In_102);
nand U664 (N_664,In_636,In_830);
nand U665 (N_665,In_933,In_671);
xor U666 (N_666,In_770,In_826);
xnor U667 (N_667,In_929,In_363);
nor U668 (N_668,In_311,In_724);
or U669 (N_669,In_920,In_134);
and U670 (N_670,In_860,In_719);
nand U671 (N_671,In_820,In_724);
or U672 (N_672,In_507,In_58);
xor U673 (N_673,In_471,In_81);
or U674 (N_674,In_160,In_983);
nor U675 (N_675,In_6,In_635);
nor U676 (N_676,In_374,In_466);
nor U677 (N_677,In_541,In_941);
xnor U678 (N_678,In_689,In_71);
and U679 (N_679,In_613,In_301);
and U680 (N_680,In_128,In_264);
and U681 (N_681,In_909,In_638);
nor U682 (N_682,In_319,In_363);
nand U683 (N_683,In_731,In_294);
nand U684 (N_684,In_267,In_500);
xor U685 (N_685,In_761,In_82);
or U686 (N_686,In_822,In_181);
or U687 (N_687,In_755,In_433);
or U688 (N_688,In_447,In_471);
or U689 (N_689,In_821,In_370);
and U690 (N_690,In_232,In_831);
nor U691 (N_691,In_850,In_668);
xor U692 (N_692,In_527,In_760);
and U693 (N_693,In_144,In_544);
nor U694 (N_694,In_5,In_648);
xor U695 (N_695,In_104,In_225);
or U696 (N_696,In_661,In_383);
nand U697 (N_697,In_708,In_79);
nand U698 (N_698,In_282,In_890);
or U699 (N_699,In_812,In_952);
xnor U700 (N_700,In_958,In_100);
xor U701 (N_701,In_107,In_455);
or U702 (N_702,In_882,In_141);
or U703 (N_703,In_462,In_596);
nand U704 (N_704,In_993,In_948);
or U705 (N_705,In_707,In_558);
or U706 (N_706,In_94,In_400);
and U707 (N_707,In_451,In_201);
xor U708 (N_708,In_884,In_506);
and U709 (N_709,In_197,In_584);
xor U710 (N_710,In_482,In_122);
xor U711 (N_711,In_866,In_863);
or U712 (N_712,In_706,In_738);
and U713 (N_713,In_663,In_664);
nor U714 (N_714,In_182,In_918);
nand U715 (N_715,In_546,In_13);
or U716 (N_716,In_646,In_298);
or U717 (N_717,In_523,In_729);
and U718 (N_718,In_377,In_230);
nor U719 (N_719,In_18,In_27);
nor U720 (N_720,In_559,In_334);
nor U721 (N_721,In_447,In_48);
xor U722 (N_722,In_10,In_930);
xor U723 (N_723,In_742,In_77);
and U724 (N_724,In_922,In_869);
or U725 (N_725,In_50,In_571);
and U726 (N_726,In_350,In_639);
nand U727 (N_727,In_443,In_202);
and U728 (N_728,In_426,In_191);
or U729 (N_729,In_502,In_521);
or U730 (N_730,In_227,In_335);
nand U731 (N_731,In_770,In_118);
xor U732 (N_732,In_950,In_174);
and U733 (N_733,In_261,In_532);
nand U734 (N_734,In_908,In_398);
xnor U735 (N_735,In_316,In_391);
and U736 (N_736,In_831,In_750);
and U737 (N_737,In_284,In_351);
or U738 (N_738,In_210,In_393);
or U739 (N_739,In_117,In_597);
xnor U740 (N_740,In_191,In_585);
and U741 (N_741,In_155,In_418);
nand U742 (N_742,In_889,In_966);
nand U743 (N_743,In_109,In_648);
xnor U744 (N_744,In_647,In_966);
nand U745 (N_745,In_461,In_673);
and U746 (N_746,In_614,In_167);
and U747 (N_747,In_960,In_913);
xnor U748 (N_748,In_941,In_642);
nor U749 (N_749,In_525,In_883);
xnor U750 (N_750,In_188,In_218);
nor U751 (N_751,In_75,In_555);
nor U752 (N_752,In_663,In_244);
or U753 (N_753,In_88,In_401);
xor U754 (N_754,In_167,In_181);
or U755 (N_755,In_623,In_672);
or U756 (N_756,In_279,In_339);
or U757 (N_757,In_93,In_390);
nand U758 (N_758,In_340,In_299);
nand U759 (N_759,In_605,In_211);
nand U760 (N_760,In_532,In_452);
nand U761 (N_761,In_181,In_750);
or U762 (N_762,In_824,In_827);
nor U763 (N_763,In_749,In_809);
or U764 (N_764,In_232,In_372);
nor U765 (N_765,In_21,In_622);
or U766 (N_766,In_863,In_943);
xnor U767 (N_767,In_481,In_112);
and U768 (N_768,In_854,In_710);
and U769 (N_769,In_687,In_664);
nor U770 (N_770,In_489,In_826);
nand U771 (N_771,In_722,In_585);
nand U772 (N_772,In_468,In_535);
and U773 (N_773,In_264,In_785);
or U774 (N_774,In_612,In_131);
and U775 (N_775,In_598,In_117);
xor U776 (N_776,In_288,In_596);
nand U777 (N_777,In_53,In_105);
xor U778 (N_778,In_730,In_99);
or U779 (N_779,In_394,In_260);
nor U780 (N_780,In_404,In_674);
and U781 (N_781,In_359,In_917);
or U782 (N_782,In_576,In_854);
and U783 (N_783,In_697,In_751);
and U784 (N_784,In_663,In_396);
nand U785 (N_785,In_56,In_417);
and U786 (N_786,In_736,In_620);
or U787 (N_787,In_482,In_19);
and U788 (N_788,In_638,In_488);
and U789 (N_789,In_51,In_31);
nand U790 (N_790,In_914,In_398);
and U791 (N_791,In_870,In_313);
nand U792 (N_792,In_860,In_637);
nand U793 (N_793,In_665,In_169);
nand U794 (N_794,In_228,In_411);
or U795 (N_795,In_319,In_961);
or U796 (N_796,In_281,In_338);
nor U797 (N_797,In_729,In_430);
nor U798 (N_798,In_20,In_733);
nand U799 (N_799,In_625,In_686);
xor U800 (N_800,In_250,In_495);
nor U801 (N_801,In_836,In_947);
nand U802 (N_802,In_351,In_515);
or U803 (N_803,In_878,In_434);
nor U804 (N_804,In_904,In_845);
and U805 (N_805,In_992,In_422);
or U806 (N_806,In_535,In_528);
nor U807 (N_807,In_7,In_806);
or U808 (N_808,In_282,In_914);
nand U809 (N_809,In_625,In_390);
xnor U810 (N_810,In_397,In_119);
or U811 (N_811,In_402,In_392);
xnor U812 (N_812,In_124,In_267);
or U813 (N_813,In_890,In_646);
nand U814 (N_814,In_568,In_194);
nor U815 (N_815,In_39,In_610);
nor U816 (N_816,In_949,In_841);
and U817 (N_817,In_817,In_712);
nand U818 (N_818,In_808,In_524);
xnor U819 (N_819,In_832,In_174);
xor U820 (N_820,In_366,In_938);
nand U821 (N_821,In_712,In_181);
nand U822 (N_822,In_743,In_540);
nand U823 (N_823,In_57,In_483);
and U824 (N_824,In_947,In_643);
nand U825 (N_825,In_106,In_177);
and U826 (N_826,In_782,In_563);
and U827 (N_827,In_368,In_306);
nor U828 (N_828,In_383,In_790);
nand U829 (N_829,In_491,In_877);
nand U830 (N_830,In_469,In_400);
nor U831 (N_831,In_957,In_130);
nand U832 (N_832,In_515,In_363);
or U833 (N_833,In_556,In_57);
nor U834 (N_834,In_53,In_636);
nand U835 (N_835,In_535,In_713);
xnor U836 (N_836,In_932,In_865);
xnor U837 (N_837,In_92,In_673);
or U838 (N_838,In_794,In_113);
and U839 (N_839,In_492,In_181);
or U840 (N_840,In_749,In_824);
xor U841 (N_841,In_399,In_968);
nand U842 (N_842,In_959,In_127);
nand U843 (N_843,In_361,In_82);
nor U844 (N_844,In_905,In_288);
xnor U845 (N_845,In_9,In_410);
and U846 (N_846,In_995,In_653);
nand U847 (N_847,In_353,In_475);
and U848 (N_848,In_757,In_276);
nand U849 (N_849,In_469,In_966);
or U850 (N_850,In_105,In_578);
or U851 (N_851,In_848,In_916);
and U852 (N_852,In_965,In_317);
or U853 (N_853,In_476,In_243);
nand U854 (N_854,In_101,In_359);
and U855 (N_855,In_728,In_753);
nand U856 (N_856,In_21,In_543);
nor U857 (N_857,In_539,In_873);
nand U858 (N_858,In_691,In_581);
nor U859 (N_859,In_520,In_392);
and U860 (N_860,In_549,In_566);
xor U861 (N_861,In_266,In_636);
nor U862 (N_862,In_716,In_626);
xor U863 (N_863,In_349,In_778);
xor U864 (N_864,In_782,In_22);
nand U865 (N_865,In_186,In_147);
and U866 (N_866,In_204,In_271);
nor U867 (N_867,In_852,In_0);
nor U868 (N_868,In_245,In_849);
nand U869 (N_869,In_484,In_194);
or U870 (N_870,In_313,In_143);
xor U871 (N_871,In_149,In_997);
or U872 (N_872,In_619,In_480);
and U873 (N_873,In_492,In_607);
and U874 (N_874,In_350,In_867);
nand U875 (N_875,In_648,In_895);
or U876 (N_876,In_13,In_396);
xnor U877 (N_877,In_517,In_855);
and U878 (N_878,In_763,In_325);
and U879 (N_879,In_938,In_513);
or U880 (N_880,In_227,In_340);
xnor U881 (N_881,In_956,In_277);
nor U882 (N_882,In_609,In_442);
or U883 (N_883,In_560,In_30);
and U884 (N_884,In_541,In_726);
and U885 (N_885,In_256,In_494);
xor U886 (N_886,In_491,In_904);
nor U887 (N_887,In_504,In_740);
nor U888 (N_888,In_986,In_403);
nor U889 (N_889,In_261,In_143);
or U890 (N_890,In_118,In_462);
nand U891 (N_891,In_119,In_845);
or U892 (N_892,In_329,In_624);
nand U893 (N_893,In_135,In_374);
xnor U894 (N_894,In_472,In_85);
xnor U895 (N_895,In_913,In_577);
nor U896 (N_896,In_948,In_794);
nor U897 (N_897,In_515,In_620);
nand U898 (N_898,In_666,In_908);
xor U899 (N_899,In_416,In_371);
xor U900 (N_900,In_489,In_991);
or U901 (N_901,In_120,In_902);
xor U902 (N_902,In_69,In_307);
nand U903 (N_903,In_173,In_786);
and U904 (N_904,In_242,In_535);
nor U905 (N_905,In_397,In_854);
and U906 (N_906,In_125,In_879);
nor U907 (N_907,In_161,In_690);
xnor U908 (N_908,In_985,In_320);
and U909 (N_909,In_363,In_181);
or U910 (N_910,In_110,In_123);
and U911 (N_911,In_6,In_53);
nor U912 (N_912,In_603,In_317);
nand U913 (N_913,In_102,In_942);
nor U914 (N_914,In_505,In_176);
or U915 (N_915,In_284,In_426);
nand U916 (N_916,In_781,In_754);
and U917 (N_917,In_776,In_946);
nor U918 (N_918,In_454,In_81);
and U919 (N_919,In_899,In_185);
nor U920 (N_920,In_353,In_792);
nand U921 (N_921,In_897,In_841);
xor U922 (N_922,In_597,In_151);
and U923 (N_923,In_317,In_453);
xor U924 (N_924,In_546,In_2);
xor U925 (N_925,In_894,In_717);
xnor U926 (N_926,In_673,In_803);
and U927 (N_927,In_383,In_296);
nand U928 (N_928,In_319,In_873);
xnor U929 (N_929,In_125,In_306);
xnor U930 (N_930,In_17,In_384);
or U931 (N_931,In_133,In_144);
nor U932 (N_932,In_380,In_38);
or U933 (N_933,In_126,In_834);
nor U934 (N_934,In_7,In_82);
and U935 (N_935,In_598,In_682);
and U936 (N_936,In_776,In_572);
xor U937 (N_937,In_26,In_745);
and U938 (N_938,In_239,In_286);
nor U939 (N_939,In_101,In_914);
xnor U940 (N_940,In_720,In_218);
xnor U941 (N_941,In_340,In_999);
nand U942 (N_942,In_20,In_528);
nand U943 (N_943,In_252,In_77);
nor U944 (N_944,In_22,In_941);
nor U945 (N_945,In_280,In_470);
nor U946 (N_946,In_289,In_988);
nor U947 (N_947,In_237,In_491);
or U948 (N_948,In_497,In_945);
and U949 (N_949,In_732,In_744);
and U950 (N_950,In_780,In_36);
or U951 (N_951,In_790,In_920);
or U952 (N_952,In_261,In_49);
and U953 (N_953,In_92,In_762);
and U954 (N_954,In_169,In_573);
xor U955 (N_955,In_429,In_21);
nor U956 (N_956,In_702,In_872);
or U957 (N_957,In_147,In_355);
nand U958 (N_958,In_157,In_651);
nor U959 (N_959,In_759,In_69);
xnor U960 (N_960,In_179,In_532);
xnor U961 (N_961,In_360,In_159);
nand U962 (N_962,In_891,In_397);
and U963 (N_963,In_764,In_994);
or U964 (N_964,In_338,In_847);
or U965 (N_965,In_439,In_25);
or U966 (N_966,In_487,In_781);
and U967 (N_967,In_15,In_260);
xnor U968 (N_968,In_847,In_725);
xnor U969 (N_969,In_537,In_787);
and U970 (N_970,In_539,In_573);
nand U971 (N_971,In_709,In_185);
and U972 (N_972,In_452,In_502);
nand U973 (N_973,In_610,In_651);
nor U974 (N_974,In_196,In_619);
nand U975 (N_975,In_227,In_883);
xnor U976 (N_976,In_753,In_471);
or U977 (N_977,In_470,In_622);
xnor U978 (N_978,In_581,In_932);
nor U979 (N_979,In_178,In_561);
nor U980 (N_980,In_704,In_782);
nand U981 (N_981,In_139,In_167);
nand U982 (N_982,In_584,In_282);
nand U983 (N_983,In_308,In_759);
nand U984 (N_984,In_357,In_483);
or U985 (N_985,In_154,In_438);
nand U986 (N_986,In_294,In_812);
xnor U987 (N_987,In_543,In_228);
and U988 (N_988,In_52,In_833);
or U989 (N_989,In_119,In_567);
or U990 (N_990,In_704,In_988);
xnor U991 (N_991,In_450,In_885);
nand U992 (N_992,In_408,In_891);
and U993 (N_993,In_551,In_696);
or U994 (N_994,In_271,In_98);
nand U995 (N_995,In_577,In_216);
nor U996 (N_996,In_533,In_521);
nand U997 (N_997,In_583,In_578);
nand U998 (N_998,In_338,In_158);
nor U999 (N_999,In_900,In_503);
or U1000 (N_1000,N_18,N_459);
nand U1001 (N_1001,N_715,N_209);
nor U1002 (N_1002,N_467,N_747);
or U1003 (N_1003,N_354,N_673);
nand U1004 (N_1004,N_306,N_776);
or U1005 (N_1005,N_170,N_668);
nor U1006 (N_1006,N_931,N_328);
xor U1007 (N_1007,N_113,N_215);
nor U1008 (N_1008,N_307,N_23);
nand U1009 (N_1009,N_378,N_800);
xnor U1010 (N_1010,N_846,N_440);
nor U1011 (N_1011,N_45,N_135);
or U1012 (N_1012,N_536,N_691);
and U1013 (N_1013,N_841,N_295);
and U1014 (N_1014,N_184,N_341);
and U1015 (N_1015,N_560,N_945);
nand U1016 (N_1016,N_842,N_855);
nor U1017 (N_1017,N_449,N_525);
nand U1018 (N_1018,N_671,N_214);
xnor U1019 (N_1019,N_227,N_516);
xnor U1020 (N_1020,N_946,N_213);
or U1021 (N_1021,N_285,N_823);
nor U1022 (N_1022,N_469,N_533);
or U1023 (N_1023,N_360,N_137);
and U1024 (N_1024,N_416,N_41);
nor U1025 (N_1025,N_350,N_557);
nor U1026 (N_1026,N_875,N_221);
xor U1027 (N_1027,N_356,N_130);
nand U1028 (N_1028,N_547,N_194);
nand U1029 (N_1029,N_476,N_95);
nand U1030 (N_1030,N_926,N_98);
xnor U1031 (N_1031,N_602,N_633);
and U1032 (N_1032,N_573,N_653);
xor U1033 (N_1033,N_826,N_25);
nand U1034 (N_1034,N_918,N_195);
xnor U1035 (N_1035,N_13,N_774);
xnor U1036 (N_1036,N_984,N_454);
nand U1037 (N_1037,N_146,N_927);
xor U1038 (N_1038,N_101,N_634);
and U1039 (N_1039,N_230,N_494);
and U1040 (N_1040,N_446,N_665);
nand U1041 (N_1041,N_973,N_364);
nand U1042 (N_1042,N_229,N_358);
nor U1043 (N_1043,N_461,N_352);
xor U1044 (N_1044,N_298,N_883);
and U1045 (N_1045,N_380,N_854);
xnor U1046 (N_1046,N_594,N_488);
or U1047 (N_1047,N_274,N_474);
nor U1048 (N_1048,N_243,N_296);
nand U1049 (N_1049,N_844,N_375);
nor U1050 (N_1050,N_152,N_735);
and U1051 (N_1051,N_753,N_637);
nor U1052 (N_1052,N_757,N_165);
nand U1053 (N_1053,N_916,N_491);
nand U1054 (N_1054,N_649,N_752);
or U1055 (N_1055,N_681,N_748);
nor U1056 (N_1056,N_845,N_124);
xnor U1057 (N_1057,N_670,N_732);
or U1058 (N_1058,N_466,N_696);
nor U1059 (N_1059,N_455,N_182);
and U1060 (N_1060,N_365,N_962);
xnor U1061 (N_1061,N_801,N_384);
nand U1062 (N_1062,N_472,N_28);
nor U1063 (N_1063,N_241,N_609);
nor U1064 (N_1064,N_911,N_54);
xor U1065 (N_1065,N_895,N_817);
xor U1066 (N_1066,N_938,N_216);
nor U1067 (N_1067,N_627,N_333);
or U1068 (N_1068,N_312,N_499);
xnor U1069 (N_1069,N_746,N_706);
xor U1070 (N_1070,N_813,N_546);
nand U1071 (N_1071,N_138,N_161);
and U1072 (N_1072,N_782,N_340);
xnor U1073 (N_1073,N_880,N_907);
xnor U1074 (N_1074,N_485,N_104);
or U1075 (N_1075,N_919,N_142);
and U1076 (N_1076,N_878,N_82);
or U1077 (N_1077,N_534,N_69);
nor U1078 (N_1078,N_55,N_798);
and U1079 (N_1079,N_27,N_397);
nand U1080 (N_1080,N_527,N_29);
xor U1081 (N_1081,N_587,N_149);
nand U1082 (N_1082,N_379,N_34);
nand U1083 (N_1083,N_596,N_551);
or U1084 (N_1084,N_92,N_768);
or U1085 (N_1085,N_711,N_954);
xor U1086 (N_1086,N_932,N_568);
xor U1087 (N_1087,N_48,N_212);
nor U1088 (N_1088,N_223,N_452);
and U1089 (N_1089,N_612,N_250);
nand U1090 (N_1090,N_120,N_30);
xnor U1091 (N_1091,N_72,N_167);
and U1092 (N_1092,N_980,N_828);
xor U1093 (N_1093,N_481,N_426);
nand U1094 (N_1094,N_299,N_97);
or U1095 (N_1095,N_924,N_122);
xnor U1096 (N_1096,N_33,N_639);
nand U1097 (N_1097,N_291,N_638);
nor U1098 (N_1098,N_871,N_503);
xor U1099 (N_1099,N_5,N_870);
xor U1100 (N_1100,N_96,N_552);
nand U1101 (N_1101,N_601,N_831);
or U1102 (N_1102,N_153,N_114);
nor U1103 (N_1103,N_884,N_190);
nand U1104 (N_1104,N_667,N_119);
nor U1105 (N_1105,N_477,N_240);
nand U1106 (N_1106,N_502,N_193);
or U1107 (N_1107,N_433,N_815);
xnor U1108 (N_1108,N_17,N_934);
xor U1109 (N_1109,N_460,N_159);
or U1110 (N_1110,N_565,N_765);
nor U1111 (N_1111,N_816,N_857);
nand U1112 (N_1112,N_660,N_260);
and U1113 (N_1113,N_548,N_94);
nand U1114 (N_1114,N_265,N_759);
nand U1115 (N_1115,N_635,N_343);
and U1116 (N_1116,N_963,N_382);
xor U1117 (N_1117,N_156,N_626);
or U1118 (N_1118,N_879,N_275);
nand U1119 (N_1119,N_834,N_991);
nor U1120 (N_1120,N_942,N_383);
nand U1121 (N_1121,N_662,N_658);
and U1122 (N_1122,N_81,N_877);
xor U1123 (N_1123,N_687,N_981);
xnor U1124 (N_1124,N_85,N_659);
or U1125 (N_1125,N_710,N_684);
and U1126 (N_1126,N_389,N_258);
nor U1127 (N_1127,N_720,N_648);
and U1128 (N_1128,N_51,N_832);
xor U1129 (N_1129,N_179,N_729);
nand U1130 (N_1130,N_914,N_654);
and U1131 (N_1131,N_308,N_31);
nand U1132 (N_1132,N_123,N_414);
xnor U1133 (N_1133,N_666,N_3);
or U1134 (N_1134,N_868,N_246);
or U1135 (N_1135,N_528,N_738);
nand U1136 (N_1136,N_22,N_707);
and U1137 (N_1137,N_779,N_725);
nor U1138 (N_1138,N_7,N_971);
xor U1139 (N_1139,N_237,N_809);
nor U1140 (N_1140,N_332,N_131);
nand U1141 (N_1141,N_37,N_901);
nor U1142 (N_1142,N_500,N_399);
xor U1143 (N_1143,N_419,N_731);
nand U1144 (N_1144,N_284,N_73);
and U1145 (N_1145,N_251,N_917);
nand U1146 (N_1146,N_592,N_524);
nand U1147 (N_1147,N_550,N_703);
nand U1148 (N_1148,N_65,N_965);
xor U1149 (N_1149,N_226,N_750);
nand U1150 (N_1150,N_559,N_583);
nand U1151 (N_1151,N_852,N_754);
nor U1152 (N_1152,N_368,N_309);
nor U1153 (N_1153,N_836,N_267);
nand U1154 (N_1154,N_283,N_994);
nand U1155 (N_1155,N_608,N_2);
and U1156 (N_1156,N_257,N_327);
xnor U1157 (N_1157,N_204,N_68);
and U1158 (N_1158,N_38,N_572);
nand U1159 (N_1159,N_238,N_764);
and U1160 (N_1160,N_58,N_522);
and U1161 (N_1161,N_960,N_886);
nor U1162 (N_1162,N_408,N_959);
nor U1163 (N_1163,N_90,N_228);
nand U1164 (N_1164,N_171,N_806);
or U1165 (N_1165,N_392,N_825);
or U1166 (N_1166,N_133,N_367);
nand U1167 (N_1167,N_144,N_713);
and U1168 (N_1168,N_763,N_644);
nand U1169 (N_1169,N_937,N_317);
nor U1170 (N_1170,N_155,N_401);
nor U1171 (N_1171,N_822,N_331);
nor U1172 (N_1172,N_0,N_890);
nand U1173 (N_1173,N_66,N_118);
nand U1174 (N_1174,N_778,N_489);
nor U1175 (N_1175,N_603,N_271);
xnor U1176 (N_1176,N_661,N_742);
nand U1177 (N_1177,N_345,N_780);
nand U1178 (N_1178,N_701,N_176);
nor U1179 (N_1179,N_617,N_514);
xnor U1180 (N_1180,N_263,N_24);
and U1181 (N_1181,N_74,N_744);
or U1182 (N_1182,N_542,N_174);
or U1183 (N_1183,N_342,N_52);
xor U1184 (N_1184,N_821,N_874);
nand U1185 (N_1185,N_132,N_346);
nor U1186 (N_1186,N_196,N_941);
nor U1187 (N_1187,N_539,N_783);
nand U1188 (N_1188,N_741,N_187);
nor U1189 (N_1189,N_108,N_43);
xor U1190 (N_1190,N_876,N_904);
and U1191 (N_1191,N_421,N_109);
nor U1192 (N_1192,N_116,N_44);
and U1193 (N_1193,N_128,N_374);
xor U1194 (N_1194,N_330,N_207);
nand U1195 (N_1195,N_575,N_898);
or U1196 (N_1196,N_554,N_409);
nand U1197 (N_1197,N_432,N_509);
or U1198 (N_1198,N_676,N_682);
or U1199 (N_1199,N_688,N_289);
nand U1200 (N_1200,N_859,N_255);
nor U1201 (N_1201,N_357,N_261);
nor U1202 (N_1202,N_789,N_812);
nor U1203 (N_1203,N_273,N_463);
or U1204 (N_1204,N_584,N_20);
xor U1205 (N_1205,N_224,N_610);
or U1206 (N_1206,N_56,N_395);
or U1207 (N_1207,N_53,N_686);
nor U1208 (N_1208,N_811,N_42);
or U1209 (N_1209,N_353,N_301);
and U1210 (N_1210,N_796,N_837);
or U1211 (N_1211,N_430,N_803);
nor U1212 (N_1212,N_833,N_791);
or U1213 (N_1213,N_264,N_785);
nor U1214 (N_1214,N_39,N_311);
nand U1215 (N_1215,N_998,N_482);
xor U1216 (N_1216,N_140,N_517);
or U1217 (N_1217,N_107,N_413);
nand U1218 (N_1218,N_287,N_699);
xor U1219 (N_1219,N_497,N_359);
xnor U1220 (N_1220,N_906,N_210);
xnor U1221 (N_1221,N_843,N_690);
xor U1222 (N_1222,N_758,N_669);
nand U1223 (N_1223,N_136,N_558);
nand U1224 (N_1224,N_473,N_751);
nand U1225 (N_1225,N_511,N_923);
nand U1226 (N_1226,N_531,N_373);
xor U1227 (N_1227,N_166,N_445);
and U1228 (N_1228,N_642,N_348);
or U1229 (N_1229,N_465,N_75);
nand U1230 (N_1230,N_675,N_254);
and U1231 (N_1231,N_967,N_724);
or U1232 (N_1232,N_288,N_436);
or U1233 (N_1233,N_700,N_145);
nor U1234 (N_1234,N_770,N_712);
nand U1235 (N_1235,N_247,N_978);
nand U1236 (N_1236,N_232,N_564);
nor U1237 (N_1237,N_570,N_974);
or U1238 (N_1238,N_944,N_304);
or U1239 (N_1239,N_698,N_405);
nand U1240 (N_1240,N_615,N_76);
nand U1241 (N_1241,N_347,N_294);
or U1242 (N_1242,N_588,N_125);
or U1243 (N_1243,N_492,N_510);
xnor U1244 (N_1244,N_537,N_89);
xor U1245 (N_1245,N_972,N_351);
nor U1246 (N_1246,N_979,N_282);
and U1247 (N_1247,N_105,N_767);
nand U1248 (N_1248,N_57,N_366);
nand U1249 (N_1249,N_189,N_929);
nand U1250 (N_1250,N_989,N_185);
nor U1251 (N_1251,N_191,N_178);
and U1252 (N_1252,N_329,N_180);
nand U1253 (N_1253,N_6,N_336);
nor U1254 (N_1254,N_958,N_672);
nor U1255 (N_1255,N_928,N_1);
and U1256 (N_1256,N_953,N_936);
or U1257 (N_1257,N_632,N_148);
and U1258 (N_1258,N_679,N_276);
nor U1259 (N_1259,N_620,N_920);
nor U1260 (N_1260,N_303,N_802);
or U1261 (N_1261,N_234,N_168);
or U1262 (N_1262,N_630,N_866);
or U1263 (N_1263,N_976,N_172);
nor U1264 (N_1264,N_211,N_434);
or U1265 (N_1265,N_899,N_4);
xor U1266 (N_1266,N_32,N_808);
xor U1267 (N_1267,N_970,N_231);
nor U1268 (N_1268,N_372,N_520);
xor U1269 (N_1269,N_723,N_49);
and U1270 (N_1270,N_158,N_253);
or U1271 (N_1271,N_427,N_292);
or U1272 (N_1272,N_93,N_850);
or U1273 (N_1273,N_252,N_614);
and U1274 (N_1274,N_412,N_504);
or U1275 (N_1275,N_100,N_36);
nor U1276 (N_1276,N_694,N_956);
and U1277 (N_1277,N_730,N_597);
nand U1278 (N_1278,N_9,N_403);
xnor U1279 (N_1279,N_636,N_456);
or U1280 (N_1280,N_745,N_396);
nand U1281 (N_1281,N_921,N_947);
and U1282 (N_1282,N_983,N_279);
nand U1283 (N_1283,N_717,N_618);
or U1284 (N_1284,N_948,N_591);
nand U1285 (N_1285,N_818,N_987);
or U1286 (N_1286,N_997,N_71);
xnor U1287 (N_1287,N_961,N_259);
and U1288 (N_1288,N_721,N_99);
or U1289 (N_1289,N_201,N_391);
nand U1290 (N_1290,N_15,N_865);
nor U1291 (N_1291,N_471,N_349);
or U1292 (N_1292,N_129,N_35);
and U1293 (N_1293,N_233,N_339);
nor U1294 (N_1294,N_840,N_869);
nand U1295 (N_1295,N_404,N_912);
nor U1296 (N_1296,N_362,N_538);
or U1297 (N_1297,N_62,N_900);
or U1298 (N_1298,N_103,N_266);
xnor U1299 (N_1299,N_950,N_88);
and U1300 (N_1300,N_77,N_208);
nor U1301 (N_1301,N_897,N_569);
nor U1302 (N_1302,N_881,N_578);
or U1303 (N_1303,N_310,N_183);
and U1304 (N_1304,N_598,N_293);
nor U1305 (N_1305,N_111,N_198);
or U1306 (N_1306,N_280,N_290);
or U1307 (N_1307,N_655,N_773);
xnor U1308 (N_1308,N_862,N_784);
or U1309 (N_1309,N_338,N_600);
nand U1310 (N_1310,N_319,N_206);
nand U1311 (N_1311,N_448,N_363);
and U1312 (N_1312,N_498,N_269);
nand U1313 (N_1313,N_361,N_739);
and U1314 (N_1314,N_415,N_164);
or U1315 (N_1315,N_512,N_930);
xnor U1316 (N_1316,N_425,N_475);
nor U1317 (N_1317,N_217,N_992);
or U1318 (N_1318,N_795,N_369);
xor U1319 (N_1319,N_487,N_444);
nor U1320 (N_1320,N_11,N_685);
nor U1321 (N_1321,N_235,N_986);
nor U1322 (N_1322,N_50,N_59);
xnor U1323 (N_1323,N_205,N_576);
nand U1324 (N_1324,N_793,N_134);
xnor U1325 (N_1325,N_996,N_589);
nor U1326 (N_1326,N_755,N_714);
nor U1327 (N_1327,N_222,N_641);
nand U1328 (N_1328,N_830,N_457);
or U1329 (N_1329,N_621,N_579);
nor U1330 (N_1330,N_272,N_86);
nand U1331 (N_1331,N_645,N_388);
nor U1332 (N_1332,N_786,N_797);
nor U1333 (N_1333,N_197,N_535);
or U1334 (N_1334,N_486,N_521);
nand U1335 (N_1335,N_628,N_438);
nor U1336 (N_1336,N_804,N_695);
or U1337 (N_1337,N_824,N_305);
xor U1338 (N_1338,N_952,N_450);
and U1339 (N_1339,N_173,N_218);
xnor U1340 (N_1340,N_67,N_417);
or U1341 (N_1341,N_422,N_657);
and U1342 (N_1342,N_16,N_507);
or U1343 (N_1343,N_483,N_902);
nor U1344 (N_1344,N_320,N_286);
and U1345 (N_1345,N_915,N_873);
xor U1346 (N_1346,N_743,N_740);
or U1347 (N_1347,N_12,N_894);
and U1348 (N_1348,N_127,N_727);
xor U1349 (N_1349,N_544,N_736);
nand U1350 (N_1350,N_545,N_799);
and U1351 (N_1351,N_19,N_313);
nor U1352 (N_1352,N_794,N_163);
and U1353 (N_1353,N_115,N_400);
nand U1354 (N_1354,N_300,N_734);
and U1355 (N_1355,N_964,N_680);
nand U1356 (N_1356,N_14,N_318);
or U1357 (N_1357,N_80,N_518);
or U1358 (N_1358,N_787,N_110);
nor U1359 (N_1359,N_624,N_849);
nand U1360 (N_1360,N_442,N_102);
and U1361 (N_1361,N_443,N_451);
and U1362 (N_1362,N_775,N_177);
or U1363 (N_1363,N_969,N_181);
and U1364 (N_1364,N_112,N_910);
or U1365 (N_1365,N_909,N_429);
nor U1366 (N_1366,N_355,N_761);
or U1367 (N_1367,N_777,N_410);
or U1368 (N_1368,N_646,N_70);
nand U1369 (N_1369,N_683,N_143);
xor U1370 (N_1370,N_623,N_322);
nor U1371 (N_1371,N_887,N_933);
and U1372 (N_1372,N_371,N_860);
and U1373 (N_1373,N_495,N_814);
xnor U1374 (N_1374,N_79,N_91);
or U1375 (N_1375,N_861,N_519);
nand U1376 (N_1376,N_175,N_402);
xnor U1377 (N_1377,N_896,N_297);
xor U1378 (N_1378,N_435,N_792);
xor U1379 (N_1379,N_493,N_447);
nand U1380 (N_1380,N_709,N_913);
nor U1381 (N_1381,N_326,N_728);
xor U1382 (N_1382,N_838,N_556);
nand U1383 (N_1383,N_394,N_737);
and U1384 (N_1384,N_561,N_398);
or U1385 (N_1385,N_480,N_506);
nor U1386 (N_1386,N_84,N_420);
or U1387 (N_1387,N_955,N_788);
or U1388 (N_1388,N_563,N_719);
or U1389 (N_1389,N_277,N_664);
nor U1390 (N_1390,N_387,N_968);
nand U1391 (N_1391,N_526,N_242);
nand U1392 (N_1392,N_428,N_622);
nor U1393 (N_1393,N_882,N_925);
xnor U1394 (N_1394,N_64,N_990);
and U1395 (N_1395,N_249,N_549);
or U1396 (N_1396,N_678,N_885);
nor U1397 (N_1397,N_982,N_771);
nand U1398 (N_1398,N_431,N_858);
nor U1399 (N_1399,N_63,N_839);
and U1400 (N_1400,N_656,N_762);
nor U1401 (N_1401,N_381,N_523);
and U1402 (N_1402,N_939,N_325);
or U1403 (N_1403,N_147,N_315);
xnor U1404 (N_1404,N_150,N_157);
nand U1405 (N_1405,N_490,N_484);
or U1406 (N_1406,N_406,N_513);
nor U1407 (N_1407,N_220,N_697);
and U1408 (N_1408,N_501,N_595);
nor U1409 (N_1409,N_46,N_708);
nand U1410 (N_1410,N_424,N_270);
nand U1411 (N_1411,N_468,N_478);
nand U1412 (N_1412,N_571,N_411);
and U1413 (N_1413,N_423,N_805);
or U1414 (N_1414,N_377,N_508);
nor U1415 (N_1415,N_693,N_203);
and U1416 (N_1416,N_625,N_169);
and U1417 (N_1417,N_581,N_335);
or U1418 (N_1418,N_236,N_10);
or U1419 (N_1419,N_692,N_117);
and U1420 (N_1420,N_772,N_139);
and U1421 (N_1421,N_541,N_949);
nand U1422 (N_1422,N_566,N_585);
and U1423 (N_1423,N_891,N_337);
xor U1424 (N_1424,N_704,N_496);
nor U1425 (N_1425,N_121,N_604);
or U1426 (N_1426,N_47,N_87);
or U1427 (N_1427,N_951,N_810);
nand U1428 (N_1428,N_733,N_458);
nand U1429 (N_1429,N_268,N_126);
and U1430 (N_1430,N_376,N_21);
nor U1431 (N_1431,N_888,N_555);
xor U1432 (N_1432,N_716,N_462);
and U1433 (N_1433,N_470,N_851);
and U1434 (N_1434,N_567,N_848);
and U1435 (N_1435,N_993,N_61);
xor U1436 (N_1436,N_940,N_199);
xor U1437 (N_1437,N_616,N_760);
or U1438 (N_1438,N_530,N_574);
or U1439 (N_1439,N_321,N_248);
nor U1440 (N_1440,N_151,N_390);
nand U1441 (N_1441,N_278,N_202);
or U1442 (N_1442,N_769,N_281);
and U1443 (N_1443,N_652,N_385);
xnor U1444 (N_1444,N_722,N_540);
or U1445 (N_1445,N_999,N_26);
and U1446 (N_1446,N_106,N_726);
xnor U1447 (N_1447,N_580,N_599);
nand U1448 (N_1448,N_829,N_872);
and U1449 (N_1449,N_864,N_543);
nand U1450 (N_1450,N_908,N_631);
nor U1451 (N_1451,N_957,N_985);
and U1452 (N_1452,N_643,N_749);
xor U1453 (N_1453,N_966,N_619);
nand U1454 (N_1454,N_532,N_141);
nand U1455 (N_1455,N_650,N_40);
nor U1456 (N_1456,N_441,N_606);
nand U1457 (N_1457,N_889,N_200);
xor U1458 (N_1458,N_651,N_386);
xnor U1459 (N_1459,N_766,N_590);
nand U1460 (N_1460,N_577,N_819);
nor U1461 (N_1461,N_479,N_605);
and U1462 (N_1462,N_867,N_316);
nor U1463 (N_1463,N_781,N_995);
nand U1464 (N_1464,N_324,N_863);
or U1465 (N_1465,N_718,N_418);
and U1466 (N_1466,N_674,N_160);
nand U1467 (N_1467,N_582,N_83);
nor U1468 (N_1468,N_856,N_437);
nand U1469 (N_1469,N_677,N_323);
or U1470 (N_1470,N_827,N_988);
nor U1471 (N_1471,N_922,N_647);
nand U1472 (N_1472,N_239,N_689);
or U1473 (N_1473,N_186,N_245);
nor U1474 (N_1474,N_407,N_935);
nor U1475 (N_1475,N_593,N_893);
or U1476 (N_1476,N_162,N_820);
nand U1477 (N_1477,N_613,N_663);
nand U1478 (N_1478,N_219,N_453);
nor U1479 (N_1479,N_314,N_256);
nor U1480 (N_1480,N_78,N_756);
xor U1481 (N_1481,N_529,N_225);
nor U1482 (N_1482,N_262,N_607);
nor U1483 (N_1483,N_705,N_439);
and U1484 (N_1484,N_807,N_629);
nor U1485 (N_1485,N_943,N_977);
xnor U1486 (N_1486,N_790,N_853);
or U1487 (N_1487,N_847,N_835);
and U1488 (N_1488,N_302,N_188);
nand U1489 (N_1489,N_515,N_975);
nand U1490 (N_1490,N_244,N_562);
nor U1491 (N_1491,N_903,N_154);
and U1492 (N_1492,N_370,N_344);
and U1493 (N_1493,N_586,N_8);
or U1494 (N_1494,N_505,N_611);
nand U1495 (N_1495,N_892,N_334);
nand U1496 (N_1496,N_702,N_464);
or U1497 (N_1497,N_393,N_640);
and U1498 (N_1498,N_553,N_192);
nor U1499 (N_1499,N_60,N_905);
or U1500 (N_1500,N_989,N_380);
nand U1501 (N_1501,N_683,N_449);
nor U1502 (N_1502,N_576,N_270);
and U1503 (N_1503,N_239,N_39);
nand U1504 (N_1504,N_201,N_950);
nand U1505 (N_1505,N_297,N_344);
nand U1506 (N_1506,N_817,N_341);
and U1507 (N_1507,N_332,N_857);
nand U1508 (N_1508,N_147,N_539);
nor U1509 (N_1509,N_218,N_913);
nand U1510 (N_1510,N_756,N_996);
and U1511 (N_1511,N_259,N_742);
nand U1512 (N_1512,N_354,N_586);
xor U1513 (N_1513,N_715,N_337);
or U1514 (N_1514,N_35,N_16);
xor U1515 (N_1515,N_895,N_959);
nand U1516 (N_1516,N_470,N_60);
xnor U1517 (N_1517,N_250,N_640);
and U1518 (N_1518,N_139,N_941);
xnor U1519 (N_1519,N_561,N_840);
xor U1520 (N_1520,N_169,N_763);
and U1521 (N_1521,N_771,N_916);
nor U1522 (N_1522,N_506,N_378);
or U1523 (N_1523,N_320,N_597);
and U1524 (N_1524,N_527,N_788);
and U1525 (N_1525,N_898,N_233);
or U1526 (N_1526,N_382,N_851);
xor U1527 (N_1527,N_255,N_640);
nor U1528 (N_1528,N_86,N_661);
nand U1529 (N_1529,N_705,N_520);
and U1530 (N_1530,N_882,N_676);
xnor U1531 (N_1531,N_476,N_263);
xnor U1532 (N_1532,N_527,N_325);
nand U1533 (N_1533,N_225,N_17);
nand U1534 (N_1534,N_762,N_214);
nor U1535 (N_1535,N_673,N_209);
nor U1536 (N_1536,N_783,N_764);
xor U1537 (N_1537,N_234,N_762);
or U1538 (N_1538,N_157,N_252);
nand U1539 (N_1539,N_772,N_368);
xnor U1540 (N_1540,N_568,N_647);
and U1541 (N_1541,N_752,N_253);
nor U1542 (N_1542,N_839,N_495);
nand U1543 (N_1543,N_661,N_574);
nor U1544 (N_1544,N_402,N_293);
and U1545 (N_1545,N_963,N_950);
or U1546 (N_1546,N_837,N_318);
or U1547 (N_1547,N_141,N_622);
and U1548 (N_1548,N_843,N_428);
nand U1549 (N_1549,N_181,N_108);
nand U1550 (N_1550,N_312,N_802);
nand U1551 (N_1551,N_753,N_247);
xnor U1552 (N_1552,N_721,N_545);
nor U1553 (N_1553,N_534,N_393);
nand U1554 (N_1554,N_154,N_304);
nand U1555 (N_1555,N_639,N_901);
nand U1556 (N_1556,N_957,N_958);
xnor U1557 (N_1557,N_830,N_237);
nand U1558 (N_1558,N_729,N_991);
and U1559 (N_1559,N_957,N_578);
and U1560 (N_1560,N_887,N_295);
and U1561 (N_1561,N_26,N_512);
xor U1562 (N_1562,N_674,N_650);
nor U1563 (N_1563,N_46,N_359);
or U1564 (N_1564,N_739,N_536);
nand U1565 (N_1565,N_22,N_791);
nor U1566 (N_1566,N_343,N_546);
nand U1567 (N_1567,N_564,N_199);
nor U1568 (N_1568,N_422,N_588);
nand U1569 (N_1569,N_711,N_382);
and U1570 (N_1570,N_444,N_922);
nor U1571 (N_1571,N_439,N_671);
xnor U1572 (N_1572,N_578,N_532);
nand U1573 (N_1573,N_934,N_805);
xnor U1574 (N_1574,N_34,N_294);
and U1575 (N_1575,N_962,N_726);
or U1576 (N_1576,N_220,N_833);
xnor U1577 (N_1577,N_47,N_575);
nand U1578 (N_1578,N_367,N_473);
or U1579 (N_1579,N_973,N_246);
nor U1580 (N_1580,N_702,N_927);
and U1581 (N_1581,N_842,N_579);
or U1582 (N_1582,N_640,N_388);
xor U1583 (N_1583,N_45,N_705);
nor U1584 (N_1584,N_642,N_312);
and U1585 (N_1585,N_895,N_477);
nand U1586 (N_1586,N_340,N_15);
and U1587 (N_1587,N_549,N_612);
nor U1588 (N_1588,N_325,N_697);
or U1589 (N_1589,N_300,N_211);
xnor U1590 (N_1590,N_47,N_431);
and U1591 (N_1591,N_663,N_754);
or U1592 (N_1592,N_78,N_903);
and U1593 (N_1593,N_545,N_708);
nand U1594 (N_1594,N_833,N_41);
nor U1595 (N_1595,N_89,N_966);
xor U1596 (N_1596,N_626,N_107);
nor U1597 (N_1597,N_269,N_929);
and U1598 (N_1598,N_813,N_132);
nor U1599 (N_1599,N_38,N_831);
nand U1600 (N_1600,N_17,N_693);
or U1601 (N_1601,N_19,N_8);
and U1602 (N_1602,N_932,N_278);
nor U1603 (N_1603,N_78,N_149);
or U1604 (N_1604,N_425,N_744);
nand U1605 (N_1605,N_588,N_456);
and U1606 (N_1606,N_538,N_732);
or U1607 (N_1607,N_446,N_703);
nand U1608 (N_1608,N_566,N_413);
nor U1609 (N_1609,N_573,N_626);
xor U1610 (N_1610,N_854,N_955);
nand U1611 (N_1611,N_919,N_768);
xnor U1612 (N_1612,N_625,N_582);
or U1613 (N_1613,N_681,N_343);
and U1614 (N_1614,N_512,N_666);
nor U1615 (N_1615,N_466,N_281);
nor U1616 (N_1616,N_943,N_639);
nand U1617 (N_1617,N_469,N_486);
or U1618 (N_1618,N_681,N_462);
nor U1619 (N_1619,N_847,N_953);
nor U1620 (N_1620,N_922,N_100);
and U1621 (N_1621,N_756,N_295);
or U1622 (N_1622,N_663,N_246);
or U1623 (N_1623,N_556,N_972);
nand U1624 (N_1624,N_818,N_568);
and U1625 (N_1625,N_471,N_210);
nand U1626 (N_1626,N_815,N_252);
and U1627 (N_1627,N_111,N_466);
or U1628 (N_1628,N_107,N_918);
or U1629 (N_1629,N_618,N_261);
xnor U1630 (N_1630,N_185,N_588);
nand U1631 (N_1631,N_352,N_167);
xnor U1632 (N_1632,N_353,N_427);
and U1633 (N_1633,N_468,N_582);
xnor U1634 (N_1634,N_517,N_7);
nor U1635 (N_1635,N_142,N_637);
nor U1636 (N_1636,N_470,N_201);
and U1637 (N_1637,N_633,N_749);
or U1638 (N_1638,N_943,N_627);
nor U1639 (N_1639,N_825,N_653);
or U1640 (N_1640,N_107,N_112);
xor U1641 (N_1641,N_215,N_503);
xor U1642 (N_1642,N_497,N_204);
nand U1643 (N_1643,N_594,N_789);
nand U1644 (N_1644,N_919,N_841);
xnor U1645 (N_1645,N_203,N_97);
and U1646 (N_1646,N_127,N_994);
xor U1647 (N_1647,N_677,N_823);
nand U1648 (N_1648,N_783,N_585);
or U1649 (N_1649,N_307,N_981);
or U1650 (N_1650,N_621,N_952);
xnor U1651 (N_1651,N_638,N_538);
and U1652 (N_1652,N_257,N_160);
xor U1653 (N_1653,N_885,N_584);
xnor U1654 (N_1654,N_289,N_851);
nor U1655 (N_1655,N_896,N_27);
xnor U1656 (N_1656,N_292,N_835);
or U1657 (N_1657,N_658,N_819);
or U1658 (N_1658,N_825,N_57);
or U1659 (N_1659,N_937,N_989);
or U1660 (N_1660,N_487,N_546);
nor U1661 (N_1661,N_524,N_326);
xor U1662 (N_1662,N_961,N_933);
and U1663 (N_1663,N_537,N_758);
or U1664 (N_1664,N_882,N_487);
and U1665 (N_1665,N_267,N_794);
nor U1666 (N_1666,N_573,N_195);
and U1667 (N_1667,N_687,N_891);
xnor U1668 (N_1668,N_347,N_955);
and U1669 (N_1669,N_174,N_479);
nand U1670 (N_1670,N_622,N_46);
and U1671 (N_1671,N_658,N_104);
or U1672 (N_1672,N_388,N_742);
or U1673 (N_1673,N_676,N_805);
and U1674 (N_1674,N_264,N_266);
or U1675 (N_1675,N_294,N_624);
and U1676 (N_1676,N_274,N_829);
xor U1677 (N_1677,N_673,N_685);
nand U1678 (N_1678,N_244,N_12);
nor U1679 (N_1679,N_997,N_447);
nand U1680 (N_1680,N_394,N_103);
and U1681 (N_1681,N_652,N_338);
or U1682 (N_1682,N_92,N_464);
or U1683 (N_1683,N_518,N_0);
xnor U1684 (N_1684,N_14,N_182);
nor U1685 (N_1685,N_918,N_733);
and U1686 (N_1686,N_93,N_241);
or U1687 (N_1687,N_474,N_198);
nor U1688 (N_1688,N_757,N_716);
or U1689 (N_1689,N_687,N_320);
nand U1690 (N_1690,N_688,N_441);
nand U1691 (N_1691,N_365,N_218);
or U1692 (N_1692,N_994,N_799);
or U1693 (N_1693,N_234,N_764);
and U1694 (N_1694,N_650,N_772);
xor U1695 (N_1695,N_781,N_36);
nor U1696 (N_1696,N_167,N_671);
xor U1697 (N_1697,N_660,N_959);
and U1698 (N_1698,N_6,N_524);
xor U1699 (N_1699,N_838,N_334);
and U1700 (N_1700,N_30,N_507);
and U1701 (N_1701,N_885,N_570);
or U1702 (N_1702,N_659,N_351);
nand U1703 (N_1703,N_776,N_419);
and U1704 (N_1704,N_556,N_74);
nor U1705 (N_1705,N_498,N_622);
xnor U1706 (N_1706,N_967,N_271);
or U1707 (N_1707,N_143,N_511);
or U1708 (N_1708,N_229,N_815);
or U1709 (N_1709,N_251,N_522);
nand U1710 (N_1710,N_983,N_446);
xor U1711 (N_1711,N_152,N_61);
and U1712 (N_1712,N_108,N_576);
xnor U1713 (N_1713,N_483,N_751);
xor U1714 (N_1714,N_52,N_293);
and U1715 (N_1715,N_638,N_363);
xnor U1716 (N_1716,N_902,N_648);
nand U1717 (N_1717,N_215,N_311);
or U1718 (N_1718,N_307,N_53);
nand U1719 (N_1719,N_211,N_345);
nor U1720 (N_1720,N_262,N_326);
and U1721 (N_1721,N_635,N_251);
and U1722 (N_1722,N_331,N_585);
or U1723 (N_1723,N_379,N_570);
nand U1724 (N_1724,N_307,N_667);
xnor U1725 (N_1725,N_50,N_351);
or U1726 (N_1726,N_58,N_698);
nor U1727 (N_1727,N_515,N_913);
and U1728 (N_1728,N_448,N_957);
nor U1729 (N_1729,N_615,N_119);
nor U1730 (N_1730,N_817,N_358);
and U1731 (N_1731,N_137,N_286);
and U1732 (N_1732,N_146,N_624);
nand U1733 (N_1733,N_147,N_949);
nor U1734 (N_1734,N_474,N_125);
xnor U1735 (N_1735,N_750,N_468);
nor U1736 (N_1736,N_438,N_390);
or U1737 (N_1737,N_714,N_534);
xnor U1738 (N_1738,N_911,N_836);
nand U1739 (N_1739,N_855,N_229);
nor U1740 (N_1740,N_398,N_364);
or U1741 (N_1741,N_127,N_487);
nand U1742 (N_1742,N_983,N_744);
and U1743 (N_1743,N_227,N_462);
or U1744 (N_1744,N_334,N_826);
xor U1745 (N_1745,N_21,N_818);
nor U1746 (N_1746,N_144,N_59);
or U1747 (N_1747,N_874,N_785);
nor U1748 (N_1748,N_353,N_588);
nand U1749 (N_1749,N_700,N_757);
xor U1750 (N_1750,N_728,N_988);
or U1751 (N_1751,N_417,N_366);
nor U1752 (N_1752,N_279,N_266);
nor U1753 (N_1753,N_703,N_939);
nor U1754 (N_1754,N_727,N_386);
xnor U1755 (N_1755,N_921,N_890);
xnor U1756 (N_1756,N_895,N_605);
or U1757 (N_1757,N_542,N_754);
nand U1758 (N_1758,N_322,N_279);
xor U1759 (N_1759,N_357,N_905);
or U1760 (N_1760,N_468,N_962);
nand U1761 (N_1761,N_844,N_380);
nor U1762 (N_1762,N_971,N_989);
and U1763 (N_1763,N_760,N_393);
nor U1764 (N_1764,N_712,N_13);
or U1765 (N_1765,N_639,N_268);
nor U1766 (N_1766,N_602,N_266);
nor U1767 (N_1767,N_668,N_566);
or U1768 (N_1768,N_145,N_662);
xor U1769 (N_1769,N_669,N_240);
and U1770 (N_1770,N_300,N_316);
nand U1771 (N_1771,N_273,N_596);
nand U1772 (N_1772,N_667,N_292);
nand U1773 (N_1773,N_44,N_619);
or U1774 (N_1774,N_507,N_63);
nand U1775 (N_1775,N_106,N_840);
or U1776 (N_1776,N_959,N_136);
nand U1777 (N_1777,N_646,N_241);
and U1778 (N_1778,N_811,N_3);
nor U1779 (N_1779,N_636,N_761);
nand U1780 (N_1780,N_393,N_710);
or U1781 (N_1781,N_379,N_742);
or U1782 (N_1782,N_322,N_679);
nand U1783 (N_1783,N_211,N_159);
and U1784 (N_1784,N_973,N_561);
and U1785 (N_1785,N_444,N_800);
nor U1786 (N_1786,N_553,N_362);
nor U1787 (N_1787,N_633,N_653);
nor U1788 (N_1788,N_102,N_306);
or U1789 (N_1789,N_992,N_766);
and U1790 (N_1790,N_628,N_155);
nand U1791 (N_1791,N_846,N_875);
nand U1792 (N_1792,N_484,N_630);
nor U1793 (N_1793,N_54,N_391);
or U1794 (N_1794,N_682,N_265);
xor U1795 (N_1795,N_615,N_431);
nand U1796 (N_1796,N_481,N_323);
nand U1797 (N_1797,N_342,N_529);
nor U1798 (N_1798,N_777,N_428);
and U1799 (N_1799,N_723,N_291);
and U1800 (N_1800,N_508,N_651);
and U1801 (N_1801,N_990,N_503);
xnor U1802 (N_1802,N_398,N_257);
nand U1803 (N_1803,N_169,N_245);
nor U1804 (N_1804,N_498,N_441);
and U1805 (N_1805,N_825,N_710);
nand U1806 (N_1806,N_443,N_134);
nor U1807 (N_1807,N_953,N_261);
and U1808 (N_1808,N_639,N_392);
and U1809 (N_1809,N_34,N_362);
and U1810 (N_1810,N_896,N_776);
and U1811 (N_1811,N_996,N_8);
and U1812 (N_1812,N_499,N_694);
or U1813 (N_1813,N_360,N_446);
or U1814 (N_1814,N_753,N_791);
or U1815 (N_1815,N_556,N_858);
nor U1816 (N_1816,N_976,N_278);
or U1817 (N_1817,N_794,N_217);
or U1818 (N_1818,N_286,N_497);
and U1819 (N_1819,N_516,N_512);
nand U1820 (N_1820,N_512,N_317);
nand U1821 (N_1821,N_83,N_231);
nand U1822 (N_1822,N_460,N_898);
nor U1823 (N_1823,N_242,N_442);
nand U1824 (N_1824,N_210,N_542);
nor U1825 (N_1825,N_197,N_792);
nor U1826 (N_1826,N_229,N_965);
nand U1827 (N_1827,N_284,N_187);
and U1828 (N_1828,N_204,N_527);
nand U1829 (N_1829,N_570,N_289);
and U1830 (N_1830,N_624,N_322);
nand U1831 (N_1831,N_7,N_728);
nor U1832 (N_1832,N_294,N_307);
and U1833 (N_1833,N_831,N_991);
nor U1834 (N_1834,N_218,N_657);
xor U1835 (N_1835,N_853,N_812);
nand U1836 (N_1836,N_938,N_43);
nand U1837 (N_1837,N_12,N_337);
xnor U1838 (N_1838,N_652,N_877);
nand U1839 (N_1839,N_391,N_327);
or U1840 (N_1840,N_403,N_545);
or U1841 (N_1841,N_493,N_251);
and U1842 (N_1842,N_540,N_930);
xnor U1843 (N_1843,N_932,N_802);
nor U1844 (N_1844,N_506,N_321);
nand U1845 (N_1845,N_218,N_163);
xor U1846 (N_1846,N_975,N_461);
or U1847 (N_1847,N_180,N_665);
or U1848 (N_1848,N_756,N_480);
nand U1849 (N_1849,N_743,N_936);
nand U1850 (N_1850,N_936,N_754);
nand U1851 (N_1851,N_446,N_522);
or U1852 (N_1852,N_584,N_637);
nor U1853 (N_1853,N_727,N_269);
xnor U1854 (N_1854,N_216,N_797);
xnor U1855 (N_1855,N_647,N_232);
and U1856 (N_1856,N_851,N_575);
nand U1857 (N_1857,N_180,N_458);
xnor U1858 (N_1858,N_936,N_468);
and U1859 (N_1859,N_166,N_883);
and U1860 (N_1860,N_160,N_764);
nand U1861 (N_1861,N_982,N_721);
and U1862 (N_1862,N_779,N_838);
and U1863 (N_1863,N_445,N_731);
xnor U1864 (N_1864,N_537,N_79);
nand U1865 (N_1865,N_343,N_994);
and U1866 (N_1866,N_392,N_314);
and U1867 (N_1867,N_463,N_348);
or U1868 (N_1868,N_271,N_140);
or U1869 (N_1869,N_202,N_920);
nand U1870 (N_1870,N_981,N_946);
nor U1871 (N_1871,N_902,N_625);
nand U1872 (N_1872,N_512,N_409);
xor U1873 (N_1873,N_581,N_729);
nor U1874 (N_1874,N_246,N_526);
nor U1875 (N_1875,N_591,N_818);
and U1876 (N_1876,N_483,N_964);
nor U1877 (N_1877,N_681,N_486);
nand U1878 (N_1878,N_353,N_387);
nand U1879 (N_1879,N_821,N_802);
nor U1880 (N_1880,N_485,N_981);
nor U1881 (N_1881,N_947,N_393);
nor U1882 (N_1882,N_1,N_282);
nand U1883 (N_1883,N_832,N_82);
or U1884 (N_1884,N_437,N_977);
xor U1885 (N_1885,N_146,N_520);
xnor U1886 (N_1886,N_759,N_241);
xnor U1887 (N_1887,N_345,N_527);
nand U1888 (N_1888,N_640,N_173);
nand U1889 (N_1889,N_710,N_700);
nand U1890 (N_1890,N_346,N_586);
or U1891 (N_1891,N_324,N_457);
or U1892 (N_1892,N_210,N_320);
or U1893 (N_1893,N_471,N_84);
nor U1894 (N_1894,N_601,N_435);
and U1895 (N_1895,N_270,N_427);
nand U1896 (N_1896,N_849,N_200);
nand U1897 (N_1897,N_44,N_92);
nand U1898 (N_1898,N_883,N_191);
xor U1899 (N_1899,N_232,N_544);
xnor U1900 (N_1900,N_560,N_990);
nor U1901 (N_1901,N_700,N_51);
or U1902 (N_1902,N_836,N_356);
xnor U1903 (N_1903,N_444,N_74);
and U1904 (N_1904,N_81,N_320);
or U1905 (N_1905,N_547,N_574);
xnor U1906 (N_1906,N_251,N_19);
nor U1907 (N_1907,N_924,N_947);
xor U1908 (N_1908,N_61,N_651);
and U1909 (N_1909,N_942,N_22);
nor U1910 (N_1910,N_773,N_350);
xnor U1911 (N_1911,N_721,N_312);
nand U1912 (N_1912,N_633,N_2);
and U1913 (N_1913,N_897,N_577);
nand U1914 (N_1914,N_329,N_275);
nand U1915 (N_1915,N_934,N_66);
and U1916 (N_1916,N_691,N_404);
or U1917 (N_1917,N_48,N_165);
nand U1918 (N_1918,N_213,N_190);
and U1919 (N_1919,N_678,N_403);
and U1920 (N_1920,N_83,N_432);
xnor U1921 (N_1921,N_289,N_572);
nand U1922 (N_1922,N_703,N_316);
nand U1923 (N_1923,N_80,N_179);
nand U1924 (N_1924,N_670,N_500);
xor U1925 (N_1925,N_736,N_55);
xor U1926 (N_1926,N_550,N_589);
nand U1927 (N_1927,N_769,N_418);
nor U1928 (N_1928,N_936,N_163);
nand U1929 (N_1929,N_279,N_965);
nand U1930 (N_1930,N_510,N_508);
or U1931 (N_1931,N_519,N_678);
and U1932 (N_1932,N_968,N_523);
or U1933 (N_1933,N_697,N_73);
and U1934 (N_1934,N_898,N_556);
nor U1935 (N_1935,N_102,N_484);
xnor U1936 (N_1936,N_381,N_190);
xnor U1937 (N_1937,N_93,N_128);
xor U1938 (N_1938,N_499,N_353);
or U1939 (N_1939,N_67,N_65);
or U1940 (N_1940,N_870,N_743);
nor U1941 (N_1941,N_752,N_469);
nand U1942 (N_1942,N_819,N_8);
xnor U1943 (N_1943,N_775,N_498);
xnor U1944 (N_1944,N_218,N_521);
nor U1945 (N_1945,N_797,N_218);
nor U1946 (N_1946,N_93,N_315);
nor U1947 (N_1947,N_913,N_884);
or U1948 (N_1948,N_728,N_266);
xnor U1949 (N_1949,N_274,N_444);
nor U1950 (N_1950,N_471,N_507);
nand U1951 (N_1951,N_886,N_789);
nor U1952 (N_1952,N_28,N_321);
nor U1953 (N_1953,N_115,N_308);
xor U1954 (N_1954,N_888,N_928);
or U1955 (N_1955,N_36,N_904);
nor U1956 (N_1956,N_270,N_467);
and U1957 (N_1957,N_780,N_703);
nand U1958 (N_1958,N_836,N_776);
nor U1959 (N_1959,N_521,N_500);
nor U1960 (N_1960,N_641,N_228);
or U1961 (N_1961,N_830,N_104);
nand U1962 (N_1962,N_457,N_980);
and U1963 (N_1963,N_557,N_649);
and U1964 (N_1964,N_761,N_184);
xnor U1965 (N_1965,N_956,N_434);
and U1966 (N_1966,N_26,N_647);
nand U1967 (N_1967,N_680,N_269);
and U1968 (N_1968,N_835,N_295);
nor U1969 (N_1969,N_572,N_202);
xor U1970 (N_1970,N_228,N_260);
xnor U1971 (N_1971,N_337,N_7);
and U1972 (N_1972,N_618,N_506);
nor U1973 (N_1973,N_27,N_9);
nand U1974 (N_1974,N_325,N_144);
or U1975 (N_1975,N_424,N_628);
nor U1976 (N_1976,N_369,N_311);
or U1977 (N_1977,N_935,N_876);
xnor U1978 (N_1978,N_595,N_91);
nand U1979 (N_1979,N_653,N_671);
xor U1980 (N_1980,N_196,N_356);
xnor U1981 (N_1981,N_811,N_850);
and U1982 (N_1982,N_834,N_926);
and U1983 (N_1983,N_683,N_924);
or U1984 (N_1984,N_699,N_473);
nand U1985 (N_1985,N_499,N_386);
and U1986 (N_1986,N_350,N_904);
xnor U1987 (N_1987,N_953,N_148);
nor U1988 (N_1988,N_994,N_338);
nand U1989 (N_1989,N_927,N_988);
nor U1990 (N_1990,N_659,N_557);
or U1991 (N_1991,N_454,N_147);
and U1992 (N_1992,N_535,N_104);
nor U1993 (N_1993,N_788,N_929);
nor U1994 (N_1994,N_767,N_230);
and U1995 (N_1995,N_962,N_79);
xnor U1996 (N_1996,N_986,N_55);
nor U1997 (N_1997,N_323,N_115);
or U1998 (N_1998,N_996,N_312);
xor U1999 (N_1999,N_708,N_103);
nand U2000 (N_2000,N_1668,N_1445);
and U2001 (N_2001,N_1629,N_1319);
xnor U2002 (N_2002,N_1791,N_1302);
and U2003 (N_2003,N_1682,N_1832);
and U2004 (N_2004,N_1997,N_1779);
or U2005 (N_2005,N_1856,N_1480);
nor U2006 (N_2006,N_1635,N_1403);
and U2007 (N_2007,N_1102,N_1667);
and U2008 (N_2008,N_1361,N_1293);
nand U2009 (N_2009,N_1487,N_1711);
xor U2010 (N_2010,N_1025,N_1378);
nand U2011 (N_2011,N_1740,N_1388);
or U2012 (N_2012,N_1287,N_1936);
or U2013 (N_2013,N_1077,N_1249);
nand U2014 (N_2014,N_1013,N_1336);
nand U2015 (N_2015,N_1631,N_1713);
xnor U2016 (N_2016,N_1289,N_1072);
and U2017 (N_2017,N_1307,N_1156);
xnor U2018 (N_2018,N_1983,N_1611);
and U2019 (N_2019,N_1773,N_1825);
xor U2020 (N_2020,N_1589,N_1954);
nor U2021 (N_2021,N_1402,N_1516);
or U2022 (N_2022,N_1597,N_1996);
or U2023 (N_2023,N_1532,N_1888);
and U2024 (N_2024,N_1309,N_1027);
nand U2025 (N_2025,N_1831,N_1883);
nor U2026 (N_2026,N_1160,N_1690);
and U2027 (N_2027,N_1397,N_1324);
nor U2028 (N_2028,N_1114,N_1626);
nand U2029 (N_2029,N_1218,N_1437);
nor U2030 (N_2030,N_1584,N_1707);
xnor U2031 (N_2031,N_1971,N_1907);
nand U2032 (N_2032,N_1733,N_1554);
or U2033 (N_2033,N_1123,N_1029);
nor U2034 (N_2034,N_1314,N_1570);
xor U2035 (N_2035,N_1693,N_1987);
xor U2036 (N_2036,N_1448,N_1199);
nand U2037 (N_2037,N_1731,N_1255);
or U2038 (N_2038,N_1219,N_1173);
nand U2039 (N_2039,N_1855,N_1952);
nor U2040 (N_2040,N_1694,N_1428);
xor U2041 (N_2041,N_1655,N_1507);
xor U2042 (N_2042,N_1572,N_1168);
or U2043 (N_2043,N_1300,N_1228);
xor U2044 (N_2044,N_1843,N_1178);
or U2045 (N_2045,N_1435,N_1038);
nor U2046 (N_2046,N_1006,N_1460);
nand U2047 (N_2047,N_1527,N_1505);
and U2048 (N_2048,N_1717,N_1250);
nor U2049 (N_2049,N_1747,N_1816);
or U2050 (N_2050,N_1652,N_1327);
and U2051 (N_2051,N_1898,N_1663);
or U2052 (N_2052,N_1468,N_1285);
nand U2053 (N_2053,N_1605,N_1356);
and U2054 (N_2054,N_1271,N_1819);
and U2055 (N_2055,N_1918,N_1879);
xnor U2056 (N_2056,N_1432,N_1761);
xnor U2057 (N_2057,N_1004,N_1782);
and U2058 (N_2058,N_1703,N_1121);
and U2059 (N_2059,N_1908,N_1175);
xnor U2060 (N_2060,N_1870,N_1363);
and U2061 (N_2061,N_1318,N_1624);
and U2062 (N_2062,N_1824,N_1512);
nor U2063 (N_2063,N_1992,N_1033);
nor U2064 (N_2064,N_1665,N_1381);
or U2065 (N_2065,N_1863,N_1009);
xor U2066 (N_2066,N_1661,N_1743);
xnor U2067 (N_2067,N_1391,N_1912);
and U2068 (N_2068,N_1645,N_1498);
and U2069 (N_2069,N_1315,N_1500);
nand U2070 (N_2070,N_1270,N_1198);
nor U2071 (N_2071,N_1808,N_1470);
or U2072 (N_2072,N_1969,N_1478);
nand U2073 (N_2073,N_1642,N_1990);
nor U2074 (N_2074,N_1764,N_1582);
and U2075 (N_2075,N_1368,N_1777);
and U2076 (N_2076,N_1654,N_1535);
nor U2077 (N_2077,N_1488,N_1347);
and U2078 (N_2078,N_1138,N_1400);
and U2079 (N_2079,N_1281,N_1973);
xnor U2080 (N_2080,N_1963,N_1162);
xor U2081 (N_2081,N_1903,N_1798);
xor U2082 (N_2082,N_1752,N_1679);
xor U2083 (N_2083,N_1510,N_1670);
nand U2084 (N_2084,N_1886,N_1538);
and U2085 (N_2085,N_1464,N_1930);
xnor U2086 (N_2086,N_1950,N_1817);
or U2087 (N_2087,N_1834,N_1949);
or U2088 (N_2088,N_1122,N_1180);
xor U2089 (N_2089,N_1265,N_1967);
and U2090 (N_2090,N_1910,N_1880);
nor U2091 (N_2091,N_1279,N_1386);
nor U2092 (N_2092,N_1951,N_1638);
and U2093 (N_2093,N_1502,N_1343);
nor U2094 (N_2094,N_1239,N_1409);
nor U2095 (N_2095,N_1277,N_1770);
nand U2096 (N_2096,N_1669,N_1687);
and U2097 (N_2097,N_1812,N_1062);
and U2098 (N_2098,N_1442,N_1842);
nand U2099 (N_2099,N_1857,N_1174);
nand U2100 (N_2100,N_1932,N_1862);
nor U2101 (N_2101,N_1795,N_1418);
nand U2102 (N_2102,N_1294,N_1905);
and U2103 (N_2103,N_1634,N_1625);
nand U2104 (N_2104,N_1349,N_1060);
nor U2105 (N_2105,N_1001,N_1758);
and U2106 (N_2106,N_1794,N_1454);
or U2107 (N_2107,N_1672,N_1833);
and U2108 (N_2108,N_1523,N_1530);
xnor U2109 (N_2109,N_1960,N_1790);
xnor U2110 (N_2110,N_1157,N_1221);
nand U2111 (N_2111,N_1933,N_1783);
xnor U2112 (N_2112,N_1734,N_1431);
nand U2113 (N_2113,N_1511,N_1709);
and U2114 (N_2114,N_1247,N_1253);
and U2115 (N_2115,N_1387,N_1389);
and U2116 (N_2116,N_1207,N_1847);
xor U2117 (N_2117,N_1142,N_1835);
or U2118 (N_2118,N_1447,N_1109);
and U2119 (N_2119,N_1374,N_1094);
or U2120 (N_2120,N_1297,N_1002);
nand U2121 (N_2121,N_1463,N_1362);
or U2122 (N_2122,N_1177,N_1684);
xnor U2123 (N_2123,N_1167,N_1022);
nand U2124 (N_2124,N_1272,N_1215);
nand U2125 (N_2125,N_1934,N_1152);
or U2126 (N_2126,N_1877,N_1131);
nand U2127 (N_2127,N_1561,N_1537);
xnor U2128 (N_2128,N_1261,N_1685);
and U2129 (N_2129,N_1268,N_1937);
nor U2130 (N_2130,N_1064,N_1686);
nand U2131 (N_2131,N_1020,N_1067);
nand U2132 (N_2132,N_1430,N_1260);
or U2133 (N_2133,N_1548,N_1774);
nand U2134 (N_2134,N_1895,N_1968);
and U2135 (N_2135,N_1039,N_1728);
nand U2136 (N_2136,N_1736,N_1964);
xor U2137 (N_2137,N_1200,N_1061);
nor U2138 (N_2138,N_1134,N_1274);
and U2139 (N_2139,N_1201,N_1225);
nand U2140 (N_2140,N_1818,N_1748);
nand U2141 (N_2141,N_1112,N_1256);
and U2142 (N_2142,N_1757,N_1034);
nand U2143 (N_2143,N_1521,N_1139);
xnor U2144 (N_2144,N_1037,N_1887);
or U2145 (N_2145,N_1931,N_1137);
and U2146 (N_2146,N_1163,N_1858);
xor U2147 (N_2147,N_1604,N_1030);
nor U2148 (N_2148,N_1110,N_1528);
nor U2149 (N_2149,N_1913,N_1775);
and U2150 (N_2150,N_1339,N_1325);
nor U2151 (N_2151,N_1415,N_1925);
xnor U2152 (N_2152,N_1036,N_1729);
or U2153 (N_2153,N_1814,N_1477);
xnor U2154 (N_2154,N_1889,N_1651);
nor U2155 (N_2155,N_1751,N_1380);
or U2156 (N_2156,N_1105,N_1191);
nor U2157 (N_2157,N_1745,N_1283);
nand U2158 (N_2158,N_1522,N_1595);
nor U2159 (N_2159,N_1312,N_1881);
and U2160 (N_2160,N_1490,N_1941);
nor U2161 (N_2161,N_1706,N_1921);
or U2162 (N_2162,N_1014,N_1737);
and U2163 (N_2163,N_1989,N_1557);
nand U2164 (N_2164,N_1227,N_1154);
xnor U2165 (N_2165,N_1508,N_1620);
or U2166 (N_2166,N_1011,N_1637);
and U2167 (N_2167,N_1536,N_1242);
nor U2168 (N_2168,N_1630,N_1308);
nor U2169 (N_2169,N_1662,N_1475);
or U2170 (N_2170,N_1248,N_1202);
or U2171 (N_2171,N_1097,N_1085);
nor U2172 (N_2172,N_1566,N_1115);
nand U2173 (N_2173,N_1063,N_1732);
xnor U2174 (N_2174,N_1130,N_1443);
nand U2175 (N_2175,N_1902,N_1041);
or U2176 (N_2176,N_1809,N_1188);
nor U2177 (N_2177,N_1906,N_1735);
and U2178 (N_2178,N_1046,N_1999);
and U2179 (N_2179,N_1826,N_1456);
nand U2180 (N_2180,N_1229,N_1723);
and U2181 (N_2181,N_1296,N_1525);
nand U2182 (N_2182,N_1111,N_1364);
nand U2183 (N_2183,N_1412,N_1216);
nand U2184 (N_2184,N_1266,N_1617);
or U2185 (N_2185,N_1223,N_1433);
xor U2186 (N_2186,N_1171,N_1853);
xor U2187 (N_2187,N_1165,N_1189);
nor U2188 (N_2188,N_1609,N_1126);
and U2189 (N_2189,N_1796,N_1799);
nor U2190 (N_2190,N_1771,N_1059);
xnor U2191 (N_2191,N_1222,N_1680);
and U2192 (N_2192,N_1158,N_1984);
nand U2193 (N_2193,N_1328,N_1196);
nor U2194 (N_2194,N_1957,N_1392);
and U2195 (N_2195,N_1859,N_1563);
xor U2196 (N_2196,N_1897,N_1514);
nand U2197 (N_2197,N_1753,N_1915);
or U2198 (N_2198,N_1534,N_1718);
nand U2199 (N_2199,N_1334,N_1243);
and U2200 (N_2200,N_1966,N_1830);
nor U2201 (N_2201,N_1854,N_1803);
and U2202 (N_2202,N_1040,N_1264);
xnor U2203 (N_2203,N_1829,N_1917);
nor U2204 (N_2204,N_1691,N_1104);
or U2205 (N_2205,N_1564,N_1822);
nor U2206 (N_2206,N_1553,N_1015);
nand U2207 (N_2207,N_1320,N_1408);
or U2208 (N_2208,N_1474,N_1452);
or U2209 (N_2209,N_1065,N_1664);
and U2210 (N_2210,N_1341,N_1410);
and U2211 (N_2211,N_1190,N_1150);
xnor U2212 (N_2212,N_1288,N_1533);
and U2213 (N_2213,N_1559,N_1153);
xnor U2214 (N_2214,N_1141,N_1575);
xnor U2215 (N_2215,N_1338,N_1252);
xnor U2216 (N_2216,N_1721,N_1100);
xnor U2217 (N_2217,N_1371,N_1186);
nor U2218 (N_2218,N_1394,N_1953);
or U2219 (N_2219,N_1568,N_1784);
or U2220 (N_2220,N_1421,N_1357);
nand U2221 (N_2221,N_1772,N_1928);
or U2222 (N_2222,N_1420,N_1018);
nor U2223 (N_2223,N_1836,N_1267);
and U2224 (N_2224,N_1519,N_1524);
and U2225 (N_2225,N_1323,N_1206);
or U2226 (N_2226,N_1440,N_1348);
nand U2227 (N_2227,N_1096,N_1689);
xor U2228 (N_2228,N_1742,N_1465);
xor U2229 (N_2229,N_1956,N_1032);
nand U2230 (N_2230,N_1867,N_1485);
xor U2231 (N_2231,N_1974,N_1923);
xor U2232 (N_2232,N_1499,N_1991);
nor U2233 (N_2233,N_1547,N_1016);
and U2234 (N_2234,N_1571,N_1346);
and U2235 (N_2235,N_1769,N_1716);
and U2236 (N_2236,N_1161,N_1768);
xor U2237 (N_2237,N_1292,N_1083);
xnor U2238 (N_2238,N_1501,N_1944);
nand U2239 (N_2239,N_1031,N_1263);
or U2240 (N_2240,N_1284,N_1466);
nand U2241 (N_2241,N_1810,N_1451);
nand U2242 (N_2242,N_1531,N_1476);
and U2243 (N_2243,N_1647,N_1237);
and U2244 (N_2244,N_1393,N_1352);
nand U2245 (N_2245,N_1070,N_1384);
or U2246 (N_2246,N_1377,N_1212);
nand U2247 (N_2247,N_1113,N_1805);
and U2248 (N_2248,N_1179,N_1606);
or U2249 (N_2249,N_1079,N_1169);
and U2250 (N_2250,N_1231,N_1955);
and U2251 (N_2251,N_1813,N_1450);
or U2252 (N_2252,N_1149,N_1708);
nor U2253 (N_2253,N_1539,N_1885);
nand U2254 (N_2254,N_1405,N_1164);
nand U2255 (N_2255,N_1765,N_1839);
nand U2256 (N_2256,N_1700,N_1351);
xnor U2257 (N_2257,N_1108,N_1172);
nand U2258 (N_2258,N_1695,N_1762);
nor U2259 (N_2259,N_1414,N_1444);
xor U2260 (N_2260,N_1714,N_1705);
nand U2261 (N_2261,N_1360,N_1492);
nor U2262 (N_2262,N_1756,N_1099);
nand U2263 (N_2263,N_1978,N_1326);
or U2264 (N_2264,N_1639,N_1439);
xnor U2265 (N_2265,N_1052,N_1995);
nand U2266 (N_2266,N_1598,N_1891);
nand U2267 (N_2267,N_1003,N_1851);
nor U2268 (N_2268,N_1927,N_1116);
xor U2269 (N_2269,N_1241,N_1176);
or U2270 (N_2270,N_1993,N_1593);
xnor U2271 (N_2271,N_1005,N_1495);
xnor U2272 (N_2272,N_1872,N_1194);
and U2273 (N_2273,N_1614,N_1453);
nand U2274 (N_2274,N_1788,N_1815);
or U2275 (N_2275,N_1980,N_1750);
nor U2276 (N_2276,N_1649,N_1419);
nand U2277 (N_2277,N_1446,N_1698);
nor U2278 (N_2278,N_1449,N_1674);
nand U2279 (N_2279,N_1778,N_1303);
and U2280 (N_2280,N_1958,N_1692);
and U2281 (N_2281,N_1940,N_1159);
nand U2282 (N_2282,N_1959,N_1573);
nand U2283 (N_2283,N_1491,N_1659);
and U2284 (N_2284,N_1939,N_1244);
and U2285 (N_2285,N_1359,N_1373);
xnor U2286 (N_2286,N_1946,N_1101);
or U2287 (N_2287,N_1311,N_1090);
nand U2288 (N_2288,N_1776,N_1683);
and U2289 (N_2289,N_1182,N_1722);
xor U2290 (N_2290,N_1413,N_1828);
xor U2291 (N_2291,N_1673,N_1755);
nand U2292 (N_2292,N_1185,N_1358);
xor U2293 (N_2293,N_1396,N_1591);
nor U2294 (N_2294,N_1429,N_1084);
xor U2295 (N_2295,N_1864,N_1633);
nand U2296 (N_2296,N_1044,N_1076);
xor U2297 (N_2297,N_1233,N_1214);
xor U2298 (N_2298,N_1354,N_1838);
or U2299 (N_2299,N_1342,N_1192);
nand U2300 (N_2300,N_1929,N_1763);
or U2301 (N_2301,N_1258,N_1896);
nor U2302 (N_2302,N_1407,N_1088);
nor U2303 (N_2303,N_1181,N_1086);
nand U2304 (N_2304,N_1807,N_1330);
xor U2305 (N_2305,N_1618,N_1074);
nor U2306 (N_2306,N_1565,N_1558);
or U2307 (N_2307,N_1837,N_1401);
or U2308 (N_2308,N_1583,N_1081);
and U2309 (N_2309,N_1560,N_1545);
nand U2310 (N_2310,N_1852,N_1120);
or U2311 (N_2311,N_1053,N_1619);
nor U2312 (N_2312,N_1376,N_1230);
xnor U2313 (N_2313,N_1471,N_1844);
or U2314 (N_2314,N_1599,N_1166);
xor U2315 (N_2315,N_1390,N_1744);
and U2316 (N_2316,N_1427,N_1213);
xnor U2317 (N_2317,N_1489,N_1472);
nand U2318 (N_2318,N_1848,N_1459);
or U2319 (N_2319,N_1576,N_1610);
nand U2320 (N_2320,N_1128,N_1304);
and U2321 (N_2321,N_1622,N_1846);
nand U2322 (N_2322,N_1726,N_1613);
or U2323 (N_2323,N_1900,N_1484);
nand U2324 (N_2324,N_1458,N_1926);
nand U2325 (N_2325,N_1197,N_1187);
xnor U2326 (N_2326,N_1259,N_1493);
and U2327 (N_2327,N_1331,N_1183);
nor U2328 (N_2328,N_1845,N_1602);
xnor U2329 (N_2329,N_1045,N_1529);
and U2330 (N_2330,N_1860,N_1416);
and U2331 (N_2331,N_1151,N_1840);
or U2332 (N_2332,N_1461,N_1656);
nand U2333 (N_2333,N_1977,N_1217);
nor U2334 (N_2334,N_1310,N_1370);
nor U2335 (N_2335,N_1496,N_1556);
xnor U2336 (N_2336,N_1073,N_1914);
nor U2337 (N_2337,N_1462,N_1549);
nor U2338 (N_2338,N_1975,N_1050);
or U2339 (N_2339,N_1793,N_1298);
or U2340 (N_2340,N_1211,N_1608);
xnor U2341 (N_2341,N_1008,N_1697);
and U2342 (N_2342,N_1766,N_1650);
nand U2343 (N_2343,N_1787,N_1892);
and U2344 (N_2344,N_1434,N_1055);
nand U2345 (N_2345,N_1517,N_1455);
and U2346 (N_2346,N_1023,N_1945);
or U2347 (N_2347,N_1585,N_1209);
or U2348 (N_2348,N_1071,N_1581);
or U2349 (N_2349,N_1486,N_1965);
nor U2350 (N_2350,N_1701,N_1098);
nor U2351 (N_2351,N_1136,N_1220);
nor U2352 (N_2352,N_1849,N_1724);
nand U2353 (N_2353,N_1603,N_1007);
or U2354 (N_2354,N_1911,N_1290);
or U2355 (N_2355,N_1155,N_1056);
xnor U2356 (N_2356,N_1286,N_1555);
and U2357 (N_2357,N_1132,N_1238);
and U2358 (N_2358,N_1916,N_1893);
and U2359 (N_2359,N_1801,N_1089);
nor U2360 (N_2360,N_1353,N_1372);
and U2361 (N_2361,N_1636,N_1621);
nor U2362 (N_2362,N_1741,N_1379);
nor U2363 (N_2363,N_1457,N_1542);
nor U2364 (N_2364,N_1026,N_1494);
or U2365 (N_2365,N_1425,N_1671);
nor U2366 (N_2366,N_1866,N_1366);
xnor U2367 (N_2367,N_1441,N_1382);
and U2368 (N_2368,N_1301,N_1666);
nor U2369 (N_2369,N_1273,N_1904);
nor U2370 (N_2370,N_1080,N_1580);
nand U2371 (N_2371,N_1337,N_1208);
or U2372 (N_2372,N_1095,N_1746);
nand U2373 (N_2373,N_1800,N_1375);
xor U2374 (N_2374,N_1106,N_1865);
and U2375 (N_2375,N_1049,N_1596);
or U2376 (N_2376,N_1543,N_1601);
nand U2377 (N_2377,N_1117,N_1497);
or U2378 (N_2378,N_1473,N_1333);
xor U2379 (N_2379,N_1607,N_1291);
and U2380 (N_2380,N_1367,N_1520);
or U2381 (N_2381,N_1979,N_1078);
nor U2382 (N_2382,N_1299,N_1562);
nor U2383 (N_2383,N_1612,N_1399);
and U2384 (N_2384,N_1240,N_1827);
nor U2385 (N_2385,N_1899,N_1234);
xor U2386 (N_2386,N_1436,N_1550);
nand U2387 (N_2387,N_1232,N_1972);
nor U2388 (N_2388,N_1119,N_1587);
nor U2389 (N_2389,N_1526,N_1658);
nor U2390 (N_2390,N_1861,N_1942);
and U2391 (N_2391,N_1600,N_1306);
nor U2392 (N_2392,N_1727,N_1785);
nor U2393 (N_2393,N_1344,N_1760);
or U2394 (N_2394,N_1019,N_1569);
or U2395 (N_2395,N_1345,N_1988);
nand U2396 (N_2396,N_1246,N_1884);
or U2397 (N_2397,N_1657,N_1012);
xnor U2398 (N_2398,N_1780,N_1592);
nand U2399 (N_2399,N_1909,N_1615);
nand U2400 (N_2400,N_1438,N_1623);
xnor U2401 (N_2401,N_1254,N_1365);
or U2402 (N_2402,N_1823,N_1143);
nand U2403 (N_2403,N_1616,N_1935);
nor U2404 (N_2404,N_1068,N_1540);
nor U2405 (N_2405,N_1515,N_1710);
nand U2406 (N_2406,N_1588,N_1125);
xnor U2407 (N_2407,N_1546,N_1043);
nor U2408 (N_2408,N_1350,N_1411);
xor U2409 (N_2409,N_1504,N_1586);
xnor U2410 (N_2410,N_1820,N_1203);
nor U2411 (N_2411,N_1193,N_1943);
xnor U2412 (N_2412,N_1469,N_1675);
nand U2413 (N_2413,N_1578,N_1329);
and U2414 (N_2414,N_1048,N_1961);
nor U2415 (N_2415,N_1875,N_1677);
and U2416 (N_2416,N_1894,N_1640);
nand U2417 (N_2417,N_1574,N_1643);
or U2418 (N_2418,N_1204,N_1146);
nor U2419 (N_2419,N_1406,N_1704);
nor U2420 (N_2420,N_1715,N_1841);
xor U2421 (N_2421,N_1148,N_1226);
xnor U2422 (N_2422,N_1797,N_1579);
and U2423 (N_2423,N_1091,N_1195);
nor U2424 (N_2424,N_1340,N_1275);
nand U2425 (N_2425,N_1424,N_1082);
xnor U2426 (N_2426,N_1135,N_1075);
or U2427 (N_2427,N_1878,N_1802);
or U2428 (N_2428,N_1107,N_1874);
and U2429 (N_2429,N_1369,N_1922);
xnor U2430 (N_2430,N_1994,N_1140);
xnor U2431 (N_2431,N_1850,N_1998);
or U2432 (N_2432,N_1947,N_1873);
and U2433 (N_2433,N_1646,N_1245);
and U2434 (N_2434,N_1092,N_1882);
and U2435 (N_2435,N_1986,N_1696);
xnor U2436 (N_2436,N_1676,N_1981);
xnor U2437 (N_2437,N_1144,N_1725);
or U2438 (N_2438,N_1127,N_1924);
and U2439 (N_2439,N_1251,N_1786);
nand U2440 (N_2440,N_1590,N_1118);
nand U2441 (N_2441,N_1481,N_1047);
or U2442 (N_2442,N_1017,N_1422);
nand U2443 (N_2443,N_1594,N_1398);
xor U2444 (N_2444,N_1901,N_1467);
and U2445 (N_2445,N_1948,N_1811);
nor U2446 (N_2446,N_1236,N_1024);
or U2447 (N_2447,N_1383,N_1257);
or U2448 (N_2448,N_1821,N_1276);
or U2449 (N_2449,N_1000,N_1042);
xor U2450 (N_2450,N_1678,N_1305);
and U2451 (N_2451,N_1321,N_1804);
xor U2452 (N_2452,N_1712,N_1976);
xnor U2453 (N_2453,N_1720,N_1057);
nor U2454 (N_2454,N_1322,N_1789);
nor U2455 (N_2455,N_1021,N_1058);
nand U2456 (N_2456,N_1035,N_1739);
or U2457 (N_2457,N_1577,N_1919);
and U2458 (N_2458,N_1509,N_1133);
nor U2459 (N_2459,N_1170,N_1210);
nand U2460 (N_2460,N_1781,N_1087);
nor U2461 (N_2461,N_1806,N_1316);
xnor U2462 (N_2462,N_1681,N_1871);
nor U2463 (N_2463,N_1567,N_1641);
and U2464 (N_2464,N_1385,N_1552);
nand U2465 (N_2465,N_1876,N_1628);
xor U2466 (N_2466,N_1404,N_1482);
xnor U2467 (N_2467,N_1145,N_1513);
and U2468 (N_2468,N_1962,N_1295);
nand U2469 (N_2469,N_1205,N_1632);
nand U2470 (N_2470,N_1627,N_1970);
nor U2471 (N_2471,N_1235,N_1868);
xnor U2472 (N_2472,N_1051,N_1648);
or U2473 (N_2473,N_1262,N_1028);
and U2474 (N_2474,N_1426,N_1551);
nor U2475 (N_2475,N_1423,N_1503);
nand U2476 (N_2476,N_1395,N_1754);
and U2477 (N_2477,N_1792,N_1280);
or U2478 (N_2478,N_1869,N_1738);
nor U2479 (N_2479,N_1129,N_1544);
xnor U2480 (N_2480,N_1103,N_1749);
nor U2481 (N_2481,N_1920,N_1184);
and U2482 (N_2482,N_1890,N_1644);
and U2483 (N_2483,N_1702,N_1317);
nor U2484 (N_2484,N_1010,N_1653);
and U2485 (N_2485,N_1767,N_1269);
nor U2486 (N_2486,N_1985,N_1054);
nor U2487 (N_2487,N_1224,N_1278);
or U2488 (N_2488,N_1483,N_1335);
xor U2489 (N_2489,N_1506,N_1417);
nor U2490 (N_2490,N_1066,N_1730);
nand U2491 (N_2491,N_1719,N_1313);
nor U2492 (N_2492,N_1355,N_1124);
or U2493 (N_2493,N_1282,N_1541);
nor U2494 (N_2494,N_1982,N_1938);
nor U2495 (N_2495,N_1069,N_1479);
nor U2496 (N_2496,N_1688,N_1759);
nand U2497 (N_2497,N_1093,N_1332);
and U2498 (N_2498,N_1660,N_1147);
and U2499 (N_2499,N_1518,N_1699);
or U2500 (N_2500,N_1751,N_1709);
xnor U2501 (N_2501,N_1686,N_1543);
or U2502 (N_2502,N_1110,N_1366);
xor U2503 (N_2503,N_1866,N_1927);
and U2504 (N_2504,N_1516,N_1092);
xnor U2505 (N_2505,N_1229,N_1537);
or U2506 (N_2506,N_1554,N_1228);
xor U2507 (N_2507,N_1401,N_1189);
and U2508 (N_2508,N_1504,N_1447);
and U2509 (N_2509,N_1526,N_1411);
nand U2510 (N_2510,N_1295,N_1425);
xnor U2511 (N_2511,N_1428,N_1960);
xor U2512 (N_2512,N_1339,N_1774);
and U2513 (N_2513,N_1159,N_1105);
or U2514 (N_2514,N_1665,N_1431);
or U2515 (N_2515,N_1502,N_1711);
xnor U2516 (N_2516,N_1504,N_1784);
nand U2517 (N_2517,N_1329,N_1012);
nand U2518 (N_2518,N_1739,N_1075);
nand U2519 (N_2519,N_1265,N_1268);
and U2520 (N_2520,N_1687,N_1760);
and U2521 (N_2521,N_1776,N_1794);
and U2522 (N_2522,N_1695,N_1561);
nand U2523 (N_2523,N_1242,N_1121);
or U2524 (N_2524,N_1275,N_1791);
nand U2525 (N_2525,N_1060,N_1476);
or U2526 (N_2526,N_1011,N_1496);
xnor U2527 (N_2527,N_1961,N_1485);
xor U2528 (N_2528,N_1741,N_1045);
or U2529 (N_2529,N_1879,N_1600);
xor U2530 (N_2530,N_1899,N_1300);
nand U2531 (N_2531,N_1363,N_1697);
nand U2532 (N_2532,N_1815,N_1029);
or U2533 (N_2533,N_1357,N_1757);
and U2534 (N_2534,N_1164,N_1001);
nor U2535 (N_2535,N_1739,N_1434);
nand U2536 (N_2536,N_1378,N_1257);
or U2537 (N_2537,N_1303,N_1428);
and U2538 (N_2538,N_1717,N_1215);
nand U2539 (N_2539,N_1234,N_1763);
nand U2540 (N_2540,N_1495,N_1192);
or U2541 (N_2541,N_1004,N_1124);
xnor U2542 (N_2542,N_1998,N_1919);
nand U2543 (N_2543,N_1787,N_1354);
xnor U2544 (N_2544,N_1180,N_1204);
xnor U2545 (N_2545,N_1904,N_1928);
and U2546 (N_2546,N_1064,N_1716);
or U2547 (N_2547,N_1380,N_1453);
xor U2548 (N_2548,N_1965,N_1582);
or U2549 (N_2549,N_1546,N_1840);
nor U2550 (N_2550,N_1812,N_1520);
nand U2551 (N_2551,N_1130,N_1031);
nor U2552 (N_2552,N_1484,N_1114);
xor U2553 (N_2553,N_1593,N_1758);
nand U2554 (N_2554,N_1901,N_1092);
or U2555 (N_2555,N_1335,N_1664);
nor U2556 (N_2556,N_1814,N_1839);
and U2557 (N_2557,N_1707,N_1905);
or U2558 (N_2558,N_1661,N_1292);
xnor U2559 (N_2559,N_1433,N_1978);
xor U2560 (N_2560,N_1721,N_1708);
or U2561 (N_2561,N_1721,N_1368);
xor U2562 (N_2562,N_1051,N_1783);
or U2563 (N_2563,N_1653,N_1628);
xor U2564 (N_2564,N_1793,N_1417);
nor U2565 (N_2565,N_1137,N_1257);
or U2566 (N_2566,N_1114,N_1666);
nor U2567 (N_2567,N_1029,N_1914);
nor U2568 (N_2568,N_1524,N_1885);
and U2569 (N_2569,N_1671,N_1616);
xor U2570 (N_2570,N_1876,N_1392);
nand U2571 (N_2571,N_1611,N_1296);
and U2572 (N_2572,N_1453,N_1701);
or U2573 (N_2573,N_1672,N_1633);
xnor U2574 (N_2574,N_1631,N_1659);
xor U2575 (N_2575,N_1498,N_1640);
nand U2576 (N_2576,N_1042,N_1088);
or U2577 (N_2577,N_1031,N_1028);
or U2578 (N_2578,N_1688,N_1484);
nor U2579 (N_2579,N_1682,N_1298);
and U2580 (N_2580,N_1770,N_1773);
or U2581 (N_2581,N_1710,N_1652);
nor U2582 (N_2582,N_1843,N_1319);
nand U2583 (N_2583,N_1025,N_1430);
nor U2584 (N_2584,N_1625,N_1791);
or U2585 (N_2585,N_1502,N_1934);
and U2586 (N_2586,N_1349,N_1950);
xor U2587 (N_2587,N_1637,N_1039);
xor U2588 (N_2588,N_1109,N_1715);
and U2589 (N_2589,N_1652,N_1558);
nand U2590 (N_2590,N_1430,N_1842);
nor U2591 (N_2591,N_1547,N_1758);
xor U2592 (N_2592,N_1857,N_1353);
nor U2593 (N_2593,N_1197,N_1611);
xnor U2594 (N_2594,N_1703,N_1054);
and U2595 (N_2595,N_1681,N_1292);
nand U2596 (N_2596,N_1955,N_1809);
or U2597 (N_2597,N_1597,N_1007);
xnor U2598 (N_2598,N_1906,N_1202);
xor U2599 (N_2599,N_1207,N_1602);
nand U2600 (N_2600,N_1069,N_1273);
xor U2601 (N_2601,N_1628,N_1895);
and U2602 (N_2602,N_1420,N_1925);
or U2603 (N_2603,N_1172,N_1083);
nor U2604 (N_2604,N_1011,N_1143);
xor U2605 (N_2605,N_1347,N_1770);
and U2606 (N_2606,N_1482,N_1499);
nor U2607 (N_2607,N_1559,N_1571);
nor U2608 (N_2608,N_1584,N_1268);
and U2609 (N_2609,N_1208,N_1486);
or U2610 (N_2610,N_1131,N_1734);
nand U2611 (N_2611,N_1464,N_1646);
nor U2612 (N_2612,N_1999,N_1161);
nand U2613 (N_2613,N_1267,N_1095);
and U2614 (N_2614,N_1913,N_1074);
and U2615 (N_2615,N_1345,N_1172);
nor U2616 (N_2616,N_1463,N_1157);
nor U2617 (N_2617,N_1911,N_1545);
xnor U2618 (N_2618,N_1444,N_1656);
xor U2619 (N_2619,N_1438,N_1984);
xor U2620 (N_2620,N_1888,N_1795);
nor U2621 (N_2621,N_1976,N_1476);
nor U2622 (N_2622,N_1043,N_1068);
or U2623 (N_2623,N_1093,N_1459);
nand U2624 (N_2624,N_1621,N_1871);
or U2625 (N_2625,N_1956,N_1280);
nand U2626 (N_2626,N_1154,N_1403);
xnor U2627 (N_2627,N_1511,N_1842);
nor U2628 (N_2628,N_1502,N_1203);
and U2629 (N_2629,N_1019,N_1502);
xor U2630 (N_2630,N_1447,N_1049);
and U2631 (N_2631,N_1916,N_1899);
nand U2632 (N_2632,N_1444,N_1324);
nand U2633 (N_2633,N_1945,N_1991);
nand U2634 (N_2634,N_1180,N_1840);
nor U2635 (N_2635,N_1782,N_1249);
and U2636 (N_2636,N_1397,N_1909);
nand U2637 (N_2637,N_1949,N_1558);
and U2638 (N_2638,N_1435,N_1997);
nor U2639 (N_2639,N_1357,N_1361);
nor U2640 (N_2640,N_1682,N_1941);
nand U2641 (N_2641,N_1954,N_1001);
and U2642 (N_2642,N_1839,N_1850);
nor U2643 (N_2643,N_1091,N_1942);
nor U2644 (N_2644,N_1758,N_1834);
and U2645 (N_2645,N_1314,N_1484);
xor U2646 (N_2646,N_1463,N_1433);
and U2647 (N_2647,N_1493,N_1749);
nor U2648 (N_2648,N_1216,N_1203);
or U2649 (N_2649,N_1720,N_1340);
xor U2650 (N_2650,N_1675,N_1701);
and U2651 (N_2651,N_1405,N_1348);
and U2652 (N_2652,N_1217,N_1181);
and U2653 (N_2653,N_1418,N_1121);
nand U2654 (N_2654,N_1744,N_1672);
nand U2655 (N_2655,N_1618,N_1519);
nand U2656 (N_2656,N_1183,N_1605);
nand U2657 (N_2657,N_1344,N_1380);
and U2658 (N_2658,N_1315,N_1243);
xnor U2659 (N_2659,N_1362,N_1942);
and U2660 (N_2660,N_1988,N_1102);
or U2661 (N_2661,N_1098,N_1459);
nand U2662 (N_2662,N_1522,N_1091);
nand U2663 (N_2663,N_1703,N_1968);
nor U2664 (N_2664,N_1390,N_1691);
nor U2665 (N_2665,N_1614,N_1178);
or U2666 (N_2666,N_1515,N_1819);
or U2667 (N_2667,N_1414,N_1229);
or U2668 (N_2668,N_1006,N_1932);
xor U2669 (N_2669,N_1647,N_1493);
nor U2670 (N_2670,N_1822,N_1584);
xor U2671 (N_2671,N_1122,N_1279);
and U2672 (N_2672,N_1734,N_1414);
or U2673 (N_2673,N_1672,N_1678);
and U2674 (N_2674,N_1227,N_1225);
nand U2675 (N_2675,N_1142,N_1312);
and U2676 (N_2676,N_1583,N_1076);
nor U2677 (N_2677,N_1179,N_1696);
xnor U2678 (N_2678,N_1858,N_1614);
xnor U2679 (N_2679,N_1810,N_1565);
nand U2680 (N_2680,N_1699,N_1511);
or U2681 (N_2681,N_1676,N_1338);
xnor U2682 (N_2682,N_1268,N_1606);
xnor U2683 (N_2683,N_1986,N_1445);
and U2684 (N_2684,N_1298,N_1617);
and U2685 (N_2685,N_1638,N_1953);
nand U2686 (N_2686,N_1612,N_1605);
nor U2687 (N_2687,N_1276,N_1604);
nand U2688 (N_2688,N_1242,N_1972);
or U2689 (N_2689,N_1131,N_1101);
xnor U2690 (N_2690,N_1810,N_1524);
or U2691 (N_2691,N_1984,N_1397);
and U2692 (N_2692,N_1749,N_1136);
nor U2693 (N_2693,N_1474,N_1140);
or U2694 (N_2694,N_1605,N_1483);
xor U2695 (N_2695,N_1986,N_1713);
xor U2696 (N_2696,N_1897,N_1091);
and U2697 (N_2697,N_1279,N_1650);
xor U2698 (N_2698,N_1097,N_1492);
xor U2699 (N_2699,N_1358,N_1299);
or U2700 (N_2700,N_1975,N_1732);
and U2701 (N_2701,N_1473,N_1335);
nand U2702 (N_2702,N_1629,N_1403);
nand U2703 (N_2703,N_1947,N_1367);
nand U2704 (N_2704,N_1116,N_1402);
or U2705 (N_2705,N_1992,N_1904);
nand U2706 (N_2706,N_1035,N_1040);
and U2707 (N_2707,N_1763,N_1237);
or U2708 (N_2708,N_1914,N_1300);
nand U2709 (N_2709,N_1801,N_1063);
nand U2710 (N_2710,N_1357,N_1411);
nand U2711 (N_2711,N_1280,N_1623);
and U2712 (N_2712,N_1460,N_1020);
and U2713 (N_2713,N_1909,N_1087);
nor U2714 (N_2714,N_1884,N_1929);
xnor U2715 (N_2715,N_1883,N_1481);
or U2716 (N_2716,N_1509,N_1069);
and U2717 (N_2717,N_1279,N_1657);
nand U2718 (N_2718,N_1728,N_1730);
xnor U2719 (N_2719,N_1707,N_1137);
or U2720 (N_2720,N_1215,N_1217);
and U2721 (N_2721,N_1233,N_1012);
and U2722 (N_2722,N_1144,N_1066);
or U2723 (N_2723,N_1366,N_1157);
or U2724 (N_2724,N_1179,N_1866);
nand U2725 (N_2725,N_1239,N_1717);
nor U2726 (N_2726,N_1341,N_1925);
xnor U2727 (N_2727,N_1649,N_1644);
nor U2728 (N_2728,N_1006,N_1494);
and U2729 (N_2729,N_1857,N_1412);
and U2730 (N_2730,N_1124,N_1472);
nand U2731 (N_2731,N_1419,N_1964);
nor U2732 (N_2732,N_1047,N_1625);
or U2733 (N_2733,N_1980,N_1473);
or U2734 (N_2734,N_1481,N_1515);
nor U2735 (N_2735,N_1491,N_1660);
and U2736 (N_2736,N_1250,N_1941);
and U2737 (N_2737,N_1260,N_1616);
nand U2738 (N_2738,N_1634,N_1852);
and U2739 (N_2739,N_1730,N_1623);
and U2740 (N_2740,N_1438,N_1463);
xnor U2741 (N_2741,N_1314,N_1410);
xor U2742 (N_2742,N_1377,N_1704);
nor U2743 (N_2743,N_1472,N_1352);
nand U2744 (N_2744,N_1961,N_1670);
nor U2745 (N_2745,N_1632,N_1900);
and U2746 (N_2746,N_1235,N_1445);
nand U2747 (N_2747,N_1890,N_1155);
nor U2748 (N_2748,N_1197,N_1179);
or U2749 (N_2749,N_1591,N_1890);
nor U2750 (N_2750,N_1193,N_1412);
xnor U2751 (N_2751,N_1986,N_1256);
and U2752 (N_2752,N_1211,N_1203);
nand U2753 (N_2753,N_1639,N_1215);
or U2754 (N_2754,N_1138,N_1030);
and U2755 (N_2755,N_1431,N_1346);
xor U2756 (N_2756,N_1458,N_1868);
and U2757 (N_2757,N_1000,N_1963);
and U2758 (N_2758,N_1202,N_1155);
or U2759 (N_2759,N_1094,N_1646);
nand U2760 (N_2760,N_1770,N_1566);
or U2761 (N_2761,N_1134,N_1204);
or U2762 (N_2762,N_1067,N_1347);
and U2763 (N_2763,N_1121,N_1171);
xor U2764 (N_2764,N_1311,N_1841);
nor U2765 (N_2765,N_1778,N_1126);
nor U2766 (N_2766,N_1829,N_1453);
nor U2767 (N_2767,N_1268,N_1017);
or U2768 (N_2768,N_1350,N_1584);
nor U2769 (N_2769,N_1334,N_1862);
xnor U2770 (N_2770,N_1932,N_1603);
and U2771 (N_2771,N_1731,N_1665);
nor U2772 (N_2772,N_1893,N_1139);
or U2773 (N_2773,N_1267,N_1333);
or U2774 (N_2774,N_1675,N_1755);
xor U2775 (N_2775,N_1687,N_1874);
nand U2776 (N_2776,N_1646,N_1115);
or U2777 (N_2777,N_1273,N_1751);
and U2778 (N_2778,N_1175,N_1274);
xnor U2779 (N_2779,N_1531,N_1362);
nand U2780 (N_2780,N_1365,N_1646);
and U2781 (N_2781,N_1751,N_1362);
nor U2782 (N_2782,N_1361,N_1989);
or U2783 (N_2783,N_1857,N_1181);
and U2784 (N_2784,N_1871,N_1271);
and U2785 (N_2785,N_1511,N_1540);
or U2786 (N_2786,N_1051,N_1840);
xnor U2787 (N_2787,N_1084,N_1944);
or U2788 (N_2788,N_1637,N_1684);
nand U2789 (N_2789,N_1182,N_1440);
xnor U2790 (N_2790,N_1062,N_1148);
nand U2791 (N_2791,N_1166,N_1979);
and U2792 (N_2792,N_1137,N_1090);
nor U2793 (N_2793,N_1070,N_1888);
or U2794 (N_2794,N_1284,N_1216);
nor U2795 (N_2795,N_1427,N_1291);
nand U2796 (N_2796,N_1600,N_1293);
nor U2797 (N_2797,N_1727,N_1154);
nor U2798 (N_2798,N_1345,N_1809);
xnor U2799 (N_2799,N_1625,N_1230);
or U2800 (N_2800,N_1370,N_1817);
or U2801 (N_2801,N_1201,N_1256);
or U2802 (N_2802,N_1994,N_1346);
nand U2803 (N_2803,N_1027,N_1204);
and U2804 (N_2804,N_1317,N_1565);
and U2805 (N_2805,N_1778,N_1904);
nand U2806 (N_2806,N_1560,N_1891);
or U2807 (N_2807,N_1373,N_1779);
nor U2808 (N_2808,N_1245,N_1181);
nor U2809 (N_2809,N_1008,N_1225);
xnor U2810 (N_2810,N_1034,N_1778);
xor U2811 (N_2811,N_1128,N_1407);
xnor U2812 (N_2812,N_1885,N_1512);
or U2813 (N_2813,N_1141,N_1989);
xor U2814 (N_2814,N_1947,N_1471);
nand U2815 (N_2815,N_1850,N_1094);
or U2816 (N_2816,N_1875,N_1758);
nand U2817 (N_2817,N_1455,N_1609);
nand U2818 (N_2818,N_1894,N_1938);
nand U2819 (N_2819,N_1890,N_1703);
nor U2820 (N_2820,N_1068,N_1677);
nor U2821 (N_2821,N_1524,N_1750);
and U2822 (N_2822,N_1208,N_1773);
and U2823 (N_2823,N_1568,N_1734);
nor U2824 (N_2824,N_1336,N_1808);
nor U2825 (N_2825,N_1443,N_1775);
nor U2826 (N_2826,N_1955,N_1313);
or U2827 (N_2827,N_1134,N_1921);
xor U2828 (N_2828,N_1945,N_1983);
nor U2829 (N_2829,N_1437,N_1076);
xor U2830 (N_2830,N_1207,N_1292);
and U2831 (N_2831,N_1851,N_1184);
nor U2832 (N_2832,N_1429,N_1274);
nor U2833 (N_2833,N_1319,N_1519);
xor U2834 (N_2834,N_1208,N_1188);
and U2835 (N_2835,N_1018,N_1811);
nand U2836 (N_2836,N_1209,N_1367);
or U2837 (N_2837,N_1465,N_1918);
nor U2838 (N_2838,N_1430,N_1130);
xor U2839 (N_2839,N_1835,N_1821);
and U2840 (N_2840,N_1238,N_1652);
nand U2841 (N_2841,N_1904,N_1345);
nor U2842 (N_2842,N_1942,N_1111);
xnor U2843 (N_2843,N_1267,N_1120);
nand U2844 (N_2844,N_1458,N_1525);
or U2845 (N_2845,N_1708,N_1208);
nor U2846 (N_2846,N_1107,N_1193);
nand U2847 (N_2847,N_1274,N_1578);
nor U2848 (N_2848,N_1671,N_1990);
xnor U2849 (N_2849,N_1291,N_1139);
xor U2850 (N_2850,N_1060,N_1064);
and U2851 (N_2851,N_1409,N_1111);
nand U2852 (N_2852,N_1618,N_1963);
nand U2853 (N_2853,N_1693,N_1794);
or U2854 (N_2854,N_1415,N_1401);
nand U2855 (N_2855,N_1042,N_1954);
nand U2856 (N_2856,N_1618,N_1032);
or U2857 (N_2857,N_1950,N_1641);
or U2858 (N_2858,N_1454,N_1026);
nor U2859 (N_2859,N_1111,N_1740);
xnor U2860 (N_2860,N_1580,N_1796);
nand U2861 (N_2861,N_1838,N_1089);
and U2862 (N_2862,N_1051,N_1883);
nor U2863 (N_2863,N_1740,N_1744);
xor U2864 (N_2864,N_1065,N_1543);
and U2865 (N_2865,N_1669,N_1560);
nor U2866 (N_2866,N_1258,N_1574);
and U2867 (N_2867,N_1591,N_1321);
and U2868 (N_2868,N_1168,N_1838);
nand U2869 (N_2869,N_1138,N_1584);
xor U2870 (N_2870,N_1701,N_1192);
nand U2871 (N_2871,N_1498,N_1610);
nand U2872 (N_2872,N_1188,N_1644);
xor U2873 (N_2873,N_1955,N_1375);
and U2874 (N_2874,N_1082,N_1464);
xor U2875 (N_2875,N_1549,N_1775);
nor U2876 (N_2876,N_1338,N_1248);
nand U2877 (N_2877,N_1821,N_1974);
xor U2878 (N_2878,N_1886,N_1252);
and U2879 (N_2879,N_1622,N_1970);
and U2880 (N_2880,N_1239,N_1632);
or U2881 (N_2881,N_1431,N_1107);
xnor U2882 (N_2882,N_1548,N_1666);
xnor U2883 (N_2883,N_1360,N_1846);
xor U2884 (N_2884,N_1262,N_1396);
and U2885 (N_2885,N_1313,N_1371);
nand U2886 (N_2886,N_1859,N_1628);
nor U2887 (N_2887,N_1785,N_1602);
nand U2888 (N_2888,N_1382,N_1572);
xnor U2889 (N_2889,N_1803,N_1616);
xor U2890 (N_2890,N_1242,N_1736);
nor U2891 (N_2891,N_1820,N_1941);
nand U2892 (N_2892,N_1823,N_1731);
or U2893 (N_2893,N_1114,N_1389);
nand U2894 (N_2894,N_1112,N_1512);
nor U2895 (N_2895,N_1536,N_1046);
and U2896 (N_2896,N_1924,N_1575);
or U2897 (N_2897,N_1417,N_1280);
and U2898 (N_2898,N_1585,N_1122);
or U2899 (N_2899,N_1170,N_1069);
nand U2900 (N_2900,N_1513,N_1029);
and U2901 (N_2901,N_1460,N_1126);
and U2902 (N_2902,N_1740,N_1360);
and U2903 (N_2903,N_1410,N_1639);
nor U2904 (N_2904,N_1753,N_1288);
xnor U2905 (N_2905,N_1479,N_1992);
xor U2906 (N_2906,N_1535,N_1205);
nand U2907 (N_2907,N_1056,N_1017);
or U2908 (N_2908,N_1569,N_1485);
nor U2909 (N_2909,N_1523,N_1914);
nor U2910 (N_2910,N_1324,N_1071);
or U2911 (N_2911,N_1829,N_1158);
nand U2912 (N_2912,N_1975,N_1150);
nand U2913 (N_2913,N_1115,N_1754);
nor U2914 (N_2914,N_1016,N_1247);
or U2915 (N_2915,N_1254,N_1897);
and U2916 (N_2916,N_1530,N_1147);
nand U2917 (N_2917,N_1691,N_1713);
xnor U2918 (N_2918,N_1985,N_1277);
or U2919 (N_2919,N_1063,N_1623);
and U2920 (N_2920,N_1508,N_1520);
nand U2921 (N_2921,N_1162,N_1221);
and U2922 (N_2922,N_1591,N_1235);
or U2923 (N_2923,N_1026,N_1344);
and U2924 (N_2924,N_1435,N_1279);
xor U2925 (N_2925,N_1659,N_1451);
xnor U2926 (N_2926,N_1794,N_1535);
or U2927 (N_2927,N_1463,N_1870);
nand U2928 (N_2928,N_1750,N_1296);
nor U2929 (N_2929,N_1198,N_1849);
or U2930 (N_2930,N_1056,N_1315);
nand U2931 (N_2931,N_1024,N_1260);
xor U2932 (N_2932,N_1994,N_1493);
or U2933 (N_2933,N_1480,N_1269);
nand U2934 (N_2934,N_1035,N_1247);
nand U2935 (N_2935,N_1997,N_1877);
nand U2936 (N_2936,N_1897,N_1618);
nand U2937 (N_2937,N_1340,N_1552);
xnor U2938 (N_2938,N_1464,N_1478);
nand U2939 (N_2939,N_1010,N_1165);
nor U2940 (N_2940,N_1855,N_1381);
xor U2941 (N_2941,N_1291,N_1096);
and U2942 (N_2942,N_1093,N_1110);
or U2943 (N_2943,N_1096,N_1722);
nor U2944 (N_2944,N_1467,N_1376);
nand U2945 (N_2945,N_1400,N_1108);
and U2946 (N_2946,N_1166,N_1516);
and U2947 (N_2947,N_1101,N_1007);
nor U2948 (N_2948,N_1578,N_1076);
nand U2949 (N_2949,N_1694,N_1425);
and U2950 (N_2950,N_1489,N_1557);
nor U2951 (N_2951,N_1025,N_1803);
or U2952 (N_2952,N_1230,N_1155);
nand U2953 (N_2953,N_1794,N_1188);
nand U2954 (N_2954,N_1992,N_1834);
or U2955 (N_2955,N_1435,N_1176);
xnor U2956 (N_2956,N_1232,N_1406);
xnor U2957 (N_2957,N_1646,N_1966);
xor U2958 (N_2958,N_1167,N_1541);
or U2959 (N_2959,N_1104,N_1491);
nand U2960 (N_2960,N_1262,N_1462);
or U2961 (N_2961,N_1061,N_1998);
nand U2962 (N_2962,N_1490,N_1964);
and U2963 (N_2963,N_1160,N_1959);
xor U2964 (N_2964,N_1512,N_1905);
nor U2965 (N_2965,N_1661,N_1442);
or U2966 (N_2966,N_1210,N_1924);
nor U2967 (N_2967,N_1226,N_1473);
xnor U2968 (N_2968,N_1233,N_1004);
and U2969 (N_2969,N_1943,N_1930);
nor U2970 (N_2970,N_1955,N_1556);
or U2971 (N_2971,N_1574,N_1014);
nand U2972 (N_2972,N_1026,N_1552);
nand U2973 (N_2973,N_1358,N_1951);
xnor U2974 (N_2974,N_1531,N_1975);
or U2975 (N_2975,N_1103,N_1563);
nand U2976 (N_2976,N_1362,N_1347);
nand U2977 (N_2977,N_1665,N_1152);
and U2978 (N_2978,N_1066,N_1687);
nand U2979 (N_2979,N_1725,N_1523);
or U2980 (N_2980,N_1939,N_1801);
xnor U2981 (N_2981,N_1041,N_1543);
and U2982 (N_2982,N_1818,N_1269);
or U2983 (N_2983,N_1352,N_1000);
nor U2984 (N_2984,N_1045,N_1130);
or U2985 (N_2985,N_1345,N_1245);
nor U2986 (N_2986,N_1743,N_1875);
nor U2987 (N_2987,N_1626,N_1878);
xnor U2988 (N_2988,N_1878,N_1478);
and U2989 (N_2989,N_1974,N_1208);
and U2990 (N_2990,N_1646,N_1861);
and U2991 (N_2991,N_1384,N_1539);
xnor U2992 (N_2992,N_1355,N_1873);
xor U2993 (N_2993,N_1004,N_1323);
nor U2994 (N_2994,N_1795,N_1122);
or U2995 (N_2995,N_1352,N_1110);
nor U2996 (N_2996,N_1965,N_1309);
xor U2997 (N_2997,N_1881,N_1541);
and U2998 (N_2998,N_1245,N_1504);
nand U2999 (N_2999,N_1340,N_1065);
nor U3000 (N_3000,N_2882,N_2492);
and U3001 (N_3001,N_2351,N_2757);
and U3002 (N_3002,N_2203,N_2145);
or U3003 (N_3003,N_2269,N_2358);
nand U3004 (N_3004,N_2515,N_2721);
and U3005 (N_3005,N_2233,N_2587);
and U3006 (N_3006,N_2905,N_2206);
xor U3007 (N_3007,N_2558,N_2644);
nor U3008 (N_3008,N_2257,N_2796);
xor U3009 (N_3009,N_2525,N_2226);
xnor U3010 (N_3010,N_2969,N_2607);
xnor U3011 (N_3011,N_2639,N_2890);
and U3012 (N_3012,N_2056,N_2496);
nor U3013 (N_3013,N_2316,N_2093);
xor U3014 (N_3014,N_2650,N_2336);
nand U3015 (N_3015,N_2262,N_2741);
and U3016 (N_3016,N_2931,N_2579);
and U3017 (N_3017,N_2772,N_2596);
and U3018 (N_3018,N_2082,N_2478);
and U3019 (N_3019,N_2410,N_2394);
or U3020 (N_3020,N_2957,N_2344);
nand U3021 (N_3021,N_2662,N_2548);
or U3022 (N_3022,N_2378,N_2227);
nor U3023 (N_3023,N_2047,N_2542);
nor U3024 (N_3024,N_2207,N_2057);
or U3025 (N_3025,N_2891,N_2723);
nand U3026 (N_3026,N_2756,N_2384);
and U3027 (N_3027,N_2967,N_2432);
and U3028 (N_3028,N_2580,N_2318);
nor U3029 (N_3029,N_2341,N_2750);
or U3030 (N_3030,N_2357,N_2068);
nand U3031 (N_3031,N_2265,N_2292);
xor U3032 (N_3032,N_2675,N_2812);
nand U3033 (N_3033,N_2865,N_2908);
nand U3034 (N_3034,N_2991,N_2470);
or U3035 (N_3035,N_2561,N_2396);
nand U3036 (N_3036,N_2011,N_2943);
or U3037 (N_3037,N_2832,N_2692);
or U3038 (N_3038,N_2286,N_2742);
nor U3039 (N_3039,N_2764,N_2331);
xor U3040 (N_3040,N_2454,N_2465);
nor U3041 (N_3041,N_2950,N_2877);
xnor U3042 (N_3042,N_2635,N_2502);
and U3043 (N_3043,N_2321,N_2523);
nand U3044 (N_3044,N_2555,N_2802);
and U3045 (N_3045,N_2980,N_2522);
xor U3046 (N_3046,N_2553,N_2346);
or U3047 (N_3047,N_2067,N_2420);
nand U3048 (N_3048,N_2114,N_2044);
xor U3049 (N_3049,N_2095,N_2317);
nor U3050 (N_3050,N_2264,N_2614);
or U3051 (N_3051,N_2792,N_2340);
nor U3052 (N_3052,N_2187,N_2472);
xor U3053 (N_3053,N_2586,N_2433);
nor U3054 (N_3054,N_2505,N_2214);
nor U3055 (N_3055,N_2213,N_2618);
xor U3056 (N_3056,N_2605,N_2874);
and U3057 (N_3057,N_2038,N_2075);
nor U3058 (N_3058,N_2304,N_2391);
and U3059 (N_3059,N_2312,N_2962);
or U3060 (N_3060,N_2245,N_2517);
nor U3061 (N_3061,N_2805,N_2685);
nor U3062 (N_3062,N_2875,N_2576);
and U3063 (N_3063,N_2965,N_2475);
nand U3064 (N_3064,N_2388,N_2694);
and U3065 (N_3065,N_2033,N_2025);
and U3066 (N_3066,N_2268,N_2134);
xor U3067 (N_3067,N_2017,N_2016);
or U3068 (N_3068,N_2857,N_2101);
nand U3069 (N_3069,N_2974,N_2275);
nor U3070 (N_3070,N_2946,N_2296);
xnor U3071 (N_3071,N_2333,N_2456);
nand U3072 (N_3072,N_2636,N_2731);
nand U3073 (N_3073,N_2012,N_2283);
xor U3074 (N_3074,N_2087,N_2199);
or U3075 (N_3075,N_2099,N_2229);
xor U3076 (N_3076,N_2904,N_2418);
xor U3077 (N_3077,N_2823,N_2246);
nor U3078 (N_3078,N_2365,N_2160);
nor U3079 (N_3079,N_2147,N_2876);
xor U3080 (N_3080,N_2574,N_2864);
nor U3081 (N_3081,N_2319,N_2055);
xor U3082 (N_3082,N_2747,N_2966);
nor U3083 (N_3083,N_2354,N_2234);
nor U3084 (N_3084,N_2191,N_2745);
and U3085 (N_3085,N_2666,N_2322);
nand U3086 (N_3086,N_2437,N_2701);
and U3087 (N_3087,N_2853,N_2704);
nor U3088 (N_3088,N_2609,N_2254);
and U3089 (N_3089,N_2440,N_2362);
nand U3090 (N_3090,N_2272,N_2842);
and U3091 (N_3091,N_2601,N_2899);
nor U3092 (N_3092,N_2273,N_2712);
nand U3093 (N_3093,N_2993,N_2421);
nand U3094 (N_3094,N_2951,N_2359);
nand U3095 (N_3095,N_2810,N_2997);
xnor U3096 (N_3096,N_2090,N_2615);
nand U3097 (N_3097,N_2276,N_2734);
nor U3098 (N_3098,N_2063,N_2473);
nor U3099 (N_3099,N_2252,N_2348);
xnor U3100 (N_3100,N_2168,N_2976);
and U3101 (N_3101,N_2474,N_2504);
nor U3102 (N_3102,N_2688,N_2451);
nor U3103 (N_3103,N_2298,N_2516);
nor U3104 (N_3104,N_2042,N_2935);
nand U3105 (N_3105,N_2487,N_2049);
and U3106 (N_3106,N_2181,N_2386);
or U3107 (N_3107,N_2933,N_2520);
nor U3108 (N_3108,N_2881,N_2441);
xor U3109 (N_3109,N_2591,N_2002);
or U3110 (N_3110,N_2198,N_2104);
nand U3111 (N_3111,N_2076,N_2807);
or U3112 (N_3112,N_2290,N_2366);
nand U3113 (N_3113,N_2611,N_2767);
and U3114 (N_3114,N_2783,N_2638);
nand U3115 (N_3115,N_2032,N_2755);
or U3116 (N_3116,N_2870,N_2142);
and U3117 (N_3117,N_2034,N_2699);
and U3118 (N_3118,N_2713,N_2886);
xor U3119 (N_3119,N_2556,N_2782);
nand U3120 (N_3120,N_2045,N_2380);
or U3121 (N_3121,N_2917,N_2236);
nand U3122 (N_3122,N_2197,N_2428);
or U3123 (N_3123,N_2249,N_2968);
or U3124 (N_3124,N_2566,N_2368);
xor U3125 (N_3125,N_2453,N_2854);
xnor U3126 (N_3126,N_2003,N_2387);
or U3127 (N_3127,N_2156,N_2061);
nand U3128 (N_3128,N_2413,N_2686);
and U3129 (N_3129,N_2578,N_2878);
and U3130 (N_3130,N_2824,N_2895);
nor U3131 (N_3131,N_2669,N_2036);
and U3132 (N_3132,N_2445,N_2221);
nand U3133 (N_3133,N_2288,N_2773);
xor U3134 (N_3134,N_2811,N_2959);
xor U3135 (N_3135,N_2927,N_2350);
and U3136 (N_3136,N_2656,N_2128);
nor U3137 (N_3137,N_2179,N_2146);
nand U3138 (N_3138,N_2948,N_2702);
and U3139 (N_3139,N_2389,N_2171);
nand U3140 (N_3140,N_2982,N_2661);
nand U3141 (N_3141,N_2758,N_2111);
and U3142 (N_3142,N_2051,N_2697);
and U3143 (N_3143,N_2008,N_2912);
nand U3144 (N_3144,N_2856,N_2964);
xnor U3145 (N_3145,N_2626,N_2488);
xor U3146 (N_3146,N_2078,N_2131);
and U3147 (N_3147,N_2289,N_2484);
nor U3148 (N_3148,N_2536,N_2715);
nand U3149 (N_3149,N_2630,N_2370);
nand U3150 (N_3150,N_2623,N_2695);
or U3151 (N_3151,N_2754,N_2508);
xnor U3152 (N_3152,N_2102,N_2161);
nand U3153 (N_3153,N_2598,N_2816);
nand U3154 (N_3154,N_2295,N_2762);
nor U3155 (N_3155,N_2294,N_2706);
or U3156 (N_3156,N_2442,N_2654);
and U3157 (N_3157,N_2983,N_2640);
nor U3158 (N_3158,N_2833,N_2521);
xnor U3159 (N_3159,N_2349,N_2200);
and U3160 (N_3160,N_2460,N_2519);
nor U3161 (N_3161,N_2390,N_2960);
nand U3162 (N_3162,N_2846,N_2159);
or U3163 (N_3163,N_2798,N_2788);
nand U3164 (N_3164,N_2172,N_2840);
xor U3165 (N_3165,N_2363,N_2914);
or U3166 (N_3166,N_2039,N_2210);
and U3167 (N_3167,N_2019,N_2732);
nor U3168 (N_3168,N_2543,N_2722);
nor U3169 (N_3169,N_2133,N_2787);
and U3170 (N_3170,N_2324,N_2896);
or U3171 (N_3171,N_2251,N_2244);
nor U3172 (N_3172,N_2961,N_2583);
nor U3173 (N_3173,N_2112,N_2415);
or U3174 (N_3174,N_2613,N_2608);
or U3175 (N_3175,N_2533,N_2748);
or U3176 (N_3176,N_2308,N_2998);
nor U3177 (N_3177,N_2205,N_2281);
nor U3178 (N_3178,N_2863,N_2549);
nand U3179 (N_3179,N_2117,N_2570);
or U3180 (N_3180,N_2115,N_2155);
xnor U3181 (N_3181,N_2060,N_2970);
or U3182 (N_3182,N_2332,N_2157);
nor U3183 (N_3183,N_2148,N_2749);
or U3184 (N_3184,N_2271,N_2633);
nor U3185 (N_3185,N_2446,N_2430);
nand U3186 (N_3186,N_2469,N_2239);
nand U3187 (N_3187,N_2778,N_2136);
nor U3188 (N_3188,N_2184,N_2270);
nor U3189 (N_3189,N_2105,N_2814);
nor U3190 (N_3190,N_2577,N_2594);
nand U3191 (N_3191,N_2023,N_2986);
nand U3192 (N_3192,N_2154,N_2676);
nand U3193 (N_3193,N_2267,N_2110);
nand U3194 (N_3194,N_2809,N_2600);
and U3195 (N_3195,N_2567,N_2373);
and U3196 (N_3196,N_2595,N_2338);
xnor U3197 (N_3197,N_2907,N_2138);
xnor U3198 (N_3198,N_2303,N_2844);
nor U3199 (N_3199,N_2506,N_2158);
and U3200 (N_3200,N_2862,N_2855);
or U3201 (N_3201,N_2660,N_2489);
nor U3202 (N_3202,N_2402,N_2301);
nand U3203 (N_3203,N_2422,N_2909);
nand U3204 (N_3204,N_2530,N_2717);
and U3205 (N_3205,N_2979,N_2637);
nand U3206 (N_3206,N_2822,N_2170);
nor U3207 (N_3207,N_2328,N_2728);
xor U3208 (N_3208,N_2375,N_2920);
and U3209 (N_3209,N_2151,N_2592);
nand U3210 (N_3210,N_2427,N_2932);
xnor U3211 (N_3211,N_2455,N_2797);
nor U3212 (N_3212,N_2382,N_2169);
and U3213 (N_3213,N_2334,N_2551);
nor U3214 (N_3214,N_2795,N_2022);
nor U3215 (N_3215,N_2524,N_2135);
and U3216 (N_3216,N_2975,N_2746);
nand U3217 (N_3217,N_2632,N_2994);
nand U3218 (N_3218,N_2072,N_2679);
nor U3219 (N_3219,N_2938,N_2237);
and U3220 (N_3220,N_2476,N_2009);
or U3221 (N_3221,N_2682,N_2235);
and U3222 (N_3222,N_2837,N_2848);
and U3223 (N_3223,N_2513,N_2144);
and U3224 (N_3224,N_2284,N_2010);
or U3225 (N_3225,N_2766,N_2841);
nor U3226 (N_3226,N_2879,N_2751);
and U3227 (N_3227,N_2510,N_2922);
nor U3228 (N_3228,N_2070,N_2497);
nand U3229 (N_3229,N_2314,N_2217);
nor U3230 (N_3230,N_2062,N_2936);
nor U3231 (N_3231,N_2569,N_2693);
xor U3232 (N_3232,N_2821,N_2597);
and U3233 (N_3233,N_2326,N_2554);
xnor U3234 (N_3234,N_2079,N_2861);
and U3235 (N_3235,N_2282,N_2691);
nand U3236 (N_3236,N_2887,N_2956);
nor U3237 (N_3237,N_2028,N_2190);
or U3238 (N_3238,N_2655,N_2176);
nand U3239 (N_3239,N_2431,N_2188);
xor U3240 (N_3240,N_2696,N_2037);
xor U3241 (N_3241,N_2174,N_2077);
nand U3242 (N_3242,N_2125,N_2836);
and U3243 (N_3243,N_2674,N_2263);
nand U3244 (N_3244,N_2483,N_2083);
nand U3245 (N_3245,N_2494,N_2645);
nand U3246 (N_3246,N_2653,N_2089);
or U3247 (N_3247,N_2371,N_2232);
xnor U3248 (N_3248,N_2582,N_2439);
and U3249 (N_3249,N_2825,N_2098);
xnor U3250 (N_3250,N_2126,N_2537);
xnor U3251 (N_3251,N_2910,N_2624);
nor U3252 (N_3252,N_2647,N_2829);
xnor U3253 (N_3253,N_2612,N_2572);
and U3254 (N_3254,N_2681,N_2992);
or U3255 (N_3255,N_2124,N_2230);
xnor U3256 (N_3256,N_2790,N_2094);
xnor U3257 (N_3257,N_2406,N_2452);
or U3258 (N_3258,N_2311,N_2310);
and U3259 (N_3259,N_2941,N_2954);
xor U3260 (N_3260,N_2779,N_2643);
nor U3261 (N_3261,N_2139,N_2564);
and U3262 (N_3262,N_2759,N_2532);
or U3263 (N_3263,N_2794,N_2163);
or U3264 (N_3264,N_2186,N_2066);
or U3265 (N_3265,N_2573,N_2627);
or U3266 (N_3266,N_2892,N_2355);
nor U3267 (N_3267,N_2784,N_2827);
nand U3268 (N_3268,N_2468,N_2765);
xor U3269 (N_3269,N_2781,N_2541);
nand U3270 (N_3270,N_2498,N_2804);
and U3271 (N_3271,N_2058,N_2086);
nand U3272 (N_3272,N_2356,N_2107);
nor U3273 (N_3273,N_2059,N_2053);
nor U3274 (N_3274,N_2625,N_2700);
and U3275 (N_3275,N_2719,N_2735);
xor U3276 (N_3276,N_2447,N_2990);
or U3277 (N_3277,N_2106,N_2806);
nor U3278 (N_3278,N_2776,N_2538);
or U3279 (N_3279,N_2622,N_2423);
nand U3280 (N_3280,N_2726,N_2031);
nor U3281 (N_3281,N_2345,N_2512);
nor U3282 (N_3282,N_2467,N_2725);
nor U3283 (N_3283,N_2118,N_2429);
xnor U3284 (N_3284,N_2074,N_2302);
nand U3285 (N_3285,N_2547,N_2557);
or U3286 (N_3286,N_2668,N_2479);
or U3287 (N_3287,N_2116,N_2999);
or U3288 (N_3288,N_2004,N_2397);
nand U3289 (N_3289,N_2540,N_2740);
nand U3290 (N_3290,N_2849,N_2934);
nand U3291 (N_3291,N_2379,N_2122);
nand U3292 (N_3292,N_2385,N_2071);
and U3293 (N_3293,N_2871,N_2720);
nand U3294 (N_3294,N_2514,N_2534);
and U3295 (N_3295,N_2733,N_2178);
nand U3296 (N_3296,N_2834,N_2684);
nor U3297 (N_3297,N_2337,N_2710);
xnor U3298 (N_3298,N_2201,N_2563);
nand U3299 (N_3299,N_2381,N_2250);
or U3300 (N_3300,N_2744,N_2021);
or U3301 (N_3301,N_2672,N_2046);
nor U3302 (N_3302,N_2973,N_2800);
xor U3303 (N_3303,N_2939,N_2589);
xnor U3304 (N_3304,N_2771,N_2243);
nand U3305 (N_3305,N_2893,N_2743);
xor U3306 (N_3306,N_2727,N_2218);
or U3307 (N_3307,N_2462,N_2565);
nand U3308 (N_3308,N_2705,N_2544);
nor U3309 (N_3309,N_2266,N_2761);
and U3310 (N_3310,N_2813,N_2480);
or U3311 (N_3311,N_2127,N_2485);
nand U3312 (N_3312,N_2546,N_2981);
and U3313 (N_3313,N_2689,N_2760);
or U3314 (N_3314,N_2277,N_2550);
nand U3315 (N_3315,N_2988,N_2223);
nor U3316 (N_3316,N_2278,N_2416);
and U3317 (N_3317,N_2924,N_2673);
nand U3318 (N_3318,N_2828,N_2121);
xnor U3319 (N_3319,N_2461,N_2539);
nor U3320 (N_3320,N_2287,N_2150);
nor U3321 (N_3321,N_2642,N_2499);
and U3322 (N_3322,N_2987,N_2211);
nor U3323 (N_3323,N_2984,N_2955);
or U3324 (N_3324,N_2323,N_2815);
and U3325 (N_3325,N_2818,N_2977);
or U3326 (N_3326,N_2606,N_2364);
or U3327 (N_3327,N_2737,N_2192);
xor U3328 (N_3328,N_2255,N_2293);
nand U3329 (N_3329,N_2738,N_2026);
or U3330 (N_3330,N_2372,N_2736);
nor U3331 (N_3331,N_2315,N_2477);
nand U3332 (N_3332,N_2216,N_2280);
nor U3333 (N_3333,N_2883,N_2043);
and U3334 (N_3334,N_2225,N_2531);
nand U3335 (N_3335,N_2353,N_2080);
or U3336 (N_3336,N_2081,N_2073);
and U3337 (N_3337,N_2763,N_2339);
nor U3338 (N_3338,N_2620,N_2527);
xor U3339 (N_3339,N_2299,N_2367);
nor U3340 (N_3340,N_2403,N_2641);
nor U3341 (N_3341,N_2360,N_2978);
and U3342 (N_3342,N_2902,N_2831);
nand U3343 (N_3343,N_2258,N_2035);
or U3344 (N_3344,N_2343,N_2667);
nor U3345 (N_3345,N_2714,N_2401);
and U3346 (N_3346,N_2392,N_2989);
xnor U3347 (N_3347,N_2166,N_2149);
or U3348 (N_3348,N_2889,N_2665);
and U3349 (N_3349,N_2325,N_2703);
and U3350 (N_3350,N_2425,N_2238);
nand U3351 (N_3351,N_2599,N_2526);
and U3352 (N_3352,N_2103,N_2953);
and U3353 (N_3353,N_2329,N_2024);
nor U3354 (N_3354,N_2119,N_2664);
and U3355 (N_3355,N_2729,N_2202);
and U3356 (N_3356,N_2867,N_2411);
nand U3357 (N_3357,N_2185,N_2459);
and U3358 (N_3358,N_2929,N_2552);
and U3359 (N_3359,N_2509,N_2069);
and U3360 (N_3360,N_2376,N_2949);
nand U3361 (N_3361,N_2224,N_2940);
and U3362 (N_3362,N_2256,N_2852);
nor U3363 (N_3363,N_2400,N_2109);
nand U3364 (N_3364,N_2130,N_2947);
xor U3365 (N_3365,N_2260,N_2436);
and U3366 (N_3366,N_2097,N_2670);
nand U3367 (N_3367,N_2786,N_2930);
or U3368 (N_3368,N_2141,N_2383);
nand U3369 (N_3369,N_2648,N_2915);
nor U3370 (N_3370,N_2231,N_2709);
xor U3371 (N_3371,N_2680,N_2830);
and U3372 (N_3372,N_2408,N_2438);
nor U3373 (N_3373,N_2851,N_2928);
and U3374 (N_3374,N_2471,N_2435);
or U3375 (N_3375,N_2054,N_2040);
or U3376 (N_3376,N_2568,N_2374);
nand U3377 (N_3377,N_2120,N_2503);
xor U3378 (N_3378,N_2405,N_2610);
nor U3379 (N_3379,N_2985,N_2604);
nand U3380 (N_3380,N_2084,N_2958);
xor U3381 (N_3381,N_2048,N_2942);
and U3382 (N_3382,N_2247,N_2657);
and U3383 (N_3383,N_2342,N_2835);
nand U3384 (N_3384,N_2528,N_2306);
and U3385 (N_3385,N_2690,N_2649);
nand U3386 (N_3386,N_2730,N_2646);
nand U3387 (N_3387,N_2228,N_2545);
xor U3388 (N_3388,N_2535,N_2937);
or U3389 (N_3389,N_2562,N_2716);
nor U3390 (N_3390,N_2361,N_2466);
and U3391 (N_3391,N_2507,N_2785);
nand U3392 (N_3392,N_2711,N_2212);
nor U3393 (N_3393,N_2511,N_2995);
and U3394 (N_3394,N_2859,N_2183);
nor U3395 (N_3395,N_2671,N_2619);
and U3396 (N_3396,N_2707,N_2219);
and U3397 (N_3397,N_2013,N_2593);
xor U3398 (N_3398,N_2193,N_2007);
xnor U3399 (N_3399,N_2585,N_2309);
xor U3400 (N_3400,N_2153,N_2843);
or U3401 (N_3401,N_2659,N_2140);
nor U3402 (N_3402,N_2189,N_2100);
nor U3403 (N_3403,N_2581,N_2651);
nand U3404 (N_3404,N_2242,N_2774);
and U3405 (N_3405,N_2501,N_2963);
nor U3406 (N_3406,N_2464,N_2096);
nand U3407 (N_3407,N_2064,N_2307);
nor U3408 (N_3408,N_2209,N_2724);
or U3409 (N_3409,N_2739,N_2913);
xor U3410 (N_3410,N_2352,N_2050);
nand U3411 (N_3411,N_2718,N_2885);
nor U3412 (N_3412,N_2793,N_2291);
and U3413 (N_3413,N_2869,N_2631);
nor U3414 (N_3414,N_2137,N_2085);
or U3415 (N_3415,N_2482,N_2327);
nor U3416 (N_3416,N_2808,N_2167);
nand U3417 (N_3417,N_2320,N_2916);
or U3418 (N_3418,N_2165,N_2698);
or U3419 (N_3419,N_2458,N_2377);
or U3420 (N_3420,N_2407,N_2888);
xor U3421 (N_3421,N_2559,N_2426);
nor U3422 (N_3422,N_2162,N_2602);
nand U3423 (N_3423,N_2708,N_2222);
or U3424 (N_3424,N_2014,N_2253);
nand U3425 (N_3425,N_2173,N_2434);
and U3426 (N_3426,N_2481,N_2872);
xor U3427 (N_3427,N_2182,N_2996);
nor U3428 (N_3428,N_2628,N_2177);
or U3429 (N_3429,N_2880,N_2241);
xnor U3430 (N_3430,N_2884,N_2018);
nor U3431 (N_3431,N_2204,N_2129);
or U3432 (N_3432,N_2030,N_2903);
xnor U3433 (N_3433,N_2108,N_2196);
and U3434 (N_3434,N_2529,N_2775);
xnor U3435 (N_3435,N_2113,N_2259);
nor U3436 (N_3436,N_2091,N_2500);
xnor U3437 (N_3437,N_2687,N_2923);
or U3438 (N_3438,N_2409,N_2588);
and U3439 (N_3439,N_2486,N_2412);
or U3440 (N_3440,N_2952,N_2005);
nand U3441 (N_3441,N_2780,N_2897);
or U3442 (N_3442,N_2819,N_2919);
nor U3443 (N_3443,N_2584,N_2015);
or U3444 (N_3444,N_2918,N_2677);
nor U3445 (N_3445,N_2838,N_2123);
nand U3446 (N_3446,N_2590,N_2457);
and U3447 (N_3447,N_2027,N_2001);
and U3448 (N_3448,N_2845,N_2925);
xor U3449 (N_3449,N_2092,N_2663);
and U3450 (N_3450,N_2395,N_2195);
nor U3451 (N_3451,N_2208,N_2041);
xnor U3452 (N_3452,N_2495,N_2777);
or U3453 (N_3453,N_2658,N_2279);
xor U3454 (N_3454,N_2000,N_2789);
nor U3455 (N_3455,N_2404,N_2448);
and U3456 (N_3456,N_2616,N_2803);
nand U3457 (N_3457,N_2490,N_2417);
and U3458 (N_3458,N_2463,N_2866);
nand U3459 (N_3459,N_2752,N_2860);
nand U3460 (N_3460,N_2029,N_2518);
nand U3461 (N_3461,N_2215,N_2399);
or U3462 (N_3462,N_2901,N_2220);
xor U3463 (N_3463,N_2906,N_2847);
xnor U3464 (N_3464,N_2799,N_2132);
nand U3465 (N_3465,N_2006,N_2152);
and U3466 (N_3466,N_2143,N_2393);
nand U3467 (N_3467,N_2493,N_2926);
xnor U3468 (N_3468,N_2305,N_2898);
and U3469 (N_3469,N_2164,N_2683);
nand U3470 (N_3470,N_2826,N_2285);
nand U3471 (N_3471,N_2180,N_2398);
or U3472 (N_3472,N_2443,N_2621);
xnor U3473 (N_3473,N_2911,N_2873);
nand U3474 (N_3474,N_2300,N_2369);
and U3475 (N_3475,N_2194,N_2652);
and U3476 (N_3476,N_2020,N_2944);
or U3477 (N_3477,N_2065,N_2839);
or U3478 (N_3478,N_2424,N_2240);
nor U3479 (N_3479,N_2575,N_2820);
and U3480 (N_3480,N_2770,N_2088);
nand U3481 (N_3481,N_2850,N_2858);
nand U3482 (N_3482,N_2678,N_2419);
nor U3483 (N_3483,N_2817,N_2335);
or U3484 (N_3484,N_2801,N_2945);
and U3485 (N_3485,N_2261,N_2791);
nand U3486 (N_3486,N_2175,N_2768);
nand U3487 (N_3487,N_2972,N_2450);
xnor U3488 (N_3488,N_2629,N_2894);
nand U3489 (N_3489,N_2868,N_2248);
nor U3490 (N_3490,N_2330,N_2491);
xor U3491 (N_3491,N_2313,N_2274);
nand U3492 (N_3492,N_2634,N_2921);
nor U3493 (N_3493,N_2617,N_2560);
and U3494 (N_3494,N_2444,N_2900);
nor U3495 (N_3495,N_2769,N_2449);
or U3496 (N_3496,N_2297,N_2753);
and U3497 (N_3497,N_2603,N_2414);
and U3498 (N_3498,N_2347,N_2571);
or U3499 (N_3499,N_2971,N_2052);
xnor U3500 (N_3500,N_2115,N_2072);
nor U3501 (N_3501,N_2949,N_2870);
nor U3502 (N_3502,N_2435,N_2812);
nand U3503 (N_3503,N_2201,N_2184);
and U3504 (N_3504,N_2490,N_2562);
nand U3505 (N_3505,N_2691,N_2053);
xnor U3506 (N_3506,N_2651,N_2574);
and U3507 (N_3507,N_2427,N_2067);
nand U3508 (N_3508,N_2393,N_2162);
nor U3509 (N_3509,N_2209,N_2012);
nor U3510 (N_3510,N_2920,N_2721);
nand U3511 (N_3511,N_2776,N_2936);
or U3512 (N_3512,N_2706,N_2672);
nand U3513 (N_3513,N_2768,N_2938);
xor U3514 (N_3514,N_2183,N_2560);
or U3515 (N_3515,N_2091,N_2031);
xnor U3516 (N_3516,N_2689,N_2124);
and U3517 (N_3517,N_2412,N_2979);
xor U3518 (N_3518,N_2998,N_2905);
nor U3519 (N_3519,N_2589,N_2761);
and U3520 (N_3520,N_2196,N_2379);
or U3521 (N_3521,N_2616,N_2988);
and U3522 (N_3522,N_2880,N_2083);
and U3523 (N_3523,N_2973,N_2469);
nor U3524 (N_3524,N_2548,N_2298);
nor U3525 (N_3525,N_2220,N_2039);
nand U3526 (N_3526,N_2341,N_2828);
nor U3527 (N_3527,N_2180,N_2120);
or U3528 (N_3528,N_2753,N_2639);
nor U3529 (N_3529,N_2425,N_2340);
and U3530 (N_3530,N_2151,N_2986);
or U3531 (N_3531,N_2704,N_2429);
nor U3532 (N_3532,N_2680,N_2790);
or U3533 (N_3533,N_2169,N_2410);
nand U3534 (N_3534,N_2994,N_2912);
and U3535 (N_3535,N_2524,N_2007);
nand U3536 (N_3536,N_2773,N_2541);
nor U3537 (N_3537,N_2469,N_2176);
xor U3538 (N_3538,N_2506,N_2307);
or U3539 (N_3539,N_2012,N_2442);
and U3540 (N_3540,N_2760,N_2363);
xor U3541 (N_3541,N_2378,N_2300);
xor U3542 (N_3542,N_2355,N_2164);
or U3543 (N_3543,N_2546,N_2185);
or U3544 (N_3544,N_2339,N_2196);
or U3545 (N_3545,N_2688,N_2470);
nand U3546 (N_3546,N_2156,N_2534);
nand U3547 (N_3547,N_2703,N_2564);
xor U3548 (N_3548,N_2513,N_2808);
or U3549 (N_3549,N_2631,N_2144);
nand U3550 (N_3550,N_2461,N_2968);
or U3551 (N_3551,N_2413,N_2605);
nor U3552 (N_3552,N_2843,N_2064);
xor U3553 (N_3553,N_2602,N_2057);
nor U3554 (N_3554,N_2237,N_2300);
xor U3555 (N_3555,N_2165,N_2129);
nor U3556 (N_3556,N_2877,N_2313);
nand U3557 (N_3557,N_2738,N_2004);
or U3558 (N_3558,N_2763,N_2005);
or U3559 (N_3559,N_2182,N_2003);
and U3560 (N_3560,N_2855,N_2084);
and U3561 (N_3561,N_2543,N_2496);
nor U3562 (N_3562,N_2037,N_2484);
or U3563 (N_3563,N_2007,N_2850);
xor U3564 (N_3564,N_2510,N_2548);
nand U3565 (N_3565,N_2250,N_2296);
and U3566 (N_3566,N_2724,N_2498);
nand U3567 (N_3567,N_2912,N_2385);
and U3568 (N_3568,N_2701,N_2598);
nor U3569 (N_3569,N_2143,N_2057);
nand U3570 (N_3570,N_2215,N_2203);
xor U3571 (N_3571,N_2060,N_2944);
nand U3572 (N_3572,N_2925,N_2359);
and U3573 (N_3573,N_2627,N_2976);
or U3574 (N_3574,N_2672,N_2375);
or U3575 (N_3575,N_2105,N_2257);
nor U3576 (N_3576,N_2911,N_2499);
or U3577 (N_3577,N_2881,N_2667);
xnor U3578 (N_3578,N_2496,N_2662);
and U3579 (N_3579,N_2239,N_2058);
nand U3580 (N_3580,N_2350,N_2677);
or U3581 (N_3581,N_2374,N_2154);
or U3582 (N_3582,N_2608,N_2041);
nand U3583 (N_3583,N_2273,N_2033);
xor U3584 (N_3584,N_2513,N_2222);
xor U3585 (N_3585,N_2647,N_2457);
nor U3586 (N_3586,N_2613,N_2389);
xnor U3587 (N_3587,N_2744,N_2043);
and U3588 (N_3588,N_2138,N_2021);
nor U3589 (N_3589,N_2904,N_2586);
nor U3590 (N_3590,N_2729,N_2805);
or U3591 (N_3591,N_2044,N_2771);
and U3592 (N_3592,N_2509,N_2094);
xnor U3593 (N_3593,N_2666,N_2923);
nand U3594 (N_3594,N_2103,N_2887);
and U3595 (N_3595,N_2506,N_2431);
nor U3596 (N_3596,N_2523,N_2207);
xnor U3597 (N_3597,N_2426,N_2715);
nand U3598 (N_3598,N_2460,N_2264);
xnor U3599 (N_3599,N_2425,N_2714);
or U3600 (N_3600,N_2533,N_2396);
xnor U3601 (N_3601,N_2015,N_2968);
nand U3602 (N_3602,N_2733,N_2601);
or U3603 (N_3603,N_2110,N_2246);
xor U3604 (N_3604,N_2622,N_2945);
and U3605 (N_3605,N_2830,N_2546);
xor U3606 (N_3606,N_2926,N_2068);
and U3607 (N_3607,N_2866,N_2077);
nor U3608 (N_3608,N_2583,N_2883);
xnor U3609 (N_3609,N_2793,N_2935);
nor U3610 (N_3610,N_2780,N_2890);
nand U3611 (N_3611,N_2535,N_2303);
and U3612 (N_3612,N_2770,N_2007);
and U3613 (N_3613,N_2681,N_2732);
xnor U3614 (N_3614,N_2286,N_2756);
xor U3615 (N_3615,N_2528,N_2840);
and U3616 (N_3616,N_2768,N_2413);
nor U3617 (N_3617,N_2128,N_2788);
and U3618 (N_3618,N_2314,N_2364);
and U3619 (N_3619,N_2984,N_2708);
nand U3620 (N_3620,N_2566,N_2372);
nand U3621 (N_3621,N_2786,N_2083);
nand U3622 (N_3622,N_2990,N_2391);
or U3623 (N_3623,N_2675,N_2176);
xor U3624 (N_3624,N_2398,N_2583);
xnor U3625 (N_3625,N_2604,N_2908);
xnor U3626 (N_3626,N_2819,N_2874);
nand U3627 (N_3627,N_2695,N_2382);
or U3628 (N_3628,N_2117,N_2688);
nand U3629 (N_3629,N_2519,N_2723);
xor U3630 (N_3630,N_2656,N_2593);
nand U3631 (N_3631,N_2924,N_2862);
or U3632 (N_3632,N_2079,N_2643);
nand U3633 (N_3633,N_2089,N_2545);
and U3634 (N_3634,N_2371,N_2867);
and U3635 (N_3635,N_2125,N_2783);
xnor U3636 (N_3636,N_2794,N_2495);
nand U3637 (N_3637,N_2693,N_2419);
nor U3638 (N_3638,N_2563,N_2776);
or U3639 (N_3639,N_2155,N_2841);
or U3640 (N_3640,N_2053,N_2953);
nor U3641 (N_3641,N_2705,N_2158);
xor U3642 (N_3642,N_2930,N_2879);
xor U3643 (N_3643,N_2127,N_2135);
nor U3644 (N_3644,N_2590,N_2837);
or U3645 (N_3645,N_2904,N_2399);
nor U3646 (N_3646,N_2974,N_2973);
nand U3647 (N_3647,N_2964,N_2780);
xor U3648 (N_3648,N_2850,N_2114);
nand U3649 (N_3649,N_2659,N_2383);
or U3650 (N_3650,N_2330,N_2049);
xor U3651 (N_3651,N_2107,N_2778);
nor U3652 (N_3652,N_2489,N_2368);
nor U3653 (N_3653,N_2882,N_2063);
nor U3654 (N_3654,N_2415,N_2627);
nand U3655 (N_3655,N_2585,N_2116);
nor U3656 (N_3656,N_2947,N_2154);
and U3657 (N_3657,N_2895,N_2173);
nand U3658 (N_3658,N_2796,N_2726);
nand U3659 (N_3659,N_2103,N_2244);
xnor U3660 (N_3660,N_2186,N_2662);
xor U3661 (N_3661,N_2830,N_2067);
and U3662 (N_3662,N_2705,N_2784);
and U3663 (N_3663,N_2636,N_2549);
nand U3664 (N_3664,N_2797,N_2785);
nand U3665 (N_3665,N_2607,N_2602);
and U3666 (N_3666,N_2369,N_2340);
and U3667 (N_3667,N_2294,N_2840);
nor U3668 (N_3668,N_2810,N_2290);
nand U3669 (N_3669,N_2915,N_2786);
and U3670 (N_3670,N_2495,N_2168);
xor U3671 (N_3671,N_2110,N_2135);
and U3672 (N_3672,N_2799,N_2832);
nor U3673 (N_3673,N_2082,N_2489);
xor U3674 (N_3674,N_2946,N_2799);
and U3675 (N_3675,N_2177,N_2185);
xor U3676 (N_3676,N_2535,N_2207);
xnor U3677 (N_3677,N_2914,N_2437);
nand U3678 (N_3678,N_2964,N_2537);
nand U3679 (N_3679,N_2539,N_2733);
and U3680 (N_3680,N_2196,N_2839);
and U3681 (N_3681,N_2934,N_2337);
xnor U3682 (N_3682,N_2927,N_2000);
and U3683 (N_3683,N_2699,N_2844);
nand U3684 (N_3684,N_2343,N_2732);
or U3685 (N_3685,N_2546,N_2603);
nand U3686 (N_3686,N_2063,N_2365);
and U3687 (N_3687,N_2559,N_2561);
nor U3688 (N_3688,N_2495,N_2609);
or U3689 (N_3689,N_2940,N_2785);
nand U3690 (N_3690,N_2298,N_2067);
or U3691 (N_3691,N_2307,N_2646);
nor U3692 (N_3692,N_2529,N_2251);
or U3693 (N_3693,N_2847,N_2720);
xnor U3694 (N_3694,N_2321,N_2770);
xor U3695 (N_3695,N_2853,N_2506);
nand U3696 (N_3696,N_2442,N_2403);
nand U3697 (N_3697,N_2636,N_2720);
xor U3698 (N_3698,N_2755,N_2649);
nor U3699 (N_3699,N_2709,N_2692);
nand U3700 (N_3700,N_2265,N_2252);
and U3701 (N_3701,N_2488,N_2286);
and U3702 (N_3702,N_2448,N_2364);
or U3703 (N_3703,N_2404,N_2706);
or U3704 (N_3704,N_2264,N_2239);
nand U3705 (N_3705,N_2587,N_2417);
nand U3706 (N_3706,N_2876,N_2707);
or U3707 (N_3707,N_2239,N_2149);
nor U3708 (N_3708,N_2948,N_2005);
or U3709 (N_3709,N_2659,N_2213);
nor U3710 (N_3710,N_2694,N_2302);
nor U3711 (N_3711,N_2333,N_2728);
and U3712 (N_3712,N_2866,N_2790);
xnor U3713 (N_3713,N_2621,N_2878);
nand U3714 (N_3714,N_2842,N_2219);
xnor U3715 (N_3715,N_2719,N_2369);
or U3716 (N_3716,N_2799,N_2201);
xnor U3717 (N_3717,N_2853,N_2718);
and U3718 (N_3718,N_2510,N_2267);
nor U3719 (N_3719,N_2004,N_2470);
nand U3720 (N_3720,N_2606,N_2466);
and U3721 (N_3721,N_2512,N_2767);
and U3722 (N_3722,N_2184,N_2175);
and U3723 (N_3723,N_2677,N_2166);
and U3724 (N_3724,N_2905,N_2915);
nor U3725 (N_3725,N_2327,N_2130);
nor U3726 (N_3726,N_2715,N_2859);
nand U3727 (N_3727,N_2867,N_2827);
nor U3728 (N_3728,N_2931,N_2612);
nor U3729 (N_3729,N_2394,N_2786);
and U3730 (N_3730,N_2109,N_2108);
xor U3731 (N_3731,N_2805,N_2370);
xor U3732 (N_3732,N_2439,N_2650);
and U3733 (N_3733,N_2569,N_2815);
and U3734 (N_3734,N_2080,N_2573);
nor U3735 (N_3735,N_2091,N_2640);
and U3736 (N_3736,N_2981,N_2021);
xnor U3737 (N_3737,N_2399,N_2547);
or U3738 (N_3738,N_2145,N_2605);
or U3739 (N_3739,N_2939,N_2433);
and U3740 (N_3740,N_2010,N_2685);
nand U3741 (N_3741,N_2477,N_2985);
and U3742 (N_3742,N_2541,N_2506);
nor U3743 (N_3743,N_2270,N_2411);
nor U3744 (N_3744,N_2060,N_2057);
nand U3745 (N_3745,N_2679,N_2655);
or U3746 (N_3746,N_2826,N_2912);
nor U3747 (N_3747,N_2600,N_2755);
xor U3748 (N_3748,N_2196,N_2179);
nand U3749 (N_3749,N_2985,N_2303);
and U3750 (N_3750,N_2774,N_2905);
or U3751 (N_3751,N_2591,N_2998);
or U3752 (N_3752,N_2446,N_2010);
nor U3753 (N_3753,N_2931,N_2491);
or U3754 (N_3754,N_2125,N_2225);
or U3755 (N_3755,N_2496,N_2371);
xnor U3756 (N_3756,N_2517,N_2220);
nand U3757 (N_3757,N_2257,N_2050);
nand U3758 (N_3758,N_2262,N_2083);
nand U3759 (N_3759,N_2768,N_2205);
or U3760 (N_3760,N_2643,N_2213);
nand U3761 (N_3761,N_2389,N_2325);
and U3762 (N_3762,N_2837,N_2932);
nor U3763 (N_3763,N_2230,N_2556);
and U3764 (N_3764,N_2624,N_2472);
and U3765 (N_3765,N_2634,N_2822);
nand U3766 (N_3766,N_2455,N_2887);
nand U3767 (N_3767,N_2774,N_2408);
or U3768 (N_3768,N_2926,N_2479);
or U3769 (N_3769,N_2172,N_2983);
and U3770 (N_3770,N_2217,N_2608);
nor U3771 (N_3771,N_2948,N_2946);
nand U3772 (N_3772,N_2452,N_2482);
nand U3773 (N_3773,N_2666,N_2478);
or U3774 (N_3774,N_2472,N_2565);
nor U3775 (N_3775,N_2378,N_2149);
xor U3776 (N_3776,N_2878,N_2224);
or U3777 (N_3777,N_2362,N_2959);
nor U3778 (N_3778,N_2581,N_2016);
and U3779 (N_3779,N_2147,N_2333);
xor U3780 (N_3780,N_2412,N_2883);
nor U3781 (N_3781,N_2332,N_2710);
or U3782 (N_3782,N_2694,N_2923);
nor U3783 (N_3783,N_2155,N_2564);
nor U3784 (N_3784,N_2642,N_2086);
xor U3785 (N_3785,N_2534,N_2885);
and U3786 (N_3786,N_2045,N_2165);
nor U3787 (N_3787,N_2952,N_2870);
xor U3788 (N_3788,N_2031,N_2955);
and U3789 (N_3789,N_2821,N_2683);
or U3790 (N_3790,N_2355,N_2622);
or U3791 (N_3791,N_2570,N_2745);
or U3792 (N_3792,N_2074,N_2082);
and U3793 (N_3793,N_2668,N_2710);
nor U3794 (N_3794,N_2466,N_2117);
nor U3795 (N_3795,N_2984,N_2783);
nand U3796 (N_3796,N_2948,N_2762);
nand U3797 (N_3797,N_2427,N_2820);
and U3798 (N_3798,N_2740,N_2093);
and U3799 (N_3799,N_2629,N_2409);
nand U3800 (N_3800,N_2930,N_2526);
and U3801 (N_3801,N_2246,N_2302);
or U3802 (N_3802,N_2362,N_2077);
or U3803 (N_3803,N_2712,N_2974);
and U3804 (N_3804,N_2937,N_2928);
and U3805 (N_3805,N_2342,N_2078);
and U3806 (N_3806,N_2036,N_2372);
nand U3807 (N_3807,N_2197,N_2024);
nor U3808 (N_3808,N_2930,N_2483);
or U3809 (N_3809,N_2759,N_2618);
nand U3810 (N_3810,N_2998,N_2347);
nor U3811 (N_3811,N_2571,N_2782);
or U3812 (N_3812,N_2807,N_2618);
and U3813 (N_3813,N_2282,N_2454);
nand U3814 (N_3814,N_2132,N_2600);
nand U3815 (N_3815,N_2274,N_2124);
or U3816 (N_3816,N_2468,N_2452);
or U3817 (N_3817,N_2748,N_2574);
nor U3818 (N_3818,N_2230,N_2353);
and U3819 (N_3819,N_2551,N_2768);
nand U3820 (N_3820,N_2475,N_2622);
xnor U3821 (N_3821,N_2190,N_2552);
and U3822 (N_3822,N_2078,N_2564);
or U3823 (N_3823,N_2616,N_2236);
or U3824 (N_3824,N_2463,N_2709);
nand U3825 (N_3825,N_2201,N_2814);
xnor U3826 (N_3826,N_2262,N_2759);
and U3827 (N_3827,N_2948,N_2012);
and U3828 (N_3828,N_2397,N_2495);
and U3829 (N_3829,N_2328,N_2115);
xnor U3830 (N_3830,N_2510,N_2296);
nor U3831 (N_3831,N_2227,N_2172);
nor U3832 (N_3832,N_2648,N_2011);
nand U3833 (N_3833,N_2836,N_2855);
nor U3834 (N_3834,N_2355,N_2926);
nand U3835 (N_3835,N_2702,N_2718);
or U3836 (N_3836,N_2547,N_2774);
xnor U3837 (N_3837,N_2450,N_2324);
and U3838 (N_3838,N_2581,N_2577);
xnor U3839 (N_3839,N_2230,N_2745);
nor U3840 (N_3840,N_2356,N_2838);
or U3841 (N_3841,N_2594,N_2247);
xor U3842 (N_3842,N_2584,N_2944);
xnor U3843 (N_3843,N_2260,N_2939);
xnor U3844 (N_3844,N_2381,N_2545);
xnor U3845 (N_3845,N_2767,N_2610);
or U3846 (N_3846,N_2581,N_2626);
or U3847 (N_3847,N_2923,N_2946);
or U3848 (N_3848,N_2950,N_2389);
nand U3849 (N_3849,N_2851,N_2476);
and U3850 (N_3850,N_2266,N_2949);
xor U3851 (N_3851,N_2456,N_2990);
nand U3852 (N_3852,N_2559,N_2147);
and U3853 (N_3853,N_2261,N_2705);
xnor U3854 (N_3854,N_2304,N_2031);
nand U3855 (N_3855,N_2603,N_2621);
nand U3856 (N_3856,N_2501,N_2838);
xnor U3857 (N_3857,N_2424,N_2597);
nand U3858 (N_3858,N_2896,N_2020);
nand U3859 (N_3859,N_2893,N_2355);
xnor U3860 (N_3860,N_2482,N_2621);
and U3861 (N_3861,N_2025,N_2375);
nor U3862 (N_3862,N_2577,N_2251);
xor U3863 (N_3863,N_2160,N_2529);
nand U3864 (N_3864,N_2398,N_2743);
and U3865 (N_3865,N_2970,N_2384);
nand U3866 (N_3866,N_2893,N_2530);
nor U3867 (N_3867,N_2588,N_2325);
xor U3868 (N_3868,N_2228,N_2580);
nand U3869 (N_3869,N_2416,N_2912);
xor U3870 (N_3870,N_2310,N_2543);
or U3871 (N_3871,N_2076,N_2432);
xor U3872 (N_3872,N_2907,N_2696);
nand U3873 (N_3873,N_2007,N_2111);
nor U3874 (N_3874,N_2224,N_2087);
xnor U3875 (N_3875,N_2857,N_2569);
nor U3876 (N_3876,N_2406,N_2734);
or U3877 (N_3877,N_2489,N_2369);
xnor U3878 (N_3878,N_2980,N_2131);
xnor U3879 (N_3879,N_2286,N_2653);
or U3880 (N_3880,N_2113,N_2937);
nor U3881 (N_3881,N_2504,N_2999);
nor U3882 (N_3882,N_2010,N_2786);
nor U3883 (N_3883,N_2378,N_2166);
nand U3884 (N_3884,N_2036,N_2139);
nor U3885 (N_3885,N_2966,N_2749);
nand U3886 (N_3886,N_2088,N_2129);
nor U3887 (N_3887,N_2803,N_2326);
or U3888 (N_3888,N_2766,N_2195);
or U3889 (N_3889,N_2668,N_2359);
nor U3890 (N_3890,N_2100,N_2225);
nor U3891 (N_3891,N_2869,N_2557);
or U3892 (N_3892,N_2243,N_2670);
or U3893 (N_3893,N_2947,N_2056);
and U3894 (N_3894,N_2181,N_2023);
and U3895 (N_3895,N_2333,N_2141);
or U3896 (N_3896,N_2911,N_2104);
and U3897 (N_3897,N_2007,N_2388);
or U3898 (N_3898,N_2217,N_2970);
nor U3899 (N_3899,N_2739,N_2256);
and U3900 (N_3900,N_2596,N_2514);
and U3901 (N_3901,N_2873,N_2294);
or U3902 (N_3902,N_2734,N_2055);
nor U3903 (N_3903,N_2301,N_2814);
nand U3904 (N_3904,N_2097,N_2190);
xnor U3905 (N_3905,N_2549,N_2752);
xor U3906 (N_3906,N_2755,N_2371);
or U3907 (N_3907,N_2759,N_2702);
or U3908 (N_3908,N_2992,N_2734);
xor U3909 (N_3909,N_2857,N_2941);
nor U3910 (N_3910,N_2200,N_2511);
xor U3911 (N_3911,N_2968,N_2797);
nor U3912 (N_3912,N_2528,N_2909);
nor U3913 (N_3913,N_2268,N_2099);
and U3914 (N_3914,N_2587,N_2269);
nand U3915 (N_3915,N_2578,N_2148);
or U3916 (N_3916,N_2464,N_2359);
nand U3917 (N_3917,N_2652,N_2923);
nand U3918 (N_3918,N_2552,N_2958);
nor U3919 (N_3919,N_2587,N_2752);
or U3920 (N_3920,N_2285,N_2130);
or U3921 (N_3921,N_2693,N_2488);
nor U3922 (N_3922,N_2447,N_2096);
nand U3923 (N_3923,N_2290,N_2572);
xor U3924 (N_3924,N_2697,N_2713);
or U3925 (N_3925,N_2586,N_2311);
or U3926 (N_3926,N_2276,N_2980);
or U3927 (N_3927,N_2281,N_2638);
nor U3928 (N_3928,N_2782,N_2854);
nand U3929 (N_3929,N_2512,N_2539);
or U3930 (N_3930,N_2042,N_2326);
or U3931 (N_3931,N_2257,N_2141);
nand U3932 (N_3932,N_2541,N_2533);
nor U3933 (N_3933,N_2802,N_2425);
or U3934 (N_3934,N_2289,N_2500);
and U3935 (N_3935,N_2927,N_2440);
and U3936 (N_3936,N_2343,N_2085);
xnor U3937 (N_3937,N_2789,N_2123);
and U3938 (N_3938,N_2451,N_2676);
or U3939 (N_3939,N_2823,N_2248);
and U3940 (N_3940,N_2800,N_2926);
xor U3941 (N_3941,N_2610,N_2696);
xor U3942 (N_3942,N_2961,N_2379);
nand U3943 (N_3943,N_2930,N_2638);
nand U3944 (N_3944,N_2580,N_2570);
nor U3945 (N_3945,N_2286,N_2743);
nor U3946 (N_3946,N_2385,N_2578);
xnor U3947 (N_3947,N_2302,N_2248);
nand U3948 (N_3948,N_2579,N_2038);
xnor U3949 (N_3949,N_2994,N_2849);
and U3950 (N_3950,N_2486,N_2969);
or U3951 (N_3951,N_2955,N_2037);
or U3952 (N_3952,N_2834,N_2533);
or U3953 (N_3953,N_2560,N_2616);
nor U3954 (N_3954,N_2382,N_2458);
nand U3955 (N_3955,N_2123,N_2051);
or U3956 (N_3956,N_2258,N_2064);
nor U3957 (N_3957,N_2050,N_2000);
nor U3958 (N_3958,N_2700,N_2181);
or U3959 (N_3959,N_2139,N_2606);
or U3960 (N_3960,N_2868,N_2376);
nand U3961 (N_3961,N_2324,N_2139);
nand U3962 (N_3962,N_2593,N_2074);
and U3963 (N_3963,N_2325,N_2062);
or U3964 (N_3964,N_2205,N_2184);
or U3965 (N_3965,N_2296,N_2009);
or U3966 (N_3966,N_2496,N_2042);
xor U3967 (N_3967,N_2420,N_2779);
xnor U3968 (N_3968,N_2401,N_2670);
xnor U3969 (N_3969,N_2407,N_2908);
or U3970 (N_3970,N_2890,N_2487);
and U3971 (N_3971,N_2989,N_2375);
and U3972 (N_3972,N_2371,N_2287);
or U3973 (N_3973,N_2607,N_2065);
and U3974 (N_3974,N_2412,N_2206);
nor U3975 (N_3975,N_2363,N_2470);
xnor U3976 (N_3976,N_2805,N_2820);
or U3977 (N_3977,N_2983,N_2154);
or U3978 (N_3978,N_2272,N_2550);
nor U3979 (N_3979,N_2836,N_2552);
nor U3980 (N_3980,N_2588,N_2690);
xor U3981 (N_3981,N_2930,N_2174);
nor U3982 (N_3982,N_2820,N_2704);
xnor U3983 (N_3983,N_2613,N_2673);
and U3984 (N_3984,N_2058,N_2917);
and U3985 (N_3985,N_2887,N_2581);
and U3986 (N_3986,N_2505,N_2085);
xnor U3987 (N_3987,N_2451,N_2483);
xnor U3988 (N_3988,N_2380,N_2325);
and U3989 (N_3989,N_2068,N_2647);
xor U3990 (N_3990,N_2587,N_2320);
or U3991 (N_3991,N_2480,N_2804);
or U3992 (N_3992,N_2795,N_2052);
and U3993 (N_3993,N_2613,N_2426);
nand U3994 (N_3994,N_2299,N_2758);
xor U3995 (N_3995,N_2296,N_2641);
or U3996 (N_3996,N_2515,N_2316);
or U3997 (N_3997,N_2250,N_2833);
or U3998 (N_3998,N_2916,N_2602);
nor U3999 (N_3999,N_2487,N_2048);
nand U4000 (N_4000,N_3072,N_3600);
or U4001 (N_4001,N_3017,N_3975);
nand U4002 (N_4002,N_3752,N_3381);
and U4003 (N_4003,N_3265,N_3134);
xor U4004 (N_4004,N_3048,N_3660);
and U4005 (N_4005,N_3662,N_3497);
nor U4006 (N_4006,N_3868,N_3152);
and U4007 (N_4007,N_3454,N_3139);
nand U4008 (N_4008,N_3615,N_3121);
and U4009 (N_4009,N_3866,N_3698);
xnor U4010 (N_4010,N_3018,N_3391);
nor U4011 (N_4011,N_3505,N_3186);
xor U4012 (N_4012,N_3861,N_3179);
xor U4013 (N_4013,N_3198,N_3478);
and U4014 (N_4014,N_3398,N_3234);
nand U4015 (N_4015,N_3718,N_3770);
and U4016 (N_4016,N_3298,N_3292);
and U4017 (N_4017,N_3098,N_3605);
or U4018 (N_4018,N_3514,N_3541);
xor U4019 (N_4019,N_3390,N_3342);
nor U4020 (N_4020,N_3372,N_3058);
or U4021 (N_4021,N_3320,N_3801);
nand U4022 (N_4022,N_3784,N_3754);
xor U4023 (N_4023,N_3189,N_3503);
and U4024 (N_4024,N_3827,N_3316);
nor U4025 (N_4025,N_3969,N_3830);
and U4026 (N_4026,N_3167,N_3879);
nor U4027 (N_4027,N_3275,N_3688);
or U4028 (N_4028,N_3252,N_3743);
and U4029 (N_4029,N_3444,N_3021);
and U4030 (N_4030,N_3011,N_3691);
nor U4031 (N_4031,N_3719,N_3218);
nor U4032 (N_4032,N_3377,N_3054);
nor U4033 (N_4033,N_3565,N_3217);
nor U4034 (N_4034,N_3838,N_3411);
and U4035 (N_4035,N_3038,N_3271);
or U4036 (N_4036,N_3985,N_3219);
nor U4037 (N_4037,N_3159,N_3279);
and U4038 (N_4038,N_3535,N_3241);
or U4039 (N_4039,N_3629,N_3183);
nor U4040 (N_4040,N_3309,N_3539);
and U4041 (N_4041,N_3091,N_3376);
nand U4042 (N_4042,N_3588,N_3124);
xor U4043 (N_4043,N_3208,N_3071);
nand U4044 (N_4044,N_3233,N_3761);
and U4045 (N_4045,N_3317,N_3482);
xnor U4046 (N_4046,N_3434,N_3191);
xnor U4047 (N_4047,N_3206,N_3773);
xor U4048 (N_4048,N_3913,N_3158);
and U4049 (N_4049,N_3424,N_3926);
or U4050 (N_4050,N_3820,N_3181);
or U4051 (N_4051,N_3173,N_3710);
xnor U4052 (N_4052,N_3070,N_3865);
nor U4053 (N_4053,N_3612,N_3287);
nor U4054 (N_4054,N_3822,N_3848);
xnor U4055 (N_4055,N_3805,N_3310);
and U4056 (N_4056,N_3966,N_3724);
nor U4057 (N_4057,N_3803,N_3509);
xor U4058 (N_4058,N_3731,N_3188);
or U4059 (N_4059,N_3350,N_3367);
nor U4060 (N_4060,N_3263,N_3560);
or U4061 (N_4061,N_3620,N_3006);
nor U4062 (N_4062,N_3751,N_3193);
nand U4063 (N_4063,N_3105,N_3380);
or U4064 (N_4064,N_3452,N_3523);
or U4065 (N_4065,N_3646,N_3516);
nand U4066 (N_4066,N_3699,N_3517);
nand U4067 (N_4067,N_3502,N_3487);
and U4068 (N_4068,N_3645,N_3543);
or U4069 (N_4069,N_3847,N_3477);
or U4070 (N_4070,N_3603,N_3997);
or U4071 (N_4071,N_3722,N_3389);
or U4072 (N_4072,N_3694,N_3468);
nor U4073 (N_4073,N_3849,N_3131);
nor U4074 (N_4074,N_3035,N_3397);
or U4075 (N_4075,N_3222,N_3932);
nor U4076 (N_4076,N_3883,N_3570);
xor U4077 (N_4077,N_3313,N_3613);
and U4078 (N_4078,N_3169,N_3409);
and U4079 (N_4079,N_3976,N_3033);
or U4080 (N_4080,N_3093,N_3163);
or U4081 (N_4081,N_3548,N_3529);
xnor U4082 (N_4082,N_3150,N_3908);
or U4083 (N_4083,N_3610,N_3851);
or U4084 (N_4084,N_3869,N_3863);
xnor U4085 (N_4085,N_3488,N_3546);
xor U4086 (N_4086,N_3427,N_3388);
nor U4087 (N_4087,N_3069,N_3671);
or U4088 (N_4088,N_3980,N_3418);
nor U4089 (N_4089,N_3775,N_3513);
or U4090 (N_4090,N_3445,N_3119);
nand U4091 (N_4091,N_3531,N_3576);
and U4092 (N_4092,N_3666,N_3571);
xnor U4093 (N_4093,N_3507,N_3165);
and U4094 (N_4094,N_3792,N_3675);
nand U4095 (N_4095,N_3184,N_3286);
and U4096 (N_4096,N_3045,N_3564);
or U4097 (N_4097,N_3392,N_3239);
or U4098 (N_4098,N_3034,N_3364);
nand U4099 (N_4099,N_3484,N_3755);
nor U4100 (N_4100,N_3542,N_3358);
nor U4101 (N_4101,N_3097,N_3850);
nand U4102 (N_4102,N_3981,N_3387);
nor U4103 (N_4103,N_3669,N_3592);
and U4104 (N_4104,N_3476,N_3986);
or U4105 (N_4105,N_3566,N_3272);
nor U4106 (N_4106,N_3261,N_3288);
or U4107 (N_4107,N_3974,N_3088);
nand U4108 (N_4108,N_3559,N_3875);
xor U4109 (N_4109,N_3510,N_3050);
xor U4110 (N_4110,N_3325,N_3324);
or U4111 (N_4111,N_3057,N_3664);
nor U4112 (N_4112,N_3900,N_3789);
xnor U4113 (N_4113,N_3899,N_3971);
xnor U4114 (N_4114,N_3927,N_3500);
and U4115 (N_4115,N_3598,N_3678);
xnor U4116 (N_4116,N_3774,N_3897);
or U4117 (N_4117,N_3228,N_3260);
nand U4118 (N_4118,N_3793,N_3352);
or U4119 (N_4119,N_3416,N_3028);
nor U4120 (N_4120,N_3084,N_3676);
nand U4121 (N_4121,N_3253,N_3151);
and U4122 (N_4122,N_3415,N_3983);
xor U4123 (N_4123,N_3022,N_3723);
nand U4124 (N_4124,N_3649,N_3878);
xnor U4125 (N_4125,N_3819,N_3037);
or U4126 (N_4126,N_3652,N_3065);
xor U4127 (N_4127,N_3496,N_3931);
or U4128 (N_4128,N_3914,N_3008);
and U4129 (N_4129,N_3683,N_3420);
and U4130 (N_4130,N_3806,N_3371);
xor U4131 (N_4131,N_3906,N_3475);
nand U4132 (N_4132,N_3385,N_3685);
nor U4133 (N_4133,N_3606,N_3696);
xor U4134 (N_4134,N_3122,N_3361);
xor U4135 (N_4135,N_3319,N_3705);
nand U4136 (N_4136,N_3891,N_3795);
nor U4137 (N_4137,N_3082,N_3378);
and U4138 (N_4138,N_3410,N_3843);
nand U4139 (N_4139,N_3277,N_3573);
xnor U4140 (N_4140,N_3032,N_3757);
and U4141 (N_4141,N_3818,N_3711);
and U4142 (N_4142,N_3280,N_3951);
or U4143 (N_4143,N_3824,N_3563);
or U4144 (N_4144,N_3758,N_3481);
xnor U4145 (N_4145,N_3704,N_3499);
nand U4146 (N_4146,N_3946,N_3817);
or U4147 (N_4147,N_3102,N_3967);
and U4148 (N_4148,N_3644,N_3010);
nand U4149 (N_4149,N_3572,N_3335);
xnor U4150 (N_4150,N_3264,N_3457);
or U4151 (N_4151,N_3024,N_3668);
xor U4152 (N_4152,N_3842,N_3489);
nor U4153 (N_4153,N_3422,N_3766);
nor U4154 (N_4154,N_3938,N_3880);
or U4155 (N_4155,N_3641,N_3905);
and U4156 (N_4156,N_3740,N_3759);
or U4157 (N_4157,N_3485,N_3903);
nor U4158 (N_4158,N_3577,N_3321);
nand U4159 (N_4159,N_3349,N_3601);
nor U4160 (N_4160,N_3407,N_3845);
nand U4161 (N_4161,N_3441,N_3658);
nor U4162 (N_4162,N_3290,N_3305);
xnor U4163 (N_4163,N_3395,N_3844);
nor U4164 (N_4164,N_3232,N_3673);
or U4165 (N_4165,N_3622,N_3994);
and U4166 (N_4166,N_3205,N_3004);
xnor U4167 (N_4167,N_3602,N_3744);
xnor U4168 (N_4168,N_3747,N_3060);
nand U4169 (N_4169,N_3061,N_3405);
nand U4170 (N_4170,N_3901,N_3709);
and U4171 (N_4171,N_3582,N_3240);
xor U4172 (N_4172,N_3968,N_3829);
or U4173 (N_4173,N_3832,N_3249);
or U4174 (N_4174,N_3810,N_3928);
xnor U4175 (N_4175,N_3142,N_3493);
and U4176 (N_4176,N_3384,N_3703);
nand U4177 (N_4177,N_3989,N_3130);
nand U4178 (N_4178,N_3254,N_3657);
nor U4179 (N_4179,N_3977,N_3632);
nor U4180 (N_4180,N_3182,N_3552);
or U4181 (N_4181,N_3778,N_3581);
nor U4182 (N_4182,N_3431,N_3465);
nor U4183 (N_4183,N_3283,N_3562);
or U4184 (N_4184,N_3874,N_3047);
nand U4185 (N_4185,N_3972,N_3929);
or U4186 (N_4186,N_3987,N_3199);
or U4187 (N_4187,N_3619,N_3939);
nor U4188 (N_4188,N_3225,N_3745);
xor U4189 (N_4189,N_3423,N_3351);
and U4190 (N_4190,N_3215,N_3170);
nor U4191 (N_4191,N_3211,N_3593);
or U4192 (N_4192,N_3715,N_3382);
and U4193 (N_4193,N_3519,N_3174);
and U4194 (N_4194,N_3790,N_3002);
nand U4195 (N_4195,N_3278,N_3196);
nor U4196 (N_4196,N_3781,N_3567);
nand U4197 (N_4197,N_3877,N_3762);
xor U4198 (N_4198,N_3144,N_3876);
xnor U4199 (N_4199,N_3052,N_3894);
xnor U4200 (N_4200,N_3295,N_3083);
and U4201 (N_4201,N_3794,N_3814);
and U4202 (N_4202,N_3628,N_3296);
xor U4203 (N_4203,N_3362,N_3648);
or U4204 (N_4204,N_3242,N_3852);
nor U4205 (N_4205,N_3544,N_3125);
nor U4206 (N_4206,N_3354,N_3412);
and U4207 (N_4207,N_3443,N_3729);
nor U4208 (N_4208,N_3005,N_3149);
nor U4209 (N_4209,N_3962,N_3432);
nor U4210 (N_4210,N_3092,N_3734);
nor U4211 (N_4211,N_3348,N_3248);
nor U4212 (N_4212,N_3360,N_3322);
xor U4213 (N_4213,N_3950,N_3727);
xnor U4214 (N_4214,N_3767,N_3433);
nand U4215 (N_4215,N_3943,N_3530);
nor U4216 (N_4216,N_3942,N_3132);
xor U4217 (N_4217,N_3802,N_3919);
or U4218 (N_4218,N_3236,N_3785);
nor U4219 (N_4219,N_3569,N_3129);
or U4220 (N_4220,N_3467,N_3937);
and U4221 (N_4221,N_3941,N_3101);
nand U4222 (N_4222,N_3428,N_3749);
xor U4223 (N_4223,N_3074,N_3138);
or U4224 (N_4224,N_3145,N_3812);
or U4225 (N_4225,N_3616,N_3210);
nor U4226 (N_4226,N_3935,N_3285);
or U4227 (N_4227,N_3627,N_3587);
xor U4228 (N_4228,N_3902,N_3608);
nor U4229 (N_4229,N_3545,N_3399);
nand U4230 (N_4230,N_3979,N_3661);
nand U4231 (N_4231,N_3365,N_3635);
nor U4232 (N_4232,N_3912,N_3995);
nor U4233 (N_4233,N_3654,N_3925);
nor U4234 (N_4234,N_3453,N_3674);
and U4235 (N_4235,N_3553,N_3959);
nor U4236 (N_4236,N_3742,N_3448);
or U4237 (N_4237,N_3659,N_3996);
or U4238 (N_4238,N_3557,N_3282);
and U4239 (N_4239,N_3156,N_3214);
xor U4240 (N_4240,N_3599,N_3194);
xor U4241 (N_4241,N_3491,N_3302);
nor U4242 (N_4242,N_3213,N_3728);
nand U4243 (N_4243,N_3117,N_3811);
or U4244 (N_4244,N_3312,N_3791);
nor U4245 (N_4245,N_3857,N_3737);
or U4246 (N_4246,N_3769,N_3164);
nand U4247 (N_4247,N_3701,N_3888);
nor U4248 (N_4248,N_3884,N_3854);
nand U4249 (N_4249,N_3595,N_3373);
xor U4250 (N_4250,N_3948,N_3345);
nor U4251 (N_4251,N_3294,N_3930);
xor U4252 (N_4252,N_3799,N_3647);
or U4253 (N_4253,N_3245,N_3259);
and U4254 (N_4254,N_3227,N_3267);
nor U4255 (N_4255,N_3561,N_3402);
xor U4256 (N_4256,N_3355,N_3999);
nand U4257 (N_4257,N_3417,N_3554);
and U4258 (N_4258,N_3575,N_3821);
nor U4259 (N_4259,N_3772,N_3687);
nand U4260 (N_4260,N_3998,N_3501);
xor U4261 (N_4261,N_3735,N_3104);
or U4262 (N_4262,N_3625,N_3515);
nor U4263 (N_4263,N_3590,N_3043);
nor U4264 (N_4264,N_3584,N_3221);
and U4265 (N_4265,N_3978,N_3089);
nand U4266 (N_4266,N_3127,N_3682);
nor U4267 (N_4267,N_3339,N_3113);
or U4268 (N_4268,N_3421,N_3695);
nor U4269 (N_4269,N_3306,N_3146);
xnor U4270 (N_4270,N_3760,N_3403);
nor U4271 (N_4271,N_3094,N_3076);
nor U4272 (N_4272,N_3116,N_3430);
xor U4273 (N_4273,N_3041,N_3859);
and U4274 (N_4274,N_3716,N_3001);
nand U4275 (N_4275,N_3436,N_3898);
nor U4276 (N_4276,N_3244,N_3965);
xor U4277 (N_4277,N_3988,N_3982);
nor U4278 (N_4278,N_3807,N_3623);
and U4279 (N_4279,N_3229,N_3640);
or U4280 (N_4280,N_3733,N_3025);
nand U4281 (N_4281,N_3585,N_3255);
nor U4282 (N_4282,N_3887,N_3956);
nor U4283 (N_4283,N_3330,N_3250);
and U4284 (N_4284,N_3702,N_3068);
and U4285 (N_4285,N_3400,N_3301);
nor U4286 (N_4286,N_3099,N_3763);
nand U4287 (N_4287,N_3200,N_3029);
or U4288 (N_4288,N_3413,N_3970);
and U4289 (N_4289,N_3141,N_3918);
xnor U4290 (N_4290,N_3708,N_3066);
or U4291 (N_4291,N_3472,N_3178);
nand U4292 (N_4292,N_3512,N_3204);
nor U4293 (N_4293,N_3356,N_3426);
nor U4294 (N_4294,N_3212,N_3090);
nor U4295 (N_4295,N_3955,N_3012);
xor U4296 (N_4296,N_3223,N_3314);
xor U4297 (N_4297,N_3009,N_3256);
xor U4298 (N_4298,N_3040,N_3787);
or U4299 (N_4299,N_3055,N_3148);
or U4300 (N_4300,N_3825,N_3527);
or U4301 (N_4301,N_3663,N_3386);
xor U4302 (N_4302,N_3934,N_3651);
and U4303 (N_4303,N_3776,N_3538);
xnor U4304 (N_4304,N_3808,N_3161);
nand U4305 (N_4305,N_3344,N_3853);
or U4306 (N_4306,N_3379,N_3308);
and U4307 (N_4307,N_3329,N_3013);
or U4308 (N_4308,N_3872,N_3521);
nor U4309 (N_4309,N_3246,N_3195);
nor U4310 (N_4310,N_3000,N_3067);
xor U4311 (N_4311,N_3408,N_3128);
nor U4312 (N_4312,N_3015,N_3536);
nor U4313 (N_4313,N_3520,N_3108);
xnor U4314 (N_4314,N_3604,N_3924);
or U4315 (N_4315,N_3534,N_3783);
nor U4316 (N_4316,N_3607,N_3257);
and U4317 (N_4317,N_3518,N_3166);
nor U4318 (N_4318,N_3079,N_3961);
or U4319 (N_4319,N_3077,N_3168);
xor U4320 (N_4320,N_3680,N_3933);
or U4321 (N_4321,N_3580,N_3780);
xnor U4322 (N_4322,N_3591,N_3419);
nand U4323 (N_4323,N_3123,N_3677);
or U4324 (N_4324,N_3732,N_3885);
nor U4325 (N_4325,N_3533,N_3450);
xor U4326 (N_4326,N_3800,N_3686);
xnor U4327 (N_4327,N_3177,N_3126);
nor U4328 (N_4328,N_3611,N_3895);
or U4329 (N_4329,N_3036,N_3464);
or U4330 (N_4330,N_3442,N_3917);
or U4331 (N_4331,N_3840,N_3023);
xor U4332 (N_4332,N_3947,N_3837);
nor U4333 (N_4333,N_3867,N_3506);
or U4334 (N_4334,N_3366,N_3638);
and U4335 (N_4335,N_3712,N_3087);
xor U4336 (N_4336,N_3637,N_3291);
nor U4337 (N_4337,N_3353,N_3369);
nor U4338 (N_4338,N_3550,N_3080);
or U4339 (N_4339,N_3782,N_3846);
nand U4340 (N_4340,N_3393,N_3266);
nand U4341 (N_4341,N_3864,N_3993);
xnor U4342 (N_4342,N_3338,N_3537);
nor U4343 (N_4343,N_3449,N_3343);
or U4344 (N_4344,N_3202,N_3268);
nand U4345 (N_4345,N_3315,N_3653);
or U4346 (N_4346,N_3307,N_3636);
nand U4347 (N_4347,N_3921,N_3007);
nand U4348 (N_4348,N_3439,N_3095);
nand U4349 (N_4349,N_3435,N_3201);
xor U4350 (N_4350,N_3336,N_3281);
nor U4351 (N_4351,N_3549,N_3765);
or U4352 (N_4352,N_3826,N_3813);
nand U4353 (N_4353,N_3331,N_3157);
or U4354 (N_4354,N_3618,N_3609);
nand U4355 (N_4355,N_3672,N_3816);
nor U4356 (N_4356,N_3190,N_3486);
and U4357 (N_4357,N_3739,N_3334);
nand U4358 (N_4358,N_3656,N_3470);
or U4359 (N_4359,N_3836,N_3870);
and U4360 (N_4360,N_3062,N_3297);
nor U4361 (N_4361,N_3140,N_3957);
nor U4362 (N_4362,N_3893,N_3624);
nand U4363 (N_4363,N_3406,N_3551);
nand U4364 (N_4364,N_3555,N_3019);
or U4365 (N_4365,N_3437,N_3289);
nand U4366 (N_4366,N_3284,N_3269);
nand U4367 (N_4367,N_3952,N_3631);
and U4368 (N_4368,N_3690,N_3230);
xnor U4369 (N_4369,N_3684,N_3238);
nor U4370 (N_4370,N_3841,N_3630);
or U4371 (N_4371,N_3954,N_3973);
xor U4372 (N_4372,N_3049,N_3171);
nor U4373 (N_4373,N_3809,N_3176);
nand U4374 (N_4374,N_3508,N_3120);
and U4375 (N_4375,N_3085,N_3910);
and U4376 (N_4376,N_3586,N_3304);
nand U4377 (N_4377,N_3707,N_3992);
nor U4378 (N_4378,N_3831,N_3958);
nor U4379 (N_4379,N_3451,N_3016);
xnor U4380 (N_4380,N_3725,N_3064);
or U4381 (N_4381,N_3788,N_3494);
nand U4382 (N_4382,N_3764,N_3337);
nor U4383 (N_4383,N_3458,N_3920);
or U4384 (N_4384,N_3429,N_3262);
xnor U4385 (N_4385,N_3990,N_3721);
nor U4386 (N_4386,N_3299,N_3368);
and U4387 (N_4387,N_3558,N_3706);
and U4388 (N_4388,N_3375,N_3796);
nand U4389 (N_4389,N_3073,N_3258);
nor U4390 (N_4390,N_3044,N_3147);
nor U4391 (N_4391,N_3614,N_3328);
nand U4392 (N_4392,N_3231,N_3495);
or U4393 (N_4393,N_3059,N_3136);
or U4394 (N_4394,N_3425,N_3110);
xnor U4395 (N_4395,N_3340,N_3003);
and U4396 (N_4396,N_3115,N_3768);
nand U4397 (N_4397,N_3882,N_3963);
or U4398 (N_4398,N_3911,N_3396);
and U4399 (N_4399,N_3143,N_3498);
xor U4400 (N_4400,N_3953,N_3480);
nor U4401 (N_4401,N_3540,N_3511);
nor U4402 (N_4402,N_3922,N_3192);
nand U4403 (N_4403,N_3700,N_3798);
xor U4404 (N_4404,N_3326,N_3078);
nor U4405 (N_4405,N_3311,N_3667);
and U4406 (N_4406,N_3858,N_3175);
nor U4407 (N_4407,N_3323,N_3135);
or U4408 (N_4408,N_3274,N_3483);
and U4409 (N_4409,N_3909,N_3626);
xor U4410 (N_4410,N_3679,N_3655);
xnor U4411 (N_4411,N_3357,N_3873);
or U4412 (N_4412,N_3945,N_3446);
or U4413 (N_4413,N_3597,N_3896);
xnor U4414 (N_4414,N_3692,N_3964);
or U4415 (N_4415,N_3860,N_3596);
xnor U4416 (N_4416,N_3689,N_3459);
nand U4417 (N_4417,N_3447,N_3293);
and U4418 (N_4418,N_3579,N_3960);
xor U4419 (N_4419,N_3461,N_3681);
or U4420 (N_4420,N_3247,N_3111);
and U4421 (N_4421,N_3779,N_3114);
or U4422 (N_4422,N_3118,N_3303);
nand U4423 (N_4423,N_3713,N_3823);
or U4424 (N_4424,N_3197,N_3463);
xnor U4425 (N_4425,N_3717,N_3492);
xor U4426 (N_4426,N_3333,N_3504);
and U4427 (N_4427,N_3916,N_3155);
nand U4428 (N_4428,N_3643,N_3904);
nand U4429 (N_4429,N_3594,N_3394);
nand U4430 (N_4430,N_3756,N_3730);
or U4431 (N_4431,N_3053,N_3318);
nand U4432 (N_4432,N_3828,N_3532);
nor U4433 (N_4433,N_3100,N_3172);
or U4434 (N_4434,N_3374,N_3634);
and U4435 (N_4435,N_3383,N_3046);
or U4436 (N_4436,N_3771,N_3226);
nand U4437 (N_4437,N_3589,N_3455);
xnor U4438 (N_4438,N_3026,N_3180);
or U4439 (N_4439,N_3528,N_3714);
nor U4440 (N_4440,N_3574,N_3438);
or U4441 (N_4441,N_3777,N_3748);
and U4442 (N_4442,N_3923,N_3490);
nand U4443 (N_4443,N_3881,N_3915);
or U4444 (N_4444,N_3466,N_3804);
nor U4445 (N_4445,N_3738,N_3273);
nand U4446 (N_4446,N_3462,N_3020);
or U4447 (N_4447,N_3359,N_3404);
or U4448 (N_4448,N_3081,N_3524);
xor U4449 (N_4449,N_3341,N_3473);
nor U4450 (N_4450,N_3991,N_3051);
nand U4451 (N_4451,N_3726,N_3621);
nor U4452 (N_4452,N_3633,N_3346);
nand U4453 (N_4453,N_3741,N_3031);
nor U4454 (N_4454,N_3871,N_3160);
and U4455 (N_4455,N_3556,N_3203);
or U4456 (N_4456,N_3209,N_3014);
nand U4457 (N_4457,N_3370,N_3525);
nor U4458 (N_4458,N_3984,N_3797);
and U4459 (N_4459,N_3456,N_3106);
xor U4460 (N_4460,N_3137,N_3665);
nor U4461 (N_4461,N_3940,N_3109);
and U4462 (N_4462,N_3890,N_3154);
and U4463 (N_4463,N_3243,N_3030);
nor U4464 (N_4464,N_3526,N_3693);
or U4465 (N_4465,N_3039,N_3522);
xnor U4466 (N_4466,N_3270,N_3642);
xor U4467 (N_4467,N_3207,N_3224);
nand U4468 (N_4468,N_3460,N_3103);
and U4469 (N_4469,N_3162,N_3086);
or U4470 (N_4470,N_3220,N_3697);
or U4471 (N_4471,N_3414,N_3056);
nor U4472 (N_4472,N_3856,N_3892);
xor U4473 (N_4473,N_3107,N_3096);
xnor U4474 (N_4474,N_3583,N_3479);
xor U4475 (N_4475,N_3835,N_3944);
and U4476 (N_4476,N_3936,N_3401);
and U4477 (N_4477,N_3886,N_3332);
or U4478 (N_4478,N_3650,N_3237);
and U4479 (N_4479,N_3815,N_3347);
and U4480 (N_4480,N_3617,N_3027);
nand U4481 (N_4481,N_3750,N_3786);
xor U4482 (N_4482,N_3063,N_3363);
nand U4483 (N_4483,N_3889,N_3949);
or U4484 (N_4484,N_3112,N_3185);
nand U4485 (N_4485,N_3720,N_3235);
or U4486 (N_4486,N_3474,N_3276);
and U4487 (N_4487,N_3471,N_3753);
nor U4488 (N_4488,N_3547,N_3907);
xor U4489 (N_4489,N_3187,N_3075);
xor U4490 (N_4490,N_3251,N_3639);
nand U4491 (N_4491,N_3833,N_3855);
xor U4492 (N_4492,N_3327,N_3578);
xor U4493 (N_4493,N_3216,N_3736);
nand U4494 (N_4494,N_3746,N_3862);
nand U4495 (N_4495,N_3670,N_3133);
nand U4496 (N_4496,N_3042,N_3153);
or U4497 (N_4497,N_3568,N_3469);
xnor U4498 (N_4498,N_3834,N_3839);
or U4499 (N_4499,N_3300,N_3440);
nand U4500 (N_4500,N_3490,N_3739);
nand U4501 (N_4501,N_3574,N_3777);
nor U4502 (N_4502,N_3623,N_3441);
or U4503 (N_4503,N_3292,N_3906);
or U4504 (N_4504,N_3781,N_3721);
nor U4505 (N_4505,N_3315,N_3235);
xnor U4506 (N_4506,N_3841,N_3439);
nor U4507 (N_4507,N_3456,N_3572);
nand U4508 (N_4508,N_3400,N_3838);
xnor U4509 (N_4509,N_3975,N_3669);
and U4510 (N_4510,N_3506,N_3343);
and U4511 (N_4511,N_3578,N_3910);
or U4512 (N_4512,N_3761,N_3262);
or U4513 (N_4513,N_3353,N_3338);
and U4514 (N_4514,N_3617,N_3959);
and U4515 (N_4515,N_3155,N_3531);
nor U4516 (N_4516,N_3912,N_3550);
nor U4517 (N_4517,N_3700,N_3420);
or U4518 (N_4518,N_3751,N_3247);
nand U4519 (N_4519,N_3101,N_3875);
and U4520 (N_4520,N_3345,N_3358);
nor U4521 (N_4521,N_3160,N_3319);
or U4522 (N_4522,N_3805,N_3049);
nor U4523 (N_4523,N_3860,N_3072);
xor U4524 (N_4524,N_3764,N_3030);
xor U4525 (N_4525,N_3494,N_3932);
and U4526 (N_4526,N_3308,N_3395);
and U4527 (N_4527,N_3981,N_3920);
nor U4528 (N_4528,N_3757,N_3345);
nor U4529 (N_4529,N_3734,N_3223);
nor U4530 (N_4530,N_3999,N_3111);
or U4531 (N_4531,N_3436,N_3063);
nand U4532 (N_4532,N_3918,N_3841);
nor U4533 (N_4533,N_3149,N_3282);
nor U4534 (N_4534,N_3574,N_3274);
nand U4535 (N_4535,N_3212,N_3668);
and U4536 (N_4536,N_3792,N_3507);
xor U4537 (N_4537,N_3746,N_3072);
nand U4538 (N_4538,N_3677,N_3251);
xnor U4539 (N_4539,N_3173,N_3107);
nand U4540 (N_4540,N_3365,N_3896);
nor U4541 (N_4541,N_3539,N_3892);
nand U4542 (N_4542,N_3763,N_3577);
xor U4543 (N_4543,N_3347,N_3768);
or U4544 (N_4544,N_3919,N_3681);
nand U4545 (N_4545,N_3281,N_3068);
or U4546 (N_4546,N_3912,N_3203);
nand U4547 (N_4547,N_3651,N_3169);
nor U4548 (N_4548,N_3827,N_3704);
and U4549 (N_4549,N_3675,N_3041);
nor U4550 (N_4550,N_3658,N_3840);
nand U4551 (N_4551,N_3244,N_3139);
xor U4552 (N_4552,N_3121,N_3403);
nand U4553 (N_4553,N_3993,N_3271);
and U4554 (N_4554,N_3420,N_3172);
xor U4555 (N_4555,N_3478,N_3651);
and U4556 (N_4556,N_3813,N_3245);
nor U4557 (N_4557,N_3685,N_3378);
and U4558 (N_4558,N_3282,N_3921);
and U4559 (N_4559,N_3093,N_3237);
nor U4560 (N_4560,N_3263,N_3529);
xnor U4561 (N_4561,N_3560,N_3859);
nor U4562 (N_4562,N_3150,N_3179);
xnor U4563 (N_4563,N_3468,N_3782);
nand U4564 (N_4564,N_3065,N_3279);
nor U4565 (N_4565,N_3089,N_3509);
nor U4566 (N_4566,N_3790,N_3593);
or U4567 (N_4567,N_3223,N_3466);
nor U4568 (N_4568,N_3904,N_3751);
nand U4569 (N_4569,N_3824,N_3549);
or U4570 (N_4570,N_3080,N_3373);
nand U4571 (N_4571,N_3435,N_3552);
xor U4572 (N_4572,N_3646,N_3715);
or U4573 (N_4573,N_3785,N_3457);
nor U4574 (N_4574,N_3645,N_3419);
or U4575 (N_4575,N_3579,N_3496);
nor U4576 (N_4576,N_3543,N_3718);
nand U4577 (N_4577,N_3392,N_3124);
nand U4578 (N_4578,N_3748,N_3594);
nor U4579 (N_4579,N_3716,N_3571);
and U4580 (N_4580,N_3739,N_3636);
and U4581 (N_4581,N_3589,N_3820);
xnor U4582 (N_4582,N_3645,N_3293);
or U4583 (N_4583,N_3336,N_3088);
nand U4584 (N_4584,N_3975,N_3526);
nand U4585 (N_4585,N_3152,N_3966);
xnor U4586 (N_4586,N_3219,N_3242);
or U4587 (N_4587,N_3007,N_3091);
nand U4588 (N_4588,N_3914,N_3484);
xnor U4589 (N_4589,N_3179,N_3760);
nand U4590 (N_4590,N_3820,N_3863);
nor U4591 (N_4591,N_3783,N_3363);
nand U4592 (N_4592,N_3326,N_3958);
or U4593 (N_4593,N_3555,N_3769);
or U4594 (N_4594,N_3273,N_3854);
and U4595 (N_4595,N_3202,N_3003);
nand U4596 (N_4596,N_3661,N_3713);
or U4597 (N_4597,N_3338,N_3743);
and U4598 (N_4598,N_3351,N_3867);
nor U4599 (N_4599,N_3946,N_3532);
nand U4600 (N_4600,N_3472,N_3405);
xnor U4601 (N_4601,N_3614,N_3247);
nor U4602 (N_4602,N_3021,N_3550);
nand U4603 (N_4603,N_3118,N_3997);
nand U4604 (N_4604,N_3798,N_3925);
or U4605 (N_4605,N_3566,N_3751);
nor U4606 (N_4606,N_3972,N_3483);
xor U4607 (N_4607,N_3162,N_3071);
xnor U4608 (N_4608,N_3284,N_3407);
or U4609 (N_4609,N_3042,N_3966);
or U4610 (N_4610,N_3097,N_3015);
nand U4611 (N_4611,N_3053,N_3010);
and U4612 (N_4612,N_3284,N_3746);
xnor U4613 (N_4613,N_3953,N_3108);
or U4614 (N_4614,N_3806,N_3567);
xor U4615 (N_4615,N_3469,N_3187);
or U4616 (N_4616,N_3245,N_3486);
nand U4617 (N_4617,N_3913,N_3628);
nor U4618 (N_4618,N_3981,N_3707);
xnor U4619 (N_4619,N_3997,N_3648);
or U4620 (N_4620,N_3854,N_3582);
xor U4621 (N_4621,N_3279,N_3665);
nand U4622 (N_4622,N_3068,N_3875);
nand U4623 (N_4623,N_3814,N_3908);
xor U4624 (N_4624,N_3727,N_3274);
xnor U4625 (N_4625,N_3408,N_3739);
or U4626 (N_4626,N_3869,N_3551);
nand U4627 (N_4627,N_3960,N_3820);
nor U4628 (N_4628,N_3277,N_3824);
or U4629 (N_4629,N_3829,N_3663);
or U4630 (N_4630,N_3017,N_3145);
xnor U4631 (N_4631,N_3158,N_3418);
or U4632 (N_4632,N_3486,N_3968);
nand U4633 (N_4633,N_3670,N_3188);
or U4634 (N_4634,N_3500,N_3624);
xnor U4635 (N_4635,N_3212,N_3079);
nand U4636 (N_4636,N_3934,N_3544);
and U4637 (N_4637,N_3621,N_3163);
xnor U4638 (N_4638,N_3195,N_3065);
and U4639 (N_4639,N_3651,N_3684);
and U4640 (N_4640,N_3009,N_3397);
nor U4641 (N_4641,N_3652,N_3498);
nand U4642 (N_4642,N_3094,N_3228);
and U4643 (N_4643,N_3031,N_3881);
nor U4644 (N_4644,N_3832,N_3298);
nand U4645 (N_4645,N_3266,N_3791);
and U4646 (N_4646,N_3659,N_3209);
or U4647 (N_4647,N_3359,N_3847);
nand U4648 (N_4648,N_3157,N_3547);
and U4649 (N_4649,N_3556,N_3694);
and U4650 (N_4650,N_3838,N_3765);
nor U4651 (N_4651,N_3514,N_3795);
or U4652 (N_4652,N_3591,N_3555);
nand U4653 (N_4653,N_3134,N_3930);
nand U4654 (N_4654,N_3131,N_3492);
xnor U4655 (N_4655,N_3728,N_3575);
nand U4656 (N_4656,N_3279,N_3510);
or U4657 (N_4657,N_3755,N_3965);
or U4658 (N_4658,N_3832,N_3023);
and U4659 (N_4659,N_3653,N_3718);
xor U4660 (N_4660,N_3173,N_3816);
or U4661 (N_4661,N_3587,N_3883);
or U4662 (N_4662,N_3871,N_3294);
or U4663 (N_4663,N_3822,N_3024);
and U4664 (N_4664,N_3834,N_3499);
xnor U4665 (N_4665,N_3291,N_3869);
or U4666 (N_4666,N_3087,N_3277);
nor U4667 (N_4667,N_3683,N_3334);
and U4668 (N_4668,N_3044,N_3686);
and U4669 (N_4669,N_3553,N_3917);
and U4670 (N_4670,N_3688,N_3285);
xnor U4671 (N_4671,N_3812,N_3517);
or U4672 (N_4672,N_3529,N_3687);
nor U4673 (N_4673,N_3929,N_3573);
xnor U4674 (N_4674,N_3864,N_3512);
nor U4675 (N_4675,N_3526,N_3213);
nand U4676 (N_4676,N_3161,N_3787);
nor U4677 (N_4677,N_3001,N_3437);
or U4678 (N_4678,N_3503,N_3035);
xnor U4679 (N_4679,N_3590,N_3777);
and U4680 (N_4680,N_3526,N_3527);
nand U4681 (N_4681,N_3517,N_3684);
nand U4682 (N_4682,N_3463,N_3362);
nor U4683 (N_4683,N_3142,N_3102);
and U4684 (N_4684,N_3329,N_3942);
xor U4685 (N_4685,N_3061,N_3793);
nand U4686 (N_4686,N_3413,N_3982);
and U4687 (N_4687,N_3764,N_3514);
and U4688 (N_4688,N_3179,N_3390);
or U4689 (N_4689,N_3238,N_3530);
or U4690 (N_4690,N_3852,N_3052);
nor U4691 (N_4691,N_3245,N_3270);
or U4692 (N_4692,N_3237,N_3585);
xor U4693 (N_4693,N_3535,N_3507);
xor U4694 (N_4694,N_3301,N_3911);
or U4695 (N_4695,N_3293,N_3590);
nand U4696 (N_4696,N_3989,N_3152);
or U4697 (N_4697,N_3459,N_3755);
or U4698 (N_4698,N_3592,N_3482);
or U4699 (N_4699,N_3478,N_3047);
or U4700 (N_4700,N_3110,N_3391);
or U4701 (N_4701,N_3578,N_3463);
nor U4702 (N_4702,N_3385,N_3332);
or U4703 (N_4703,N_3127,N_3234);
nor U4704 (N_4704,N_3862,N_3392);
xnor U4705 (N_4705,N_3577,N_3547);
nand U4706 (N_4706,N_3654,N_3169);
and U4707 (N_4707,N_3282,N_3689);
or U4708 (N_4708,N_3725,N_3001);
and U4709 (N_4709,N_3918,N_3738);
or U4710 (N_4710,N_3673,N_3857);
nor U4711 (N_4711,N_3576,N_3551);
xnor U4712 (N_4712,N_3773,N_3878);
and U4713 (N_4713,N_3584,N_3002);
nand U4714 (N_4714,N_3068,N_3822);
nand U4715 (N_4715,N_3501,N_3290);
and U4716 (N_4716,N_3301,N_3368);
nand U4717 (N_4717,N_3901,N_3164);
or U4718 (N_4718,N_3251,N_3987);
nor U4719 (N_4719,N_3026,N_3781);
xnor U4720 (N_4720,N_3882,N_3465);
nand U4721 (N_4721,N_3037,N_3849);
and U4722 (N_4722,N_3756,N_3115);
nor U4723 (N_4723,N_3634,N_3925);
or U4724 (N_4724,N_3516,N_3438);
nor U4725 (N_4725,N_3276,N_3179);
and U4726 (N_4726,N_3303,N_3588);
and U4727 (N_4727,N_3347,N_3575);
and U4728 (N_4728,N_3565,N_3460);
nor U4729 (N_4729,N_3369,N_3967);
and U4730 (N_4730,N_3349,N_3312);
and U4731 (N_4731,N_3243,N_3838);
nor U4732 (N_4732,N_3100,N_3964);
nor U4733 (N_4733,N_3614,N_3274);
xnor U4734 (N_4734,N_3260,N_3241);
nor U4735 (N_4735,N_3495,N_3880);
nand U4736 (N_4736,N_3122,N_3553);
or U4737 (N_4737,N_3325,N_3829);
xor U4738 (N_4738,N_3401,N_3667);
nor U4739 (N_4739,N_3807,N_3573);
nor U4740 (N_4740,N_3353,N_3715);
nor U4741 (N_4741,N_3206,N_3979);
nor U4742 (N_4742,N_3239,N_3540);
nand U4743 (N_4743,N_3255,N_3127);
and U4744 (N_4744,N_3665,N_3228);
or U4745 (N_4745,N_3804,N_3644);
nor U4746 (N_4746,N_3038,N_3836);
and U4747 (N_4747,N_3242,N_3170);
xor U4748 (N_4748,N_3863,N_3077);
nor U4749 (N_4749,N_3656,N_3126);
and U4750 (N_4750,N_3501,N_3593);
and U4751 (N_4751,N_3365,N_3685);
and U4752 (N_4752,N_3494,N_3135);
and U4753 (N_4753,N_3611,N_3082);
and U4754 (N_4754,N_3619,N_3820);
nor U4755 (N_4755,N_3070,N_3134);
nor U4756 (N_4756,N_3575,N_3277);
and U4757 (N_4757,N_3227,N_3482);
nand U4758 (N_4758,N_3966,N_3427);
nor U4759 (N_4759,N_3534,N_3672);
or U4760 (N_4760,N_3811,N_3103);
nor U4761 (N_4761,N_3037,N_3636);
or U4762 (N_4762,N_3772,N_3710);
nand U4763 (N_4763,N_3387,N_3794);
and U4764 (N_4764,N_3495,N_3029);
nor U4765 (N_4765,N_3513,N_3168);
nand U4766 (N_4766,N_3295,N_3345);
and U4767 (N_4767,N_3412,N_3776);
or U4768 (N_4768,N_3475,N_3382);
and U4769 (N_4769,N_3598,N_3814);
nand U4770 (N_4770,N_3774,N_3671);
and U4771 (N_4771,N_3357,N_3908);
nor U4772 (N_4772,N_3223,N_3178);
nor U4773 (N_4773,N_3934,N_3836);
nand U4774 (N_4774,N_3014,N_3874);
xnor U4775 (N_4775,N_3922,N_3861);
nand U4776 (N_4776,N_3842,N_3189);
and U4777 (N_4777,N_3496,N_3946);
and U4778 (N_4778,N_3349,N_3204);
or U4779 (N_4779,N_3425,N_3397);
nand U4780 (N_4780,N_3403,N_3778);
nand U4781 (N_4781,N_3310,N_3881);
nand U4782 (N_4782,N_3110,N_3271);
nand U4783 (N_4783,N_3485,N_3717);
or U4784 (N_4784,N_3246,N_3582);
xor U4785 (N_4785,N_3710,N_3495);
xnor U4786 (N_4786,N_3921,N_3456);
or U4787 (N_4787,N_3330,N_3273);
or U4788 (N_4788,N_3939,N_3853);
or U4789 (N_4789,N_3558,N_3784);
xor U4790 (N_4790,N_3838,N_3784);
nor U4791 (N_4791,N_3258,N_3886);
xor U4792 (N_4792,N_3565,N_3693);
and U4793 (N_4793,N_3650,N_3813);
and U4794 (N_4794,N_3243,N_3439);
nor U4795 (N_4795,N_3331,N_3449);
xnor U4796 (N_4796,N_3761,N_3620);
nand U4797 (N_4797,N_3245,N_3083);
xor U4798 (N_4798,N_3779,N_3982);
nand U4799 (N_4799,N_3281,N_3182);
or U4800 (N_4800,N_3563,N_3641);
or U4801 (N_4801,N_3192,N_3350);
nand U4802 (N_4802,N_3887,N_3785);
or U4803 (N_4803,N_3720,N_3400);
nor U4804 (N_4804,N_3872,N_3902);
xor U4805 (N_4805,N_3626,N_3911);
and U4806 (N_4806,N_3617,N_3921);
nand U4807 (N_4807,N_3637,N_3450);
or U4808 (N_4808,N_3492,N_3428);
and U4809 (N_4809,N_3351,N_3352);
and U4810 (N_4810,N_3662,N_3382);
or U4811 (N_4811,N_3610,N_3218);
nor U4812 (N_4812,N_3107,N_3574);
xor U4813 (N_4813,N_3740,N_3245);
nor U4814 (N_4814,N_3478,N_3051);
or U4815 (N_4815,N_3552,N_3100);
nand U4816 (N_4816,N_3752,N_3264);
or U4817 (N_4817,N_3529,N_3993);
nor U4818 (N_4818,N_3331,N_3054);
or U4819 (N_4819,N_3084,N_3746);
nand U4820 (N_4820,N_3836,N_3666);
nand U4821 (N_4821,N_3709,N_3905);
xnor U4822 (N_4822,N_3617,N_3233);
or U4823 (N_4823,N_3401,N_3049);
nand U4824 (N_4824,N_3220,N_3322);
nand U4825 (N_4825,N_3812,N_3473);
and U4826 (N_4826,N_3862,N_3261);
nand U4827 (N_4827,N_3238,N_3526);
nand U4828 (N_4828,N_3756,N_3074);
nor U4829 (N_4829,N_3246,N_3625);
or U4830 (N_4830,N_3910,N_3603);
or U4831 (N_4831,N_3863,N_3456);
xnor U4832 (N_4832,N_3291,N_3917);
or U4833 (N_4833,N_3344,N_3286);
or U4834 (N_4834,N_3464,N_3092);
nand U4835 (N_4835,N_3345,N_3689);
nor U4836 (N_4836,N_3045,N_3789);
nand U4837 (N_4837,N_3073,N_3225);
nand U4838 (N_4838,N_3478,N_3807);
nand U4839 (N_4839,N_3364,N_3236);
and U4840 (N_4840,N_3679,N_3925);
or U4841 (N_4841,N_3117,N_3137);
or U4842 (N_4842,N_3139,N_3256);
nand U4843 (N_4843,N_3332,N_3612);
nor U4844 (N_4844,N_3044,N_3111);
xnor U4845 (N_4845,N_3459,N_3051);
nor U4846 (N_4846,N_3893,N_3702);
nand U4847 (N_4847,N_3593,N_3484);
and U4848 (N_4848,N_3644,N_3005);
nand U4849 (N_4849,N_3738,N_3441);
nor U4850 (N_4850,N_3060,N_3179);
nand U4851 (N_4851,N_3516,N_3330);
xor U4852 (N_4852,N_3739,N_3634);
nand U4853 (N_4853,N_3198,N_3001);
nand U4854 (N_4854,N_3464,N_3381);
xnor U4855 (N_4855,N_3620,N_3287);
nor U4856 (N_4856,N_3141,N_3082);
and U4857 (N_4857,N_3701,N_3522);
nand U4858 (N_4858,N_3030,N_3598);
nand U4859 (N_4859,N_3178,N_3158);
xnor U4860 (N_4860,N_3533,N_3017);
and U4861 (N_4861,N_3088,N_3439);
xor U4862 (N_4862,N_3079,N_3056);
xor U4863 (N_4863,N_3905,N_3630);
nor U4864 (N_4864,N_3794,N_3067);
xor U4865 (N_4865,N_3452,N_3995);
nor U4866 (N_4866,N_3638,N_3041);
nor U4867 (N_4867,N_3382,N_3355);
nand U4868 (N_4868,N_3373,N_3542);
and U4869 (N_4869,N_3537,N_3500);
xor U4870 (N_4870,N_3820,N_3729);
nand U4871 (N_4871,N_3434,N_3328);
nor U4872 (N_4872,N_3992,N_3576);
xnor U4873 (N_4873,N_3303,N_3878);
nand U4874 (N_4874,N_3321,N_3062);
nor U4875 (N_4875,N_3959,N_3589);
and U4876 (N_4876,N_3849,N_3650);
and U4877 (N_4877,N_3167,N_3595);
nor U4878 (N_4878,N_3924,N_3629);
xnor U4879 (N_4879,N_3726,N_3821);
nand U4880 (N_4880,N_3863,N_3970);
nor U4881 (N_4881,N_3774,N_3979);
nand U4882 (N_4882,N_3108,N_3252);
nor U4883 (N_4883,N_3671,N_3273);
nor U4884 (N_4884,N_3718,N_3079);
xor U4885 (N_4885,N_3677,N_3347);
xnor U4886 (N_4886,N_3729,N_3066);
or U4887 (N_4887,N_3630,N_3944);
and U4888 (N_4888,N_3740,N_3481);
or U4889 (N_4889,N_3382,N_3455);
nor U4890 (N_4890,N_3718,N_3010);
nand U4891 (N_4891,N_3095,N_3999);
nand U4892 (N_4892,N_3473,N_3620);
or U4893 (N_4893,N_3839,N_3439);
nor U4894 (N_4894,N_3059,N_3475);
xnor U4895 (N_4895,N_3712,N_3314);
nor U4896 (N_4896,N_3949,N_3277);
and U4897 (N_4897,N_3355,N_3075);
nand U4898 (N_4898,N_3125,N_3952);
and U4899 (N_4899,N_3670,N_3499);
xor U4900 (N_4900,N_3260,N_3125);
nand U4901 (N_4901,N_3357,N_3638);
xnor U4902 (N_4902,N_3298,N_3469);
and U4903 (N_4903,N_3006,N_3994);
and U4904 (N_4904,N_3895,N_3679);
nor U4905 (N_4905,N_3062,N_3764);
nor U4906 (N_4906,N_3362,N_3581);
or U4907 (N_4907,N_3752,N_3642);
or U4908 (N_4908,N_3008,N_3852);
or U4909 (N_4909,N_3129,N_3683);
and U4910 (N_4910,N_3961,N_3918);
nand U4911 (N_4911,N_3843,N_3021);
or U4912 (N_4912,N_3719,N_3784);
and U4913 (N_4913,N_3188,N_3425);
and U4914 (N_4914,N_3129,N_3739);
and U4915 (N_4915,N_3833,N_3222);
and U4916 (N_4916,N_3354,N_3790);
nand U4917 (N_4917,N_3497,N_3332);
or U4918 (N_4918,N_3364,N_3035);
or U4919 (N_4919,N_3180,N_3416);
nand U4920 (N_4920,N_3691,N_3182);
and U4921 (N_4921,N_3601,N_3201);
nor U4922 (N_4922,N_3707,N_3300);
and U4923 (N_4923,N_3457,N_3055);
xor U4924 (N_4924,N_3702,N_3597);
or U4925 (N_4925,N_3739,N_3175);
nand U4926 (N_4926,N_3485,N_3068);
xnor U4927 (N_4927,N_3034,N_3706);
nor U4928 (N_4928,N_3973,N_3767);
and U4929 (N_4929,N_3601,N_3481);
nor U4930 (N_4930,N_3628,N_3388);
xnor U4931 (N_4931,N_3865,N_3956);
or U4932 (N_4932,N_3768,N_3032);
and U4933 (N_4933,N_3034,N_3262);
nand U4934 (N_4934,N_3465,N_3129);
xnor U4935 (N_4935,N_3795,N_3298);
and U4936 (N_4936,N_3735,N_3267);
nor U4937 (N_4937,N_3347,N_3192);
nor U4938 (N_4938,N_3073,N_3108);
nor U4939 (N_4939,N_3167,N_3221);
nor U4940 (N_4940,N_3019,N_3333);
nor U4941 (N_4941,N_3289,N_3619);
and U4942 (N_4942,N_3147,N_3957);
and U4943 (N_4943,N_3212,N_3406);
and U4944 (N_4944,N_3166,N_3718);
or U4945 (N_4945,N_3789,N_3765);
xor U4946 (N_4946,N_3301,N_3513);
xnor U4947 (N_4947,N_3546,N_3110);
and U4948 (N_4948,N_3889,N_3162);
and U4949 (N_4949,N_3833,N_3414);
and U4950 (N_4950,N_3899,N_3576);
and U4951 (N_4951,N_3671,N_3203);
xor U4952 (N_4952,N_3742,N_3246);
and U4953 (N_4953,N_3781,N_3242);
nor U4954 (N_4954,N_3015,N_3276);
and U4955 (N_4955,N_3981,N_3178);
and U4956 (N_4956,N_3588,N_3543);
nand U4957 (N_4957,N_3277,N_3000);
or U4958 (N_4958,N_3508,N_3849);
or U4959 (N_4959,N_3573,N_3074);
or U4960 (N_4960,N_3667,N_3031);
nor U4961 (N_4961,N_3311,N_3162);
and U4962 (N_4962,N_3588,N_3694);
or U4963 (N_4963,N_3148,N_3484);
nand U4964 (N_4964,N_3055,N_3417);
or U4965 (N_4965,N_3300,N_3546);
xnor U4966 (N_4966,N_3591,N_3463);
nor U4967 (N_4967,N_3457,N_3270);
or U4968 (N_4968,N_3612,N_3085);
xnor U4969 (N_4969,N_3175,N_3539);
xor U4970 (N_4970,N_3140,N_3706);
xor U4971 (N_4971,N_3095,N_3897);
nand U4972 (N_4972,N_3343,N_3367);
nor U4973 (N_4973,N_3630,N_3258);
or U4974 (N_4974,N_3090,N_3159);
and U4975 (N_4975,N_3672,N_3968);
xor U4976 (N_4976,N_3714,N_3935);
nor U4977 (N_4977,N_3632,N_3719);
nand U4978 (N_4978,N_3506,N_3709);
nor U4979 (N_4979,N_3251,N_3112);
xnor U4980 (N_4980,N_3525,N_3457);
xnor U4981 (N_4981,N_3035,N_3012);
nor U4982 (N_4982,N_3535,N_3832);
and U4983 (N_4983,N_3675,N_3369);
and U4984 (N_4984,N_3270,N_3359);
or U4985 (N_4985,N_3636,N_3101);
or U4986 (N_4986,N_3997,N_3002);
and U4987 (N_4987,N_3888,N_3578);
nand U4988 (N_4988,N_3569,N_3410);
or U4989 (N_4989,N_3188,N_3295);
nand U4990 (N_4990,N_3793,N_3314);
xor U4991 (N_4991,N_3814,N_3168);
nand U4992 (N_4992,N_3027,N_3202);
nand U4993 (N_4993,N_3182,N_3214);
or U4994 (N_4994,N_3487,N_3199);
and U4995 (N_4995,N_3760,N_3849);
or U4996 (N_4996,N_3914,N_3514);
nor U4997 (N_4997,N_3661,N_3243);
and U4998 (N_4998,N_3339,N_3719);
nor U4999 (N_4999,N_3778,N_3359);
nand U5000 (N_5000,N_4040,N_4150);
nand U5001 (N_5001,N_4919,N_4543);
and U5002 (N_5002,N_4342,N_4743);
nand U5003 (N_5003,N_4384,N_4748);
xnor U5004 (N_5004,N_4464,N_4922);
nand U5005 (N_5005,N_4727,N_4959);
and U5006 (N_5006,N_4846,N_4976);
xor U5007 (N_5007,N_4447,N_4954);
or U5008 (N_5008,N_4062,N_4492);
nand U5009 (N_5009,N_4803,N_4430);
nand U5010 (N_5010,N_4100,N_4310);
xnor U5011 (N_5011,N_4847,N_4592);
and U5012 (N_5012,N_4224,N_4608);
and U5013 (N_5013,N_4419,N_4963);
or U5014 (N_5014,N_4518,N_4788);
and U5015 (N_5015,N_4547,N_4532);
nand U5016 (N_5016,N_4501,N_4413);
and U5017 (N_5017,N_4321,N_4577);
and U5018 (N_5018,N_4170,N_4314);
or U5019 (N_5019,N_4990,N_4636);
and U5020 (N_5020,N_4266,N_4587);
nor U5021 (N_5021,N_4367,N_4439);
and U5022 (N_5022,N_4039,N_4763);
nor U5023 (N_5023,N_4120,N_4907);
xor U5024 (N_5024,N_4979,N_4397);
or U5025 (N_5025,N_4682,N_4565);
and U5026 (N_5026,N_4362,N_4662);
or U5027 (N_5027,N_4685,N_4752);
or U5028 (N_5028,N_4920,N_4791);
or U5029 (N_5029,N_4630,N_4677);
or U5030 (N_5030,N_4722,N_4036);
nand U5031 (N_5031,N_4940,N_4533);
and U5032 (N_5032,N_4667,N_4134);
nor U5033 (N_5033,N_4719,N_4725);
and U5034 (N_5034,N_4228,N_4023);
or U5035 (N_5035,N_4034,N_4481);
nand U5036 (N_5036,N_4307,N_4506);
or U5037 (N_5037,N_4472,N_4042);
and U5038 (N_5038,N_4640,N_4840);
xor U5039 (N_5039,N_4179,N_4790);
and U5040 (N_5040,N_4552,N_4912);
or U5041 (N_5041,N_4969,N_4379);
nand U5042 (N_5042,N_4328,N_4096);
nand U5043 (N_5043,N_4766,N_4869);
and U5044 (N_5044,N_4054,N_4015);
nand U5045 (N_5045,N_4626,N_4204);
nor U5046 (N_5046,N_4888,N_4541);
nor U5047 (N_5047,N_4581,N_4002);
xnor U5048 (N_5048,N_4848,N_4388);
xnor U5049 (N_5049,N_4897,N_4390);
xnor U5050 (N_5050,N_4807,N_4122);
or U5051 (N_5051,N_4461,N_4595);
nor U5052 (N_5052,N_4793,N_4285);
xnor U5053 (N_5053,N_4065,N_4038);
nor U5054 (N_5054,N_4841,N_4730);
xor U5055 (N_5055,N_4649,N_4312);
nor U5056 (N_5056,N_4918,N_4851);
or U5057 (N_5057,N_4381,N_4945);
nor U5058 (N_5058,N_4875,N_4911);
and U5059 (N_5059,N_4905,N_4024);
nand U5060 (N_5060,N_4915,N_4811);
and U5061 (N_5061,N_4427,N_4988);
nand U5062 (N_5062,N_4396,N_4659);
and U5063 (N_5063,N_4200,N_4726);
xnor U5064 (N_5064,N_4966,N_4297);
and U5065 (N_5065,N_4782,N_4870);
nor U5066 (N_5066,N_4765,N_4816);
nand U5067 (N_5067,N_4434,N_4070);
or U5068 (N_5068,N_4099,N_4267);
xor U5069 (N_5069,N_4776,N_4638);
and U5070 (N_5070,N_4562,N_4681);
xor U5071 (N_5071,N_4044,N_4859);
nor U5072 (N_5072,N_4928,N_4814);
or U5073 (N_5073,N_4942,N_4639);
nand U5074 (N_5074,N_4000,N_4197);
and U5075 (N_5075,N_4061,N_4718);
nor U5076 (N_5076,N_4475,N_4889);
and U5077 (N_5077,N_4697,N_4670);
and U5078 (N_5078,N_4291,N_4346);
or U5079 (N_5079,N_4029,N_4713);
or U5080 (N_5080,N_4391,N_4850);
xnor U5081 (N_5081,N_4190,N_4611);
nand U5082 (N_5082,N_4056,N_4523);
or U5083 (N_5083,N_4927,N_4806);
nand U5084 (N_5084,N_4265,N_4799);
nand U5085 (N_5085,N_4019,N_4779);
and U5086 (N_5086,N_4570,N_4855);
nor U5087 (N_5087,N_4223,N_4978);
nand U5088 (N_5088,N_4967,N_4206);
and U5089 (N_5089,N_4690,N_4633);
xnor U5090 (N_5090,N_4074,N_4237);
nand U5091 (N_5091,N_4524,N_4904);
xor U5092 (N_5092,N_4892,N_4354);
and U5093 (N_5093,N_4734,N_4508);
nand U5094 (N_5094,N_4196,N_4613);
nor U5095 (N_5095,N_4130,N_4972);
and U5096 (N_5096,N_4385,N_4449);
or U5097 (N_5097,N_4553,N_4288);
or U5098 (N_5098,N_4446,N_4195);
nor U5099 (N_5099,N_4324,N_4064);
and U5100 (N_5100,N_4631,N_4091);
nor U5101 (N_5101,N_4025,N_4094);
nor U5102 (N_5102,N_4331,N_4490);
nor U5103 (N_5103,N_4171,N_4836);
nand U5104 (N_5104,N_4345,N_4079);
or U5105 (N_5105,N_4704,N_4637);
or U5106 (N_5106,N_4135,N_4746);
nor U5107 (N_5107,N_4699,N_4764);
and U5108 (N_5108,N_4383,N_4977);
nand U5109 (N_5109,N_4934,N_4035);
nor U5110 (N_5110,N_4401,N_4620);
and U5111 (N_5111,N_4937,N_4634);
xnor U5112 (N_5112,N_4377,N_4256);
xnor U5113 (N_5113,N_4526,N_4232);
or U5114 (N_5114,N_4466,N_4548);
nor U5115 (N_5115,N_4674,N_4672);
or U5116 (N_5116,N_4465,N_4833);
and U5117 (N_5117,N_4047,N_4772);
nand U5118 (N_5118,N_4077,N_4832);
nor U5119 (N_5119,N_4497,N_4045);
or U5120 (N_5120,N_4629,N_4879);
nor U5121 (N_5121,N_4917,N_4360);
nor U5122 (N_5122,N_4794,N_4320);
or U5123 (N_5123,N_4231,N_4758);
or U5124 (N_5124,N_4160,N_4365);
and U5125 (N_5125,N_4088,N_4111);
or U5126 (N_5126,N_4557,N_4169);
nor U5127 (N_5127,N_4805,N_4392);
and U5128 (N_5128,N_4189,N_4353);
xnor U5129 (N_5129,N_4612,N_4175);
nand U5130 (N_5130,N_4361,N_4106);
nor U5131 (N_5131,N_4031,N_4624);
nor U5132 (N_5132,N_4753,N_4487);
xor U5133 (N_5133,N_4780,N_4105);
nand U5134 (N_5134,N_4226,N_4368);
nand U5135 (N_5135,N_4380,N_4366);
xnor U5136 (N_5136,N_4123,N_4184);
xnor U5137 (N_5137,N_4375,N_4341);
or U5138 (N_5138,N_4452,N_4902);
xor U5139 (N_5139,N_4866,N_4738);
nand U5140 (N_5140,N_4510,N_4652);
nand U5141 (N_5141,N_4731,N_4117);
and U5142 (N_5142,N_4217,N_4474);
nor U5143 (N_5143,N_4589,N_4132);
xnor U5144 (N_5144,N_4207,N_4350);
xor U5145 (N_5145,N_4334,N_4315);
xor U5146 (N_5146,N_4948,N_4787);
and U5147 (N_5147,N_4899,N_4454);
nand U5148 (N_5148,N_4711,N_4133);
or U5149 (N_5149,N_4403,N_4268);
nand U5150 (N_5150,N_4568,N_4894);
xor U5151 (N_5151,N_4947,N_4839);
nand U5152 (N_5152,N_4322,N_4477);
nor U5153 (N_5153,N_4534,N_4095);
nor U5154 (N_5154,N_4571,N_4168);
nor U5155 (N_5155,N_4293,N_4614);
nor U5156 (N_5156,N_4673,N_4276);
nor U5157 (N_5157,N_4212,N_4826);
nor U5158 (N_5158,N_4149,N_4984);
or U5159 (N_5159,N_4248,N_4389);
xnor U5160 (N_5160,N_4574,N_4873);
and U5161 (N_5161,N_4273,N_4622);
or U5162 (N_5162,N_4828,N_4253);
nor U5163 (N_5163,N_4411,N_4163);
or U5164 (N_5164,N_4946,N_4137);
nor U5165 (N_5165,N_4973,N_4340);
nor U5166 (N_5166,N_4191,N_4643);
xor U5167 (N_5167,N_4882,N_4777);
nor U5168 (N_5168,N_4529,N_4668);
nor U5169 (N_5169,N_4060,N_4156);
or U5170 (N_5170,N_4438,N_4692);
nor U5171 (N_5171,N_4255,N_4710);
or U5172 (N_5172,N_4834,N_4617);
nor U5173 (N_5173,N_4759,N_4337);
or U5174 (N_5174,N_4081,N_4615);
or U5175 (N_5175,N_4559,N_4644);
or U5176 (N_5176,N_4657,N_4856);
nand U5177 (N_5177,N_4233,N_4049);
nand U5178 (N_5178,N_4220,N_4625);
nand U5179 (N_5179,N_4483,N_4586);
and U5180 (N_5180,N_4116,N_4198);
nand U5181 (N_5181,N_4043,N_4603);
or U5182 (N_5182,N_4003,N_4304);
xnor U5183 (N_5183,N_4087,N_4671);
nand U5184 (N_5184,N_4511,N_4660);
nand U5185 (N_5185,N_4240,N_4602);
xnor U5186 (N_5186,N_4496,N_4502);
or U5187 (N_5187,N_4445,N_4563);
nor U5188 (N_5188,N_4909,N_4999);
and U5189 (N_5189,N_4838,N_4386);
nor U5190 (N_5190,N_4970,N_4621);
and U5191 (N_5191,N_4732,N_4144);
or U5192 (N_5192,N_4022,N_4742);
nor U5193 (N_5193,N_4818,N_4645);
nor U5194 (N_5194,N_4263,N_4952);
and U5195 (N_5195,N_4844,N_4352);
nor U5196 (N_5196,N_4303,N_4279);
nor U5197 (N_5197,N_4605,N_4247);
xnor U5198 (N_5198,N_4961,N_4802);
and U5199 (N_5199,N_4417,N_4527);
xor U5200 (N_5200,N_4323,N_4333);
xnor U5201 (N_5201,N_4488,N_4230);
nand U5202 (N_5202,N_4102,N_4891);
nand U5203 (N_5203,N_4306,N_4716);
or U5204 (N_5204,N_4507,N_4789);
and U5205 (N_5205,N_4878,N_4264);
and U5206 (N_5206,N_4830,N_4183);
and U5207 (N_5207,N_4141,N_4578);
xor U5208 (N_5208,N_4050,N_4867);
nand U5209 (N_5209,N_4080,N_4299);
nand U5210 (N_5210,N_4103,N_4126);
nor U5211 (N_5211,N_4600,N_4989);
nand U5212 (N_5212,N_4118,N_4319);
nand U5213 (N_5213,N_4257,N_4254);
and U5214 (N_5214,N_4119,N_4845);
nand U5215 (N_5215,N_4355,N_4654);
and U5216 (N_5216,N_4332,N_4741);
nand U5217 (N_5217,N_4618,N_4462);
xor U5218 (N_5218,N_4679,N_4001);
or U5219 (N_5219,N_4317,N_4701);
and U5220 (N_5220,N_4278,N_4715);
or U5221 (N_5221,N_4075,N_4837);
nand U5222 (N_5222,N_4085,N_4028);
or U5223 (N_5223,N_4041,N_4140);
or U5224 (N_5224,N_4486,N_4033);
nand U5225 (N_5225,N_4347,N_4953);
nor U5226 (N_5226,N_4986,N_4274);
or U5227 (N_5227,N_4338,N_4610);
nor U5228 (N_5228,N_4167,N_4641);
xor U5229 (N_5229,N_4480,N_4456);
nand U5230 (N_5230,N_4046,N_4992);
or U5231 (N_5231,N_4583,N_4755);
and U5232 (N_5232,N_4712,N_4053);
and U5233 (N_5233,N_4343,N_4164);
or U5234 (N_5234,N_4709,N_4162);
nor U5235 (N_5235,N_4286,N_4604);
xor U5236 (N_5236,N_4262,N_4647);
xor U5237 (N_5237,N_4313,N_4418);
or U5238 (N_5238,N_4993,N_4406);
and U5239 (N_5239,N_4903,N_4877);
nand U5240 (N_5240,N_4261,N_4567);
or U5241 (N_5241,N_4180,N_4745);
and U5242 (N_5242,N_4093,N_4305);
and U5243 (N_5243,N_4975,N_4271);
or U5244 (N_5244,N_4363,N_4289);
nor U5245 (N_5245,N_4139,N_4051);
nand U5246 (N_5246,N_4211,N_4166);
and U5247 (N_5247,N_4635,N_4723);
nand U5248 (N_5248,N_4017,N_4359);
and U5249 (N_5249,N_4728,N_4576);
nand U5250 (N_5250,N_4440,N_4714);
or U5251 (N_5251,N_4251,N_4747);
and U5252 (N_5252,N_4235,N_4072);
xor U5253 (N_5253,N_4590,N_4298);
nor U5254 (N_5254,N_4098,N_4933);
and U5255 (N_5255,N_4720,N_4284);
nand U5256 (N_5256,N_4227,N_4415);
nor U5257 (N_5257,N_4512,N_4757);
nand U5258 (N_5258,N_4736,N_4376);
and U5259 (N_5259,N_4407,N_4357);
and U5260 (N_5260,N_4177,N_4213);
xnor U5261 (N_5261,N_4517,N_4750);
nor U5262 (N_5262,N_4535,N_4925);
xnor U5263 (N_5263,N_4683,N_4965);
or U5264 (N_5264,N_4702,N_4356);
and U5265 (N_5265,N_4857,N_4831);
nand U5266 (N_5266,N_4244,N_4619);
and U5267 (N_5267,N_4016,N_4426);
nand U5268 (N_5268,N_4863,N_4199);
or U5269 (N_5269,N_4436,N_4402);
and U5270 (N_5270,N_4358,N_4971);
nor U5271 (N_5271,N_4494,N_4459);
or U5272 (N_5272,N_4405,N_4784);
nand U5273 (N_5273,N_4455,N_4404);
xor U5274 (N_5274,N_4229,N_4883);
and U5275 (N_5275,N_4387,N_4063);
nor U5276 (N_5276,N_4400,N_4296);
nor U5277 (N_5277,N_4393,N_4804);
or U5278 (N_5278,N_4152,N_4594);
or U5279 (N_5279,N_4964,N_4020);
or U5280 (N_5280,N_4431,N_4127);
and U5281 (N_5281,N_4210,N_4537);
nand U5282 (N_5282,N_4371,N_4658);
nor U5283 (N_5283,N_4822,N_4239);
or U5284 (N_5284,N_4243,N_4173);
nand U5285 (N_5285,N_4269,N_4890);
or U5286 (N_5286,N_4409,N_4009);
and U5287 (N_5287,N_4691,N_4069);
and U5288 (N_5288,N_4258,N_4032);
or U5289 (N_5289,N_4203,N_4185);
xor U5290 (N_5290,N_4842,N_4663);
nor U5291 (N_5291,N_4008,N_4339);
or U5292 (N_5292,N_4187,N_4145);
xnor U5293 (N_5293,N_4007,N_4491);
and U5294 (N_5294,N_4650,N_4982);
xor U5295 (N_5295,N_4071,N_4944);
nand U5296 (N_5296,N_4129,N_4374);
nor U5297 (N_5297,N_4378,N_4991);
nand U5298 (N_5298,N_4495,N_4048);
or U5299 (N_5299,N_4572,N_4216);
or U5300 (N_5300,N_4423,N_4528);
and U5301 (N_5301,N_4694,N_4451);
or U5302 (N_5302,N_4525,N_4432);
or U5303 (N_5303,N_4215,N_4735);
or U5304 (N_5304,N_4573,N_4287);
or U5305 (N_5305,N_4778,N_4609);
nand U5306 (N_5306,N_4695,N_4225);
or U5307 (N_5307,N_4154,N_4756);
or U5308 (N_5308,N_4868,N_4536);
nand U5309 (N_5309,N_4740,N_4078);
nor U5310 (N_5310,N_4272,N_4458);
and U5311 (N_5311,N_4656,N_4142);
nand U5312 (N_5312,N_4148,N_4951);
xor U5313 (N_5313,N_4700,N_4941);
nor U5314 (N_5314,N_4428,N_4484);
nand U5315 (N_5315,N_4770,N_4936);
and U5316 (N_5316,N_4914,N_4675);
and U5317 (N_5317,N_4550,N_4467);
and U5318 (N_5318,N_4880,N_4027);
or U5319 (N_5319,N_4957,N_4579);
and U5320 (N_5320,N_4131,N_4479);
or U5321 (N_5321,N_4194,N_4884);
xor U5322 (N_5322,N_4538,N_4083);
nor U5323 (N_5323,N_4901,N_4294);
nor U5324 (N_5324,N_4739,N_4018);
nand U5325 (N_5325,N_4013,N_4968);
nand U5326 (N_5326,N_4921,N_4886);
and U5327 (N_5327,N_4666,N_4761);
xor U5328 (N_5328,N_4703,N_4509);
nor U5329 (N_5329,N_4939,N_4798);
xor U5330 (N_5330,N_4448,N_4689);
nor U5331 (N_5331,N_4607,N_4531);
or U5332 (N_5332,N_4737,N_4995);
nand U5333 (N_5333,N_4935,N_4113);
xor U5334 (N_5334,N_4012,N_4121);
and U5335 (N_5335,N_4218,N_4336);
nor U5336 (N_5336,N_4311,N_4327);
nor U5337 (N_5337,N_4566,N_4792);
nand U5338 (N_5338,N_4478,N_4569);
nand U5339 (N_5339,N_4249,N_4707);
nor U5340 (N_5340,N_4364,N_4316);
nor U5341 (N_5341,N_4862,N_4962);
nand U5342 (N_5342,N_4955,N_4208);
xor U5343 (N_5343,N_4059,N_4530);
and U5344 (N_5344,N_4623,N_4923);
and U5345 (N_5345,N_4282,N_4290);
xnor U5346 (N_5346,N_4275,N_4539);
or U5347 (N_5347,N_4853,N_4544);
and U5348 (N_5348,N_4176,N_4949);
or U5349 (N_5349,N_4030,N_4242);
or U5350 (N_5350,N_4433,N_4596);
and U5351 (N_5351,N_4522,N_4421);
xnor U5352 (N_5352,N_4651,N_4760);
xor U5353 (N_5353,N_4412,N_4416);
xor U5354 (N_5354,N_4885,N_4414);
nand U5355 (N_5355,N_4835,N_4125);
xnor U5356 (N_5356,N_4956,N_4829);
nor U5357 (N_5357,N_4724,N_4205);
and U5358 (N_5358,N_4021,N_4549);
nand U5359 (N_5359,N_4010,N_4706);
xnor U5360 (N_5360,N_4514,N_4422);
nand U5361 (N_5361,N_4705,N_4781);
and U5362 (N_5362,N_4687,N_4108);
and U5363 (N_5363,N_4561,N_4219);
xor U5364 (N_5364,N_4241,N_4006);
nor U5365 (N_5365,N_4329,N_4283);
nor U5366 (N_5366,N_4498,N_4676);
nor U5367 (N_5367,N_4819,N_4221);
nor U5368 (N_5368,N_4994,N_4599);
xor U5369 (N_5369,N_4037,N_4097);
nor U5370 (N_5370,N_4473,N_4926);
xor U5371 (N_5371,N_4186,N_4774);
nor U5372 (N_5372,N_4153,N_4864);
or U5373 (N_5373,N_4545,N_4688);
xor U5374 (N_5374,N_4066,N_4733);
nor U5375 (N_5375,N_4786,N_4515);
or U5376 (N_5376,N_4082,N_4849);
and U5377 (N_5377,N_4178,N_4112);
xor U5378 (N_5378,N_4906,N_4147);
or U5379 (N_5379,N_4542,N_4398);
xnor U5380 (N_5380,N_4820,N_4058);
nor U5381 (N_5381,N_4500,N_4852);
xor U5382 (N_5382,N_4564,N_4335);
xnor U5383 (N_5383,N_4974,N_4678);
xnor U5384 (N_5384,N_4751,N_4591);
nand U5385 (N_5385,N_4504,N_4420);
and U5386 (N_5386,N_4245,N_4874);
nand U5387 (N_5387,N_4827,N_4214);
or U5388 (N_5388,N_4182,N_4084);
nor U5389 (N_5389,N_4181,N_4128);
and U5390 (N_5390,N_4372,N_4696);
nor U5391 (N_5391,N_4540,N_4554);
or U5392 (N_5392,N_4252,N_4382);
nor U5393 (N_5393,N_4938,N_4309);
xor U5394 (N_5394,N_4192,N_4410);
xnor U5395 (N_5395,N_4399,N_4513);
and U5396 (N_5396,N_4987,N_4916);
and U5397 (N_5397,N_4895,N_4664);
nand U5398 (N_5398,N_4238,N_4680);
nor U5399 (N_5399,N_4876,N_4468);
nand U5400 (N_5400,N_4825,N_4520);
or U5401 (N_5401,N_4246,N_4823);
or U5402 (N_5402,N_4913,N_4435);
xor U5403 (N_5403,N_4260,N_4370);
nand U5404 (N_5404,N_4642,N_4717);
nor U5405 (N_5405,N_4499,N_4089);
or U5406 (N_5406,N_4797,N_4301);
nand U5407 (N_5407,N_4998,N_4172);
or U5408 (N_5408,N_4773,N_4151);
or U5409 (N_5409,N_4136,N_4429);
nand U5410 (N_5410,N_4295,N_4767);
xnor U5411 (N_5411,N_4929,N_4908);
or U5412 (N_5412,N_4887,N_4158);
or U5413 (N_5413,N_4302,N_4146);
or U5414 (N_5414,N_4860,N_4161);
nand U5415 (N_5415,N_4476,N_4808);
and U5416 (N_5416,N_4107,N_4555);
nor U5417 (N_5417,N_4344,N_4632);
xor U5418 (N_5418,N_4110,N_4983);
nand U5419 (N_5419,N_4985,N_4960);
nor U5420 (N_5420,N_4308,N_4470);
or U5421 (N_5421,N_4157,N_4373);
and U5422 (N_5422,N_4521,N_4597);
and U5423 (N_5423,N_4057,N_4950);
and U5424 (N_5424,N_4585,N_4646);
and U5425 (N_5425,N_4444,N_4684);
xor U5426 (N_5426,N_4351,N_4783);
xor U5427 (N_5427,N_4943,N_4785);
nand U5428 (N_5428,N_4014,N_4234);
nor U5429 (N_5429,N_4281,N_4924);
and U5430 (N_5430,N_4930,N_4560);
and U5431 (N_5431,N_4661,N_4815);
nor U5432 (N_5432,N_4114,N_4768);
nand U5433 (N_5433,N_4721,N_4813);
xor U5434 (N_5434,N_4068,N_4729);
or U5435 (N_5435,N_4858,N_4115);
or U5436 (N_5436,N_4004,N_4865);
and U5437 (N_5437,N_4588,N_4222);
xnor U5438 (N_5438,N_4073,N_4277);
or U5439 (N_5439,N_4067,N_4698);
xnor U5440 (N_5440,N_4425,N_4669);
and U5441 (N_5441,N_4582,N_4469);
or U5442 (N_5442,N_4627,N_4159);
or U5443 (N_5443,N_4749,N_4980);
xnor U5444 (N_5444,N_4871,N_4580);
or U5445 (N_5445,N_4408,N_4101);
or U5446 (N_5446,N_4861,N_4872);
nand U5447 (N_5447,N_4109,N_4809);
nand U5448 (N_5448,N_4817,N_4708);
nor U5449 (N_5449,N_4898,N_4188);
nor U5450 (N_5450,N_4450,N_4686);
xor U5451 (N_5451,N_4086,N_4598);
nand U5452 (N_5452,N_4824,N_4318);
nor U5453 (N_5453,N_4369,N_4325);
and U5454 (N_5454,N_4665,N_4259);
xor U5455 (N_5455,N_4812,N_4910);
or U5456 (N_5456,N_4503,N_4394);
nand U5457 (N_5457,N_4485,N_4326);
nor U5458 (N_5458,N_4174,N_4996);
or U5459 (N_5459,N_4593,N_4843);
or U5460 (N_5460,N_4443,N_4460);
nand U5461 (N_5461,N_4300,N_4958);
and U5462 (N_5462,N_4005,N_4349);
xor U5463 (N_5463,N_4775,N_4202);
nand U5464 (N_5464,N_4546,N_4801);
xnor U5465 (N_5465,N_4463,N_4981);
and U5466 (N_5466,N_4292,N_4796);
xnor U5467 (N_5467,N_4437,N_4584);
nor U5468 (N_5468,N_4471,N_4997);
or U5469 (N_5469,N_4011,N_4896);
or U5470 (N_5470,N_4026,N_4900);
or U5471 (N_5471,N_4893,N_4104);
nor U5472 (N_5472,N_4453,N_4575);
and U5473 (N_5473,N_4653,N_4800);
xnor U5474 (N_5474,N_4209,N_4395);
nand U5475 (N_5475,N_4881,N_4754);
and U5476 (N_5476,N_4201,N_4744);
or U5477 (N_5477,N_4270,N_4441);
and U5478 (N_5478,N_4931,N_4655);
and U5479 (N_5479,N_4493,N_4092);
nor U5480 (N_5480,N_4769,N_4482);
nor U5481 (N_5481,N_4519,N_4052);
or U5482 (N_5482,N_4348,N_4143);
xor U5483 (N_5483,N_4424,N_4854);
xor U5484 (N_5484,N_4236,N_4551);
or U5485 (N_5485,N_4558,N_4193);
xor U5486 (N_5486,N_4165,N_4601);
and U5487 (N_5487,N_4442,N_4556);
nand U5488 (N_5488,N_4155,N_4250);
nor U5489 (N_5489,N_4330,N_4628);
or U5490 (N_5490,N_4810,N_4516);
xnor U5491 (N_5491,N_4648,N_4606);
xnor U5492 (N_5492,N_4124,N_4693);
xnor U5493 (N_5493,N_4457,N_4762);
xor U5494 (N_5494,N_4280,N_4055);
nor U5495 (N_5495,N_4771,N_4090);
or U5496 (N_5496,N_4821,N_4616);
nand U5497 (N_5497,N_4505,N_4489);
xor U5498 (N_5498,N_4932,N_4138);
nand U5499 (N_5499,N_4795,N_4076);
nand U5500 (N_5500,N_4566,N_4774);
nand U5501 (N_5501,N_4808,N_4317);
nand U5502 (N_5502,N_4065,N_4199);
xnor U5503 (N_5503,N_4284,N_4509);
or U5504 (N_5504,N_4471,N_4776);
xor U5505 (N_5505,N_4190,N_4096);
nand U5506 (N_5506,N_4624,N_4802);
or U5507 (N_5507,N_4073,N_4539);
nor U5508 (N_5508,N_4997,N_4616);
and U5509 (N_5509,N_4525,N_4933);
and U5510 (N_5510,N_4418,N_4871);
and U5511 (N_5511,N_4197,N_4079);
xor U5512 (N_5512,N_4605,N_4558);
and U5513 (N_5513,N_4003,N_4328);
xor U5514 (N_5514,N_4570,N_4625);
nor U5515 (N_5515,N_4418,N_4958);
and U5516 (N_5516,N_4633,N_4911);
nor U5517 (N_5517,N_4606,N_4088);
xor U5518 (N_5518,N_4365,N_4701);
nor U5519 (N_5519,N_4472,N_4567);
nor U5520 (N_5520,N_4409,N_4350);
nor U5521 (N_5521,N_4524,N_4762);
xor U5522 (N_5522,N_4147,N_4786);
nand U5523 (N_5523,N_4667,N_4057);
nand U5524 (N_5524,N_4334,N_4120);
and U5525 (N_5525,N_4131,N_4429);
or U5526 (N_5526,N_4953,N_4548);
or U5527 (N_5527,N_4721,N_4456);
nor U5528 (N_5528,N_4067,N_4952);
nor U5529 (N_5529,N_4757,N_4722);
nand U5530 (N_5530,N_4176,N_4595);
or U5531 (N_5531,N_4661,N_4940);
nand U5532 (N_5532,N_4473,N_4681);
and U5533 (N_5533,N_4632,N_4880);
and U5534 (N_5534,N_4737,N_4720);
nor U5535 (N_5535,N_4882,N_4873);
nand U5536 (N_5536,N_4689,N_4799);
nand U5537 (N_5537,N_4900,N_4739);
xnor U5538 (N_5538,N_4176,N_4358);
and U5539 (N_5539,N_4960,N_4388);
nor U5540 (N_5540,N_4019,N_4079);
nand U5541 (N_5541,N_4692,N_4904);
xnor U5542 (N_5542,N_4061,N_4057);
and U5543 (N_5543,N_4593,N_4642);
or U5544 (N_5544,N_4183,N_4116);
xor U5545 (N_5545,N_4957,N_4445);
xnor U5546 (N_5546,N_4798,N_4732);
nor U5547 (N_5547,N_4901,N_4196);
or U5548 (N_5548,N_4277,N_4248);
and U5549 (N_5549,N_4686,N_4077);
xnor U5550 (N_5550,N_4081,N_4980);
xnor U5551 (N_5551,N_4822,N_4509);
nor U5552 (N_5552,N_4363,N_4249);
nand U5553 (N_5553,N_4515,N_4642);
and U5554 (N_5554,N_4268,N_4699);
or U5555 (N_5555,N_4602,N_4639);
or U5556 (N_5556,N_4773,N_4474);
or U5557 (N_5557,N_4809,N_4521);
nand U5558 (N_5558,N_4607,N_4026);
nor U5559 (N_5559,N_4895,N_4174);
nor U5560 (N_5560,N_4414,N_4325);
nor U5561 (N_5561,N_4268,N_4331);
xnor U5562 (N_5562,N_4273,N_4755);
or U5563 (N_5563,N_4479,N_4617);
and U5564 (N_5564,N_4874,N_4453);
xor U5565 (N_5565,N_4474,N_4563);
and U5566 (N_5566,N_4924,N_4235);
nor U5567 (N_5567,N_4676,N_4674);
nand U5568 (N_5568,N_4189,N_4919);
nor U5569 (N_5569,N_4111,N_4509);
or U5570 (N_5570,N_4306,N_4024);
nand U5571 (N_5571,N_4166,N_4250);
nor U5572 (N_5572,N_4148,N_4503);
xnor U5573 (N_5573,N_4211,N_4174);
xnor U5574 (N_5574,N_4133,N_4225);
nand U5575 (N_5575,N_4153,N_4028);
xor U5576 (N_5576,N_4833,N_4316);
xor U5577 (N_5577,N_4599,N_4363);
and U5578 (N_5578,N_4864,N_4962);
nand U5579 (N_5579,N_4965,N_4496);
and U5580 (N_5580,N_4702,N_4321);
and U5581 (N_5581,N_4400,N_4244);
and U5582 (N_5582,N_4950,N_4230);
and U5583 (N_5583,N_4747,N_4312);
and U5584 (N_5584,N_4825,N_4795);
or U5585 (N_5585,N_4954,N_4086);
nor U5586 (N_5586,N_4024,N_4788);
nand U5587 (N_5587,N_4709,N_4999);
and U5588 (N_5588,N_4533,N_4653);
or U5589 (N_5589,N_4606,N_4253);
xor U5590 (N_5590,N_4012,N_4685);
or U5591 (N_5591,N_4252,N_4110);
nor U5592 (N_5592,N_4035,N_4908);
nor U5593 (N_5593,N_4268,N_4201);
or U5594 (N_5594,N_4437,N_4442);
and U5595 (N_5595,N_4664,N_4773);
or U5596 (N_5596,N_4428,N_4998);
nand U5597 (N_5597,N_4880,N_4944);
xnor U5598 (N_5598,N_4017,N_4316);
nor U5599 (N_5599,N_4693,N_4152);
nand U5600 (N_5600,N_4232,N_4060);
xnor U5601 (N_5601,N_4919,N_4885);
or U5602 (N_5602,N_4257,N_4144);
nor U5603 (N_5603,N_4354,N_4468);
and U5604 (N_5604,N_4288,N_4438);
xor U5605 (N_5605,N_4353,N_4942);
and U5606 (N_5606,N_4404,N_4565);
or U5607 (N_5607,N_4487,N_4654);
xnor U5608 (N_5608,N_4157,N_4748);
nor U5609 (N_5609,N_4180,N_4473);
nor U5610 (N_5610,N_4720,N_4217);
nand U5611 (N_5611,N_4646,N_4099);
nand U5612 (N_5612,N_4758,N_4436);
xnor U5613 (N_5613,N_4816,N_4113);
or U5614 (N_5614,N_4775,N_4510);
and U5615 (N_5615,N_4182,N_4243);
and U5616 (N_5616,N_4148,N_4335);
xnor U5617 (N_5617,N_4165,N_4179);
or U5618 (N_5618,N_4447,N_4819);
or U5619 (N_5619,N_4500,N_4038);
and U5620 (N_5620,N_4066,N_4448);
or U5621 (N_5621,N_4232,N_4138);
or U5622 (N_5622,N_4747,N_4337);
or U5623 (N_5623,N_4451,N_4541);
nor U5624 (N_5624,N_4355,N_4111);
and U5625 (N_5625,N_4457,N_4650);
nor U5626 (N_5626,N_4641,N_4309);
and U5627 (N_5627,N_4288,N_4958);
nand U5628 (N_5628,N_4808,N_4377);
or U5629 (N_5629,N_4095,N_4235);
or U5630 (N_5630,N_4738,N_4410);
or U5631 (N_5631,N_4998,N_4262);
xnor U5632 (N_5632,N_4429,N_4106);
xor U5633 (N_5633,N_4746,N_4788);
or U5634 (N_5634,N_4621,N_4377);
and U5635 (N_5635,N_4383,N_4661);
nand U5636 (N_5636,N_4188,N_4638);
or U5637 (N_5637,N_4799,N_4951);
nand U5638 (N_5638,N_4681,N_4277);
xor U5639 (N_5639,N_4158,N_4400);
and U5640 (N_5640,N_4549,N_4683);
nand U5641 (N_5641,N_4063,N_4215);
xor U5642 (N_5642,N_4660,N_4594);
xnor U5643 (N_5643,N_4852,N_4404);
nor U5644 (N_5644,N_4724,N_4225);
or U5645 (N_5645,N_4734,N_4263);
or U5646 (N_5646,N_4706,N_4890);
xor U5647 (N_5647,N_4164,N_4282);
nand U5648 (N_5648,N_4006,N_4513);
nor U5649 (N_5649,N_4995,N_4581);
and U5650 (N_5650,N_4303,N_4894);
nor U5651 (N_5651,N_4028,N_4957);
nand U5652 (N_5652,N_4355,N_4475);
nor U5653 (N_5653,N_4765,N_4414);
nor U5654 (N_5654,N_4400,N_4067);
or U5655 (N_5655,N_4402,N_4895);
nor U5656 (N_5656,N_4689,N_4073);
or U5657 (N_5657,N_4378,N_4710);
nor U5658 (N_5658,N_4946,N_4198);
or U5659 (N_5659,N_4250,N_4464);
nand U5660 (N_5660,N_4247,N_4631);
or U5661 (N_5661,N_4082,N_4716);
nor U5662 (N_5662,N_4309,N_4985);
nand U5663 (N_5663,N_4944,N_4892);
xnor U5664 (N_5664,N_4653,N_4902);
nand U5665 (N_5665,N_4531,N_4192);
or U5666 (N_5666,N_4044,N_4227);
and U5667 (N_5667,N_4705,N_4028);
or U5668 (N_5668,N_4924,N_4297);
nand U5669 (N_5669,N_4258,N_4767);
nand U5670 (N_5670,N_4312,N_4021);
and U5671 (N_5671,N_4229,N_4727);
and U5672 (N_5672,N_4096,N_4830);
xor U5673 (N_5673,N_4357,N_4945);
and U5674 (N_5674,N_4179,N_4495);
and U5675 (N_5675,N_4248,N_4569);
nand U5676 (N_5676,N_4703,N_4863);
xor U5677 (N_5677,N_4936,N_4593);
nor U5678 (N_5678,N_4830,N_4660);
or U5679 (N_5679,N_4713,N_4400);
xnor U5680 (N_5680,N_4927,N_4070);
nand U5681 (N_5681,N_4281,N_4581);
or U5682 (N_5682,N_4255,N_4026);
and U5683 (N_5683,N_4819,N_4300);
nor U5684 (N_5684,N_4747,N_4053);
and U5685 (N_5685,N_4340,N_4771);
or U5686 (N_5686,N_4620,N_4071);
nor U5687 (N_5687,N_4315,N_4087);
and U5688 (N_5688,N_4299,N_4466);
or U5689 (N_5689,N_4696,N_4806);
and U5690 (N_5690,N_4861,N_4772);
or U5691 (N_5691,N_4155,N_4646);
and U5692 (N_5692,N_4058,N_4351);
nor U5693 (N_5693,N_4956,N_4262);
nor U5694 (N_5694,N_4213,N_4206);
nor U5695 (N_5695,N_4507,N_4370);
nand U5696 (N_5696,N_4760,N_4311);
or U5697 (N_5697,N_4439,N_4946);
nand U5698 (N_5698,N_4396,N_4612);
or U5699 (N_5699,N_4000,N_4666);
or U5700 (N_5700,N_4266,N_4049);
and U5701 (N_5701,N_4696,N_4015);
xnor U5702 (N_5702,N_4786,N_4102);
or U5703 (N_5703,N_4566,N_4357);
and U5704 (N_5704,N_4823,N_4047);
nor U5705 (N_5705,N_4327,N_4881);
xor U5706 (N_5706,N_4202,N_4615);
xor U5707 (N_5707,N_4662,N_4525);
or U5708 (N_5708,N_4438,N_4686);
nor U5709 (N_5709,N_4289,N_4692);
nor U5710 (N_5710,N_4752,N_4710);
and U5711 (N_5711,N_4237,N_4350);
or U5712 (N_5712,N_4561,N_4932);
nor U5713 (N_5713,N_4386,N_4365);
xor U5714 (N_5714,N_4297,N_4728);
xor U5715 (N_5715,N_4520,N_4655);
and U5716 (N_5716,N_4841,N_4848);
and U5717 (N_5717,N_4737,N_4841);
xor U5718 (N_5718,N_4647,N_4750);
and U5719 (N_5719,N_4903,N_4516);
nand U5720 (N_5720,N_4467,N_4701);
nor U5721 (N_5721,N_4024,N_4654);
nand U5722 (N_5722,N_4420,N_4619);
nand U5723 (N_5723,N_4882,N_4912);
xnor U5724 (N_5724,N_4183,N_4720);
nor U5725 (N_5725,N_4046,N_4759);
and U5726 (N_5726,N_4293,N_4202);
or U5727 (N_5727,N_4133,N_4497);
nand U5728 (N_5728,N_4473,N_4182);
or U5729 (N_5729,N_4329,N_4247);
or U5730 (N_5730,N_4323,N_4745);
or U5731 (N_5731,N_4530,N_4181);
or U5732 (N_5732,N_4779,N_4856);
and U5733 (N_5733,N_4105,N_4475);
nand U5734 (N_5734,N_4767,N_4391);
or U5735 (N_5735,N_4188,N_4576);
and U5736 (N_5736,N_4217,N_4091);
xor U5737 (N_5737,N_4773,N_4095);
nand U5738 (N_5738,N_4740,N_4312);
nand U5739 (N_5739,N_4228,N_4389);
or U5740 (N_5740,N_4922,N_4814);
nor U5741 (N_5741,N_4968,N_4682);
or U5742 (N_5742,N_4830,N_4146);
nor U5743 (N_5743,N_4820,N_4851);
xnor U5744 (N_5744,N_4907,N_4594);
or U5745 (N_5745,N_4192,N_4667);
nand U5746 (N_5746,N_4004,N_4796);
xor U5747 (N_5747,N_4610,N_4423);
and U5748 (N_5748,N_4849,N_4393);
xnor U5749 (N_5749,N_4539,N_4591);
nor U5750 (N_5750,N_4501,N_4443);
or U5751 (N_5751,N_4633,N_4277);
or U5752 (N_5752,N_4086,N_4704);
xor U5753 (N_5753,N_4709,N_4144);
and U5754 (N_5754,N_4656,N_4444);
or U5755 (N_5755,N_4139,N_4965);
nor U5756 (N_5756,N_4103,N_4016);
and U5757 (N_5757,N_4518,N_4846);
and U5758 (N_5758,N_4399,N_4667);
or U5759 (N_5759,N_4908,N_4457);
or U5760 (N_5760,N_4479,N_4021);
nand U5761 (N_5761,N_4151,N_4393);
and U5762 (N_5762,N_4261,N_4634);
nand U5763 (N_5763,N_4932,N_4069);
xnor U5764 (N_5764,N_4920,N_4832);
and U5765 (N_5765,N_4840,N_4187);
and U5766 (N_5766,N_4071,N_4160);
and U5767 (N_5767,N_4265,N_4008);
or U5768 (N_5768,N_4388,N_4341);
nor U5769 (N_5769,N_4130,N_4943);
nor U5770 (N_5770,N_4437,N_4708);
and U5771 (N_5771,N_4273,N_4930);
or U5772 (N_5772,N_4085,N_4474);
and U5773 (N_5773,N_4460,N_4547);
or U5774 (N_5774,N_4516,N_4153);
xnor U5775 (N_5775,N_4376,N_4655);
or U5776 (N_5776,N_4694,N_4631);
nor U5777 (N_5777,N_4935,N_4408);
xor U5778 (N_5778,N_4699,N_4060);
xnor U5779 (N_5779,N_4650,N_4608);
and U5780 (N_5780,N_4063,N_4788);
nand U5781 (N_5781,N_4610,N_4350);
xor U5782 (N_5782,N_4780,N_4011);
nand U5783 (N_5783,N_4356,N_4123);
and U5784 (N_5784,N_4667,N_4715);
or U5785 (N_5785,N_4359,N_4814);
and U5786 (N_5786,N_4021,N_4719);
nor U5787 (N_5787,N_4155,N_4046);
xor U5788 (N_5788,N_4008,N_4507);
nor U5789 (N_5789,N_4571,N_4718);
or U5790 (N_5790,N_4060,N_4285);
nand U5791 (N_5791,N_4284,N_4771);
nand U5792 (N_5792,N_4767,N_4329);
xnor U5793 (N_5793,N_4854,N_4585);
nor U5794 (N_5794,N_4518,N_4307);
nand U5795 (N_5795,N_4781,N_4588);
and U5796 (N_5796,N_4707,N_4487);
or U5797 (N_5797,N_4912,N_4389);
nor U5798 (N_5798,N_4606,N_4760);
nand U5799 (N_5799,N_4200,N_4835);
xor U5800 (N_5800,N_4573,N_4955);
xnor U5801 (N_5801,N_4024,N_4334);
or U5802 (N_5802,N_4354,N_4212);
xor U5803 (N_5803,N_4513,N_4719);
and U5804 (N_5804,N_4362,N_4182);
and U5805 (N_5805,N_4637,N_4148);
or U5806 (N_5806,N_4436,N_4596);
nand U5807 (N_5807,N_4778,N_4023);
and U5808 (N_5808,N_4052,N_4354);
nand U5809 (N_5809,N_4846,N_4517);
and U5810 (N_5810,N_4887,N_4572);
and U5811 (N_5811,N_4986,N_4293);
xor U5812 (N_5812,N_4691,N_4817);
and U5813 (N_5813,N_4944,N_4874);
nand U5814 (N_5814,N_4788,N_4351);
xor U5815 (N_5815,N_4947,N_4932);
or U5816 (N_5816,N_4852,N_4104);
xnor U5817 (N_5817,N_4519,N_4143);
nand U5818 (N_5818,N_4375,N_4689);
or U5819 (N_5819,N_4156,N_4984);
and U5820 (N_5820,N_4156,N_4919);
nor U5821 (N_5821,N_4975,N_4489);
nor U5822 (N_5822,N_4237,N_4225);
xnor U5823 (N_5823,N_4034,N_4602);
and U5824 (N_5824,N_4566,N_4647);
xor U5825 (N_5825,N_4340,N_4628);
nor U5826 (N_5826,N_4861,N_4161);
nand U5827 (N_5827,N_4646,N_4225);
and U5828 (N_5828,N_4986,N_4502);
nor U5829 (N_5829,N_4578,N_4525);
or U5830 (N_5830,N_4929,N_4670);
nor U5831 (N_5831,N_4210,N_4601);
xor U5832 (N_5832,N_4227,N_4331);
nand U5833 (N_5833,N_4732,N_4358);
or U5834 (N_5834,N_4916,N_4343);
or U5835 (N_5835,N_4697,N_4662);
or U5836 (N_5836,N_4953,N_4638);
or U5837 (N_5837,N_4989,N_4243);
and U5838 (N_5838,N_4459,N_4771);
nor U5839 (N_5839,N_4489,N_4909);
xor U5840 (N_5840,N_4003,N_4438);
xnor U5841 (N_5841,N_4180,N_4349);
and U5842 (N_5842,N_4106,N_4844);
nor U5843 (N_5843,N_4397,N_4758);
xor U5844 (N_5844,N_4553,N_4965);
xnor U5845 (N_5845,N_4254,N_4569);
nand U5846 (N_5846,N_4901,N_4845);
xor U5847 (N_5847,N_4750,N_4753);
or U5848 (N_5848,N_4912,N_4837);
or U5849 (N_5849,N_4909,N_4464);
xor U5850 (N_5850,N_4539,N_4375);
xnor U5851 (N_5851,N_4405,N_4346);
xnor U5852 (N_5852,N_4037,N_4505);
nand U5853 (N_5853,N_4099,N_4476);
or U5854 (N_5854,N_4155,N_4662);
nand U5855 (N_5855,N_4486,N_4771);
and U5856 (N_5856,N_4738,N_4300);
nand U5857 (N_5857,N_4525,N_4463);
and U5858 (N_5858,N_4817,N_4065);
and U5859 (N_5859,N_4814,N_4154);
nand U5860 (N_5860,N_4244,N_4160);
xnor U5861 (N_5861,N_4104,N_4265);
and U5862 (N_5862,N_4829,N_4467);
nand U5863 (N_5863,N_4108,N_4992);
or U5864 (N_5864,N_4011,N_4023);
and U5865 (N_5865,N_4589,N_4090);
nor U5866 (N_5866,N_4763,N_4289);
xnor U5867 (N_5867,N_4631,N_4784);
nand U5868 (N_5868,N_4420,N_4068);
and U5869 (N_5869,N_4505,N_4914);
xor U5870 (N_5870,N_4062,N_4596);
or U5871 (N_5871,N_4326,N_4338);
and U5872 (N_5872,N_4770,N_4997);
or U5873 (N_5873,N_4014,N_4997);
xnor U5874 (N_5874,N_4939,N_4933);
nand U5875 (N_5875,N_4792,N_4082);
and U5876 (N_5876,N_4130,N_4282);
and U5877 (N_5877,N_4457,N_4636);
and U5878 (N_5878,N_4692,N_4352);
xor U5879 (N_5879,N_4913,N_4981);
and U5880 (N_5880,N_4197,N_4717);
and U5881 (N_5881,N_4304,N_4464);
or U5882 (N_5882,N_4685,N_4772);
nand U5883 (N_5883,N_4050,N_4418);
xnor U5884 (N_5884,N_4234,N_4989);
and U5885 (N_5885,N_4935,N_4904);
nor U5886 (N_5886,N_4262,N_4414);
nand U5887 (N_5887,N_4279,N_4041);
xnor U5888 (N_5888,N_4799,N_4622);
or U5889 (N_5889,N_4788,N_4860);
nor U5890 (N_5890,N_4286,N_4352);
or U5891 (N_5891,N_4005,N_4350);
nand U5892 (N_5892,N_4736,N_4286);
and U5893 (N_5893,N_4478,N_4142);
and U5894 (N_5894,N_4873,N_4162);
xnor U5895 (N_5895,N_4978,N_4106);
and U5896 (N_5896,N_4723,N_4795);
nor U5897 (N_5897,N_4767,N_4440);
xor U5898 (N_5898,N_4328,N_4700);
xor U5899 (N_5899,N_4351,N_4121);
or U5900 (N_5900,N_4687,N_4735);
xor U5901 (N_5901,N_4647,N_4358);
or U5902 (N_5902,N_4820,N_4370);
or U5903 (N_5903,N_4643,N_4902);
or U5904 (N_5904,N_4475,N_4118);
nand U5905 (N_5905,N_4405,N_4379);
or U5906 (N_5906,N_4245,N_4901);
nand U5907 (N_5907,N_4435,N_4933);
nand U5908 (N_5908,N_4685,N_4414);
and U5909 (N_5909,N_4874,N_4189);
or U5910 (N_5910,N_4840,N_4090);
or U5911 (N_5911,N_4197,N_4458);
xor U5912 (N_5912,N_4741,N_4066);
and U5913 (N_5913,N_4871,N_4215);
and U5914 (N_5914,N_4337,N_4615);
and U5915 (N_5915,N_4179,N_4690);
nand U5916 (N_5916,N_4697,N_4532);
xor U5917 (N_5917,N_4631,N_4725);
and U5918 (N_5918,N_4919,N_4529);
nand U5919 (N_5919,N_4167,N_4964);
and U5920 (N_5920,N_4326,N_4450);
or U5921 (N_5921,N_4545,N_4939);
nor U5922 (N_5922,N_4066,N_4388);
nor U5923 (N_5923,N_4186,N_4855);
xor U5924 (N_5924,N_4591,N_4146);
nand U5925 (N_5925,N_4227,N_4673);
and U5926 (N_5926,N_4389,N_4172);
or U5927 (N_5927,N_4894,N_4958);
nand U5928 (N_5928,N_4742,N_4354);
xnor U5929 (N_5929,N_4733,N_4877);
nor U5930 (N_5930,N_4031,N_4301);
xor U5931 (N_5931,N_4450,N_4575);
or U5932 (N_5932,N_4744,N_4506);
and U5933 (N_5933,N_4653,N_4750);
xnor U5934 (N_5934,N_4788,N_4185);
or U5935 (N_5935,N_4383,N_4410);
xnor U5936 (N_5936,N_4403,N_4340);
or U5937 (N_5937,N_4135,N_4116);
nor U5938 (N_5938,N_4829,N_4488);
nor U5939 (N_5939,N_4429,N_4542);
xor U5940 (N_5940,N_4996,N_4555);
or U5941 (N_5941,N_4448,N_4458);
nand U5942 (N_5942,N_4317,N_4243);
nor U5943 (N_5943,N_4318,N_4725);
or U5944 (N_5944,N_4923,N_4997);
xnor U5945 (N_5945,N_4922,N_4490);
nand U5946 (N_5946,N_4065,N_4608);
or U5947 (N_5947,N_4635,N_4831);
and U5948 (N_5948,N_4471,N_4867);
xor U5949 (N_5949,N_4660,N_4849);
or U5950 (N_5950,N_4787,N_4905);
and U5951 (N_5951,N_4417,N_4020);
xnor U5952 (N_5952,N_4514,N_4671);
nor U5953 (N_5953,N_4561,N_4951);
and U5954 (N_5954,N_4201,N_4672);
and U5955 (N_5955,N_4683,N_4966);
xnor U5956 (N_5956,N_4183,N_4355);
nand U5957 (N_5957,N_4107,N_4765);
nor U5958 (N_5958,N_4288,N_4756);
nand U5959 (N_5959,N_4389,N_4318);
or U5960 (N_5960,N_4097,N_4384);
xnor U5961 (N_5961,N_4791,N_4457);
and U5962 (N_5962,N_4582,N_4715);
or U5963 (N_5963,N_4788,N_4211);
nand U5964 (N_5964,N_4394,N_4674);
and U5965 (N_5965,N_4425,N_4304);
and U5966 (N_5966,N_4858,N_4766);
nand U5967 (N_5967,N_4030,N_4457);
or U5968 (N_5968,N_4960,N_4257);
nor U5969 (N_5969,N_4522,N_4367);
and U5970 (N_5970,N_4207,N_4759);
xnor U5971 (N_5971,N_4116,N_4686);
or U5972 (N_5972,N_4638,N_4995);
nor U5973 (N_5973,N_4847,N_4200);
or U5974 (N_5974,N_4190,N_4518);
and U5975 (N_5975,N_4407,N_4087);
nor U5976 (N_5976,N_4034,N_4429);
and U5977 (N_5977,N_4419,N_4101);
nor U5978 (N_5978,N_4098,N_4387);
and U5979 (N_5979,N_4094,N_4340);
or U5980 (N_5980,N_4020,N_4403);
xnor U5981 (N_5981,N_4726,N_4844);
nand U5982 (N_5982,N_4880,N_4600);
and U5983 (N_5983,N_4599,N_4141);
nor U5984 (N_5984,N_4131,N_4908);
xnor U5985 (N_5985,N_4455,N_4537);
xnor U5986 (N_5986,N_4537,N_4502);
or U5987 (N_5987,N_4019,N_4645);
xnor U5988 (N_5988,N_4990,N_4289);
or U5989 (N_5989,N_4852,N_4802);
nand U5990 (N_5990,N_4068,N_4117);
nand U5991 (N_5991,N_4697,N_4321);
nand U5992 (N_5992,N_4963,N_4137);
xor U5993 (N_5993,N_4896,N_4766);
nor U5994 (N_5994,N_4628,N_4980);
or U5995 (N_5995,N_4631,N_4855);
nand U5996 (N_5996,N_4212,N_4535);
nand U5997 (N_5997,N_4836,N_4183);
nand U5998 (N_5998,N_4711,N_4169);
and U5999 (N_5999,N_4350,N_4033);
nand U6000 (N_6000,N_5064,N_5015);
or U6001 (N_6001,N_5002,N_5327);
nand U6002 (N_6002,N_5631,N_5340);
xor U6003 (N_6003,N_5962,N_5928);
xnor U6004 (N_6004,N_5828,N_5841);
xnor U6005 (N_6005,N_5212,N_5537);
or U6006 (N_6006,N_5087,N_5813);
nand U6007 (N_6007,N_5436,N_5502);
or U6008 (N_6008,N_5782,N_5716);
nor U6009 (N_6009,N_5923,N_5777);
nand U6010 (N_6010,N_5945,N_5377);
nor U6011 (N_6011,N_5897,N_5235);
or U6012 (N_6012,N_5872,N_5299);
nor U6013 (N_6013,N_5698,N_5362);
nand U6014 (N_6014,N_5198,N_5162);
xor U6015 (N_6015,N_5544,N_5428);
or U6016 (N_6016,N_5865,N_5637);
nand U6017 (N_6017,N_5839,N_5425);
or U6018 (N_6018,N_5925,N_5219);
or U6019 (N_6019,N_5496,N_5338);
or U6020 (N_6020,N_5442,N_5969);
xor U6021 (N_6021,N_5846,N_5430);
xor U6022 (N_6022,N_5244,N_5313);
nor U6023 (N_6023,N_5890,N_5439);
xnor U6024 (N_6024,N_5447,N_5385);
xnor U6025 (N_6025,N_5984,N_5312);
nor U6026 (N_6026,N_5184,N_5337);
nor U6027 (N_6027,N_5717,N_5729);
nor U6028 (N_6028,N_5810,N_5909);
or U6029 (N_6029,N_5226,N_5167);
nand U6030 (N_6030,N_5530,N_5268);
nand U6031 (N_6031,N_5180,N_5793);
and U6032 (N_6032,N_5787,N_5613);
nor U6033 (N_6033,N_5424,N_5001);
or U6034 (N_6034,N_5189,N_5014);
and U6035 (N_6035,N_5382,N_5889);
nand U6036 (N_6036,N_5566,N_5645);
and U6037 (N_6037,N_5205,N_5141);
nand U6038 (N_6038,N_5877,N_5641);
nand U6039 (N_6039,N_5917,N_5241);
xor U6040 (N_6040,N_5183,N_5927);
and U6041 (N_6041,N_5310,N_5602);
and U6042 (N_6042,N_5368,N_5719);
nor U6043 (N_6043,N_5517,N_5375);
nand U6044 (N_6044,N_5459,N_5868);
or U6045 (N_6045,N_5685,N_5123);
nand U6046 (N_6046,N_5915,N_5239);
nor U6047 (N_6047,N_5990,N_5113);
xnor U6048 (N_6048,N_5900,N_5343);
or U6049 (N_6049,N_5253,N_5630);
nand U6050 (N_6050,N_5161,N_5030);
nor U6051 (N_6051,N_5888,N_5831);
nor U6052 (N_6052,N_5472,N_5699);
nor U6053 (N_6053,N_5899,N_5781);
or U6054 (N_6054,N_5947,N_5484);
and U6055 (N_6055,N_5832,N_5322);
nand U6056 (N_6056,N_5732,N_5379);
or U6057 (N_6057,N_5309,N_5154);
and U6058 (N_6058,N_5854,N_5657);
or U6059 (N_6059,N_5245,N_5640);
nor U6060 (N_6060,N_5743,N_5512);
xor U6061 (N_6061,N_5153,N_5911);
nor U6062 (N_6062,N_5993,N_5648);
xnor U6063 (N_6063,N_5039,N_5125);
nand U6064 (N_6064,N_5871,N_5879);
nand U6065 (N_6065,N_5936,N_5274);
nand U6066 (N_6066,N_5816,N_5258);
nor U6067 (N_6067,N_5776,N_5429);
or U6068 (N_6068,N_5407,N_5821);
nor U6069 (N_6069,N_5131,N_5187);
xor U6070 (N_6070,N_5966,N_5228);
or U6071 (N_6071,N_5427,N_5804);
or U6072 (N_6072,N_5778,N_5000);
or U6073 (N_6073,N_5214,N_5220);
xnor U6074 (N_6074,N_5022,N_5599);
and U6075 (N_6075,N_5166,N_5453);
nand U6076 (N_6076,N_5152,N_5088);
or U6077 (N_6077,N_5119,N_5647);
xnor U6078 (N_6078,N_5702,N_5934);
nor U6079 (N_6079,N_5878,N_5416);
and U6080 (N_6080,N_5977,N_5838);
nand U6081 (N_6081,N_5133,N_5972);
or U6082 (N_6082,N_5792,N_5315);
nand U6083 (N_6083,N_5417,N_5097);
and U6084 (N_6084,N_5513,N_5096);
nor U6085 (N_6085,N_5789,N_5948);
nand U6086 (N_6086,N_5823,N_5847);
xnor U6087 (N_6087,N_5303,N_5500);
and U6088 (N_6088,N_5297,N_5869);
xnor U6089 (N_6089,N_5882,N_5651);
nor U6090 (N_6090,N_5745,N_5819);
or U6091 (N_6091,N_5277,N_5979);
xor U6092 (N_6092,N_5388,N_5485);
nor U6093 (N_6093,N_5255,N_5207);
or U6094 (N_6094,N_5766,N_5373);
nor U6095 (N_6095,N_5494,N_5815);
or U6096 (N_6096,N_5861,N_5107);
xnor U6097 (N_6097,N_5524,N_5558);
or U6098 (N_6098,N_5314,N_5506);
nor U6099 (N_6099,N_5486,N_5068);
nor U6100 (N_6100,N_5089,N_5413);
nand U6101 (N_6101,N_5720,N_5755);
or U6102 (N_6102,N_5772,N_5455);
or U6103 (N_6103,N_5248,N_5907);
and U6104 (N_6104,N_5072,N_5522);
and U6105 (N_6105,N_5985,N_5626);
xor U6106 (N_6106,N_5468,N_5686);
nor U6107 (N_6107,N_5604,N_5767);
nor U6108 (N_6108,N_5067,N_5175);
or U6109 (N_6109,N_5176,N_5643);
nand U6110 (N_6110,N_5148,N_5996);
xnor U6111 (N_6111,N_5735,N_5572);
and U6112 (N_6112,N_5462,N_5234);
xnor U6113 (N_6113,N_5760,N_5177);
xor U6114 (N_6114,N_5901,N_5935);
nand U6115 (N_6115,N_5575,N_5178);
and U6116 (N_6116,N_5858,N_5197);
nand U6117 (N_6117,N_5667,N_5902);
nor U6118 (N_6118,N_5445,N_5045);
xor U6119 (N_6119,N_5510,N_5862);
and U6120 (N_6120,N_5672,N_5357);
nand U6121 (N_6121,N_5393,N_5541);
nand U6122 (N_6122,N_5024,N_5655);
nor U6123 (N_6123,N_5976,N_5543);
nor U6124 (N_6124,N_5712,N_5975);
xnor U6125 (N_6125,N_5098,N_5264);
nand U6126 (N_6126,N_5301,N_5344);
and U6127 (N_6127,N_5050,N_5689);
nand U6128 (N_6128,N_5551,N_5389);
xor U6129 (N_6129,N_5267,N_5801);
xor U6130 (N_6130,N_5112,N_5329);
nand U6131 (N_6131,N_5079,N_5086);
nand U6132 (N_6132,N_5070,N_5246);
or U6133 (N_6133,N_5055,N_5281);
xnor U6134 (N_6134,N_5955,N_5908);
nor U6135 (N_6135,N_5798,N_5155);
nor U6136 (N_6136,N_5412,N_5761);
xor U6137 (N_6137,N_5410,N_5342);
nor U6138 (N_6138,N_5678,N_5031);
nand U6139 (N_6139,N_5283,N_5179);
nor U6140 (N_6140,N_5880,N_5622);
nor U6141 (N_6141,N_5632,N_5276);
nor U6142 (N_6142,N_5608,N_5538);
or U6143 (N_6143,N_5010,N_5914);
or U6144 (N_6144,N_5399,N_5415);
and U6145 (N_6145,N_5690,N_5949);
xnor U6146 (N_6146,N_5104,N_5581);
or U6147 (N_6147,N_5919,N_5674);
nand U6148 (N_6148,N_5922,N_5762);
nor U6149 (N_6149,N_5250,N_5953);
or U6150 (N_6150,N_5479,N_5036);
xor U6151 (N_6151,N_5033,N_5043);
nand U6152 (N_6152,N_5095,N_5998);
nand U6153 (N_6153,N_5252,N_5597);
and U6154 (N_6154,N_5066,N_5443);
nand U6155 (N_6155,N_5094,N_5291);
xor U6156 (N_6156,N_5595,N_5426);
nand U6157 (N_6157,N_5741,N_5017);
nand U6158 (N_6158,N_5654,N_5611);
xnor U6159 (N_6159,N_5929,N_5147);
xor U6160 (N_6160,N_5691,N_5421);
and U6161 (N_6161,N_5403,N_5193);
nor U6162 (N_6162,N_5225,N_5444);
and U6163 (N_6163,N_5649,N_5232);
and U6164 (N_6164,N_5652,N_5783);
xnor U6165 (N_6165,N_5826,N_5169);
or U6166 (N_6166,N_5114,N_5320);
nand U6167 (N_6167,N_5511,N_5186);
and U6168 (N_6168,N_5116,N_5319);
nor U6169 (N_6169,N_5653,N_5780);
or U6170 (N_6170,N_5628,N_5432);
xor U6171 (N_6171,N_5898,N_5749);
and U6172 (N_6172,N_5339,N_5701);
and U6173 (N_6173,N_5011,N_5156);
and U6174 (N_6174,N_5202,N_5324);
and U6175 (N_6175,N_5400,N_5675);
nor U6176 (N_6176,N_5129,N_5090);
nand U6177 (N_6177,N_5848,N_5361);
or U6178 (N_6178,N_5822,N_5397);
and U6179 (N_6179,N_5534,N_5005);
and U6180 (N_6180,N_5884,N_5693);
or U6181 (N_6181,N_5620,N_5335);
nand U6182 (N_6182,N_5845,N_5224);
nand U6183 (N_6183,N_5788,N_5886);
xnor U6184 (N_6184,N_5292,N_5333);
nand U6185 (N_6185,N_5041,N_5082);
nor U6186 (N_6186,N_5296,N_5895);
nand U6187 (N_6187,N_5531,N_5683);
nand U6188 (N_6188,N_5495,N_5600);
nor U6189 (N_6189,N_5547,N_5768);
nand U6190 (N_6190,N_5380,N_5109);
nor U6191 (N_6191,N_5466,N_5265);
or U6192 (N_6192,N_5091,N_5330);
or U6193 (N_6193,N_5542,N_5709);
xnor U6194 (N_6194,N_5211,N_5074);
and U6195 (N_6195,N_5032,N_5995);
nand U6196 (N_6196,N_5223,N_5487);
nand U6197 (N_6197,N_5028,N_5217);
nand U6198 (N_6198,N_5085,N_5243);
xor U6199 (N_6199,N_5765,N_5564);
or U6200 (N_6200,N_5325,N_5229);
xnor U6201 (N_6201,N_5584,N_5124);
xor U6202 (N_6202,N_5565,N_5062);
and U6203 (N_6203,N_5920,N_5199);
and U6204 (N_6204,N_5944,N_5295);
and U6205 (N_6205,N_5351,N_5257);
xor U6206 (N_6206,N_5151,N_5203);
nand U6207 (N_6207,N_5278,N_5288);
xnor U6208 (N_6208,N_5249,N_5606);
nand U6209 (N_6209,N_5130,N_5004);
nor U6210 (N_6210,N_5300,N_5710);
or U6211 (N_6211,N_5118,N_5594);
or U6212 (N_6212,N_5681,N_5573);
nor U6213 (N_6213,N_5744,N_5590);
and U6214 (N_6214,N_5019,N_5827);
and U6215 (N_6215,N_5857,N_5834);
xnor U6216 (N_6216,N_5891,N_5579);
nor U6217 (N_6217,N_5025,N_5692);
nand U6218 (N_6218,N_5121,N_5931);
and U6219 (N_6219,N_5306,N_5058);
xor U6220 (N_6220,N_5951,N_5808);
xor U6221 (N_6221,N_5746,N_5673);
and U6222 (N_6222,N_5809,N_5163);
xnor U6223 (N_6223,N_5038,N_5509);
nor U6224 (N_6224,N_5478,N_5658);
nor U6225 (N_6225,N_5568,N_5730);
xnor U6226 (N_6226,N_5470,N_5231);
nor U6227 (N_6227,N_5318,N_5601);
or U6228 (N_6228,N_5610,N_5964);
and U6229 (N_6229,N_5135,N_5077);
or U6230 (N_6230,N_5963,N_5974);
or U6231 (N_6231,N_5504,N_5639);
or U6232 (N_6232,N_5738,N_5759);
nand U6233 (N_6233,N_5795,N_5073);
xor U6234 (N_6234,N_5422,N_5609);
nor U6235 (N_6235,N_5773,N_5864);
xor U6236 (N_6236,N_5589,N_5555);
and U6237 (N_6237,N_5520,N_5275);
or U6238 (N_6238,N_5127,N_5616);
nor U6239 (N_6239,N_5605,N_5725);
and U6240 (N_6240,N_5668,N_5515);
nand U6241 (N_6241,N_5254,N_5614);
xnor U6242 (N_6242,N_5896,N_5401);
or U6243 (N_6243,N_5866,N_5438);
or U6244 (N_6244,N_5458,N_5802);
or U6245 (N_6245,N_5941,N_5190);
nand U6246 (N_6246,N_5930,N_5987);
or U6247 (N_6247,N_5218,N_5836);
xor U6248 (N_6248,N_5063,N_5483);
nand U6249 (N_6249,N_5950,N_5469);
nor U6250 (N_6250,N_5539,N_5806);
or U6251 (N_6251,N_5587,N_5285);
xor U6252 (N_6252,N_5684,N_5892);
and U6253 (N_6253,N_5341,N_5856);
xnor U6254 (N_6254,N_5536,N_5835);
or U6255 (N_6255,N_5618,N_5302);
xor U6256 (N_6256,N_5394,N_5800);
nand U6257 (N_6257,N_5259,N_5409);
and U6258 (N_6258,N_5546,N_5820);
and U6259 (N_6259,N_5859,N_5978);
nor U6260 (N_6260,N_5707,N_5192);
or U6261 (N_6261,N_5446,N_5697);
and U6262 (N_6262,N_5700,N_5591);
and U6263 (N_6263,N_5867,N_5336);
xor U6264 (N_6264,N_5726,N_5607);
and U6265 (N_6265,N_5290,N_5172);
and U6266 (N_6266,N_5364,N_5983);
nor U6267 (N_6267,N_5100,N_5560);
or U6268 (N_6268,N_5386,N_5279);
xor U6269 (N_6269,N_5791,N_5957);
xor U6270 (N_6270,N_5662,N_5044);
and U6271 (N_6271,N_5465,N_5794);
xnor U6272 (N_6272,N_5742,N_5260);
xor U6273 (N_6273,N_5824,N_5261);
nand U6274 (N_6274,N_5499,N_5818);
or U6275 (N_6275,N_5905,N_5840);
and U6276 (N_6276,N_5661,N_5814);
nand U6277 (N_6277,N_5311,N_5185);
nor U6278 (N_6278,N_5384,N_5076);
or U6279 (N_6279,N_5830,N_5181);
nor U6280 (N_6280,N_5474,N_5482);
xnor U6281 (N_6281,N_5708,N_5441);
nor U6282 (N_6282,N_5355,N_5092);
and U6283 (N_6283,N_5870,N_5454);
or U6284 (N_6284,N_5450,N_5334);
nand U6285 (N_6285,N_5567,N_5576);
or U6286 (N_6286,N_5695,N_5775);
and U6287 (N_6287,N_5040,N_5305);
xor U6288 (N_6288,N_5149,N_5347);
or U6289 (N_6289,N_5664,N_5110);
xor U6290 (N_6290,N_5885,N_5803);
nor U6291 (N_6291,N_5408,N_5020);
and U6292 (N_6292,N_5215,N_5256);
and U6293 (N_6293,N_5376,N_5621);
xor U6294 (N_6294,N_5390,N_5753);
xnor U6295 (N_6295,N_5863,N_5665);
or U6296 (N_6296,N_5206,N_5904);
nand U6297 (N_6297,N_5514,N_5646);
xnor U6298 (N_6298,N_5208,N_5769);
and U6299 (N_6299,N_5307,N_5578);
nor U6300 (N_6300,N_5728,N_5122);
nor U6301 (N_6301,N_5293,N_5704);
and U6302 (N_6302,N_5140,N_5563);
or U6303 (N_6303,N_5222,N_5739);
xnor U6304 (N_6304,N_5706,N_5102);
and U6305 (N_6305,N_5182,N_5851);
nor U6306 (N_6306,N_5237,N_5282);
and U6307 (N_6307,N_5023,N_5433);
and U6308 (N_6308,N_5965,N_5894);
or U6309 (N_6309,N_5298,N_5049);
and U6310 (N_6310,N_5736,N_5492);
or U6311 (N_6311,N_5997,N_5940);
and U6312 (N_6312,N_5916,N_5881);
xnor U6313 (N_6313,N_5523,N_5372);
nand U6314 (N_6314,N_5569,N_5120);
nor U6315 (N_6315,N_5529,N_5727);
or U6316 (N_6316,N_5532,N_5317);
xnor U6317 (N_6317,N_5677,N_5754);
and U6318 (N_6318,N_5526,N_5849);
xnor U6319 (N_6319,N_5924,N_5843);
xnor U6320 (N_6320,N_5046,N_5272);
nor U6321 (N_6321,N_5047,N_5910);
nor U6322 (N_6322,N_5431,N_5942);
xnor U6323 (N_6323,N_5266,N_5503);
nand U6324 (N_6324,N_5304,N_5946);
xnor U6325 (N_6325,N_5491,N_5345);
and U6326 (N_6326,N_5037,N_5475);
or U6327 (N_6327,N_5021,N_5718);
and U6328 (N_6328,N_5939,N_5134);
nor U6329 (N_6329,N_5687,N_5406);
and U6330 (N_6330,N_5696,N_5461);
nand U6331 (N_6331,N_5026,N_5638);
nand U6332 (N_6332,N_5540,N_5423);
xnor U6333 (N_6333,N_5713,N_5751);
nand U6334 (N_6334,N_5932,N_5173);
nor U6335 (N_6335,N_5918,N_5233);
xor U6336 (N_6336,N_5138,N_5799);
nor U6337 (N_6337,N_5093,N_5842);
xnor U6338 (N_6338,N_5016,N_5570);
or U6339 (N_6339,N_5952,N_5533);
nand U6340 (N_6340,N_5352,N_5853);
nand U6341 (N_6341,N_5750,N_5111);
and U6342 (N_6342,N_5680,N_5006);
xor U6343 (N_6343,N_5968,N_5132);
nor U6344 (N_6344,N_5350,N_5060);
xnor U6345 (N_6345,N_5262,N_5013);
or U6346 (N_6346,N_5644,N_5508);
nand U6347 (N_6347,N_5785,N_5634);
or U6348 (N_6348,N_5624,N_5786);
and U6349 (N_6349,N_5764,N_5195);
nor U6350 (N_6350,N_5585,N_5489);
xnor U6351 (N_6351,N_5269,N_5703);
xnor U6352 (N_6352,N_5053,N_5556);
nor U6353 (N_6353,N_5369,N_5194);
nand U6354 (N_6354,N_5081,N_5381);
nand U6355 (N_6355,N_5770,N_5906);
nor U6356 (N_6356,N_5926,N_5117);
nor U6357 (N_6357,N_5378,N_5771);
or U6358 (N_6358,N_5108,N_5498);
nand U6359 (N_6359,N_5370,N_5629);
nand U6360 (N_6360,N_5286,N_5747);
nand U6361 (N_6361,N_5844,N_5165);
or U6362 (N_6362,N_5876,N_5559);
or U6363 (N_6363,N_5405,N_5577);
nand U6364 (N_6364,N_5061,N_5733);
and U6365 (N_6365,N_5497,N_5142);
or U6366 (N_6366,N_5656,N_5724);
or U6367 (N_6367,N_5273,N_5420);
and U6368 (N_6368,N_5490,N_5812);
xor U6369 (N_6369,N_5358,N_5383);
nand U6370 (N_6370,N_5535,N_5280);
xor U6371 (N_6371,N_5580,N_5583);
and U6372 (N_6372,N_5694,N_5582);
nor U6373 (N_6373,N_5501,N_5457);
and U6374 (N_6374,N_5128,N_5071);
and U6375 (N_6375,N_5164,N_5105);
nand U6376 (N_6376,N_5137,N_5054);
nand U6377 (N_6377,N_5065,N_5271);
nor U6378 (N_6378,N_5052,N_5227);
and U6379 (N_6379,N_5238,N_5528);
or U6380 (N_6380,N_5221,N_5797);
nand U6381 (N_6381,N_5270,N_5817);
nand U6382 (N_6382,N_5938,N_5009);
xor U6383 (N_6383,N_5715,N_5852);
nand U6384 (N_6384,N_5912,N_5346);
nor U6385 (N_6385,N_5991,N_5463);
xnor U6386 (N_6386,N_5230,N_5332);
and U6387 (N_6387,N_5737,N_5236);
or U6388 (N_6388,N_5360,N_5174);
or U6389 (N_6389,N_5242,N_5402);
nand U6390 (N_6390,N_5359,N_5115);
nor U6391 (N_6391,N_5434,N_5168);
and U6392 (N_6392,N_5722,N_5196);
nand U6393 (N_6393,N_5452,N_5603);
and U6394 (N_6394,N_5615,N_5561);
nor U6395 (N_6395,N_5519,N_5660);
and U6396 (N_6396,N_5850,N_5103);
nor U6397 (N_6397,N_5075,N_5748);
nand U6398 (N_6398,N_5464,N_5612);
nor U6399 (N_6399,N_5903,N_5552);
nand U6400 (N_6400,N_5171,N_5449);
nand U6401 (N_6401,N_5411,N_5588);
nand U6402 (N_6402,N_5807,N_5619);
xnor U6403 (N_6403,N_5099,N_5811);
or U6404 (N_6404,N_5679,N_5959);
nand U6405 (N_6405,N_5213,N_5471);
nand U6406 (N_6406,N_5825,N_5981);
or U6407 (N_6407,N_5057,N_5209);
nor U6408 (N_6408,N_5967,N_5414);
nand U6409 (N_6409,N_5170,N_5042);
nand U6410 (N_6410,N_5636,N_5893);
or U6411 (N_6411,N_5855,N_5160);
or U6412 (N_6412,N_5507,N_5545);
nor U6413 (N_6413,N_5982,N_5035);
nor U6414 (N_6414,N_5525,N_5883);
xor U6415 (N_6415,N_5451,N_5437);
and U6416 (N_6416,N_5711,N_5549);
and U6417 (N_6417,N_5200,N_5007);
or U6418 (N_6418,N_5933,N_5456);
or U6419 (N_6419,N_5617,N_5666);
nor U6420 (N_6420,N_5106,N_5083);
xor U6421 (N_6421,N_5029,N_5650);
nand U6422 (N_6422,N_5937,N_5860);
and U6423 (N_6423,N_5371,N_5574);
or U6424 (N_6424,N_5986,N_5363);
xor U6425 (N_6425,N_5973,N_5837);
nand U6426 (N_6426,N_5516,N_5159);
nor U6427 (N_6427,N_5596,N_5349);
nor U6428 (N_6428,N_5136,N_5505);
and U6429 (N_6429,N_5488,N_5476);
or U6430 (N_6430,N_5240,N_5374);
nand U6431 (N_6431,N_5988,N_5779);
or U6432 (N_6432,N_5078,N_5027);
and U6433 (N_6433,N_5460,N_5048);
nor U6434 (N_6434,N_5144,N_5731);
xor U6435 (N_6435,N_5008,N_5682);
or U6436 (N_6436,N_5473,N_5418);
nand U6437 (N_6437,N_5586,N_5287);
nor U6438 (N_6438,N_5875,N_5676);
or U6439 (N_6439,N_5557,N_5714);
or U6440 (N_6440,N_5326,N_5404);
or U6441 (N_6441,N_5913,N_5763);
or U6442 (N_6442,N_5999,N_5150);
and U6443 (N_6443,N_5734,N_5518);
and U6444 (N_6444,N_5158,N_5623);
nand U6445 (N_6445,N_5954,N_5805);
or U6446 (N_6446,N_5659,N_5308);
nand U6447 (N_6447,N_5018,N_5774);
and U6448 (N_6448,N_5921,N_5356);
nor U6449 (N_6449,N_5328,N_5034);
or U6450 (N_6450,N_5440,N_5396);
or U6451 (N_6451,N_5669,N_5387);
nor U6452 (N_6452,N_5080,N_5201);
xnor U6453 (N_6453,N_5012,N_5980);
and U6454 (N_6454,N_5887,N_5084);
or U6455 (N_6455,N_5874,N_5247);
and U6456 (N_6456,N_5527,N_5493);
and U6457 (N_6457,N_5989,N_5956);
nor U6458 (N_6458,N_5958,N_5671);
xnor U6459 (N_6459,N_5592,N_5331);
xnor U6460 (N_6460,N_5353,N_5598);
or U6461 (N_6461,N_5548,N_5126);
or U6462 (N_6462,N_5571,N_5670);
or U6463 (N_6463,N_5992,N_5289);
and U6464 (N_6464,N_5633,N_5971);
xor U6465 (N_6465,N_5391,N_5553);
and U6466 (N_6466,N_5191,N_5435);
or U6467 (N_6467,N_5593,N_5143);
nor U6468 (N_6468,N_5365,N_5284);
or U6469 (N_6469,N_5663,N_5784);
or U6470 (N_6470,N_5398,N_5480);
nand U6471 (N_6471,N_5635,N_5757);
nor U6472 (N_6472,N_5796,N_5139);
xor U6473 (N_6473,N_5521,N_5467);
or U6474 (N_6474,N_5216,N_5146);
nand U6475 (N_6475,N_5294,N_5145);
nand U6476 (N_6476,N_5961,N_5723);
nand U6477 (N_6477,N_5392,N_5970);
or U6478 (N_6478,N_5873,N_5448);
nor U6479 (N_6479,N_5752,N_5263);
and U6480 (N_6480,N_5188,N_5419);
xor U6481 (N_6481,N_5316,N_5003);
nand U6482 (N_6482,N_5354,N_5627);
xor U6483 (N_6483,N_5756,N_5790);
nand U6484 (N_6484,N_5321,N_5758);
nor U6485 (N_6485,N_5943,N_5366);
or U6486 (N_6486,N_5210,N_5157);
xor U6487 (N_6487,N_5481,N_5204);
or U6488 (N_6488,N_5562,N_5367);
xnor U6489 (N_6489,N_5721,N_5688);
xor U6490 (N_6490,N_5994,N_5642);
nand U6491 (N_6491,N_5348,N_5251);
nand U6492 (N_6492,N_5395,N_5740);
or U6493 (N_6493,N_5554,N_5059);
nor U6494 (N_6494,N_5477,N_5323);
nor U6495 (N_6495,N_5069,N_5550);
xor U6496 (N_6496,N_5056,N_5705);
nor U6497 (N_6497,N_5829,N_5625);
and U6498 (N_6498,N_5051,N_5833);
xor U6499 (N_6499,N_5101,N_5960);
nor U6500 (N_6500,N_5243,N_5436);
or U6501 (N_6501,N_5993,N_5515);
and U6502 (N_6502,N_5229,N_5285);
nand U6503 (N_6503,N_5205,N_5268);
xor U6504 (N_6504,N_5573,N_5175);
nand U6505 (N_6505,N_5078,N_5373);
or U6506 (N_6506,N_5302,N_5167);
xnor U6507 (N_6507,N_5476,N_5157);
xnor U6508 (N_6508,N_5786,N_5773);
nand U6509 (N_6509,N_5487,N_5989);
nor U6510 (N_6510,N_5661,N_5650);
and U6511 (N_6511,N_5616,N_5609);
or U6512 (N_6512,N_5008,N_5859);
or U6513 (N_6513,N_5130,N_5502);
or U6514 (N_6514,N_5697,N_5369);
nand U6515 (N_6515,N_5898,N_5527);
and U6516 (N_6516,N_5207,N_5187);
or U6517 (N_6517,N_5232,N_5472);
or U6518 (N_6518,N_5402,N_5796);
xor U6519 (N_6519,N_5827,N_5157);
nor U6520 (N_6520,N_5130,N_5414);
or U6521 (N_6521,N_5989,N_5160);
nor U6522 (N_6522,N_5352,N_5959);
and U6523 (N_6523,N_5727,N_5687);
or U6524 (N_6524,N_5833,N_5519);
nor U6525 (N_6525,N_5726,N_5047);
or U6526 (N_6526,N_5786,N_5460);
or U6527 (N_6527,N_5489,N_5713);
nor U6528 (N_6528,N_5050,N_5991);
and U6529 (N_6529,N_5361,N_5890);
or U6530 (N_6530,N_5568,N_5455);
or U6531 (N_6531,N_5769,N_5114);
xor U6532 (N_6532,N_5293,N_5686);
and U6533 (N_6533,N_5065,N_5610);
and U6534 (N_6534,N_5383,N_5626);
nor U6535 (N_6535,N_5169,N_5537);
nor U6536 (N_6536,N_5299,N_5405);
and U6537 (N_6537,N_5848,N_5298);
or U6538 (N_6538,N_5813,N_5919);
xor U6539 (N_6539,N_5522,N_5496);
nand U6540 (N_6540,N_5659,N_5778);
nand U6541 (N_6541,N_5292,N_5294);
and U6542 (N_6542,N_5353,N_5344);
nor U6543 (N_6543,N_5799,N_5196);
nor U6544 (N_6544,N_5752,N_5350);
nor U6545 (N_6545,N_5118,N_5861);
nor U6546 (N_6546,N_5959,N_5626);
nand U6547 (N_6547,N_5251,N_5062);
and U6548 (N_6548,N_5192,N_5062);
xor U6549 (N_6549,N_5700,N_5680);
xor U6550 (N_6550,N_5078,N_5872);
nor U6551 (N_6551,N_5810,N_5745);
nand U6552 (N_6552,N_5298,N_5598);
xor U6553 (N_6553,N_5746,N_5920);
and U6554 (N_6554,N_5375,N_5916);
xor U6555 (N_6555,N_5797,N_5612);
and U6556 (N_6556,N_5934,N_5118);
and U6557 (N_6557,N_5524,N_5412);
nand U6558 (N_6558,N_5581,N_5750);
and U6559 (N_6559,N_5755,N_5256);
nor U6560 (N_6560,N_5279,N_5907);
or U6561 (N_6561,N_5437,N_5610);
nand U6562 (N_6562,N_5533,N_5780);
and U6563 (N_6563,N_5905,N_5700);
or U6564 (N_6564,N_5860,N_5870);
and U6565 (N_6565,N_5880,N_5576);
and U6566 (N_6566,N_5040,N_5093);
xnor U6567 (N_6567,N_5038,N_5991);
nor U6568 (N_6568,N_5324,N_5258);
nand U6569 (N_6569,N_5067,N_5324);
nor U6570 (N_6570,N_5343,N_5318);
and U6571 (N_6571,N_5624,N_5968);
nand U6572 (N_6572,N_5223,N_5128);
nor U6573 (N_6573,N_5045,N_5188);
or U6574 (N_6574,N_5290,N_5352);
nor U6575 (N_6575,N_5862,N_5703);
nand U6576 (N_6576,N_5230,N_5808);
xnor U6577 (N_6577,N_5839,N_5604);
nor U6578 (N_6578,N_5402,N_5653);
or U6579 (N_6579,N_5378,N_5118);
xnor U6580 (N_6580,N_5543,N_5018);
xnor U6581 (N_6581,N_5051,N_5986);
xor U6582 (N_6582,N_5788,N_5378);
nand U6583 (N_6583,N_5562,N_5385);
nand U6584 (N_6584,N_5835,N_5813);
and U6585 (N_6585,N_5571,N_5860);
xor U6586 (N_6586,N_5136,N_5190);
nand U6587 (N_6587,N_5210,N_5320);
xnor U6588 (N_6588,N_5911,N_5424);
nor U6589 (N_6589,N_5589,N_5362);
nand U6590 (N_6590,N_5722,N_5530);
xnor U6591 (N_6591,N_5744,N_5166);
nand U6592 (N_6592,N_5004,N_5512);
and U6593 (N_6593,N_5856,N_5499);
and U6594 (N_6594,N_5453,N_5417);
xor U6595 (N_6595,N_5366,N_5756);
nor U6596 (N_6596,N_5786,N_5915);
or U6597 (N_6597,N_5976,N_5750);
or U6598 (N_6598,N_5927,N_5806);
xnor U6599 (N_6599,N_5844,N_5365);
xnor U6600 (N_6600,N_5188,N_5096);
xnor U6601 (N_6601,N_5839,N_5883);
or U6602 (N_6602,N_5729,N_5146);
and U6603 (N_6603,N_5175,N_5174);
and U6604 (N_6604,N_5266,N_5375);
nor U6605 (N_6605,N_5313,N_5393);
or U6606 (N_6606,N_5638,N_5649);
and U6607 (N_6607,N_5729,N_5434);
nor U6608 (N_6608,N_5726,N_5738);
xnor U6609 (N_6609,N_5924,N_5650);
xor U6610 (N_6610,N_5404,N_5130);
or U6611 (N_6611,N_5417,N_5105);
and U6612 (N_6612,N_5963,N_5069);
nand U6613 (N_6613,N_5885,N_5849);
and U6614 (N_6614,N_5292,N_5417);
nand U6615 (N_6615,N_5081,N_5958);
nor U6616 (N_6616,N_5115,N_5832);
nand U6617 (N_6617,N_5056,N_5159);
and U6618 (N_6618,N_5496,N_5289);
nor U6619 (N_6619,N_5872,N_5450);
nand U6620 (N_6620,N_5470,N_5882);
nand U6621 (N_6621,N_5509,N_5631);
nand U6622 (N_6622,N_5855,N_5841);
nor U6623 (N_6623,N_5694,N_5745);
or U6624 (N_6624,N_5883,N_5603);
and U6625 (N_6625,N_5961,N_5375);
or U6626 (N_6626,N_5152,N_5970);
and U6627 (N_6627,N_5737,N_5715);
nand U6628 (N_6628,N_5836,N_5308);
nor U6629 (N_6629,N_5265,N_5874);
and U6630 (N_6630,N_5009,N_5652);
nor U6631 (N_6631,N_5878,N_5760);
nor U6632 (N_6632,N_5353,N_5911);
xnor U6633 (N_6633,N_5321,N_5124);
nand U6634 (N_6634,N_5175,N_5364);
and U6635 (N_6635,N_5295,N_5112);
xor U6636 (N_6636,N_5745,N_5665);
and U6637 (N_6637,N_5468,N_5829);
nor U6638 (N_6638,N_5118,N_5583);
or U6639 (N_6639,N_5917,N_5643);
xor U6640 (N_6640,N_5570,N_5322);
xnor U6641 (N_6641,N_5724,N_5695);
or U6642 (N_6642,N_5016,N_5685);
xor U6643 (N_6643,N_5606,N_5512);
or U6644 (N_6644,N_5331,N_5859);
or U6645 (N_6645,N_5265,N_5675);
nor U6646 (N_6646,N_5548,N_5328);
nor U6647 (N_6647,N_5131,N_5597);
or U6648 (N_6648,N_5135,N_5581);
or U6649 (N_6649,N_5717,N_5033);
and U6650 (N_6650,N_5812,N_5777);
nand U6651 (N_6651,N_5393,N_5845);
xor U6652 (N_6652,N_5353,N_5959);
and U6653 (N_6653,N_5536,N_5733);
xor U6654 (N_6654,N_5488,N_5774);
or U6655 (N_6655,N_5397,N_5350);
xnor U6656 (N_6656,N_5541,N_5038);
or U6657 (N_6657,N_5590,N_5185);
nand U6658 (N_6658,N_5005,N_5720);
and U6659 (N_6659,N_5150,N_5334);
nand U6660 (N_6660,N_5077,N_5503);
nand U6661 (N_6661,N_5990,N_5935);
and U6662 (N_6662,N_5024,N_5874);
or U6663 (N_6663,N_5408,N_5386);
and U6664 (N_6664,N_5499,N_5855);
or U6665 (N_6665,N_5664,N_5659);
xnor U6666 (N_6666,N_5880,N_5437);
xor U6667 (N_6667,N_5092,N_5772);
or U6668 (N_6668,N_5935,N_5932);
nor U6669 (N_6669,N_5372,N_5844);
or U6670 (N_6670,N_5654,N_5518);
nor U6671 (N_6671,N_5618,N_5805);
xor U6672 (N_6672,N_5929,N_5057);
xnor U6673 (N_6673,N_5948,N_5087);
nor U6674 (N_6674,N_5416,N_5338);
and U6675 (N_6675,N_5879,N_5372);
xor U6676 (N_6676,N_5940,N_5305);
and U6677 (N_6677,N_5206,N_5055);
and U6678 (N_6678,N_5654,N_5849);
xor U6679 (N_6679,N_5964,N_5144);
and U6680 (N_6680,N_5236,N_5477);
nand U6681 (N_6681,N_5658,N_5975);
nand U6682 (N_6682,N_5822,N_5633);
and U6683 (N_6683,N_5707,N_5920);
or U6684 (N_6684,N_5276,N_5816);
or U6685 (N_6685,N_5268,N_5348);
xor U6686 (N_6686,N_5173,N_5345);
and U6687 (N_6687,N_5418,N_5253);
or U6688 (N_6688,N_5681,N_5164);
xor U6689 (N_6689,N_5001,N_5548);
xor U6690 (N_6690,N_5116,N_5350);
or U6691 (N_6691,N_5841,N_5676);
and U6692 (N_6692,N_5814,N_5430);
nand U6693 (N_6693,N_5073,N_5733);
xor U6694 (N_6694,N_5373,N_5003);
nand U6695 (N_6695,N_5830,N_5679);
or U6696 (N_6696,N_5745,N_5926);
or U6697 (N_6697,N_5497,N_5923);
nor U6698 (N_6698,N_5507,N_5625);
nor U6699 (N_6699,N_5348,N_5755);
nand U6700 (N_6700,N_5944,N_5215);
nand U6701 (N_6701,N_5291,N_5477);
nand U6702 (N_6702,N_5609,N_5603);
xor U6703 (N_6703,N_5385,N_5739);
or U6704 (N_6704,N_5346,N_5249);
xnor U6705 (N_6705,N_5654,N_5432);
xor U6706 (N_6706,N_5664,N_5937);
or U6707 (N_6707,N_5204,N_5596);
or U6708 (N_6708,N_5628,N_5370);
nand U6709 (N_6709,N_5454,N_5902);
nand U6710 (N_6710,N_5637,N_5007);
xor U6711 (N_6711,N_5752,N_5216);
xnor U6712 (N_6712,N_5032,N_5540);
xor U6713 (N_6713,N_5530,N_5470);
nand U6714 (N_6714,N_5439,N_5310);
and U6715 (N_6715,N_5671,N_5389);
nor U6716 (N_6716,N_5487,N_5736);
or U6717 (N_6717,N_5192,N_5957);
nand U6718 (N_6718,N_5256,N_5728);
or U6719 (N_6719,N_5832,N_5084);
xnor U6720 (N_6720,N_5157,N_5361);
xor U6721 (N_6721,N_5478,N_5992);
and U6722 (N_6722,N_5354,N_5456);
nor U6723 (N_6723,N_5141,N_5236);
and U6724 (N_6724,N_5605,N_5295);
and U6725 (N_6725,N_5106,N_5014);
or U6726 (N_6726,N_5147,N_5992);
xor U6727 (N_6727,N_5762,N_5410);
nor U6728 (N_6728,N_5021,N_5161);
and U6729 (N_6729,N_5957,N_5439);
xnor U6730 (N_6730,N_5205,N_5301);
nor U6731 (N_6731,N_5591,N_5761);
xnor U6732 (N_6732,N_5421,N_5837);
xor U6733 (N_6733,N_5978,N_5408);
or U6734 (N_6734,N_5062,N_5884);
nor U6735 (N_6735,N_5097,N_5131);
or U6736 (N_6736,N_5998,N_5973);
nand U6737 (N_6737,N_5781,N_5327);
or U6738 (N_6738,N_5579,N_5147);
and U6739 (N_6739,N_5385,N_5654);
nand U6740 (N_6740,N_5078,N_5891);
nor U6741 (N_6741,N_5286,N_5047);
nand U6742 (N_6742,N_5516,N_5374);
nand U6743 (N_6743,N_5392,N_5372);
and U6744 (N_6744,N_5127,N_5467);
xor U6745 (N_6745,N_5283,N_5878);
or U6746 (N_6746,N_5190,N_5057);
and U6747 (N_6747,N_5842,N_5646);
or U6748 (N_6748,N_5933,N_5044);
and U6749 (N_6749,N_5077,N_5228);
xor U6750 (N_6750,N_5972,N_5844);
or U6751 (N_6751,N_5689,N_5075);
nand U6752 (N_6752,N_5677,N_5081);
or U6753 (N_6753,N_5738,N_5454);
nand U6754 (N_6754,N_5068,N_5164);
nor U6755 (N_6755,N_5301,N_5743);
and U6756 (N_6756,N_5803,N_5156);
nor U6757 (N_6757,N_5134,N_5334);
nor U6758 (N_6758,N_5469,N_5650);
xnor U6759 (N_6759,N_5999,N_5315);
nor U6760 (N_6760,N_5533,N_5402);
xor U6761 (N_6761,N_5269,N_5071);
nand U6762 (N_6762,N_5406,N_5828);
xnor U6763 (N_6763,N_5165,N_5829);
nor U6764 (N_6764,N_5410,N_5101);
and U6765 (N_6765,N_5233,N_5577);
nor U6766 (N_6766,N_5244,N_5266);
and U6767 (N_6767,N_5611,N_5363);
and U6768 (N_6768,N_5492,N_5036);
nand U6769 (N_6769,N_5390,N_5125);
nor U6770 (N_6770,N_5753,N_5810);
nor U6771 (N_6771,N_5613,N_5376);
or U6772 (N_6772,N_5050,N_5332);
xnor U6773 (N_6773,N_5009,N_5532);
or U6774 (N_6774,N_5787,N_5362);
or U6775 (N_6775,N_5861,N_5310);
nor U6776 (N_6776,N_5158,N_5696);
xnor U6777 (N_6777,N_5258,N_5081);
nor U6778 (N_6778,N_5423,N_5545);
or U6779 (N_6779,N_5503,N_5991);
and U6780 (N_6780,N_5127,N_5841);
or U6781 (N_6781,N_5308,N_5145);
or U6782 (N_6782,N_5848,N_5868);
and U6783 (N_6783,N_5767,N_5827);
or U6784 (N_6784,N_5150,N_5111);
and U6785 (N_6785,N_5139,N_5330);
nand U6786 (N_6786,N_5909,N_5451);
and U6787 (N_6787,N_5205,N_5682);
or U6788 (N_6788,N_5102,N_5332);
xnor U6789 (N_6789,N_5397,N_5352);
nor U6790 (N_6790,N_5973,N_5957);
xor U6791 (N_6791,N_5501,N_5247);
nor U6792 (N_6792,N_5077,N_5410);
xor U6793 (N_6793,N_5798,N_5137);
and U6794 (N_6794,N_5031,N_5967);
and U6795 (N_6795,N_5018,N_5531);
or U6796 (N_6796,N_5704,N_5897);
xor U6797 (N_6797,N_5804,N_5519);
nand U6798 (N_6798,N_5497,N_5749);
nand U6799 (N_6799,N_5757,N_5320);
nand U6800 (N_6800,N_5015,N_5441);
or U6801 (N_6801,N_5571,N_5431);
and U6802 (N_6802,N_5514,N_5394);
xor U6803 (N_6803,N_5046,N_5224);
nor U6804 (N_6804,N_5811,N_5269);
or U6805 (N_6805,N_5521,N_5519);
and U6806 (N_6806,N_5222,N_5241);
xor U6807 (N_6807,N_5387,N_5218);
or U6808 (N_6808,N_5053,N_5101);
nand U6809 (N_6809,N_5451,N_5175);
nor U6810 (N_6810,N_5766,N_5400);
nand U6811 (N_6811,N_5774,N_5625);
nand U6812 (N_6812,N_5038,N_5740);
and U6813 (N_6813,N_5783,N_5999);
nor U6814 (N_6814,N_5443,N_5159);
or U6815 (N_6815,N_5847,N_5472);
xor U6816 (N_6816,N_5222,N_5421);
and U6817 (N_6817,N_5702,N_5339);
and U6818 (N_6818,N_5197,N_5033);
and U6819 (N_6819,N_5715,N_5900);
nor U6820 (N_6820,N_5036,N_5987);
or U6821 (N_6821,N_5485,N_5158);
or U6822 (N_6822,N_5026,N_5305);
nand U6823 (N_6823,N_5969,N_5936);
or U6824 (N_6824,N_5336,N_5373);
nor U6825 (N_6825,N_5347,N_5718);
and U6826 (N_6826,N_5560,N_5433);
nor U6827 (N_6827,N_5580,N_5466);
xor U6828 (N_6828,N_5942,N_5809);
or U6829 (N_6829,N_5682,N_5801);
nand U6830 (N_6830,N_5736,N_5090);
or U6831 (N_6831,N_5703,N_5825);
or U6832 (N_6832,N_5005,N_5258);
nand U6833 (N_6833,N_5357,N_5602);
xnor U6834 (N_6834,N_5747,N_5362);
and U6835 (N_6835,N_5794,N_5668);
and U6836 (N_6836,N_5903,N_5224);
and U6837 (N_6837,N_5702,N_5022);
xnor U6838 (N_6838,N_5720,N_5570);
and U6839 (N_6839,N_5416,N_5779);
nand U6840 (N_6840,N_5988,N_5220);
or U6841 (N_6841,N_5862,N_5804);
nand U6842 (N_6842,N_5271,N_5563);
xor U6843 (N_6843,N_5167,N_5200);
and U6844 (N_6844,N_5468,N_5836);
and U6845 (N_6845,N_5062,N_5790);
or U6846 (N_6846,N_5888,N_5950);
nor U6847 (N_6847,N_5825,N_5008);
nand U6848 (N_6848,N_5172,N_5857);
nand U6849 (N_6849,N_5049,N_5263);
and U6850 (N_6850,N_5709,N_5950);
or U6851 (N_6851,N_5958,N_5660);
nand U6852 (N_6852,N_5007,N_5010);
xnor U6853 (N_6853,N_5538,N_5999);
or U6854 (N_6854,N_5524,N_5783);
nor U6855 (N_6855,N_5394,N_5759);
nor U6856 (N_6856,N_5481,N_5556);
nand U6857 (N_6857,N_5232,N_5444);
nand U6858 (N_6858,N_5186,N_5034);
xor U6859 (N_6859,N_5143,N_5688);
or U6860 (N_6860,N_5961,N_5376);
and U6861 (N_6861,N_5921,N_5945);
and U6862 (N_6862,N_5209,N_5785);
and U6863 (N_6863,N_5578,N_5182);
and U6864 (N_6864,N_5642,N_5205);
nand U6865 (N_6865,N_5584,N_5311);
or U6866 (N_6866,N_5478,N_5972);
or U6867 (N_6867,N_5607,N_5155);
or U6868 (N_6868,N_5166,N_5971);
xor U6869 (N_6869,N_5005,N_5654);
nand U6870 (N_6870,N_5461,N_5814);
xnor U6871 (N_6871,N_5843,N_5317);
nor U6872 (N_6872,N_5812,N_5775);
and U6873 (N_6873,N_5963,N_5150);
and U6874 (N_6874,N_5778,N_5883);
xnor U6875 (N_6875,N_5340,N_5329);
or U6876 (N_6876,N_5549,N_5152);
nor U6877 (N_6877,N_5800,N_5031);
and U6878 (N_6878,N_5021,N_5191);
xor U6879 (N_6879,N_5973,N_5875);
nand U6880 (N_6880,N_5443,N_5851);
nand U6881 (N_6881,N_5065,N_5703);
and U6882 (N_6882,N_5414,N_5310);
and U6883 (N_6883,N_5488,N_5171);
nor U6884 (N_6884,N_5421,N_5777);
nor U6885 (N_6885,N_5975,N_5292);
nor U6886 (N_6886,N_5331,N_5403);
or U6887 (N_6887,N_5741,N_5537);
and U6888 (N_6888,N_5935,N_5720);
xnor U6889 (N_6889,N_5713,N_5992);
or U6890 (N_6890,N_5313,N_5240);
nor U6891 (N_6891,N_5360,N_5248);
nand U6892 (N_6892,N_5243,N_5721);
nor U6893 (N_6893,N_5288,N_5051);
and U6894 (N_6894,N_5526,N_5782);
nand U6895 (N_6895,N_5243,N_5145);
nand U6896 (N_6896,N_5718,N_5956);
and U6897 (N_6897,N_5701,N_5564);
and U6898 (N_6898,N_5590,N_5836);
or U6899 (N_6899,N_5780,N_5277);
or U6900 (N_6900,N_5694,N_5497);
nor U6901 (N_6901,N_5440,N_5677);
nor U6902 (N_6902,N_5004,N_5909);
and U6903 (N_6903,N_5019,N_5748);
nand U6904 (N_6904,N_5588,N_5286);
xor U6905 (N_6905,N_5226,N_5014);
and U6906 (N_6906,N_5261,N_5591);
nor U6907 (N_6907,N_5281,N_5384);
or U6908 (N_6908,N_5062,N_5533);
nor U6909 (N_6909,N_5916,N_5001);
and U6910 (N_6910,N_5550,N_5459);
or U6911 (N_6911,N_5323,N_5250);
nor U6912 (N_6912,N_5986,N_5764);
nand U6913 (N_6913,N_5732,N_5715);
nand U6914 (N_6914,N_5913,N_5494);
nand U6915 (N_6915,N_5710,N_5234);
or U6916 (N_6916,N_5238,N_5456);
nand U6917 (N_6917,N_5145,N_5558);
or U6918 (N_6918,N_5699,N_5131);
xnor U6919 (N_6919,N_5041,N_5416);
and U6920 (N_6920,N_5107,N_5657);
or U6921 (N_6921,N_5414,N_5637);
nor U6922 (N_6922,N_5752,N_5046);
and U6923 (N_6923,N_5886,N_5512);
xnor U6924 (N_6924,N_5852,N_5220);
nor U6925 (N_6925,N_5176,N_5835);
nand U6926 (N_6926,N_5655,N_5116);
xor U6927 (N_6927,N_5851,N_5592);
nor U6928 (N_6928,N_5387,N_5326);
xnor U6929 (N_6929,N_5774,N_5947);
and U6930 (N_6930,N_5622,N_5401);
or U6931 (N_6931,N_5666,N_5798);
nand U6932 (N_6932,N_5628,N_5451);
xor U6933 (N_6933,N_5206,N_5929);
xnor U6934 (N_6934,N_5191,N_5215);
and U6935 (N_6935,N_5206,N_5663);
nor U6936 (N_6936,N_5815,N_5781);
and U6937 (N_6937,N_5703,N_5071);
nand U6938 (N_6938,N_5953,N_5132);
or U6939 (N_6939,N_5672,N_5957);
xnor U6940 (N_6940,N_5420,N_5516);
xor U6941 (N_6941,N_5763,N_5857);
nand U6942 (N_6942,N_5910,N_5418);
xor U6943 (N_6943,N_5449,N_5578);
nor U6944 (N_6944,N_5908,N_5685);
nor U6945 (N_6945,N_5897,N_5787);
and U6946 (N_6946,N_5643,N_5415);
nand U6947 (N_6947,N_5844,N_5261);
and U6948 (N_6948,N_5814,N_5785);
and U6949 (N_6949,N_5609,N_5121);
xnor U6950 (N_6950,N_5836,N_5379);
nand U6951 (N_6951,N_5042,N_5450);
and U6952 (N_6952,N_5307,N_5693);
xnor U6953 (N_6953,N_5472,N_5167);
nor U6954 (N_6954,N_5941,N_5999);
nand U6955 (N_6955,N_5237,N_5394);
or U6956 (N_6956,N_5657,N_5219);
xor U6957 (N_6957,N_5122,N_5036);
and U6958 (N_6958,N_5415,N_5206);
or U6959 (N_6959,N_5345,N_5365);
nor U6960 (N_6960,N_5634,N_5609);
nand U6961 (N_6961,N_5448,N_5845);
or U6962 (N_6962,N_5271,N_5386);
xor U6963 (N_6963,N_5644,N_5536);
nor U6964 (N_6964,N_5282,N_5170);
or U6965 (N_6965,N_5924,N_5506);
nor U6966 (N_6966,N_5159,N_5064);
xnor U6967 (N_6967,N_5695,N_5025);
xnor U6968 (N_6968,N_5347,N_5876);
or U6969 (N_6969,N_5736,N_5099);
xnor U6970 (N_6970,N_5341,N_5407);
xor U6971 (N_6971,N_5739,N_5602);
xor U6972 (N_6972,N_5193,N_5165);
or U6973 (N_6973,N_5469,N_5642);
and U6974 (N_6974,N_5229,N_5745);
xor U6975 (N_6975,N_5729,N_5207);
and U6976 (N_6976,N_5445,N_5602);
and U6977 (N_6977,N_5788,N_5120);
and U6978 (N_6978,N_5141,N_5178);
and U6979 (N_6979,N_5040,N_5460);
nor U6980 (N_6980,N_5587,N_5229);
and U6981 (N_6981,N_5925,N_5436);
or U6982 (N_6982,N_5555,N_5492);
or U6983 (N_6983,N_5217,N_5731);
and U6984 (N_6984,N_5337,N_5697);
nand U6985 (N_6985,N_5139,N_5148);
xnor U6986 (N_6986,N_5970,N_5257);
nor U6987 (N_6987,N_5787,N_5791);
nand U6988 (N_6988,N_5797,N_5573);
and U6989 (N_6989,N_5196,N_5935);
nor U6990 (N_6990,N_5146,N_5159);
nor U6991 (N_6991,N_5888,N_5649);
nor U6992 (N_6992,N_5913,N_5038);
nor U6993 (N_6993,N_5961,N_5208);
or U6994 (N_6994,N_5429,N_5761);
or U6995 (N_6995,N_5167,N_5190);
or U6996 (N_6996,N_5249,N_5933);
xor U6997 (N_6997,N_5453,N_5508);
or U6998 (N_6998,N_5996,N_5516);
or U6999 (N_6999,N_5292,N_5585);
nor U7000 (N_7000,N_6450,N_6532);
nor U7001 (N_7001,N_6157,N_6358);
nor U7002 (N_7002,N_6688,N_6136);
nor U7003 (N_7003,N_6365,N_6918);
nand U7004 (N_7004,N_6772,N_6910);
and U7005 (N_7005,N_6721,N_6329);
or U7006 (N_7006,N_6602,N_6463);
or U7007 (N_7007,N_6300,N_6205);
nand U7008 (N_7008,N_6481,N_6742);
nand U7009 (N_7009,N_6440,N_6891);
nor U7010 (N_7010,N_6022,N_6853);
xnor U7011 (N_7011,N_6550,N_6207);
nor U7012 (N_7012,N_6869,N_6786);
or U7013 (N_7013,N_6752,N_6023);
nor U7014 (N_7014,N_6055,N_6222);
nor U7015 (N_7015,N_6650,N_6925);
and U7016 (N_7016,N_6470,N_6792);
and U7017 (N_7017,N_6027,N_6405);
nor U7018 (N_7018,N_6283,N_6050);
or U7019 (N_7019,N_6131,N_6421);
nor U7020 (N_7020,N_6590,N_6195);
or U7021 (N_7021,N_6194,N_6780);
xnor U7022 (N_7022,N_6956,N_6635);
nand U7023 (N_7023,N_6821,N_6731);
nand U7024 (N_7024,N_6913,N_6390);
nand U7025 (N_7025,N_6460,N_6416);
and U7026 (N_7026,N_6293,N_6709);
nor U7027 (N_7027,N_6434,N_6989);
or U7028 (N_7028,N_6630,N_6690);
nor U7029 (N_7029,N_6503,N_6746);
and U7030 (N_7030,N_6987,N_6920);
and U7031 (N_7031,N_6980,N_6156);
or U7032 (N_7032,N_6308,N_6148);
nor U7033 (N_7033,N_6596,N_6897);
nand U7034 (N_7034,N_6697,N_6419);
or U7035 (N_7035,N_6408,N_6342);
nand U7036 (N_7036,N_6519,N_6095);
xnor U7037 (N_7037,N_6739,N_6415);
xnor U7038 (N_7038,N_6998,N_6243);
or U7039 (N_7039,N_6430,N_6474);
or U7040 (N_7040,N_6379,N_6391);
xnor U7041 (N_7041,N_6042,N_6097);
and U7042 (N_7042,N_6587,N_6737);
and U7043 (N_7043,N_6318,N_6583);
or U7044 (N_7044,N_6571,N_6139);
nand U7045 (N_7045,N_6830,N_6996);
xnor U7046 (N_7046,N_6132,N_6137);
and U7047 (N_7047,N_6158,N_6109);
nand U7048 (N_7048,N_6842,N_6193);
or U7049 (N_7049,N_6225,N_6727);
and U7050 (N_7050,N_6764,N_6404);
and U7051 (N_7051,N_6327,N_6932);
nor U7052 (N_7052,N_6570,N_6025);
nor U7053 (N_7053,N_6502,N_6791);
and U7054 (N_7054,N_6620,N_6685);
or U7055 (N_7055,N_6217,N_6312);
or U7056 (N_7056,N_6352,N_6089);
xnor U7057 (N_7057,N_6304,N_6058);
and U7058 (N_7058,N_6941,N_6281);
and U7059 (N_7059,N_6829,N_6515);
or U7060 (N_7060,N_6238,N_6950);
nand U7061 (N_7061,N_6972,N_6862);
and U7062 (N_7062,N_6107,N_6494);
nand U7063 (N_7063,N_6591,N_6401);
nand U7064 (N_7064,N_6499,N_6579);
nand U7065 (N_7065,N_6744,N_6464);
nor U7066 (N_7066,N_6264,N_6626);
and U7067 (N_7067,N_6256,N_6751);
nand U7068 (N_7068,N_6654,N_6868);
nor U7069 (N_7069,N_6334,N_6483);
nor U7070 (N_7070,N_6728,N_6310);
and U7071 (N_7071,N_6576,N_6274);
and U7072 (N_7072,N_6533,N_6858);
and U7073 (N_7073,N_6625,N_6134);
and U7074 (N_7074,N_6065,N_6230);
nand U7075 (N_7075,N_6767,N_6438);
nor U7076 (N_7076,N_6774,N_6954);
xnor U7077 (N_7077,N_6554,N_6114);
and U7078 (N_7078,N_6497,N_6926);
and U7079 (N_7079,N_6616,N_6286);
or U7080 (N_7080,N_6878,N_6290);
xor U7081 (N_7081,N_6796,N_6066);
nor U7082 (N_7082,N_6899,N_6078);
nor U7083 (N_7083,N_6660,N_6810);
or U7084 (N_7084,N_6642,N_6967);
nand U7085 (N_7085,N_6944,N_6887);
or U7086 (N_7086,N_6738,N_6825);
nand U7087 (N_7087,N_6113,N_6611);
nand U7088 (N_7088,N_6766,N_6695);
nor U7089 (N_7089,N_6258,N_6455);
or U7090 (N_7090,N_6535,N_6407);
or U7091 (N_7091,N_6666,N_6511);
nor U7092 (N_7092,N_6229,N_6876);
nand U7093 (N_7093,N_6632,N_6002);
xor U7094 (N_7094,N_6668,N_6553);
or U7095 (N_7095,N_6387,N_6296);
xor U7096 (N_7096,N_6990,N_6043);
xor U7097 (N_7097,N_6127,N_6513);
nor U7098 (N_7098,N_6077,N_6924);
nor U7099 (N_7099,N_6565,N_6558);
or U7100 (N_7100,N_6277,N_6729);
and U7101 (N_7101,N_6867,N_6453);
xnor U7102 (N_7102,N_6209,N_6595);
nor U7103 (N_7103,N_6098,N_6566);
xnor U7104 (N_7104,N_6272,N_6561);
nor U7105 (N_7105,N_6382,N_6469);
nor U7106 (N_7106,N_6864,N_6601);
xor U7107 (N_7107,N_6659,N_6241);
xnor U7108 (N_7108,N_6639,N_6377);
xnor U7109 (N_7109,N_6907,N_6017);
and U7110 (N_7110,N_6273,N_6648);
nor U7111 (N_7111,N_6613,N_6444);
xnor U7112 (N_7112,N_6108,N_6619);
nand U7113 (N_7113,N_6348,N_6894);
xnor U7114 (N_7114,N_6573,N_6201);
and U7115 (N_7115,N_6458,N_6734);
nor U7116 (N_7116,N_6933,N_6884);
nand U7117 (N_7117,N_6009,N_6640);
xor U7118 (N_7118,N_6285,N_6518);
and U7119 (N_7119,N_6543,N_6331);
nand U7120 (N_7120,N_6152,N_6768);
nand U7121 (N_7121,N_6784,N_6992);
xor U7122 (N_7122,N_6054,N_6865);
nor U7123 (N_7123,N_6577,N_6046);
and U7124 (N_7124,N_6653,N_6788);
or U7125 (N_7125,N_6008,N_6180);
or U7126 (N_7126,N_6551,N_6722);
xnor U7127 (N_7127,N_6983,N_6999);
nor U7128 (N_7128,N_6720,N_6667);
xor U7129 (N_7129,N_6889,N_6384);
nor U7130 (N_7130,N_6643,N_6228);
nor U7131 (N_7131,N_6362,N_6257);
nand U7132 (N_7132,N_6112,N_6445);
nor U7133 (N_7133,N_6208,N_6517);
and U7134 (N_7134,N_6693,N_6824);
or U7135 (N_7135,N_6614,N_6586);
xnor U7136 (N_7136,N_6725,N_6656);
nand U7137 (N_7137,N_6147,N_6185);
and U7138 (N_7138,N_6429,N_6875);
nor U7139 (N_7139,N_6339,N_6366);
nor U7140 (N_7140,N_6712,N_6846);
or U7141 (N_7141,N_6530,N_6874);
nor U7142 (N_7142,N_6756,N_6520);
nor U7143 (N_7143,N_6588,N_6462);
nand U7144 (N_7144,N_6562,N_6947);
nand U7145 (N_7145,N_6930,N_6549);
nor U7146 (N_7146,N_6169,N_6350);
nand U7147 (N_7147,N_6968,N_6014);
or U7148 (N_7148,N_6188,N_6291);
nand U7149 (N_7149,N_6809,N_6432);
nand U7150 (N_7150,N_6982,N_6634);
nand U7151 (N_7151,N_6580,N_6710);
or U7152 (N_7152,N_6206,N_6093);
nand U7153 (N_7153,N_6378,N_6370);
and U7154 (N_7154,N_6593,N_6584);
and U7155 (N_7155,N_6397,N_6904);
nor U7156 (N_7156,N_6969,N_6509);
xor U7157 (N_7157,N_6822,N_6942);
or U7158 (N_7158,N_6603,N_6957);
xor U7159 (N_7159,N_6371,N_6182);
nor U7160 (N_7160,N_6548,N_6563);
nand U7161 (N_7161,N_6399,N_6317);
or U7162 (N_7162,N_6485,N_6605);
nor U7163 (N_7163,N_6525,N_6164);
nand U7164 (N_7164,N_6841,N_6029);
nor U7165 (N_7165,N_6087,N_6016);
and U7166 (N_7166,N_6010,N_6198);
nand U7167 (N_7167,N_6504,N_6376);
xnor U7168 (N_7168,N_6001,N_6321);
xnor U7169 (N_7169,N_6447,N_6231);
xor U7170 (N_7170,N_6121,N_6964);
nand U7171 (N_7171,N_6621,N_6070);
xnor U7172 (N_7172,N_6383,N_6675);
or U7173 (N_7173,N_6528,N_6105);
xor U7174 (N_7174,N_6807,N_6475);
and U7175 (N_7175,N_6467,N_6030);
and U7176 (N_7176,N_6978,N_6024);
or U7177 (N_7177,N_6575,N_6159);
nand U7178 (N_7178,N_6993,N_6816);
nor U7179 (N_7179,N_6388,N_6119);
nor U7180 (N_7180,N_6946,N_6249);
and U7181 (N_7181,N_6879,N_6961);
and U7182 (N_7182,N_6804,N_6628);
or U7183 (N_7183,N_6117,N_6615);
and U7184 (N_7184,N_6314,N_6820);
nor U7185 (N_7185,N_6326,N_6911);
nand U7186 (N_7186,N_6179,N_6624);
or U7187 (N_7187,N_6652,N_6330);
nand U7188 (N_7188,N_6202,N_6061);
or U7189 (N_7189,N_6236,N_6880);
nand U7190 (N_7190,N_6689,N_6958);
xnor U7191 (N_7191,N_6790,N_6817);
or U7192 (N_7192,N_6902,N_6457);
and U7193 (N_7193,N_6110,N_6263);
nor U7194 (N_7194,N_6364,N_6507);
nor U7195 (N_7195,N_6482,N_6031);
or U7196 (N_7196,N_6995,N_6336);
nor U7197 (N_7197,N_6120,N_6698);
nand U7198 (N_7198,N_6071,N_6232);
or U7199 (N_7199,N_6011,N_6204);
xor U7200 (N_7200,N_6569,N_6522);
or U7201 (N_7201,N_6765,N_6026);
xnor U7202 (N_7202,N_6333,N_6191);
or U7203 (N_7203,N_6403,N_6374);
xnor U7204 (N_7204,N_6048,N_6708);
xnor U7205 (N_7205,N_6092,N_6262);
xnor U7206 (N_7206,N_6715,N_6612);
and U7207 (N_7207,N_6960,N_6800);
and U7208 (N_7208,N_6437,N_6581);
nand U7209 (N_7209,N_6045,N_6053);
or U7210 (N_7210,N_6498,N_6610);
and U7211 (N_7211,N_6069,N_6349);
xor U7212 (N_7212,N_6711,N_6510);
nand U7213 (N_7213,N_6559,N_6177);
xor U7214 (N_7214,N_6673,N_6245);
and U7215 (N_7215,N_6276,N_6707);
nor U7216 (N_7216,N_6854,N_6325);
nor U7217 (N_7217,N_6776,N_6490);
or U7218 (N_7218,N_6672,N_6724);
nor U7219 (N_7219,N_6931,N_6417);
nor U7220 (N_7220,N_6948,N_6135);
nor U7221 (N_7221,N_6372,N_6815);
xor U7222 (N_7222,N_6090,N_6893);
and U7223 (N_7223,N_6827,N_6056);
xor U7224 (N_7224,N_6699,N_6221);
or U7225 (N_7225,N_6622,N_6847);
and U7226 (N_7226,N_6541,N_6051);
or U7227 (N_7227,N_6203,N_6487);
xor U7228 (N_7228,N_6844,N_6898);
xnor U7229 (N_7229,N_6523,N_6637);
or U7230 (N_7230,N_6534,N_6919);
or U7231 (N_7231,N_6736,N_6289);
xnor U7232 (N_7232,N_6977,N_6723);
nor U7233 (N_7233,N_6446,N_6126);
nor U7234 (N_7234,N_6769,N_6848);
xor U7235 (N_7235,N_6934,N_6338);
nor U7236 (N_7236,N_6044,N_6828);
xnor U7237 (N_7237,N_6890,N_6806);
or U7238 (N_7238,N_6428,N_6020);
or U7239 (N_7239,N_6861,N_6812);
and U7240 (N_7240,N_6315,N_6150);
nor U7241 (N_7241,N_6213,N_6261);
xor U7242 (N_7242,N_6718,N_6521);
or U7243 (N_7243,N_6545,N_6211);
and U7244 (N_7244,N_6060,N_6531);
and U7245 (N_7245,N_6166,N_6857);
nand U7246 (N_7246,N_6655,N_6514);
and U7247 (N_7247,N_6702,N_6785);
nor U7248 (N_7248,N_6970,N_6955);
or U7249 (N_7249,N_6818,N_6441);
and U7250 (N_7250,N_6067,N_6813);
xnor U7251 (N_7251,N_6162,N_6381);
nor U7252 (N_7252,N_6142,N_6538);
or U7253 (N_7253,N_6552,N_6762);
nor U7254 (N_7254,N_6295,N_6560);
xnor U7255 (N_7255,N_6100,N_6091);
and U7256 (N_7256,N_6599,N_6248);
xor U7257 (N_7257,N_6268,N_6086);
xnor U7258 (N_7258,N_6506,N_6598);
and U7259 (N_7259,N_6294,N_6665);
or U7260 (N_7260,N_6369,N_6837);
nor U7261 (N_7261,N_6251,N_6811);
or U7262 (N_7262,N_6144,N_6354);
xnor U7263 (N_7263,N_6988,N_6224);
xnor U7264 (N_7264,N_6781,N_6540);
xor U7265 (N_7265,N_6787,N_6396);
and U7266 (N_7266,N_6214,N_6143);
nand U7267 (N_7267,N_6465,N_6075);
xor U7268 (N_7268,N_6883,N_6505);
or U7269 (N_7269,N_6491,N_6305);
or U7270 (N_7270,N_6351,N_6081);
nor U7271 (N_7271,N_6994,N_6705);
nor U7272 (N_7272,N_6280,N_6892);
nand U7273 (N_7273,N_6963,N_6840);
nand U7274 (N_7274,N_6122,N_6471);
nand U7275 (N_7275,N_6420,N_6319);
or U7276 (N_7276,N_6937,N_6452);
nor U7277 (N_7277,N_6151,N_6129);
xor U7278 (N_7278,N_6753,N_6664);
and U7279 (N_7279,N_6448,N_6244);
and U7280 (N_7280,N_6782,N_6138);
xor U7281 (N_7281,N_6473,N_6917);
nor U7282 (N_7282,N_6976,N_6145);
xnor U7283 (N_7283,N_6835,N_6353);
xnor U7284 (N_7284,N_6476,N_6537);
or U7285 (N_7285,N_6116,N_6466);
or U7286 (N_7286,N_6442,N_6953);
or U7287 (N_7287,N_6409,N_6539);
nor U7288 (N_7288,N_6343,N_6716);
nor U7289 (N_7289,N_6860,N_6758);
and U7290 (N_7290,N_6508,N_6971);
nor U7291 (N_7291,N_6922,N_6704);
nand U7292 (N_7292,N_6747,N_6255);
and U7293 (N_7293,N_6410,N_6219);
nand U7294 (N_7294,N_6076,N_6657);
xnor U7295 (N_7295,N_6808,N_6297);
and U7296 (N_7296,N_6123,N_6984);
xor U7297 (N_7297,N_6269,N_6555);
or U7298 (N_7298,N_6717,N_6527);
xnor U7299 (N_7299,N_6423,N_6082);
or U7300 (N_7300,N_6303,N_6355);
nor U7301 (N_7301,N_6775,N_6233);
or U7302 (N_7302,N_6028,N_6052);
xnor U7303 (N_7303,N_6335,N_6951);
or U7304 (N_7304,N_6118,N_6085);
and U7305 (N_7305,N_6265,N_6083);
and U7306 (N_7306,N_6160,N_6801);
or U7307 (N_7307,N_6062,N_6627);
nand U7308 (N_7308,N_6492,N_6478);
or U7309 (N_7309,N_6703,N_6341);
nand U7310 (N_7310,N_6111,N_6823);
xor U7311 (N_7311,N_6495,N_6174);
xnor U7312 (N_7312,N_6568,N_6037);
nor U7313 (N_7313,N_6006,N_6748);
or U7314 (N_7314,N_6877,N_6005);
nand U7315 (N_7315,N_6146,N_6683);
nand U7316 (N_7316,N_6176,N_6965);
nand U7317 (N_7317,N_6885,N_6674);
nor U7318 (N_7318,N_6328,N_6099);
nand U7319 (N_7319,N_6018,N_6292);
or U7320 (N_7320,N_6658,N_6484);
and U7321 (N_7321,N_6400,N_6344);
or U7322 (N_7322,N_6691,N_6713);
nand U7323 (N_7323,N_6459,N_6451);
or U7324 (N_7324,N_6102,N_6638);
nor U7325 (N_7325,N_6168,N_6313);
or U7326 (N_7326,N_6536,N_6866);
nor U7327 (N_7327,N_6896,N_6486);
nor U7328 (N_7328,N_6803,N_6585);
nor U7329 (N_7329,N_6247,N_6743);
and U7330 (N_7330,N_6914,N_6124);
and U7331 (N_7331,N_6629,N_6080);
and U7332 (N_7332,N_6216,N_6088);
or U7333 (N_7333,N_6493,N_6196);
nor U7334 (N_7334,N_6049,N_6929);
or U7335 (N_7335,N_6959,N_6347);
xor U7336 (N_7336,N_6516,N_6385);
xor U7337 (N_7337,N_6337,N_6719);
nand U7338 (N_7338,N_6849,N_6443);
or U7339 (N_7339,N_6242,N_6661);
nand U7340 (N_7340,N_6461,N_6073);
nor U7341 (N_7341,N_6836,N_6427);
and U7342 (N_7342,N_6171,N_6740);
and U7343 (N_7343,N_6367,N_6794);
nand U7344 (N_7344,N_6906,N_6912);
xor U7345 (N_7345,N_6418,N_6096);
or U7346 (N_7346,N_6477,N_6047);
nand U7347 (N_7347,N_6547,N_6870);
xor U7348 (N_7348,N_6040,N_6278);
or U7349 (N_7349,N_6745,N_6797);
nand U7350 (N_7350,N_6072,N_6680);
nor U7351 (N_7351,N_6212,N_6732);
nand U7352 (N_7352,N_6838,N_6940);
and U7353 (N_7353,N_6340,N_6411);
xnor U7354 (N_7354,N_6104,N_6750);
nor U7355 (N_7355,N_6007,N_6299);
nand U7356 (N_7356,N_6155,N_6019);
nand U7357 (N_7357,N_6240,N_6163);
xnor U7358 (N_7358,N_6927,N_6760);
or U7359 (N_7359,N_6036,N_6633);
nor U7360 (N_7360,N_6597,N_6779);
nor U7361 (N_7361,N_6239,N_6015);
and U7362 (N_7362,N_6345,N_6210);
xor U7363 (N_7363,N_6192,N_6393);
nand U7364 (N_7364,N_6275,N_6033);
xor U7365 (N_7365,N_6886,N_6952);
nand U7366 (N_7366,N_6454,N_6916);
or U7367 (N_7367,N_6644,N_6422);
and U7368 (N_7368,N_6153,N_6662);
and U7369 (N_7369,N_6677,N_6681);
and U7370 (N_7370,N_6394,N_6701);
or U7371 (N_7371,N_6714,N_6623);
and U7372 (N_7372,N_6363,N_6903);
nor U7373 (N_7373,N_6754,N_6641);
and U7374 (N_7374,N_6449,N_6755);
or U7375 (N_7375,N_6309,N_6106);
or U7376 (N_7376,N_6572,N_6636);
or U7377 (N_7377,N_6395,N_6252);
xnor U7378 (N_7378,N_6426,N_6981);
xor U7379 (N_7379,N_6288,N_6939);
nand U7380 (N_7380,N_6359,N_6564);
xor U7381 (N_7381,N_6038,N_6798);
xor U7382 (N_7382,N_6094,N_6021);
xnor U7383 (N_7383,N_6424,N_6831);
nand U7384 (N_7384,N_6068,N_6279);
or U7385 (N_7385,N_6472,N_6512);
and U7386 (N_7386,N_6253,N_6175);
nand U7387 (N_7387,N_6556,N_6726);
nand U7388 (N_7388,N_6189,N_6749);
nor U7389 (N_7389,N_6041,N_6489);
nand U7390 (N_7390,N_6413,N_6425);
and U7391 (N_7391,N_6928,N_6997);
and U7392 (N_7392,N_6852,N_6479);
nor U7393 (N_7393,N_6901,N_6183);
nor U7394 (N_7394,N_6979,N_6406);
and U7395 (N_7395,N_6582,N_6500);
or U7396 (N_7396,N_6872,N_6735);
and U7397 (N_7397,N_6307,N_6819);
nor U7398 (N_7398,N_6943,N_6684);
xor U7399 (N_7399,N_6435,N_6254);
xnor U7400 (N_7400,N_6003,N_6687);
and U7401 (N_7401,N_6199,N_6607);
or U7402 (N_7402,N_6480,N_6266);
nor U7403 (N_7403,N_6834,N_6115);
nand U7404 (N_7404,N_6973,N_6215);
xor U7405 (N_7405,N_6084,N_6696);
or U7406 (N_7406,N_6935,N_6287);
or U7407 (N_7407,N_6170,N_6074);
nand U7408 (N_7408,N_6826,N_6686);
nor U7409 (N_7409,N_6012,N_6799);
nor U7410 (N_7410,N_6647,N_6227);
or U7411 (N_7411,N_6789,N_6671);
xnor U7412 (N_7412,N_6682,N_6373);
and U7413 (N_7413,N_6140,N_6496);
and U7414 (N_7414,N_6649,N_6133);
nor U7415 (N_7415,N_6759,N_6356);
nand U7416 (N_7416,N_6234,N_6375);
nand U7417 (N_7417,N_6845,N_6246);
xor U7418 (N_7418,N_6962,N_6154);
nor U7419 (N_7419,N_6832,N_6778);
nand U7420 (N_7420,N_6368,N_6795);
or U7421 (N_7421,N_6173,N_6197);
or U7422 (N_7422,N_6178,N_6802);
nand U7423 (N_7423,N_6915,N_6125);
nor U7424 (N_7424,N_6524,N_6574);
xnor U7425 (N_7425,N_6311,N_6346);
and U7426 (N_7426,N_6592,N_6035);
or U7427 (N_7427,N_6651,N_6167);
nor U7428 (N_7428,N_6617,N_6600);
or U7429 (N_7429,N_6439,N_6161);
nand U7430 (N_7430,N_6526,N_6186);
or U7431 (N_7431,N_6398,N_6986);
and U7432 (N_7432,N_6850,N_6900);
and U7433 (N_7433,N_6895,N_6670);
nand U7434 (N_7434,N_6360,N_6282);
nand U7435 (N_7435,N_6646,N_6678);
and U7436 (N_7436,N_6361,N_6057);
xor U7437 (N_7437,N_6542,N_6267);
xnor U7438 (N_7438,N_6730,N_6908);
xnor U7439 (N_7439,N_6783,N_6706);
nor U7440 (N_7440,N_6320,N_6260);
nor U7441 (N_7441,N_6259,N_6284);
xor U7442 (N_7442,N_6606,N_6034);
or U7443 (N_7443,N_6488,N_6692);
xnor U7444 (N_7444,N_6851,N_6843);
nor U7445 (N_7445,N_6814,N_6544);
nor U7446 (N_7446,N_6546,N_6389);
nor U7447 (N_7447,N_6676,N_6468);
and U7448 (N_7448,N_6921,N_6936);
xor U7449 (N_7449,N_6141,N_6741);
and U7450 (N_7450,N_6966,N_6187);
nor U7451 (N_7451,N_6863,N_6763);
or U7452 (N_7452,N_6923,N_6985);
nand U7453 (N_7453,N_6032,N_6000);
xnor U7454 (N_7454,N_6529,N_6975);
nor U7455 (N_7455,N_6223,N_6700);
nand U7456 (N_7456,N_6130,N_6938);
xor U7457 (N_7457,N_6905,N_6380);
xor U7458 (N_7458,N_6101,N_6805);
or U7459 (N_7459,N_6190,N_6645);
nor U7460 (N_7460,N_6589,N_6298);
and U7461 (N_7461,N_6103,N_6172);
and U7462 (N_7462,N_6433,N_6039);
nand U7463 (N_7463,N_6250,N_6679);
and U7464 (N_7464,N_6501,N_6974);
and U7465 (N_7465,N_6833,N_6608);
nor U7466 (N_7466,N_6306,N_6200);
and U7467 (N_7467,N_6873,N_6567);
nor U7468 (N_7468,N_6165,N_6557);
nor U7469 (N_7469,N_6324,N_6436);
nand U7470 (N_7470,N_6059,N_6323);
or U7471 (N_7471,N_6063,N_6149);
and U7472 (N_7472,N_6064,N_6386);
or U7473 (N_7473,N_6856,N_6663);
nand U7474 (N_7474,N_6322,N_6332);
nor U7475 (N_7475,N_6316,N_6237);
or U7476 (N_7476,N_6609,N_6909);
xnor U7477 (N_7477,N_6773,N_6301);
nor U7478 (N_7478,N_6757,N_6181);
nand U7479 (N_7479,N_6694,N_6226);
nand U7480 (N_7480,N_6184,N_6218);
nor U7481 (N_7481,N_6235,N_6949);
nand U7482 (N_7482,N_6604,N_6357);
or U7483 (N_7483,N_6128,N_6855);
nor U7484 (N_7484,N_6013,N_6412);
xnor U7485 (N_7485,N_6392,N_6402);
nor U7486 (N_7486,N_6882,N_6594);
and U7487 (N_7487,N_6302,N_6991);
nand U7488 (N_7488,N_6669,N_6004);
nor U7489 (N_7489,N_6079,N_6881);
xor U7490 (N_7490,N_6871,N_6761);
and U7491 (N_7491,N_6431,N_6771);
nor U7492 (N_7492,N_6733,N_6859);
and U7493 (N_7493,N_6793,N_6839);
nor U7494 (N_7494,N_6271,N_6770);
or U7495 (N_7495,N_6456,N_6220);
xor U7496 (N_7496,N_6888,N_6945);
nand U7497 (N_7497,N_6631,N_6414);
nand U7498 (N_7498,N_6618,N_6578);
or U7499 (N_7499,N_6270,N_6777);
nand U7500 (N_7500,N_6994,N_6932);
or U7501 (N_7501,N_6210,N_6025);
or U7502 (N_7502,N_6418,N_6065);
nor U7503 (N_7503,N_6397,N_6207);
and U7504 (N_7504,N_6254,N_6720);
xor U7505 (N_7505,N_6698,N_6048);
xnor U7506 (N_7506,N_6280,N_6541);
nor U7507 (N_7507,N_6598,N_6582);
or U7508 (N_7508,N_6218,N_6291);
and U7509 (N_7509,N_6734,N_6704);
and U7510 (N_7510,N_6112,N_6487);
and U7511 (N_7511,N_6226,N_6657);
or U7512 (N_7512,N_6168,N_6470);
nor U7513 (N_7513,N_6725,N_6862);
nand U7514 (N_7514,N_6714,N_6955);
xor U7515 (N_7515,N_6101,N_6620);
or U7516 (N_7516,N_6344,N_6706);
nor U7517 (N_7517,N_6022,N_6143);
nand U7518 (N_7518,N_6635,N_6287);
and U7519 (N_7519,N_6948,N_6041);
xor U7520 (N_7520,N_6151,N_6303);
xor U7521 (N_7521,N_6490,N_6686);
xor U7522 (N_7522,N_6008,N_6145);
xor U7523 (N_7523,N_6183,N_6353);
or U7524 (N_7524,N_6001,N_6006);
and U7525 (N_7525,N_6833,N_6847);
xnor U7526 (N_7526,N_6349,N_6774);
nor U7527 (N_7527,N_6160,N_6688);
and U7528 (N_7528,N_6249,N_6484);
and U7529 (N_7529,N_6765,N_6683);
nand U7530 (N_7530,N_6706,N_6286);
xnor U7531 (N_7531,N_6568,N_6246);
and U7532 (N_7532,N_6916,N_6185);
xor U7533 (N_7533,N_6017,N_6395);
and U7534 (N_7534,N_6076,N_6618);
and U7535 (N_7535,N_6420,N_6565);
nand U7536 (N_7536,N_6585,N_6282);
nand U7537 (N_7537,N_6214,N_6201);
nor U7538 (N_7538,N_6427,N_6494);
or U7539 (N_7539,N_6218,N_6622);
and U7540 (N_7540,N_6604,N_6725);
nand U7541 (N_7541,N_6577,N_6318);
nor U7542 (N_7542,N_6399,N_6446);
nand U7543 (N_7543,N_6625,N_6180);
xor U7544 (N_7544,N_6580,N_6610);
or U7545 (N_7545,N_6043,N_6400);
nor U7546 (N_7546,N_6941,N_6098);
nor U7547 (N_7547,N_6856,N_6379);
and U7548 (N_7548,N_6188,N_6276);
nand U7549 (N_7549,N_6564,N_6996);
and U7550 (N_7550,N_6725,N_6097);
nand U7551 (N_7551,N_6963,N_6441);
xor U7552 (N_7552,N_6321,N_6011);
xor U7553 (N_7553,N_6580,N_6653);
xor U7554 (N_7554,N_6921,N_6137);
nand U7555 (N_7555,N_6233,N_6931);
nand U7556 (N_7556,N_6987,N_6178);
xor U7557 (N_7557,N_6243,N_6985);
or U7558 (N_7558,N_6824,N_6888);
or U7559 (N_7559,N_6863,N_6261);
or U7560 (N_7560,N_6711,N_6642);
nand U7561 (N_7561,N_6124,N_6572);
nand U7562 (N_7562,N_6509,N_6578);
nand U7563 (N_7563,N_6940,N_6184);
xor U7564 (N_7564,N_6362,N_6232);
nand U7565 (N_7565,N_6449,N_6946);
or U7566 (N_7566,N_6719,N_6081);
nor U7567 (N_7567,N_6012,N_6307);
nor U7568 (N_7568,N_6148,N_6848);
or U7569 (N_7569,N_6168,N_6749);
and U7570 (N_7570,N_6011,N_6777);
xnor U7571 (N_7571,N_6056,N_6210);
xor U7572 (N_7572,N_6025,N_6369);
or U7573 (N_7573,N_6450,N_6056);
nand U7574 (N_7574,N_6680,N_6149);
xor U7575 (N_7575,N_6708,N_6924);
and U7576 (N_7576,N_6227,N_6039);
and U7577 (N_7577,N_6250,N_6629);
nor U7578 (N_7578,N_6657,N_6532);
and U7579 (N_7579,N_6617,N_6807);
nand U7580 (N_7580,N_6287,N_6076);
nor U7581 (N_7581,N_6941,N_6890);
or U7582 (N_7582,N_6766,N_6945);
xor U7583 (N_7583,N_6293,N_6743);
nand U7584 (N_7584,N_6658,N_6049);
nor U7585 (N_7585,N_6876,N_6372);
xor U7586 (N_7586,N_6721,N_6692);
and U7587 (N_7587,N_6802,N_6717);
nand U7588 (N_7588,N_6482,N_6973);
xnor U7589 (N_7589,N_6575,N_6045);
or U7590 (N_7590,N_6718,N_6967);
and U7591 (N_7591,N_6036,N_6494);
xor U7592 (N_7592,N_6877,N_6312);
nand U7593 (N_7593,N_6494,N_6570);
xor U7594 (N_7594,N_6849,N_6166);
or U7595 (N_7595,N_6636,N_6427);
or U7596 (N_7596,N_6278,N_6739);
nand U7597 (N_7597,N_6356,N_6171);
or U7598 (N_7598,N_6344,N_6683);
nor U7599 (N_7599,N_6511,N_6186);
xnor U7600 (N_7600,N_6081,N_6821);
nand U7601 (N_7601,N_6585,N_6661);
nor U7602 (N_7602,N_6204,N_6701);
nand U7603 (N_7603,N_6088,N_6821);
xnor U7604 (N_7604,N_6874,N_6942);
or U7605 (N_7605,N_6691,N_6383);
and U7606 (N_7606,N_6049,N_6751);
nor U7607 (N_7607,N_6343,N_6795);
nand U7608 (N_7608,N_6365,N_6199);
nor U7609 (N_7609,N_6055,N_6775);
xor U7610 (N_7610,N_6730,N_6781);
or U7611 (N_7611,N_6996,N_6130);
or U7612 (N_7612,N_6875,N_6331);
xor U7613 (N_7613,N_6697,N_6839);
and U7614 (N_7614,N_6281,N_6098);
and U7615 (N_7615,N_6214,N_6473);
xnor U7616 (N_7616,N_6842,N_6313);
or U7617 (N_7617,N_6675,N_6440);
nor U7618 (N_7618,N_6465,N_6242);
nand U7619 (N_7619,N_6115,N_6511);
nor U7620 (N_7620,N_6222,N_6326);
xor U7621 (N_7621,N_6130,N_6684);
xnor U7622 (N_7622,N_6401,N_6342);
and U7623 (N_7623,N_6982,N_6461);
nor U7624 (N_7624,N_6359,N_6553);
and U7625 (N_7625,N_6428,N_6699);
nand U7626 (N_7626,N_6521,N_6128);
xnor U7627 (N_7627,N_6227,N_6648);
nand U7628 (N_7628,N_6847,N_6384);
nand U7629 (N_7629,N_6976,N_6670);
xnor U7630 (N_7630,N_6277,N_6837);
and U7631 (N_7631,N_6707,N_6105);
and U7632 (N_7632,N_6090,N_6418);
nand U7633 (N_7633,N_6048,N_6178);
xnor U7634 (N_7634,N_6169,N_6033);
nor U7635 (N_7635,N_6774,N_6958);
xnor U7636 (N_7636,N_6169,N_6466);
nand U7637 (N_7637,N_6169,N_6734);
nor U7638 (N_7638,N_6026,N_6173);
nand U7639 (N_7639,N_6497,N_6313);
nor U7640 (N_7640,N_6562,N_6676);
and U7641 (N_7641,N_6328,N_6829);
nor U7642 (N_7642,N_6260,N_6560);
or U7643 (N_7643,N_6082,N_6969);
or U7644 (N_7644,N_6421,N_6659);
nand U7645 (N_7645,N_6312,N_6168);
nor U7646 (N_7646,N_6651,N_6553);
xnor U7647 (N_7647,N_6236,N_6304);
and U7648 (N_7648,N_6072,N_6785);
nand U7649 (N_7649,N_6947,N_6675);
and U7650 (N_7650,N_6474,N_6482);
nor U7651 (N_7651,N_6818,N_6690);
nand U7652 (N_7652,N_6014,N_6244);
nand U7653 (N_7653,N_6046,N_6372);
nand U7654 (N_7654,N_6555,N_6408);
nor U7655 (N_7655,N_6557,N_6586);
and U7656 (N_7656,N_6956,N_6479);
xor U7657 (N_7657,N_6853,N_6824);
xnor U7658 (N_7658,N_6581,N_6419);
nand U7659 (N_7659,N_6366,N_6667);
or U7660 (N_7660,N_6407,N_6525);
and U7661 (N_7661,N_6213,N_6490);
nor U7662 (N_7662,N_6549,N_6513);
or U7663 (N_7663,N_6165,N_6474);
nand U7664 (N_7664,N_6255,N_6568);
nand U7665 (N_7665,N_6391,N_6903);
or U7666 (N_7666,N_6215,N_6004);
and U7667 (N_7667,N_6649,N_6551);
and U7668 (N_7668,N_6301,N_6108);
or U7669 (N_7669,N_6531,N_6490);
nor U7670 (N_7670,N_6554,N_6657);
or U7671 (N_7671,N_6396,N_6459);
xnor U7672 (N_7672,N_6523,N_6150);
xnor U7673 (N_7673,N_6812,N_6207);
and U7674 (N_7674,N_6276,N_6253);
xor U7675 (N_7675,N_6125,N_6291);
nor U7676 (N_7676,N_6495,N_6241);
or U7677 (N_7677,N_6951,N_6704);
or U7678 (N_7678,N_6088,N_6085);
and U7679 (N_7679,N_6552,N_6435);
or U7680 (N_7680,N_6630,N_6624);
nor U7681 (N_7681,N_6567,N_6589);
xnor U7682 (N_7682,N_6553,N_6912);
nor U7683 (N_7683,N_6956,N_6330);
xor U7684 (N_7684,N_6004,N_6992);
and U7685 (N_7685,N_6279,N_6447);
nor U7686 (N_7686,N_6481,N_6112);
and U7687 (N_7687,N_6303,N_6498);
nand U7688 (N_7688,N_6998,N_6200);
or U7689 (N_7689,N_6647,N_6927);
and U7690 (N_7690,N_6996,N_6089);
xor U7691 (N_7691,N_6910,N_6969);
xnor U7692 (N_7692,N_6281,N_6755);
or U7693 (N_7693,N_6762,N_6709);
xnor U7694 (N_7694,N_6422,N_6281);
or U7695 (N_7695,N_6313,N_6201);
or U7696 (N_7696,N_6436,N_6930);
and U7697 (N_7697,N_6090,N_6323);
nand U7698 (N_7698,N_6267,N_6593);
nand U7699 (N_7699,N_6712,N_6559);
xnor U7700 (N_7700,N_6555,N_6492);
nand U7701 (N_7701,N_6109,N_6308);
xor U7702 (N_7702,N_6284,N_6745);
nand U7703 (N_7703,N_6278,N_6053);
nor U7704 (N_7704,N_6699,N_6478);
nand U7705 (N_7705,N_6152,N_6980);
xor U7706 (N_7706,N_6409,N_6805);
xnor U7707 (N_7707,N_6746,N_6415);
and U7708 (N_7708,N_6975,N_6026);
nor U7709 (N_7709,N_6901,N_6740);
nand U7710 (N_7710,N_6094,N_6251);
xnor U7711 (N_7711,N_6411,N_6495);
or U7712 (N_7712,N_6848,N_6884);
nand U7713 (N_7713,N_6038,N_6919);
nor U7714 (N_7714,N_6835,N_6173);
nor U7715 (N_7715,N_6635,N_6060);
or U7716 (N_7716,N_6669,N_6792);
and U7717 (N_7717,N_6302,N_6844);
nand U7718 (N_7718,N_6312,N_6933);
or U7719 (N_7719,N_6883,N_6930);
nor U7720 (N_7720,N_6429,N_6651);
nand U7721 (N_7721,N_6198,N_6795);
and U7722 (N_7722,N_6194,N_6958);
nand U7723 (N_7723,N_6675,N_6927);
xor U7724 (N_7724,N_6402,N_6690);
nor U7725 (N_7725,N_6668,N_6251);
nand U7726 (N_7726,N_6112,N_6028);
and U7727 (N_7727,N_6379,N_6908);
or U7728 (N_7728,N_6567,N_6161);
or U7729 (N_7729,N_6511,N_6854);
and U7730 (N_7730,N_6306,N_6932);
xnor U7731 (N_7731,N_6314,N_6134);
xnor U7732 (N_7732,N_6349,N_6914);
nor U7733 (N_7733,N_6393,N_6432);
and U7734 (N_7734,N_6518,N_6006);
nor U7735 (N_7735,N_6491,N_6338);
and U7736 (N_7736,N_6500,N_6911);
and U7737 (N_7737,N_6215,N_6380);
and U7738 (N_7738,N_6504,N_6168);
or U7739 (N_7739,N_6110,N_6793);
xnor U7740 (N_7740,N_6016,N_6838);
nand U7741 (N_7741,N_6144,N_6427);
xor U7742 (N_7742,N_6390,N_6300);
nor U7743 (N_7743,N_6036,N_6952);
and U7744 (N_7744,N_6799,N_6471);
xor U7745 (N_7745,N_6320,N_6475);
or U7746 (N_7746,N_6364,N_6694);
nor U7747 (N_7747,N_6862,N_6101);
and U7748 (N_7748,N_6392,N_6106);
xnor U7749 (N_7749,N_6617,N_6903);
or U7750 (N_7750,N_6745,N_6016);
and U7751 (N_7751,N_6616,N_6086);
nand U7752 (N_7752,N_6430,N_6649);
or U7753 (N_7753,N_6342,N_6081);
or U7754 (N_7754,N_6764,N_6489);
nand U7755 (N_7755,N_6478,N_6227);
nand U7756 (N_7756,N_6839,N_6691);
nor U7757 (N_7757,N_6688,N_6403);
and U7758 (N_7758,N_6371,N_6670);
xnor U7759 (N_7759,N_6267,N_6207);
nor U7760 (N_7760,N_6559,N_6545);
or U7761 (N_7761,N_6684,N_6926);
nor U7762 (N_7762,N_6454,N_6466);
xor U7763 (N_7763,N_6369,N_6955);
nor U7764 (N_7764,N_6299,N_6755);
xor U7765 (N_7765,N_6178,N_6945);
nand U7766 (N_7766,N_6334,N_6790);
or U7767 (N_7767,N_6615,N_6575);
and U7768 (N_7768,N_6834,N_6125);
nand U7769 (N_7769,N_6623,N_6353);
xor U7770 (N_7770,N_6290,N_6560);
or U7771 (N_7771,N_6088,N_6994);
nand U7772 (N_7772,N_6235,N_6192);
or U7773 (N_7773,N_6116,N_6469);
and U7774 (N_7774,N_6119,N_6080);
nand U7775 (N_7775,N_6994,N_6752);
or U7776 (N_7776,N_6531,N_6907);
nor U7777 (N_7777,N_6257,N_6421);
and U7778 (N_7778,N_6432,N_6777);
xnor U7779 (N_7779,N_6331,N_6608);
nand U7780 (N_7780,N_6335,N_6719);
xnor U7781 (N_7781,N_6820,N_6735);
nand U7782 (N_7782,N_6679,N_6803);
or U7783 (N_7783,N_6777,N_6428);
nand U7784 (N_7784,N_6390,N_6850);
nand U7785 (N_7785,N_6531,N_6969);
and U7786 (N_7786,N_6074,N_6791);
nor U7787 (N_7787,N_6166,N_6564);
xor U7788 (N_7788,N_6439,N_6916);
or U7789 (N_7789,N_6503,N_6289);
xor U7790 (N_7790,N_6442,N_6234);
nor U7791 (N_7791,N_6216,N_6473);
or U7792 (N_7792,N_6091,N_6584);
or U7793 (N_7793,N_6604,N_6753);
and U7794 (N_7794,N_6762,N_6174);
and U7795 (N_7795,N_6436,N_6169);
and U7796 (N_7796,N_6257,N_6814);
nor U7797 (N_7797,N_6905,N_6459);
or U7798 (N_7798,N_6037,N_6189);
or U7799 (N_7799,N_6159,N_6481);
or U7800 (N_7800,N_6343,N_6597);
or U7801 (N_7801,N_6440,N_6342);
or U7802 (N_7802,N_6121,N_6859);
or U7803 (N_7803,N_6033,N_6415);
or U7804 (N_7804,N_6921,N_6150);
nand U7805 (N_7805,N_6328,N_6243);
nor U7806 (N_7806,N_6530,N_6347);
and U7807 (N_7807,N_6912,N_6463);
nor U7808 (N_7808,N_6480,N_6682);
xor U7809 (N_7809,N_6714,N_6300);
or U7810 (N_7810,N_6885,N_6374);
xnor U7811 (N_7811,N_6599,N_6091);
nand U7812 (N_7812,N_6147,N_6507);
nor U7813 (N_7813,N_6782,N_6557);
nor U7814 (N_7814,N_6012,N_6352);
and U7815 (N_7815,N_6969,N_6947);
nor U7816 (N_7816,N_6378,N_6604);
nor U7817 (N_7817,N_6249,N_6045);
xnor U7818 (N_7818,N_6076,N_6596);
nor U7819 (N_7819,N_6013,N_6717);
nand U7820 (N_7820,N_6466,N_6890);
and U7821 (N_7821,N_6969,N_6254);
and U7822 (N_7822,N_6620,N_6607);
or U7823 (N_7823,N_6641,N_6240);
nand U7824 (N_7824,N_6320,N_6750);
xnor U7825 (N_7825,N_6153,N_6159);
xor U7826 (N_7826,N_6618,N_6686);
or U7827 (N_7827,N_6903,N_6609);
nand U7828 (N_7828,N_6908,N_6315);
nor U7829 (N_7829,N_6501,N_6257);
nand U7830 (N_7830,N_6774,N_6372);
xor U7831 (N_7831,N_6628,N_6477);
xnor U7832 (N_7832,N_6801,N_6031);
or U7833 (N_7833,N_6413,N_6993);
or U7834 (N_7834,N_6443,N_6733);
nor U7835 (N_7835,N_6559,N_6144);
nor U7836 (N_7836,N_6051,N_6463);
xor U7837 (N_7837,N_6061,N_6022);
xnor U7838 (N_7838,N_6323,N_6216);
nand U7839 (N_7839,N_6442,N_6301);
and U7840 (N_7840,N_6819,N_6516);
nor U7841 (N_7841,N_6589,N_6508);
and U7842 (N_7842,N_6551,N_6261);
nand U7843 (N_7843,N_6609,N_6802);
and U7844 (N_7844,N_6444,N_6250);
nand U7845 (N_7845,N_6478,N_6621);
and U7846 (N_7846,N_6062,N_6725);
nand U7847 (N_7847,N_6855,N_6258);
nand U7848 (N_7848,N_6454,N_6785);
or U7849 (N_7849,N_6020,N_6129);
xnor U7850 (N_7850,N_6271,N_6356);
xor U7851 (N_7851,N_6034,N_6182);
nand U7852 (N_7852,N_6287,N_6937);
nor U7853 (N_7853,N_6318,N_6362);
or U7854 (N_7854,N_6708,N_6813);
nor U7855 (N_7855,N_6792,N_6199);
and U7856 (N_7856,N_6092,N_6151);
or U7857 (N_7857,N_6399,N_6129);
nand U7858 (N_7858,N_6514,N_6682);
and U7859 (N_7859,N_6534,N_6175);
nand U7860 (N_7860,N_6717,N_6263);
nand U7861 (N_7861,N_6922,N_6070);
nand U7862 (N_7862,N_6389,N_6937);
xor U7863 (N_7863,N_6122,N_6802);
xnor U7864 (N_7864,N_6728,N_6430);
nor U7865 (N_7865,N_6747,N_6294);
nand U7866 (N_7866,N_6536,N_6076);
nor U7867 (N_7867,N_6699,N_6932);
and U7868 (N_7868,N_6170,N_6856);
xor U7869 (N_7869,N_6639,N_6630);
or U7870 (N_7870,N_6994,N_6315);
and U7871 (N_7871,N_6861,N_6462);
and U7872 (N_7872,N_6998,N_6204);
nor U7873 (N_7873,N_6327,N_6513);
and U7874 (N_7874,N_6873,N_6799);
nor U7875 (N_7875,N_6045,N_6889);
and U7876 (N_7876,N_6044,N_6400);
or U7877 (N_7877,N_6388,N_6823);
nor U7878 (N_7878,N_6933,N_6741);
nor U7879 (N_7879,N_6900,N_6235);
xnor U7880 (N_7880,N_6936,N_6331);
and U7881 (N_7881,N_6787,N_6605);
xor U7882 (N_7882,N_6436,N_6874);
or U7883 (N_7883,N_6410,N_6836);
or U7884 (N_7884,N_6478,N_6351);
nor U7885 (N_7885,N_6464,N_6134);
nand U7886 (N_7886,N_6569,N_6946);
nor U7887 (N_7887,N_6971,N_6181);
xor U7888 (N_7888,N_6543,N_6248);
nand U7889 (N_7889,N_6131,N_6370);
nor U7890 (N_7890,N_6684,N_6646);
nor U7891 (N_7891,N_6893,N_6702);
nand U7892 (N_7892,N_6821,N_6480);
xor U7893 (N_7893,N_6916,N_6324);
nor U7894 (N_7894,N_6350,N_6379);
or U7895 (N_7895,N_6812,N_6691);
or U7896 (N_7896,N_6745,N_6634);
xnor U7897 (N_7897,N_6844,N_6458);
nand U7898 (N_7898,N_6689,N_6960);
and U7899 (N_7899,N_6239,N_6526);
nand U7900 (N_7900,N_6755,N_6197);
nand U7901 (N_7901,N_6108,N_6234);
nand U7902 (N_7902,N_6500,N_6565);
and U7903 (N_7903,N_6059,N_6567);
nand U7904 (N_7904,N_6433,N_6162);
nand U7905 (N_7905,N_6330,N_6463);
and U7906 (N_7906,N_6931,N_6278);
nand U7907 (N_7907,N_6875,N_6945);
xor U7908 (N_7908,N_6899,N_6670);
and U7909 (N_7909,N_6446,N_6105);
and U7910 (N_7910,N_6525,N_6214);
or U7911 (N_7911,N_6965,N_6664);
nor U7912 (N_7912,N_6581,N_6667);
nand U7913 (N_7913,N_6906,N_6365);
or U7914 (N_7914,N_6153,N_6338);
xnor U7915 (N_7915,N_6406,N_6443);
xnor U7916 (N_7916,N_6879,N_6804);
nor U7917 (N_7917,N_6228,N_6054);
nand U7918 (N_7918,N_6377,N_6596);
and U7919 (N_7919,N_6762,N_6462);
or U7920 (N_7920,N_6138,N_6747);
or U7921 (N_7921,N_6846,N_6023);
xnor U7922 (N_7922,N_6635,N_6639);
or U7923 (N_7923,N_6255,N_6322);
nand U7924 (N_7924,N_6286,N_6255);
and U7925 (N_7925,N_6063,N_6134);
or U7926 (N_7926,N_6950,N_6928);
xnor U7927 (N_7927,N_6029,N_6738);
nand U7928 (N_7928,N_6707,N_6261);
nand U7929 (N_7929,N_6008,N_6069);
xnor U7930 (N_7930,N_6539,N_6500);
and U7931 (N_7931,N_6976,N_6542);
and U7932 (N_7932,N_6073,N_6302);
or U7933 (N_7933,N_6589,N_6496);
nor U7934 (N_7934,N_6807,N_6517);
xnor U7935 (N_7935,N_6061,N_6527);
and U7936 (N_7936,N_6610,N_6786);
nor U7937 (N_7937,N_6951,N_6774);
and U7938 (N_7938,N_6871,N_6906);
and U7939 (N_7939,N_6801,N_6784);
nand U7940 (N_7940,N_6466,N_6637);
or U7941 (N_7941,N_6281,N_6354);
nand U7942 (N_7942,N_6849,N_6915);
xnor U7943 (N_7943,N_6889,N_6450);
or U7944 (N_7944,N_6398,N_6774);
nor U7945 (N_7945,N_6749,N_6481);
and U7946 (N_7946,N_6001,N_6507);
nand U7947 (N_7947,N_6396,N_6871);
or U7948 (N_7948,N_6436,N_6247);
and U7949 (N_7949,N_6079,N_6476);
nand U7950 (N_7950,N_6430,N_6476);
nand U7951 (N_7951,N_6869,N_6462);
nor U7952 (N_7952,N_6433,N_6058);
or U7953 (N_7953,N_6510,N_6788);
xnor U7954 (N_7954,N_6119,N_6205);
xnor U7955 (N_7955,N_6786,N_6795);
nand U7956 (N_7956,N_6119,N_6731);
or U7957 (N_7957,N_6573,N_6438);
xor U7958 (N_7958,N_6556,N_6420);
nor U7959 (N_7959,N_6733,N_6446);
nand U7960 (N_7960,N_6710,N_6752);
or U7961 (N_7961,N_6766,N_6240);
and U7962 (N_7962,N_6856,N_6893);
and U7963 (N_7963,N_6344,N_6982);
xnor U7964 (N_7964,N_6839,N_6253);
nor U7965 (N_7965,N_6192,N_6806);
xnor U7966 (N_7966,N_6479,N_6608);
or U7967 (N_7967,N_6870,N_6469);
and U7968 (N_7968,N_6629,N_6269);
nor U7969 (N_7969,N_6522,N_6702);
or U7970 (N_7970,N_6887,N_6249);
or U7971 (N_7971,N_6257,N_6533);
and U7972 (N_7972,N_6197,N_6448);
nor U7973 (N_7973,N_6334,N_6127);
and U7974 (N_7974,N_6216,N_6515);
and U7975 (N_7975,N_6496,N_6557);
and U7976 (N_7976,N_6252,N_6661);
or U7977 (N_7977,N_6793,N_6749);
nor U7978 (N_7978,N_6569,N_6568);
xnor U7979 (N_7979,N_6040,N_6103);
nand U7980 (N_7980,N_6743,N_6926);
nand U7981 (N_7981,N_6631,N_6290);
nor U7982 (N_7982,N_6225,N_6541);
nand U7983 (N_7983,N_6664,N_6605);
xor U7984 (N_7984,N_6152,N_6245);
nor U7985 (N_7985,N_6296,N_6902);
or U7986 (N_7986,N_6533,N_6158);
nor U7987 (N_7987,N_6383,N_6971);
xor U7988 (N_7988,N_6778,N_6831);
nor U7989 (N_7989,N_6914,N_6291);
nor U7990 (N_7990,N_6492,N_6406);
and U7991 (N_7991,N_6193,N_6267);
nand U7992 (N_7992,N_6551,N_6753);
xnor U7993 (N_7993,N_6695,N_6153);
xnor U7994 (N_7994,N_6168,N_6984);
nand U7995 (N_7995,N_6190,N_6521);
xnor U7996 (N_7996,N_6601,N_6328);
or U7997 (N_7997,N_6180,N_6030);
xnor U7998 (N_7998,N_6733,N_6438);
or U7999 (N_7999,N_6754,N_6070);
nand U8000 (N_8000,N_7717,N_7322);
or U8001 (N_8001,N_7591,N_7381);
nand U8002 (N_8002,N_7655,N_7302);
nand U8003 (N_8003,N_7305,N_7395);
nand U8004 (N_8004,N_7827,N_7782);
and U8005 (N_8005,N_7466,N_7756);
or U8006 (N_8006,N_7124,N_7257);
or U8007 (N_8007,N_7231,N_7248);
nor U8008 (N_8008,N_7706,N_7028);
or U8009 (N_8009,N_7375,N_7668);
nand U8010 (N_8010,N_7829,N_7673);
nand U8011 (N_8011,N_7404,N_7823);
or U8012 (N_8012,N_7414,N_7025);
nor U8013 (N_8013,N_7748,N_7621);
nor U8014 (N_8014,N_7749,N_7581);
nand U8015 (N_8015,N_7413,N_7502);
or U8016 (N_8016,N_7079,N_7891);
nor U8017 (N_8017,N_7491,N_7670);
nand U8018 (N_8018,N_7604,N_7196);
nor U8019 (N_8019,N_7134,N_7232);
xnor U8020 (N_8020,N_7901,N_7968);
nand U8021 (N_8021,N_7431,N_7836);
nand U8022 (N_8022,N_7427,N_7315);
and U8023 (N_8023,N_7443,N_7368);
xnor U8024 (N_8024,N_7189,N_7695);
nand U8025 (N_8025,N_7721,N_7486);
nand U8026 (N_8026,N_7663,N_7826);
or U8027 (N_8027,N_7985,N_7720);
and U8028 (N_8028,N_7074,N_7037);
xor U8029 (N_8029,N_7547,N_7928);
nor U8030 (N_8030,N_7949,N_7813);
nand U8031 (N_8031,N_7109,N_7053);
nor U8032 (N_8032,N_7635,N_7878);
or U8033 (N_8033,N_7843,N_7336);
or U8034 (N_8034,N_7541,N_7816);
and U8035 (N_8035,N_7108,N_7538);
nand U8036 (N_8036,N_7871,N_7235);
or U8037 (N_8037,N_7275,N_7995);
or U8038 (N_8038,N_7849,N_7214);
xnor U8039 (N_8039,N_7952,N_7485);
nor U8040 (N_8040,N_7434,N_7613);
and U8041 (N_8041,N_7961,N_7210);
or U8042 (N_8042,N_7258,N_7910);
nand U8043 (N_8043,N_7505,N_7060);
nand U8044 (N_8044,N_7340,N_7701);
and U8045 (N_8045,N_7744,N_7306);
nor U8046 (N_8046,N_7153,N_7144);
nand U8047 (N_8047,N_7730,N_7239);
or U8048 (N_8048,N_7742,N_7441);
nand U8049 (N_8049,N_7941,N_7353);
and U8050 (N_8050,N_7372,N_7161);
xor U8051 (N_8051,N_7154,N_7810);
nand U8052 (N_8052,N_7379,N_7068);
and U8053 (N_8053,N_7927,N_7200);
or U8054 (N_8054,N_7295,N_7680);
or U8055 (N_8055,N_7298,N_7609);
nor U8056 (N_8056,N_7997,N_7128);
or U8057 (N_8057,N_7692,N_7796);
nand U8058 (N_8058,N_7082,N_7240);
and U8059 (N_8059,N_7480,N_7216);
or U8060 (N_8060,N_7640,N_7935);
nand U8061 (N_8061,N_7840,N_7360);
nand U8062 (N_8062,N_7634,N_7664);
or U8063 (N_8063,N_7030,N_7512);
nand U8064 (N_8064,N_7837,N_7533);
nand U8065 (N_8065,N_7960,N_7387);
xnor U8066 (N_8066,N_7100,N_7608);
nand U8067 (N_8067,N_7571,N_7758);
nand U8068 (N_8068,N_7909,N_7637);
or U8069 (N_8069,N_7435,N_7267);
nand U8070 (N_8070,N_7054,N_7081);
xor U8071 (N_8071,N_7430,N_7967);
nand U8072 (N_8072,N_7000,N_7033);
or U8073 (N_8073,N_7352,N_7553);
or U8074 (N_8074,N_7755,N_7204);
nand U8075 (N_8075,N_7982,N_7511);
nand U8076 (N_8076,N_7882,N_7069);
or U8077 (N_8077,N_7130,N_7363);
or U8078 (N_8078,N_7408,N_7019);
and U8079 (N_8079,N_7580,N_7078);
or U8080 (N_8080,N_7627,N_7099);
nor U8081 (N_8081,N_7133,N_7474);
nand U8082 (N_8082,N_7517,N_7510);
nand U8083 (N_8083,N_7316,N_7654);
nand U8084 (N_8084,N_7661,N_7606);
nand U8085 (N_8085,N_7051,N_7162);
or U8086 (N_8086,N_7278,N_7526);
nor U8087 (N_8087,N_7531,N_7650);
and U8088 (N_8088,N_7179,N_7209);
or U8089 (N_8089,N_7243,N_7999);
xor U8090 (N_8090,N_7217,N_7550);
and U8091 (N_8091,N_7897,N_7940);
or U8092 (N_8092,N_7681,N_7065);
nor U8093 (N_8093,N_7432,N_7539);
nand U8094 (N_8094,N_7147,N_7064);
nor U8095 (N_8095,N_7947,N_7605);
nor U8096 (N_8096,N_7975,N_7679);
nand U8097 (N_8097,N_7088,N_7333);
xnor U8098 (N_8098,N_7097,N_7715);
and U8099 (N_8099,N_7981,N_7921);
nand U8100 (N_8100,N_7791,N_7788);
xnor U8101 (N_8101,N_7471,N_7991);
nand U8102 (N_8102,N_7260,N_7419);
nand U8103 (N_8103,N_7906,N_7058);
and U8104 (N_8104,N_7366,N_7215);
xnor U8105 (N_8105,N_7916,N_7674);
and U8106 (N_8106,N_7031,N_7197);
or U8107 (N_8107,N_7032,N_7672);
xnor U8108 (N_8108,N_7345,N_7804);
xnor U8109 (N_8109,N_7318,N_7422);
xnor U8110 (N_8110,N_7190,N_7610);
and U8111 (N_8111,N_7175,N_7966);
or U8112 (N_8112,N_7176,N_7020);
xor U8113 (N_8113,N_7980,N_7855);
nand U8114 (N_8114,N_7726,N_7898);
xor U8115 (N_8115,N_7457,N_7439);
nor U8116 (N_8116,N_7110,N_7561);
nor U8117 (N_8117,N_7396,N_7022);
nor U8118 (N_8118,N_7518,N_7202);
xor U8119 (N_8119,N_7743,N_7090);
nand U8120 (N_8120,N_7957,N_7631);
xor U8121 (N_8121,N_7467,N_7818);
or U8122 (N_8122,N_7135,N_7753);
nor U8123 (N_8123,N_7630,N_7913);
and U8124 (N_8124,N_7310,N_7174);
or U8125 (N_8125,N_7713,N_7639);
nand U8126 (N_8126,N_7040,N_7993);
nor U8127 (N_8127,N_7436,N_7010);
xnor U8128 (N_8128,N_7005,N_7615);
nor U8129 (N_8129,N_7955,N_7114);
or U8130 (N_8130,N_7814,N_7208);
xnor U8131 (N_8131,N_7786,N_7218);
nand U8132 (N_8132,N_7475,N_7567);
nor U8133 (N_8133,N_7867,N_7455);
nor U8134 (N_8134,N_7568,N_7973);
nand U8135 (N_8135,N_7905,N_7309);
or U8136 (N_8136,N_7223,N_7537);
xnor U8137 (N_8137,N_7164,N_7481);
nand U8138 (N_8138,N_7798,N_7984);
and U8139 (N_8139,N_7833,N_7647);
nor U8140 (N_8140,N_7237,N_7464);
and U8141 (N_8141,N_7018,N_7771);
and U8142 (N_8142,N_7374,N_7719);
and U8143 (N_8143,N_7564,N_7091);
and U8144 (N_8144,N_7026,N_7596);
and U8145 (N_8145,N_7930,N_7902);
nor U8146 (N_8146,N_7354,N_7429);
nand U8147 (N_8147,N_7462,N_7657);
nor U8148 (N_8148,N_7041,N_7887);
xor U8149 (N_8149,N_7038,N_7712);
xor U8150 (N_8150,N_7762,N_7344);
and U8151 (N_8151,N_7899,N_7588);
nand U8152 (N_8152,N_7084,N_7582);
or U8153 (N_8153,N_7220,N_7625);
nand U8154 (N_8154,N_7401,N_7165);
or U8155 (N_8155,N_7769,N_7917);
nor U8156 (N_8156,N_7977,N_7280);
xnor U8157 (N_8157,N_7219,N_7250);
nor U8158 (N_8158,N_7183,N_7676);
and U8159 (N_8159,N_7983,N_7620);
and U8160 (N_8160,N_7272,N_7854);
nor U8161 (N_8161,N_7448,N_7076);
nor U8162 (N_8162,N_7566,N_7397);
nand U8163 (N_8163,N_7754,N_7382);
or U8164 (N_8164,N_7127,N_7346);
or U8165 (N_8165,N_7044,N_7407);
and U8166 (N_8166,N_7013,N_7888);
nand U8167 (N_8167,N_7492,N_7934);
nor U8168 (N_8168,N_7277,N_7416);
or U8169 (N_8169,N_7619,N_7884);
nand U8170 (N_8170,N_7875,N_7111);
xnor U8171 (N_8171,N_7385,N_7137);
and U8172 (N_8172,N_7781,N_7320);
xor U8173 (N_8173,N_7686,N_7299);
and U8174 (N_8174,N_7574,N_7483);
nand U8175 (N_8175,N_7528,N_7498);
nor U8176 (N_8176,N_7508,N_7711);
nand U8177 (N_8177,N_7349,N_7118);
nand U8178 (N_8178,N_7107,N_7314);
xnor U8179 (N_8179,N_7392,N_7131);
or U8180 (N_8180,N_7583,N_7002);
xor U8181 (N_8181,N_7168,N_7515);
xnor U8182 (N_8182,N_7113,N_7468);
and U8183 (N_8183,N_7872,N_7778);
nor U8184 (N_8184,N_7103,N_7722);
or U8185 (N_8185,N_7746,N_7367);
xnor U8186 (N_8186,N_7597,N_7115);
nand U8187 (N_8187,N_7045,N_7487);
and U8188 (N_8188,N_7188,N_7669);
and U8189 (N_8189,N_7181,N_7992);
or U8190 (N_8190,N_7834,N_7688);
nor U8191 (N_8191,N_7914,N_7546);
and U8192 (N_8192,N_7739,N_7645);
and U8193 (N_8193,N_7595,N_7159);
and U8194 (N_8194,N_7572,N_7766);
or U8195 (N_8195,N_7042,N_7251);
nand U8196 (N_8196,N_7536,N_7732);
nor U8197 (N_8197,N_7842,N_7009);
or U8198 (N_8198,N_7415,N_7924);
and U8199 (N_8199,N_7171,N_7911);
and U8200 (N_8200,N_7832,N_7281);
xor U8201 (N_8201,N_7029,N_7438);
or U8202 (N_8202,N_7342,N_7105);
xor U8203 (N_8203,N_7093,N_7417);
or U8204 (N_8204,N_7794,N_7723);
nor U8205 (N_8205,N_7555,N_7761);
nor U8206 (N_8206,N_7229,N_7007);
or U8207 (N_8207,N_7101,N_7021);
nor U8208 (N_8208,N_7760,N_7864);
or U8209 (N_8209,N_7501,N_7256);
nor U8210 (N_8210,N_7186,N_7643);
xnor U8211 (N_8211,N_7557,N_7365);
or U8212 (N_8212,N_7835,N_7141);
xnor U8213 (N_8213,N_7741,N_7425);
and U8214 (N_8214,N_7249,N_7612);
xnor U8215 (N_8215,N_7377,N_7587);
nor U8216 (N_8216,N_7184,N_7073);
and U8217 (N_8217,N_7907,N_7287);
nor U8218 (N_8218,N_7638,N_7389);
or U8219 (N_8219,N_7750,N_7851);
nor U8220 (N_8220,N_7230,N_7169);
xor U8221 (N_8221,N_7173,N_7912);
or U8222 (N_8222,N_7160,N_7540);
nand U8223 (N_8223,N_7323,N_7241);
xor U8224 (N_8224,N_7034,N_7759);
xnor U8225 (N_8225,N_7881,N_7187);
nor U8226 (N_8226,N_7974,N_7332);
nor U8227 (N_8227,N_7877,N_7954);
xor U8228 (N_8228,N_7611,N_7773);
nor U8229 (N_8229,N_7861,N_7452);
or U8230 (N_8230,N_7682,N_7560);
nor U8231 (N_8231,N_7733,N_7048);
or U8232 (N_8232,N_7312,N_7570);
xnor U8233 (N_8233,N_7433,N_7626);
nand U8234 (N_8234,N_7211,N_7055);
nand U8235 (N_8235,N_7805,N_7521);
nor U8236 (N_8236,N_7563,N_7378);
and U8237 (N_8237,N_7089,N_7482);
nor U8238 (N_8238,N_7112,N_7863);
nor U8239 (N_8239,N_7569,N_7710);
nor U8240 (N_8240,N_7070,N_7269);
and U8241 (N_8241,N_7494,N_7972);
nand U8242 (N_8242,N_7602,N_7558);
xnor U8243 (N_8243,N_7848,N_7338);
or U8244 (N_8244,N_7490,N_7789);
nand U8245 (N_8245,N_7283,N_7694);
xnor U8246 (N_8246,N_7503,N_7592);
or U8247 (N_8247,N_7347,N_7282);
and U8248 (N_8248,N_7227,N_7700);
or U8249 (N_8249,N_7166,N_7325);
xor U8250 (N_8250,N_7205,N_7117);
xnor U8251 (N_8251,N_7554,N_7327);
or U8252 (N_8252,N_7776,N_7406);
and U8253 (N_8253,N_7303,N_7775);
or U8254 (N_8254,N_7659,N_7932);
and U8255 (N_8255,N_7057,N_7268);
and U8256 (N_8256,N_7463,N_7262);
xnor U8257 (N_8257,N_7915,N_7129);
xnor U8258 (N_8258,N_7520,N_7524);
nand U8259 (N_8259,N_7527,N_7800);
xor U8260 (N_8260,N_7274,N_7270);
nor U8261 (N_8261,N_7601,N_7530);
nand U8262 (N_8262,N_7145,N_7203);
xnor U8263 (N_8263,N_7092,N_7472);
or U8264 (N_8264,N_7535,N_7850);
nand U8265 (N_8265,N_7194,N_7066);
xor U8266 (N_8266,N_7138,N_7976);
or U8267 (N_8267,N_7224,N_7576);
and U8268 (N_8268,N_7459,N_7445);
and U8269 (N_8269,N_7324,N_7649);
xor U8270 (N_8270,N_7265,N_7437);
and U8271 (N_8271,N_7987,N_7326);
nor U8272 (N_8272,N_7087,N_7370);
and U8273 (N_8273,N_7962,N_7933);
xnor U8274 (N_8274,N_7618,N_7542);
or U8275 (N_8275,N_7357,N_7461);
and U8276 (N_8276,N_7290,N_7736);
and U8277 (N_8277,N_7157,N_7506);
xor U8278 (N_8278,N_7622,N_7691);
nand U8279 (N_8279,N_7651,N_7361);
xnor U8280 (N_8280,N_7399,N_7390);
or U8281 (N_8281,N_7096,N_7644);
or U8282 (N_8282,N_7683,N_7348);
or U8283 (N_8283,N_7291,N_7543);
nor U8284 (N_8284,N_7628,N_7125);
or U8285 (N_8285,N_7255,N_7892);
xnor U8286 (N_8286,N_7737,N_7132);
or U8287 (N_8287,N_7499,N_7339);
nor U8288 (N_8288,N_7938,N_7920);
xor U8289 (N_8289,N_7095,N_7411);
or U8290 (N_8290,N_7388,N_7319);
and U8291 (N_8291,N_7321,N_7085);
nor U8292 (N_8292,N_7684,N_7446);
and U8293 (N_8293,N_7516,N_7246);
and U8294 (N_8294,N_7945,N_7793);
or U8295 (N_8295,N_7971,N_7594);
nor U8296 (N_8296,N_7412,N_7895);
nor U8297 (N_8297,N_7696,N_7247);
or U8298 (N_8298,N_7136,N_7394);
and U8299 (N_8299,N_7293,N_7155);
or U8300 (N_8300,N_7629,N_7725);
nor U8301 (N_8301,N_7802,N_7104);
and U8302 (N_8302,N_7534,N_7192);
and U8303 (N_8303,N_7213,N_7106);
nor U8304 (N_8304,N_7652,N_7690);
or U8305 (N_8305,N_7146,N_7469);
or U8306 (N_8306,N_7944,N_7244);
nand U8307 (N_8307,N_7350,N_7328);
xor U8308 (N_8308,N_7820,N_7641);
and U8309 (N_8309,N_7261,N_7886);
and U8310 (N_8310,N_7885,N_7442);
or U8311 (N_8311,N_7708,N_7440);
nor U8312 (N_8312,N_7740,N_7685);
nand U8313 (N_8313,N_7236,N_7838);
nand U8314 (N_8314,N_7986,N_7552);
or U8315 (N_8315,N_7573,N_7632);
nand U8316 (N_8316,N_7918,N_7263);
nand U8317 (N_8317,N_7825,N_7799);
or U8318 (N_8318,N_7121,N_7273);
nand U8319 (N_8319,N_7598,N_7853);
xnor U8320 (N_8320,N_7012,N_7059);
or U8321 (N_8321,N_7116,N_7286);
or U8322 (N_8322,N_7653,N_7646);
and U8323 (N_8323,N_7772,N_7948);
and U8324 (N_8324,N_7364,N_7102);
or U8325 (N_8325,N_7167,N_7617);
nor U8326 (N_8326,N_7790,N_7083);
nor U8327 (N_8327,N_7815,N_7035);
or U8328 (N_8328,N_7784,N_7678);
nor U8329 (N_8329,N_7925,N_7479);
or U8330 (N_8330,N_7424,N_7666);
nor U8331 (N_8331,N_7509,N_7234);
xor U8332 (N_8332,N_7774,N_7964);
nand U8333 (N_8333,N_7391,N_7063);
nor U8334 (N_8334,N_7857,N_7585);
or U8335 (N_8335,N_7279,N_7812);
nand U8336 (N_8336,N_7264,N_7050);
and U8337 (N_8337,N_7398,N_7845);
and U8338 (N_8338,N_7454,N_7824);
and U8339 (N_8339,N_7195,N_7317);
nor U8340 (N_8340,N_7809,N_7006);
or U8341 (N_8341,N_7797,N_7225);
or U8342 (N_8342,N_7470,N_7151);
xor U8343 (N_8343,N_7817,N_7787);
nand U8344 (N_8344,N_7900,N_7728);
nand U8345 (N_8345,N_7926,N_7525);
xnor U8346 (N_8346,N_7245,N_7359);
xnor U8347 (N_8347,N_7889,N_7052);
or U8348 (N_8348,N_7942,N_7697);
or U8349 (N_8349,N_7072,N_7616);
nor U8350 (N_8350,N_7946,N_7636);
and U8351 (N_8351,N_7376,N_7514);
xor U8352 (N_8352,N_7094,N_7329);
nand U8353 (N_8353,N_7599,N_7831);
nand U8354 (N_8354,N_7017,N_7577);
or U8355 (N_8355,N_7402,N_7497);
nor U8356 (N_8356,N_7768,N_7705);
and U8357 (N_8357,N_7201,N_7075);
nor U8358 (N_8358,N_7830,N_7709);
and U8359 (N_8359,N_7170,N_7355);
or U8360 (N_8360,N_7633,N_7400);
xnor U8361 (N_8361,N_7767,N_7667);
and U8362 (N_8362,N_7988,N_7969);
and U8363 (N_8363,N_7142,N_7004);
and U8364 (N_8364,N_7562,N_7228);
nand U8365 (N_8365,N_7724,N_7529);
xor U8366 (N_8366,N_7098,N_7575);
xor U8367 (N_8367,N_7671,N_7253);
xnor U8368 (N_8368,N_7545,N_7801);
nand U8369 (N_8369,N_7254,N_7893);
and U8370 (N_8370,N_7420,N_7143);
nor U8371 (N_8371,N_7222,N_7036);
nand U8372 (N_8372,N_7806,N_7308);
nor U8373 (N_8373,N_7233,N_7660);
and U8374 (N_8374,N_7177,N_7334);
xnor U8375 (N_8375,N_7642,N_7819);
nand U8376 (N_8376,N_7444,N_7873);
nor U8377 (N_8377,N_7858,N_7047);
nor U8378 (N_8378,N_7880,N_7702);
and U8379 (N_8379,N_7297,N_7965);
xor U8380 (N_8380,N_7285,N_7731);
or U8381 (N_8381,N_7453,N_7311);
nor U8382 (N_8382,N_7123,N_7484);
nand U8383 (N_8383,N_7792,N_7500);
or U8384 (N_8384,N_7386,N_7996);
nor U8385 (N_8385,N_7903,N_7939);
nor U8386 (N_8386,N_7959,N_7276);
and U8387 (N_8387,N_7665,N_7008);
and U8388 (N_8388,N_7846,N_7745);
and U8389 (N_8389,N_7590,N_7623);
nand U8390 (N_8390,N_7953,N_7296);
nor U8391 (N_8391,N_7931,N_7752);
and U8392 (N_8392,N_7238,N_7341);
xor U8393 (N_8393,N_7313,N_7689);
nand U8394 (N_8394,N_7699,N_7504);
and U8395 (N_8395,N_7062,N_7380);
xnor U8396 (N_8396,N_7693,N_7152);
xor U8397 (N_8397,N_7199,N_7158);
and U8398 (N_8398,N_7191,N_7207);
nor U8399 (N_8399,N_7393,N_7777);
nor U8400 (N_8400,N_7067,N_7593);
xor U8401 (N_8401,N_7304,N_7292);
nand U8402 (N_8402,N_7140,N_7356);
nor U8403 (N_8403,N_7016,N_7765);
and U8404 (N_8404,N_7879,N_7783);
nand U8405 (N_8405,N_7023,N_7493);
nor U8406 (N_8406,N_7704,N_7727);
xor U8407 (N_8407,N_7841,N_7936);
xor U8408 (N_8408,N_7757,N_7549);
nand U8409 (N_8409,N_7738,N_7923);
nand U8410 (N_8410,N_7001,N_7011);
nand U8411 (N_8411,N_7478,N_7330);
and U8412 (N_8412,N_7015,N_7584);
and U8413 (N_8413,N_7014,N_7770);
or U8414 (N_8414,N_7149,N_7148);
nand U8415 (N_8415,N_7271,N_7603);
nand U8416 (N_8416,N_7734,N_7077);
xnor U8417 (N_8417,N_7922,N_7351);
nand U8418 (N_8418,N_7126,N_7476);
nor U8419 (N_8419,N_7779,N_7495);
nor U8420 (N_8420,N_7465,N_7300);
and U8421 (N_8421,N_7206,N_7156);
nand U8422 (N_8422,N_7747,N_7556);
and U8423 (N_8423,N_7894,N_7428);
or U8424 (N_8424,N_7859,N_7384);
or U8425 (N_8425,N_7221,N_7648);
nand U8426 (N_8426,N_7703,N_7822);
nor U8427 (N_8427,N_7658,N_7288);
xor U8428 (N_8428,N_7343,N_7865);
nor U8429 (N_8429,N_7410,N_7551);
nand U8430 (N_8430,N_7226,N_7523);
and U8431 (N_8431,N_7544,N_7828);
nand U8432 (N_8432,N_7994,N_7335);
nand U8433 (N_8433,N_7139,N_7716);
or U8434 (N_8434,N_7839,N_7473);
nor U8435 (N_8435,N_7447,N_7337);
or U8436 (N_8436,N_7056,N_7607);
and U8437 (N_8437,N_7426,N_7450);
or U8438 (N_8438,N_7908,N_7212);
nor U8439 (N_8439,N_7120,N_7003);
or U8440 (N_8440,N_7198,N_7373);
xnor U8441 (N_8441,N_7943,N_7458);
and U8442 (N_8442,N_7489,N_7252);
or U8443 (N_8443,N_7751,N_7624);
nor U8444 (N_8444,N_7869,N_7718);
and U8445 (N_8445,N_7405,N_7043);
xor U8446 (N_8446,N_7423,N_7958);
or U8447 (N_8447,N_7714,N_7662);
and U8448 (N_8448,N_7507,N_7027);
nand U8449 (N_8449,N_7856,N_7477);
xor U8450 (N_8450,N_7795,N_7409);
nor U8451 (N_8451,N_7488,N_7513);
xor U8452 (N_8452,N_7532,N_7785);
nand U8453 (N_8453,N_7421,N_7970);
and U8454 (N_8454,N_7919,N_7519);
nor U8455 (N_8455,N_7956,N_7565);
xnor U8456 (N_8456,N_7086,N_7821);
and U8457 (N_8457,N_7950,N_7687);
or U8458 (N_8458,N_7866,N_7456);
nor U8459 (N_8459,N_7371,N_7698);
nand U8460 (N_8460,N_7451,N_7049);
nor U8461 (N_8461,N_7522,N_7811);
and U8462 (N_8462,N_7808,N_7046);
nor U8463 (N_8463,N_7847,N_7182);
nand U8464 (N_8464,N_7496,N_7600);
nand U8465 (N_8465,N_7862,N_7331);
and U8466 (N_8466,N_7266,N_7193);
nor U8467 (N_8467,N_7071,N_7735);
or U8468 (N_8468,N_7729,N_7870);
or U8469 (N_8469,N_7172,N_7807);
nor U8470 (N_8470,N_7929,N_7119);
nand U8471 (N_8471,N_7242,N_7579);
nand U8472 (N_8472,N_7763,N_7061);
xor U8473 (N_8473,N_7874,N_7852);
nor U8474 (N_8474,N_7301,N_7369);
nor U8475 (N_8475,N_7998,N_7868);
or U8476 (N_8476,N_7362,N_7978);
xnor U8477 (N_8477,N_7284,N_7860);
or U8478 (N_8478,N_7039,N_7178);
or U8479 (N_8479,N_7289,N_7896);
nor U8480 (N_8480,N_7559,N_7656);
nor U8481 (N_8481,N_7990,N_7675);
nor U8482 (N_8482,N_7979,N_7307);
and U8483 (N_8483,N_7403,N_7150);
nor U8484 (N_8484,N_7951,N_7180);
nor U8485 (N_8485,N_7963,N_7989);
and U8486 (N_8486,N_7803,N_7122);
nand U8487 (N_8487,N_7904,N_7844);
and U8488 (N_8488,N_7707,N_7764);
or U8489 (N_8489,N_7677,N_7586);
or U8490 (N_8490,N_7418,N_7876);
nand U8491 (N_8491,N_7294,N_7589);
or U8492 (N_8492,N_7883,N_7185);
or U8493 (N_8493,N_7890,N_7163);
or U8494 (N_8494,N_7024,N_7548);
and U8495 (N_8495,N_7614,N_7358);
and U8496 (N_8496,N_7460,N_7383);
or U8497 (N_8497,N_7259,N_7080);
or U8498 (N_8498,N_7780,N_7937);
or U8499 (N_8499,N_7449,N_7578);
or U8500 (N_8500,N_7017,N_7615);
nand U8501 (N_8501,N_7602,N_7403);
nor U8502 (N_8502,N_7797,N_7879);
or U8503 (N_8503,N_7812,N_7723);
and U8504 (N_8504,N_7183,N_7320);
nand U8505 (N_8505,N_7861,N_7899);
xnor U8506 (N_8506,N_7058,N_7778);
nor U8507 (N_8507,N_7029,N_7624);
xnor U8508 (N_8508,N_7151,N_7020);
or U8509 (N_8509,N_7715,N_7031);
and U8510 (N_8510,N_7925,N_7165);
xor U8511 (N_8511,N_7257,N_7076);
or U8512 (N_8512,N_7578,N_7805);
nand U8513 (N_8513,N_7078,N_7758);
nand U8514 (N_8514,N_7352,N_7747);
or U8515 (N_8515,N_7224,N_7420);
and U8516 (N_8516,N_7394,N_7340);
nand U8517 (N_8517,N_7844,N_7550);
and U8518 (N_8518,N_7640,N_7576);
and U8519 (N_8519,N_7094,N_7940);
nor U8520 (N_8520,N_7683,N_7061);
nand U8521 (N_8521,N_7477,N_7556);
nor U8522 (N_8522,N_7676,N_7974);
or U8523 (N_8523,N_7555,N_7797);
and U8524 (N_8524,N_7377,N_7097);
nor U8525 (N_8525,N_7100,N_7758);
or U8526 (N_8526,N_7710,N_7803);
or U8527 (N_8527,N_7613,N_7518);
or U8528 (N_8528,N_7824,N_7261);
nor U8529 (N_8529,N_7819,N_7080);
or U8530 (N_8530,N_7315,N_7894);
xor U8531 (N_8531,N_7361,N_7393);
nor U8532 (N_8532,N_7983,N_7787);
xnor U8533 (N_8533,N_7674,N_7523);
and U8534 (N_8534,N_7112,N_7617);
or U8535 (N_8535,N_7835,N_7693);
and U8536 (N_8536,N_7440,N_7084);
or U8537 (N_8537,N_7114,N_7815);
nand U8538 (N_8538,N_7454,N_7081);
or U8539 (N_8539,N_7089,N_7552);
nor U8540 (N_8540,N_7766,N_7600);
nor U8541 (N_8541,N_7795,N_7579);
and U8542 (N_8542,N_7020,N_7773);
or U8543 (N_8543,N_7104,N_7884);
and U8544 (N_8544,N_7389,N_7166);
nor U8545 (N_8545,N_7518,N_7583);
or U8546 (N_8546,N_7500,N_7605);
nor U8547 (N_8547,N_7161,N_7129);
nor U8548 (N_8548,N_7168,N_7479);
xor U8549 (N_8549,N_7610,N_7896);
or U8550 (N_8550,N_7414,N_7033);
xnor U8551 (N_8551,N_7563,N_7553);
or U8552 (N_8552,N_7370,N_7354);
and U8553 (N_8553,N_7531,N_7612);
nand U8554 (N_8554,N_7651,N_7658);
and U8555 (N_8555,N_7097,N_7515);
nand U8556 (N_8556,N_7535,N_7467);
nand U8557 (N_8557,N_7463,N_7909);
or U8558 (N_8558,N_7070,N_7000);
nand U8559 (N_8559,N_7461,N_7324);
and U8560 (N_8560,N_7798,N_7749);
or U8561 (N_8561,N_7583,N_7158);
nand U8562 (N_8562,N_7160,N_7259);
and U8563 (N_8563,N_7130,N_7998);
nand U8564 (N_8564,N_7642,N_7980);
xnor U8565 (N_8565,N_7595,N_7594);
or U8566 (N_8566,N_7535,N_7328);
nand U8567 (N_8567,N_7651,N_7985);
or U8568 (N_8568,N_7164,N_7025);
and U8569 (N_8569,N_7108,N_7328);
and U8570 (N_8570,N_7963,N_7361);
xnor U8571 (N_8571,N_7340,N_7473);
nand U8572 (N_8572,N_7288,N_7143);
or U8573 (N_8573,N_7997,N_7551);
and U8574 (N_8574,N_7182,N_7259);
or U8575 (N_8575,N_7990,N_7459);
or U8576 (N_8576,N_7213,N_7620);
or U8577 (N_8577,N_7664,N_7423);
and U8578 (N_8578,N_7843,N_7231);
nand U8579 (N_8579,N_7093,N_7696);
xnor U8580 (N_8580,N_7084,N_7882);
or U8581 (N_8581,N_7440,N_7685);
or U8582 (N_8582,N_7904,N_7114);
nand U8583 (N_8583,N_7315,N_7194);
xnor U8584 (N_8584,N_7946,N_7835);
xor U8585 (N_8585,N_7447,N_7622);
or U8586 (N_8586,N_7004,N_7112);
nor U8587 (N_8587,N_7667,N_7734);
or U8588 (N_8588,N_7837,N_7762);
xor U8589 (N_8589,N_7067,N_7069);
or U8590 (N_8590,N_7728,N_7329);
or U8591 (N_8591,N_7424,N_7590);
xor U8592 (N_8592,N_7614,N_7980);
nand U8593 (N_8593,N_7105,N_7040);
and U8594 (N_8594,N_7781,N_7783);
and U8595 (N_8595,N_7289,N_7806);
xor U8596 (N_8596,N_7493,N_7220);
or U8597 (N_8597,N_7758,N_7811);
nand U8598 (N_8598,N_7733,N_7675);
xnor U8599 (N_8599,N_7886,N_7838);
and U8600 (N_8600,N_7359,N_7341);
xnor U8601 (N_8601,N_7796,N_7546);
xor U8602 (N_8602,N_7272,N_7985);
nand U8603 (N_8603,N_7443,N_7469);
xor U8604 (N_8604,N_7252,N_7972);
nand U8605 (N_8605,N_7292,N_7921);
or U8606 (N_8606,N_7082,N_7164);
nor U8607 (N_8607,N_7639,N_7522);
and U8608 (N_8608,N_7364,N_7039);
xnor U8609 (N_8609,N_7021,N_7194);
nand U8610 (N_8610,N_7487,N_7872);
nand U8611 (N_8611,N_7824,N_7740);
and U8612 (N_8612,N_7703,N_7341);
nand U8613 (N_8613,N_7990,N_7543);
nor U8614 (N_8614,N_7099,N_7003);
or U8615 (N_8615,N_7978,N_7079);
xnor U8616 (N_8616,N_7142,N_7425);
and U8617 (N_8617,N_7962,N_7754);
nor U8618 (N_8618,N_7712,N_7789);
xnor U8619 (N_8619,N_7055,N_7137);
nor U8620 (N_8620,N_7404,N_7534);
nor U8621 (N_8621,N_7161,N_7997);
nand U8622 (N_8622,N_7016,N_7161);
or U8623 (N_8623,N_7926,N_7507);
and U8624 (N_8624,N_7741,N_7057);
and U8625 (N_8625,N_7821,N_7455);
nor U8626 (N_8626,N_7436,N_7865);
nand U8627 (N_8627,N_7303,N_7519);
xnor U8628 (N_8628,N_7093,N_7127);
or U8629 (N_8629,N_7910,N_7883);
and U8630 (N_8630,N_7868,N_7389);
nand U8631 (N_8631,N_7291,N_7393);
nand U8632 (N_8632,N_7779,N_7970);
and U8633 (N_8633,N_7783,N_7417);
nand U8634 (N_8634,N_7009,N_7211);
nor U8635 (N_8635,N_7007,N_7525);
and U8636 (N_8636,N_7057,N_7998);
xnor U8637 (N_8637,N_7547,N_7341);
and U8638 (N_8638,N_7916,N_7707);
and U8639 (N_8639,N_7065,N_7576);
nand U8640 (N_8640,N_7870,N_7769);
nor U8641 (N_8641,N_7449,N_7129);
nor U8642 (N_8642,N_7213,N_7662);
or U8643 (N_8643,N_7498,N_7182);
nor U8644 (N_8644,N_7024,N_7196);
or U8645 (N_8645,N_7230,N_7180);
nor U8646 (N_8646,N_7422,N_7310);
nand U8647 (N_8647,N_7574,N_7510);
nor U8648 (N_8648,N_7994,N_7876);
xnor U8649 (N_8649,N_7595,N_7561);
or U8650 (N_8650,N_7193,N_7239);
nor U8651 (N_8651,N_7756,N_7736);
nand U8652 (N_8652,N_7377,N_7438);
nor U8653 (N_8653,N_7896,N_7611);
xor U8654 (N_8654,N_7460,N_7393);
or U8655 (N_8655,N_7243,N_7718);
nor U8656 (N_8656,N_7908,N_7378);
nand U8657 (N_8657,N_7055,N_7063);
nand U8658 (N_8658,N_7267,N_7931);
nand U8659 (N_8659,N_7650,N_7642);
and U8660 (N_8660,N_7808,N_7199);
nor U8661 (N_8661,N_7057,N_7069);
nand U8662 (N_8662,N_7910,N_7731);
nand U8663 (N_8663,N_7977,N_7537);
xnor U8664 (N_8664,N_7703,N_7102);
nor U8665 (N_8665,N_7601,N_7739);
xnor U8666 (N_8666,N_7766,N_7723);
xnor U8667 (N_8667,N_7359,N_7093);
or U8668 (N_8668,N_7536,N_7247);
nor U8669 (N_8669,N_7044,N_7204);
and U8670 (N_8670,N_7919,N_7397);
nor U8671 (N_8671,N_7130,N_7044);
or U8672 (N_8672,N_7783,N_7283);
and U8673 (N_8673,N_7268,N_7986);
nor U8674 (N_8674,N_7697,N_7512);
xor U8675 (N_8675,N_7089,N_7058);
nand U8676 (N_8676,N_7357,N_7603);
nor U8677 (N_8677,N_7011,N_7087);
nand U8678 (N_8678,N_7993,N_7028);
nand U8679 (N_8679,N_7679,N_7805);
and U8680 (N_8680,N_7045,N_7603);
or U8681 (N_8681,N_7479,N_7094);
nor U8682 (N_8682,N_7723,N_7565);
or U8683 (N_8683,N_7427,N_7656);
and U8684 (N_8684,N_7541,N_7542);
nor U8685 (N_8685,N_7642,N_7875);
nor U8686 (N_8686,N_7713,N_7527);
or U8687 (N_8687,N_7391,N_7169);
or U8688 (N_8688,N_7429,N_7663);
and U8689 (N_8689,N_7759,N_7123);
nand U8690 (N_8690,N_7136,N_7329);
xor U8691 (N_8691,N_7162,N_7783);
nor U8692 (N_8692,N_7750,N_7592);
or U8693 (N_8693,N_7683,N_7571);
nor U8694 (N_8694,N_7824,N_7335);
or U8695 (N_8695,N_7301,N_7522);
and U8696 (N_8696,N_7960,N_7937);
and U8697 (N_8697,N_7436,N_7115);
or U8698 (N_8698,N_7970,N_7930);
and U8699 (N_8699,N_7299,N_7959);
xor U8700 (N_8700,N_7111,N_7114);
nor U8701 (N_8701,N_7400,N_7547);
and U8702 (N_8702,N_7214,N_7019);
nand U8703 (N_8703,N_7798,N_7796);
nand U8704 (N_8704,N_7634,N_7828);
and U8705 (N_8705,N_7492,N_7487);
or U8706 (N_8706,N_7111,N_7584);
nor U8707 (N_8707,N_7367,N_7253);
xor U8708 (N_8708,N_7948,N_7136);
xnor U8709 (N_8709,N_7360,N_7882);
xor U8710 (N_8710,N_7618,N_7030);
xor U8711 (N_8711,N_7631,N_7468);
nor U8712 (N_8712,N_7330,N_7337);
and U8713 (N_8713,N_7364,N_7176);
nand U8714 (N_8714,N_7510,N_7370);
and U8715 (N_8715,N_7785,N_7263);
xor U8716 (N_8716,N_7364,N_7962);
xor U8717 (N_8717,N_7643,N_7984);
and U8718 (N_8718,N_7049,N_7483);
and U8719 (N_8719,N_7617,N_7966);
nand U8720 (N_8720,N_7281,N_7363);
nand U8721 (N_8721,N_7271,N_7207);
or U8722 (N_8722,N_7374,N_7583);
and U8723 (N_8723,N_7183,N_7809);
xor U8724 (N_8724,N_7065,N_7277);
xnor U8725 (N_8725,N_7497,N_7224);
or U8726 (N_8726,N_7795,N_7144);
and U8727 (N_8727,N_7498,N_7895);
or U8728 (N_8728,N_7674,N_7976);
xor U8729 (N_8729,N_7471,N_7162);
xnor U8730 (N_8730,N_7865,N_7797);
xor U8731 (N_8731,N_7626,N_7662);
or U8732 (N_8732,N_7820,N_7609);
xor U8733 (N_8733,N_7060,N_7309);
nor U8734 (N_8734,N_7904,N_7994);
nand U8735 (N_8735,N_7749,N_7263);
xor U8736 (N_8736,N_7465,N_7459);
nor U8737 (N_8737,N_7137,N_7226);
or U8738 (N_8738,N_7726,N_7163);
nand U8739 (N_8739,N_7675,N_7776);
nor U8740 (N_8740,N_7127,N_7597);
or U8741 (N_8741,N_7036,N_7936);
and U8742 (N_8742,N_7037,N_7484);
or U8743 (N_8743,N_7973,N_7232);
or U8744 (N_8744,N_7270,N_7939);
xor U8745 (N_8745,N_7720,N_7725);
or U8746 (N_8746,N_7115,N_7277);
xor U8747 (N_8747,N_7542,N_7013);
and U8748 (N_8748,N_7507,N_7135);
xnor U8749 (N_8749,N_7263,N_7237);
and U8750 (N_8750,N_7309,N_7691);
or U8751 (N_8751,N_7428,N_7008);
or U8752 (N_8752,N_7724,N_7607);
xnor U8753 (N_8753,N_7323,N_7468);
nor U8754 (N_8754,N_7434,N_7628);
or U8755 (N_8755,N_7590,N_7428);
nor U8756 (N_8756,N_7698,N_7162);
and U8757 (N_8757,N_7028,N_7603);
nor U8758 (N_8758,N_7525,N_7357);
or U8759 (N_8759,N_7628,N_7655);
or U8760 (N_8760,N_7044,N_7783);
and U8761 (N_8761,N_7100,N_7982);
xnor U8762 (N_8762,N_7731,N_7138);
or U8763 (N_8763,N_7375,N_7777);
nor U8764 (N_8764,N_7784,N_7723);
xor U8765 (N_8765,N_7179,N_7068);
xnor U8766 (N_8766,N_7198,N_7503);
or U8767 (N_8767,N_7082,N_7476);
nor U8768 (N_8768,N_7738,N_7371);
nand U8769 (N_8769,N_7125,N_7752);
nand U8770 (N_8770,N_7102,N_7593);
and U8771 (N_8771,N_7810,N_7940);
xor U8772 (N_8772,N_7072,N_7680);
xnor U8773 (N_8773,N_7171,N_7412);
nand U8774 (N_8774,N_7171,N_7561);
and U8775 (N_8775,N_7823,N_7612);
nor U8776 (N_8776,N_7613,N_7081);
xnor U8777 (N_8777,N_7102,N_7709);
and U8778 (N_8778,N_7893,N_7208);
or U8779 (N_8779,N_7453,N_7438);
nand U8780 (N_8780,N_7479,N_7601);
and U8781 (N_8781,N_7180,N_7741);
nand U8782 (N_8782,N_7662,N_7556);
xnor U8783 (N_8783,N_7798,N_7443);
or U8784 (N_8784,N_7700,N_7310);
xor U8785 (N_8785,N_7029,N_7318);
and U8786 (N_8786,N_7320,N_7039);
nand U8787 (N_8787,N_7412,N_7827);
nor U8788 (N_8788,N_7312,N_7785);
nor U8789 (N_8789,N_7700,N_7006);
nor U8790 (N_8790,N_7558,N_7026);
or U8791 (N_8791,N_7764,N_7319);
xor U8792 (N_8792,N_7932,N_7153);
nor U8793 (N_8793,N_7900,N_7972);
and U8794 (N_8794,N_7012,N_7424);
and U8795 (N_8795,N_7939,N_7482);
and U8796 (N_8796,N_7166,N_7604);
nand U8797 (N_8797,N_7981,N_7321);
or U8798 (N_8798,N_7552,N_7601);
nor U8799 (N_8799,N_7711,N_7273);
or U8800 (N_8800,N_7777,N_7164);
xnor U8801 (N_8801,N_7183,N_7272);
nand U8802 (N_8802,N_7141,N_7296);
nor U8803 (N_8803,N_7280,N_7558);
nor U8804 (N_8804,N_7189,N_7316);
nand U8805 (N_8805,N_7538,N_7387);
xnor U8806 (N_8806,N_7949,N_7936);
nand U8807 (N_8807,N_7245,N_7322);
and U8808 (N_8808,N_7240,N_7317);
and U8809 (N_8809,N_7713,N_7600);
or U8810 (N_8810,N_7775,N_7024);
and U8811 (N_8811,N_7473,N_7998);
nor U8812 (N_8812,N_7815,N_7758);
or U8813 (N_8813,N_7176,N_7679);
or U8814 (N_8814,N_7268,N_7571);
or U8815 (N_8815,N_7161,N_7943);
nand U8816 (N_8816,N_7274,N_7842);
nand U8817 (N_8817,N_7893,N_7579);
nor U8818 (N_8818,N_7913,N_7778);
or U8819 (N_8819,N_7596,N_7627);
nor U8820 (N_8820,N_7140,N_7013);
xor U8821 (N_8821,N_7332,N_7903);
or U8822 (N_8822,N_7047,N_7079);
xnor U8823 (N_8823,N_7669,N_7243);
or U8824 (N_8824,N_7690,N_7837);
or U8825 (N_8825,N_7092,N_7412);
xor U8826 (N_8826,N_7039,N_7370);
nor U8827 (N_8827,N_7646,N_7921);
and U8828 (N_8828,N_7314,N_7411);
nor U8829 (N_8829,N_7536,N_7606);
nand U8830 (N_8830,N_7154,N_7540);
nand U8831 (N_8831,N_7471,N_7789);
and U8832 (N_8832,N_7554,N_7929);
nand U8833 (N_8833,N_7240,N_7518);
and U8834 (N_8834,N_7737,N_7317);
nand U8835 (N_8835,N_7021,N_7036);
and U8836 (N_8836,N_7430,N_7495);
nand U8837 (N_8837,N_7144,N_7897);
xnor U8838 (N_8838,N_7942,N_7327);
nor U8839 (N_8839,N_7549,N_7243);
or U8840 (N_8840,N_7355,N_7478);
and U8841 (N_8841,N_7263,N_7310);
nand U8842 (N_8842,N_7687,N_7977);
nor U8843 (N_8843,N_7843,N_7827);
nand U8844 (N_8844,N_7175,N_7241);
nand U8845 (N_8845,N_7169,N_7934);
and U8846 (N_8846,N_7786,N_7844);
or U8847 (N_8847,N_7261,N_7312);
and U8848 (N_8848,N_7815,N_7136);
and U8849 (N_8849,N_7488,N_7041);
nor U8850 (N_8850,N_7715,N_7748);
nand U8851 (N_8851,N_7498,N_7671);
xor U8852 (N_8852,N_7931,N_7496);
xor U8853 (N_8853,N_7004,N_7621);
or U8854 (N_8854,N_7591,N_7625);
nor U8855 (N_8855,N_7810,N_7167);
xnor U8856 (N_8856,N_7696,N_7673);
nor U8857 (N_8857,N_7435,N_7830);
or U8858 (N_8858,N_7271,N_7262);
nand U8859 (N_8859,N_7778,N_7301);
nand U8860 (N_8860,N_7544,N_7212);
or U8861 (N_8861,N_7951,N_7946);
and U8862 (N_8862,N_7468,N_7035);
nand U8863 (N_8863,N_7466,N_7714);
nand U8864 (N_8864,N_7036,N_7385);
or U8865 (N_8865,N_7184,N_7903);
nand U8866 (N_8866,N_7650,N_7952);
nand U8867 (N_8867,N_7290,N_7203);
and U8868 (N_8868,N_7581,N_7483);
nand U8869 (N_8869,N_7049,N_7061);
nand U8870 (N_8870,N_7612,N_7254);
nor U8871 (N_8871,N_7525,N_7047);
nand U8872 (N_8872,N_7406,N_7971);
nand U8873 (N_8873,N_7265,N_7815);
nand U8874 (N_8874,N_7311,N_7743);
nand U8875 (N_8875,N_7781,N_7088);
xnor U8876 (N_8876,N_7199,N_7654);
or U8877 (N_8877,N_7735,N_7277);
xnor U8878 (N_8878,N_7674,N_7929);
or U8879 (N_8879,N_7808,N_7946);
or U8880 (N_8880,N_7849,N_7662);
and U8881 (N_8881,N_7328,N_7013);
xor U8882 (N_8882,N_7888,N_7684);
xnor U8883 (N_8883,N_7730,N_7748);
or U8884 (N_8884,N_7224,N_7167);
and U8885 (N_8885,N_7518,N_7172);
nand U8886 (N_8886,N_7484,N_7977);
nand U8887 (N_8887,N_7424,N_7334);
or U8888 (N_8888,N_7652,N_7228);
nor U8889 (N_8889,N_7613,N_7591);
nor U8890 (N_8890,N_7925,N_7498);
nor U8891 (N_8891,N_7702,N_7877);
xnor U8892 (N_8892,N_7155,N_7242);
and U8893 (N_8893,N_7056,N_7732);
nand U8894 (N_8894,N_7396,N_7332);
nor U8895 (N_8895,N_7388,N_7315);
or U8896 (N_8896,N_7434,N_7726);
and U8897 (N_8897,N_7537,N_7761);
and U8898 (N_8898,N_7586,N_7810);
xnor U8899 (N_8899,N_7692,N_7529);
or U8900 (N_8900,N_7395,N_7527);
nor U8901 (N_8901,N_7262,N_7378);
or U8902 (N_8902,N_7514,N_7701);
and U8903 (N_8903,N_7103,N_7374);
nor U8904 (N_8904,N_7520,N_7123);
nand U8905 (N_8905,N_7250,N_7258);
xnor U8906 (N_8906,N_7183,N_7094);
or U8907 (N_8907,N_7171,N_7991);
or U8908 (N_8908,N_7448,N_7775);
and U8909 (N_8909,N_7387,N_7094);
nor U8910 (N_8910,N_7716,N_7106);
nor U8911 (N_8911,N_7806,N_7279);
nor U8912 (N_8912,N_7391,N_7013);
xnor U8913 (N_8913,N_7669,N_7203);
xor U8914 (N_8914,N_7765,N_7761);
and U8915 (N_8915,N_7388,N_7889);
xor U8916 (N_8916,N_7184,N_7763);
xor U8917 (N_8917,N_7919,N_7076);
and U8918 (N_8918,N_7088,N_7707);
nand U8919 (N_8919,N_7653,N_7343);
xor U8920 (N_8920,N_7120,N_7579);
nand U8921 (N_8921,N_7662,N_7642);
and U8922 (N_8922,N_7982,N_7396);
nor U8923 (N_8923,N_7015,N_7473);
xor U8924 (N_8924,N_7022,N_7148);
and U8925 (N_8925,N_7648,N_7226);
and U8926 (N_8926,N_7964,N_7801);
nor U8927 (N_8927,N_7296,N_7635);
or U8928 (N_8928,N_7321,N_7489);
nor U8929 (N_8929,N_7808,N_7973);
xnor U8930 (N_8930,N_7448,N_7221);
xnor U8931 (N_8931,N_7844,N_7420);
nand U8932 (N_8932,N_7378,N_7770);
and U8933 (N_8933,N_7712,N_7970);
xnor U8934 (N_8934,N_7048,N_7362);
and U8935 (N_8935,N_7365,N_7747);
xnor U8936 (N_8936,N_7964,N_7458);
or U8937 (N_8937,N_7619,N_7980);
nand U8938 (N_8938,N_7083,N_7547);
or U8939 (N_8939,N_7050,N_7192);
or U8940 (N_8940,N_7633,N_7991);
and U8941 (N_8941,N_7829,N_7320);
nor U8942 (N_8942,N_7681,N_7010);
and U8943 (N_8943,N_7792,N_7129);
xnor U8944 (N_8944,N_7107,N_7458);
or U8945 (N_8945,N_7907,N_7839);
and U8946 (N_8946,N_7443,N_7459);
or U8947 (N_8947,N_7975,N_7033);
or U8948 (N_8948,N_7748,N_7783);
nor U8949 (N_8949,N_7128,N_7528);
or U8950 (N_8950,N_7963,N_7801);
xnor U8951 (N_8951,N_7002,N_7088);
nor U8952 (N_8952,N_7005,N_7823);
and U8953 (N_8953,N_7006,N_7630);
nand U8954 (N_8954,N_7375,N_7647);
nor U8955 (N_8955,N_7015,N_7868);
nor U8956 (N_8956,N_7556,N_7429);
or U8957 (N_8957,N_7346,N_7004);
nand U8958 (N_8958,N_7398,N_7337);
or U8959 (N_8959,N_7823,N_7873);
nor U8960 (N_8960,N_7334,N_7090);
nor U8961 (N_8961,N_7119,N_7225);
or U8962 (N_8962,N_7387,N_7445);
xor U8963 (N_8963,N_7247,N_7795);
nand U8964 (N_8964,N_7211,N_7717);
or U8965 (N_8965,N_7437,N_7894);
xor U8966 (N_8966,N_7406,N_7279);
nand U8967 (N_8967,N_7313,N_7325);
nor U8968 (N_8968,N_7551,N_7446);
and U8969 (N_8969,N_7514,N_7893);
nand U8970 (N_8970,N_7540,N_7963);
nor U8971 (N_8971,N_7941,N_7257);
nand U8972 (N_8972,N_7894,N_7617);
or U8973 (N_8973,N_7425,N_7628);
nand U8974 (N_8974,N_7755,N_7419);
xnor U8975 (N_8975,N_7429,N_7823);
xor U8976 (N_8976,N_7447,N_7712);
nor U8977 (N_8977,N_7821,N_7221);
nor U8978 (N_8978,N_7382,N_7560);
or U8979 (N_8979,N_7759,N_7951);
nand U8980 (N_8980,N_7662,N_7401);
or U8981 (N_8981,N_7192,N_7393);
and U8982 (N_8982,N_7793,N_7622);
or U8983 (N_8983,N_7197,N_7492);
or U8984 (N_8984,N_7702,N_7129);
xor U8985 (N_8985,N_7088,N_7816);
or U8986 (N_8986,N_7012,N_7226);
nor U8987 (N_8987,N_7934,N_7811);
nand U8988 (N_8988,N_7583,N_7101);
nor U8989 (N_8989,N_7796,N_7111);
nor U8990 (N_8990,N_7217,N_7415);
nand U8991 (N_8991,N_7422,N_7092);
and U8992 (N_8992,N_7085,N_7092);
nand U8993 (N_8993,N_7951,N_7625);
or U8994 (N_8994,N_7367,N_7454);
and U8995 (N_8995,N_7263,N_7596);
or U8996 (N_8996,N_7964,N_7968);
and U8997 (N_8997,N_7390,N_7610);
xnor U8998 (N_8998,N_7239,N_7433);
nor U8999 (N_8999,N_7225,N_7044);
xor U9000 (N_9000,N_8368,N_8841);
nor U9001 (N_9001,N_8164,N_8316);
or U9002 (N_9002,N_8623,N_8653);
nand U9003 (N_9003,N_8165,N_8639);
xnor U9004 (N_9004,N_8763,N_8394);
or U9005 (N_9005,N_8185,N_8967);
xor U9006 (N_9006,N_8644,N_8279);
and U9007 (N_9007,N_8170,N_8908);
xnor U9008 (N_9008,N_8740,N_8940);
and U9009 (N_9009,N_8097,N_8010);
and U9010 (N_9010,N_8152,N_8003);
or U9011 (N_9011,N_8609,N_8166);
nor U9012 (N_9012,N_8598,N_8899);
and U9013 (N_9013,N_8002,N_8363);
nand U9014 (N_9014,N_8517,N_8074);
nor U9015 (N_9015,N_8100,N_8017);
nand U9016 (N_9016,N_8088,N_8746);
nor U9017 (N_9017,N_8918,N_8086);
nand U9018 (N_9018,N_8527,N_8221);
nor U9019 (N_9019,N_8193,N_8705);
nand U9020 (N_9020,N_8791,N_8075);
xor U9021 (N_9021,N_8933,N_8982);
or U9022 (N_9022,N_8134,N_8927);
nor U9023 (N_9023,N_8347,N_8469);
nor U9024 (N_9024,N_8364,N_8774);
nor U9025 (N_9025,N_8237,N_8958);
and U9026 (N_9026,N_8851,N_8895);
nor U9027 (N_9027,N_8235,N_8995);
nor U9028 (N_9028,N_8884,N_8489);
or U9029 (N_9029,N_8990,N_8832);
nand U9030 (N_9030,N_8762,N_8563);
nand U9031 (N_9031,N_8341,N_8069);
and U9032 (N_9032,N_8696,N_8058);
or U9033 (N_9033,N_8050,N_8182);
or U9034 (N_9034,N_8189,N_8425);
and U9035 (N_9035,N_8478,N_8970);
xnor U9036 (N_9036,N_8616,N_8750);
and U9037 (N_9037,N_8805,N_8808);
xor U9038 (N_9038,N_8466,N_8124);
xor U9039 (N_9039,N_8225,N_8876);
and U9040 (N_9040,N_8168,N_8637);
and U9041 (N_9041,N_8145,N_8892);
xor U9042 (N_9042,N_8391,N_8550);
xnor U9043 (N_9043,N_8029,N_8379);
nand U9044 (N_9044,N_8471,N_8272);
nand U9045 (N_9045,N_8125,N_8813);
xor U9046 (N_9046,N_8630,N_8670);
and U9047 (N_9047,N_8321,N_8187);
and U9048 (N_9048,N_8085,N_8101);
or U9049 (N_9049,N_8936,N_8757);
or U9050 (N_9050,N_8869,N_8251);
xnor U9051 (N_9051,N_8719,N_8676);
or U9052 (N_9052,N_8924,N_8194);
nor U9053 (N_9053,N_8518,N_8432);
or U9054 (N_9054,N_8686,N_8360);
nand U9055 (N_9055,N_8349,N_8463);
and U9056 (N_9056,N_8872,N_8255);
and U9057 (N_9057,N_8092,N_8838);
xnor U9058 (N_9058,N_8036,N_8577);
and U9059 (N_9059,N_8589,N_8862);
or U9060 (N_9060,N_8878,N_8430);
nand U9061 (N_9061,N_8618,N_8094);
nor U9062 (N_9062,N_8604,N_8893);
nor U9063 (N_9063,N_8376,N_8662);
and U9064 (N_9064,N_8461,N_8373);
nand U9065 (N_9065,N_8392,N_8912);
or U9066 (N_9066,N_8920,N_8421);
xor U9067 (N_9067,N_8888,N_8938);
xnor U9068 (N_9068,N_8723,N_8283);
xor U9069 (N_9069,N_8555,N_8254);
nand U9070 (N_9070,N_8603,N_8239);
nand U9071 (N_9071,N_8181,N_8177);
and U9072 (N_9072,N_8742,N_8118);
or U9073 (N_9073,N_8854,N_8222);
xor U9074 (N_9074,N_8782,N_8687);
nor U9075 (N_9075,N_8693,N_8999);
and U9076 (N_9076,N_8579,N_8611);
xor U9077 (N_9077,N_8840,N_8848);
nand U9078 (N_9078,N_8004,N_8184);
or U9079 (N_9079,N_8792,N_8610);
nand U9080 (N_9080,N_8234,N_8881);
nor U9081 (N_9081,N_8491,N_8492);
and U9082 (N_9082,N_8262,N_8437);
xor U9083 (N_9083,N_8939,N_8581);
or U9084 (N_9084,N_8426,N_8103);
nand U9085 (N_9085,N_8093,N_8508);
nand U9086 (N_9086,N_8299,N_8830);
or U9087 (N_9087,N_8046,N_8901);
xor U9088 (N_9088,N_8654,N_8091);
nor U9089 (N_9089,N_8021,N_8119);
nor U9090 (N_9090,N_8132,N_8675);
nand U9091 (N_9091,N_8227,N_8714);
nor U9092 (N_9092,N_8057,N_8340);
or U9093 (N_9093,N_8820,N_8697);
xnor U9094 (N_9094,N_8751,N_8482);
and U9095 (N_9095,N_8907,N_8565);
or U9096 (N_9096,N_8343,N_8411);
xnor U9097 (N_9097,N_8336,N_8151);
nor U9098 (N_9098,N_8388,N_8951);
and U9099 (N_9099,N_8528,N_8290);
nand U9100 (N_9100,N_8301,N_8405);
xnor U9101 (N_9101,N_8498,N_8667);
xor U9102 (N_9102,N_8486,N_8906);
or U9103 (N_9103,N_8904,N_8961);
nor U9104 (N_9104,N_8738,N_8156);
nand U9105 (N_9105,N_8464,N_8249);
xor U9106 (N_9106,N_8393,N_8631);
or U9107 (N_9107,N_8784,N_8733);
nor U9108 (N_9108,N_8770,N_8329);
xor U9109 (N_9109,N_8661,N_8326);
and U9110 (N_9110,N_8828,N_8633);
xor U9111 (N_9111,N_8764,N_8042);
and U9112 (N_9112,N_8547,N_8732);
or U9113 (N_9113,N_8573,N_8263);
nand U9114 (N_9114,N_8073,N_8771);
xor U9115 (N_9115,N_8768,N_8082);
xor U9116 (N_9116,N_8059,N_8865);
nand U9117 (N_9117,N_8692,N_8044);
nand U9118 (N_9118,N_8399,N_8745);
and U9119 (N_9119,N_8699,N_8776);
nand U9120 (N_9120,N_8981,N_8704);
nand U9121 (N_9121,N_8846,N_8445);
nor U9122 (N_9122,N_8407,N_8635);
xor U9123 (N_9123,N_8372,N_8176);
and U9124 (N_9124,N_8921,N_8588);
and U9125 (N_9125,N_8160,N_8236);
nand U9126 (N_9126,N_8210,N_8790);
nand U9127 (N_9127,N_8355,N_8896);
xnor U9128 (N_9128,N_8837,N_8146);
xnor U9129 (N_9129,N_8529,N_8669);
and U9130 (N_9130,N_8408,N_8726);
xor U9131 (N_9131,N_8291,N_8987);
xnor U9132 (N_9132,N_8395,N_8709);
and U9133 (N_9133,N_8657,N_8700);
nand U9134 (N_9134,N_8996,N_8858);
nand U9135 (N_9135,N_8087,N_8309);
and U9136 (N_9136,N_8114,N_8035);
or U9137 (N_9137,N_8083,N_8992);
nand U9138 (N_9138,N_8931,N_8335);
nand U9139 (N_9139,N_8226,N_8576);
nor U9140 (N_9140,N_8244,N_8538);
nand U9141 (N_9141,N_8428,N_8459);
and U9142 (N_9142,N_8925,N_8786);
and U9143 (N_9143,N_8889,N_8256);
or U9144 (N_9144,N_8874,N_8328);
nor U9145 (N_9145,N_8246,N_8070);
xor U9146 (N_9146,N_8033,N_8542);
nor U9147 (N_9147,N_8135,N_8231);
nor U9148 (N_9148,N_8980,N_8849);
or U9149 (N_9149,N_8084,N_8539);
and U9150 (N_9150,N_8436,N_8624);
nand U9151 (N_9151,N_8178,N_8941);
nor U9152 (N_9152,N_8072,N_8416);
and U9153 (N_9153,N_8250,N_8449);
and U9154 (N_9154,N_8608,N_8208);
and U9155 (N_9155,N_8040,N_8883);
nand U9156 (N_9156,N_8803,N_8900);
xor U9157 (N_9157,N_8873,N_8451);
nand U9158 (N_9158,N_8795,N_8351);
or U9159 (N_9159,N_8398,N_8174);
nor U9160 (N_9160,N_8026,N_8544);
nor U9161 (N_9161,N_8983,N_8928);
xnor U9162 (N_9162,N_8270,N_8105);
nor U9163 (N_9163,N_8051,N_8028);
or U9164 (N_9164,N_8061,N_8600);
xor U9165 (N_9165,N_8822,N_8045);
nand U9166 (N_9166,N_8870,N_8626);
xor U9167 (N_9167,N_8014,N_8622);
nor U9168 (N_9168,N_8257,N_8859);
or U9169 (N_9169,N_8937,N_8882);
nand U9170 (N_9170,N_8886,N_8020);
nor U9171 (N_9171,N_8460,N_8754);
and U9172 (N_9172,N_8739,N_8488);
nand U9173 (N_9173,N_8636,N_8831);
and U9174 (N_9174,N_8023,N_8098);
nand U9175 (N_9175,N_8997,N_8671);
nand U9176 (N_9176,N_8485,N_8868);
nor U9177 (N_9177,N_8056,N_8013);
and U9178 (N_9178,N_8801,N_8140);
or U9179 (N_9179,N_8157,N_8505);
nand U9180 (N_9180,N_8298,N_8276);
and U9181 (N_9181,N_8802,N_8971);
nor U9182 (N_9182,N_8413,N_8549);
or U9183 (N_9183,N_8965,N_8747);
xor U9184 (N_9184,N_8366,N_8541);
nor U9185 (N_9185,N_8755,N_8656);
and U9186 (N_9186,N_8229,N_8816);
nor U9187 (N_9187,N_8914,N_8568);
or U9188 (N_9188,N_8897,N_8323);
nor U9189 (N_9189,N_8382,N_8294);
and U9190 (N_9190,N_8019,N_8159);
nand U9191 (N_9191,N_8613,N_8141);
or U9192 (N_9192,N_8520,N_8524);
nor U9193 (N_9193,N_8844,N_8041);
or U9194 (N_9194,N_8108,N_8353);
nor U9195 (N_9195,N_8607,N_8192);
nor U9196 (N_9196,N_8348,N_8734);
and U9197 (N_9197,N_8730,N_8111);
nor U9198 (N_9198,N_8037,N_8439);
nand U9199 (N_9199,N_8672,N_8810);
xor U9200 (N_9200,N_8409,N_8203);
nor U9201 (N_9201,N_8503,N_8556);
or U9202 (N_9202,N_8137,N_8905);
xnor U9203 (N_9203,N_8664,N_8695);
xor U9204 (N_9204,N_8259,N_8663);
xnor U9205 (N_9205,N_8233,N_8396);
and U9206 (N_9206,N_8102,N_8443);
and U9207 (N_9207,N_8964,N_8238);
and U9208 (N_9208,N_8496,N_8337);
or U9209 (N_9209,N_8817,N_8619);
nand U9210 (N_9210,N_8359,N_8674);
or U9211 (N_9211,N_8718,N_8206);
or U9212 (N_9212,N_8963,N_8902);
xnor U9213 (N_9213,N_8150,N_8659);
nand U9214 (N_9214,N_8717,N_8839);
nor U9215 (N_9215,N_8129,N_8295);
xnor U9216 (N_9216,N_8253,N_8377);
or U9217 (N_9217,N_8668,N_8324);
nor U9218 (N_9218,N_8296,N_8758);
xor U9219 (N_9219,N_8949,N_8501);
nand U9220 (N_9220,N_8632,N_8089);
and U9221 (N_9221,N_8646,N_8487);
nor U9222 (N_9222,N_8606,N_8499);
xor U9223 (N_9223,N_8153,N_8247);
xnor U9224 (N_9224,N_8712,N_8325);
nor U9225 (N_9225,N_8306,N_8318);
and U9226 (N_9226,N_8954,N_8480);
or U9227 (N_9227,N_8205,N_8665);
xnor U9228 (N_9228,N_8689,N_8476);
nand U9229 (N_9229,N_8106,N_8678);
xor U9230 (N_9230,N_8142,N_8123);
xor U9231 (N_9231,N_8063,N_8216);
nand U9232 (N_9232,N_8500,N_8648);
and U9233 (N_9233,N_8079,N_8064);
and U9234 (N_9234,N_8196,N_8371);
or U9235 (N_9235,N_8861,N_8453);
nand U9236 (N_9236,N_8344,N_8922);
or U9237 (N_9237,N_8991,N_8047);
nand U9238 (N_9238,N_8575,N_8587);
and U9239 (N_9239,N_8077,N_8209);
xnor U9240 (N_9240,N_8545,N_8759);
nor U9241 (N_9241,N_8456,N_8287);
nand U9242 (N_9242,N_8595,N_8448);
nand U9243 (N_9243,N_8877,N_8752);
nand U9244 (N_9244,N_8681,N_8357);
xor U9245 (N_9245,N_8030,N_8331);
nand U9246 (N_9246,N_8429,N_8374);
nand U9247 (N_9247,N_8702,N_8444);
and U9248 (N_9248,N_8711,N_8519);
or U9249 (N_9249,N_8024,N_8773);
nor U9250 (N_9250,N_8978,N_8826);
nor U9251 (N_9251,N_8945,N_8953);
nor U9252 (N_9252,N_8799,N_8959);
nand U9253 (N_9253,N_8943,N_8032);
nor U9254 (N_9254,N_8879,N_8475);
nand U9255 (N_9255,N_8947,N_8811);
nor U9256 (N_9256,N_8989,N_8973);
nor U9257 (N_9257,N_8628,N_8855);
or U9258 (N_9258,N_8144,N_8852);
nand U9259 (N_9259,N_8199,N_8787);
or U9260 (N_9260,N_8634,N_8120);
nand U9261 (N_9261,N_8890,N_8966);
xnor U9262 (N_9262,N_8362,N_8190);
nand U9263 (N_9263,N_8264,N_8268);
and U9264 (N_9264,N_8525,N_8706);
or U9265 (N_9265,N_8666,N_8638);
xnor U9266 (N_9266,N_8923,N_8113);
nand U9267 (N_9267,N_8490,N_8006);
nor U9268 (N_9268,N_8521,N_8725);
or U9269 (N_9269,N_8305,N_8558);
and U9270 (N_9270,N_8809,N_8812);
and U9271 (N_9271,N_8748,N_8001);
and U9272 (N_9272,N_8380,N_8412);
nand U9273 (N_9273,N_8284,N_8440);
nand U9274 (N_9274,N_8288,N_8200);
xor U9275 (N_9275,N_8384,N_8880);
and U9276 (N_9276,N_8258,N_8614);
xnor U9277 (N_9277,N_8116,N_8005);
and U9278 (N_9278,N_8772,N_8775);
xnor U9279 (N_9279,N_8853,N_8418);
nor U9280 (N_9280,N_8946,N_8683);
nor U9281 (N_9281,N_8320,N_8154);
nand U9282 (N_9282,N_8162,N_8452);
and U9283 (N_9283,N_8293,N_8167);
or U9284 (N_9284,N_8979,N_8969);
nand U9285 (N_9285,N_8076,N_8582);
nand U9286 (N_9286,N_8903,N_8169);
xor U9287 (N_9287,N_8282,N_8078);
nor U9288 (N_9288,N_8561,N_8300);
nand U9289 (N_9289,N_8535,N_8218);
xor U9290 (N_9290,N_8522,N_8333);
xnor U9291 (N_9291,N_8245,N_8534);
nor U9292 (N_9292,N_8701,N_8495);
nor U9293 (N_9293,N_8220,N_8891);
nor U9294 (N_9294,N_8578,N_8212);
nand U9295 (N_9295,N_8126,N_8523);
nor U9296 (N_9296,N_8800,N_8994);
nor U9297 (N_9297,N_8378,N_8186);
xor U9298 (N_9298,N_8000,N_8266);
or U9299 (N_9299,N_8427,N_8310);
or U9300 (N_9300,N_8562,N_8875);
nand U9301 (N_9301,N_8898,N_8984);
and U9302 (N_9302,N_8956,N_8179);
and U9303 (N_9303,N_8957,N_8807);
or U9304 (N_9304,N_8419,N_8660);
xor U9305 (N_9305,N_8474,N_8885);
nor U9306 (N_9306,N_8438,N_8531);
and U9307 (N_9307,N_8934,N_8916);
and U9308 (N_9308,N_8117,N_8548);
or U9309 (N_9309,N_8479,N_8560);
xor U9310 (N_9310,N_8369,N_8248);
nand U9311 (N_9311,N_8269,N_8338);
or U9312 (N_9312,N_8819,N_8652);
xnor U9313 (N_9313,N_8842,N_8833);
nor U9314 (N_9314,N_8365,N_8804);
and U9315 (N_9315,N_8756,N_8728);
or U9316 (N_9316,N_8798,N_8570);
or U9317 (N_9317,N_8494,N_8736);
and U9318 (N_9318,N_8617,N_8716);
nor U9319 (N_9319,N_8721,N_8434);
xor U9320 (N_9320,N_8769,N_8308);
nand U9321 (N_9321,N_8053,N_8415);
nor U9322 (N_9322,N_8387,N_8462);
or U9323 (N_9323,N_8188,N_8275);
and U9324 (N_9324,N_8009,N_8537);
xor U9325 (N_9325,N_8090,N_8055);
and U9326 (N_9326,N_8864,N_8974);
and U9327 (N_9327,N_8319,N_8354);
or U9328 (N_9328,N_8847,N_8155);
nor U9329 (N_9329,N_8691,N_8096);
nand U9330 (N_9330,N_8467,N_8385);
xnor U9331 (N_9331,N_8647,N_8694);
or U9332 (N_9332,N_8497,N_8629);
or U9333 (N_9333,N_8677,N_8332);
nor U9334 (N_9334,N_8420,N_8857);
and U9335 (N_9335,N_8417,N_8713);
and U9336 (N_9336,N_8446,N_8601);
and U9337 (N_9337,N_8223,N_8640);
xnor U9338 (N_9338,N_8099,N_8143);
and U9339 (N_9339,N_8410,N_8228);
nand U9340 (N_9340,N_8944,N_8596);
xnor U9341 (N_9341,N_8793,N_8133);
and U9342 (N_9342,N_8066,N_8543);
nand U9343 (N_9343,N_8011,N_8095);
nor U9344 (N_9344,N_8127,N_8345);
or U9345 (N_9345,N_8131,N_8825);
and U9346 (N_9346,N_8242,N_8753);
or U9347 (N_9347,N_8559,N_8115);
xor U9348 (N_9348,N_8972,N_8403);
nand U9349 (N_9349,N_8850,N_8285);
nand U9350 (N_9350,N_8472,N_8370);
and U9351 (N_9351,N_8530,N_8224);
nor U9352 (N_9352,N_8313,N_8243);
xnor U9353 (N_9353,N_8330,N_8926);
nor U9354 (N_9354,N_8381,N_8815);
or U9355 (N_9355,N_8557,N_8546);
nand U9356 (N_9356,N_8361,N_8511);
nor U9357 (N_9357,N_8690,N_8468);
nand U9358 (N_9358,N_8553,N_8625);
nor U9359 (N_9359,N_8346,N_8867);
nand U9360 (N_9360,N_8685,N_8230);
nand U9361 (N_9361,N_8955,N_8433);
or U9362 (N_9362,N_8599,N_8201);
xnor U9363 (N_9363,N_8180,N_8533);
xor U9364 (N_9364,N_8265,N_8367);
nor U9365 (N_9365,N_8767,N_8504);
and U9366 (N_9366,N_8516,N_8375);
nand U9367 (N_9367,N_8281,N_8191);
nor U9368 (N_9368,N_8483,N_8993);
or U9369 (N_9369,N_8173,N_8147);
xor U9370 (N_9370,N_8986,N_8441);
nand U9371 (N_9371,N_8240,N_8917);
nand U9372 (N_9372,N_8703,N_8871);
nor U9373 (N_9373,N_8386,N_8569);
nor U9374 (N_9374,N_8827,N_8473);
or U9375 (N_9375,N_8402,N_8679);
or U9376 (N_9376,N_8317,N_8829);
nand U9377 (N_9377,N_8797,N_8651);
xnor U9378 (N_9378,N_8593,N_8022);
and U9379 (N_9379,N_8856,N_8836);
or U9380 (N_9380,N_8860,N_8252);
or U9381 (N_9381,N_8110,N_8552);
xnor U9382 (N_9382,N_8975,N_8292);
nor U9383 (N_9383,N_8390,N_8139);
nor U9384 (N_9384,N_8735,N_8389);
nor U9385 (N_9385,N_8406,N_8835);
xor U9386 (N_9386,N_8356,N_8602);
and U9387 (N_9387,N_8650,N_8477);
nand U9388 (N_9388,N_8450,N_8779);
or U9389 (N_9389,N_8314,N_8722);
nand U9390 (N_9390,N_8457,N_8404);
xnor U9391 (N_9391,N_8303,N_8334);
nand U9392 (N_9392,N_8315,N_8038);
xor U9393 (N_9393,N_8778,N_8311);
and U9394 (N_9394,N_8514,N_8031);
nand U9395 (N_9395,N_8824,N_8271);
nand U9396 (N_9396,N_8605,N_8027);
or U9397 (N_9397,N_8590,N_8149);
or U9398 (N_9398,N_8350,N_8952);
and U9399 (N_9399,N_8863,N_8688);
xnor U9400 (N_9400,N_8585,N_8976);
xor U9401 (N_9401,N_8788,N_8148);
xnor U9402 (N_9402,N_8327,N_8278);
nand U9403 (N_9403,N_8777,N_8554);
and U9404 (N_9404,N_8136,N_8307);
xor U9405 (N_9405,N_8929,N_8458);
nand U9406 (N_9406,N_8067,N_8358);
or U9407 (N_9407,N_8304,N_8109);
or U9408 (N_9408,N_8536,N_8195);
nor U9409 (N_9409,N_8684,N_8071);
nor U9410 (N_9410,N_8007,N_8513);
nor U9411 (N_9411,N_8707,N_8540);
and U9412 (N_9412,N_8615,N_8470);
or U9413 (N_9413,N_8724,N_8729);
nor U9414 (N_9414,N_8509,N_8081);
nand U9415 (N_9415,N_8597,N_8049);
nor U9416 (N_9416,N_8698,N_8054);
nor U9417 (N_9417,N_8016,N_8274);
nor U9418 (N_9418,N_8502,N_8814);
xor U9419 (N_9419,N_8998,N_8507);
or U9420 (N_9420,N_8621,N_8232);
xor U9421 (N_9421,N_8708,N_8138);
nand U9422 (N_9422,N_8197,N_8765);
nand U9423 (N_9423,N_8977,N_8204);
or U9424 (N_9424,N_8080,N_8025);
or U9425 (N_9425,N_8175,N_8202);
xor U9426 (N_9426,N_8400,N_8062);
and U9427 (N_9427,N_8806,N_8104);
and U9428 (N_9428,N_8780,N_8731);
xor U9429 (N_9429,N_8183,N_8060);
nand U9430 (N_9430,N_8465,N_8942);
nor U9431 (N_9431,N_8919,N_8985);
xor U9432 (N_9432,N_8442,N_8214);
xnor U9433 (N_9433,N_8018,N_8423);
or U9434 (N_9434,N_8642,N_8641);
or U9435 (N_9435,N_8012,N_8068);
nand U9436 (N_9436,N_8526,N_8794);
nor U9437 (N_9437,N_8843,N_8107);
and U9438 (N_9438,N_8130,N_8715);
nor U9439 (N_9439,N_8112,N_8781);
nor U9440 (N_9440,N_8342,N_8566);
nand U9441 (N_9441,N_8273,N_8655);
nand U9442 (N_9442,N_8572,N_8785);
nand U9443 (N_9443,N_8962,N_8894);
xor U9444 (N_9444,N_8217,N_8789);
nand U9445 (N_9445,N_8761,N_8760);
or U9446 (N_9446,N_8834,N_8506);
xor U9447 (N_9447,N_8352,N_8414);
nor U9448 (N_9448,N_8213,N_8909);
nor U9449 (N_9449,N_8551,N_8571);
xnor U9450 (N_9450,N_8818,N_8484);
nor U9451 (N_9451,N_8988,N_8737);
nor U9452 (N_9452,N_8741,N_8720);
and U9453 (N_9453,N_8454,N_8915);
and U9454 (N_9454,N_8383,N_8821);
nor U9455 (N_9455,N_8493,N_8643);
nand U9456 (N_9456,N_8911,N_8215);
xor U9457 (N_9457,N_8866,N_8574);
nor U9458 (N_9458,N_8455,N_8960);
xor U9459 (N_9459,N_8749,N_8649);
nor U9460 (N_9460,N_8645,N_8567);
nor U9461 (N_9461,N_8682,N_8161);
nor U9462 (N_9462,N_8008,N_8039);
or U9463 (N_9463,N_8783,N_8289);
nand U9464 (N_9464,N_8302,N_8339);
xnor U9465 (N_9465,N_8401,N_8532);
nor U9466 (N_9466,N_8211,N_8122);
or U9467 (N_9467,N_8932,N_8207);
nor U9468 (N_9468,N_8297,N_8673);
xnor U9469 (N_9469,N_8743,N_8620);
nor U9470 (N_9470,N_8172,N_8680);
xnor U9471 (N_9471,N_8887,N_8043);
or U9472 (N_9472,N_8910,N_8286);
xor U9473 (N_9473,N_8397,N_8261);
xor U9474 (N_9474,N_8564,N_8515);
nor U9475 (N_9475,N_8796,N_8612);
and U9476 (N_9476,N_8158,N_8580);
and U9477 (N_9477,N_8198,N_8424);
xnor U9478 (N_9478,N_8948,N_8065);
and U9479 (N_9479,N_8930,N_8447);
nor U9480 (N_9480,N_8322,N_8913);
nor U9481 (N_9481,N_8766,N_8312);
nand U9482 (N_9482,N_8727,N_8052);
nor U9483 (N_9483,N_8422,N_8744);
nand U9484 (N_9484,N_8845,N_8586);
or U9485 (N_9485,N_8591,N_8241);
nor U9486 (N_9486,N_8510,N_8950);
nand U9487 (N_9487,N_8627,N_8594);
or U9488 (N_9488,N_8823,N_8034);
nand U9489 (N_9489,N_8583,N_8968);
or U9490 (N_9490,N_8481,N_8260);
nand U9491 (N_9491,N_8015,N_8935);
or U9492 (N_9492,N_8584,N_8128);
and U9493 (N_9493,N_8658,N_8267);
or U9494 (N_9494,N_8592,N_8219);
nand U9495 (N_9495,N_8048,N_8277);
nor U9496 (N_9496,N_8121,N_8280);
and U9497 (N_9497,N_8171,N_8163);
and U9498 (N_9498,N_8710,N_8512);
and U9499 (N_9499,N_8431,N_8435);
nor U9500 (N_9500,N_8155,N_8353);
xor U9501 (N_9501,N_8923,N_8674);
nor U9502 (N_9502,N_8249,N_8509);
and U9503 (N_9503,N_8949,N_8329);
and U9504 (N_9504,N_8871,N_8738);
nand U9505 (N_9505,N_8714,N_8506);
nand U9506 (N_9506,N_8743,N_8703);
xor U9507 (N_9507,N_8300,N_8610);
nor U9508 (N_9508,N_8159,N_8975);
nor U9509 (N_9509,N_8933,N_8431);
xnor U9510 (N_9510,N_8658,N_8458);
nor U9511 (N_9511,N_8293,N_8162);
nor U9512 (N_9512,N_8695,N_8349);
xnor U9513 (N_9513,N_8350,N_8541);
nor U9514 (N_9514,N_8281,N_8145);
or U9515 (N_9515,N_8688,N_8468);
and U9516 (N_9516,N_8403,N_8045);
and U9517 (N_9517,N_8438,N_8181);
xnor U9518 (N_9518,N_8488,N_8524);
or U9519 (N_9519,N_8033,N_8607);
nand U9520 (N_9520,N_8959,N_8161);
nor U9521 (N_9521,N_8106,N_8804);
nor U9522 (N_9522,N_8401,N_8533);
nand U9523 (N_9523,N_8123,N_8061);
and U9524 (N_9524,N_8204,N_8863);
xnor U9525 (N_9525,N_8422,N_8167);
xnor U9526 (N_9526,N_8638,N_8152);
xnor U9527 (N_9527,N_8224,N_8172);
nor U9528 (N_9528,N_8411,N_8905);
nor U9529 (N_9529,N_8828,N_8566);
or U9530 (N_9530,N_8523,N_8847);
and U9531 (N_9531,N_8810,N_8946);
and U9532 (N_9532,N_8096,N_8680);
xor U9533 (N_9533,N_8976,N_8266);
xnor U9534 (N_9534,N_8806,N_8801);
nand U9535 (N_9535,N_8691,N_8240);
xor U9536 (N_9536,N_8582,N_8460);
nor U9537 (N_9537,N_8257,N_8486);
xor U9538 (N_9538,N_8965,N_8653);
or U9539 (N_9539,N_8111,N_8023);
or U9540 (N_9540,N_8292,N_8313);
xnor U9541 (N_9541,N_8490,N_8421);
xnor U9542 (N_9542,N_8053,N_8553);
xor U9543 (N_9543,N_8888,N_8314);
and U9544 (N_9544,N_8218,N_8987);
nor U9545 (N_9545,N_8338,N_8212);
or U9546 (N_9546,N_8775,N_8516);
nand U9547 (N_9547,N_8575,N_8978);
xnor U9548 (N_9548,N_8099,N_8623);
nand U9549 (N_9549,N_8649,N_8091);
nand U9550 (N_9550,N_8563,N_8554);
or U9551 (N_9551,N_8660,N_8527);
nand U9552 (N_9552,N_8137,N_8237);
and U9553 (N_9553,N_8620,N_8590);
nand U9554 (N_9554,N_8904,N_8172);
nor U9555 (N_9555,N_8541,N_8030);
and U9556 (N_9556,N_8538,N_8557);
xor U9557 (N_9557,N_8714,N_8911);
nor U9558 (N_9558,N_8294,N_8746);
nand U9559 (N_9559,N_8026,N_8819);
or U9560 (N_9560,N_8399,N_8153);
nor U9561 (N_9561,N_8287,N_8639);
nand U9562 (N_9562,N_8533,N_8774);
xor U9563 (N_9563,N_8038,N_8873);
or U9564 (N_9564,N_8658,N_8518);
nand U9565 (N_9565,N_8690,N_8864);
nor U9566 (N_9566,N_8137,N_8437);
nor U9567 (N_9567,N_8420,N_8575);
xor U9568 (N_9568,N_8562,N_8934);
nor U9569 (N_9569,N_8084,N_8782);
or U9570 (N_9570,N_8497,N_8616);
nand U9571 (N_9571,N_8743,N_8903);
nor U9572 (N_9572,N_8924,N_8747);
nor U9573 (N_9573,N_8119,N_8925);
nand U9574 (N_9574,N_8721,N_8291);
nor U9575 (N_9575,N_8894,N_8474);
nor U9576 (N_9576,N_8867,N_8143);
nand U9577 (N_9577,N_8678,N_8737);
nor U9578 (N_9578,N_8286,N_8926);
and U9579 (N_9579,N_8999,N_8618);
xor U9580 (N_9580,N_8127,N_8830);
or U9581 (N_9581,N_8143,N_8874);
nor U9582 (N_9582,N_8730,N_8009);
or U9583 (N_9583,N_8807,N_8566);
and U9584 (N_9584,N_8939,N_8591);
nor U9585 (N_9585,N_8127,N_8460);
nor U9586 (N_9586,N_8021,N_8391);
and U9587 (N_9587,N_8165,N_8313);
nor U9588 (N_9588,N_8354,N_8458);
and U9589 (N_9589,N_8033,N_8177);
or U9590 (N_9590,N_8950,N_8210);
and U9591 (N_9591,N_8298,N_8283);
nand U9592 (N_9592,N_8333,N_8387);
and U9593 (N_9593,N_8164,N_8243);
xnor U9594 (N_9594,N_8282,N_8112);
nor U9595 (N_9595,N_8481,N_8723);
nand U9596 (N_9596,N_8868,N_8186);
nor U9597 (N_9597,N_8322,N_8042);
nor U9598 (N_9598,N_8791,N_8472);
or U9599 (N_9599,N_8351,N_8607);
nand U9600 (N_9600,N_8073,N_8209);
nor U9601 (N_9601,N_8354,N_8717);
and U9602 (N_9602,N_8052,N_8949);
nand U9603 (N_9603,N_8950,N_8585);
or U9604 (N_9604,N_8605,N_8373);
nor U9605 (N_9605,N_8590,N_8174);
and U9606 (N_9606,N_8720,N_8340);
and U9607 (N_9607,N_8275,N_8433);
nand U9608 (N_9608,N_8228,N_8646);
nand U9609 (N_9609,N_8238,N_8898);
or U9610 (N_9610,N_8669,N_8931);
or U9611 (N_9611,N_8867,N_8454);
xnor U9612 (N_9612,N_8007,N_8506);
nand U9613 (N_9613,N_8106,N_8949);
and U9614 (N_9614,N_8904,N_8754);
or U9615 (N_9615,N_8864,N_8111);
nor U9616 (N_9616,N_8908,N_8997);
nor U9617 (N_9617,N_8107,N_8050);
nor U9618 (N_9618,N_8006,N_8903);
nor U9619 (N_9619,N_8631,N_8637);
and U9620 (N_9620,N_8910,N_8608);
nor U9621 (N_9621,N_8424,N_8757);
nand U9622 (N_9622,N_8023,N_8774);
xnor U9623 (N_9623,N_8117,N_8409);
and U9624 (N_9624,N_8721,N_8894);
nand U9625 (N_9625,N_8867,N_8880);
or U9626 (N_9626,N_8802,N_8219);
nand U9627 (N_9627,N_8230,N_8515);
nor U9628 (N_9628,N_8130,N_8477);
and U9629 (N_9629,N_8547,N_8164);
nor U9630 (N_9630,N_8503,N_8881);
nor U9631 (N_9631,N_8978,N_8062);
xnor U9632 (N_9632,N_8519,N_8839);
and U9633 (N_9633,N_8629,N_8386);
or U9634 (N_9634,N_8622,N_8380);
nand U9635 (N_9635,N_8003,N_8434);
or U9636 (N_9636,N_8158,N_8389);
or U9637 (N_9637,N_8643,N_8006);
xor U9638 (N_9638,N_8203,N_8485);
and U9639 (N_9639,N_8797,N_8371);
and U9640 (N_9640,N_8002,N_8245);
nor U9641 (N_9641,N_8196,N_8225);
xor U9642 (N_9642,N_8378,N_8355);
nand U9643 (N_9643,N_8033,N_8949);
and U9644 (N_9644,N_8672,N_8902);
or U9645 (N_9645,N_8550,N_8760);
nor U9646 (N_9646,N_8095,N_8625);
xnor U9647 (N_9647,N_8267,N_8310);
and U9648 (N_9648,N_8878,N_8992);
and U9649 (N_9649,N_8003,N_8668);
nor U9650 (N_9650,N_8394,N_8284);
nor U9651 (N_9651,N_8745,N_8956);
or U9652 (N_9652,N_8108,N_8288);
or U9653 (N_9653,N_8830,N_8130);
nand U9654 (N_9654,N_8362,N_8485);
xor U9655 (N_9655,N_8488,N_8725);
or U9656 (N_9656,N_8203,N_8293);
xor U9657 (N_9657,N_8545,N_8279);
nor U9658 (N_9658,N_8396,N_8460);
or U9659 (N_9659,N_8053,N_8625);
or U9660 (N_9660,N_8060,N_8640);
and U9661 (N_9661,N_8647,N_8411);
and U9662 (N_9662,N_8643,N_8005);
xor U9663 (N_9663,N_8118,N_8165);
and U9664 (N_9664,N_8308,N_8609);
xnor U9665 (N_9665,N_8013,N_8490);
nand U9666 (N_9666,N_8890,N_8223);
nor U9667 (N_9667,N_8009,N_8487);
or U9668 (N_9668,N_8122,N_8947);
xor U9669 (N_9669,N_8529,N_8452);
or U9670 (N_9670,N_8973,N_8927);
nor U9671 (N_9671,N_8243,N_8130);
and U9672 (N_9672,N_8930,N_8333);
nor U9673 (N_9673,N_8588,N_8105);
xor U9674 (N_9674,N_8664,N_8851);
and U9675 (N_9675,N_8491,N_8945);
and U9676 (N_9676,N_8990,N_8117);
xor U9677 (N_9677,N_8667,N_8467);
or U9678 (N_9678,N_8277,N_8999);
and U9679 (N_9679,N_8007,N_8146);
nor U9680 (N_9680,N_8666,N_8025);
or U9681 (N_9681,N_8386,N_8766);
or U9682 (N_9682,N_8735,N_8005);
xnor U9683 (N_9683,N_8484,N_8201);
xnor U9684 (N_9684,N_8036,N_8441);
xor U9685 (N_9685,N_8258,N_8823);
or U9686 (N_9686,N_8010,N_8935);
and U9687 (N_9687,N_8152,N_8220);
xor U9688 (N_9688,N_8702,N_8092);
nor U9689 (N_9689,N_8412,N_8363);
or U9690 (N_9690,N_8541,N_8469);
nand U9691 (N_9691,N_8062,N_8254);
and U9692 (N_9692,N_8904,N_8740);
or U9693 (N_9693,N_8609,N_8218);
xor U9694 (N_9694,N_8470,N_8355);
nor U9695 (N_9695,N_8802,N_8349);
nor U9696 (N_9696,N_8957,N_8855);
and U9697 (N_9697,N_8010,N_8420);
nor U9698 (N_9698,N_8417,N_8608);
or U9699 (N_9699,N_8851,N_8436);
xor U9700 (N_9700,N_8892,N_8425);
and U9701 (N_9701,N_8327,N_8726);
nor U9702 (N_9702,N_8732,N_8284);
xor U9703 (N_9703,N_8463,N_8241);
nand U9704 (N_9704,N_8611,N_8170);
or U9705 (N_9705,N_8920,N_8558);
nand U9706 (N_9706,N_8154,N_8629);
and U9707 (N_9707,N_8070,N_8447);
nand U9708 (N_9708,N_8865,N_8107);
and U9709 (N_9709,N_8603,N_8931);
nor U9710 (N_9710,N_8567,N_8950);
and U9711 (N_9711,N_8742,N_8825);
or U9712 (N_9712,N_8374,N_8337);
nor U9713 (N_9713,N_8557,N_8483);
nand U9714 (N_9714,N_8302,N_8018);
xnor U9715 (N_9715,N_8841,N_8165);
nor U9716 (N_9716,N_8916,N_8711);
nand U9717 (N_9717,N_8217,N_8422);
xnor U9718 (N_9718,N_8511,N_8948);
nand U9719 (N_9719,N_8817,N_8612);
and U9720 (N_9720,N_8775,N_8356);
xor U9721 (N_9721,N_8589,N_8876);
nor U9722 (N_9722,N_8109,N_8497);
xor U9723 (N_9723,N_8584,N_8179);
nand U9724 (N_9724,N_8209,N_8897);
xnor U9725 (N_9725,N_8535,N_8974);
nor U9726 (N_9726,N_8634,N_8111);
nor U9727 (N_9727,N_8926,N_8387);
nor U9728 (N_9728,N_8991,N_8868);
and U9729 (N_9729,N_8908,N_8470);
xnor U9730 (N_9730,N_8601,N_8952);
xnor U9731 (N_9731,N_8092,N_8968);
xor U9732 (N_9732,N_8710,N_8742);
and U9733 (N_9733,N_8198,N_8277);
and U9734 (N_9734,N_8450,N_8968);
and U9735 (N_9735,N_8254,N_8830);
xor U9736 (N_9736,N_8168,N_8792);
and U9737 (N_9737,N_8982,N_8620);
nor U9738 (N_9738,N_8051,N_8508);
nor U9739 (N_9739,N_8942,N_8812);
or U9740 (N_9740,N_8069,N_8929);
and U9741 (N_9741,N_8130,N_8979);
nand U9742 (N_9742,N_8401,N_8404);
nor U9743 (N_9743,N_8547,N_8679);
xnor U9744 (N_9744,N_8664,N_8382);
nand U9745 (N_9745,N_8525,N_8654);
nand U9746 (N_9746,N_8760,N_8357);
or U9747 (N_9747,N_8039,N_8776);
and U9748 (N_9748,N_8583,N_8555);
nor U9749 (N_9749,N_8157,N_8799);
nand U9750 (N_9750,N_8772,N_8871);
or U9751 (N_9751,N_8864,N_8171);
or U9752 (N_9752,N_8345,N_8257);
nand U9753 (N_9753,N_8643,N_8064);
nor U9754 (N_9754,N_8500,N_8436);
and U9755 (N_9755,N_8975,N_8006);
and U9756 (N_9756,N_8258,N_8316);
and U9757 (N_9757,N_8226,N_8266);
nand U9758 (N_9758,N_8871,N_8222);
and U9759 (N_9759,N_8590,N_8037);
xor U9760 (N_9760,N_8350,N_8967);
nand U9761 (N_9761,N_8787,N_8198);
and U9762 (N_9762,N_8687,N_8385);
or U9763 (N_9763,N_8325,N_8273);
xor U9764 (N_9764,N_8906,N_8677);
or U9765 (N_9765,N_8900,N_8440);
and U9766 (N_9766,N_8932,N_8559);
nor U9767 (N_9767,N_8088,N_8296);
or U9768 (N_9768,N_8515,N_8504);
nor U9769 (N_9769,N_8605,N_8970);
xor U9770 (N_9770,N_8785,N_8409);
or U9771 (N_9771,N_8782,N_8938);
nand U9772 (N_9772,N_8823,N_8162);
or U9773 (N_9773,N_8020,N_8537);
and U9774 (N_9774,N_8867,N_8423);
and U9775 (N_9775,N_8860,N_8248);
and U9776 (N_9776,N_8205,N_8170);
xor U9777 (N_9777,N_8212,N_8692);
xor U9778 (N_9778,N_8968,N_8125);
and U9779 (N_9779,N_8995,N_8091);
nand U9780 (N_9780,N_8854,N_8331);
and U9781 (N_9781,N_8101,N_8380);
nand U9782 (N_9782,N_8261,N_8111);
nand U9783 (N_9783,N_8518,N_8495);
or U9784 (N_9784,N_8234,N_8026);
xnor U9785 (N_9785,N_8856,N_8116);
and U9786 (N_9786,N_8269,N_8478);
xnor U9787 (N_9787,N_8992,N_8974);
xnor U9788 (N_9788,N_8953,N_8857);
or U9789 (N_9789,N_8069,N_8416);
nand U9790 (N_9790,N_8953,N_8966);
nor U9791 (N_9791,N_8692,N_8056);
nand U9792 (N_9792,N_8824,N_8541);
nor U9793 (N_9793,N_8880,N_8570);
or U9794 (N_9794,N_8959,N_8089);
xor U9795 (N_9795,N_8997,N_8079);
and U9796 (N_9796,N_8206,N_8391);
or U9797 (N_9797,N_8651,N_8072);
xnor U9798 (N_9798,N_8445,N_8195);
and U9799 (N_9799,N_8359,N_8533);
nand U9800 (N_9800,N_8654,N_8038);
nor U9801 (N_9801,N_8077,N_8555);
nor U9802 (N_9802,N_8484,N_8263);
or U9803 (N_9803,N_8306,N_8448);
nor U9804 (N_9804,N_8074,N_8399);
or U9805 (N_9805,N_8425,N_8629);
and U9806 (N_9806,N_8585,N_8113);
nor U9807 (N_9807,N_8045,N_8722);
or U9808 (N_9808,N_8200,N_8775);
nand U9809 (N_9809,N_8443,N_8911);
or U9810 (N_9810,N_8363,N_8257);
xor U9811 (N_9811,N_8941,N_8106);
xnor U9812 (N_9812,N_8827,N_8731);
nor U9813 (N_9813,N_8418,N_8164);
nor U9814 (N_9814,N_8787,N_8004);
xnor U9815 (N_9815,N_8497,N_8041);
xnor U9816 (N_9816,N_8714,N_8209);
and U9817 (N_9817,N_8706,N_8229);
and U9818 (N_9818,N_8331,N_8911);
or U9819 (N_9819,N_8357,N_8998);
xnor U9820 (N_9820,N_8227,N_8390);
or U9821 (N_9821,N_8498,N_8064);
xnor U9822 (N_9822,N_8695,N_8908);
nor U9823 (N_9823,N_8571,N_8356);
or U9824 (N_9824,N_8718,N_8515);
or U9825 (N_9825,N_8822,N_8586);
or U9826 (N_9826,N_8349,N_8318);
nand U9827 (N_9827,N_8168,N_8897);
xor U9828 (N_9828,N_8894,N_8905);
or U9829 (N_9829,N_8425,N_8825);
nand U9830 (N_9830,N_8716,N_8911);
or U9831 (N_9831,N_8292,N_8173);
nand U9832 (N_9832,N_8168,N_8458);
nor U9833 (N_9833,N_8750,N_8191);
or U9834 (N_9834,N_8550,N_8476);
nand U9835 (N_9835,N_8140,N_8788);
nand U9836 (N_9836,N_8602,N_8913);
nand U9837 (N_9837,N_8689,N_8841);
xnor U9838 (N_9838,N_8949,N_8553);
xor U9839 (N_9839,N_8083,N_8336);
xnor U9840 (N_9840,N_8178,N_8450);
and U9841 (N_9841,N_8079,N_8798);
nand U9842 (N_9842,N_8110,N_8741);
and U9843 (N_9843,N_8597,N_8894);
or U9844 (N_9844,N_8696,N_8680);
or U9845 (N_9845,N_8490,N_8880);
and U9846 (N_9846,N_8004,N_8468);
or U9847 (N_9847,N_8058,N_8903);
or U9848 (N_9848,N_8521,N_8284);
and U9849 (N_9849,N_8183,N_8764);
xor U9850 (N_9850,N_8783,N_8566);
nand U9851 (N_9851,N_8724,N_8461);
nor U9852 (N_9852,N_8541,N_8840);
or U9853 (N_9853,N_8898,N_8671);
nor U9854 (N_9854,N_8024,N_8735);
and U9855 (N_9855,N_8436,N_8165);
nand U9856 (N_9856,N_8479,N_8546);
nor U9857 (N_9857,N_8569,N_8670);
xnor U9858 (N_9858,N_8503,N_8957);
xor U9859 (N_9859,N_8151,N_8968);
or U9860 (N_9860,N_8246,N_8307);
nor U9861 (N_9861,N_8928,N_8289);
nor U9862 (N_9862,N_8261,N_8843);
xnor U9863 (N_9863,N_8088,N_8789);
nand U9864 (N_9864,N_8307,N_8757);
or U9865 (N_9865,N_8618,N_8491);
xnor U9866 (N_9866,N_8422,N_8166);
xnor U9867 (N_9867,N_8597,N_8077);
or U9868 (N_9868,N_8135,N_8884);
nor U9869 (N_9869,N_8835,N_8980);
nand U9870 (N_9870,N_8506,N_8604);
nor U9871 (N_9871,N_8751,N_8214);
xor U9872 (N_9872,N_8483,N_8730);
or U9873 (N_9873,N_8873,N_8010);
nor U9874 (N_9874,N_8252,N_8476);
xor U9875 (N_9875,N_8822,N_8015);
and U9876 (N_9876,N_8330,N_8034);
xnor U9877 (N_9877,N_8043,N_8175);
xnor U9878 (N_9878,N_8048,N_8340);
xnor U9879 (N_9879,N_8340,N_8342);
nor U9880 (N_9880,N_8037,N_8748);
nor U9881 (N_9881,N_8313,N_8020);
nor U9882 (N_9882,N_8175,N_8281);
xnor U9883 (N_9883,N_8040,N_8822);
or U9884 (N_9884,N_8220,N_8959);
or U9885 (N_9885,N_8908,N_8492);
xor U9886 (N_9886,N_8373,N_8862);
or U9887 (N_9887,N_8295,N_8851);
nand U9888 (N_9888,N_8239,N_8830);
and U9889 (N_9889,N_8290,N_8877);
or U9890 (N_9890,N_8324,N_8512);
and U9891 (N_9891,N_8263,N_8487);
and U9892 (N_9892,N_8863,N_8014);
xor U9893 (N_9893,N_8398,N_8004);
xor U9894 (N_9894,N_8846,N_8210);
nand U9895 (N_9895,N_8541,N_8887);
nand U9896 (N_9896,N_8145,N_8434);
or U9897 (N_9897,N_8102,N_8552);
nor U9898 (N_9898,N_8716,N_8816);
nor U9899 (N_9899,N_8229,N_8098);
and U9900 (N_9900,N_8293,N_8096);
and U9901 (N_9901,N_8523,N_8608);
nand U9902 (N_9902,N_8835,N_8636);
nor U9903 (N_9903,N_8521,N_8530);
xor U9904 (N_9904,N_8157,N_8805);
nand U9905 (N_9905,N_8926,N_8907);
and U9906 (N_9906,N_8970,N_8723);
and U9907 (N_9907,N_8250,N_8965);
or U9908 (N_9908,N_8797,N_8707);
xnor U9909 (N_9909,N_8669,N_8569);
or U9910 (N_9910,N_8644,N_8123);
and U9911 (N_9911,N_8951,N_8622);
and U9912 (N_9912,N_8653,N_8107);
nand U9913 (N_9913,N_8121,N_8155);
nand U9914 (N_9914,N_8281,N_8576);
xor U9915 (N_9915,N_8407,N_8979);
nand U9916 (N_9916,N_8968,N_8720);
nand U9917 (N_9917,N_8498,N_8189);
or U9918 (N_9918,N_8347,N_8404);
nor U9919 (N_9919,N_8536,N_8869);
nand U9920 (N_9920,N_8976,N_8252);
nand U9921 (N_9921,N_8851,N_8178);
nor U9922 (N_9922,N_8801,N_8729);
nand U9923 (N_9923,N_8489,N_8292);
and U9924 (N_9924,N_8523,N_8535);
nor U9925 (N_9925,N_8389,N_8475);
nor U9926 (N_9926,N_8566,N_8114);
or U9927 (N_9927,N_8142,N_8477);
nor U9928 (N_9928,N_8660,N_8475);
nor U9929 (N_9929,N_8082,N_8702);
and U9930 (N_9930,N_8305,N_8910);
nand U9931 (N_9931,N_8303,N_8567);
and U9932 (N_9932,N_8867,N_8377);
or U9933 (N_9933,N_8161,N_8481);
nand U9934 (N_9934,N_8156,N_8802);
nand U9935 (N_9935,N_8490,N_8825);
nor U9936 (N_9936,N_8986,N_8242);
or U9937 (N_9937,N_8797,N_8031);
nor U9938 (N_9938,N_8503,N_8912);
nor U9939 (N_9939,N_8665,N_8196);
nand U9940 (N_9940,N_8508,N_8961);
or U9941 (N_9941,N_8286,N_8050);
xnor U9942 (N_9942,N_8189,N_8374);
and U9943 (N_9943,N_8949,N_8076);
and U9944 (N_9944,N_8144,N_8042);
nor U9945 (N_9945,N_8787,N_8594);
or U9946 (N_9946,N_8614,N_8321);
xnor U9947 (N_9947,N_8677,N_8782);
and U9948 (N_9948,N_8745,N_8813);
or U9949 (N_9949,N_8335,N_8786);
nand U9950 (N_9950,N_8835,N_8728);
xor U9951 (N_9951,N_8610,N_8542);
nor U9952 (N_9952,N_8906,N_8648);
xor U9953 (N_9953,N_8684,N_8642);
or U9954 (N_9954,N_8401,N_8021);
nor U9955 (N_9955,N_8760,N_8474);
or U9956 (N_9956,N_8281,N_8949);
nor U9957 (N_9957,N_8432,N_8467);
nand U9958 (N_9958,N_8166,N_8552);
nor U9959 (N_9959,N_8987,N_8299);
or U9960 (N_9960,N_8107,N_8136);
or U9961 (N_9961,N_8432,N_8475);
or U9962 (N_9962,N_8428,N_8606);
nor U9963 (N_9963,N_8572,N_8079);
and U9964 (N_9964,N_8479,N_8987);
nand U9965 (N_9965,N_8520,N_8194);
or U9966 (N_9966,N_8836,N_8994);
xor U9967 (N_9967,N_8224,N_8783);
and U9968 (N_9968,N_8219,N_8035);
nor U9969 (N_9969,N_8498,N_8629);
and U9970 (N_9970,N_8968,N_8838);
and U9971 (N_9971,N_8030,N_8606);
or U9972 (N_9972,N_8913,N_8748);
xnor U9973 (N_9973,N_8196,N_8083);
or U9974 (N_9974,N_8031,N_8078);
xor U9975 (N_9975,N_8861,N_8025);
or U9976 (N_9976,N_8650,N_8962);
or U9977 (N_9977,N_8479,N_8856);
and U9978 (N_9978,N_8264,N_8452);
or U9979 (N_9979,N_8417,N_8836);
xor U9980 (N_9980,N_8929,N_8088);
nor U9981 (N_9981,N_8745,N_8682);
and U9982 (N_9982,N_8908,N_8689);
and U9983 (N_9983,N_8776,N_8649);
or U9984 (N_9984,N_8573,N_8204);
nand U9985 (N_9985,N_8862,N_8982);
nor U9986 (N_9986,N_8704,N_8197);
and U9987 (N_9987,N_8621,N_8995);
nor U9988 (N_9988,N_8363,N_8986);
or U9989 (N_9989,N_8087,N_8515);
xor U9990 (N_9990,N_8145,N_8634);
xnor U9991 (N_9991,N_8111,N_8393);
nand U9992 (N_9992,N_8627,N_8415);
nand U9993 (N_9993,N_8589,N_8453);
nand U9994 (N_9994,N_8851,N_8542);
xor U9995 (N_9995,N_8918,N_8392);
or U9996 (N_9996,N_8115,N_8705);
nor U9997 (N_9997,N_8546,N_8564);
and U9998 (N_9998,N_8644,N_8259);
or U9999 (N_9999,N_8616,N_8140);
xor UO_0 (O_0,N_9390,N_9688);
and UO_1 (O_1,N_9391,N_9776);
nand UO_2 (O_2,N_9584,N_9811);
nor UO_3 (O_3,N_9227,N_9257);
nand UO_4 (O_4,N_9942,N_9752);
or UO_5 (O_5,N_9235,N_9480);
and UO_6 (O_6,N_9302,N_9279);
and UO_7 (O_7,N_9578,N_9101);
xnor UO_8 (O_8,N_9907,N_9184);
xnor UO_9 (O_9,N_9309,N_9087);
nor UO_10 (O_10,N_9926,N_9543);
and UO_11 (O_11,N_9135,N_9167);
nor UO_12 (O_12,N_9594,N_9016);
nand UO_13 (O_13,N_9654,N_9422);
and UO_14 (O_14,N_9367,N_9321);
and UO_15 (O_15,N_9627,N_9557);
nor UO_16 (O_16,N_9721,N_9779);
nor UO_17 (O_17,N_9045,N_9361);
nor UO_18 (O_18,N_9298,N_9676);
xor UO_19 (O_19,N_9568,N_9802);
and UO_20 (O_20,N_9365,N_9673);
nand UO_21 (O_21,N_9879,N_9248);
or UO_22 (O_22,N_9807,N_9079);
nor UO_23 (O_23,N_9659,N_9446);
and UO_24 (O_24,N_9270,N_9326);
nor UO_25 (O_25,N_9155,N_9509);
or UO_26 (O_26,N_9465,N_9404);
or UO_27 (O_27,N_9768,N_9751);
and UO_28 (O_28,N_9088,N_9878);
nand UO_29 (O_29,N_9950,N_9967);
and UO_30 (O_30,N_9136,N_9975);
or UO_31 (O_31,N_9370,N_9631);
nand UO_32 (O_32,N_9012,N_9359);
or UO_33 (O_33,N_9418,N_9352);
and UO_34 (O_34,N_9702,N_9318);
nor UO_35 (O_35,N_9420,N_9691);
nand UO_36 (O_36,N_9201,N_9396);
nor UO_37 (O_37,N_9571,N_9819);
and UO_38 (O_38,N_9484,N_9667);
nor UO_39 (O_39,N_9372,N_9804);
or UO_40 (O_40,N_9905,N_9392);
xor UO_41 (O_41,N_9362,N_9683);
nor UO_42 (O_42,N_9853,N_9173);
nand UO_43 (O_43,N_9221,N_9407);
or UO_44 (O_44,N_9430,N_9250);
or UO_45 (O_45,N_9389,N_9314);
xor UO_46 (O_46,N_9160,N_9320);
xor UO_47 (O_47,N_9093,N_9939);
and UO_48 (O_48,N_9928,N_9463);
nor UO_49 (O_49,N_9954,N_9948);
and UO_50 (O_50,N_9639,N_9836);
nand UO_51 (O_51,N_9742,N_9785);
or UO_52 (O_52,N_9979,N_9888);
nor UO_53 (O_53,N_9215,N_9598);
nor UO_54 (O_54,N_9202,N_9771);
or UO_55 (O_55,N_9708,N_9044);
xor UO_56 (O_56,N_9651,N_9798);
or UO_57 (O_57,N_9360,N_9025);
and UO_58 (O_58,N_9374,N_9382);
and UO_59 (O_59,N_9772,N_9019);
nor UO_60 (O_60,N_9066,N_9006);
nor UO_61 (O_61,N_9086,N_9762);
nor UO_62 (O_62,N_9253,N_9722);
nand UO_63 (O_63,N_9514,N_9517);
and UO_64 (O_64,N_9901,N_9337);
xor UO_65 (O_65,N_9440,N_9100);
xor UO_66 (O_66,N_9706,N_9805);
or UO_67 (O_67,N_9255,N_9075);
nand UO_68 (O_68,N_9756,N_9870);
nor UO_69 (O_69,N_9048,N_9511);
nand UO_70 (O_70,N_9355,N_9628);
xor UO_71 (O_71,N_9774,N_9063);
nand UO_72 (O_72,N_9696,N_9941);
nor UO_73 (O_73,N_9497,N_9451);
nor UO_74 (O_74,N_9229,N_9765);
nand UO_75 (O_75,N_9653,N_9648);
nor UO_76 (O_76,N_9183,N_9922);
xnor UO_77 (O_77,N_9633,N_9748);
or UO_78 (O_78,N_9476,N_9310);
and UO_79 (O_79,N_9014,N_9992);
and UO_80 (O_80,N_9040,N_9490);
xnor UO_81 (O_81,N_9474,N_9307);
or UO_82 (O_82,N_9123,N_9760);
nor UO_83 (O_83,N_9290,N_9620);
xor UO_84 (O_84,N_9634,N_9029);
nor UO_85 (O_85,N_9055,N_9472);
nor UO_86 (O_86,N_9658,N_9577);
and UO_87 (O_87,N_9550,N_9883);
xnor UO_88 (O_88,N_9137,N_9458);
nand UO_89 (O_89,N_9234,N_9711);
or UO_90 (O_90,N_9138,N_9127);
xor UO_91 (O_91,N_9993,N_9512);
and UO_92 (O_92,N_9991,N_9064);
and UO_93 (O_93,N_9985,N_9946);
xnor UO_94 (O_94,N_9876,N_9847);
nor UO_95 (O_95,N_9841,N_9013);
and UO_96 (O_96,N_9723,N_9099);
and UO_97 (O_97,N_9333,N_9850);
nor UO_98 (O_98,N_9328,N_9945);
and UO_99 (O_99,N_9304,N_9165);
nor UO_100 (O_100,N_9397,N_9377);
and UO_101 (O_101,N_9564,N_9986);
or UO_102 (O_102,N_9583,N_9913);
nor UO_103 (O_103,N_9956,N_9289);
nor UO_104 (O_104,N_9726,N_9828);
nand UO_105 (O_105,N_9582,N_9505);
and UO_106 (O_106,N_9761,N_9146);
nand UO_107 (O_107,N_9910,N_9720);
and UO_108 (O_108,N_9800,N_9325);
nand UO_109 (O_109,N_9518,N_9830);
or UO_110 (O_110,N_9506,N_9741);
nand UO_111 (O_111,N_9553,N_9534);
and UO_112 (O_112,N_9070,N_9097);
nand UO_113 (O_113,N_9117,N_9790);
nand UO_114 (O_114,N_9996,N_9107);
or UO_115 (O_115,N_9252,N_9153);
or UO_116 (O_116,N_9411,N_9102);
nor UO_117 (O_117,N_9834,N_9461);
nor UO_118 (O_118,N_9031,N_9781);
and UO_119 (O_119,N_9695,N_9504);
xor UO_120 (O_120,N_9799,N_9116);
and UO_121 (O_121,N_9464,N_9664);
nand UO_122 (O_122,N_9618,N_9145);
xnor UO_123 (O_123,N_9849,N_9867);
nor UO_124 (O_124,N_9181,N_9965);
or UO_125 (O_125,N_9516,N_9459);
xnor UO_126 (O_126,N_9624,N_9424);
xnor UO_127 (O_127,N_9174,N_9533);
nand UO_128 (O_128,N_9488,N_9872);
and UO_129 (O_129,N_9258,N_9681);
nor UO_130 (O_130,N_9010,N_9990);
nor UO_131 (O_131,N_9843,N_9275);
nand UO_132 (O_132,N_9049,N_9570);
or UO_133 (O_133,N_9169,N_9077);
or UO_134 (O_134,N_9881,N_9487);
xnor UO_135 (O_135,N_9431,N_9644);
or UO_136 (O_136,N_9384,N_9429);
or UO_137 (O_137,N_9874,N_9749);
or UO_138 (O_138,N_9943,N_9230);
nor UO_139 (O_139,N_9225,N_9846);
and UO_140 (O_140,N_9262,N_9526);
and UO_141 (O_141,N_9053,N_9247);
nor UO_142 (O_142,N_9483,N_9052);
nand UO_143 (O_143,N_9192,N_9902);
nand UO_144 (O_144,N_9898,N_9311);
or UO_145 (O_145,N_9812,N_9606);
nand UO_146 (O_146,N_9890,N_9393);
nand UO_147 (O_147,N_9626,N_9641);
nand UO_148 (O_148,N_9560,N_9637);
xor UO_149 (O_149,N_9323,N_9629);
and UO_150 (O_150,N_9647,N_9441);
and UO_151 (O_151,N_9562,N_9338);
nor UO_152 (O_152,N_9635,N_9278);
nor UO_153 (O_153,N_9216,N_9521);
nor UO_154 (O_154,N_9203,N_9030);
and UO_155 (O_155,N_9886,N_9875);
xor UO_156 (O_156,N_9595,N_9095);
and UO_157 (O_157,N_9515,N_9732);
and UO_158 (O_158,N_9636,N_9468);
nand UO_159 (O_159,N_9575,N_9682);
nand UO_160 (O_160,N_9074,N_9198);
and UO_161 (O_161,N_9238,N_9873);
nand UO_162 (O_162,N_9957,N_9082);
or UO_163 (O_163,N_9027,N_9132);
nand UO_164 (O_164,N_9981,N_9940);
and UO_165 (O_165,N_9267,N_9037);
and UO_166 (O_166,N_9605,N_9232);
nor UO_167 (O_167,N_9268,N_9838);
and UO_168 (O_168,N_9880,N_9347);
nand UO_169 (O_169,N_9668,N_9690);
xor UO_170 (O_170,N_9306,N_9034);
xnor UO_171 (O_171,N_9661,N_9987);
nand UO_172 (O_172,N_9371,N_9716);
xnor UO_173 (O_173,N_9916,N_9108);
nand UO_174 (O_174,N_9921,N_9046);
and UO_175 (O_175,N_9477,N_9705);
or UO_176 (O_176,N_9851,N_9660);
nor UO_177 (O_177,N_9276,N_9535);
xnor UO_178 (O_178,N_9224,N_9241);
and UO_179 (O_179,N_9866,N_9433);
xnor UO_180 (O_180,N_9170,N_9735);
and UO_181 (O_181,N_9450,N_9601);
and UO_182 (O_182,N_9780,N_9909);
and UO_183 (O_183,N_9856,N_9000);
nand UO_184 (O_184,N_9933,N_9481);
nand UO_185 (O_185,N_9923,N_9291);
xor UO_186 (O_186,N_9822,N_9373);
xor UO_187 (O_187,N_9317,N_9151);
nand UO_188 (O_188,N_9150,N_9292);
xor UO_189 (O_189,N_9657,N_9508);
xor UO_190 (O_190,N_9500,N_9427);
nand UO_191 (O_191,N_9345,N_9071);
and UO_192 (O_192,N_9294,N_9689);
and UO_193 (O_193,N_9949,N_9194);
nor UO_194 (O_194,N_9478,N_9700);
nand UO_195 (O_195,N_9596,N_9211);
or UO_196 (O_196,N_9801,N_9630);
xor UO_197 (O_197,N_9810,N_9694);
nand UO_198 (O_198,N_9266,N_9817);
and UO_199 (O_199,N_9900,N_9640);
and UO_200 (O_200,N_9056,N_9593);
nor UO_201 (O_201,N_9114,N_9354);
and UO_202 (O_202,N_9832,N_9265);
xnor UO_203 (O_203,N_9784,N_9715);
or UO_204 (O_204,N_9416,N_9200);
nor UO_205 (O_205,N_9793,N_9914);
nand UO_206 (O_206,N_9861,N_9473);
xnor UO_207 (O_207,N_9541,N_9178);
nand UO_208 (O_208,N_9995,N_9316);
or UO_209 (O_209,N_9809,N_9558);
or UO_210 (O_210,N_9597,N_9662);
xor UO_211 (O_211,N_9513,N_9067);
nor UO_212 (O_212,N_9054,N_9960);
or UO_213 (O_213,N_9693,N_9523);
or UO_214 (O_214,N_9972,N_9971);
or UO_215 (O_215,N_9443,N_9161);
nor UO_216 (O_216,N_9962,N_9520);
xor UO_217 (O_217,N_9725,N_9144);
nor UO_218 (O_218,N_9764,N_9346);
or UO_219 (O_219,N_9091,N_9530);
xnor UO_220 (O_220,N_9754,N_9273);
and UO_221 (O_221,N_9296,N_9899);
or UO_222 (O_222,N_9281,N_9154);
or UO_223 (O_223,N_9727,N_9023);
xor UO_224 (O_224,N_9988,N_9588);
nor UO_225 (O_225,N_9061,N_9084);
nor UO_226 (O_226,N_9402,N_9669);
xor UO_227 (O_227,N_9206,N_9332);
xor UO_228 (O_228,N_9356,N_9134);
or UO_229 (O_229,N_9501,N_9112);
nor UO_230 (O_230,N_9747,N_9018);
xor UO_231 (O_231,N_9643,N_9894);
or UO_232 (O_232,N_9222,N_9058);
or UO_233 (O_233,N_9493,N_9042);
and UO_234 (O_234,N_9403,N_9120);
and UO_235 (O_235,N_9240,N_9139);
and UO_236 (O_236,N_9734,N_9237);
nand UO_237 (O_237,N_9287,N_9329);
or UO_238 (O_238,N_9001,N_9769);
or UO_239 (O_239,N_9563,N_9622);
xnor UO_240 (O_240,N_9740,N_9953);
nor UO_241 (O_241,N_9554,N_9891);
or UO_242 (O_242,N_9692,N_9341);
nor UO_243 (O_243,N_9005,N_9565);
and UO_244 (O_244,N_9621,N_9759);
nand UO_245 (O_245,N_9586,N_9024);
xnor UO_246 (O_246,N_9567,N_9831);
xnor UO_247 (O_247,N_9714,N_9090);
nand UO_248 (O_248,N_9409,N_9572);
xnor UO_249 (O_249,N_9439,N_9806);
and UO_250 (O_250,N_9701,N_9911);
nand UO_251 (O_251,N_9897,N_9434);
or UO_252 (O_252,N_9984,N_9531);
and UO_253 (O_253,N_9590,N_9816);
xor UO_254 (O_254,N_9186,N_9792);
and UO_255 (O_255,N_9363,N_9955);
nand UO_256 (O_256,N_9733,N_9111);
xnor UO_257 (O_257,N_9185,N_9105);
nor UO_258 (O_258,N_9686,N_9193);
xor UO_259 (O_259,N_9475,N_9813);
nand UO_260 (O_260,N_9350,N_9574);
and UO_261 (O_261,N_9286,N_9863);
nand UO_262 (O_262,N_9896,N_9918);
or UO_263 (O_263,N_9730,N_9188);
nor UO_264 (O_264,N_9315,N_9978);
xnor UO_265 (O_265,N_9348,N_9226);
xor UO_266 (O_266,N_9724,N_9118);
nor UO_267 (O_267,N_9983,N_9495);
nand UO_268 (O_268,N_9825,N_9743);
nand UO_269 (O_269,N_9162,N_9398);
or UO_270 (O_270,N_9094,N_9213);
nand UO_271 (O_271,N_9655,N_9786);
or UO_272 (O_272,N_9164,N_9449);
xnor UO_273 (O_273,N_9559,N_9737);
nor UO_274 (O_274,N_9426,N_9448);
nor UO_275 (O_275,N_9613,N_9524);
xor UO_276 (O_276,N_9770,N_9710);
nor UO_277 (O_277,N_9994,N_9645);
and UO_278 (O_278,N_9608,N_9915);
nor UO_279 (O_279,N_9158,N_9674);
xnor UO_280 (O_280,N_9085,N_9378);
nor UO_281 (O_281,N_9002,N_9947);
xnor UO_282 (O_282,N_9050,N_9453);
nor UO_283 (O_283,N_9189,N_9904);
nor UO_284 (O_284,N_9125,N_9297);
and UO_285 (O_285,N_9435,N_9794);
nor UO_286 (O_286,N_9385,N_9833);
or UO_287 (O_287,N_9078,N_9231);
nor UO_288 (O_288,N_9197,N_9652);
or UO_289 (O_289,N_9376,N_9157);
nor UO_290 (O_290,N_9103,N_9903);
xor UO_291 (O_291,N_9322,N_9854);
and UO_292 (O_292,N_9489,N_9869);
or UO_293 (O_293,N_9339,N_9199);
or UO_294 (O_294,N_9062,N_9815);
nor UO_295 (O_295,N_9998,N_9485);
nor UO_296 (O_296,N_9386,N_9599);
xor UO_297 (O_297,N_9457,N_9379);
and UO_298 (O_298,N_9060,N_9209);
or UO_299 (O_299,N_9412,N_9142);
nor UO_300 (O_300,N_9930,N_9579);
and UO_301 (O_301,N_9607,N_9961);
nor UO_302 (O_302,N_9039,N_9491);
xnor UO_303 (O_303,N_9739,N_9351);
and UO_304 (O_304,N_9387,N_9619);
and UO_305 (O_305,N_9728,N_9008);
nand UO_306 (O_306,N_9551,N_9542);
or UO_307 (O_307,N_9456,N_9499);
nand UO_308 (O_308,N_9009,N_9210);
and UO_309 (O_309,N_9228,N_9602);
or UO_310 (O_310,N_9697,N_9340);
or UO_311 (O_311,N_9750,N_9038);
and UO_312 (O_312,N_9395,N_9835);
or UO_313 (O_313,N_9823,N_9787);
nor UO_314 (O_314,N_9121,N_9207);
or UO_315 (O_315,N_9249,N_9783);
xnor UO_316 (O_316,N_9122,N_9791);
and UO_317 (O_317,N_9445,N_9581);
xor UO_318 (O_318,N_9217,N_9358);
nand UO_319 (O_319,N_9180,N_9679);
and UO_320 (O_320,N_9140,N_9587);
and UO_321 (O_321,N_9410,N_9566);
nand UO_322 (O_322,N_9591,N_9615);
and UO_323 (O_323,N_9452,N_9096);
nor UO_324 (O_324,N_9623,N_9130);
or UO_325 (O_325,N_9738,N_9803);
and UO_326 (O_326,N_9980,N_9080);
or UO_327 (O_327,N_9388,N_9383);
nand UO_328 (O_328,N_9663,N_9036);
nor UO_329 (O_329,N_9280,N_9131);
nand UO_330 (O_330,N_9935,N_9442);
nand UO_331 (O_331,N_9343,N_9007);
nand UO_332 (O_332,N_9758,N_9646);
nand UO_333 (O_333,N_9889,N_9254);
or UO_334 (O_334,N_9149,N_9675);
and UO_335 (O_335,N_9011,N_9471);
nor UO_336 (O_336,N_9503,N_9952);
nor UO_337 (O_337,N_9767,N_9892);
nor UO_338 (O_338,N_9380,N_9614);
and UO_339 (O_339,N_9908,N_9126);
xnor UO_340 (O_340,N_9507,N_9537);
nor UO_341 (O_341,N_9244,N_9982);
xnor UO_342 (O_342,N_9642,N_9366);
or UO_343 (O_343,N_9844,N_9604);
nand UO_344 (O_344,N_9245,N_9865);
nor UO_345 (O_345,N_9305,N_9919);
or UO_346 (O_346,N_9437,N_9405);
nand UO_347 (O_347,N_9837,N_9788);
or UO_348 (O_348,N_9552,N_9147);
nand UO_349 (O_349,N_9677,N_9089);
nand UO_350 (O_350,N_9617,N_9547);
xor UO_351 (O_351,N_9110,N_9576);
or UO_352 (O_352,N_9818,N_9482);
or UO_353 (O_353,N_9035,N_9109);
xnor UO_354 (O_354,N_9059,N_9375);
and UO_355 (O_355,N_9494,N_9775);
nand UO_356 (O_356,N_9808,N_9492);
and UO_357 (O_357,N_9033,N_9589);
xnor UO_358 (O_358,N_9745,N_9707);
xor UO_359 (O_359,N_9649,N_9616);
xnor UO_360 (O_360,N_9303,N_9274);
nor UO_361 (O_361,N_9580,N_9549);
nor UO_362 (O_362,N_9444,N_9187);
or UO_363 (O_363,N_9143,N_9729);
xnor UO_364 (O_364,N_9428,N_9963);
and UO_365 (O_365,N_9133,N_9288);
nor UO_366 (O_366,N_9259,N_9974);
nor UO_367 (O_367,N_9795,N_9083);
xor UO_368 (O_368,N_9295,N_9319);
xor UO_369 (O_369,N_9864,N_9666);
nor UO_370 (O_370,N_9308,N_9330);
xor UO_371 (O_371,N_9251,N_9175);
nor UO_372 (O_372,N_9796,N_9717);
nand UO_373 (O_373,N_9842,N_9709);
nor UO_374 (O_374,N_9284,N_9736);
xnor UO_375 (O_375,N_9032,N_9855);
and UO_376 (O_376,N_9797,N_9260);
or UO_377 (O_377,N_9124,N_9313);
or UO_378 (O_378,N_9882,N_9051);
or UO_379 (O_379,N_9925,N_9525);
and UO_380 (O_380,N_9196,N_9519);
nor UO_381 (O_381,N_9092,N_9191);
or UO_382 (O_382,N_9585,N_9219);
and UO_383 (O_383,N_9934,N_9968);
and UO_384 (O_384,N_9556,N_9753);
and UO_385 (O_385,N_9177,N_9532);
nand UO_386 (O_386,N_9827,N_9159);
nand UO_387 (O_387,N_9885,N_9282);
nand UO_388 (O_388,N_9684,N_9166);
xor UO_389 (O_389,N_9859,N_9069);
xor UO_390 (O_390,N_9421,N_9415);
or UO_391 (O_391,N_9858,N_9912);
nor UO_392 (O_392,N_9073,N_9182);
nor UO_393 (O_393,N_9924,N_9820);
xnor UO_394 (O_394,N_9205,N_9043);
and UO_395 (O_395,N_9357,N_9269);
nand UO_396 (O_396,N_9824,N_9301);
xor UO_397 (O_397,N_9964,N_9068);
xnor UO_398 (O_398,N_9632,N_9862);
nor UO_399 (O_399,N_9293,N_9777);
nor UO_400 (O_400,N_9003,N_9860);
or UO_401 (O_401,N_9168,N_9335);
and UO_402 (O_402,N_9680,N_9746);
nor UO_403 (O_403,N_9171,N_9821);
nand UO_404 (O_404,N_9573,N_9528);
or UO_405 (O_405,N_9406,N_9522);
or UO_406 (O_406,N_9264,N_9973);
xor UO_407 (O_407,N_9022,N_9479);
or UO_408 (O_408,N_9977,N_9413);
xnor UO_409 (O_409,N_9208,N_9462);
xor UO_410 (O_410,N_9119,N_9256);
or UO_411 (O_411,N_9243,N_9713);
nor UO_412 (O_412,N_9277,N_9929);
or UO_413 (O_413,N_9546,N_9454);
nor UO_414 (O_414,N_9047,N_9312);
and UO_415 (O_415,N_9129,N_9887);
xnor UO_416 (O_416,N_9218,N_9331);
xnor UO_417 (O_417,N_9283,N_9246);
nor UO_418 (O_418,N_9938,N_9538);
xor UO_419 (O_419,N_9195,N_9015);
nor UO_420 (O_420,N_9778,N_9712);
xnor UO_421 (O_421,N_9300,N_9755);
xnor UO_422 (O_422,N_9381,N_9271);
and UO_423 (O_423,N_9204,N_9327);
and UO_424 (O_424,N_9937,N_9017);
or UO_425 (O_425,N_9906,N_9704);
nor UO_426 (O_426,N_9414,N_9212);
xor UO_427 (O_427,N_9757,N_9496);
or UO_428 (O_428,N_9455,N_9561);
nand UO_429 (O_429,N_9612,N_9344);
nand UO_430 (O_430,N_9555,N_9104);
and UO_431 (O_431,N_9460,N_9970);
nand UO_432 (O_432,N_9285,N_9548);
xnor UO_433 (O_433,N_9242,N_9239);
or UO_434 (O_434,N_9163,N_9076);
or UO_435 (O_435,N_9884,N_9467);
or UO_436 (O_436,N_9400,N_9877);
and UO_437 (O_437,N_9544,N_9098);
xor UO_438 (O_438,N_9951,N_9917);
xnor UO_439 (O_439,N_9419,N_9026);
or UO_440 (O_440,N_9141,N_9510);
xor UO_441 (O_441,N_9190,N_9976);
nor UO_442 (O_442,N_9353,N_9703);
and UO_443 (O_443,N_9057,N_9447);
xnor UO_444 (O_444,N_9600,N_9028);
xor UO_445 (O_445,N_9021,N_9172);
nand UO_446 (O_446,N_9364,N_9789);
and UO_447 (O_447,N_9368,N_9272);
nand UO_448 (O_448,N_9989,N_9152);
or UO_449 (O_449,N_9678,N_9650);
and UO_450 (O_450,N_9936,N_9969);
nand UO_451 (O_451,N_9698,N_9502);
nand UO_452 (O_452,N_9004,N_9081);
and UO_453 (O_453,N_9763,N_9438);
and UO_454 (O_454,N_9719,N_9625);
and UO_455 (O_455,N_9826,N_9603);
and UO_456 (O_456,N_9656,N_9020);
and UO_457 (O_457,N_9672,N_9671);
or UO_458 (O_458,N_9334,N_9773);
xor UO_459 (O_459,N_9148,N_9432);
nor UO_460 (O_460,N_9932,N_9113);
nor UO_461 (O_461,N_9927,N_9744);
or UO_462 (O_462,N_9857,N_9299);
xnor UO_463 (O_463,N_9766,N_9342);
nand UO_464 (O_464,N_9220,N_9944);
and UO_465 (O_465,N_9638,N_9718);
and UO_466 (O_466,N_9699,N_9156);
or UO_467 (O_467,N_9399,N_9106);
xnor UO_468 (O_468,N_9997,N_9840);
and UO_469 (O_469,N_9423,N_9569);
nand UO_470 (O_470,N_9839,N_9336);
or UO_471 (O_471,N_9417,N_9115);
xnor UO_472 (O_472,N_9895,N_9999);
xnor UO_473 (O_473,N_9369,N_9609);
xor UO_474 (O_474,N_9687,N_9041);
and UO_475 (O_475,N_9394,N_9782);
nor UO_476 (O_476,N_9233,N_9868);
and UO_477 (O_477,N_9665,N_9236);
xor UO_478 (O_478,N_9469,N_9261);
xnor UO_479 (O_479,N_9470,N_9931);
xor UO_480 (O_480,N_9436,N_9425);
and UO_481 (O_481,N_9959,N_9128);
and UO_482 (O_482,N_9829,N_9610);
and UO_483 (O_483,N_9486,N_9324);
nor UO_484 (O_484,N_9545,N_9065);
nor UO_485 (O_485,N_9871,N_9611);
nand UO_486 (O_486,N_9685,N_9401);
nor UO_487 (O_487,N_9527,N_9349);
nor UO_488 (O_488,N_9920,N_9845);
or UO_489 (O_489,N_9852,N_9670);
and UO_490 (O_490,N_9072,N_9539);
or UO_491 (O_491,N_9536,N_9814);
or UO_492 (O_492,N_9731,N_9529);
nand UO_493 (O_493,N_9592,N_9958);
xor UO_494 (O_494,N_9263,N_9179);
nor UO_495 (O_495,N_9466,N_9966);
nor UO_496 (O_496,N_9176,N_9848);
xnor UO_497 (O_497,N_9498,N_9214);
xnor UO_498 (O_498,N_9540,N_9408);
xor UO_499 (O_499,N_9893,N_9223);
and UO_500 (O_500,N_9554,N_9475);
nand UO_501 (O_501,N_9713,N_9266);
and UO_502 (O_502,N_9220,N_9741);
nand UO_503 (O_503,N_9538,N_9940);
nor UO_504 (O_504,N_9068,N_9347);
or UO_505 (O_505,N_9460,N_9785);
and UO_506 (O_506,N_9913,N_9320);
xnor UO_507 (O_507,N_9344,N_9531);
nand UO_508 (O_508,N_9200,N_9782);
nor UO_509 (O_509,N_9810,N_9547);
nor UO_510 (O_510,N_9502,N_9650);
or UO_511 (O_511,N_9909,N_9479);
and UO_512 (O_512,N_9491,N_9185);
or UO_513 (O_513,N_9084,N_9320);
or UO_514 (O_514,N_9677,N_9845);
nor UO_515 (O_515,N_9860,N_9668);
xnor UO_516 (O_516,N_9015,N_9530);
xnor UO_517 (O_517,N_9564,N_9298);
nor UO_518 (O_518,N_9895,N_9067);
nand UO_519 (O_519,N_9966,N_9753);
xor UO_520 (O_520,N_9288,N_9261);
and UO_521 (O_521,N_9010,N_9287);
and UO_522 (O_522,N_9425,N_9910);
or UO_523 (O_523,N_9540,N_9641);
xor UO_524 (O_524,N_9748,N_9696);
and UO_525 (O_525,N_9489,N_9478);
and UO_526 (O_526,N_9532,N_9295);
nor UO_527 (O_527,N_9303,N_9923);
and UO_528 (O_528,N_9517,N_9267);
nor UO_529 (O_529,N_9653,N_9168);
nor UO_530 (O_530,N_9064,N_9449);
and UO_531 (O_531,N_9074,N_9578);
or UO_532 (O_532,N_9937,N_9778);
xnor UO_533 (O_533,N_9494,N_9541);
or UO_534 (O_534,N_9508,N_9616);
or UO_535 (O_535,N_9578,N_9127);
and UO_536 (O_536,N_9523,N_9941);
nand UO_537 (O_537,N_9931,N_9286);
nand UO_538 (O_538,N_9831,N_9974);
xor UO_539 (O_539,N_9129,N_9621);
xnor UO_540 (O_540,N_9725,N_9762);
nand UO_541 (O_541,N_9277,N_9354);
nand UO_542 (O_542,N_9380,N_9876);
xor UO_543 (O_543,N_9520,N_9001);
or UO_544 (O_544,N_9917,N_9520);
and UO_545 (O_545,N_9909,N_9296);
xnor UO_546 (O_546,N_9579,N_9055);
or UO_547 (O_547,N_9422,N_9574);
nand UO_548 (O_548,N_9930,N_9359);
nand UO_549 (O_549,N_9992,N_9199);
and UO_550 (O_550,N_9716,N_9302);
or UO_551 (O_551,N_9135,N_9774);
or UO_552 (O_552,N_9460,N_9653);
nor UO_553 (O_553,N_9755,N_9008);
xnor UO_554 (O_554,N_9736,N_9902);
and UO_555 (O_555,N_9409,N_9441);
nand UO_556 (O_556,N_9460,N_9673);
or UO_557 (O_557,N_9234,N_9743);
nor UO_558 (O_558,N_9817,N_9690);
xor UO_559 (O_559,N_9616,N_9101);
or UO_560 (O_560,N_9645,N_9150);
xor UO_561 (O_561,N_9510,N_9519);
or UO_562 (O_562,N_9103,N_9348);
nor UO_563 (O_563,N_9648,N_9340);
nand UO_564 (O_564,N_9289,N_9584);
nand UO_565 (O_565,N_9230,N_9459);
nand UO_566 (O_566,N_9676,N_9412);
nor UO_567 (O_567,N_9511,N_9545);
or UO_568 (O_568,N_9782,N_9282);
or UO_569 (O_569,N_9664,N_9441);
nor UO_570 (O_570,N_9916,N_9873);
or UO_571 (O_571,N_9777,N_9207);
or UO_572 (O_572,N_9404,N_9098);
nand UO_573 (O_573,N_9200,N_9216);
or UO_574 (O_574,N_9727,N_9990);
xnor UO_575 (O_575,N_9763,N_9437);
nor UO_576 (O_576,N_9232,N_9730);
nor UO_577 (O_577,N_9152,N_9490);
or UO_578 (O_578,N_9990,N_9717);
nor UO_579 (O_579,N_9900,N_9776);
and UO_580 (O_580,N_9855,N_9931);
and UO_581 (O_581,N_9298,N_9427);
or UO_582 (O_582,N_9875,N_9390);
nor UO_583 (O_583,N_9972,N_9773);
nor UO_584 (O_584,N_9756,N_9941);
xor UO_585 (O_585,N_9157,N_9413);
and UO_586 (O_586,N_9362,N_9364);
nor UO_587 (O_587,N_9265,N_9994);
nor UO_588 (O_588,N_9164,N_9465);
nand UO_589 (O_589,N_9325,N_9951);
xnor UO_590 (O_590,N_9340,N_9910);
or UO_591 (O_591,N_9105,N_9268);
nand UO_592 (O_592,N_9008,N_9306);
xor UO_593 (O_593,N_9233,N_9990);
or UO_594 (O_594,N_9721,N_9976);
or UO_595 (O_595,N_9271,N_9308);
nor UO_596 (O_596,N_9023,N_9504);
nor UO_597 (O_597,N_9331,N_9696);
nand UO_598 (O_598,N_9948,N_9150);
nand UO_599 (O_599,N_9229,N_9183);
xnor UO_600 (O_600,N_9030,N_9177);
and UO_601 (O_601,N_9976,N_9354);
nand UO_602 (O_602,N_9791,N_9261);
xnor UO_603 (O_603,N_9430,N_9830);
or UO_604 (O_604,N_9603,N_9052);
xor UO_605 (O_605,N_9305,N_9535);
and UO_606 (O_606,N_9630,N_9070);
xor UO_607 (O_607,N_9167,N_9688);
xnor UO_608 (O_608,N_9842,N_9765);
and UO_609 (O_609,N_9484,N_9406);
and UO_610 (O_610,N_9012,N_9081);
and UO_611 (O_611,N_9784,N_9996);
or UO_612 (O_612,N_9944,N_9321);
and UO_613 (O_613,N_9275,N_9197);
or UO_614 (O_614,N_9929,N_9549);
nand UO_615 (O_615,N_9233,N_9712);
nor UO_616 (O_616,N_9630,N_9960);
and UO_617 (O_617,N_9803,N_9971);
and UO_618 (O_618,N_9254,N_9394);
and UO_619 (O_619,N_9564,N_9550);
xor UO_620 (O_620,N_9569,N_9682);
xor UO_621 (O_621,N_9911,N_9402);
nand UO_622 (O_622,N_9421,N_9325);
nor UO_623 (O_623,N_9824,N_9852);
nor UO_624 (O_624,N_9416,N_9858);
and UO_625 (O_625,N_9683,N_9881);
nor UO_626 (O_626,N_9165,N_9665);
xor UO_627 (O_627,N_9180,N_9028);
nand UO_628 (O_628,N_9955,N_9683);
and UO_629 (O_629,N_9054,N_9738);
or UO_630 (O_630,N_9239,N_9314);
and UO_631 (O_631,N_9610,N_9341);
or UO_632 (O_632,N_9971,N_9097);
nand UO_633 (O_633,N_9086,N_9930);
or UO_634 (O_634,N_9752,N_9615);
nor UO_635 (O_635,N_9828,N_9387);
or UO_636 (O_636,N_9456,N_9415);
nand UO_637 (O_637,N_9370,N_9629);
nand UO_638 (O_638,N_9026,N_9853);
xnor UO_639 (O_639,N_9251,N_9124);
nor UO_640 (O_640,N_9862,N_9137);
and UO_641 (O_641,N_9641,N_9093);
and UO_642 (O_642,N_9101,N_9823);
nor UO_643 (O_643,N_9541,N_9654);
nand UO_644 (O_644,N_9560,N_9511);
xnor UO_645 (O_645,N_9849,N_9394);
and UO_646 (O_646,N_9106,N_9991);
and UO_647 (O_647,N_9149,N_9789);
nor UO_648 (O_648,N_9968,N_9340);
or UO_649 (O_649,N_9048,N_9200);
and UO_650 (O_650,N_9599,N_9087);
nand UO_651 (O_651,N_9138,N_9129);
and UO_652 (O_652,N_9993,N_9214);
or UO_653 (O_653,N_9413,N_9920);
nor UO_654 (O_654,N_9815,N_9634);
nand UO_655 (O_655,N_9162,N_9674);
xor UO_656 (O_656,N_9623,N_9371);
nand UO_657 (O_657,N_9597,N_9710);
xor UO_658 (O_658,N_9200,N_9342);
or UO_659 (O_659,N_9411,N_9812);
nor UO_660 (O_660,N_9861,N_9864);
xor UO_661 (O_661,N_9485,N_9261);
nor UO_662 (O_662,N_9137,N_9592);
nand UO_663 (O_663,N_9071,N_9594);
nor UO_664 (O_664,N_9323,N_9843);
nand UO_665 (O_665,N_9972,N_9621);
xnor UO_666 (O_666,N_9984,N_9209);
or UO_667 (O_667,N_9416,N_9744);
or UO_668 (O_668,N_9083,N_9945);
or UO_669 (O_669,N_9972,N_9912);
nor UO_670 (O_670,N_9749,N_9038);
and UO_671 (O_671,N_9782,N_9256);
nor UO_672 (O_672,N_9879,N_9393);
or UO_673 (O_673,N_9696,N_9736);
xor UO_674 (O_674,N_9047,N_9768);
nor UO_675 (O_675,N_9643,N_9594);
xor UO_676 (O_676,N_9805,N_9702);
xor UO_677 (O_677,N_9152,N_9583);
or UO_678 (O_678,N_9670,N_9082);
xor UO_679 (O_679,N_9362,N_9681);
and UO_680 (O_680,N_9876,N_9043);
xnor UO_681 (O_681,N_9255,N_9114);
xnor UO_682 (O_682,N_9505,N_9718);
nor UO_683 (O_683,N_9749,N_9847);
xnor UO_684 (O_684,N_9819,N_9017);
or UO_685 (O_685,N_9464,N_9205);
xnor UO_686 (O_686,N_9313,N_9705);
xnor UO_687 (O_687,N_9825,N_9653);
and UO_688 (O_688,N_9410,N_9795);
xnor UO_689 (O_689,N_9301,N_9705);
or UO_690 (O_690,N_9501,N_9937);
nand UO_691 (O_691,N_9277,N_9827);
or UO_692 (O_692,N_9910,N_9372);
or UO_693 (O_693,N_9948,N_9504);
nand UO_694 (O_694,N_9704,N_9079);
or UO_695 (O_695,N_9409,N_9828);
or UO_696 (O_696,N_9507,N_9320);
or UO_697 (O_697,N_9940,N_9212);
nor UO_698 (O_698,N_9110,N_9977);
or UO_699 (O_699,N_9610,N_9276);
xor UO_700 (O_700,N_9285,N_9807);
nor UO_701 (O_701,N_9910,N_9719);
xnor UO_702 (O_702,N_9722,N_9836);
or UO_703 (O_703,N_9853,N_9952);
and UO_704 (O_704,N_9792,N_9282);
or UO_705 (O_705,N_9434,N_9824);
and UO_706 (O_706,N_9634,N_9098);
nor UO_707 (O_707,N_9321,N_9436);
nor UO_708 (O_708,N_9995,N_9781);
and UO_709 (O_709,N_9441,N_9328);
xor UO_710 (O_710,N_9429,N_9005);
nand UO_711 (O_711,N_9605,N_9456);
and UO_712 (O_712,N_9291,N_9157);
or UO_713 (O_713,N_9337,N_9597);
xor UO_714 (O_714,N_9666,N_9931);
and UO_715 (O_715,N_9742,N_9017);
xor UO_716 (O_716,N_9478,N_9886);
nor UO_717 (O_717,N_9182,N_9476);
xor UO_718 (O_718,N_9580,N_9481);
and UO_719 (O_719,N_9203,N_9105);
nor UO_720 (O_720,N_9089,N_9771);
and UO_721 (O_721,N_9767,N_9184);
xor UO_722 (O_722,N_9161,N_9249);
xnor UO_723 (O_723,N_9530,N_9589);
or UO_724 (O_724,N_9554,N_9500);
or UO_725 (O_725,N_9526,N_9458);
or UO_726 (O_726,N_9880,N_9580);
nor UO_727 (O_727,N_9626,N_9829);
xor UO_728 (O_728,N_9507,N_9312);
xor UO_729 (O_729,N_9074,N_9489);
and UO_730 (O_730,N_9403,N_9847);
and UO_731 (O_731,N_9954,N_9484);
or UO_732 (O_732,N_9503,N_9939);
nor UO_733 (O_733,N_9826,N_9751);
or UO_734 (O_734,N_9549,N_9403);
nor UO_735 (O_735,N_9951,N_9139);
nand UO_736 (O_736,N_9397,N_9287);
or UO_737 (O_737,N_9099,N_9805);
xor UO_738 (O_738,N_9788,N_9533);
or UO_739 (O_739,N_9009,N_9459);
nor UO_740 (O_740,N_9158,N_9675);
and UO_741 (O_741,N_9125,N_9777);
and UO_742 (O_742,N_9218,N_9961);
xor UO_743 (O_743,N_9134,N_9667);
nor UO_744 (O_744,N_9341,N_9850);
nor UO_745 (O_745,N_9741,N_9201);
xor UO_746 (O_746,N_9513,N_9535);
or UO_747 (O_747,N_9297,N_9732);
nor UO_748 (O_748,N_9357,N_9028);
nor UO_749 (O_749,N_9575,N_9195);
nor UO_750 (O_750,N_9717,N_9627);
nand UO_751 (O_751,N_9914,N_9390);
xnor UO_752 (O_752,N_9973,N_9351);
xor UO_753 (O_753,N_9994,N_9129);
xor UO_754 (O_754,N_9075,N_9249);
or UO_755 (O_755,N_9288,N_9371);
nand UO_756 (O_756,N_9016,N_9631);
nand UO_757 (O_757,N_9789,N_9628);
nor UO_758 (O_758,N_9897,N_9191);
or UO_759 (O_759,N_9738,N_9466);
xor UO_760 (O_760,N_9034,N_9510);
or UO_761 (O_761,N_9979,N_9052);
or UO_762 (O_762,N_9867,N_9283);
or UO_763 (O_763,N_9220,N_9236);
nand UO_764 (O_764,N_9287,N_9016);
and UO_765 (O_765,N_9604,N_9938);
and UO_766 (O_766,N_9552,N_9604);
or UO_767 (O_767,N_9359,N_9508);
nor UO_768 (O_768,N_9878,N_9152);
or UO_769 (O_769,N_9607,N_9753);
and UO_770 (O_770,N_9437,N_9585);
or UO_771 (O_771,N_9699,N_9487);
xor UO_772 (O_772,N_9507,N_9533);
or UO_773 (O_773,N_9241,N_9732);
or UO_774 (O_774,N_9037,N_9232);
xnor UO_775 (O_775,N_9393,N_9588);
and UO_776 (O_776,N_9416,N_9755);
or UO_777 (O_777,N_9021,N_9537);
nor UO_778 (O_778,N_9156,N_9584);
xnor UO_779 (O_779,N_9184,N_9651);
nor UO_780 (O_780,N_9225,N_9210);
nand UO_781 (O_781,N_9952,N_9339);
xor UO_782 (O_782,N_9743,N_9178);
nor UO_783 (O_783,N_9628,N_9669);
nand UO_784 (O_784,N_9782,N_9776);
nor UO_785 (O_785,N_9569,N_9269);
nor UO_786 (O_786,N_9833,N_9267);
or UO_787 (O_787,N_9898,N_9771);
nor UO_788 (O_788,N_9898,N_9620);
nand UO_789 (O_789,N_9961,N_9684);
xnor UO_790 (O_790,N_9026,N_9569);
or UO_791 (O_791,N_9329,N_9105);
or UO_792 (O_792,N_9569,N_9927);
xor UO_793 (O_793,N_9994,N_9089);
and UO_794 (O_794,N_9652,N_9568);
and UO_795 (O_795,N_9383,N_9607);
or UO_796 (O_796,N_9630,N_9738);
xnor UO_797 (O_797,N_9129,N_9598);
and UO_798 (O_798,N_9562,N_9505);
and UO_799 (O_799,N_9406,N_9695);
nor UO_800 (O_800,N_9033,N_9925);
or UO_801 (O_801,N_9828,N_9020);
or UO_802 (O_802,N_9445,N_9885);
xor UO_803 (O_803,N_9077,N_9563);
and UO_804 (O_804,N_9906,N_9957);
xnor UO_805 (O_805,N_9564,N_9657);
xnor UO_806 (O_806,N_9141,N_9659);
nor UO_807 (O_807,N_9793,N_9046);
xor UO_808 (O_808,N_9008,N_9251);
nand UO_809 (O_809,N_9097,N_9333);
or UO_810 (O_810,N_9010,N_9930);
and UO_811 (O_811,N_9747,N_9243);
nor UO_812 (O_812,N_9685,N_9980);
nor UO_813 (O_813,N_9530,N_9182);
nor UO_814 (O_814,N_9377,N_9612);
and UO_815 (O_815,N_9228,N_9387);
nand UO_816 (O_816,N_9016,N_9695);
nor UO_817 (O_817,N_9418,N_9632);
nor UO_818 (O_818,N_9612,N_9917);
nor UO_819 (O_819,N_9663,N_9912);
or UO_820 (O_820,N_9911,N_9743);
nor UO_821 (O_821,N_9532,N_9523);
nor UO_822 (O_822,N_9685,N_9145);
nor UO_823 (O_823,N_9966,N_9831);
xor UO_824 (O_824,N_9012,N_9730);
nand UO_825 (O_825,N_9388,N_9178);
nand UO_826 (O_826,N_9922,N_9896);
nor UO_827 (O_827,N_9096,N_9465);
or UO_828 (O_828,N_9112,N_9091);
and UO_829 (O_829,N_9855,N_9662);
and UO_830 (O_830,N_9781,N_9065);
nor UO_831 (O_831,N_9974,N_9779);
nor UO_832 (O_832,N_9683,N_9191);
xor UO_833 (O_833,N_9308,N_9558);
nor UO_834 (O_834,N_9729,N_9454);
or UO_835 (O_835,N_9613,N_9705);
and UO_836 (O_836,N_9776,N_9537);
xor UO_837 (O_837,N_9161,N_9054);
nor UO_838 (O_838,N_9776,N_9945);
nor UO_839 (O_839,N_9466,N_9139);
nand UO_840 (O_840,N_9238,N_9396);
or UO_841 (O_841,N_9972,N_9055);
xor UO_842 (O_842,N_9481,N_9795);
or UO_843 (O_843,N_9288,N_9173);
nand UO_844 (O_844,N_9485,N_9427);
and UO_845 (O_845,N_9003,N_9891);
nor UO_846 (O_846,N_9263,N_9958);
or UO_847 (O_847,N_9976,N_9307);
and UO_848 (O_848,N_9309,N_9186);
nand UO_849 (O_849,N_9073,N_9054);
nand UO_850 (O_850,N_9293,N_9970);
nand UO_851 (O_851,N_9406,N_9355);
nor UO_852 (O_852,N_9092,N_9599);
and UO_853 (O_853,N_9296,N_9442);
and UO_854 (O_854,N_9572,N_9603);
xnor UO_855 (O_855,N_9726,N_9632);
nand UO_856 (O_856,N_9510,N_9642);
xnor UO_857 (O_857,N_9440,N_9579);
nor UO_858 (O_858,N_9223,N_9651);
or UO_859 (O_859,N_9661,N_9441);
and UO_860 (O_860,N_9931,N_9099);
or UO_861 (O_861,N_9884,N_9451);
and UO_862 (O_862,N_9372,N_9218);
nor UO_863 (O_863,N_9890,N_9622);
xnor UO_864 (O_864,N_9470,N_9670);
nor UO_865 (O_865,N_9831,N_9335);
or UO_866 (O_866,N_9232,N_9239);
nand UO_867 (O_867,N_9442,N_9652);
or UO_868 (O_868,N_9432,N_9921);
nand UO_869 (O_869,N_9906,N_9813);
and UO_870 (O_870,N_9206,N_9308);
or UO_871 (O_871,N_9436,N_9379);
and UO_872 (O_872,N_9329,N_9688);
and UO_873 (O_873,N_9131,N_9215);
nor UO_874 (O_874,N_9741,N_9429);
nand UO_875 (O_875,N_9796,N_9154);
nor UO_876 (O_876,N_9877,N_9656);
or UO_877 (O_877,N_9238,N_9781);
nor UO_878 (O_878,N_9082,N_9063);
and UO_879 (O_879,N_9235,N_9210);
nand UO_880 (O_880,N_9817,N_9841);
or UO_881 (O_881,N_9454,N_9713);
nor UO_882 (O_882,N_9671,N_9483);
xor UO_883 (O_883,N_9126,N_9751);
nor UO_884 (O_884,N_9263,N_9829);
xnor UO_885 (O_885,N_9658,N_9017);
nor UO_886 (O_886,N_9820,N_9703);
nand UO_887 (O_887,N_9190,N_9966);
and UO_888 (O_888,N_9025,N_9960);
or UO_889 (O_889,N_9055,N_9816);
or UO_890 (O_890,N_9965,N_9784);
xnor UO_891 (O_891,N_9832,N_9827);
nand UO_892 (O_892,N_9060,N_9598);
or UO_893 (O_893,N_9757,N_9367);
nand UO_894 (O_894,N_9653,N_9420);
or UO_895 (O_895,N_9751,N_9872);
xor UO_896 (O_896,N_9957,N_9699);
nand UO_897 (O_897,N_9521,N_9675);
nand UO_898 (O_898,N_9500,N_9524);
or UO_899 (O_899,N_9169,N_9687);
xnor UO_900 (O_900,N_9161,N_9712);
or UO_901 (O_901,N_9602,N_9043);
or UO_902 (O_902,N_9858,N_9337);
xnor UO_903 (O_903,N_9168,N_9953);
nand UO_904 (O_904,N_9837,N_9311);
nand UO_905 (O_905,N_9171,N_9969);
or UO_906 (O_906,N_9786,N_9444);
nand UO_907 (O_907,N_9585,N_9032);
and UO_908 (O_908,N_9611,N_9022);
and UO_909 (O_909,N_9046,N_9665);
and UO_910 (O_910,N_9268,N_9543);
nand UO_911 (O_911,N_9316,N_9037);
nand UO_912 (O_912,N_9188,N_9196);
or UO_913 (O_913,N_9176,N_9896);
or UO_914 (O_914,N_9644,N_9058);
or UO_915 (O_915,N_9874,N_9543);
nor UO_916 (O_916,N_9154,N_9750);
and UO_917 (O_917,N_9872,N_9757);
nand UO_918 (O_918,N_9055,N_9101);
nor UO_919 (O_919,N_9376,N_9484);
nand UO_920 (O_920,N_9679,N_9036);
nand UO_921 (O_921,N_9591,N_9659);
xor UO_922 (O_922,N_9206,N_9281);
or UO_923 (O_923,N_9399,N_9473);
or UO_924 (O_924,N_9968,N_9054);
and UO_925 (O_925,N_9748,N_9952);
and UO_926 (O_926,N_9427,N_9454);
nand UO_927 (O_927,N_9512,N_9626);
nand UO_928 (O_928,N_9012,N_9690);
and UO_929 (O_929,N_9630,N_9243);
or UO_930 (O_930,N_9530,N_9199);
nand UO_931 (O_931,N_9954,N_9735);
xor UO_932 (O_932,N_9614,N_9641);
or UO_933 (O_933,N_9245,N_9198);
xor UO_934 (O_934,N_9249,N_9787);
or UO_935 (O_935,N_9078,N_9212);
and UO_936 (O_936,N_9824,N_9307);
nor UO_937 (O_937,N_9845,N_9628);
nor UO_938 (O_938,N_9943,N_9208);
xnor UO_939 (O_939,N_9212,N_9953);
nor UO_940 (O_940,N_9186,N_9471);
and UO_941 (O_941,N_9997,N_9209);
nand UO_942 (O_942,N_9990,N_9166);
and UO_943 (O_943,N_9812,N_9828);
or UO_944 (O_944,N_9110,N_9747);
or UO_945 (O_945,N_9770,N_9517);
or UO_946 (O_946,N_9906,N_9746);
and UO_947 (O_947,N_9107,N_9103);
nor UO_948 (O_948,N_9270,N_9750);
xor UO_949 (O_949,N_9845,N_9934);
nor UO_950 (O_950,N_9885,N_9830);
and UO_951 (O_951,N_9190,N_9524);
xor UO_952 (O_952,N_9098,N_9777);
or UO_953 (O_953,N_9745,N_9547);
or UO_954 (O_954,N_9799,N_9111);
xor UO_955 (O_955,N_9595,N_9888);
and UO_956 (O_956,N_9120,N_9144);
or UO_957 (O_957,N_9155,N_9078);
or UO_958 (O_958,N_9747,N_9429);
nand UO_959 (O_959,N_9530,N_9205);
nand UO_960 (O_960,N_9007,N_9905);
nand UO_961 (O_961,N_9926,N_9254);
nand UO_962 (O_962,N_9619,N_9419);
xor UO_963 (O_963,N_9288,N_9247);
xnor UO_964 (O_964,N_9637,N_9186);
nand UO_965 (O_965,N_9745,N_9181);
and UO_966 (O_966,N_9586,N_9452);
and UO_967 (O_967,N_9880,N_9500);
nor UO_968 (O_968,N_9922,N_9809);
nand UO_969 (O_969,N_9322,N_9183);
and UO_970 (O_970,N_9436,N_9241);
or UO_971 (O_971,N_9300,N_9306);
xor UO_972 (O_972,N_9879,N_9472);
or UO_973 (O_973,N_9233,N_9100);
and UO_974 (O_974,N_9680,N_9164);
xor UO_975 (O_975,N_9202,N_9384);
nor UO_976 (O_976,N_9564,N_9580);
nor UO_977 (O_977,N_9080,N_9433);
nor UO_978 (O_978,N_9701,N_9991);
xnor UO_979 (O_979,N_9389,N_9494);
and UO_980 (O_980,N_9554,N_9818);
or UO_981 (O_981,N_9799,N_9268);
or UO_982 (O_982,N_9965,N_9688);
nand UO_983 (O_983,N_9557,N_9568);
nand UO_984 (O_984,N_9529,N_9656);
xor UO_985 (O_985,N_9867,N_9139);
nor UO_986 (O_986,N_9661,N_9213);
and UO_987 (O_987,N_9350,N_9400);
nand UO_988 (O_988,N_9934,N_9168);
or UO_989 (O_989,N_9034,N_9687);
nand UO_990 (O_990,N_9648,N_9554);
or UO_991 (O_991,N_9408,N_9403);
and UO_992 (O_992,N_9156,N_9671);
nor UO_993 (O_993,N_9936,N_9094);
or UO_994 (O_994,N_9808,N_9976);
xnor UO_995 (O_995,N_9886,N_9206);
nor UO_996 (O_996,N_9620,N_9581);
and UO_997 (O_997,N_9977,N_9085);
nand UO_998 (O_998,N_9389,N_9917);
nor UO_999 (O_999,N_9707,N_9471);
or UO_1000 (O_1000,N_9527,N_9466);
nor UO_1001 (O_1001,N_9750,N_9955);
nor UO_1002 (O_1002,N_9245,N_9345);
xnor UO_1003 (O_1003,N_9747,N_9943);
xor UO_1004 (O_1004,N_9907,N_9190);
and UO_1005 (O_1005,N_9198,N_9516);
xnor UO_1006 (O_1006,N_9803,N_9226);
nor UO_1007 (O_1007,N_9876,N_9262);
or UO_1008 (O_1008,N_9765,N_9538);
xor UO_1009 (O_1009,N_9323,N_9831);
nor UO_1010 (O_1010,N_9489,N_9471);
and UO_1011 (O_1011,N_9835,N_9542);
and UO_1012 (O_1012,N_9106,N_9935);
nor UO_1013 (O_1013,N_9070,N_9262);
xor UO_1014 (O_1014,N_9378,N_9187);
and UO_1015 (O_1015,N_9644,N_9280);
nand UO_1016 (O_1016,N_9603,N_9860);
nand UO_1017 (O_1017,N_9042,N_9240);
and UO_1018 (O_1018,N_9186,N_9125);
xnor UO_1019 (O_1019,N_9313,N_9521);
or UO_1020 (O_1020,N_9999,N_9744);
xnor UO_1021 (O_1021,N_9744,N_9124);
nor UO_1022 (O_1022,N_9325,N_9291);
and UO_1023 (O_1023,N_9432,N_9640);
xor UO_1024 (O_1024,N_9868,N_9607);
xor UO_1025 (O_1025,N_9693,N_9182);
xnor UO_1026 (O_1026,N_9222,N_9734);
nand UO_1027 (O_1027,N_9100,N_9536);
xor UO_1028 (O_1028,N_9283,N_9063);
or UO_1029 (O_1029,N_9264,N_9663);
or UO_1030 (O_1030,N_9988,N_9741);
xor UO_1031 (O_1031,N_9161,N_9822);
nand UO_1032 (O_1032,N_9201,N_9966);
and UO_1033 (O_1033,N_9039,N_9434);
or UO_1034 (O_1034,N_9755,N_9985);
nor UO_1035 (O_1035,N_9761,N_9201);
nor UO_1036 (O_1036,N_9867,N_9901);
nand UO_1037 (O_1037,N_9723,N_9769);
or UO_1038 (O_1038,N_9447,N_9452);
xor UO_1039 (O_1039,N_9345,N_9664);
nand UO_1040 (O_1040,N_9854,N_9375);
xnor UO_1041 (O_1041,N_9277,N_9850);
xnor UO_1042 (O_1042,N_9787,N_9488);
and UO_1043 (O_1043,N_9508,N_9626);
and UO_1044 (O_1044,N_9738,N_9833);
and UO_1045 (O_1045,N_9304,N_9193);
nand UO_1046 (O_1046,N_9392,N_9248);
xor UO_1047 (O_1047,N_9566,N_9960);
or UO_1048 (O_1048,N_9622,N_9880);
or UO_1049 (O_1049,N_9030,N_9049);
nor UO_1050 (O_1050,N_9835,N_9557);
nor UO_1051 (O_1051,N_9967,N_9819);
xor UO_1052 (O_1052,N_9511,N_9093);
nand UO_1053 (O_1053,N_9892,N_9342);
xor UO_1054 (O_1054,N_9505,N_9151);
nor UO_1055 (O_1055,N_9630,N_9602);
or UO_1056 (O_1056,N_9338,N_9365);
nor UO_1057 (O_1057,N_9414,N_9422);
and UO_1058 (O_1058,N_9470,N_9453);
xor UO_1059 (O_1059,N_9350,N_9886);
nand UO_1060 (O_1060,N_9543,N_9808);
xor UO_1061 (O_1061,N_9158,N_9533);
nor UO_1062 (O_1062,N_9133,N_9940);
and UO_1063 (O_1063,N_9288,N_9612);
nor UO_1064 (O_1064,N_9514,N_9134);
nor UO_1065 (O_1065,N_9884,N_9173);
and UO_1066 (O_1066,N_9682,N_9210);
nand UO_1067 (O_1067,N_9030,N_9723);
nand UO_1068 (O_1068,N_9705,N_9491);
xnor UO_1069 (O_1069,N_9633,N_9044);
nand UO_1070 (O_1070,N_9764,N_9538);
or UO_1071 (O_1071,N_9117,N_9662);
nand UO_1072 (O_1072,N_9960,N_9108);
xor UO_1073 (O_1073,N_9673,N_9551);
nand UO_1074 (O_1074,N_9277,N_9371);
xnor UO_1075 (O_1075,N_9141,N_9075);
xor UO_1076 (O_1076,N_9214,N_9030);
or UO_1077 (O_1077,N_9328,N_9125);
xnor UO_1078 (O_1078,N_9444,N_9917);
and UO_1079 (O_1079,N_9408,N_9880);
nand UO_1080 (O_1080,N_9313,N_9103);
and UO_1081 (O_1081,N_9830,N_9609);
nand UO_1082 (O_1082,N_9751,N_9006);
nand UO_1083 (O_1083,N_9490,N_9343);
and UO_1084 (O_1084,N_9783,N_9261);
xnor UO_1085 (O_1085,N_9672,N_9670);
nor UO_1086 (O_1086,N_9398,N_9903);
nand UO_1087 (O_1087,N_9251,N_9044);
and UO_1088 (O_1088,N_9034,N_9289);
and UO_1089 (O_1089,N_9605,N_9542);
and UO_1090 (O_1090,N_9102,N_9039);
or UO_1091 (O_1091,N_9182,N_9542);
and UO_1092 (O_1092,N_9579,N_9033);
xnor UO_1093 (O_1093,N_9985,N_9966);
nor UO_1094 (O_1094,N_9749,N_9688);
or UO_1095 (O_1095,N_9742,N_9046);
or UO_1096 (O_1096,N_9271,N_9959);
xnor UO_1097 (O_1097,N_9151,N_9120);
nor UO_1098 (O_1098,N_9507,N_9354);
nand UO_1099 (O_1099,N_9883,N_9998);
or UO_1100 (O_1100,N_9926,N_9685);
nor UO_1101 (O_1101,N_9473,N_9263);
nand UO_1102 (O_1102,N_9180,N_9283);
xor UO_1103 (O_1103,N_9784,N_9871);
or UO_1104 (O_1104,N_9735,N_9864);
and UO_1105 (O_1105,N_9997,N_9254);
and UO_1106 (O_1106,N_9311,N_9022);
and UO_1107 (O_1107,N_9724,N_9283);
or UO_1108 (O_1108,N_9241,N_9820);
and UO_1109 (O_1109,N_9963,N_9467);
nor UO_1110 (O_1110,N_9325,N_9258);
xor UO_1111 (O_1111,N_9106,N_9604);
nor UO_1112 (O_1112,N_9214,N_9797);
and UO_1113 (O_1113,N_9522,N_9952);
nand UO_1114 (O_1114,N_9569,N_9700);
and UO_1115 (O_1115,N_9269,N_9564);
xor UO_1116 (O_1116,N_9805,N_9787);
xnor UO_1117 (O_1117,N_9622,N_9968);
xnor UO_1118 (O_1118,N_9304,N_9261);
nand UO_1119 (O_1119,N_9959,N_9545);
nand UO_1120 (O_1120,N_9804,N_9024);
or UO_1121 (O_1121,N_9309,N_9601);
xor UO_1122 (O_1122,N_9913,N_9398);
xor UO_1123 (O_1123,N_9784,N_9832);
and UO_1124 (O_1124,N_9478,N_9649);
and UO_1125 (O_1125,N_9581,N_9500);
xnor UO_1126 (O_1126,N_9871,N_9126);
nand UO_1127 (O_1127,N_9786,N_9867);
nor UO_1128 (O_1128,N_9623,N_9154);
nand UO_1129 (O_1129,N_9544,N_9018);
or UO_1130 (O_1130,N_9884,N_9337);
or UO_1131 (O_1131,N_9335,N_9475);
xor UO_1132 (O_1132,N_9196,N_9571);
and UO_1133 (O_1133,N_9966,N_9487);
nand UO_1134 (O_1134,N_9559,N_9632);
and UO_1135 (O_1135,N_9026,N_9079);
xor UO_1136 (O_1136,N_9598,N_9968);
nand UO_1137 (O_1137,N_9351,N_9863);
and UO_1138 (O_1138,N_9378,N_9697);
nor UO_1139 (O_1139,N_9452,N_9844);
xnor UO_1140 (O_1140,N_9071,N_9779);
nand UO_1141 (O_1141,N_9057,N_9883);
xnor UO_1142 (O_1142,N_9463,N_9869);
or UO_1143 (O_1143,N_9205,N_9916);
and UO_1144 (O_1144,N_9353,N_9309);
nand UO_1145 (O_1145,N_9790,N_9630);
and UO_1146 (O_1146,N_9124,N_9428);
xor UO_1147 (O_1147,N_9434,N_9351);
nor UO_1148 (O_1148,N_9369,N_9707);
and UO_1149 (O_1149,N_9683,N_9704);
nor UO_1150 (O_1150,N_9546,N_9733);
or UO_1151 (O_1151,N_9699,N_9163);
or UO_1152 (O_1152,N_9162,N_9130);
nor UO_1153 (O_1153,N_9477,N_9372);
xor UO_1154 (O_1154,N_9936,N_9767);
nand UO_1155 (O_1155,N_9178,N_9788);
and UO_1156 (O_1156,N_9308,N_9422);
or UO_1157 (O_1157,N_9215,N_9486);
and UO_1158 (O_1158,N_9321,N_9558);
nor UO_1159 (O_1159,N_9491,N_9943);
nand UO_1160 (O_1160,N_9205,N_9290);
nand UO_1161 (O_1161,N_9625,N_9702);
nor UO_1162 (O_1162,N_9738,N_9810);
nor UO_1163 (O_1163,N_9569,N_9897);
or UO_1164 (O_1164,N_9429,N_9109);
nand UO_1165 (O_1165,N_9699,N_9242);
nand UO_1166 (O_1166,N_9700,N_9286);
or UO_1167 (O_1167,N_9336,N_9957);
and UO_1168 (O_1168,N_9779,N_9447);
or UO_1169 (O_1169,N_9571,N_9259);
and UO_1170 (O_1170,N_9917,N_9161);
nand UO_1171 (O_1171,N_9922,N_9271);
xnor UO_1172 (O_1172,N_9764,N_9780);
xor UO_1173 (O_1173,N_9728,N_9628);
nor UO_1174 (O_1174,N_9225,N_9399);
xor UO_1175 (O_1175,N_9828,N_9829);
nand UO_1176 (O_1176,N_9387,N_9781);
or UO_1177 (O_1177,N_9838,N_9163);
nor UO_1178 (O_1178,N_9290,N_9450);
nand UO_1179 (O_1179,N_9841,N_9327);
and UO_1180 (O_1180,N_9526,N_9686);
xor UO_1181 (O_1181,N_9822,N_9747);
nor UO_1182 (O_1182,N_9235,N_9917);
xor UO_1183 (O_1183,N_9658,N_9206);
nor UO_1184 (O_1184,N_9029,N_9227);
or UO_1185 (O_1185,N_9366,N_9569);
or UO_1186 (O_1186,N_9869,N_9157);
nor UO_1187 (O_1187,N_9313,N_9488);
nor UO_1188 (O_1188,N_9973,N_9719);
nor UO_1189 (O_1189,N_9442,N_9819);
nand UO_1190 (O_1190,N_9091,N_9842);
nand UO_1191 (O_1191,N_9497,N_9150);
and UO_1192 (O_1192,N_9990,N_9816);
or UO_1193 (O_1193,N_9449,N_9147);
nor UO_1194 (O_1194,N_9097,N_9398);
and UO_1195 (O_1195,N_9562,N_9711);
nand UO_1196 (O_1196,N_9447,N_9459);
nand UO_1197 (O_1197,N_9774,N_9538);
nand UO_1198 (O_1198,N_9768,N_9502);
xnor UO_1199 (O_1199,N_9831,N_9301);
nor UO_1200 (O_1200,N_9340,N_9332);
nand UO_1201 (O_1201,N_9439,N_9698);
and UO_1202 (O_1202,N_9583,N_9673);
nand UO_1203 (O_1203,N_9288,N_9990);
xnor UO_1204 (O_1204,N_9031,N_9251);
nand UO_1205 (O_1205,N_9256,N_9298);
nor UO_1206 (O_1206,N_9176,N_9729);
or UO_1207 (O_1207,N_9826,N_9100);
and UO_1208 (O_1208,N_9323,N_9832);
nand UO_1209 (O_1209,N_9226,N_9406);
nor UO_1210 (O_1210,N_9728,N_9832);
or UO_1211 (O_1211,N_9384,N_9026);
or UO_1212 (O_1212,N_9664,N_9031);
nor UO_1213 (O_1213,N_9881,N_9950);
nor UO_1214 (O_1214,N_9513,N_9878);
xor UO_1215 (O_1215,N_9752,N_9873);
nand UO_1216 (O_1216,N_9476,N_9797);
nor UO_1217 (O_1217,N_9489,N_9140);
xor UO_1218 (O_1218,N_9527,N_9515);
nand UO_1219 (O_1219,N_9469,N_9430);
xnor UO_1220 (O_1220,N_9659,N_9432);
or UO_1221 (O_1221,N_9376,N_9760);
xnor UO_1222 (O_1222,N_9976,N_9504);
or UO_1223 (O_1223,N_9887,N_9485);
nor UO_1224 (O_1224,N_9634,N_9969);
or UO_1225 (O_1225,N_9673,N_9731);
and UO_1226 (O_1226,N_9463,N_9707);
xnor UO_1227 (O_1227,N_9693,N_9240);
or UO_1228 (O_1228,N_9345,N_9861);
and UO_1229 (O_1229,N_9820,N_9087);
nand UO_1230 (O_1230,N_9227,N_9592);
nor UO_1231 (O_1231,N_9793,N_9394);
nor UO_1232 (O_1232,N_9945,N_9010);
nand UO_1233 (O_1233,N_9603,N_9912);
or UO_1234 (O_1234,N_9436,N_9551);
nor UO_1235 (O_1235,N_9653,N_9949);
or UO_1236 (O_1236,N_9130,N_9140);
nand UO_1237 (O_1237,N_9402,N_9188);
nand UO_1238 (O_1238,N_9637,N_9006);
nand UO_1239 (O_1239,N_9549,N_9002);
and UO_1240 (O_1240,N_9343,N_9433);
or UO_1241 (O_1241,N_9174,N_9774);
xor UO_1242 (O_1242,N_9822,N_9048);
nor UO_1243 (O_1243,N_9958,N_9262);
xor UO_1244 (O_1244,N_9812,N_9440);
nor UO_1245 (O_1245,N_9155,N_9992);
xnor UO_1246 (O_1246,N_9121,N_9015);
or UO_1247 (O_1247,N_9132,N_9335);
xor UO_1248 (O_1248,N_9023,N_9236);
and UO_1249 (O_1249,N_9402,N_9260);
nor UO_1250 (O_1250,N_9844,N_9573);
xnor UO_1251 (O_1251,N_9257,N_9117);
and UO_1252 (O_1252,N_9817,N_9070);
and UO_1253 (O_1253,N_9285,N_9276);
or UO_1254 (O_1254,N_9236,N_9450);
and UO_1255 (O_1255,N_9522,N_9148);
nor UO_1256 (O_1256,N_9061,N_9305);
xnor UO_1257 (O_1257,N_9428,N_9366);
or UO_1258 (O_1258,N_9807,N_9639);
xor UO_1259 (O_1259,N_9125,N_9253);
xor UO_1260 (O_1260,N_9588,N_9501);
and UO_1261 (O_1261,N_9430,N_9427);
xor UO_1262 (O_1262,N_9663,N_9432);
nor UO_1263 (O_1263,N_9846,N_9794);
or UO_1264 (O_1264,N_9489,N_9749);
xnor UO_1265 (O_1265,N_9766,N_9680);
xor UO_1266 (O_1266,N_9481,N_9281);
xor UO_1267 (O_1267,N_9635,N_9376);
nand UO_1268 (O_1268,N_9742,N_9545);
and UO_1269 (O_1269,N_9844,N_9023);
nor UO_1270 (O_1270,N_9500,N_9609);
nor UO_1271 (O_1271,N_9483,N_9389);
nor UO_1272 (O_1272,N_9434,N_9554);
and UO_1273 (O_1273,N_9759,N_9855);
or UO_1274 (O_1274,N_9763,N_9013);
nand UO_1275 (O_1275,N_9395,N_9836);
xnor UO_1276 (O_1276,N_9783,N_9917);
xor UO_1277 (O_1277,N_9835,N_9915);
nand UO_1278 (O_1278,N_9774,N_9747);
and UO_1279 (O_1279,N_9119,N_9002);
or UO_1280 (O_1280,N_9775,N_9028);
or UO_1281 (O_1281,N_9652,N_9336);
xnor UO_1282 (O_1282,N_9899,N_9418);
or UO_1283 (O_1283,N_9777,N_9779);
nor UO_1284 (O_1284,N_9971,N_9503);
nor UO_1285 (O_1285,N_9275,N_9484);
xnor UO_1286 (O_1286,N_9860,N_9166);
xnor UO_1287 (O_1287,N_9472,N_9744);
nor UO_1288 (O_1288,N_9804,N_9841);
xnor UO_1289 (O_1289,N_9631,N_9427);
or UO_1290 (O_1290,N_9603,N_9511);
xnor UO_1291 (O_1291,N_9376,N_9099);
nor UO_1292 (O_1292,N_9165,N_9912);
or UO_1293 (O_1293,N_9554,N_9748);
nand UO_1294 (O_1294,N_9203,N_9204);
and UO_1295 (O_1295,N_9304,N_9691);
or UO_1296 (O_1296,N_9412,N_9333);
or UO_1297 (O_1297,N_9121,N_9291);
and UO_1298 (O_1298,N_9702,N_9255);
nor UO_1299 (O_1299,N_9996,N_9097);
or UO_1300 (O_1300,N_9498,N_9958);
xor UO_1301 (O_1301,N_9691,N_9674);
nor UO_1302 (O_1302,N_9664,N_9940);
and UO_1303 (O_1303,N_9167,N_9121);
nor UO_1304 (O_1304,N_9936,N_9598);
nand UO_1305 (O_1305,N_9295,N_9904);
nor UO_1306 (O_1306,N_9559,N_9929);
nand UO_1307 (O_1307,N_9620,N_9489);
nand UO_1308 (O_1308,N_9150,N_9748);
and UO_1309 (O_1309,N_9699,N_9597);
xor UO_1310 (O_1310,N_9905,N_9151);
and UO_1311 (O_1311,N_9391,N_9221);
and UO_1312 (O_1312,N_9940,N_9378);
xnor UO_1313 (O_1313,N_9611,N_9679);
xnor UO_1314 (O_1314,N_9774,N_9350);
nor UO_1315 (O_1315,N_9759,N_9871);
nand UO_1316 (O_1316,N_9475,N_9374);
nor UO_1317 (O_1317,N_9239,N_9779);
nor UO_1318 (O_1318,N_9401,N_9515);
nor UO_1319 (O_1319,N_9559,N_9973);
nor UO_1320 (O_1320,N_9203,N_9216);
nor UO_1321 (O_1321,N_9617,N_9929);
and UO_1322 (O_1322,N_9004,N_9976);
xnor UO_1323 (O_1323,N_9204,N_9628);
nor UO_1324 (O_1324,N_9872,N_9761);
nor UO_1325 (O_1325,N_9112,N_9122);
or UO_1326 (O_1326,N_9871,N_9193);
nand UO_1327 (O_1327,N_9722,N_9877);
or UO_1328 (O_1328,N_9080,N_9001);
nor UO_1329 (O_1329,N_9151,N_9927);
xnor UO_1330 (O_1330,N_9901,N_9188);
nand UO_1331 (O_1331,N_9883,N_9678);
nor UO_1332 (O_1332,N_9064,N_9846);
or UO_1333 (O_1333,N_9722,N_9307);
or UO_1334 (O_1334,N_9194,N_9819);
and UO_1335 (O_1335,N_9445,N_9415);
nor UO_1336 (O_1336,N_9832,N_9754);
nor UO_1337 (O_1337,N_9509,N_9695);
and UO_1338 (O_1338,N_9400,N_9627);
nand UO_1339 (O_1339,N_9863,N_9430);
nor UO_1340 (O_1340,N_9236,N_9871);
and UO_1341 (O_1341,N_9340,N_9764);
or UO_1342 (O_1342,N_9219,N_9898);
or UO_1343 (O_1343,N_9550,N_9204);
nand UO_1344 (O_1344,N_9757,N_9960);
nor UO_1345 (O_1345,N_9075,N_9960);
nand UO_1346 (O_1346,N_9669,N_9558);
and UO_1347 (O_1347,N_9824,N_9513);
xor UO_1348 (O_1348,N_9562,N_9796);
xnor UO_1349 (O_1349,N_9695,N_9537);
nand UO_1350 (O_1350,N_9902,N_9616);
nor UO_1351 (O_1351,N_9599,N_9277);
nand UO_1352 (O_1352,N_9814,N_9547);
xnor UO_1353 (O_1353,N_9434,N_9664);
xor UO_1354 (O_1354,N_9623,N_9011);
or UO_1355 (O_1355,N_9097,N_9019);
nand UO_1356 (O_1356,N_9216,N_9811);
and UO_1357 (O_1357,N_9614,N_9424);
nand UO_1358 (O_1358,N_9225,N_9060);
xnor UO_1359 (O_1359,N_9736,N_9808);
xnor UO_1360 (O_1360,N_9564,N_9216);
nand UO_1361 (O_1361,N_9326,N_9928);
nand UO_1362 (O_1362,N_9221,N_9993);
xnor UO_1363 (O_1363,N_9355,N_9072);
or UO_1364 (O_1364,N_9571,N_9208);
and UO_1365 (O_1365,N_9489,N_9448);
xor UO_1366 (O_1366,N_9804,N_9110);
and UO_1367 (O_1367,N_9805,N_9358);
and UO_1368 (O_1368,N_9028,N_9200);
nor UO_1369 (O_1369,N_9350,N_9729);
or UO_1370 (O_1370,N_9283,N_9051);
xnor UO_1371 (O_1371,N_9472,N_9662);
and UO_1372 (O_1372,N_9993,N_9595);
and UO_1373 (O_1373,N_9272,N_9873);
and UO_1374 (O_1374,N_9768,N_9381);
xor UO_1375 (O_1375,N_9754,N_9606);
nand UO_1376 (O_1376,N_9735,N_9692);
nand UO_1377 (O_1377,N_9085,N_9694);
and UO_1378 (O_1378,N_9157,N_9837);
xor UO_1379 (O_1379,N_9720,N_9478);
and UO_1380 (O_1380,N_9162,N_9571);
or UO_1381 (O_1381,N_9568,N_9566);
or UO_1382 (O_1382,N_9437,N_9220);
or UO_1383 (O_1383,N_9449,N_9718);
and UO_1384 (O_1384,N_9662,N_9764);
xnor UO_1385 (O_1385,N_9396,N_9601);
nor UO_1386 (O_1386,N_9185,N_9250);
or UO_1387 (O_1387,N_9802,N_9264);
nand UO_1388 (O_1388,N_9542,N_9016);
nand UO_1389 (O_1389,N_9685,N_9408);
nand UO_1390 (O_1390,N_9962,N_9589);
nor UO_1391 (O_1391,N_9359,N_9194);
and UO_1392 (O_1392,N_9894,N_9923);
nand UO_1393 (O_1393,N_9725,N_9092);
nand UO_1394 (O_1394,N_9878,N_9620);
xnor UO_1395 (O_1395,N_9538,N_9653);
xnor UO_1396 (O_1396,N_9430,N_9225);
nand UO_1397 (O_1397,N_9410,N_9115);
nor UO_1398 (O_1398,N_9265,N_9398);
nand UO_1399 (O_1399,N_9837,N_9927);
or UO_1400 (O_1400,N_9117,N_9417);
or UO_1401 (O_1401,N_9198,N_9363);
and UO_1402 (O_1402,N_9440,N_9551);
xor UO_1403 (O_1403,N_9952,N_9786);
and UO_1404 (O_1404,N_9418,N_9820);
xnor UO_1405 (O_1405,N_9846,N_9160);
nor UO_1406 (O_1406,N_9716,N_9879);
nor UO_1407 (O_1407,N_9413,N_9788);
or UO_1408 (O_1408,N_9657,N_9004);
or UO_1409 (O_1409,N_9313,N_9947);
and UO_1410 (O_1410,N_9145,N_9769);
nor UO_1411 (O_1411,N_9799,N_9897);
xor UO_1412 (O_1412,N_9571,N_9598);
or UO_1413 (O_1413,N_9598,N_9860);
nand UO_1414 (O_1414,N_9683,N_9984);
nand UO_1415 (O_1415,N_9960,N_9494);
or UO_1416 (O_1416,N_9211,N_9103);
or UO_1417 (O_1417,N_9823,N_9148);
or UO_1418 (O_1418,N_9383,N_9854);
or UO_1419 (O_1419,N_9422,N_9000);
xnor UO_1420 (O_1420,N_9698,N_9899);
or UO_1421 (O_1421,N_9052,N_9504);
and UO_1422 (O_1422,N_9827,N_9985);
xnor UO_1423 (O_1423,N_9472,N_9893);
xnor UO_1424 (O_1424,N_9829,N_9086);
xor UO_1425 (O_1425,N_9324,N_9361);
xnor UO_1426 (O_1426,N_9159,N_9282);
xnor UO_1427 (O_1427,N_9940,N_9116);
and UO_1428 (O_1428,N_9881,N_9751);
and UO_1429 (O_1429,N_9574,N_9203);
nand UO_1430 (O_1430,N_9630,N_9431);
and UO_1431 (O_1431,N_9784,N_9226);
or UO_1432 (O_1432,N_9423,N_9976);
xnor UO_1433 (O_1433,N_9109,N_9008);
nor UO_1434 (O_1434,N_9143,N_9535);
nand UO_1435 (O_1435,N_9232,N_9845);
xor UO_1436 (O_1436,N_9748,N_9829);
xor UO_1437 (O_1437,N_9555,N_9873);
and UO_1438 (O_1438,N_9668,N_9366);
nor UO_1439 (O_1439,N_9589,N_9478);
nand UO_1440 (O_1440,N_9004,N_9014);
xor UO_1441 (O_1441,N_9588,N_9762);
or UO_1442 (O_1442,N_9131,N_9200);
nor UO_1443 (O_1443,N_9176,N_9278);
and UO_1444 (O_1444,N_9023,N_9103);
or UO_1445 (O_1445,N_9226,N_9700);
nand UO_1446 (O_1446,N_9521,N_9084);
or UO_1447 (O_1447,N_9696,N_9571);
nand UO_1448 (O_1448,N_9582,N_9438);
nor UO_1449 (O_1449,N_9394,N_9501);
and UO_1450 (O_1450,N_9525,N_9489);
or UO_1451 (O_1451,N_9468,N_9004);
xnor UO_1452 (O_1452,N_9458,N_9642);
nor UO_1453 (O_1453,N_9603,N_9568);
nand UO_1454 (O_1454,N_9900,N_9236);
nor UO_1455 (O_1455,N_9492,N_9726);
or UO_1456 (O_1456,N_9356,N_9420);
nand UO_1457 (O_1457,N_9997,N_9366);
nor UO_1458 (O_1458,N_9693,N_9356);
and UO_1459 (O_1459,N_9507,N_9413);
and UO_1460 (O_1460,N_9637,N_9350);
xor UO_1461 (O_1461,N_9785,N_9368);
nor UO_1462 (O_1462,N_9892,N_9949);
xor UO_1463 (O_1463,N_9823,N_9845);
and UO_1464 (O_1464,N_9959,N_9054);
xor UO_1465 (O_1465,N_9773,N_9816);
xor UO_1466 (O_1466,N_9883,N_9521);
xor UO_1467 (O_1467,N_9535,N_9175);
nor UO_1468 (O_1468,N_9671,N_9334);
xnor UO_1469 (O_1469,N_9144,N_9217);
or UO_1470 (O_1470,N_9724,N_9281);
nand UO_1471 (O_1471,N_9525,N_9571);
or UO_1472 (O_1472,N_9225,N_9369);
or UO_1473 (O_1473,N_9754,N_9331);
and UO_1474 (O_1474,N_9434,N_9675);
and UO_1475 (O_1475,N_9737,N_9463);
nand UO_1476 (O_1476,N_9825,N_9965);
nand UO_1477 (O_1477,N_9186,N_9429);
xor UO_1478 (O_1478,N_9678,N_9847);
xnor UO_1479 (O_1479,N_9188,N_9265);
and UO_1480 (O_1480,N_9506,N_9606);
nand UO_1481 (O_1481,N_9956,N_9221);
nand UO_1482 (O_1482,N_9041,N_9844);
nand UO_1483 (O_1483,N_9087,N_9877);
nor UO_1484 (O_1484,N_9371,N_9998);
nand UO_1485 (O_1485,N_9611,N_9016);
or UO_1486 (O_1486,N_9892,N_9465);
and UO_1487 (O_1487,N_9448,N_9827);
nor UO_1488 (O_1488,N_9304,N_9280);
and UO_1489 (O_1489,N_9152,N_9589);
nand UO_1490 (O_1490,N_9766,N_9594);
and UO_1491 (O_1491,N_9405,N_9606);
or UO_1492 (O_1492,N_9640,N_9253);
or UO_1493 (O_1493,N_9639,N_9533);
or UO_1494 (O_1494,N_9915,N_9645);
or UO_1495 (O_1495,N_9248,N_9533);
or UO_1496 (O_1496,N_9781,N_9989);
nand UO_1497 (O_1497,N_9423,N_9882);
nor UO_1498 (O_1498,N_9314,N_9879);
nor UO_1499 (O_1499,N_9667,N_9223);
endmodule