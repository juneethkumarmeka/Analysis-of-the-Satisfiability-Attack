module basic_2500_25000_3000_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_648,In_1784);
xor U1 (N_1,In_1783,In_543);
or U2 (N_2,In_1411,In_1785);
nand U3 (N_3,In_1687,In_2448);
nand U4 (N_4,In_1600,In_1035);
and U5 (N_5,In_2048,In_1336);
and U6 (N_6,In_1234,In_318);
and U7 (N_7,In_1678,In_1960);
nor U8 (N_8,In_97,In_148);
and U9 (N_9,In_1535,In_1114);
xnor U10 (N_10,In_904,In_1185);
xnor U11 (N_11,In_1342,In_2489);
xor U12 (N_12,In_253,In_176);
xnor U13 (N_13,In_1400,In_1349);
and U14 (N_14,In_1584,In_175);
or U15 (N_15,In_2,In_1103);
or U16 (N_16,In_2292,In_2400);
xnor U17 (N_17,In_290,In_902);
nor U18 (N_18,In_735,In_1454);
or U19 (N_19,In_716,In_820);
and U20 (N_20,In_1686,In_1746);
nand U21 (N_21,In_146,In_1860);
nor U22 (N_22,In_1504,In_27);
or U23 (N_23,In_1436,In_50);
or U24 (N_24,In_342,In_2162);
or U25 (N_25,In_2161,In_600);
nor U26 (N_26,In_534,In_1953);
or U27 (N_27,In_495,In_2117);
xor U28 (N_28,In_951,In_1346);
nand U29 (N_29,In_1542,In_0);
and U30 (N_30,In_2398,In_2253);
xor U31 (N_31,In_911,In_255);
and U32 (N_32,In_1474,In_1972);
or U33 (N_33,In_1494,In_1961);
and U34 (N_34,In_326,In_2209);
or U35 (N_35,In_237,In_168);
or U36 (N_36,In_354,In_2471);
or U37 (N_37,In_1318,In_1227);
or U38 (N_38,In_1423,In_394);
and U39 (N_39,In_461,In_1782);
xnor U40 (N_40,In_1105,In_2174);
or U41 (N_41,In_330,In_179);
nor U42 (N_42,In_378,In_494);
nand U43 (N_43,In_2127,In_2077);
and U44 (N_44,In_340,In_935);
nor U45 (N_45,In_1196,In_1232);
xnor U46 (N_46,In_1138,In_2222);
nor U47 (N_47,In_1485,In_2337);
nand U48 (N_48,In_2334,In_42);
or U49 (N_49,In_65,In_1191);
and U50 (N_50,In_2439,In_421);
and U51 (N_51,In_391,In_630);
and U52 (N_52,In_214,In_196);
and U53 (N_53,In_1226,In_476);
nor U54 (N_54,In_818,In_1266);
xnor U55 (N_55,In_2455,In_35);
nor U56 (N_56,In_635,In_1689);
nor U57 (N_57,In_1399,In_287);
and U58 (N_58,In_1479,In_1999);
nand U59 (N_59,In_762,In_445);
nand U60 (N_60,In_103,In_22);
nor U61 (N_61,In_186,In_1541);
nor U62 (N_62,In_2086,In_440);
nor U63 (N_63,In_2373,In_450);
or U64 (N_64,In_142,In_1493);
xor U65 (N_65,In_104,In_769);
and U66 (N_66,In_869,In_133);
and U67 (N_67,In_1666,In_344);
or U68 (N_68,In_2223,In_966);
nand U69 (N_69,In_134,In_687);
nor U70 (N_70,In_560,In_953);
and U71 (N_71,In_386,In_541);
or U72 (N_72,In_1507,In_1367);
nor U73 (N_73,In_2025,In_2258);
nand U74 (N_74,In_279,In_1895);
and U75 (N_75,In_1768,In_1052);
xor U76 (N_76,In_1863,In_1016);
or U77 (N_77,In_2112,In_137);
nand U78 (N_78,In_2148,In_162);
or U79 (N_79,In_2172,In_699);
and U80 (N_80,In_791,In_976);
nand U81 (N_81,In_598,In_1045);
xor U82 (N_82,In_2121,In_1492);
nand U83 (N_83,In_45,In_1024);
or U84 (N_84,In_633,In_167);
nor U85 (N_85,In_1853,In_264);
nand U86 (N_86,In_2377,In_1833);
or U87 (N_87,In_1491,In_434);
or U88 (N_88,In_428,In_901);
nand U89 (N_89,In_2485,In_513);
or U90 (N_90,In_907,In_2040);
or U91 (N_91,In_449,In_2273);
nand U92 (N_92,In_1630,In_602);
nor U93 (N_93,In_1156,In_2453);
xor U94 (N_94,In_1903,In_20);
nand U95 (N_95,In_2323,In_945);
or U96 (N_96,In_2220,In_2217);
xor U97 (N_97,In_1550,In_388);
nand U98 (N_98,In_2319,In_1617);
and U99 (N_99,In_319,In_2108);
xnor U100 (N_100,In_1740,In_1308);
and U101 (N_101,In_207,In_788);
and U102 (N_102,In_532,In_1446);
or U103 (N_103,In_2457,In_1183);
nand U104 (N_104,In_2451,In_78);
xnor U105 (N_105,In_1119,In_2277);
nor U106 (N_106,In_718,In_1332);
nand U107 (N_107,In_928,In_644);
xor U108 (N_108,In_1095,In_229);
and U109 (N_109,In_2213,In_570);
nor U110 (N_110,In_1927,In_462);
nand U111 (N_111,In_1090,In_2085);
and U112 (N_112,In_180,In_2327);
or U113 (N_113,In_1819,In_91);
or U114 (N_114,In_135,In_372);
xnor U115 (N_115,In_1324,In_2286);
nand U116 (N_116,In_1847,In_830);
and U117 (N_117,In_1606,In_2308);
xnor U118 (N_118,In_203,In_161);
and U119 (N_119,In_31,In_2016);
nand U120 (N_120,In_566,In_550);
or U121 (N_121,In_2297,In_1518);
nor U122 (N_122,In_251,In_1078);
and U123 (N_123,In_1533,In_1592);
or U124 (N_124,In_1247,In_1300);
or U125 (N_125,In_812,In_777);
xnor U126 (N_126,In_136,In_2134);
and U127 (N_127,In_2126,In_1495);
xnor U128 (N_128,In_1030,In_359);
or U129 (N_129,In_517,In_46);
nand U130 (N_130,In_1951,In_2461);
and U131 (N_131,In_1874,In_683);
and U132 (N_132,In_86,In_2272);
and U133 (N_133,In_384,In_1403);
nand U134 (N_134,In_554,In_518);
and U135 (N_135,In_1309,In_1167);
nand U136 (N_136,In_800,In_525);
and U137 (N_137,In_1829,In_2071);
xor U138 (N_138,In_1994,In_1458);
or U139 (N_139,In_1339,In_1820);
and U140 (N_140,In_831,In_2135);
nor U141 (N_141,In_888,In_1886);
xnor U142 (N_142,In_511,In_2477);
or U143 (N_143,In_341,In_1422);
and U144 (N_144,In_510,In_2046);
or U145 (N_145,In_2452,In_1778);
xor U146 (N_146,In_1735,In_2190);
nor U147 (N_147,In_744,In_987);
xnor U148 (N_148,In_1418,In_1622);
nand U149 (N_149,In_1073,In_159);
nand U150 (N_150,In_2459,In_1276);
or U151 (N_151,In_1758,In_677);
nand U152 (N_152,In_194,In_631);
and U153 (N_153,In_1798,In_2359);
nand U154 (N_154,In_1851,In_924);
and U155 (N_155,In_2371,In_2491);
xnor U156 (N_156,In_256,In_530);
nand U157 (N_157,In_1182,In_1110);
nor U158 (N_158,In_2120,In_559);
and U159 (N_159,In_1553,In_1770);
xor U160 (N_160,In_1958,In_746);
and U161 (N_161,In_929,In_742);
nand U162 (N_162,In_34,In_2275);
and U163 (N_163,In_1811,In_2106);
nor U164 (N_164,In_1051,In_1814);
xor U165 (N_165,In_1831,In_268);
nand U166 (N_166,In_1169,In_1189);
nand U167 (N_167,In_569,In_958);
nor U168 (N_168,In_1369,In_1616);
and U169 (N_169,In_1857,In_1765);
xnor U170 (N_170,In_1982,In_2429);
and U171 (N_171,In_944,In_2151);
and U172 (N_172,In_1433,In_451);
or U173 (N_173,In_927,In_1229);
nand U174 (N_174,In_1161,In_866);
and U175 (N_175,In_975,In_850);
nor U176 (N_176,In_1194,In_387);
or U177 (N_177,In_2476,In_620);
xnor U178 (N_178,In_1567,In_2235);
nand U179 (N_179,In_2283,In_1228);
nand U180 (N_180,In_1426,In_1712);
nand U181 (N_181,In_258,In_1685);
xnor U182 (N_182,In_1887,In_712);
nand U183 (N_183,In_2437,In_509);
and U184 (N_184,In_422,In_1801);
and U185 (N_185,In_1395,In_1179);
nand U186 (N_186,In_1866,In_2160);
and U187 (N_187,In_2414,In_1481);
and U188 (N_188,In_2008,In_343);
and U189 (N_189,In_2043,In_516);
nor U190 (N_190,In_1421,In_1467);
nor U191 (N_191,In_969,In_899);
and U192 (N_192,In_1896,In_1291);
nor U193 (N_193,In_1304,In_1737);
nand U194 (N_194,In_1050,In_2236);
nand U195 (N_195,In_874,In_1718);
or U196 (N_196,In_1576,In_1926);
nand U197 (N_197,In_2279,In_708);
xnor U198 (N_198,In_299,In_2208);
nand U199 (N_199,In_2200,In_26);
xnor U200 (N_200,In_2203,In_601);
or U201 (N_201,In_720,In_1713);
nand U202 (N_202,In_1466,In_2354);
and U203 (N_203,In_700,In_1835);
or U204 (N_204,In_1190,In_363);
or U205 (N_205,In_1027,In_1230);
nand U206 (N_206,In_860,In_1);
nand U207 (N_207,In_412,In_123);
nor U208 (N_208,In_2364,In_2247);
xor U209 (N_209,In_1094,In_2311);
xnor U210 (N_210,In_627,In_7);
or U211 (N_211,In_932,In_819);
and U212 (N_212,In_723,In_333);
xnor U213 (N_213,In_2079,In_2341);
xor U214 (N_214,In_1599,In_727);
xor U215 (N_215,In_1539,In_1744);
nor U216 (N_216,In_2144,In_713);
nand U217 (N_217,In_1377,In_2034);
xor U218 (N_218,In_1343,In_1430);
nand U219 (N_219,In_1813,In_2069);
nand U220 (N_220,In_871,In_521);
nor U221 (N_221,In_2047,In_182);
nor U222 (N_222,In_2038,In_918);
nand U223 (N_223,In_2321,In_471);
xnor U224 (N_224,In_2231,In_2234);
or U225 (N_225,In_1021,In_1872);
xnor U226 (N_226,In_2122,In_124);
nor U227 (N_227,In_2284,In_2210);
xor U228 (N_228,In_581,In_1112);
nand U229 (N_229,In_1294,In_1483);
nor U230 (N_230,In_2405,In_841);
nor U231 (N_231,In_2224,In_415);
nor U232 (N_232,In_1379,In_1134);
xor U233 (N_233,In_1205,In_1011);
and U234 (N_234,In_1405,In_1463);
xor U235 (N_235,In_349,In_325);
and U236 (N_236,In_1544,In_2076);
or U237 (N_237,In_2496,In_590);
nand U238 (N_238,In_284,In_961);
nor U239 (N_239,In_155,In_1626);
nand U240 (N_240,In_611,In_671);
nand U241 (N_241,In_417,In_441);
nor U242 (N_242,In_2153,In_347);
nand U243 (N_243,In_2003,In_593);
or U244 (N_244,In_2299,In_295);
nor U245 (N_245,In_1524,In_2374);
and U246 (N_246,In_1509,In_1143);
nand U247 (N_247,In_1407,In_315);
nand U248 (N_248,In_992,In_1231);
nor U249 (N_249,In_974,In_1575);
or U250 (N_250,In_2061,In_529);
xnor U251 (N_251,In_1873,In_1184);
xor U252 (N_252,In_565,In_1916);
nor U253 (N_253,In_1545,In_1233);
or U254 (N_254,In_1681,In_1918);
nor U255 (N_255,In_174,In_1139);
and U256 (N_256,In_858,In_1036);
nor U257 (N_257,In_353,In_235);
nand U258 (N_258,In_2152,In_1669);
and U259 (N_259,In_770,In_1163);
and U260 (N_260,In_67,In_416);
nand U261 (N_261,In_887,In_1675);
nor U262 (N_262,In_1260,In_2394);
or U263 (N_263,In_2406,In_896);
or U264 (N_264,In_2417,In_1155);
or U265 (N_265,In_1906,In_1448);
xor U266 (N_266,In_1450,In_982);
or U267 (N_267,In_1314,In_1146);
nand U268 (N_268,In_1838,In_1453);
and U269 (N_269,In_626,In_1564);
or U270 (N_270,In_970,In_783);
nor U271 (N_271,In_863,In_2198);
and U272 (N_272,In_1128,In_1827);
or U273 (N_273,In_1353,In_539);
nor U274 (N_274,In_583,In_813);
xnor U275 (N_275,In_307,In_1644);
nor U276 (N_276,In_1216,In_51);
and U277 (N_277,In_1655,In_681);
nand U278 (N_278,In_2011,In_1312);
nor U279 (N_279,In_1743,In_609);
nor U280 (N_280,In_1284,In_2166);
and U281 (N_281,In_1736,In_154);
or U282 (N_282,In_1614,In_526);
nor U283 (N_283,In_1009,In_389);
or U284 (N_284,In_2212,In_2178);
nor U285 (N_285,In_1836,In_1135);
nand U286 (N_286,In_212,In_1749);
or U287 (N_287,In_1325,In_675);
or U288 (N_288,In_955,In_789);
or U289 (N_289,In_2466,In_2487);
xor U290 (N_290,In_2099,In_938);
or U291 (N_291,In_195,In_247);
or U292 (N_292,In_2328,In_2310);
nand U293 (N_293,In_2395,In_678);
nand U294 (N_294,In_220,In_647);
xnor U295 (N_295,In_972,In_694);
nor U296 (N_296,In_1580,In_2221);
nor U297 (N_297,In_243,In_38);
nand U298 (N_298,In_2369,In_2347);
nand U299 (N_299,In_456,In_37);
and U300 (N_300,In_170,In_1307);
and U301 (N_301,In_192,In_1549);
xor U302 (N_302,In_1883,In_538);
xnor U303 (N_303,In_1417,In_1597);
xnor U304 (N_304,In_2019,In_2020);
and U305 (N_305,In_2419,In_1047);
nand U306 (N_306,In_385,In_773);
nor U307 (N_307,In_2484,In_2475);
and U308 (N_308,In_990,In_920);
nor U309 (N_309,In_1438,In_952);
nor U310 (N_310,In_2449,In_1933);
or U311 (N_311,In_2467,In_301);
nand U312 (N_312,In_1511,In_1610);
nor U313 (N_313,In_2396,In_407);
and U314 (N_314,In_823,In_439);
nor U315 (N_315,In_1396,In_891);
or U316 (N_316,In_573,In_715);
xor U317 (N_317,In_1968,In_352);
or U318 (N_318,In_2165,In_1975);
nand U319 (N_319,In_743,In_1442);
nor U320 (N_320,In_1757,In_2114);
or U321 (N_321,In_1480,In_1728);
or U322 (N_322,In_14,In_1899);
xnor U323 (N_323,In_100,In_2344);
xor U324 (N_324,In_1251,In_2101);
xor U325 (N_325,In_956,In_1322);
xnor U326 (N_326,In_2097,In_2133);
and U327 (N_327,In_2193,In_2167);
nor U328 (N_328,In_759,In_122);
and U329 (N_329,In_2123,In_1427);
nor U330 (N_330,In_758,In_150);
xor U331 (N_331,In_1796,In_1026);
and U332 (N_332,In_1250,In_2256);
xnor U333 (N_333,In_676,In_651);
nor U334 (N_334,In_971,In_87);
nor U335 (N_335,In_1013,In_1374);
nor U336 (N_336,In_588,In_1520);
and U337 (N_337,In_906,In_184);
and U338 (N_338,In_2062,In_807);
and U339 (N_339,In_1805,In_41);
and U340 (N_340,In_483,In_2052);
nor U341 (N_341,In_1213,In_1240);
and U342 (N_342,In_74,In_1653);
xnor U343 (N_343,In_586,In_963);
or U344 (N_344,In_2239,In_838);
or U345 (N_345,In_1077,In_1419);
nand U346 (N_346,In_1745,In_291);
nor U347 (N_347,In_1780,In_1629);
nand U348 (N_348,In_1921,In_2156);
or U349 (N_349,In_499,In_1131);
and U350 (N_350,In_851,In_166);
and U351 (N_351,In_147,In_2353);
or U352 (N_352,In_81,In_981);
nor U353 (N_353,In_2228,In_616);
xor U354 (N_354,In_3,In_1341);
nand U355 (N_355,In_1772,In_1748);
nor U356 (N_356,In_139,In_473);
xnor U357 (N_357,In_1262,In_1787);
or U358 (N_358,In_2237,In_2257);
or U359 (N_359,In_1905,In_2051);
and U360 (N_360,In_1708,In_1282);
or U361 (N_361,In_2331,In_1969);
nor U362 (N_362,In_1996,In_10);
nand U363 (N_363,In_726,In_1941);
nand U364 (N_364,In_1547,In_2492);
nand U365 (N_365,In_1086,In_1651);
or U366 (N_366,In_1362,In_2107);
nor U367 (N_367,In_2074,In_316);
xor U368 (N_368,In_1605,In_1832);
xor U369 (N_369,In_1596,In_2497);
or U370 (N_370,In_331,In_221);
xor U371 (N_371,In_1673,In_701);
and U372 (N_372,In_364,In_1537);
nand U373 (N_373,In_1197,In_77);
nand U374 (N_374,In_2180,In_115);
and U375 (N_375,In_2088,In_1007);
nor U376 (N_376,In_520,In_185);
nor U377 (N_377,In_1409,In_1038);
and U378 (N_378,In_210,In_1044);
xor U379 (N_379,In_374,In_898);
and U380 (N_380,In_259,In_1674);
nor U381 (N_381,In_1789,In_397);
or U382 (N_382,In_2057,In_877);
and U383 (N_383,In_1102,In_2171);
xnor U384 (N_384,In_829,In_774);
or U385 (N_385,In_2169,In_1410);
or U386 (N_386,In_1634,In_444);
xor U387 (N_387,In_979,In_1841);
and U388 (N_388,In_504,In_469);
or U389 (N_389,In_1637,In_1145);
nand U390 (N_390,In_2176,In_2488);
xor U391 (N_391,In_1350,In_1729);
and U392 (N_392,In_747,In_1812);
nor U393 (N_393,In_1107,In_1366);
nor U394 (N_394,In_1486,In_890);
and U395 (N_395,In_1852,In_266);
xnor U396 (N_396,In_1048,In_413);
nor U397 (N_397,In_578,In_1122);
or U398 (N_398,In_2211,In_382);
nor U399 (N_399,In_973,In_490);
xor U400 (N_400,In_2118,In_276);
nor U401 (N_401,In_492,In_197);
nor U402 (N_402,In_1693,In_1619);
nand U403 (N_403,In_1572,In_47);
nand U404 (N_404,In_481,In_643);
or U405 (N_405,In_1313,In_1710);
nor U406 (N_406,In_2241,In_1907);
nand U407 (N_407,In_505,In_2454);
nor U408 (N_408,In_1053,In_1130);
or U409 (N_409,In_1791,In_1816);
nor U410 (N_410,In_114,In_872);
nor U411 (N_411,In_1581,In_1159);
nor U412 (N_412,In_628,In_2370);
nor U413 (N_413,In_2482,In_2443);
or U414 (N_414,In_638,In_1397);
or U415 (N_415,In_1691,In_1255);
and U416 (N_416,In_1297,In_2407);
xnor U417 (N_417,In_1747,In_1447);
xnor U418 (N_418,In_1931,In_33);
nand U419 (N_419,In_423,In_2262);
and U420 (N_420,In_668,In_926);
or U421 (N_421,In_1611,In_2330);
and U422 (N_422,In_817,In_1557);
or U423 (N_423,In_908,In_612);
nand U424 (N_424,In_1010,In_905);
nor U425 (N_425,In_1187,In_191);
nor U426 (N_426,In_1040,In_1929);
nand U427 (N_427,In_2430,In_664);
xnor U428 (N_428,In_393,In_1168);
xnor U429 (N_429,In_2070,In_1914);
nand U430 (N_430,In_1759,In_582);
or U431 (N_431,In_1897,In_1003);
nand U432 (N_432,In_1242,In_1064);
xor U433 (N_433,In_1781,In_1721);
or U434 (N_434,In_2143,In_1225);
and U435 (N_435,In_2197,In_592);
and U436 (N_436,In_1437,In_121);
or U437 (N_437,In_1265,In_2059);
xor U438 (N_438,In_2030,In_2316);
and U439 (N_439,In_790,In_355);
nand U440 (N_440,In_1404,In_1657);
nor U441 (N_441,In_1711,In_886);
nor U442 (N_442,In_2304,In_502);
nor U443 (N_443,In_1137,In_356);
and U444 (N_444,In_361,In_1270);
and U445 (N_445,In_362,In_1849);
nor U446 (N_446,In_2137,In_1915);
or U447 (N_447,In_1683,In_2087);
xnor U448 (N_448,In_1360,In_2179);
nand U449 (N_449,In_719,In_54);
nand U450 (N_450,In_2177,In_1104);
nor U451 (N_451,In_2105,In_2296);
or U452 (N_452,In_875,In_674);
nand U453 (N_453,In_833,In_1152);
or U454 (N_454,In_2246,In_795);
nand U455 (N_455,In_1525,In_1058);
or U456 (N_456,In_728,In_105);
xor U457 (N_457,In_2206,In_1706);
or U458 (N_458,In_1971,In_500);
xnor U459 (N_459,In_470,In_2339);
nand U460 (N_460,In_2032,In_1980);
xnor U461 (N_461,In_870,In_64);
xnor U462 (N_462,In_1761,In_2072);
and U463 (N_463,In_2157,In_561);
nand U464 (N_464,In_2267,In_556);
nor U465 (N_465,In_1659,In_1219);
xnor U466 (N_466,In_320,In_2078);
nor U467 (N_467,In_1217,In_1002);
nand U468 (N_468,In_1371,In_732);
or U469 (N_469,In_766,In_1793);
and U470 (N_470,In_661,In_2291);
nor U471 (N_471,In_1393,In_607);
nor U472 (N_472,In_442,In_563);
and U473 (N_473,In_729,In_277);
xnor U474 (N_474,In_1725,In_2100);
xor U475 (N_475,In_1337,In_1821);
xnor U476 (N_476,In_1286,In_1967);
nand U477 (N_477,In_405,In_1662);
nand U478 (N_478,In_986,In_937);
and U479 (N_479,In_1856,In_360);
and U480 (N_480,In_1456,In_327);
and U481 (N_481,In_1583,In_2124);
or U482 (N_482,In_1985,In_1331);
or U483 (N_483,In_1638,In_2004);
nand U484 (N_484,In_2149,In_1259);
and U485 (N_485,In_408,In_1862);
nand U486 (N_486,In_1425,In_2205);
nand U487 (N_487,In_910,In_1936);
xnor U488 (N_488,In_682,In_1876);
or U489 (N_489,In_2384,In_216);
nor U490 (N_490,In_655,In_29);
and U491 (N_491,In_2438,In_248);
nor U492 (N_492,In_1954,In_357);
xor U493 (N_493,In_1815,In_269);
nor U494 (N_494,In_16,In_508);
xnor U495 (N_495,In_1977,In_1904);
or U496 (N_496,In_1382,In_1976);
or U497 (N_497,In_1753,In_1800);
or U498 (N_498,In_980,In_1316);
xnor U499 (N_499,In_99,In_250);
or U500 (N_500,In_1722,In_1513);
nor U501 (N_501,In_751,In_1641);
nor U502 (N_502,In_844,In_545);
xnor U503 (N_503,In_1556,In_24);
or U504 (N_504,In_2456,In_231);
xnor U505 (N_505,In_2372,In_76);
and U506 (N_506,In_2442,In_1540);
or U507 (N_507,In_426,In_60);
nand U508 (N_508,In_1528,In_597);
xor U509 (N_509,In_2010,In_656);
and U510 (N_510,In_300,In_2064);
or U511 (N_511,In_2468,In_515);
nand U512 (N_512,In_1001,In_272);
or U513 (N_513,In_171,In_1519);
nor U514 (N_514,In_2306,In_465);
nand U515 (N_515,In_772,In_2066);
nand U516 (N_516,In_1413,In_1786);
nor U517 (N_517,In_479,In_1111);
and U518 (N_518,In_1069,In_2365);
nor U519 (N_519,In_988,In_2302);
xnor U520 (N_520,In_1472,In_1521);
nand U521 (N_521,In_32,In_2392);
nor U522 (N_522,In_2240,In_1505);
nand U523 (N_523,In_1285,In_215);
and U524 (N_524,In_615,In_1279);
xnor U525 (N_525,In_261,In_1172);
xor U526 (N_526,In_1806,In_2060);
nor U527 (N_527,In_1075,In_825);
nand U528 (N_528,In_488,In_533);
nor U529 (N_529,In_1245,In_959);
xnor U530 (N_530,In_1434,In_1560);
nand U531 (N_531,In_1473,In_1955);
nor U532 (N_532,In_1115,In_1699);
and U533 (N_533,In_172,In_2028);
or U534 (N_534,In_1888,In_1223);
nand U535 (N_535,In_757,In_63);
or U536 (N_536,In_780,In_1202);
xor U537 (N_537,In_707,In_2068);
or U538 (N_538,In_1484,In_798);
nand U539 (N_539,In_1804,In_157);
or U540 (N_540,In_884,In_983);
and U541 (N_541,In_1526,In_760);
and U542 (N_542,In_2287,In_1558);
nor U543 (N_543,In_400,In_2441);
nand U544 (N_544,In_1534,In_535);
and U545 (N_545,In_839,In_257);
xnor U546 (N_546,In_1877,In_1731);
nand U547 (N_547,In_206,In_940);
or U548 (N_548,In_234,In_1054);
xnor U549 (N_549,In_1664,In_1153);
nor U550 (N_550,In_1607,In_1500);
nand U551 (N_551,In_1057,In_1354);
and U552 (N_552,In_1773,In_25);
nor U553 (N_553,In_619,In_1884);
nand U554 (N_554,In_2042,In_8);
or U555 (N_555,In_1679,In_1807);
and U556 (N_556,In_690,In_1970);
xnor U557 (N_557,In_1068,In_828);
nand U558 (N_558,In_1650,In_547);
nand U559 (N_559,In_1858,In_1997);
or U560 (N_560,In_2188,In_740);
xor U561 (N_561,In_1628,In_85);
nor U562 (N_562,In_662,In_836);
and U563 (N_563,In_116,In_190);
or U564 (N_564,In_209,In_1497);
xnor U565 (N_565,In_1998,In_419);
nor U566 (N_566,In_2138,In_1963);
or U567 (N_567,In_429,In_454);
or U568 (N_568,In_1506,In_125);
or U569 (N_569,In_965,In_585);
and U570 (N_570,In_140,In_6);
nor U571 (N_571,In_1272,In_1741);
or U572 (N_572,In_2164,In_2199);
nand U573 (N_573,In_282,In_1633);
nand U574 (N_574,In_1571,In_1351);
nand U575 (N_575,In_1615,In_1444);
and U576 (N_576,In_1253,In_477);
nor U577 (N_577,In_1656,In_2252);
nor U578 (N_578,In_548,In_126);
nand U579 (N_579,In_1319,In_1375);
and U580 (N_580,In_596,In_1522);
nor U581 (N_581,In_768,In_2014);
nor U582 (N_582,In_934,In_2140);
or U583 (N_583,In_158,In_1660);
and U584 (N_584,In_460,In_2248);
or U585 (N_585,In_1140,In_1952);
nand U586 (N_586,In_1859,In_1871);
or U587 (N_587,In_109,In_418);
nor U588 (N_588,In_572,In_1563);
or U589 (N_589,In_1452,In_1165);
nor U590 (N_590,In_2404,In_1823);
or U591 (N_591,In_1097,In_2387);
xnor U592 (N_592,In_1333,In_1917);
and U593 (N_593,In_2196,In_1697);
and U594 (N_594,In_2368,In_79);
and U595 (N_595,In_1116,In_2412);
and U596 (N_596,In_1890,In_335);
nand U597 (N_597,In_1578,In_649);
and U598 (N_598,In_2096,In_2402);
nor U599 (N_599,In_112,In_985);
nand U600 (N_600,In_2204,In_1764);
or U601 (N_601,In_1141,In_2464);
nand U602 (N_602,In_663,In_799);
xor U603 (N_603,In_373,In_2173);
or U604 (N_604,In_1142,In_1386);
nor U605 (N_605,In_1277,In_1364);
or U606 (N_606,In_2300,In_1992);
xnor U607 (N_607,In_1973,In_2063);
nor U608 (N_608,In_1698,In_1039);
xnor U609 (N_609,In_1676,In_653);
and U610 (N_610,In_1006,In_285);
nand U611 (N_611,In_2481,In_297);
or U612 (N_612,In_802,In_913);
or U613 (N_613,In_324,In_1586);
nand U614 (N_614,In_443,In_2447);
nor U615 (N_615,In_198,In_2145);
or U616 (N_616,In_323,In_1603);
xnor U617 (N_617,In_2425,In_1885);
and U618 (N_618,In_13,In_540);
nor U619 (N_619,In_1278,In_809);
xnor U620 (N_620,In_424,In_2293);
xor U621 (N_621,In_263,In_1878);
nor U622 (N_622,In_2343,In_44);
or U623 (N_623,In_1739,In_2378);
nor U624 (N_624,In_1210,In_463);
and U625 (N_625,In_9,In_2480);
nor U626 (N_626,In_1029,In_1944);
xnor U627 (N_627,In_1964,In_1625);
and U628 (N_628,In_62,In_2390);
nor U629 (N_629,In_2288,In_1212);
and U630 (N_630,In_302,In_57);
xor U631 (N_631,In_2181,In_2309);
nand U632 (N_632,In_623,In_1388);
xor U633 (N_633,In_1546,In_219);
nand U634 (N_634,In_1591,In_1910);
xnor U635 (N_635,In_512,In_2381);
or U636 (N_636,In_2215,In_278);
or U637 (N_637,In_296,In_665);
and U638 (N_638,In_688,In_2150);
nand U639 (N_639,In_903,In_754);
or U640 (N_640,In_1471,In_679);
and U641 (N_641,In_120,In_1704);
xor U642 (N_642,In_2058,In_1109);
or U643 (N_643,In_1175,In_856);
and U644 (N_644,In_689,In_200);
xnor U645 (N_645,In_936,In_2029);
and U646 (N_646,In_1275,In_2281);
and U647 (N_647,In_281,In_2254);
nand U648 (N_648,In_1032,In_1258);
nor U649 (N_649,In_1093,In_2393);
nand U650 (N_650,In_2420,In_2201);
or U651 (N_651,In_1767,In_2345);
and U652 (N_652,In_2278,In_1482);
nor U653 (N_653,In_111,In_599);
nand U654 (N_654,In_181,In_1428);
xor U655 (N_655,In_2261,In_2495);
nor U656 (N_656,In_645,In_1527);
nand U657 (N_657,In_1694,In_23);
or U658 (N_658,In_1236,In_2397);
nor U659 (N_659,In_1986,In_1199);
and U660 (N_660,In_1120,In_1512);
xor U661 (N_661,In_1935,In_2294);
nor U662 (N_662,In_309,In_1293);
or U663 (N_663,In_11,In_1329);
nor U664 (N_664,In_1306,In_366);
or U665 (N_665,In_218,In_897);
nand U666 (N_666,In_474,In_1652);
nor U667 (N_667,In_245,In_332);
xor U668 (N_668,In_267,In_2080);
or U669 (N_669,In_2023,In_552);
nand U670 (N_670,In_2486,In_1406);
nor U671 (N_671,In_1352,In_646);
and U672 (N_672,In_59,In_2233);
nor U673 (N_673,In_1488,In_1632);
xor U674 (N_674,In_1464,In_1356);
nor U675 (N_675,In_553,In_1844);
nor U676 (N_676,In_650,In_1569);
and U677 (N_677,In_1649,In_178);
or U678 (N_678,In_2093,In_1498);
and U679 (N_679,In_2110,In_1854);
and U680 (N_680,In_1192,In_204);
xor U681 (N_681,In_1752,In_1948);
nor U682 (N_682,In_2168,In_1671);
and U683 (N_683,In_1588,In_1357);
nand U684 (N_684,In_193,In_4);
and U685 (N_685,In_1991,In_98);
and U686 (N_686,In_2342,In_916);
xor U687 (N_687,In_503,In_336);
nand U688 (N_688,In_2363,In_605);
and U689 (N_689,In_1340,In_537);
xor U690 (N_690,In_1431,In_1151);
nor U691 (N_691,In_2355,In_1802);
xor U692 (N_692,In_2358,In_1837);
nor U693 (N_693,In_1566,In_670);
nand U694 (N_694,In_92,In_236);
nor U695 (N_695,In_827,In_283);
and U696 (N_696,In_262,In_1449);
nand U697 (N_697,In_317,In_1593);
nor U698 (N_698,In_227,In_1870);
xnor U699 (N_699,In_1620,In_430);
xor U700 (N_700,In_2426,In_188);
or U701 (N_701,In_1370,In_1777);
nor U702 (N_702,In_2401,In_314);
nor U703 (N_703,In_1174,In_1389);
and U704 (N_704,In_1113,In_1330);
nor U705 (N_705,In_922,In_293);
nor U706 (N_706,In_1020,In_1328);
or U707 (N_707,In_238,In_351);
xnor U708 (N_708,In_2013,In_923);
and U709 (N_709,In_776,In_1939);
nor U710 (N_710,In_1320,In_478);
or U711 (N_711,In_2285,In_2472);
xnor U712 (N_712,In_1987,In_1451);
and U713 (N_713,In_1281,In_1984);
and U714 (N_714,In_1461,In_1195);
nand U715 (N_715,In_2104,In_1923);
nor U716 (N_716,In_968,In_156);
and U717 (N_717,In_654,In_70);
xnor U718 (N_718,In_834,In_1303);
nand U719 (N_719,In_1269,In_2431);
xor U720 (N_720,In_427,In_1623);
nor U721 (N_721,In_2115,In_497);
and U722 (N_722,In_1532,In_2335);
and U723 (N_723,In_816,In_365);
or U724 (N_724,In_370,In_66);
or U725 (N_725,In_1928,In_1724);
and U726 (N_726,In_991,In_1298);
nor U727 (N_727,In_733,In_2082);
or U728 (N_728,In_939,In_475);
nand U729 (N_729,In_1919,In_2380);
nor U730 (N_730,In_82,In_1372);
xnor U731 (N_731,In_2348,In_1469);
nand U732 (N_732,In_420,In_2416);
nor U733 (N_733,In_19,In_40);
nor U734 (N_734,In_1125,In_2245);
nand U735 (N_735,In_893,In_2130);
nand U736 (N_736,In_1076,In_1088);
nand U737 (N_737,In_549,In_2490);
or U738 (N_738,In_367,In_854);
nor U739 (N_739,In_917,In_2053);
xnor U740 (N_740,In_695,In_2015);
xnor U741 (N_741,In_1631,In_173);
and U742 (N_742,In_814,In_1663);
nand U743 (N_743,In_848,In_1703);
and U744 (N_744,In_704,In_1643);
nand U745 (N_745,In_1670,In_837);
xnor U746 (N_746,In_487,In_1925);
or U747 (N_747,In_2409,In_2450);
and U748 (N_748,In_2375,In_1760);
xor U749 (N_749,In_1966,In_1668);
or U750 (N_750,In_821,In_2427);
and U751 (N_751,In_1123,In_624);
nand U752 (N_752,In_714,In_177);
nor U753 (N_753,In_1311,In_30);
nand U754 (N_754,In_310,In_2317);
xor U755 (N_755,In_328,In_1263);
nand U756 (N_756,In_1178,In_1268);
nor U757 (N_757,In_1264,In_1274);
or U758 (N_758,In_2022,In_840);
and U759 (N_759,In_1391,In_1239);
xnor U760 (N_760,In_1684,In_528);
and U761 (N_761,In_738,In_693);
nor U762 (N_762,In_152,In_1609);
xor U763 (N_763,In_1771,In_1273);
and U764 (N_764,In_350,In_1401);
nor U765 (N_765,In_201,In_1126);
and U766 (N_766,In_1574,In_1083);
xor U767 (N_767,In_2142,In_2090);
nor U768 (N_768,In_1408,In_2113);
xor U769 (N_769,In_977,In_1589);
nor U770 (N_770,In_1750,In_294);
xnor U771 (N_771,In_1790,In_1538);
and U772 (N_772,In_52,In_1769);
or U773 (N_773,In_1289,In_5);
xor U774 (N_774,In_1074,In_778);
xnor U775 (N_775,In_202,In_960);
and U776 (N_776,In_1665,In_141);
nor U777 (N_777,In_2154,In_2089);
nor U778 (N_778,In_1658,In_1733);
nor U779 (N_779,In_402,In_2194);
nor U780 (N_780,In_1487,In_996);
or U781 (N_781,In_1612,In_1795);
nand U782 (N_782,In_409,In_334);
nand U783 (N_783,In_2413,In_943);
nor U784 (N_784,In_1173,In_2483);
or U785 (N_785,In_1490,In_1127);
and U786 (N_786,In_1701,In_189);
nor U787 (N_787,In_89,In_446);
xnor U788 (N_788,In_1515,In_1106);
xor U789 (N_789,In_617,In_447);
nand U790 (N_790,In_1734,In_2183);
xor U791 (N_791,In_1420,In_1635);
xnor U792 (N_792,In_949,In_692);
xnor U793 (N_793,In_2470,In_610);
xor U794 (N_794,In_1717,In_2024);
xnor U795 (N_795,In_1440,In_2315);
nand U796 (N_796,In_1302,In_767);
nor U797 (N_797,In_2329,In_2050);
or U798 (N_798,In_1066,In_1705);
xnor U799 (N_799,In_964,In_2187);
and U800 (N_800,In_1296,In_1121);
nor U801 (N_801,In_950,In_2009);
xor U802 (N_802,In_801,In_575);
and U803 (N_803,In_542,In_587);
nand U804 (N_804,In_1868,In_1280);
or U805 (N_805,In_997,In_1157);
or U806 (N_806,In_1496,In_2360);
nand U807 (N_807,In_80,In_249);
nor U808 (N_808,In_1347,In_603);
nand U809 (N_809,In_93,In_2421);
or U810 (N_810,In_73,In_2189);
nand U811 (N_811,In_339,In_810);
nand U812 (N_812,In_1742,In_993);
xor U813 (N_813,In_1938,In_1180);
xnor U814 (N_814,In_794,In_1091);
or U815 (N_815,In_2349,In_226);
nand U816 (N_816,In_1946,In_346);
nor U817 (N_817,In_2175,In_1869);
nand U818 (N_818,In_867,In_1412);
nand U819 (N_819,In_1014,In_205);
xnor U820 (N_820,In_270,In_1774);
nor U821 (N_821,In_1220,In_1085);
nand U822 (N_822,In_999,In_882);
and U823 (N_823,In_1166,In_223);
or U824 (N_824,In_1056,In_629);
or U825 (N_825,In_1435,In_1714);
nor U826 (N_826,In_1894,In_2039);
nor U827 (N_827,In_1716,In_804);
nand U828 (N_828,In_2035,In_792);
xor U829 (N_829,In_1443,In_576);
xnor U830 (N_830,In_594,In_145);
xnor U831 (N_831,In_1033,In_1214);
and U832 (N_832,In_233,In_2081);
or U833 (N_833,In_672,In_2435);
nor U834 (N_834,In_1875,In_524);
and U835 (N_835,In_787,In_390);
nand U836 (N_836,In_571,In_2276);
and U837 (N_837,In_117,In_1315);
nand U838 (N_838,In_1133,In_1775);
nand U839 (N_839,In_1709,In_2147);
nor U840 (N_840,In_48,In_1517);
nand U841 (N_841,In_2465,In_304);
nor U842 (N_842,In_2436,In_667);
and U843 (N_843,In_1602,In_1305);
xnor U844 (N_844,In_1082,In_604);
xor U845 (N_845,In_536,In_1667);
or U846 (N_846,In_224,In_306);
xnor U847 (N_847,In_921,In_919);
or U848 (N_848,In_1101,In_1956);
xor U849 (N_849,In_1818,In_1840);
xor U850 (N_850,In_1261,In_2065);
and U851 (N_851,In_1015,In_1358);
or U852 (N_852,In_1457,In_730);
and U853 (N_853,In_868,In_1063);
nand U854 (N_854,In_1055,In_2129);
xnor U855 (N_855,In_1042,In_2226);
xnor U856 (N_856,In_2218,In_1957);
or U857 (N_857,In_544,In_2289);
nor U858 (N_858,In_595,In_1695);
nand U859 (N_859,In_1920,In_895);
and U860 (N_860,In_2251,In_358);
nor U861 (N_861,In_1299,In_1865);
and U862 (N_862,In_2391,In_217);
nand U863 (N_863,In_2445,In_75);
and U864 (N_864,In_2214,In_2295);
nor U865 (N_865,In_1335,In_1881);
nor U866 (N_866,In_2139,In_466);
or U867 (N_867,In_1640,In_1004);
nor U868 (N_868,In_684,In_1902);
nand U869 (N_869,In_797,In_1879);
nand U870 (N_870,In_242,In_1414);
nor U871 (N_871,In_311,In_2001);
xnor U872 (N_872,In_2128,In_1502);
nor U873 (N_873,In_1924,In_771);
nand U874 (N_874,In_431,In_1732);
or U875 (N_875,In_1776,In_1025);
xnor U876 (N_876,In_2202,In_1950);
nand U877 (N_877,In_2033,In_2192);
nor U878 (N_878,In_639,In_2242);
xor U879 (N_879,In_1891,In_467);
nand U880 (N_880,In_724,In_784);
nand U881 (N_881,In_660,In_1642);
and U882 (N_882,In_614,In_2389);
or U883 (N_883,In_1061,In_2026);
xor U884 (N_884,In_632,In_1892);
xor U885 (N_885,In_2158,In_1079);
xnor U886 (N_886,In_1154,In_1508);
nor U887 (N_887,In_2229,In_618);
and U888 (N_888,In_1824,In_691);
xnor U889 (N_889,In_435,In_1394);
or U890 (N_890,In_1845,In_1424);
nor U891 (N_891,In_2270,In_1613);
nand U892 (N_892,In_1150,In_842);
nand U893 (N_893,In_739,In_786);
nand U894 (N_894,In_862,In_994);
nand U895 (N_895,In_577,In_2049);
or U896 (N_896,In_71,In_1049);
xor U897 (N_897,In_2367,In_119);
xor U898 (N_898,In_748,In_706);
and U899 (N_899,In_849,In_225);
or U900 (N_900,In_2225,In_1937);
nor U901 (N_901,In_2109,In_398);
nor U902 (N_902,In_1200,In_1646);
or U903 (N_903,In_574,In_1995);
and U904 (N_904,In_1661,In_1392);
or U905 (N_905,In_289,In_1246);
nor U906 (N_906,In_1565,In_793);
nand U907 (N_907,In_2102,In_815);
and U908 (N_908,In_2132,In_562);
nor U909 (N_909,In_1072,In_567);
nand U910 (N_910,In_954,In_2054);
and U911 (N_911,In_239,In_811);
nor U912 (N_912,In_636,In_1149);
nor U913 (N_913,In_1046,In_1080);
xnor U914 (N_914,In_931,In_2324);
xnor U915 (N_915,In_379,In_241);
nor U916 (N_916,In_621,In_1445);
nor U917 (N_917,In_734,In_657);
and U918 (N_918,In_1834,In_433);
and U919 (N_919,In_1911,In_2386);
nor U920 (N_920,In_1402,In_1327);
and U921 (N_921,In_2422,In_2131);
nor U922 (N_922,In_1244,In_1019);
nor U923 (N_923,In_160,In_425);
nor U924 (N_924,In_2493,In_345);
or U925 (N_925,In_2170,In_2083);
or U926 (N_926,In_94,In_1204);
nand U927 (N_927,In_113,In_1730);
nand U928 (N_928,In_2357,In_404);
nor U929 (N_929,In_2238,In_702);
and U930 (N_930,In_1548,In_1562);
nor U931 (N_931,In_613,In_2325);
and U932 (N_932,In_1531,In_2340);
xnor U933 (N_933,In_1476,In_1794);
nand U934 (N_934,In_2041,In_1751);
and U935 (N_935,In_491,In_806);
xor U936 (N_936,In_2095,In_2182);
nor U937 (N_937,In_685,In_1283);
nand U938 (N_938,In_132,In_2444);
xnor U939 (N_939,In_673,In_2027);
nand U940 (N_940,In_12,In_1803);
nand U941 (N_941,In_169,In_380);
or U942 (N_942,In_1715,In_1882);
or U943 (N_943,In_1348,In_1181);
and U944 (N_944,In_222,In_2075);
or U945 (N_945,In_1828,In_915);
or U946 (N_946,In_1568,In_1779);
and U947 (N_947,In_1810,In_2055);
nor U948 (N_948,In_1489,In_1383);
and U949 (N_949,In_1287,In_102);
or U950 (N_950,In_482,In_995);
nor U951 (N_951,In_1552,In_464);
nor U952 (N_952,In_1688,In_1624);
or U953 (N_953,In_455,In_637);
or U954 (N_954,In_711,In_2411);
xor U955 (N_955,In_2250,In_1385);
nor U956 (N_956,In_680,In_1084);
nor U957 (N_957,In_2399,In_376);
xnor U958 (N_958,In_322,In_1808);
nor U959 (N_959,In_1071,In_1201);
nor U960 (N_960,In_1922,In_1477);
nor U961 (N_961,In_1645,In_1989);
nor U962 (N_962,In_414,In_1459);
xor U963 (N_963,In_883,In_2376);
xor U964 (N_964,In_2006,In_208);
nor U965 (N_965,In_2191,In_1355);
xor U966 (N_966,In_2067,In_2031);
xor U967 (N_967,In_1237,In_1365);
or U968 (N_968,In_925,In_240);
or U969 (N_969,In_1763,In_2044);
nor U970 (N_970,In_1754,In_1059);
nand U971 (N_971,In_978,In_436);
xor U972 (N_972,In_1387,In_2230);
nand U973 (N_973,In_666,In_557);
nor U974 (N_974,In_348,In_2274);
nor U975 (N_975,In_18,In_110);
nor U976 (N_976,In_1416,In_1700);
nor U977 (N_977,In_912,In_2271);
or U978 (N_978,In_496,In_1672);
or U979 (N_979,In_1060,In_808);
and U980 (N_980,In_805,In_1164);
nand U981 (N_981,In_1012,In_375);
nor U982 (N_982,In_377,In_1792);
or U983 (N_983,In_1290,In_705);
and U984 (N_984,In_1983,In_1825);
or U985 (N_985,In_2428,In_2264);
nand U986 (N_986,In_1380,In_775);
and U987 (N_987,In_2383,In_1108);
nor U988 (N_988,In_1608,In_371);
xor U989 (N_989,In_2094,In_2056);
nor U990 (N_990,In_634,In_853);
xor U991 (N_991,In_697,In_2232);
or U992 (N_992,In_303,In_881);
nor U993 (N_993,In_1218,In_1846);
or U994 (N_994,In_755,In_880);
nor U995 (N_995,In_709,In_1398);
nand U996 (N_996,In_527,In_1727);
or U997 (N_997,In_271,In_2379);
or U998 (N_998,In_1468,In_2362);
and U999 (N_999,In_1842,In_1208);
nand U1000 (N_1000,In_308,In_1543);
xnor U1001 (N_1001,In_514,In_165);
or U1002 (N_1002,In_131,In_2432);
xor U1003 (N_1003,In_1981,In_480);
and U1004 (N_1004,In_1034,In_1317);
and U1005 (N_1005,In_321,In_659);
nor U1006 (N_1006,In_211,In_1067);
nand U1007 (N_1007,In_579,In_752);
xnor U1008 (N_1008,In_1209,In_551);
nor U1009 (N_1009,In_1696,In_753);
or U1010 (N_1010,In_2332,In_83);
or U1011 (N_1011,In_489,In_1177);
xnor U1012 (N_1012,In_130,In_2307);
nor U1013 (N_1013,In_1363,In_1974);
nor U1014 (N_1014,In_1719,In_845);
nand U1015 (N_1015,In_2249,In_889);
nand U1016 (N_1016,In_163,In_1618);
nand U1017 (N_1017,In_2463,In_313);
and U1018 (N_1018,In_1117,In_1323);
or U1019 (N_1019,In_1222,In_1788);
nand U1020 (N_1020,In_584,In_1850);
or U1021 (N_1021,In_859,In_832);
xor U1022 (N_1022,In_337,In_1211);
nand U1023 (N_1023,In_2111,In_383);
nor U1024 (N_1024,In_522,In_312);
xnor U1025 (N_1025,In_1587,In_2352);
nand U1026 (N_1026,In_1594,In_909);
nor U1027 (N_1027,In_2007,In_106);
and U1028 (N_1028,In_1092,In_1901);
or U1029 (N_1029,In_1198,In_2136);
nand U1030 (N_1030,In_941,In_1017);
or U1031 (N_1031,In_2458,In_957);
nor U1032 (N_1032,In_1334,In_2478);
or U1033 (N_1033,In_914,In_305);
nor U1034 (N_1034,In_1310,In_17);
xor U1035 (N_1035,In_1585,In_2408);
nand U1036 (N_1036,In_608,In_396);
nand U1037 (N_1037,In_1373,In_1241);
nor U1038 (N_1038,In_852,In_857);
nand U1039 (N_1039,In_750,In_1018);
or U1040 (N_1040,In_2498,In_1692);
nor U1041 (N_1041,In_1439,In_669);
nand U1042 (N_1042,In_260,In_138);
and U1043 (N_1043,In_2045,In_824);
nor U1044 (N_1044,In_1132,In_1799);
xnor U1045 (N_1045,In_1965,In_1147);
nand U1046 (N_1046,In_1880,In_1171);
nor U1047 (N_1047,In_2346,In_72);
nor U1048 (N_1048,In_468,In_153);
or U1049 (N_1049,In_1390,In_213);
xnor U1050 (N_1050,In_288,In_2351);
nor U1051 (N_1051,In_1037,In_2320);
nor U1052 (N_1052,In_2312,In_507);
xnor U1053 (N_1053,In_1359,In_855);
or U1054 (N_1054,In_894,In_457);
xnor U1055 (N_1055,In_625,In_2469);
xor U1056 (N_1056,In_721,In_580);
xnor U1057 (N_1057,In_2474,In_2195);
and U1058 (N_1058,In_1462,In_1893);
xnor U1059 (N_1059,In_273,In_2012);
xor U1060 (N_1060,In_1826,In_1470);
or U1061 (N_1061,In_546,In_1932);
nand U1062 (N_1062,In_1288,In_2000);
and U1063 (N_1063,In_1690,In_1707);
xor U1064 (N_1064,In_2403,In_1755);
nand U1065 (N_1065,In_401,In_761);
xor U1066 (N_1066,In_1160,In_1243);
nor U1067 (N_1067,In_1536,In_199);
and U1068 (N_1068,In_55,In_2440);
nor U1069 (N_1069,In_764,In_1344);
xor U1070 (N_1070,In_53,In_438);
or U1071 (N_1071,In_1176,In_2073);
xnor U1072 (N_1072,In_2002,In_1949);
and U1073 (N_1073,In_2303,In_292);
nor U1074 (N_1074,In_1162,In_501);
xnor U1075 (N_1075,In_1582,In_741);
xor U1076 (N_1076,In_686,In_1990);
nor U1077 (N_1077,In_1215,In_606);
xnor U1078 (N_1078,In_1947,In_1124);
xnor U1079 (N_1079,In_1158,In_2255);
nor U1080 (N_1080,In_2350,In_2219);
nor U1081 (N_1081,In_1766,In_641);
nand U1082 (N_1082,In_2473,In_1942);
nand U1083 (N_1083,In_1510,In_2338);
or U1084 (N_1084,In_2216,In_1889);
nand U1085 (N_1085,In_392,In_696);
nor U1086 (N_1086,In_745,In_1988);
xnor U1087 (N_1087,In_2159,In_1070);
and U1088 (N_1088,In_558,In_1000);
and U1089 (N_1089,In_432,In_164);
or U1090 (N_1090,In_2037,In_2298);
nor U1091 (N_1091,In_1945,In_523);
or U1092 (N_1092,In_1702,In_2305);
nand U1093 (N_1093,In_1136,In_1908);
xnor U1094 (N_1094,In_406,In_763);
or U1095 (N_1095,In_129,In_2207);
nor U1096 (N_1096,In_1415,In_2227);
xor U1097 (N_1097,In_2361,In_2084);
nand U1098 (N_1098,In_2268,In_2116);
or U1099 (N_1099,In_1555,In_1579);
nor U1100 (N_1100,In_892,In_1809);
and U1101 (N_1101,In_1008,In_826);
nor U1102 (N_1102,In_1680,In_1148);
nand U1103 (N_1103,In_2460,In_1913);
nor U1104 (N_1104,In_1514,In_1848);
and U1105 (N_1105,In_280,In_1203);
nand U1106 (N_1106,In_1224,In_998);
nor U1107 (N_1107,In_1930,In_564);
or U1108 (N_1108,In_2314,In_39);
and U1109 (N_1109,In_2017,In_1186);
nand U1110 (N_1110,In_127,In_485);
xor U1111 (N_1111,In_411,In_717);
or U1112 (N_1112,In_96,In_2244);
nand U1113 (N_1113,In_591,In_1028);
or U1114 (N_1114,In_246,In_2098);
or U1115 (N_1115,In_1129,In_2005);
or U1116 (N_1116,In_1249,In_1441);
and U1117 (N_1117,In_2103,In_1267);
nand U1118 (N_1118,In_1978,In_143);
xor U1119 (N_1119,In_68,In_1590);
or U1120 (N_1120,In_835,In_1738);
and U1121 (N_1121,In_2146,In_1503);
nand U1122 (N_1122,In_183,In_1756);
or U1123 (N_1123,In_1551,In_846);
xnor U1124 (N_1124,In_2423,In_1465);
and U1125 (N_1125,In_2424,In_2322);
nand U1126 (N_1126,In_1654,In_1720);
nand U1127 (N_1127,In_1096,In_2290);
or U1128 (N_1128,In_876,In_1043);
or U1129 (N_1129,In_2163,In_803);
nor U1130 (N_1130,In_118,In_1499);
xnor U1131 (N_1131,In_101,In_1081);
or U1132 (N_1132,In_484,In_1381);
nor U1133 (N_1133,In_1604,In_781);
xnor U1134 (N_1134,In_2036,In_589);
or U1135 (N_1135,In_252,In_710);
and U1136 (N_1136,In_1432,In_61);
xor U1137 (N_1137,In_2301,In_1235);
nor U1138 (N_1138,In_1648,In_36);
xor U1139 (N_1139,In_459,In_58);
nand U1140 (N_1140,In_2141,In_2155);
nor U1141 (N_1141,In_989,In_1238);
or U1142 (N_1142,In_2280,In_1959);
nand U1143 (N_1143,In_1723,In_84);
nand U1144 (N_1144,In_736,In_796);
nor U1145 (N_1145,In_493,In_519);
and U1146 (N_1146,In_395,In_878);
nor U1147 (N_1147,In_1221,In_1475);
nor U1148 (N_1148,In_298,In_1601);
and U1149 (N_1149,In_2385,In_900);
and U1150 (N_1150,In_1943,In_1188);
nor U1151 (N_1151,In_1639,In_967);
and U1152 (N_1152,In_947,In_1256);
nand U1153 (N_1153,In_1062,In_642);
xor U1154 (N_1154,In_2326,In_2263);
xnor U1155 (N_1155,In_1843,In_368);
or U1156 (N_1156,In_1861,In_1338);
nor U1157 (N_1157,In_640,In_399);
xnor U1158 (N_1158,In_1912,In_1561);
xor U1159 (N_1159,In_95,In_1898);
or U1160 (N_1160,In_1979,In_2356);
nand U1161 (N_1161,In_1516,In_1301);
nor U1162 (N_1162,In_149,In_948);
or U1163 (N_1163,In_1762,In_2125);
nor U1164 (N_1164,In_21,In_1065);
nor U1165 (N_1165,In_1361,In_749);
and U1166 (N_1166,In_822,In_785);
xor U1167 (N_1167,In_1501,In_2119);
nor U1168 (N_1168,In_1254,In_448);
nand U1169 (N_1169,In_1797,In_1099);
or U1170 (N_1170,In_1193,In_486);
nor U1171 (N_1171,In_1993,In_2259);
nor U1172 (N_1172,In_1934,In_187);
and U1173 (N_1173,In_2446,In_2479);
xnor U1174 (N_1174,In_1022,In_56);
nor U1175 (N_1175,In_2282,In_2265);
xor U1176 (N_1176,In_1554,In_873);
nor U1177 (N_1177,In_28,In_1830);
xor U1178 (N_1178,In_2336,In_254);
nor U1179 (N_1179,In_381,In_756);
xnor U1180 (N_1180,In_1855,In_329);
and U1181 (N_1181,In_1170,In_1529);
and U1182 (N_1182,In_437,In_1636);
nor U1183 (N_1183,In_1726,In_658);
xnor U1184 (N_1184,In_1595,In_128);
and U1185 (N_1185,In_847,In_2418);
xor U1186 (N_1186,In_2091,In_1087);
xnor U1187 (N_1187,In_88,In_1005);
and U1188 (N_1188,In_2366,In_275);
nor U1189 (N_1189,In_1321,In_2434);
xnor U1190 (N_1190,In_2433,In_2260);
xnor U1191 (N_1191,In_265,In_452);
nand U1192 (N_1192,In_2462,In_782);
nor U1193 (N_1193,In_731,In_2092);
nor U1194 (N_1194,In_1326,In_151);
xor U1195 (N_1195,In_843,In_2243);
xnor U1196 (N_1196,In_2186,In_1909);
nand U1197 (N_1197,In_765,In_453);
and U1198 (N_1198,In_1839,In_232);
nor U1199 (N_1199,In_1023,In_410);
nor U1200 (N_1200,In_942,In_43);
nand U1201 (N_1201,In_555,In_472);
and U1202 (N_1202,In_568,In_1962);
xnor U1203 (N_1203,In_144,In_722);
xor U1204 (N_1204,In_2333,In_946);
and U1205 (N_1205,In_1577,In_885);
nand U1206 (N_1206,In_1345,In_506);
or U1207 (N_1207,In_2018,In_779);
xnor U1208 (N_1208,In_2318,In_962);
xor U1209 (N_1209,In_1682,In_1041);
nor U1210 (N_1210,In_1207,In_1252);
and U1211 (N_1211,In_1570,In_879);
and U1212 (N_1212,In_1559,In_1867);
and U1213 (N_1213,In_244,In_1248);
and U1214 (N_1214,In_1378,In_1573);
nor U1215 (N_1215,In_1817,In_1118);
nor U1216 (N_1216,In_1460,In_622);
xnor U1217 (N_1217,In_984,In_1206);
nand U1218 (N_1218,In_2184,In_286);
nand U1219 (N_1219,In_2266,In_698);
nor U1220 (N_1220,In_1940,In_458);
xnor U1221 (N_1221,In_933,In_1455);
xor U1222 (N_1222,In_1677,In_1864);
and U1223 (N_1223,In_1478,In_531);
nand U1224 (N_1224,In_498,In_2499);
xor U1225 (N_1225,In_2021,In_2185);
and U1226 (N_1226,In_930,In_1089);
and U1227 (N_1227,In_2269,In_107);
and U1228 (N_1228,In_1900,In_49);
and U1229 (N_1229,In_864,In_1098);
or U1230 (N_1230,In_2382,In_2388);
nor U1231 (N_1231,In_1295,In_403);
and U1232 (N_1232,In_1647,In_1384);
nand U1233 (N_1233,In_1031,In_2313);
nand U1234 (N_1234,In_865,In_15);
xor U1235 (N_1235,In_274,In_737);
and U1236 (N_1236,In_369,In_108);
nand U1237 (N_1237,In_338,In_1621);
and U1238 (N_1238,In_1523,In_2415);
and U1239 (N_1239,In_1530,In_69);
nor U1240 (N_1240,In_1144,In_230);
and U1241 (N_1241,In_1822,In_228);
xor U1242 (N_1242,In_90,In_1627);
xnor U1243 (N_1243,In_1257,In_1376);
nor U1244 (N_1244,In_1368,In_725);
nor U1245 (N_1245,In_2410,In_1429);
and U1246 (N_1246,In_1100,In_2494);
and U1247 (N_1247,In_652,In_1271);
or U1248 (N_1248,In_861,In_1598);
or U1249 (N_1249,In_703,In_1292);
or U1250 (N_1250,In_1597,In_63);
nand U1251 (N_1251,In_1371,In_641);
and U1252 (N_1252,In_104,In_92);
nand U1253 (N_1253,In_1630,In_2280);
or U1254 (N_1254,In_1932,In_334);
nand U1255 (N_1255,In_2048,In_6);
nor U1256 (N_1256,In_336,In_1080);
nor U1257 (N_1257,In_383,In_962);
nor U1258 (N_1258,In_1217,In_1869);
nor U1259 (N_1259,In_1827,In_1860);
nor U1260 (N_1260,In_2274,In_2072);
xor U1261 (N_1261,In_1336,In_1219);
and U1262 (N_1262,In_1103,In_1949);
xor U1263 (N_1263,In_594,In_245);
or U1264 (N_1264,In_302,In_287);
nand U1265 (N_1265,In_1578,In_2245);
or U1266 (N_1266,In_2380,In_1732);
xnor U1267 (N_1267,In_333,In_2328);
or U1268 (N_1268,In_458,In_1530);
nor U1269 (N_1269,In_344,In_432);
and U1270 (N_1270,In_2495,In_40);
nor U1271 (N_1271,In_1454,In_683);
nor U1272 (N_1272,In_324,In_1358);
nand U1273 (N_1273,In_1114,In_199);
xor U1274 (N_1274,In_1930,In_1649);
and U1275 (N_1275,In_350,In_351);
and U1276 (N_1276,In_1568,In_125);
xor U1277 (N_1277,In_1173,In_977);
or U1278 (N_1278,In_1608,In_1953);
and U1279 (N_1279,In_1230,In_296);
xor U1280 (N_1280,In_273,In_120);
nand U1281 (N_1281,In_1449,In_1957);
nand U1282 (N_1282,In_2446,In_1432);
nand U1283 (N_1283,In_298,In_57);
nor U1284 (N_1284,In_2430,In_854);
or U1285 (N_1285,In_1469,In_695);
and U1286 (N_1286,In_1347,In_1264);
or U1287 (N_1287,In_1469,In_155);
nand U1288 (N_1288,In_1912,In_960);
or U1289 (N_1289,In_2108,In_1996);
and U1290 (N_1290,In_1728,In_1240);
nand U1291 (N_1291,In_1763,In_1771);
or U1292 (N_1292,In_2400,In_507);
xor U1293 (N_1293,In_638,In_1636);
or U1294 (N_1294,In_587,In_12);
nand U1295 (N_1295,In_883,In_2080);
nor U1296 (N_1296,In_66,In_2082);
and U1297 (N_1297,In_82,In_590);
or U1298 (N_1298,In_1510,In_1772);
or U1299 (N_1299,In_1412,In_2449);
xnor U1300 (N_1300,In_489,In_249);
or U1301 (N_1301,In_2402,In_333);
nand U1302 (N_1302,In_1219,In_2077);
nand U1303 (N_1303,In_1521,In_1456);
and U1304 (N_1304,In_1248,In_947);
or U1305 (N_1305,In_306,In_1525);
xor U1306 (N_1306,In_82,In_1469);
or U1307 (N_1307,In_1813,In_981);
xnor U1308 (N_1308,In_1704,In_1875);
and U1309 (N_1309,In_76,In_228);
nand U1310 (N_1310,In_471,In_920);
nand U1311 (N_1311,In_604,In_2047);
xnor U1312 (N_1312,In_1031,In_759);
nand U1313 (N_1313,In_1952,In_2229);
xnor U1314 (N_1314,In_151,In_621);
nor U1315 (N_1315,In_9,In_1461);
nor U1316 (N_1316,In_108,In_2491);
nor U1317 (N_1317,In_1843,In_486);
or U1318 (N_1318,In_2399,In_365);
xor U1319 (N_1319,In_325,In_439);
xor U1320 (N_1320,In_613,In_1282);
nand U1321 (N_1321,In_1343,In_126);
nand U1322 (N_1322,In_321,In_722);
or U1323 (N_1323,In_187,In_142);
xor U1324 (N_1324,In_2019,In_1324);
nor U1325 (N_1325,In_1207,In_1523);
nand U1326 (N_1326,In_1398,In_1854);
nand U1327 (N_1327,In_1707,In_886);
or U1328 (N_1328,In_1148,In_1111);
xor U1329 (N_1329,In_1916,In_170);
or U1330 (N_1330,In_1643,In_73);
nor U1331 (N_1331,In_852,In_14);
nand U1332 (N_1332,In_1695,In_1240);
xnor U1333 (N_1333,In_1596,In_46);
nor U1334 (N_1334,In_1924,In_2495);
and U1335 (N_1335,In_2496,In_1186);
or U1336 (N_1336,In_2093,In_2109);
or U1337 (N_1337,In_150,In_729);
or U1338 (N_1338,In_682,In_2350);
nor U1339 (N_1339,In_375,In_616);
nand U1340 (N_1340,In_993,In_2048);
nor U1341 (N_1341,In_1186,In_2356);
nand U1342 (N_1342,In_1820,In_1120);
nand U1343 (N_1343,In_851,In_1591);
xnor U1344 (N_1344,In_1517,In_2350);
or U1345 (N_1345,In_1837,In_2052);
or U1346 (N_1346,In_2162,In_1264);
xor U1347 (N_1347,In_1351,In_930);
and U1348 (N_1348,In_346,In_2037);
and U1349 (N_1349,In_1453,In_2048);
and U1350 (N_1350,In_32,In_2311);
nor U1351 (N_1351,In_163,In_1311);
and U1352 (N_1352,In_1203,In_2005);
nor U1353 (N_1353,In_688,In_1030);
and U1354 (N_1354,In_1137,In_1976);
or U1355 (N_1355,In_1606,In_327);
and U1356 (N_1356,In_89,In_1884);
or U1357 (N_1357,In_1083,In_1033);
and U1358 (N_1358,In_1637,In_789);
xnor U1359 (N_1359,In_663,In_513);
or U1360 (N_1360,In_2276,In_1194);
nand U1361 (N_1361,In_2253,In_8);
nor U1362 (N_1362,In_262,In_2062);
xnor U1363 (N_1363,In_2397,In_2216);
and U1364 (N_1364,In_444,In_808);
nand U1365 (N_1365,In_1298,In_597);
xnor U1366 (N_1366,In_1319,In_2338);
nor U1367 (N_1367,In_1502,In_223);
and U1368 (N_1368,In_1886,In_1129);
nor U1369 (N_1369,In_2203,In_716);
nor U1370 (N_1370,In_195,In_593);
or U1371 (N_1371,In_675,In_527);
and U1372 (N_1372,In_206,In_2074);
and U1373 (N_1373,In_1106,In_1891);
or U1374 (N_1374,In_76,In_247);
nand U1375 (N_1375,In_409,In_189);
xor U1376 (N_1376,In_2178,In_1351);
and U1377 (N_1377,In_1167,In_1771);
and U1378 (N_1378,In_883,In_2244);
nand U1379 (N_1379,In_2359,In_502);
nor U1380 (N_1380,In_1490,In_1484);
nor U1381 (N_1381,In_2406,In_2420);
xor U1382 (N_1382,In_2141,In_1717);
or U1383 (N_1383,In_2014,In_1509);
and U1384 (N_1384,In_2199,In_1389);
or U1385 (N_1385,In_68,In_59);
nand U1386 (N_1386,In_1679,In_393);
nor U1387 (N_1387,In_1288,In_1255);
xor U1388 (N_1388,In_956,In_1424);
nand U1389 (N_1389,In_159,In_342);
nor U1390 (N_1390,In_113,In_1240);
and U1391 (N_1391,In_192,In_1014);
or U1392 (N_1392,In_2228,In_1261);
and U1393 (N_1393,In_1768,In_1328);
or U1394 (N_1394,In_1024,In_2466);
nor U1395 (N_1395,In_1676,In_1210);
nor U1396 (N_1396,In_1597,In_949);
or U1397 (N_1397,In_507,In_1092);
nor U1398 (N_1398,In_125,In_1447);
xor U1399 (N_1399,In_1603,In_2167);
or U1400 (N_1400,In_509,In_2264);
nor U1401 (N_1401,In_357,In_14);
nor U1402 (N_1402,In_1153,In_399);
nand U1403 (N_1403,In_1599,In_2334);
xor U1404 (N_1404,In_2231,In_772);
nor U1405 (N_1405,In_617,In_1768);
nor U1406 (N_1406,In_519,In_1085);
nand U1407 (N_1407,In_2211,In_1520);
nor U1408 (N_1408,In_1481,In_2298);
nand U1409 (N_1409,In_2177,In_1925);
or U1410 (N_1410,In_1556,In_574);
nor U1411 (N_1411,In_2245,In_2261);
and U1412 (N_1412,In_2344,In_176);
or U1413 (N_1413,In_782,In_1811);
nand U1414 (N_1414,In_1013,In_1659);
or U1415 (N_1415,In_619,In_1071);
nand U1416 (N_1416,In_1311,In_316);
nand U1417 (N_1417,In_398,In_1930);
xnor U1418 (N_1418,In_643,In_579);
xnor U1419 (N_1419,In_1860,In_553);
xnor U1420 (N_1420,In_66,In_1218);
nor U1421 (N_1421,In_1700,In_1816);
nand U1422 (N_1422,In_1490,In_594);
nand U1423 (N_1423,In_1873,In_47);
nor U1424 (N_1424,In_109,In_1010);
nor U1425 (N_1425,In_2217,In_190);
and U1426 (N_1426,In_388,In_1853);
nor U1427 (N_1427,In_2216,In_1860);
and U1428 (N_1428,In_838,In_1623);
nor U1429 (N_1429,In_2478,In_2268);
xor U1430 (N_1430,In_2319,In_737);
or U1431 (N_1431,In_237,In_2022);
nor U1432 (N_1432,In_433,In_2468);
or U1433 (N_1433,In_1759,In_899);
and U1434 (N_1434,In_861,In_556);
xnor U1435 (N_1435,In_879,In_600);
nor U1436 (N_1436,In_1901,In_1842);
or U1437 (N_1437,In_2061,In_1396);
or U1438 (N_1438,In_2256,In_2001);
or U1439 (N_1439,In_653,In_1341);
and U1440 (N_1440,In_1506,In_1520);
xor U1441 (N_1441,In_1274,In_2349);
or U1442 (N_1442,In_551,In_772);
xor U1443 (N_1443,In_1838,In_151);
xor U1444 (N_1444,In_2318,In_1324);
nand U1445 (N_1445,In_124,In_1596);
nor U1446 (N_1446,In_529,In_637);
nor U1447 (N_1447,In_154,In_1863);
or U1448 (N_1448,In_274,In_228);
and U1449 (N_1449,In_1449,In_294);
or U1450 (N_1450,In_1193,In_2455);
or U1451 (N_1451,In_1915,In_2316);
nor U1452 (N_1452,In_1294,In_1370);
xor U1453 (N_1453,In_1069,In_1306);
nor U1454 (N_1454,In_1051,In_1433);
nor U1455 (N_1455,In_1267,In_840);
or U1456 (N_1456,In_1811,In_891);
and U1457 (N_1457,In_1257,In_419);
nand U1458 (N_1458,In_1322,In_2492);
nand U1459 (N_1459,In_1213,In_969);
nand U1460 (N_1460,In_640,In_1443);
nand U1461 (N_1461,In_1528,In_1360);
and U1462 (N_1462,In_598,In_262);
xnor U1463 (N_1463,In_341,In_1199);
xnor U1464 (N_1464,In_1884,In_1408);
nor U1465 (N_1465,In_197,In_520);
nor U1466 (N_1466,In_0,In_2369);
nand U1467 (N_1467,In_545,In_2312);
and U1468 (N_1468,In_2426,In_691);
nor U1469 (N_1469,In_474,In_2244);
or U1470 (N_1470,In_988,In_1078);
nor U1471 (N_1471,In_468,In_552);
xor U1472 (N_1472,In_1371,In_7);
xor U1473 (N_1473,In_2327,In_1736);
and U1474 (N_1474,In_423,In_2176);
nand U1475 (N_1475,In_2352,In_265);
or U1476 (N_1476,In_396,In_805);
xor U1477 (N_1477,In_808,In_1833);
xnor U1478 (N_1478,In_533,In_2394);
and U1479 (N_1479,In_681,In_2241);
or U1480 (N_1480,In_2387,In_1647);
nor U1481 (N_1481,In_602,In_738);
nand U1482 (N_1482,In_1852,In_1310);
nand U1483 (N_1483,In_2026,In_972);
xnor U1484 (N_1484,In_1730,In_1832);
or U1485 (N_1485,In_1568,In_507);
nand U1486 (N_1486,In_1626,In_97);
xnor U1487 (N_1487,In_36,In_2401);
xnor U1488 (N_1488,In_967,In_194);
nand U1489 (N_1489,In_2064,In_1128);
xor U1490 (N_1490,In_769,In_152);
nor U1491 (N_1491,In_1878,In_2299);
xnor U1492 (N_1492,In_975,In_1279);
nand U1493 (N_1493,In_812,In_1615);
nand U1494 (N_1494,In_1217,In_2154);
nand U1495 (N_1495,In_592,In_134);
and U1496 (N_1496,In_206,In_106);
nor U1497 (N_1497,In_2498,In_835);
nor U1498 (N_1498,In_702,In_19);
xor U1499 (N_1499,In_2371,In_1404);
and U1500 (N_1500,In_1725,In_2475);
xor U1501 (N_1501,In_530,In_822);
xor U1502 (N_1502,In_2352,In_2030);
nand U1503 (N_1503,In_2015,In_704);
and U1504 (N_1504,In_42,In_2138);
xor U1505 (N_1505,In_2446,In_1297);
xor U1506 (N_1506,In_1779,In_2447);
or U1507 (N_1507,In_2005,In_988);
or U1508 (N_1508,In_2075,In_150);
nand U1509 (N_1509,In_1030,In_2019);
and U1510 (N_1510,In_1361,In_1675);
nor U1511 (N_1511,In_1107,In_736);
nor U1512 (N_1512,In_2014,In_1968);
nor U1513 (N_1513,In_2032,In_1597);
or U1514 (N_1514,In_1866,In_1229);
nand U1515 (N_1515,In_304,In_755);
nor U1516 (N_1516,In_607,In_1845);
xor U1517 (N_1517,In_1499,In_855);
xnor U1518 (N_1518,In_2101,In_1287);
or U1519 (N_1519,In_854,In_945);
and U1520 (N_1520,In_2251,In_526);
nand U1521 (N_1521,In_27,In_404);
xor U1522 (N_1522,In_1989,In_729);
and U1523 (N_1523,In_2188,In_1159);
nor U1524 (N_1524,In_2213,In_1387);
and U1525 (N_1525,In_2499,In_1843);
nand U1526 (N_1526,In_2246,In_55);
nand U1527 (N_1527,In_298,In_1052);
and U1528 (N_1528,In_525,In_2361);
and U1529 (N_1529,In_513,In_767);
or U1530 (N_1530,In_2072,In_1536);
nor U1531 (N_1531,In_423,In_1025);
nor U1532 (N_1532,In_1229,In_1440);
and U1533 (N_1533,In_1634,In_764);
xor U1534 (N_1534,In_2048,In_1400);
nor U1535 (N_1535,In_877,In_1263);
xnor U1536 (N_1536,In_2313,In_2497);
or U1537 (N_1537,In_341,In_1942);
xnor U1538 (N_1538,In_319,In_1620);
and U1539 (N_1539,In_1322,In_1309);
and U1540 (N_1540,In_5,In_953);
and U1541 (N_1541,In_2245,In_1989);
and U1542 (N_1542,In_2369,In_2236);
and U1543 (N_1543,In_1432,In_2098);
nand U1544 (N_1544,In_820,In_304);
nor U1545 (N_1545,In_1084,In_1115);
xnor U1546 (N_1546,In_17,In_1651);
xor U1547 (N_1547,In_75,In_270);
or U1548 (N_1548,In_1079,In_2153);
xor U1549 (N_1549,In_1371,In_616);
nand U1550 (N_1550,In_634,In_2010);
nor U1551 (N_1551,In_2386,In_676);
or U1552 (N_1552,In_2208,In_10);
nor U1553 (N_1553,In_2299,In_874);
nor U1554 (N_1554,In_921,In_1684);
nor U1555 (N_1555,In_1284,In_1160);
nand U1556 (N_1556,In_2301,In_428);
nor U1557 (N_1557,In_2047,In_1039);
nor U1558 (N_1558,In_253,In_2002);
nor U1559 (N_1559,In_337,In_756);
nand U1560 (N_1560,In_1558,In_828);
nor U1561 (N_1561,In_77,In_159);
nand U1562 (N_1562,In_971,In_2241);
or U1563 (N_1563,In_1674,In_1954);
nor U1564 (N_1564,In_537,In_1292);
nor U1565 (N_1565,In_381,In_623);
xnor U1566 (N_1566,In_2423,In_239);
and U1567 (N_1567,In_56,In_163);
nand U1568 (N_1568,In_765,In_2217);
or U1569 (N_1569,In_2452,In_2313);
and U1570 (N_1570,In_1263,In_1567);
nand U1571 (N_1571,In_814,In_1757);
nor U1572 (N_1572,In_607,In_2371);
or U1573 (N_1573,In_1800,In_1958);
nand U1574 (N_1574,In_1353,In_2360);
nand U1575 (N_1575,In_261,In_136);
nor U1576 (N_1576,In_829,In_1737);
nor U1577 (N_1577,In_1457,In_1355);
nand U1578 (N_1578,In_2189,In_913);
xnor U1579 (N_1579,In_683,In_1226);
and U1580 (N_1580,In_902,In_1665);
nand U1581 (N_1581,In_173,In_2233);
nor U1582 (N_1582,In_1047,In_1469);
or U1583 (N_1583,In_134,In_460);
xor U1584 (N_1584,In_980,In_1421);
nand U1585 (N_1585,In_1359,In_72);
or U1586 (N_1586,In_2336,In_11);
nor U1587 (N_1587,In_2287,In_1089);
nor U1588 (N_1588,In_837,In_845);
nor U1589 (N_1589,In_2009,In_1627);
nand U1590 (N_1590,In_610,In_693);
or U1591 (N_1591,In_1736,In_253);
and U1592 (N_1592,In_1322,In_267);
nor U1593 (N_1593,In_1926,In_2018);
or U1594 (N_1594,In_374,In_8);
nor U1595 (N_1595,In_236,In_1487);
nor U1596 (N_1596,In_2242,In_1773);
nor U1597 (N_1597,In_22,In_2036);
xnor U1598 (N_1598,In_413,In_2484);
nand U1599 (N_1599,In_2331,In_1472);
nor U1600 (N_1600,In_1099,In_345);
and U1601 (N_1601,In_637,In_877);
nor U1602 (N_1602,In_883,In_2273);
xnor U1603 (N_1603,In_2173,In_2442);
or U1604 (N_1604,In_1630,In_497);
or U1605 (N_1605,In_901,In_1467);
and U1606 (N_1606,In_828,In_2369);
or U1607 (N_1607,In_2410,In_42);
and U1608 (N_1608,In_360,In_1240);
nand U1609 (N_1609,In_1827,In_709);
nor U1610 (N_1610,In_707,In_1001);
or U1611 (N_1611,In_1736,In_2220);
xor U1612 (N_1612,In_1472,In_613);
or U1613 (N_1613,In_276,In_383);
or U1614 (N_1614,In_136,In_403);
and U1615 (N_1615,In_222,In_1221);
xnor U1616 (N_1616,In_2181,In_1614);
nand U1617 (N_1617,In_60,In_1078);
nand U1618 (N_1618,In_936,In_850);
and U1619 (N_1619,In_1236,In_82);
xor U1620 (N_1620,In_599,In_2345);
nor U1621 (N_1621,In_931,In_2291);
and U1622 (N_1622,In_1569,In_180);
xor U1623 (N_1623,In_2476,In_1039);
nand U1624 (N_1624,In_55,In_1373);
and U1625 (N_1625,In_1244,In_1618);
or U1626 (N_1626,In_1796,In_1907);
nor U1627 (N_1627,In_1077,In_1129);
nor U1628 (N_1628,In_778,In_2177);
or U1629 (N_1629,In_136,In_282);
nor U1630 (N_1630,In_1876,In_2293);
and U1631 (N_1631,In_1387,In_1546);
nor U1632 (N_1632,In_957,In_2481);
xor U1633 (N_1633,In_1901,In_653);
and U1634 (N_1634,In_1838,In_1539);
and U1635 (N_1635,In_978,In_1304);
and U1636 (N_1636,In_2403,In_1950);
or U1637 (N_1637,In_1062,In_1984);
nor U1638 (N_1638,In_574,In_1205);
and U1639 (N_1639,In_2250,In_74);
nor U1640 (N_1640,In_1871,In_1075);
xnor U1641 (N_1641,In_2085,In_1916);
or U1642 (N_1642,In_472,In_1050);
nor U1643 (N_1643,In_155,In_923);
nand U1644 (N_1644,In_2414,In_1489);
or U1645 (N_1645,In_373,In_881);
nand U1646 (N_1646,In_1696,In_234);
xor U1647 (N_1647,In_2411,In_144);
and U1648 (N_1648,In_771,In_1271);
or U1649 (N_1649,In_1328,In_702);
nor U1650 (N_1650,In_2210,In_1051);
nand U1651 (N_1651,In_602,In_540);
or U1652 (N_1652,In_1331,In_799);
nor U1653 (N_1653,In_993,In_1523);
and U1654 (N_1654,In_1670,In_223);
and U1655 (N_1655,In_2302,In_820);
or U1656 (N_1656,In_1903,In_1602);
nand U1657 (N_1657,In_2059,In_1470);
nor U1658 (N_1658,In_1253,In_571);
or U1659 (N_1659,In_95,In_1044);
and U1660 (N_1660,In_89,In_1205);
xnor U1661 (N_1661,In_2178,In_2033);
xor U1662 (N_1662,In_692,In_860);
and U1663 (N_1663,In_820,In_1931);
nand U1664 (N_1664,In_972,In_1696);
nor U1665 (N_1665,In_388,In_833);
and U1666 (N_1666,In_683,In_151);
or U1667 (N_1667,In_1671,In_1397);
and U1668 (N_1668,In_175,In_898);
nor U1669 (N_1669,In_1136,In_656);
xor U1670 (N_1670,In_1466,In_1040);
nand U1671 (N_1671,In_340,In_334);
and U1672 (N_1672,In_1676,In_979);
nand U1673 (N_1673,In_2142,In_1617);
or U1674 (N_1674,In_778,In_697);
xor U1675 (N_1675,In_1775,In_1396);
nor U1676 (N_1676,In_2070,In_1573);
or U1677 (N_1677,In_333,In_274);
or U1678 (N_1678,In_404,In_1055);
nand U1679 (N_1679,In_1507,In_323);
xor U1680 (N_1680,In_1411,In_2080);
or U1681 (N_1681,In_76,In_2122);
xor U1682 (N_1682,In_431,In_2163);
and U1683 (N_1683,In_1593,In_1206);
nand U1684 (N_1684,In_1664,In_1052);
and U1685 (N_1685,In_1115,In_529);
xor U1686 (N_1686,In_2171,In_2499);
nor U1687 (N_1687,In_1621,In_1839);
and U1688 (N_1688,In_1965,In_893);
nand U1689 (N_1689,In_107,In_2426);
nor U1690 (N_1690,In_337,In_2185);
xnor U1691 (N_1691,In_1458,In_480);
or U1692 (N_1692,In_1582,In_28);
xor U1693 (N_1693,In_112,In_662);
and U1694 (N_1694,In_1475,In_308);
nor U1695 (N_1695,In_102,In_537);
or U1696 (N_1696,In_1089,In_791);
or U1697 (N_1697,In_481,In_1029);
nand U1698 (N_1698,In_650,In_1405);
xnor U1699 (N_1699,In_1162,In_1447);
nand U1700 (N_1700,In_1592,In_2250);
nor U1701 (N_1701,In_1985,In_554);
and U1702 (N_1702,In_316,In_17);
nand U1703 (N_1703,In_1964,In_1124);
or U1704 (N_1704,In_731,In_2070);
nor U1705 (N_1705,In_314,In_2241);
xor U1706 (N_1706,In_2336,In_1885);
nor U1707 (N_1707,In_605,In_570);
and U1708 (N_1708,In_1148,In_724);
xor U1709 (N_1709,In_1651,In_1406);
and U1710 (N_1710,In_1294,In_271);
or U1711 (N_1711,In_1302,In_506);
nor U1712 (N_1712,In_2291,In_1575);
nand U1713 (N_1713,In_866,In_2);
nor U1714 (N_1714,In_1788,In_761);
nand U1715 (N_1715,In_2226,In_125);
nor U1716 (N_1716,In_1915,In_1113);
xor U1717 (N_1717,In_2222,In_1593);
nor U1718 (N_1718,In_921,In_985);
xnor U1719 (N_1719,In_1707,In_1581);
xnor U1720 (N_1720,In_2068,In_1455);
nand U1721 (N_1721,In_2137,In_613);
or U1722 (N_1722,In_1754,In_1921);
nand U1723 (N_1723,In_1551,In_2066);
nand U1724 (N_1724,In_739,In_2408);
nor U1725 (N_1725,In_48,In_682);
nand U1726 (N_1726,In_2055,In_773);
or U1727 (N_1727,In_1489,In_343);
nor U1728 (N_1728,In_230,In_1363);
or U1729 (N_1729,In_2013,In_2217);
and U1730 (N_1730,In_2009,In_411);
or U1731 (N_1731,In_107,In_551);
and U1732 (N_1732,In_1794,In_603);
nand U1733 (N_1733,In_586,In_7);
or U1734 (N_1734,In_1203,In_568);
nor U1735 (N_1735,In_499,In_804);
xor U1736 (N_1736,In_2123,In_1160);
nand U1737 (N_1737,In_346,In_921);
xnor U1738 (N_1738,In_897,In_188);
nor U1739 (N_1739,In_1577,In_140);
xor U1740 (N_1740,In_634,In_1664);
xnor U1741 (N_1741,In_1984,In_1130);
nor U1742 (N_1742,In_1066,In_182);
nor U1743 (N_1743,In_1986,In_2046);
and U1744 (N_1744,In_857,In_1147);
and U1745 (N_1745,In_1,In_863);
nor U1746 (N_1746,In_350,In_456);
nand U1747 (N_1747,In_584,In_1270);
nand U1748 (N_1748,In_106,In_357);
or U1749 (N_1749,In_228,In_902);
xor U1750 (N_1750,In_2278,In_614);
xnor U1751 (N_1751,In_761,In_1686);
nor U1752 (N_1752,In_2351,In_1557);
nand U1753 (N_1753,In_177,In_1445);
or U1754 (N_1754,In_2292,In_794);
xor U1755 (N_1755,In_342,In_2473);
and U1756 (N_1756,In_1360,In_1603);
xnor U1757 (N_1757,In_2296,In_1928);
or U1758 (N_1758,In_917,In_841);
nand U1759 (N_1759,In_1718,In_1132);
or U1760 (N_1760,In_2324,In_478);
nand U1761 (N_1761,In_2262,In_1185);
and U1762 (N_1762,In_1941,In_1683);
nor U1763 (N_1763,In_1241,In_1785);
and U1764 (N_1764,In_1149,In_1800);
xor U1765 (N_1765,In_32,In_1276);
nor U1766 (N_1766,In_913,In_1050);
and U1767 (N_1767,In_403,In_525);
and U1768 (N_1768,In_222,In_821);
or U1769 (N_1769,In_780,In_471);
or U1770 (N_1770,In_1187,In_1410);
xor U1771 (N_1771,In_782,In_270);
and U1772 (N_1772,In_837,In_2403);
nor U1773 (N_1773,In_800,In_765);
nor U1774 (N_1774,In_2044,In_819);
xor U1775 (N_1775,In_2320,In_770);
and U1776 (N_1776,In_1096,In_2457);
xor U1777 (N_1777,In_683,In_1337);
nor U1778 (N_1778,In_734,In_1370);
nand U1779 (N_1779,In_419,In_2399);
and U1780 (N_1780,In_608,In_393);
or U1781 (N_1781,In_1273,In_788);
nand U1782 (N_1782,In_659,In_1909);
xor U1783 (N_1783,In_753,In_1273);
nand U1784 (N_1784,In_900,In_2251);
xnor U1785 (N_1785,In_1970,In_2057);
nand U1786 (N_1786,In_1613,In_1796);
nor U1787 (N_1787,In_2225,In_191);
and U1788 (N_1788,In_1642,In_1595);
xor U1789 (N_1789,In_541,In_694);
xnor U1790 (N_1790,In_41,In_1414);
and U1791 (N_1791,In_532,In_979);
nand U1792 (N_1792,In_2011,In_2474);
nand U1793 (N_1793,In_1248,In_1685);
xor U1794 (N_1794,In_466,In_1112);
nor U1795 (N_1795,In_797,In_2344);
and U1796 (N_1796,In_1673,In_500);
and U1797 (N_1797,In_94,In_1207);
and U1798 (N_1798,In_1779,In_2088);
nor U1799 (N_1799,In_1773,In_1135);
xor U1800 (N_1800,In_148,In_1348);
nand U1801 (N_1801,In_216,In_1988);
nand U1802 (N_1802,In_29,In_2002);
xnor U1803 (N_1803,In_1588,In_629);
nor U1804 (N_1804,In_277,In_2136);
nor U1805 (N_1805,In_2017,In_1667);
and U1806 (N_1806,In_1960,In_20);
xnor U1807 (N_1807,In_1883,In_1474);
xor U1808 (N_1808,In_1827,In_918);
or U1809 (N_1809,In_281,In_1989);
nand U1810 (N_1810,In_696,In_634);
and U1811 (N_1811,In_1149,In_138);
nand U1812 (N_1812,In_864,In_1870);
xor U1813 (N_1813,In_231,In_2049);
xor U1814 (N_1814,In_43,In_721);
and U1815 (N_1815,In_1467,In_586);
and U1816 (N_1816,In_660,In_830);
or U1817 (N_1817,In_692,In_455);
nand U1818 (N_1818,In_1174,In_2228);
nor U1819 (N_1819,In_801,In_910);
nand U1820 (N_1820,In_1134,In_283);
and U1821 (N_1821,In_626,In_2165);
or U1822 (N_1822,In_579,In_702);
xnor U1823 (N_1823,In_456,In_0);
or U1824 (N_1824,In_891,In_1575);
or U1825 (N_1825,In_593,In_833);
xnor U1826 (N_1826,In_2353,In_1839);
xnor U1827 (N_1827,In_2199,In_2297);
and U1828 (N_1828,In_573,In_1328);
or U1829 (N_1829,In_430,In_2227);
nand U1830 (N_1830,In_129,In_425);
xor U1831 (N_1831,In_981,In_1699);
or U1832 (N_1832,In_246,In_1376);
xnor U1833 (N_1833,In_1752,In_317);
nor U1834 (N_1834,In_1994,In_1930);
xnor U1835 (N_1835,In_2101,In_1737);
nand U1836 (N_1836,In_1824,In_2418);
nor U1837 (N_1837,In_1439,In_684);
or U1838 (N_1838,In_1103,In_1844);
xor U1839 (N_1839,In_434,In_2154);
xor U1840 (N_1840,In_1641,In_54);
xor U1841 (N_1841,In_87,In_1469);
nand U1842 (N_1842,In_399,In_1382);
and U1843 (N_1843,In_593,In_1854);
nor U1844 (N_1844,In_1736,In_1808);
or U1845 (N_1845,In_1100,In_549);
and U1846 (N_1846,In_1270,In_2049);
and U1847 (N_1847,In_809,In_1194);
and U1848 (N_1848,In_2352,In_988);
xor U1849 (N_1849,In_1242,In_2013);
or U1850 (N_1850,In_1318,In_2053);
or U1851 (N_1851,In_84,In_372);
nand U1852 (N_1852,In_1090,In_1348);
xor U1853 (N_1853,In_720,In_1416);
nand U1854 (N_1854,In_2389,In_1712);
or U1855 (N_1855,In_1234,In_1214);
or U1856 (N_1856,In_432,In_951);
or U1857 (N_1857,In_2157,In_1738);
xnor U1858 (N_1858,In_765,In_986);
and U1859 (N_1859,In_2352,In_838);
nand U1860 (N_1860,In_611,In_2229);
nor U1861 (N_1861,In_311,In_2099);
nor U1862 (N_1862,In_389,In_1145);
xor U1863 (N_1863,In_255,In_2037);
nand U1864 (N_1864,In_1668,In_56);
and U1865 (N_1865,In_2365,In_974);
nor U1866 (N_1866,In_147,In_1326);
nor U1867 (N_1867,In_857,In_543);
nand U1868 (N_1868,In_669,In_1390);
or U1869 (N_1869,In_2419,In_2273);
xnor U1870 (N_1870,In_1136,In_1124);
xor U1871 (N_1871,In_2178,In_704);
nor U1872 (N_1872,In_1823,In_471);
nor U1873 (N_1873,In_688,In_1657);
and U1874 (N_1874,In_1619,In_547);
xnor U1875 (N_1875,In_2384,In_1785);
nor U1876 (N_1876,In_2116,In_277);
and U1877 (N_1877,In_872,In_2450);
or U1878 (N_1878,In_1973,In_1704);
or U1879 (N_1879,In_1771,In_568);
xnor U1880 (N_1880,In_273,In_859);
nor U1881 (N_1881,In_105,In_970);
nand U1882 (N_1882,In_628,In_828);
xnor U1883 (N_1883,In_2094,In_1856);
and U1884 (N_1884,In_2411,In_1567);
xnor U1885 (N_1885,In_1695,In_1951);
nor U1886 (N_1886,In_449,In_997);
or U1887 (N_1887,In_1161,In_1441);
xnor U1888 (N_1888,In_142,In_1584);
nor U1889 (N_1889,In_1644,In_477);
xor U1890 (N_1890,In_1887,In_586);
xnor U1891 (N_1891,In_2083,In_2101);
xnor U1892 (N_1892,In_2011,In_1186);
xor U1893 (N_1893,In_583,In_1958);
and U1894 (N_1894,In_905,In_2143);
xnor U1895 (N_1895,In_272,In_2224);
and U1896 (N_1896,In_900,In_2058);
xnor U1897 (N_1897,In_1971,In_281);
and U1898 (N_1898,In_93,In_1484);
xnor U1899 (N_1899,In_1910,In_152);
xnor U1900 (N_1900,In_653,In_1090);
or U1901 (N_1901,In_1876,In_2070);
xnor U1902 (N_1902,In_868,In_567);
nor U1903 (N_1903,In_1840,In_2046);
xor U1904 (N_1904,In_104,In_1462);
nand U1905 (N_1905,In_25,In_334);
nor U1906 (N_1906,In_1730,In_1333);
or U1907 (N_1907,In_149,In_1298);
and U1908 (N_1908,In_14,In_620);
or U1909 (N_1909,In_1222,In_523);
nor U1910 (N_1910,In_2215,In_1274);
nand U1911 (N_1911,In_1984,In_2129);
and U1912 (N_1912,In_1367,In_681);
nor U1913 (N_1913,In_1931,In_147);
nand U1914 (N_1914,In_2303,In_1848);
nand U1915 (N_1915,In_1261,In_247);
or U1916 (N_1916,In_798,In_783);
or U1917 (N_1917,In_1823,In_961);
or U1918 (N_1918,In_1791,In_1952);
nand U1919 (N_1919,In_785,In_2217);
or U1920 (N_1920,In_1557,In_1912);
nand U1921 (N_1921,In_589,In_1812);
nand U1922 (N_1922,In_1188,In_2235);
and U1923 (N_1923,In_930,In_1729);
and U1924 (N_1924,In_2469,In_421);
or U1925 (N_1925,In_275,In_2132);
nand U1926 (N_1926,In_1672,In_446);
nand U1927 (N_1927,In_1294,In_724);
nor U1928 (N_1928,In_2422,In_1739);
nor U1929 (N_1929,In_456,In_1946);
or U1930 (N_1930,In_2138,In_1325);
xnor U1931 (N_1931,In_2095,In_1631);
and U1932 (N_1932,In_265,In_1343);
or U1933 (N_1933,In_1709,In_1921);
or U1934 (N_1934,In_1289,In_677);
and U1935 (N_1935,In_2148,In_1984);
nor U1936 (N_1936,In_92,In_779);
nor U1937 (N_1937,In_746,In_2111);
or U1938 (N_1938,In_1358,In_47);
and U1939 (N_1939,In_190,In_1899);
and U1940 (N_1940,In_2442,In_673);
xor U1941 (N_1941,In_1458,In_1950);
or U1942 (N_1942,In_1911,In_284);
nor U1943 (N_1943,In_1216,In_2162);
and U1944 (N_1944,In_1427,In_319);
or U1945 (N_1945,In_1578,In_1878);
xnor U1946 (N_1946,In_1253,In_794);
or U1947 (N_1947,In_2392,In_399);
and U1948 (N_1948,In_1522,In_1350);
nand U1949 (N_1949,In_2195,In_1095);
nor U1950 (N_1950,In_2473,In_1124);
and U1951 (N_1951,In_1254,In_614);
or U1952 (N_1952,In_1282,In_729);
nand U1953 (N_1953,In_2141,In_1719);
or U1954 (N_1954,In_739,In_445);
nand U1955 (N_1955,In_710,In_2053);
nand U1956 (N_1956,In_217,In_444);
xor U1957 (N_1957,In_1258,In_1105);
nor U1958 (N_1958,In_1194,In_754);
nand U1959 (N_1959,In_1603,In_918);
or U1960 (N_1960,In_588,In_1894);
or U1961 (N_1961,In_952,In_62);
nor U1962 (N_1962,In_2055,In_144);
nand U1963 (N_1963,In_1830,In_132);
xnor U1964 (N_1964,In_1780,In_363);
or U1965 (N_1965,In_1315,In_2440);
or U1966 (N_1966,In_1595,In_1212);
xor U1967 (N_1967,In_845,In_209);
xnor U1968 (N_1968,In_448,In_2140);
xor U1969 (N_1969,In_2398,In_1819);
nor U1970 (N_1970,In_587,In_285);
nand U1971 (N_1971,In_2172,In_880);
xnor U1972 (N_1972,In_428,In_327);
nor U1973 (N_1973,In_1168,In_1601);
nor U1974 (N_1974,In_760,In_910);
or U1975 (N_1975,In_2033,In_137);
nor U1976 (N_1976,In_1709,In_2347);
xor U1977 (N_1977,In_94,In_2042);
and U1978 (N_1978,In_364,In_2061);
nand U1979 (N_1979,In_1891,In_1098);
or U1980 (N_1980,In_954,In_311);
nor U1981 (N_1981,In_2299,In_1854);
nand U1982 (N_1982,In_270,In_1890);
nor U1983 (N_1983,In_2129,In_1491);
or U1984 (N_1984,In_1766,In_1926);
or U1985 (N_1985,In_2399,In_1546);
and U1986 (N_1986,In_1113,In_697);
and U1987 (N_1987,In_551,In_1260);
or U1988 (N_1988,In_169,In_2195);
and U1989 (N_1989,In_1288,In_1741);
and U1990 (N_1990,In_2352,In_1908);
and U1991 (N_1991,In_484,In_1307);
or U1992 (N_1992,In_1736,In_2421);
nor U1993 (N_1993,In_896,In_1999);
nand U1994 (N_1994,In_134,In_1486);
nand U1995 (N_1995,In_576,In_1722);
nor U1996 (N_1996,In_2296,In_1522);
nand U1997 (N_1997,In_1232,In_483);
xor U1998 (N_1998,In_1937,In_364);
nor U1999 (N_1999,In_1612,In_1627);
or U2000 (N_2000,In_220,In_2238);
xnor U2001 (N_2001,In_2462,In_152);
and U2002 (N_2002,In_1974,In_409);
or U2003 (N_2003,In_838,In_985);
and U2004 (N_2004,In_2434,In_967);
and U2005 (N_2005,In_1079,In_1716);
nand U2006 (N_2006,In_1700,In_1300);
xnor U2007 (N_2007,In_1968,In_71);
nor U2008 (N_2008,In_287,In_1756);
xor U2009 (N_2009,In_1507,In_838);
xor U2010 (N_2010,In_1189,In_1631);
xor U2011 (N_2011,In_195,In_1226);
nand U2012 (N_2012,In_959,In_720);
or U2013 (N_2013,In_1044,In_1086);
nand U2014 (N_2014,In_357,In_112);
xor U2015 (N_2015,In_872,In_2380);
nand U2016 (N_2016,In_298,In_2422);
or U2017 (N_2017,In_1064,In_2293);
xnor U2018 (N_2018,In_967,In_673);
and U2019 (N_2019,In_979,In_882);
and U2020 (N_2020,In_142,In_1912);
xor U2021 (N_2021,In_1277,In_951);
and U2022 (N_2022,In_1554,In_2265);
and U2023 (N_2023,In_1057,In_183);
xnor U2024 (N_2024,In_1655,In_1759);
nand U2025 (N_2025,In_1116,In_1404);
nand U2026 (N_2026,In_2393,In_1418);
xnor U2027 (N_2027,In_997,In_1861);
and U2028 (N_2028,In_573,In_1702);
nor U2029 (N_2029,In_188,In_275);
nor U2030 (N_2030,In_1980,In_283);
xor U2031 (N_2031,In_348,In_1742);
nor U2032 (N_2032,In_1527,In_1617);
nor U2033 (N_2033,In_1378,In_734);
xnor U2034 (N_2034,In_1799,In_704);
xor U2035 (N_2035,In_1988,In_1635);
xor U2036 (N_2036,In_1812,In_2299);
nor U2037 (N_2037,In_1184,In_811);
nand U2038 (N_2038,In_1035,In_771);
nor U2039 (N_2039,In_1280,In_2295);
and U2040 (N_2040,In_886,In_1319);
nor U2041 (N_2041,In_1178,In_683);
and U2042 (N_2042,In_2374,In_2442);
nand U2043 (N_2043,In_1367,In_1284);
xnor U2044 (N_2044,In_1342,In_235);
nor U2045 (N_2045,In_849,In_86);
nor U2046 (N_2046,In_1957,In_1592);
or U2047 (N_2047,In_1904,In_1719);
nand U2048 (N_2048,In_645,In_1065);
xor U2049 (N_2049,In_843,In_389);
nor U2050 (N_2050,In_344,In_767);
and U2051 (N_2051,In_2109,In_873);
nand U2052 (N_2052,In_815,In_1082);
xor U2053 (N_2053,In_1057,In_1734);
and U2054 (N_2054,In_1434,In_718);
nor U2055 (N_2055,In_1797,In_1869);
nor U2056 (N_2056,In_327,In_187);
and U2057 (N_2057,In_1717,In_872);
nor U2058 (N_2058,In_750,In_1144);
and U2059 (N_2059,In_1858,In_1028);
and U2060 (N_2060,In_786,In_1137);
or U2061 (N_2061,In_1252,In_58);
and U2062 (N_2062,In_380,In_952);
and U2063 (N_2063,In_1188,In_257);
or U2064 (N_2064,In_649,In_2257);
xnor U2065 (N_2065,In_1341,In_1643);
and U2066 (N_2066,In_2263,In_565);
xor U2067 (N_2067,In_820,In_2177);
or U2068 (N_2068,In_27,In_1876);
and U2069 (N_2069,In_2111,In_1708);
nor U2070 (N_2070,In_218,In_1201);
or U2071 (N_2071,In_821,In_2227);
or U2072 (N_2072,In_2329,In_2226);
xor U2073 (N_2073,In_1760,In_1649);
xor U2074 (N_2074,In_521,In_130);
nand U2075 (N_2075,In_1761,In_1949);
or U2076 (N_2076,In_738,In_902);
and U2077 (N_2077,In_65,In_1035);
xnor U2078 (N_2078,In_2487,In_1451);
or U2079 (N_2079,In_2098,In_897);
or U2080 (N_2080,In_966,In_2457);
xor U2081 (N_2081,In_2486,In_898);
nor U2082 (N_2082,In_638,In_2126);
nand U2083 (N_2083,In_2392,In_1617);
nor U2084 (N_2084,In_447,In_2352);
nand U2085 (N_2085,In_2311,In_795);
and U2086 (N_2086,In_1030,In_81);
nand U2087 (N_2087,In_1631,In_1717);
xnor U2088 (N_2088,In_2303,In_1104);
nand U2089 (N_2089,In_2138,In_454);
xnor U2090 (N_2090,In_574,In_796);
xnor U2091 (N_2091,In_1288,In_371);
and U2092 (N_2092,In_877,In_1876);
or U2093 (N_2093,In_2119,In_74);
nor U2094 (N_2094,In_835,In_1774);
nor U2095 (N_2095,In_1509,In_563);
nor U2096 (N_2096,In_856,In_1832);
or U2097 (N_2097,In_1754,In_1927);
nor U2098 (N_2098,In_140,In_829);
or U2099 (N_2099,In_2146,In_2247);
nor U2100 (N_2100,In_1432,In_1654);
or U2101 (N_2101,In_1507,In_1699);
and U2102 (N_2102,In_2011,In_66);
nand U2103 (N_2103,In_1804,In_1935);
nor U2104 (N_2104,In_2073,In_993);
nand U2105 (N_2105,In_610,In_692);
nor U2106 (N_2106,In_2368,In_1351);
xnor U2107 (N_2107,In_2106,In_60);
xnor U2108 (N_2108,In_346,In_1374);
xor U2109 (N_2109,In_1091,In_566);
or U2110 (N_2110,In_1217,In_654);
nand U2111 (N_2111,In_1829,In_2220);
or U2112 (N_2112,In_243,In_929);
xnor U2113 (N_2113,In_413,In_361);
nor U2114 (N_2114,In_33,In_955);
and U2115 (N_2115,In_2498,In_1788);
xor U2116 (N_2116,In_1762,In_111);
nand U2117 (N_2117,In_1752,In_1141);
or U2118 (N_2118,In_317,In_1804);
or U2119 (N_2119,In_607,In_1223);
nand U2120 (N_2120,In_1368,In_2052);
nand U2121 (N_2121,In_2099,In_1341);
and U2122 (N_2122,In_500,In_702);
nand U2123 (N_2123,In_1407,In_1306);
nor U2124 (N_2124,In_2287,In_375);
or U2125 (N_2125,In_1709,In_429);
nor U2126 (N_2126,In_182,In_266);
nand U2127 (N_2127,In_2235,In_1281);
or U2128 (N_2128,In_1415,In_2098);
or U2129 (N_2129,In_818,In_948);
or U2130 (N_2130,In_161,In_2374);
xor U2131 (N_2131,In_2314,In_2176);
and U2132 (N_2132,In_2214,In_58);
and U2133 (N_2133,In_1787,In_648);
nor U2134 (N_2134,In_1032,In_525);
nor U2135 (N_2135,In_234,In_2168);
and U2136 (N_2136,In_778,In_1557);
nor U2137 (N_2137,In_2194,In_1886);
or U2138 (N_2138,In_681,In_92);
or U2139 (N_2139,In_1713,In_48);
and U2140 (N_2140,In_2481,In_2033);
and U2141 (N_2141,In_2187,In_1806);
nor U2142 (N_2142,In_2240,In_1072);
xor U2143 (N_2143,In_1308,In_2210);
or U2144 (N_2144,In_216,In_1883);
nand U2145 (N_2145,In_704,In_933);
xor U2146 (N_2146,In_1387,In_1849);
xnor U2147 (N_2147,In_2291,In_493);
xnor U2148 (N_2148,In_522,In_503);
and U2149 (N_2149,In_1086,In_2318);
xor U2150 (N_2150,In_854,In_2001);
or U2151 (N_2151,In_2009,In_2132);
nand U2152 (N_2152,In_2351,In_2048);
xnor U2153 (N_2153,In_1644,In_1288);
nor U2154 (N_2154,In_541,In_617);
and U2155 (N_2155,In_259,In_1062);
nor U2156 (N_2156,In_893,In_166);
or U2157 (N_2157,In_1892,In_1008);
and U2158 (N_2158,In_2433,In_1860);
or U2159 (N_2159,In_1353,In_580);
nand U2160 (N_2160,In_471,In_1662);
or U2161 (N_2161,In_864,In_265);
and U2162 (N_2162,In_2358,In_918);
and U2163 (N_2163,In_2355,In_861);
nand U2164 (N_2164,In_1769,In_298);
or U2165 (N_2165,In_1856,In_2183);
xnor U2166 (N_2166,In_2295,In_1775);
or U2167 (N_2167,In_1071,In_2042);
nor U2168 (N_2168,In_814,In_874);
xor U2169 (N_2169,In_1620,In_447);
nor U2170 (N_2170,In_1534,In_1623);
and U2171 (N_2171,In_702,In_2430);
xor U2172 (N_2172,In_38,In_1635);
xnor U2173 (N_2173,In_199,In_413);
xor U2174 (N_2174,In_2178,In_841);
xnor U2175 (N_2175,In_2439,In_1962);
or U2176 (N_2176,In_342,In_264);
nor U2177 (N_2177,In_899,In_106);
nor U2178 (N_2178,In_812,In_1857);
nand U2179 (N_2179,In_2264,In_2422);
and U2180 (N_2180,In_533,In_766);
or U2181 (N_2181,In_1850,In_1922);
nor U2182 (N_2182,In_1189,In_1270);
nand U2183 (N_2183,In_2028,In_553);
xnor U2184 (N_2184,In_379,In_1727);
nand U2185 (N_2185,In_503,In_1777);
nor U2186 (N_2186,In_1805,In_2203);
and U2187 (N_2187,In_1441,In_1826);
or U2188 (N_2188,In_2486,In_749);
and U2189 (N_2189,In_342,In_511);
xor U2190 (N_2190,In_582,In_1243);
xor U2191 (N_2191,In_1612,In_2450);
or U2192 (N_2192,In_1170,In_827);
nor U2193 (N_2193,In_1128,In_1534);
nor U2194 (N_2194,In_553,In_1781);
or U2195 (N_2195,In_659,In_472);
xor U2196 (N_2196,In_2493,In_956);
or U2197 (N_2197,In_176,In_192);
and U2198 (N_2198,In_1118,In_1882);
xnor U2199 (N_2199,In_1018,In_1765);
nor U2200 (N_2200,In_784,In_76);
and U2201 (N_2201,In_697,In_364);
xnor U2202 (N_2202,In_405,In_539);
and U2203 (N_2203,In_3,In_627);
nand U2204 (N_2204,In_14,In_362);
and U2205 (N_2205,In_59,In_2147);
nor U2206 (N_2206,In_495,In_176);
and U2207 (N_2207,In_633,In_2132);
or U2208 (N_2208,In_24,In_2458);
and U2209 (N_2209,In_2465,In_2053);
nor U2210 (N_2210,In_785,In_936);
or U2211 (N_2211,In_667,In_1893);
nor U2212 (N_2212,In_579,In_67);
xnor U2213 (N_2213,In_2004,In_101);
xnor U2214 (N_2214,In_1116,In_2060);
nor U2215 (N_2215,In_2129,In_778);
nor U2216 (N_2216,In_323,In_2146);
or U2217 (N_2217,In_329,In_1391);
and U2218 (N_2218,In_724,In_2142);
xor U2219 (N_2219,In_862,In_180);
or U2220 (N_2220,In_523,In_1575);
nor U2221 (N_2221,In_316,In_1079);
nor U2222 (N_2222,In_1697,In_239);
xor U2223 (N_2223,In_2424,In_543);
nor U2224 (N_2224,In_1614,In_1300);
and U2225 (N_2225,In_2397,In_2000);
and U2226 (N_2226,In_986,In_2069);
or U2227 (N_2227,In_1103,In_1572);
xor U2228 (N_2228,In_2423,In_2155);
xnor U2229 (N_2229,In_1473,In_2386);
xnor U2230 (N_2230,In_1665,In_499);
and U2231 (N_2231,In_2315,In_333);
nand U2232 (N_2232,In_943,In_2256);
nor U2233 (N_2233,In_1239,In_1380);
and U2234 (N_2234,In_1320,In_2356);
nor U2235 (N_2235,In_3,In_851);
nor U2236 (N_2236,In_1818,In_383);
xor U2237 (N_2237,In_1691,In_1550);
or U2238 (N_2238,In_2136,In_1390);
nor U2239 (N_2239,In_61,In_1357);
and U2240 (N_2240,In_1076,In_693);
or U2241 (N_2241,In_2464,In_1849);
nand U2242 (N_2242,In_1428,In_2276);
or U2243 (N_2243,In_1940,In_1012);
nand U2244 (N_2244,In_1605,In_2127);
or U2245 (N_2245,In_680,In_1357);
xnor U2246 (N_2246,In_1014,In_677);
xor U2247 (N_2247,In_1218,In_2395);
xnor U2248 (N_2248,In_1179,In_1452);
and U2249 (N_2249,In_2190,In_2270);
and U2250 (N_2250,In_2085,In_1848);
nor U2251 (N_2251,In_1187,In_23);
xor U2252 (N_2252,In_2058,In_1742);
or U2253 (N_2253,In_1368,In_1011);
xor U2254 (N_2254,In_155,In_1769);
nor U2255 (N_2255,In_1292,In_351);
nor U2256 (N_2256,In_1868,In_639);
or U2257 (N_2257,In_877,In_943);
nor U2258 (N_2258,In_1951,In_2203);
or U2259 (N_2259,In_1035,In_2012);
nor U2260 (N_2260,In_488,In_1664);
and U2261 (N_2261,In_651,In_742);
and U2262 (N_2262,In_1503,In_210);
nor U2263 (N_2263,In_1377,In_650);
or U2264 (N_2264,In_425,In_2483);
nor U2265 (N_2265,In_627,In_623);
nor U2266 (N_2266,In_1060,In_1977);
or U2267 (N_2267,In_921,In_1264);
xnor U2268 (N_2268,In_1582,In_1164);
and U2269 (N_2269,In_565,In_1556);
nor U2270 (N_2270,In_1325,In_2071);
nand U2271 (N_2271,In_705,In_1047);
nor U2272 (N_2272,In_2027,In_1597);
and U2273 (N_2273,In_1437,In_687);
nor U2274 (N_2274,In_2461,In_2499);
and U2275 (N_2275,In_2196,In_992);
nand U2276 (N_2276,In_845,In_1166);
xnor U2277 (N_2277,In_687,In_547);
or U2278 (N_2278,In_1966,In_611);
nand U2279 (N_2279,In_1540,In_440);
and U2280 (N_2280,In_1679,In_1174);
and U2281 (N_2281,In_1389,In_2072);
and U2282 (N_2282,In_251,In_2349);
nor U2283 (N_2283,In_907,In_2316);
or U2284 (N_2284,In_31,In_621);
xnor U2285 (N_2285,In_1733,In_2404);
nor U2286 (N_2286,In_1434,In_1685);
or U2287 (N_2287,In_449,In_1412);
xor U2288 (N_2288,In_2203,In_2352);
or U2289 (N_2289,In_312,In_929);
nor U2290 (N_2290,In_702,In_288);
nor U2291 (N_2291,In_2238,In_1234);
nand U2292 (N_2292,In_398,In_1371);
and U2293 (N_2293,In_456,In_2041);
and U2294 (N_2294,In_2416,In_500);
or U2295 (N_2295,In_1997,In_345);
and U2296 (N_2296,In_2267,In_272);
nor U2297 (N_2297,In_2031,In_2013);
nand U2298 (N_2298,In_1230,In_2131);
or U2299 (N_2299,In_1153,In_920);
nand U2300 (N_2300,In_2163,In_708);
nor U2301 (N_2301,In_337,In_931);
nand U2302 (N_2302,In_1084,In_59);
nand U2303 (N_2303,In_405,In_2244);
nor U2304 (N_2304,In_1021,In_1585);
or U2305 (N_2305,In_1604,In_1904);
and U2306 (N_2306,In_776,In_68);
nand U2307 (N_2307,In_1275,In_814);
nand U2308 (N_2308,In_2156,In_362);
xnor U2309 (N_2309,In_1540,In_1506);
and U2310 (N_2310,In_2361,In_1578);
nor U2311 (N_2311,In_1226,In_158);
nand U2312 (N_2312,In_1373,In_1212);
and U2313 (N_2313,In_998,In_981);
nand U2314 (N_2314,In_2298,In_1099);
nor U2315 (N_2315,In_1982,In_750);
xor U2316 (N_2316,In_1151,In_1873);
or U2317 (N_2317,In_1857,In_2136);
xnor U2318 (N_2318,In_2084,In_187);
nor U2319 (N_2319,In_1535,In_275);
nor U2320 (N_2320,In_785,In_414);
nor U2321 (N_2321,In_1152,In_2200);
nor U2322 (N_2322,In_1066,In_2230);
nor U2323 (N_2323,In_1672,In_1898);
nand U2324 (N_2324,In_2288,In_1902);
nand U2325 (N_2325,In_2099,In_1551);
nor U2326 (N_2326,In_1160,In_1835);
and U2327 (N_2327,In_217,In_161);
nand U2328 (N_2328,In_1004,In_2232);
nor U2329 (N_2329,In_1876,In_667);
nor U2330 (N_2330,In_860,In_584);
xnor U2331 (N_2331,In_451,In_1079);
xnor U2332 (N_2332,In_59,In_286);
xor U2333 (N_2333,In_2497,In_1960);
nor U2334 (N_2334,In_779,In_1499);
xor U2335 (N_2335,In_1421,In_2372);
or U2336 (N_2336,In_1499,In_638);
xor U2337 (N_2337,In_32,In_1775);
or U2338 (N_2338,In_2198,In_126);
or U2339 (N_2339,In_284,In_1412);
or U2340 (N_2340,In_1581,In_1148);
or U2341 (N_2341,In_996,In_1469);
or U2342 (N_2342,In_46,In_735);
nand U2343 (N_2343,In_2336,In_1756);
xnor U2344 (N_2344,In_468,In_163);
xor U2345 (N_2345,In_2233,In_2064);
xor U2346 (N_2346,In_972,In_1562);
nor U2347 (N_2347,In_2286,In_920);
xor U2348 (N_2348,In_84,In_2111);
or U2349 (N_2349,In_2125,In_795);
nor U2350 (N_2350,In_2443,In_393);
xnor U2351 (N_2351,In_697,In_1395);
xor U2352 (N_2352,In_173,In_1021);
nand U2353 (N_2353,In_341,In_1060);
nor U2354 (N_2354,In_2182,In_379);
nand U2355 (N_2355,In_1934,In_2298);
xor U2356 (N_2356,In_1069,In_929);
or U2357 (N_2357,In_2311,In_73);
or U2358 (N_2358,In_2390,In_1625);
nor U2359 (N_2359,In_1463,In_2049);
xnor U2360 (N_2360,In_1154,In_1763);
and U2361 (N_2361,In_1194,In_1742);
and U2362 (N_2362,In_233,In_983);
nor U2363 (N_2363,In_2215,In_508);
nand U2364 (N_2364,In_1079,In_767);
xor U2365 (N_2365,In_545,In_2271);
xor U2366 (N_2366,In_137,In_1700);
or U2367 (N_2367,In_974,In_1398);
nor U2368 (N_2368,In_927,In_1055);
xor U2369 (N_2369,In_1401,In_1835);
xnor U2370 (N_2370,In_2275,In_1952);
and U2371 (N_2371,In_1059,In_747);
or U2372 (N_2372,In_1614,In_2449);
or U2373 (N_2373,In_647,In_1168);
nand U2374 (N_2374,In_2342,In_544);
or U2375 (N_2375,In_325,In_799);
and U2376 (N_2376,In_1255,In_1273);
or U2377 (N_2377,In_59,In_523);
nand U2378 (N_2378,In_2274,In_2497);
xor U2379 (N_2379,In_2137,In_1954);
or U2380 (N_2380,In_759,In_1994);
nand U2381 (N_2381,In_1308,In_1047);
or U2382 (N_2382,In_21,In_2111);
and U2383 (N_2383,In_1137,In_985);
xor U2384 (N_2384,In_1857,In_22);
xnor U2385 (N_2385,In_1854,In_791);
nor U2386 (N_2386,In_1277,In_1804);
nand U2387 (N_2387,In_1450,In_1796);
nor U2388 (N_2388,In_2090,In_1724);
nor U2389 (N_2389,In_1314,In_1872);
xor U2390 (N_2390,In_1877,In_590);
nor U2391 (N_2391,In_833,In_2468);
xor U2392 (N_2392,In_1247,In_850);
or U2393 (N_2393,In_1988,In_1495);
nor U2394 (N_2394,In_678,In_1288);
and U2395 (N_2395,In_606,In_1776);
xor U2396 (N_2396,In_1433,In_2380);
or U2397 (N_2397,In_155,In_1919);
and U2398 (N_2398,In_196,In_1846);
and U2399 (N_2399,In_1810,In_35);
nand U2400 (N_2400,In_623,In_473);
or U2401 (N_2401,In_209,In_1532);
or U2402 (N_2402,In_317,In_2268);
xor U2403 (N_2403,In_493,In_2262);
and U2404 (N_2404,In_5,In_2056);
or U2405 (N_2405,In_1337,In_1936);
nor U2406 (N_2406,In_1107,In_2121);
xor U2407 (N_2407,In_210,In_1414);
and U2408 (N_2408,In_160,In_1211);
xor U2409 (N_2409,In_615,In_1407);
and U2410 (N_2410,In_2386,In_1978);
nand U2411 (N_2411,In_804,In_284);
or U2412 (N_2412,In_170,In_2255);
or U2413 (N_2413,In_2026,In_1048);
or U2414 (N_2414,In_1703,In_921);
xnor U2415 (N_2415,In_696,In_141);
nand U2416 (N_2416,In_1587,In_1090);
and U2417 (N_2417,In_860,In_656);
xor U2418 (N_2418,In_1631,In_2372);
or U2419 (N_2419,In_1378,In_1656);
nor U2420 (N_2420,In_1045,In_2054);
nor U2421 (N_2421,In_825,In_1978);
and U2422 (N_2422,In_2497,In_1184);
nand U2423 (N_2423,In_205,In_1437);
nand U2424 (N_2424,In_1167,In_894);
or U2425 (N_2425,In_2495,In_289);
nor U2426 (N_2426,In_2076,In_9);
and U2427 (N_2427,In_1358,In_1077);
and U2428 (N_2428,In_2401,In_1385);
or U2429 (N_2429,In_1503,In_2343);
and U2430 (N_2430,In_1025,In_467);
or U2431 (N_2431,In_2236,In_2223);
or U2432 (N_2432,In_1551,In_1150);
and U2433 (N_2433,In_445,In_1514);
or U2434 (N_2434,In_490,In_433);
nor U2435 (N_2435,In_1217,In_853);
and U2436 (N_2436,In_1246,In_2156);
or U2437 (N_2437,In_651,In_811);
nor U2438 (N_2438,In_246,In_1129);
xor U2439 (N_2439,In_1653,In_1352);
nand U2440 (N_2440,In_2177,In_999);
xor U2441 (N_2441,In_1280,In_2434);
nand U2442 (N_2442,In_1044,In_453);
or U2443 (N_2443,In_119,In_808);
xor U2444 (N_2444,In_801,In_267);
xor U2445 (N_2445,In_734,In_1198);
nand U2446 (N_2446,In_464,In_897);
and U2447 (N_2447,In_612,In_2173);
or U2448 (N_2448,In_1695,In_556);
nor U2449 (N_2449,In_1535,In_704);
or U2450 (N_2450,In_849,In_2187);
nor U2451 (N_2451,In_1521,In_987);
and U2452 (N_2452,In_1710,In_2431);
and U2453 (N_2453,In_1204,In_2136);
nand U2454 (N_2454,In_149,In_759);
nor U2455 (N_2455,In_2154,In_1922);
nand U2456 (N_2456,In_960,In_2436);
xnor U2457 (N_2457,In_1019,In_946);
and U2458 (N_2458,In_278,In_882);
nand U2459 (N_2459,In_75,In_1483);
nor U2460 (N_2460,In_2075,In_2300);
and U2461 (N_2461,In_1804,In_2424);
xnor U2462 (N_2462,In_130,In_37);
nor U2463 (N_2463,In_548,In_2003);
nand U2464 (N_2464,In_901,In_1720);
and U2465 (N_2465,In_1426,In_706);
or U2466 (N_2466,In_1843,In_2272);
or U2467 (N_2467,In_2130,In_1855);
or U2468 (N_2468,In_1893,In_617);
xor U2469 (N_2469,In_411,In_395);
or U2470 (N_2470,In_349,In_1324);
nor U2471 (N_2471,In_2239,In_1371);
or U2472 (N_2472,In_1454,In_853);
nor U2473 (N_2473,In_1257,In_2473);
or U2474 (N_2474,In_60,In_750);
xnor U2475 (N_2475,In_2357,In_1036);
and U2476 (N_2476,In_369,In_2011);
nor U2477 (N_2477,In_2253,In_1264);
nand U2478 (N_2478,In_793,In_563);
and U2479 (N_2479,In_641,In_1051);
or U2480 (N_2480,In_1757,In_2090);
xor U2481 (N_2481,In_354,In_1962);
nor U2482 (N_2482,In_93,In_354);
or U2483 (N_2483,In_57,In_252);
xor U2484 (N_2484,In_36,In_980);
and U2485 (N_2485,In_1648,In_1786);
xnor U2486 (N_2486,In_625,In_963);
and U2487 (N_2487,In_224,In_534);
nand U2488 (N_2488,In_326,In_1087);
nor U2489 (N_2489,In_150,In_49);
nor U2490 (N_2490,In_1052,In_2430);
nor U2491 (N_2491,In_760,In_148);
xnor U2492 (N_2492,In_821,In_2399);
and U2493 (N_2493,In_895,In_1048);
nand U2494 (N_2494,In_236,In_2078);
nand U2495 (N_2495,In_2400,In_1561);
or U2496 (N_2496,In_2385,In_144);
xnor U2497 (N_2497,In_112,In_1785);
and U2498 (N_2498,In_44,In_2239);
or U2499 (N_2499,In_1441,In_1260);
nand U2500 (N_2500,N_1275,N_846);
and U2501 (N_2501,N_1942,N_1084);
or U2502 (N_2502,N_100,N_2161);
nand U2503 (N_2503,N_40,N_2486);
xor U2504 (N_2504,N_130,N_1531);
or U2505 (N_2505,N_1310,N_494);
nand U2506 (N_2506,N_430,N_306);
or U2507 (N_2507,N_2068,N_2412);
xnor U2508 (N_2508,N_75,N_13);
and U2509 (N_2509,N_890,N_800);
nor U2510 (N_2510,N_1500,N_2299);
nand U2511 (N_2511,N_401,N_756);
nand U2512 (N_2512,N_286,N_1219);
and U2513 (N_2513,N_266,N_499);
and U2514 (N_2514,N_1938,N_455);
or U2515 (N_2515,N_1273,N_625);
xnor U2516 (N_2516,N_438,N_1998);
nor U2517 (N_2517,N_2078,N_1544);
nand U2518 (N_2518,N_4,N_281);
and U2519 (N_2519,N_1792,N_2131);
and U2520 (N_2520,N_1511,N_26);
xnor U2521 (N_2521,N_2401,N_1873);
xnor U2522 (N_2522,N_956,N_757);
nand U2523 (N_2523,N_1695,N_1237);
and U2524 (N_2524,N_1823,N_2357);
nor U2525 (N_2525,N_1699,N_360);
xnor U2526 (N_2526,N_1917,N_791);
xor U2527 (N_2527,N_2134,N_1092);
and U2528 (N_2528,N_1952,N_2102);
nand U2529 (N_2529,N_18,N_63);
and U2530 (N_2530,N_1152,N_146);
nand U2531 (N_2531,N_2145,N_1067);
xor U2532 (N_2532,N_802,N_2167);
and U2533 (N_2533,N_312,N_763);
and U2534 (N_2534,N_1814,N_1257);
xnor U2535 (N_2535,N_1741,N_553);
nand U2536 (N_2536,N_1181,N_2154);
and U2537 (N_2537,N_876,N_1553);
nand U2538 (N_2538,N_285,N_2436);
or U2539 (N_2539,N_1651,N_79);
nor U2540 (N_2540,N_1317,N_969);
or U2541 (N_2541,N_886,N_2090);
nand U2542 (N_2542,N_1510,N_2282);
nor U2543 (N_2543,N_664,N_1159);
nand U2544 (N_2544,N_1138,N_2229);
nand U2545 (N_2545,N_443,N_1689);
xnor U2546 (N_2546,N_138,N_234);
and U2547 (N_2547,N_2247,N_1588);
nor U2548 (N_2548,N_1516,N_1345);
and U2549 (N_2549,N_1327,N_177);
nor U2550 (N_2550,N_399,N_538);
and U2551 (N_2551,N_69,N_1812);
and U2552 (N_2552,N_2253,N_477);
and U2553 (N_2553,N_1660,N_1635);
and U2554 (N_2554,N_900,N_423);
nand U2555 (N_2555,N_2328,N_261);
and U2556 (N_2556,N_920,N_2136);
nand U2557 (N_2557,N_1491,N_987);
or U2558 (N_2558,N_1734,N_1796);
and U2559 (N_2559,N_482,N_2203);
and U2560 (N_2560,N_2392,N_916);
xnor U2561 (N_2561,N_2112,N_774);
nand U2562 (N_2562,N_1527,N_684);
and U2563 (N_2563,N_1529,N_1183);
xnor U2564 (N_2564,N_772,N_996);
and U2565 (N_2565,N_682,N_1535);
nand U2566 (N_2566,N_1150,N_1973);
or U2567 (N_2567,N_2406,N_1398);
and U2568 (N_2568,N_391,N_2245);
or U2569 (N_2569,N_2016,N_822);
or U2570 (N_2570,N_2346,N_2219);
and U2571 (N_2571,N_2121,N_1871);
nand U2572 (N_2572,N_1013,N_1051);
xnor U2573 (N_2573,N_2238,N_1528);
and U2574 (N_2574,N_583,N_1819);
and U2575 (N_2575,N_354,N_1655);
and U2576 (N_2576,N_1388,N_1820);
and U2577 (N_2577,N_2296,N_1808);
nor U2578 (N_2578,N_831,N_631);
and U2579 (N_2579,N_677,N_1561);
and U2580 (N_2580,N_1109,N_1639);
and U2581 (N_2581,N_135,N_357);
and U2582 (N_2582,N_2276,N_1321);
xor U2583 (N_2583,N_1936,N_2028);
or U2584 (N_2584,N_27,N_2051);
xnor U2585 (N_2585,N_1851,N_47);
xor U2586 (N_2586,N_1996,N_2073);
nor U2587 (N_2587,N_781,N_1986);
and U2588 (N_2588,N_1427,N_850);
nand U2589 (N_2589,N_983,N_1867);
nand U2590 (N_2590,N_191,N_1991);
or U2591 (N_2591,N_137,N_979);
nand U2592 (N_2592,N_1325,N_1073);
and U2593 (N_2593,N_2023,N_1049);
and U2594 (N_2594,N_1974,N_673);
xnor U2595 (N_2595,N_291,N_1633);
nand U2596 (N_2596,N_1941,N_1171);
and U2597 (N_2597,N_1676,N_1293);
nand U2598 (N_2598,N_168,N_2224);
nor U2599 (N_2599,N_1570,N_1057);
xnor U2600 (N_2600,N_2222,N_1626);
nand U2601 (N_2601,N_595,N_1962);
nand U2602 (N_2602,N_1857,N_1059);
nor U2603 (N_2603,N_1415,N_628);
nor U2604 (N_2604,N_1311,N_1536);
nand U2605 (N_2605,N_1967,N_1198);
xnor U2606 (N_2606,N_990,N_2140);
nor U2607 (N_2607,N_1196,N_1399);
nand U2608 (N_2608,N_1368,N_1855);
nand U2609 (N_2609,N_542,N_816);
nand U2610 (N_2610,N_2092,N_340);
nor U2611 (N_2611,N_1740,N_1730);
and U2612 (N_2612,N_671,N_158);
nor U2613 (N_2613,N_1680,N_435);
and U2614 (N_2614,N_2309,N_2065);
and U2615 (N_2615,N_726,N_374);
and U2616 (N_2616,N_2302,N_1443);
nand U2617 (N_2617,N_1961,N_2223);
and U2618 (N_2618,N_1687,N_372);
and U2619 (N_2619,N_1424,N_1296);
xor U2620 (N_2620,N_1753,N_777);
xnor U2621 (N_2621,N_1397,N_1620);
or U2622 (N_2622,N_106,N_200);
nand U2623 (N_2623,N_1297,N_1457);
or U2624 (N_2624,N_1582,N_12);
nor U2625 (N_2625,N_2054,N_195);
nor U2626 (N_2626,N_276,N_2288);
and U2627 (N_2627,N_641,N_43);
and U2628 (N_2628,N_814,N_97);
nand U2629 (N_2629,N_761,N_919);
or U2630 (N_2630,N_141,N_1675);
nand U2631 (N_2631,N_2022,N_730);
or U2632 (N_2632,N_714,N_743);
and U2633 (N_2633,N_1343,N_2189);
nor U2634 (N_2634,N_38,N_1971);
nand U2635 (N_2635,N_1475,N_269);
or U2636 (N_2636,N_1357,N_1050);
nand U2637 (N_2637,N_2158,N_2368);
nand U2638 (N_2638,N_186,N_1265);
nor U2639 (N_2639,N_1909,N_1579);
nor U2640 (N_2640,N_390,N_1141);
nor U2641 (N_2641,N_944,N_1173);
or U2642 (N_2642,N_363,N_2106);
nand U2643 (N_2643,N_1509,N_1117);
or U2644 (N_2644,N_505,N_1768);
or U2645 (N_2645,N_1701,N_835);
nor U2646 (N_2646,N_2211,N_84);
nand U2647 (N_2647,N_635,N_1568);
nor U2648 (N_2648,N_790,N_1503);
nand U2649 (N_2649,N_1764,N_2059);
xnor U2650 (N_2650,N_984,N_2495);
and U2651 (N_2651,N_2002,N_744);
or U2652 (N_2652,N_1713,N_87);
nand U2653 (N_2653,N_806,N_1774);
nor U2654 (N_2654,N_907,N_1664);
nor U2655 (N_2655,N_1682,N_96);
nor U2656 (N_2656,N_2149,N_2294);
nand U2657 (N_2657,N_819,N_532);
and U2658 (N_2658,N_2297,N_1284);
nand U2659 (N_2659,N_1733,N_895);
and U2660 (N_2660,N_1889,N_1100);
or U2661 (N_2661,N_828,N_1672);
xor U2662 (N_2662,N_1677,N_1720);
nand U2663 (N_2663,N_1088,N_842);
xor U2664 (N_2664,N_1476,N_782);
nand U2665 (N_2665,N_597,N_1316);
and U2666 (N_2666,N_1641,N_1959);
xor U2667 (N_2667,N_145,N_1209);
and U2668 (N_2668,N_1391,N_2034);
xnor U2669 (N_2669,N_1806,N_860);
xnor U2670 (N_2670,N_105,N_1665);
nor U2671 (N_2671,N_2267,N_2234);
nand U2672 (N_2672,N_1018,N_1069);
nor U2673 (N_2673,N_844,N_1776);
nand U2674 (N_2674,N_3,N_1216);
xnor U2675 (N_2675,N_1251,N_1935);
nand U2676 (N_2676,N_1156,N_1371);
nand U2677 (N_2677,N_1172,N_1132);
or U2678 (N_2678,N_325,N_1353);
or U2679 (N_2679,N_210,N_1471);
nand U2680 (N_2680,N_1188,N_1167);
and U2681 (N_2681,N_924,N_2340);
and U2682 (N_2682,N_2487,N_1349);
nand U2683 (N_2683,N_1356,N_115);
nand U2684 (N_2684,N_2115,N_1289);
xor U2685 (N_2685,N_2249,N_1473);
and U2686 (N_2686,N_1389,N_2411);
or U2687 (N_2687,N_273,N_1148);
nand U2688 (N_2688,N_849,N_299);
and U2689 (N_2689,N_787,N_1339);
xnor U2690 (N_2690,N_676,N_20);
nor U2691 (N_2691,N_1915,N_974);
nor U2692 (N_2692,N_174,N_859);
xnor U2693 (N_2693,N_1605,N_2334);
and U2694 (N_2694,N_1179,N_1609);
nand U2695 (N_2695,N_1763,N_2263);
xnor U2696 (N_2696,N_652,N_927);
nand U2697 (N_2697,N_509,N_1124);
or U2698 (N_2698,N_2186,N_2165);
and U2699 (N_2699,N_301,N_1691);
nor U2700 (N_2700,N_446,N_598);
or U2701 (N_2701,N_466,N_2349);
or U2702 (N_2702,N_2385,N_1824);
or U2703 (N_2703,N_1143,N_1032);
or U2704 (N_2704,N_1187,N_656);
nor U2705 (N_2705,N_1233,N_552);
or U2706 (N_2706,N_386,N_793);
xnor U2707 (N_2707,N_2491,N_897);
nor U2708 (N_2708,N_1850,N_508);
nand U2709 (N_2709,N_1432,N_1074);
xnor U2710 (N_2710,N_1557,N_1523);
xnor U2711 (N_2711,N_522,N_929);
nor U2712 (N_2712,N_2183,N_856);
or U2713 (N_2713,N_1186,N_609);
nand U2714 (N_2714,N_140,N_2422);
nand U2715 (N_2715,N_1817,N_1895);
nand U2716 (N_2716,N_563,N_175);
nand U2717 (N_2717,N_1797,N_884);
xnor U2718 (N_2718,N_1359,N_39);
nor U2719 (N_2719,N_231,N_2152);
nand U2720 (N_2720,N_236,N_588);
xor U2721 (N_2721,N_537,N_1494);
xor U2722 (N_2722,N_881,N_2470);
and U2723 (N_2723,N_1872,N_392);
or U2724 (N_2724,N_573,N_2004);
xor U2725 (N_2725,N_948,N_1882);
nor U2726 (N_2726,N_975,N_1087);
nor U2727 (N_2727,N_2235,N_2440);
or U2728 (N_2728,N_1136,N_2214);
and U2729 (N_2729,N_1309,N_1006);
xor U2730 (N_2730,N_836,N_1847);
or U2731 (N_2731,N_2450,N_6);
nor U2732 (N_2732,N_1449,N_1694);
xnor U2733 (N_2733,N_674,N_2315);
nand U2734 (N_2734,N_1729,N_300);
nor U2735 (N_2735,N_998,N_720);
or U2736 (N_2736,N_1906,N_621);
nand U2737 (N_2737,N_440,N_2494);
or U2738 (N_2738,N_1843,N_1052);
and U2739 (N_2739,N_2147,N_1910);
xnor U2740 (N_2740,N_1990,N_2182);
or U2741 (N_2741,N_1684,N_1461);
nor U2742 (N_2742,N_1184,N_35);
nor U2743 (N_2743,N_288,N_81);
or U2744 (N_2744,N_449,N_10);
and U2745 (N_2745,N_2415,N_1394);
xnor U2746 (N_2746,N_578,N_2482);
nand U2747 (N_2747,N_1728,N_2321);
or U2748 (N_2748,N_955,N_1418);
and U2749 (N_2749,N_544,N_1279);
xor U2750 (N_2750,N_1189,N_2025);
nor U2751 (N_2751,N_855,N_205);
or U2752 (N_2752,N_259,N_2118);
or U2753 (N_2753,N_1539,N_1900);
nand U2754 (N_2754,N_1381,N_507);
nand U2755 (N_2755,N_820,N_993);
and U2756 (N_2756,N_1893,N_478);
xnor U2757 (N_2757,N_1395,N_1761);
xor U2758 (N_2758,N_1769,N_208);
and U2759 (N_2759,N_2373,N_1315);
xor U2760 (N_2760,N_610,N_89);
nor U2761 (N_2761,N_420,N_1506);
xnor U2762 (N_2762,N_1744,N_870);
and U2763 (N_2763,N_464,N_1408);
nor U2764 (N_2764,N_556,N_502);
or U2765 (N_2765,N_1295,N_1624);
or U2766 (N_2766,N_2421,N_1592);
nor U2767 (N_2767,N_1656,N_1319);
nor U2768 (N_2768,N_1426,N_701);
xnor U2769 (N_2769,N_190,N_1521);
or U2770 (N_2770,N_1147,N_2383);
nand U2771 (N_2771,N_214,N_2089);
nor U2772 (N_2772,N_2286,N_416);
nand U2773 (N_2773,N_2451,N_2259);
xor U2774 (N_2774,N_1280,N_1618);
nand U2775 (N_2775,N_144,N_1463);
or U2776 (N_2776,N_1590,N_1256);
or U2777 (N_2777,N_1888,N_1501);
xor U2778 (N_2778,N_1305,N_2379);
and U2779 (N_2779,N_873,N_1331);
nor U2780 (N_2780,N_471,N_2017);
nand U2781 (N_2781,N_2105,N_2339);
nand U2782 (N_2782,N_773,N_1870);
nor U2783 (N_2783,N_131,N_1925);
and U2784 (N_2784,N_1780,N_2413);
xnor U2785 (N_2785,N_1993,N_219);
and U2786 (N_2786,N_933,N_1487);
nor U2787 (N_2787,N_2326,N_558);
nand U2788 (N_2788,N_1286,N_344);
nand U2789 (N_2789,N_1572,N_810);
xor U2790 (N_2790,N_2003,N_2208);
nor U2791 (N_2791,N_1621,N_167);
nand U2792 (N_2792,N_1164,N_910);
nand U2793 (N_2793,N_2039,N_1229);
xor U2794 (N_2794,N_909,N_1044);
xnor U2795 (N_2795,N_465,N_1596);
and U2796 (N_2796,N_541,N_104);
xnor U2797 (N_2797,N_1243,N_1362);
nand U2798 (N_2798,N_21,N_692);
nor U2799 (N_2799,N_798,N_603);
or U2800 (N_2800,N_1272,N_1522);
and U2801 (N_2801,N_808,N_687);
or U2802 (N_2802,N_2046,N_48);
nand U2803 (N_2803,N_415,N_1448);
nand U2804 (N_2804,N_2418,N_862);
nand U2805 (N_2805,N_1116,N_2081);
nand U2806 (N_2806,N_1122,N_1901);
or U2807 (N_2807,N_706,N_338);
and U2808 (N_2808,N_1988,N_5);
or U2809 (N_2809,N_2175,N_162);
xnor U2810 (N_2810,N_1025,N_62);
nor U2811 (N_2811,N_1799,N_945);
and U2812 (N_2812,N_2497,N_1745);
and U2813 (N_2813,N_143,N_217);
nor U2814 (N_2814,N_2327,N_258);
or U2815 (N_2815,N_2159,N_150);
nand U2816 (N_2816,N_2100,N_837);
nand U2817 (N_2817,N_437,N_2367);
nor U2818 (N_2818,N_1790,N_1913);
nor U2819 (N_2819,N_758,N_616);
or U2820 (N_2820,N_294,N_1079);
xnor U2821 (N_2821,N_973,N_1829);
xnor U2822 (N_2822,N_2481,N_1930);
nor U2823 (N_2823,N_2384,N_1789);
and U2824 (N_2824,N_2292,N_1028);
nor U2825 (N_2825,N_123,N_848);
nor U2826 (N_2826,N_1844,N_302);
and U2827 (N_2827,N_657,N_1003);
nor U2828 (N_2828,N_1840,N_1948);
xnor U2829 (N_2829,N_1169,N_2466);
and U2830 (N_2830,N_712,N_1224);
xor U2831 (N_2831,N_2213,N_2344);
nand U2832 (N_2832,N_2428,N_1578);
xor U2833 (N_2833,N_1390,N_982);
nor U2834 (N_2834,N_1340,N_683);
nor U2835 (N_2835,N_2362,N_1354);
nand U2836 (N_2836,N_1751,N_645);
or U2837 (N_2837,N_1520,N_1538);
nor U2838 (N_2838,N_1543,N_1098);
nand U2839 (N_2839,N_1704,N_2166);
nand U2840 (N_2840,N_1387,N_2433);
nand U2841 (N_2841,N_11,N_847);
nand U2842 (N_2842,N_1756,N_2129);
and U2843 (N_2843,N_1153,N_218);
xor U2844 (N_2844,N_1249,N_569);
or U2845 (N_2845,N_659,N_1194);
xnor U2846 (N_2846,N_2289,N_1940);
nor U2847 (N_2847,N_1903,N_232);
and U2848 (N_2848,N_711,N_2255);
nor U2849 (N_2849,N_606,N_93);
or U2850 (N_2850,N_2067,N_918);
or U2851 (N_2851,N_602,N_1377);
xnor U2852 (N_2852,N_1615,N_2021);
nor U2853 (N_2853,N_2431,N_2236);
nor U2854 (N_2854,N_2132,N_270);
nor U2855 (N_2855,N_1593,N_1640);
nor U2856 (N_2856,N_579,N_1671);
xor U2857 (N_2857,N_1920,N_361);
nand U2858 (N_2858,N_1165,N_1746);
nand U2859 (N_2859,N_125,N_1031);
nor U2860 (N_2860,N_2047,N_752);
nand U2861 (N_2861,N_871,N_1253);
nand U2862 (N_2862,N_1496,N_738);
and U2863 (N_2863,N_1658,N_2419);
or U2864 (N_2864,N_380,N_1055);
nor U2865 (N_2865,N_1770,N_335);
nand U2866 (N_2866,N_1337,N_393);
or U2867 (N_2867,N_1541,N_995);
xor U2868 (N_2868,N_2285,N_1804);
nand U2869 (N_2869,N_1139,N_1046);
nand U2870 (N_2870,N_2133,N_129);
nor U2871 (N_2871,N_2071,N_230);
or U2872 (N_2872,N_575,N_364);
or U2873 (N_2873,N_2416,N_412);
or U2874 (N_2874,N_1897,N_1162);
and U2875 (N_2875,N_2232,N_2478);
nor U2876 (N_2876,N_592,N_193);
and U2877 (N_2877,N_126,N_1569);
nor U2878 (N_2878,N_1191,N_1679);
or U2879 (N_2879,N_2192,N_1404);
or U2880 (N_2880,N_1502,N_500);
nand U2881 (N_2881,N_2455,N_348);
and U2882 (N_2882,N_1382,N_1118);
nor U2883 (N_2883,N_1213,N_452);
or U2884 (N_2884,N_53,N_362);
nand U2885 (N_2885,N_2389,N_572);
or U2886 (N_2886,N_1488,N_1029);
and U2887 (N_2887,N_695,N_2432);
nor U2888 (N_2888,N_2391,N_1396);
nor U2889 (N_2889,N_1841,N_1452);
nor U2890 (N_2890,N_2142,N_986);
nor U2891 (N_2891,N_785,N_2057);
xnor U2892 (N_2892,N_665,N_794);
or U2893 (N_2893,N_874,N_932);
or U2894 (N_2894,N_1619,N_462);
or U2895 (N_2895,N_483,N_2269);
or U2896 (N_2896,N_2030,N_1137);
nand U2897 (N_2897,N_506,N_1324);
nor U2898 (N_2898,N_289,N_1722);
or U2899 (N_2899,N_1782,N_957);
nor U2900 (N_2900,N_2493,N_426);
xor U2901 (N_2901,N_2246,N_1423);
nor U2902 (N_2902,N_142,N_282);
nor U2903 (N_2903,N_2029,N_2113);
or U2904 (N_2904,N_1105,N_2280);
or U2905 (N_2905,N_1760,N_1886);
or U2906 (N_2906,N_334,N_257);
nand U2907 (N_2907,N_1831,N_1364);
nor U2908 (N_2908,N_1956,N_283);
and U2909 (N_2909,N_1946,N_1208);
and U2910 (N_2910,N_1083,N_1195);
nor U2911 (N_2911,N_2007,N_2194);
or U2912 (N_2912,N_562,N_428);
nand U2913 (N_2913,N_1185,N_1955);
xnor U2914 (N_2914,N_1921,N_2460);
nor U2915 (N_2915,N_1375,N_2061);
nand U2916 (N_2916,N_718,N_1612);
xor U2917 (N_2917,N_680,N_1202);
nor U2918 (N_2918,N_1560,N_663);
xor U2919 (N_2919,N_1611,N_868);
or U2920 (N_2920,N_1261,N_463);
or U2921 (N_2921,N_1931,N_1009);
nand U2922 (N_2922,N_2171,N_2104);
nand U2923 (N_2923,N_1786,N_1772);
and U2924 (N_2924,N_1458,N_1863);
nand U2925 (N_2925,N_1113,N_2448);
nand U2926 (N_2926,N_134,N_830);
nor U2927 (N_2927,N_1735,N_2143);
nor U2928 (N_2928,N_1053,N_702);
or U2929 (N_2929,N_98,N_1222);
xnor U2930 (N_2930,N_1647,N_1042);
nand U2931 (N_2931,N_1657,N_1292);
and U2932 (N_2932,N_57,N_1795);
nand U2933 (N_2933,N_804,N_235);
nor U2934 (N_2934,N_1126,N_1468);
nor U2935 (N_2935,N_764,N_1530);
nor U2936 (N_2936,N_404,N_2086);
nor U2937 (N_2937,N_1777,N_1258);
nand U2938 (N_2938,N_2170,N_171);
or U2939 (N_2939,N_1816,N_807);
nor U2940 (N_2940,N_342,N_1532);
nand U2941 (N_2941,N_169,N_166);
nor U2942 (N_2942,N_894,N_1016);
nand U2943 (N_2943,N_1944,N_1235);
or U2944 (N_2944,N_1610,N_2045);
xor U2945 (N_2945,N_182,N_2172);
or U2946 (N_2946,N_2241,N_1800);
and U2947 (N_2947,N_1607,N_1373);
nor U2948 (N_2948,N_1697,N_124);
and U2949 (N_2949,N_333,N_337);
xor U2950 (N_2950,N_2434,N_2402);
and U2951 (N_2951,N_2014,N_1163);
nand U2952 (N_2952,N_1827,N_1552);
and U2953 (N_2953,N_1849,N_1548);
xnor U2954 (N_2954,N_533,N_295);
or U2955 (N_2955,N_2008,N_133);
nor U2956 (N_2956,N_2283,N_2011);
and U2957 (N_2957,N_1815,N_2414);
nand U2958 (N_2958,N_2496,N_1645);
xnor U2959 (N_2959,N_1393,N_554);
nand U2960 (N_2960,N_574,N_2403);
nor U2961 (N_2961,N_265,N_77);
and U2962 (N_2962,N_2453,N_1158);
nand U2963 (N_2963,N_1039,N_1864);
nand U2964 (N_2964,N_2128,N_2366);
nand U2965 (N_2965,N_189,N_1563);
and U2966 (N_2966,N_1743,N_1600);
or U2967 (N_2967,N_2336,N_2323);
xnor U2968 (N_2968,N_2271,N_1040);
nand U2969 (N_2969,N_978,N_959);
or U2970 (N_2970,N_1033,N_345);
nand U2971 (N_2971,N_940,N_2409);
nand U2972 (N_2972,N_580,N_318);
and U2973 (N_2973,N_1914,N_1818);
and U2974 (N_2974,N_118,N_1145);
nand U2975 (N_2975,N_604,N_748);
or U2976 (N_2976,N_2010,N_1230);
and U2977 (N_2977,N_1747,N_2228);
and U2978 (N_2978,N_1771,N_1589);
and U2979 (N_2979,N_1259,N_433);
or U2980 (N_2980,N_103,N_1101);
nand U2981 (N_2981,N_1830,N_1160);
xnor U2982 (N_2982,N_587,N_1702);
xor U2983 (N_2983,N_893,N_866);
xnor U2984 (N_2984,N_905,N_1778);
and U2985 (N_2985,N_1628,N_2405);
nand U2986 (N_2986,N_1833,N_2187);
xor U2987 (N_2987,N_127,N_225);
xor U2988 (N_2988,N_2097,N_2343);
or U2989 (N_2989,N_1455,N_1947);
nand U2990 (N_2990,N_691,N_1178);
nand U2991 (N_2991,N_2215,N_2079);
nor U2992 (N_2992,N_1,N_1919);
and U2993 (N_2993,N_626,N_1866);
xor U2994 (N_2994,N_1670,N_1080);
nor U2995 (N_2995,N_891,N_1933);
and U2996 (N_2996,N_1451,N_1303);
xnor U2997 (N_2997,N_1631,N_1762);
nor U2998 (N_2998,N_1215,N_1810);
and U2999 (N_2999,N_2160,N_963);
or U3000 (N_3000,N_1710,N_1887);
and U3001 (N_3001,N_408,N_703);
nor U3002 (N_3002,N_148,N_1976);
nor U3003 (N_3003,N_1547,N_25);
nand U3004 (N_3004,N_2274,N_267);
nand U3005 (N_3005,N_54,N_2185);
nor U3006 (N_3006,N_489,N_2430);
nand U3007 (N_3007,N_1836,N_1681);
nand U3008 (N_3008,N_369,N_2137);
nand U3009 (N_3009,N_593,N_184);
or U3010 (N_3010,N_1922,N_34);
nor U3011 (N_3011,N_519,N_398);
nand U3012 (N_3012,N_728,N_2225);
nand U3013 (N_3013,N_1878,N_2168);
xnor U3014 (N_3014,N_530,N_2290);
nor U3015 (N_3015,N_490,N_678);
nor U3016 (N_3016,N_101,N_1446);
or U3017 (N_3017,N_989,N_424);
nand U3018 (N_3018,N_2048,N_926);
nor U3019 (N_3019,N_2324,N_853);
nor U3020 (N_3020,N_1420,N_2459);
or U3021 (N_3021,N_1964,N_1436);
xnor U3022 (N_3022,N_1350,N_1963);
or U3023 (N_3023,N_2355,N_2144);
or U3024 (N_3024,N_1274,N_727);
nand U3025 (N_3025,N_1926,N_1608);
nor U3026 (N_3026,N_1248,N_1322);
or U3027 (N_3027,N_2188,N_459);
or U3028 (N_3028,N_2209,N_296);
nor U3029 (N_3029,N_2120,N_52);
nor U3030 (N_3030,N_947,N_1246);
nor U3031 (N_3031,N_840,N_2477);
or U3032 (N_3032,N_805,N_2301);
xnor U3033 (N_3033,N_476,N_1546);
nand U3034 (N_3034,N_612,N_699);
nand U3035 (N_3035,N_2268,N_1234);
xor U3036 (N_3036,N_1034,N_74);
nor U3037 (N_3037,N_1417,N_1707);
nand U3038 (N_3038,N_343,N_359);
and U3039 (N_3039,N_461,N_1135);
xor U3040 (N_3040,N_2020,N_546);
or U3041 (N_3041,N_821,N_2439);
and U3042 (N_3042,N_2244,N_1278);
or U3043 (N_3043,N_2123,N_568);
xor U3044 (N_3044,N_637,N_733);
xnor U3045 (N_3045,N_1037,N_1659);
xnor U3046 (N_3046,N_2135,N_584);
xnor U3047 (N_3047,N_551,N_739);
nand U3048 (N_3048,N_776,N_2108);
xor U3049 (N_3049,N_834,N_2488);
and U3050 (N_3050,N_2353,N_934);
and U3051 (N_3051,N_2126,N_1678);
xor U3052 (N_3052,N_936,N_293);
nand U3053 (N_3053,N_2060,N_72);
or U3054 (N_3054,N_1282,N_2337);
nand U3055 (N_3055,N_2125,N_1430);
or U3056 (N_3056,N_260,N_517);
nand U3057 (N_3057,N_419,N_1663);
or U3058 (N_3058,N_2040,N_1992);
xor U3059 (N_3059,N_1606,N_1437);
and U3060 (N_3060,N_434,N_1960);
nor U3061 (N_3061,N_2417,N_2218);
and U3062 (N_3062,N_441,N_365);
nand U3063 (N_3063,N_863,N_1070);
nor U3064 (N_3064,N_1858,N_1419);
xnor U3065 (N_3065,N_1114,N_1587);
or U3066 (N_3066,N_2293,N_1128);
or U3067 (N_3067,N_474,N_1308);
and U3068 (N_3068,N_322,N_2342);
nor U3069 (N_3069,N_1537,N_561);
or U3070 (N_3070,N_1716,N_857);
or U3071 (N_3071,N_1241,N_686);
or U3072 (N_3072,N_784,N_1149);
or U3073 (N_3073,N_1787,N_2365);
or U3074 (N_3074,N_305,N_425);
and U3075 (N_3075,N_740,N_99);
and U3076 (N_3076,N_1307,N_514);
or U3077 (N_3077,N_1724,N_762);
and U3078 (N_3078,N_116,N_248);
xnor U3079 (N_3079,N_467,N_1483);
nand U3080 (N_3080,N_321,N_2258);
nand U3081 (N_3081,N_350,N_2354);
and U3082 (N_3082,N_1591,N_539);
and U3083 (N_3083,N_1512,N_1103);
or U3084 (N_3084,N_86,N_747);
nor U3085 (N_3085,N_930,N_7);
or U3086 (N_3086,N_1081,N_1244);
or U3087 (N_3087,N_615,N_1472);
xnor U3088 (N_3088,N_937,N_1048);
xnor U3089 (N_3089,N_503,N_1466);
xor U3090 (N_3090,N_1068,N_1482);
and U3091 (N_3091,N_180,N_2457);
nor U3092 (N_3092,N_16,N_1428);
or U3093 (N_3093,N_58,N_409);
or U3094 (N_3094,N_368,N_2371);
nand U3095 (N_3095,N_36,N_442);
or U3096 (N_3096,N_1444,N_2084);
xor U3097 (N_3097,N_60,N_721);
nor U3098 (N_3098,N_256,N_2109);
nand U3099 (N_3099,N_65,N_889);
or U3100 (N_3100,N_1805,N_2099);
or U3101 (N_3101,N_2250,N_2427);
nor U3102 (N_3102,N_997,N_2447);
and U3103 (N_3103,N_1486,N_1203);
nand U3104 (N_3104,N_661,N_2278);
xnor U3105 (N_3105,N_29,N_1416);
xnor U3106 (N_3106,N_1700,N_705);
nor U3107 (N_3107,N_1879,N_576);
and U3108 (N_3108,N_1749,N_1965);
nand U3109 (N_3109,N_1868,N_1004);
nor U3110 (N_3110,N_2499,N_2077);
nand U3111 (N_3111,N_548,N_222);
nand U3112 (N_3112,N_971,N_405);
or U3113 (N_3113,N_2445,N_2360);
or U3114 (N_3114,N_1999,N_1885);
or U3115 (N_3115,N_154,N_486);
xnor U3116 (N_3116,N_2390,N_668);
xnor U3117 (N_3117,N_1983,N_778);
or U3118 (N_3118,N_759,N_1065);
nand U3119 (N_3119,N_594,N_484);
nor U3120 (N_3120,N_2303,N_2429);
xnor U3121 (N_3121,N_1650,N_94);
nand U3122 (N_3122,N_1376,N_825);
and U3123 (N_3123,N_1406,N_1407);
nor U3124 (N_3124,N_1228,N_414);
and U3125 (N_3125,N_741,N_681);
nor U3126 (N_3126,N_22,N_2333);
xnor U3127 (N_3127,N_811,N_1997);
or U3128 (N_3128,N_1554,N_287);
xnor U3129 (N_3129,N_2012,N_2318);
and U3130 (N_3130,N_1839,N_2374);
nand U3131 (N_3131,N_1927,N_187);
nor U3132 (N_3132,N_151,N_2243);
xnor U3133 (N_3133,N_2375,N_928);
xnor U3134 (N_3134,N_1062,N_2070);
and U3135 (N_3135,N_2284,N_2031);
nor U3136 (N_3136,N_1283,N_1685);
nor U3137 (N_3137,N_970,N_1063);
nand U3138 (N_3138,N_2181,N_643);
and U3139 (N_3139,N_670,N_2240);
or U3140 (N_3140,N_2304,N_339);
or U3141 (N_3141,N_896,N_2329);
and U3142 (N_3142,N_967,N_327);
xnor U3143 (N_3143,N_450,N_277);
or U3144 (N_3144,N_1540,N_64);
or U3145 (N_3145,N_326,N_1845);
nor U3146 (N_3146,N_1518,N_962);
nor U3147 (N_3147,N_1168,N_1525);
nor U3148 (N_3148,N_1586,N_2387);
nand U3149 (N_3149,N_1023,N_525);
nand U3150 (N_3150,N_2273,N_207);
and U3151 (N_3151,N_722,N_1214);
xnor U3152 (N_3152,N_2449,N_388);
nor U3153 (N_3153,N_1111,N_17);
xor U3154 (N_3154,N_1616,N_1255);
nand U3155 (N_3155,N_90,N_1583);
nor U3156 (N_3156,N_2013,N_107);
nor U3157 (N_3157,N_2179,N_253);
nor U3158 (N_3158,N_349,N_1690);
and U3159 (N_3159,N_1412,N_2242);
xnor U3160 (N_3160,N_1314,N_698);
xnor U3161 (N_3161,N_2358,N_201);
or U3162 (N_3162,N_1212,N_1134);
nor U3163 (N_3163,N_961,N_753);
nor U3164 (N_3164,N_155,N_966);
nand U3165 (N_3165,N_445,N_624);
nor U3166 (N_3166,N_843,N_1066);
nor U3167 (N_3167,N_1798,N_1456);
xnor U3168 (N_3168,N_2026,N_1803);
and U3169 (N_3169,N_617,N_198);
or U3170 (N_3170,N_566,N_1975);
or U3171 (N_3171,N_66,N_2338);
and U3172 (N_3172,N_2206,N_456);
nor U3173 (N_3173,N_2141,N_451);
or U3174 (N_3174,N_988,N_2042);
nor U3175 (N_3175,N_2093,N_119);
and U3176 (N_3176,N_358,N_220);
nor U3177 (N_3177,N_599,N_1060);
nor U3178 (N_3178,N_324,N_949);
nand U3179 (N_3179,N_902,N_2216);
and U3180 (N_3180,N_1860,N_278);
and U3181 (N_3181,N_2207,N_1240);
nor U3182 (N_3182,N_245,N_212);
xor U3183 (N_3183,N_496,N_355);
nand U3184 (N_3184,N_1218,N_1642);
xor U3185 (N_3185,N_1431,N_2062);
and U3186 (N_3186,N_1958,N_865);
nor U3187 (N_3187,N_470,N_2437);
and U3188 (N_3188,N_2176,N_2396);
or U3189 (N_3189,N_383,N_0);
xor U3190 (N_3190,N_2441,N_73);
or U3191 (N_3191,N_877,N_2361);
xnor U3192 (N_3192,N_1043,N_2322);
nor U3193 (N_3193,N_1365,N_1698);
nor U3194 (N_3194,N_213,N_745);
or U3195 (N_3195,N_1577,N_2404);
xnor U3196 (N_3196,N_1811,N_824);
and U3197 (N_3197,N_2277,N_1688);
nor U3198 (N_3198,N_185,N_1328);
and U3199 (N_3199,N_2483,N_136);
xnor U3200 (N_3200,N_2096,N_724);
or U3201 (N_3201,N_454,N_173);
nor U3202 (N_3202,N_172,N_799);
or U3203 (N_3203,N_1464,N_1320);
nand U3204 (N_3204,N_1559,N_1517);
xnor U3205 (N_3205,N_1759,N_2049);
xor U3206 (N_3206,N_1791,N_262);
xnor U3207 (N_3207,N_2484,N_1355);
or U3208 (N_3208,N_526,N_475);
nand U3209 (N_3209,N_1928,N_1211);
xor U3210 (N_3210,N_238,N_1422);
nor U3211 (N_3211,N_429,N_2180);
nand U3212 (N_3212,N_249,N_1719);
and U3213 (N_3213,N_2130,N_1932);
nand U3214 (N_3214,N_654,N_1576);
nor U3215 (N_3215,N_742,N_619);
xnor U3216 (N_3216,N_2066,N_1299);
and U3217 (N_3217,N_2220,N_2015);
nand U3218 (N_3218,N_1155,N_427);
nand U3219 (N_3219,N_2107,N_1144);
or U3220 (N_3220,N_1584,N_534);
nand U3221 (N_3221,N_1978,N_448);
or U3222 (N_3222,N_1231,N_492);
and U3223 (N_3223,N_1773,N_585);
nand U3224 (N_3224,N_1302,N_246);
and U3225 (N_3225,N_2111,N_2256);
xor U3226 (N_3226,N_2000,N_1549);
xor U3227 (N_3227,N_2264,N_1351);
or U3228 (N_3228,N_1479,N_1598);
xnor U3229 (N_3229,N_1200,N_2058);
nor U3230 (N_3230,N_943,N_1788);
xor U3231 (N_3231,N_161,N_1112);
nor U3232 (N_3232,N_2019,N_1953);
or U3233 (N_3233,N_1545,N_203);
and U3234 (N_3234,N_292,N_1467);
or U3235 (N_3235,N_2064,N_268);
xor U3236 (N_3236,N_31,N_622);
nand U3237 (N_3237,N_725,N_2435);
nand U3238 (N_3238,N_1939,N_1573);
or U3239 (N_3239,N_1714,N_170);
or U3240 (N_3240,N_2452,N_1951);
and U3241 (N_3241,N_2476,N_1378);
and U3242 (N_3242,N_2056,N_76);
xnor U3243 (N_3243,N_1347,N_1266);
or U3244 (N_3244,N_994,N_113);
nand U3245 (N_3245,N_275,N_1727);
nor U3246 (N_3246,N_1924,N_1477);
nor U3247 (N_3247,N_1638,N_1190);
and U3248 (N_3248,N_216,N_2410);
and U3249 (N_3249,N_1905,N_1329);
and U3250 (N_3250,N_112,N_1174);
xnor U3251 (N_3251,N_2356,N_1085);
or U3252 (N_3252,N_1968,N_1825);
nor U3253 (N_3253,N_1784,N_555);
xor U3254 (N_3254,N_178,N_2043);
nor U3255 (N_3255,N_223,N_550);
xor U3256 (N_3256,N_1110,N_826);
or U3257 (N_3257,N_620,N_1071);
or U3258 (N_3258,N_736,N_1410);
nor U3259 (N_3259,N_523,N_2461);
or U3260 (N_3260,N_1669,N_1835);
nor U3261 (N_3261,N_2300,N_1270);
or U3262 (N_3262,N_1891,N_1752);
or U3263 (N_3263,N_2308,N_264);
and U3264 (N_3264,N_1041,N_690);
nand U3265 (N_3265,N_1564,N_1950);
nor U3266 (N_3266,N_1054,N_1846);
nor U3267 (N_3267,N_2178,N_1721);
xor U3268 (N_3268,N_1180,N_1748);
xnor U3269 (N_3269,N_1562,N_1341);
nor U3270 (N_3270,N_2202,N_241);
nand U3271 (N_3271,N_164,N_2173);
xnor U3272 (N_3272,N_1493,N_352);
xor U3273 (N_3273,N_1984,N_1038);
and U3274 (N_3274,N_1595,N_310);
or U3275 (N_3275,N_2272,N_1750);
xnor U3276 (N_3276,N_1474,N_627);
or U3277 (N_3277,N_608,N_30);
xor U3278 (N_3278,N_1000,N_1332);
nand U3279 (N_3279,N_2261,N_1492);
and U3280 (N_3280,N_1813,N_640);
or U3281 (N_3281,N_951,N_2098);
and U3282 (N_3282,N_2,N_1090);
nor U3283 (N_3283,N_1654,N_1193);
xnor U3284 (N_3284,N_760,N_1045);
or U3285 (N_3285,N_1182,N_1366);
xnor U3286 (N_3286,N_491,N_1385);
or U3287 (N_3287,N_1252,N_328);
or U3288 (N_3288,N_2239,N_1630);
or U3289 (N_3289,N_252,N_1957);
and U3290 (N_3290,N_571,N_1227);
xor U3291 (N_3291,N_1097,N_2210);
nor U3292 (N_3292,N_1409,N_224);
nor U3293 (N_3293,N_1465,N_817);
and U3294 (N_3294,N_1338,N_1923);
nand U3295 (N_3295,N_1015,N_42);
xnor U3296 (N_3296,N_1089,N_51);
and U3297 (N_3297,N_1985,N_524);
xnor U3298 (N_3298,N_653,N_1604);
nor U3299 (N_3299,N_875,N_829);
xor U3300 (N_3300,N_1515,N_308);
nor U3301 (N_3301,N_2083,N_1358);
xor U3302 (N_3302,N_1285,N_655);
and U3303 (N_3303,N_2398,N_1462);
or U3304 (N_3304,N_176,N_2291);
xor U3305 (N_3305,N_1489,N_1614);
nor U3306 (N_3306,N_50,N_1597);
and U3307 (N_3307,N_271,N_396);
nor U3308 (N_3308,N_394,N_1142);
and U3309 (N_3309,N_1306,N_83);
or U3310 (N_3310,N_1715,N_735);
nor U3311 (N_3311,N_729,N_766);
nand U3312 (N_3312,N_2307,N_1333);
or U3313 (N_3313,N_279,N_2162);
nor U3314 (N_3314,N_823,N_215);
and U3315 (N_3315,N_1565,N_1326);
nor U3316 (N_3316,N_1551,N_2443);
xor U3317 (N_3317,N_1021,N_1078);
xor U3318 (N_3318,N_2230,N_403);
nor U3319 (N_3319,N_1267,N_1929);
xnor U3320 (N_3320,N_547,N_968);
or U3321 (N_3321,N_1705,N_1807);
nand U3322 (N_3322,N_2101,N_28);
nand U3323 (N_3323,N_1880,N_1342);
nand U3324 (N_3324,N_2316,N_2088);
and U3325 (N_3325,N_2407,N_1683);
nand U3326 (N_3326,N_431,N_809);
or U3327 (N_3327,N_1225,N_1627);
nor U3328 (N_3328,N_67,N_1361);
or U3329 (N_3329,N_567,N_801);
xnor U3330 (N_3330,N_1581,N_513);
nand U3331 (N_3331,N_1856,N_1107);
or U3332 (N_3332,N_1439,N_1892);
xor U3333 (N_3333,N_878,N_543);
nand U3334 (N_3334,N_750,N_410);
and U3335 (N_3335,N_2226,N_2347);
and U3336 (N_3336,N_1842,N_1086);
nand U3337 (N_3337,N_1459,N_347);
nor U3338 (N_3338,N_1401,N_239);
and U3339 (N_3339,N_540,N_1011);
or U3340 (N_3340,N_2227,N_950);
and U3341 (N_3341,N_1869,N_999);
nand U3342 (N_3342,N_2024,N_2050);
or U3343 (N_3343,N_2378,N_192);
and U3344 (N_3344,N_2442,N_2345);
or U3345 (N_3345,N_1005,N_1121);
nand U3346 (N_3346,N_2204,N_880);
nand U3347 (N_3347,N_2036,N_2251);
or U3348 (N_3348,N_1667,N_2076);
and U3349 (N_3349,N_1732,N_660);
and U3350 (N_3350,N_44,N_24);
nand U3351 (N_3351,N_188,N_765);
xnor U3352 (N_3352,N_648,N_1413);
or U3353 (N_3353,N_1881,N_869);
xnor U3354 (N_3354,N_976,N_715);
nor U3355 (N_3355,N_1429,N_2380);
nand U3356 (N_3356,N_2155,N_159);
and U3357 (N_3357,N_110,N_1091);
nand U3358 (N_3358,N_2005,N_1236);
nand U3359 (N_3359,N_479,N_1653);
xor U3360 (N_3360,N_2424,N_1120);
nand U3361 (N_3361,N_2369,N_1036);
nand U3362 (N_3362,N_356,N_102);
nand U3363 (N_3363,N_613,N_709);
nand U3364 (N_3364,N_1505,N_2472);
and U3365 (N_3365,N_1766,N_229);
nand U3366 (N_3366,N_196,N_713);
xor U3367 (N_3367,N_1890,N_2196);
nand U3368 (N_3368,N_2169,N_1352);
xnor U3369 (N_3369,N_770,N_2471);
nand U3370 (N_3370,N_2468,N_1300);
and U3371 (N_3371,N_1802,N_1556);
and U3372 (N_3372,N_376,N_2212);
or U3373 (N_3373,N_2311,N_303);
xor U3374 (N_3374,N_734,N_1247);
and U3375 (N_3375,N_1106,N_549);
and U3376 (N_3376,N_1896,N_160);
nand U3377 (N_3377,N_1832,N_1674);
or U3378 (N_3378,N_1022,N_1865);
or U3379 (N_3379,N_1852,N_70);
and U3380 (N_3380,N_1268,N_977);
and U3381 (N_3381,N_833,N_373);
and U3382 (N_3382,N_651,N_1130);
xor U3383 (N_3383,N_669,N_1686);
nand U3384 (N_3384,N_367,N_679);
nand U3385 (N_3385,N_560,N_59);
xor U3386 (N_3386,N_1898,N_1754);
xnor U3387 (N_3387,N_911,N_2372);
nor U3388 (N_3388,N_795,N_557);
nor U3389 (N_3389,N_2217,N_2364);
or U3390 (N_3390,N_1826,N_1970);
and U3391 (N_3391,N_1904,N_2116);
nor U3392 (N_3392,N_2423,N_1767);
and U3393 (N_3393,N_1392,N_1637);
nand U3394 (N_3394,N_710,N_2492);
xnor U3395 (N_3395,N_769,N_611);
xnor U3396 (N_3396,N_2462,N_444);
nand U3397 (N_3397,N_1223,N_2119);
xnor U3398 (N_3398,N_2426,N_1498);
xnor U3399 (N_3399,N_1076,N_1271);
nand U3400 (N_3400,N_80,N_1056);
and U3401 (N_3401,N_1012,N_242);
and U3402 (N_3402,N_1911,N_1199);
or U3403 (N_3403,N_1019,N_2341);
nand U3404 (N_3404,N_1064,N_2151);
or U3405 (N_3405,N_1907,N_1558);
nor U3406 (N_3406,N_1411,N_2464);
xnor U3407 (N_3407,N_1058,N_1969);
or U3408 (N_3408,N_2146,N_1383);
and U3409 (N_3409,N_2265,N_2153);
nand U3410 (N_3410,N_2331,N_1166);
xnor U3411 (N_3411,N_632,N_2127);
and U3412 (N_3412,N_520,N_942);
nand U3413 (N_3413,N_389,N_1372);
nor U3414 (N_3414,N_307,N_792);
nand U3415 (N_3415,N_697,N_1853);
nand U3416 (N_3416,N_511,N_577);
and U3417 (N_3417,N_879,N_1571);
and U3418 (N_3418,N_458,N_1151);
or U3419 (N_3419,N_867,N_1603);
nor U3420 (N_3420,N_1738,N_45);
or U3421 (N_3421,N_1717,N_582);
nor U3422 (N_3422,N_211,N_1217);
nand U3423 (N_3423,N_400,N_2069);
or U3424 (N_3424,N_746,N_2150);
or U3425 (N_3425,N_316,N_1708);
nor U3426 (N_3426,N_2306,N_280);
or U3427 (N_3427,N_309,N_330);
nor U3428 (N_3428,N_2052,N_480);
and U3429 (N_3429,N_1433,N_1644);
nand U3430 (N_3430,N_1238,N_737);
or U3431 (N_3431,N_323,N_1775);
or U3432 (N_3432,N_2310,N_1312);
nand U3433 (N_3433,N_1623,N_1104);
xor U3434 (N_3434,N_1131,N_1441);
nor U3435 (N_3435,N_1575,N_468);
nand U3436 (N_3436,N_382,N_139);
nand U3437 (N_3437,N_958,N_1402);
xnor U3438 (N_3438,N_675,N_314);
or U3439 (N_3439,N_1526,N_1507);
or U3440 (N_3440,N_1755,N_841);
and U3441 (N_3441,N_1014,N_68);
or U3442 (N_3442,N_1594,N_1989);
or U3443 (N_3443,N_1912,N_263);
or U3444 (N_3444,N_1490,N_827);
or U3445 (N_3445,N_331,N_1636);
nand U3446 (N_3446,N_925,N_2197);
and U3447 (N_3447,N_788,N_1908);
nand U3448 (N_3448,N_1793,N_1837);
and U3449 (N_3449,N_589,N_1709);
and U3450 (N_3450,N_732,N_436);
nand U3451 (N_3451,N_935,N_1226);
or U3452 (N_3452,N_650,N_2475);
and U3453 (N_3453,N_387,N_2386);
and U3454 (N_3454,N_590,N_2425);
and U3455 (N_3455,N_845,N_605);
or U3456 (N_3456,N_2091,N_2174);
nand U3457 (N_3457,N_1533,N_377);
and U3458 (N_3458,N_917,N_46);
or U3459 (N_3459,N_2382,N_2352);
and U3460 (N_3460,N_1652,N_319);
xor U3461 (N_3461,N_636,N_1403);
and U3462 (N_3462,N_2094,N_883);
and U3463 (N_3463,N_469,N_1723);
nor U3464 (N_3464,N_1007,N_1294);
and U3465 (N_3465,N_780,N_941);
and U3466 (N_3466,N_1972,N_1096);
xnor U3467 (N_3467,N_596,N_646);
or U3468 (N_3468,N_749,N_818);
nand U3469 (N_3469,N_1779,N_1862);
and U3470 (N_3470,N_2221,N_147);
xnor U3471 (N_3471,N_1077,N_2397);
nand U3472 (N_3472,N_953,N_1119);
or U3473 (N_3473,N_892,N_422);
xnor U3474 (N_3474,N_2095,N_912);
nor U3475 (N_3475,N_2320,N_1484);
xor U3476 (N_3476,N_233,N_700);
or U3477 (N_3477,N_1822,N_1232);
xnor U3478 (N_3478,N_341,N_317);
nor U3479 (N_3479,N_2195,N_1260);
nor U3480 (N_3480,N_666,N_473);
nand U3481 (N_3481,N_1980,N_251);
or U3482 (N_3482,N_786,N_1937);
nor U3483 (N_3483,N_1757,N_723);
xor U3484 (N_3484,N_228,N_1061);
and U3485 (N_3485,N_2032,N_2394);
nor U3486 (N_3486,N_1008,N_854);
xnor U3487 (N_3487,N_1739,N_2124);
or U3488 (N_3488,N_1662,N_2164);
nand U3489 (N_3489,N_1414,N_1334);
xor U3490 (N_3490,N_501,N_1288);
nor U3491 (N_3491,N_1176,N_696);
or U3492 (N_3492,N_521,N_1438);
or U3493 (N_3493,N_2103,N_903);
xor U3494 (N_3494,N_2314,N_614);
or U3495 (N_3495,N_694,N_2074);
nand U3496 (N_3496,N_1742,N_667);
nor U3497 (N_3497,N_243,N_2163);
nand U3498 (N_3498,N_904,N_1450);
or U3499 (N_3499,N_2270,N_1301);
nor U3500 (N_3500,N_1206,N_1666);
nand U3501 (N_3501,N_1336,N_375);
or U3502 (N_3502,N_2044,N_1916);
nor U3503 (N_3503,N_564,N_1072);
xnor U3504 (N_3504,N_1877,N_642);
nor U3505 (N_3505,N_2313,N_1726);
nor U3506 (N_3506,N_152,N_545);
nor U3507 (N_3507,N_1981,N_755);
nor U3508 (N_3508,N_407,N_516);
nand U3509 (N_3509,N_250,N_379);
and U3510 (N_3510,N_284,N_885);
nand U3511 (N_3511,N_1453,N_320);
and U3512 (N_3512,N_2376,N_797);
nor U3513 (N_3513,N_2370,N_512);
and U3514 (N_3514,N_931,N_1883);
nand U3515 (N_3515,N_2156,N_2275);
nor U3516 (N_3516,N_2469,N_1207);
or U3517 (N_3517,N_1379,N_601);
xnor U3518 (N_3518,N_2231,N_872);
nor U3519 (N_3519,N_413,N_1555);
nor U3520 (N_3520,N_274,N_2018);
nand U3521 (N_3521,N_1445,N_2473);
and U3522 (N_3522,N_2467,N_1934);
nor U3523 (N_3523,N_1170,N_861);
or U3524 (N_3524,N_1269,N_2122);
or U3525 (N_3525,N_1369,N_1601);
nor U3526 (N_3526,N_226,N_565);
or U3527 (N_3527,N_1024,N_1047);
nand U3528 (N_3528,N_2458,N_2199);
nor U3529 (N_3529,N_1123,N_132);
and U3530 (N_3530,N_1712,N_915);
nor U3531 (N_3531,N_2350,N_2260);
and U3532 (N_3532,N_1629,N_1017);
and U3533 (N_3533,N_1262,N_1010);
nand U3534 (N_3534,N_1838,N_858);
or U3535 (N_3535,N_1649,N_332);
xor U3536 (N_3536,N_395,N_570);
or U3537 (N_3537,N_887,N_623);
nand U3538 (N_3538,N_1696,N_1161);
nand U3539 (N_3539,N_1370,N_41);
and U3540 (N_3540,N_689,N_529);
or U3541 (N_3541,N_254,N_1095);
nand U3542 (N_3542,N_2298,N_353);
xnor U3543 (N_3543,N_1668,N_19);
xor U3544 (N_3544,N_647,N_980);
nor U3545 (N_3545,N_1513,N_1384);
nor U3546 (N_3546,N_447,N_1648);
nor U3547 (N_3547,N_965,N_2055);
nand U3548 (N_3548,N_638,N_633);
and U3549 (N_3549,N_227,N_1140);
xor U3550 (N_3550,N_402,N_23);
nor U3551 (N_3551,N_156,N_906);
nor U3552 (N_3552,N_586,N_939);
nand U3553 (N_3553,N_120,N_1602);
xnor U3554 (N_3554,N_2465,N_901);
nand U3555 (N_3555,N_992,N_1859);
nor U3556 (N_3556,N_179,N_1133);
and U3557 (N_3557,N_1945,N_1440);
or U3558 (N_3558,N_1899,N_370);
nor U3559 (N_3559,N_708,N_964);
and U3560 (N_3560,N_149,N_1154);
nor U3561 (N_3561,N_1470,N_1204);
or U3562 (N_3562,N_1478,N_2191);
nor U3563 (N_3563,N_1380,N_1504);
and U3564 (N_3564,N_55,N_1197);
or U3565 (N_3565,N_411,N_1982);
xor U3566 (N_3566,N_812,N_346);
or U3567 (N_3567,N_1093,N_2305);
or U3568 (N_3568,N_591,N_181);
or U3569 (N_3569,N_1026,N_2480);
xor U3570 (N_3570,N_1030,N_1966);
xor U3571 (N_3571,N_153,N_630);
or U3572 (N_3572,N_1861,N_92);
or U3573 (N_3573,N_1177,N_2456);
xor U3574 (N_3574,N_2395,N_1661);
nand U3575 (N_3575,N_1348,N_1622);
and U3576 (N_3576,N_2248,N_1693);
and U3577 (N_3577,N_2193,N_1514);
or U3578 (N_3578,N_1574,N_495);
xnor U3579 (N_3579,N_32,N_1298);
xor U3580 (N_3580,N_2139,N_488);
and U3581 (N_3581,N_1239,N_1585);
xnor U3582 (N_3582,N_2075,N_1876);
nor U3583 (N_3583,N_767,N_1421);
nor U3584 (N_3584,N_453,N_607);
or U3585 (N_3585,N_9,N_2184);
nand U3586 (N_3586,N_1994,N_832);
nor U3587 (N_3587,N_255,N_2393);
or U3588 (N_3588,N_1002,N_1821);
or U3589 (N_3589,N_1146,N_1542);
nor U3590 (N_3590,N_649,N_381);
xnor U3591 (N_3591,N_1454,N_2381);
and U3592 (N_3592,N_56,N_1281);
xor U3593 (N_3593,N_78,N_1534);
and U3594 (N_3594,N_688,N_1460);
nand U3595 (N_3595,N_1854,N_1809);
nor U3596 (N_3596,N_2035,N_1725);
and U3597 (N_3597,N_2444,N_2454);
or U3598 (N_3598,N_672,N_2080);
nand U3599 (N_3599,N_888,N_49);
nor U3600 (N_3600,N_1783,N_33);
nor U3601 (N_3601,N_2485,N_2053);
nand U3602 (N_3602,N_290,N_1099);
nand U3603 (N_3603,N_2319,N_2377);
or U3604 (N_3604,N_2489,N_2201);
nand U3605 (N_3605,N_938,N_384);
xnor U3606 (N_3606,N_2287,N_1884);
nand U3607 (N_3607,N_518,N_244);
nor U3608 (N_3608,N_1485,N_972);
nand U3609 (N_3609,N_685,N_771);
nor U3610 (N_3610,N_803,N_91);
xor U3611 (N_3611,N_2351,N_2295);
xor U3612 (N_3612,N_1617,N_1221);
or U3613 (N_3613,N_779,N_1801);
nand U3614 (N_3614,N_385,N_117);
or U3615 (N_3615,N_1291,N_1367);
xnor U3616 (N_3616,N_1205,N_204);
nand U3617 (N_3617,N_421,N_202);
nand U3618 (N_3618,N_2463,N_313);
and U3619 (N_3619,N_2325,N_95);
nand U3620 (N_3620,N_1692,N_981);
nand U3621 (N_3621,N_1758,N_1400);
nor U3622 (N_3622,N_2085,N_1363);
xor U3623 (N_3623,N_432,N_1330);
nand U3624 (N_3624,N_2198,N_2446);
nand U3625 (N_3625,N_1094,N_2408);
nor U3626 (N_3626,N_329,N_1495);
and U3627 (N_3627,N_88,N_61);
xor U3628 (N_3628,N_2033,N_1848);
xor U3629 (N_3629,N_946,N_1220);
nor U3630 (N_3630,N_8,N_1318);
nor U3631 (N_3631,N_371,N_1949);
nand U3632 (N_3632,N_1632,N_237);
xnor U3633 (N_3633,N_1125,N_2335);
nor U3634 (N_3634,N_1129,N_1175);
xor U3635 (N_3635,N_629,N_707);
or U3636 (N_3636,N_717,N_1442);
nand U3637 (N_3637,N_864,N_2317);
or U3638 (N_3638,N_297,N_581);
or U3639 (N_3639,N_1718,N_460);
or U3640 (N_3640,N_1977,N_2027);
nor U3641 (N_3641,N_2348,N_481);
xor U3642 (N_3642,N_796,N_1613);
nor U3643 (N_3643,N_504,N_2438);
or U3644 (N_3644,N_2330,N_2072);
nor U3645 (N_3645,N_2148,N_439);
nor U3646 (N_3646,N_183,N_1082);
xnor U3647 (N_3647,N_1027,N_2254);
and U3648 (N_3648,N_1020,N_704);
xnor U3649 (N_3649,N_515,N_2237);
nor U3650 (N_3650,N_1346,N_1192);
nand U3651 (N_3651,N_768,N_2037);
nand U3652 (N_3652,N_2009,N_406);
and U3653 (N_3653,N_14,N_2001);
nor U3654 (N_3654,N_1736,N_1323);
or U3655 (N_3655,N_472,N_852);
xor U3656 (N_3656,N_1781,N_1304);
nor U3657 (N_3657,N_1254,N_2110);
and U3658 (N_3658,N_1954,N_815);
and U3659 (N_3659,N_2266,N_693);
xor U3660 (N_3660,N_366,N_716);
or U3661 (N_3661,N_493,N_952);
nand U3662 (N_3662,N_1127,N_639);
xor U3663 (N_3663,N_487,N_1075);
nand U3664 (N_3664,N_240,N_1731);
nor U3665 (N_3665,N_618,N_1035);
xnor U3666 (N_3666,N_1794,N_247);
xor U3667 (N_3667,N_315,N_2233);
or U3668 (N_3668,N_719,N_457);
xnor U3669 (N_3669,N_378,N_2200);
nand U3670 (N_3670,N_922,N_71);
nand U3671 (N_3671,N_1646,N_985);
nor U3672 (N_3672,N_789,N_15);
or U3673 (N_3673,N_1447,N_2138);
and U3674 (N_3674,N_913,N_1711);
nand U3675 (N_3675,N_1276,N_1481);
nor U3676 (N_3676,N_882,N_1599);
and U3677 (N_3677,N_1115,N_2041);
nand U3678 (N_3678,N_2177,N_206);
and U3679 (N_3679,N_1566,N_1264);
nand U3680 (N_3680,N_157,N_1335);
and U3681 (N_3681,N_1987,N_1210);
nand U3682 (N_3682,N_1567,N_1201);
nor U3683 (N_3683,N_1703,N_1245);
nand U3684 (N_3684,N_108,N_1634);
xor U3685 (N_3685,N_1737,N_109);
nor U3686 (N_3686,N_1242,N_1550);
nand U3687 (N_3687,N_2359,N_731);
or U3688 (N_3688,N_498,N_1001);
xnor U3689 (N_3689,N_1102,N_221);
nor U3690 (N_3690,N_851,N_1508);
xor U3691 (N_3691,N_1386,N_1277);
or U3692 (N_3692,N_960,N_114);
and U3693 (N_3693,N_1313,N_2474);
and U3694 (N_3694,N_1360,N_304);
and U3695 (N_3695,N_1785,N_535);
nand U3696 (N_3696,N_2114,N_2262);
or U3697 (N_3697,N_813,N_2399);
nand U3698 (N_3698,N_1157,N_197);
nand U3699 (N_3699,N_1374,N_2420);
and U3700 (N_3700,N_921,N_2498);
nor U3701 (N_3701,N_85,N_163);
nand U3702 (N_3702,N_37,N_2400);
or U3703 (N_3703,N_2038,N_644);
xor U3704 (N_3704,N_1405,N_1480);
nand U3705 (N_3705,N_662,N_1108);
nor U3706 (N_3706,N_1524,N_2312);
nand U3707 (N_3707,N_1519,N_1344);
nor U3708 (N_3708,N_2087,N_1673);
nand U3709 (N_3709,N_783,N_2117);
or U3710 (N_3710,N_954,N_1875);
and U3711 (N_3711,N_1874,N_1499);
nand U3712 (N_3712,N_1765,N_1706);
and U3713 (N_3713,N_634,N_1995);
or U3714 (N_3714,N_1287,N_1263);
or U3715 (N_3715,N_898,N_128);
or U3716 (N_3716,N_2190,N_527);
xnor U3717 (N_3717,N_1834,N_82);
nand U3718 (N_3718,N_1250,N_397);
and U3719 (N_3719,N_531,N_528);
or U3720 (N_3720,N_510,N_311);
or U3721 (N_3721,N_1918,N_1902);
and U3722 (N_3722,N_1943,N_2082);
and U3723 (N_3723,N_2363,N_2388);
xnor U3724 (N_3724,N_1828,N_417);
or U3725 (N_3725,N_485,N_600);
xor U3726 (N_3726,N_838,N_923);
or U3727 (N_3727,N_1425,N_2252);
or U3728 (N_3728,N_2479,N_536);
xor U3729 (N_3729,N_775,N_1643);
or U3730 (N_3730,N_754,N_1625);
or U3731 (N_3731,N_991,N_351);
and U3732 (N_3732,N_2157,N_194);
nor U3733 (N_3733,N_298,N_121);
xnor U3734 (N_3734,N_1580,N_2332);
nor U3735 (N_3735,N_2257,N_658);
and U3736 (N_3736,N_2205,N_418);
xor U3737 (N_3737,N_2279,N_914);
and U3738 (N_3738,N_908,N_2490);
and U3739 (N_3739,N_839,N_272);
nor U3740 (N_3740,N_1497,N_899);
nand U3741 (N_3741,N_165,N_2063);
and U3742 (N_3742,N_1894,N_1979);
or U3743 (N_3743,N_336,N_111);
and U3744 (N_3744,N_2006,N_751);
nor U3745 (N_3745,N_497,N_122);
xor U3746 (N_3746,N_209,N_2281);
nor U3747 (N_3747,N_1469,N_1435);
or U3748 (N_3748,N_1290,N_559);
and U3749 (N_3749,N_1434,N_199);
or U3750 (N_3750,N_1960,N_822);
or U3751 (N_3751,N_1360,N_684);
or U3752 (N_3752,N_1439,N_2374);
nor U3753 (N_3753,N_2447,N_665);
nor U3754 (N_3754,N_85,N_906);
and U3755 (N_3755,N_127,N_1401);
nor U3756 (N_3756,N_1397,N_58);
nand U3757 (N_3757,N_1640,N_372);
nor U3758 (N_3758,N_376,N_1001);
nor U3759 (N_3759,N_1445,N_10);
nor U3760 (N_3760,N_1140,N_2314);
xor U3761 (N_3761,N_829,N_1357);
xor U3762 (N_3762,N_1078,N_2043);
nor U3763 (N_3763,N_2135,N_1315);
or U3764 (N_3764,N_560,N_1173);
nand U3765 (N_3765,N_1460,N_2431);
nor U3766 (N_3766,N_1876,N_2320);
xnor U3767 (N_3767,N_1289,N_1195);
and U3768 (N_3768,N_2212,N_2456);
xnor U3769 (N_3769,N_1132,N_2338);
and U3770 (N_3770,N_818,N_1545);
xor U3771 (N_3771,N_1336,N_204);
nor U3772 (N_3772,N_2252,N_2123);
nor U3773 (N_3773,N_1153,N_932);
and U3774 (N_3774,N_116,N_2299);
or U3775 (N_3775,N_2024,N_1160);
xnor U3776 (N_3776,N_2468,N_1143);
xor U3777 (N_3777,N_896,N_1361);
nor U3778 (N_3778,N_762,N_1143);
nand U3779 (N_3779,N_968,N_672);
nand U3780 (N_3780,N_1986,N_1489);
nor U3781 (N_3781,N_1526,N_1282);
or U3782 (N_3782,N_1448,N_2428);
and U3783 (N_3783,N_645,N_1511);
xnor U3784 (N_3784,N_1899,N_1249);
and U3785 (N_3785,N_507,N_252);
or U3786 (N_3786,N_1046,N_1109);
xnor U3787 (N_3787,N_1571,N_1235);
xnor U3788 (N_3788,N_1987,N_2453);
or U3789 (N_3789,N_2013,N_1760);
and U3790 (N_3790,N_1101,N_2312);
or U3791 (N_3791,N_2216,N_1796);
or U3792 (N_3792,N_841,N_1540);
nor U3793 (N_3793,N_817,N_765);
and U3794 (N_3794,N_1255,N_1224);
and U3795 (N_3795,N_1629,N_1199);
and U3796 (N_3796,N_384,N_1978);
nand U3797 (N_3797,N_677,N_2396);
xnor U3798 (N_3798,N_543,N_1020);
or U3799 (N_3799,N_1830,N_207);
nor U3800 (N_3800,N_463,N_1424);
or U3801 (N_3801,N_1541,N_1027);
and U3802 (N_3802,N_1515,N_1833);
xnor U3803 (N_3803,N_1618,N_1499);
nor U3804 (N_3804,N_2157,N_1096);
or U3805 (N_3805,N_1580,N_2018);
nor U3806 (N_3806,N_2054,N_1072);
and U3807 (N_3807,N_1783,N_103);
or U3808 (N_3808,N_381,N_2211);
xnor U3809 (N_3809,N_1548,N_599);
xor U3810 (N_3810,N_1909,N_546);
nor U3811 (N_3811,N_2489,N_1318);
xnor U3812 (N_3812,N_1160,N_1685);
nand U3813 (N_3813,N_686,N_1757);
xor U3814 (N_3814,N_1116,N_925);
and U3815 (N_3815,N_743,N_1687);
nand U3816 (N_3816,N_1723,N_1870);
xor U3817 (N_3817,N_78,N_2021);
xnor U3818 (N_3818,N_2063,N_642);
and U3819 (N_3819,N_1230,N_2199);
and U3820 (N_3820,N_1037,N_923);
and U3821 (N_3821,N_1674,N_36);
nor U3822 (N_3822,N_2496,N_802);
nand U3823 (N_3823,N_1749,N_30);
nor U3824 (N_3824,N_551,N_388);
nand U3825 (N_3825,N_862,N_717);
xor U3826 (N_3826,N_1669,N_1002);
and U3827 (N_3827,N_2101,N_2346);
xor U3828 (N_3828,N_1739,N_616);
nor U3829 (N_3829,N_180,N_858);
nand U3830 (N_3830,N_200,N_1734);
or U3831 (N_3831,N_126,N_1825);
nor U3832 (N_3832,N_1462,N_2203);
xnor U3833 (N_3833,N_2401,N_1767);
and U3834 (N_3834,N_1411,N_1867);
xnor U3835 (N_3835,N_778,N_668);
nor U3836 (N_3836,N_1785,N_560);
nor U3837 (N_3837,N_1147,N_1086);
and U3838 (N_3838,N_1330,N_339);
and U3839 (N_3839,N_547,N_1078);
nand U3840 (N_3840,N_1848,N_288);
and U3841 (N_3841,N_1383,N_859);
and U3842 (N_3842,N_306,N_1428);
nand U3843 (N_3843,N_1620,N_200);
xnor U3844 (N_3844,N_330,N_951);
xnor U3845 (N_3845,N_1182,N_226);
or U3846 (N_3846,N_1820,N_450);
or U3847 (N_3847,N_1386,N_9);
and U3848 (N_3848,N_790,N_1899);
nor U3849 (N_3849,N_959,N_2152);
nor U3850 (N_3850,N_2149,N_2156);
xor U3851 (N_3851,N_669,N_349);
and U3852 (N_3852,N_2028,N_1495);
and U3853 (N_3853,N_103,N_1953);
and U3854 (N_3854,N_1554,N_883);
and U3855 (N_3855,N_2259,N_372);
xnor U3856 (N_3856,N_350,N_2172);
nor U3857 (N_3857,N_2226,N_1946);
nor U3858 (N_3858,N_1521,N_47);
nor U3859 (N_3859,N_1164,N_504);
xnor U3860 (N_3860,N_1005,N_386);
nand U3861 (N_3861,N_2431,N_283);
nand U3862 (N_3862,N_407,N_2146);
nor U3863 (N_3863,N_597,N_1768);
nand U3864 (N_3864,N_1213,N_781);
xor U3865 (N_3865,N_2276,N_2139);
and U3866 (N_3866,N_1087,N_1528);
and U3867 (N_3867,N_2291,N_181);
xnor U3868 (N_3868,N_2407,N_2175);
xnor U3869 (N_3869,N_458,N_2425);
nand U3870 (N_3870,N_455,N_1424);
xnor U3871 (N_3871,N_142,N_107);
nand U3872 (N_3872,N_2397,N_268);
or U3873 (N_3873,N_627,N_2284);
nor U3874 (N_3874,N_1362,N_402);
and U3875 (N_3875,N_2097,N_1310);
nor U3876 (N_3876,N_1996,N_937);
xor U3877 (N_3877,N_1943,N_1059);
nand U3878 (N_3878,N_518,N_852);
and U3879 (N_3879,N_687,N_1130);
and U3880 (N_3880,N_449,N_969);
or U3881 (N_3881,N_321,N_1475);
nor U3882 (N_3882,N_1798,N_2009);
or U3883 (N_3883,N_1295,N_921);
nand U3884 (N_3884,N_66,N_1486);
xor U3885 (N_3885,N_1206,N_2132);
xor U3886 (N_3886,N_726,N_2171);
or U3887 (N_3887,N_2167,N_1040);
or U3888 (N_3888,N_1984,N_918);
xor U3889 (N_3889,N_1809,N_1559);
nand U3890 (N_3890,N_417,N_267);
or U3891 (N_3891,N_971,N_1916);
nand U3892 (N_3892,N_2298,N_525);
nor U3893 (N_3893,N_2344,N_941);
nand U3894 (N_3894,N_1082,N_2277);
and U3895 (N_3895,N_819,N_2167);
nor U3896 (N_3896,N_579,N_1100);
and U3897 (N_3897,N_1134,N_1069);
nor U3898 (N_3898,N_84,N_2455);
xor U3899 (N_3899,N_2144,N_825);
and U3900 (N_3900,N_2014,N_2280);
nand U3901 (N_3901,N_621,N_933);
and U3902 (N_3902,N_1174,N_1979);
xor U3903 (N_3903,N_1629,N_1941);
nor U3904 (N_3904,N_1406,N_1429);
and U3905 (N_3905,N_889,N_2009);
and U3906 (N_3906,N_1901,N_604);
and U3907 (N_3907,N_361,N_1693);
nor U3908 (N_3908,N_1741,N_828);
or U3909 (N_3909,N_1358,N_215);
and U3910 (N_3910,N_211,N_1955);
nor U3911 (N_3911,N_2482,N_2195);
or U3912 (N_3912,N_1158,N_1951);
nand U3913 (N_3913,N_1327,N_1606);
and U3914 (N_3914,N_556,N_2364);
nor U3915 (N_3915,N_1135,N_1903);
nor U3916 (N_3916,N_2419,N_1230);
or U3917 (N_3917,N_732,N_2190);
nand U3918 (N_3918,N_2238,N_1265);
and U3919 (N_3919,N_398,N_261);
nand U3920 (N_3920,N_2060,N_57);
and U3921 (N_3921,N_106,N_469);
and U3922 (N_3922,N_262,N_465);
xnor U3923 (N_3923,N_278,N_1078);
nand U3924 (N_3924,N_1145,N_603);
nand U3925 (N_3925,N_1413,N_1526);
or U3926 (N_3926,N_1348,N_2355);
or U3927 (N_3927,N_1543,N_613);
and U3928 (N_3928,N_1174,N_299);
nand U3929 (N_3929,N_2379,N_1717);
xnor U3930 (N_3930,N_1849,N_1919);
nor U3931 (N_3931,N_2052,N_1273);
and U3932 (N_3932,N_2026,N_1342);
or U3933 (N_3933,N_782,N_237);
xor U3934 (N_3934,N_2041,N_1466);
nor U3935 (N_3935,N_123,N_183);
or U3936 (N_3936,N_837,N_2165);
and U3937 (N_3937,N_321,N_2163);
or U3938 (N_3938,N_1760,N_1831);
and U3939 (N_3939,N_1524,N_73);
xnor U3940 (N_3940,N_1603,N_1989);
nand U3941 (N_3941,N_343,N_1921);
nor U3942 (N_3942,N_1916,N_2075);
nand U3943 (N_3943,N_1837,N_208);
nor U3944 (N_3944,N_1008,N_1964);
or U3945 (N_3945,N_1767,N_858);
or U3946 (N_3946,N_1147,N_356);
xor U3947 (N_3947,N_297,N_1576);
and U3948 (N_3948,N_2078,N_2338);
or U3949 (N_3949,N_1161,N_1528);
nand U3950 (N_3950,N_1012,N_973);
and U3951 (N_3951,N_1712,N_435);
and U3952 (N_3952,N_1488,N_1638);
and U3953 (N_3953,N_2434,N_1878);
and U3954 (N_3954,N_1788,N_2045);
nor U3955 (N_3955,N_624,N_326);
nand U3956 (N_3956,N_676,N_1873);
and U3957 (N_3957,N_2452,N_1989);
nand U3958 (N_3958,N_279,N_82);
nor U3959 (N_3959,N_2198,N_1388);
xor U3960 (N_3960,N_2407,N_847);
nor U3961 (N_3961,N_1541,N_2360);
and U3962 (N_3962,N_1723,N_2468);
or U3963 (N_3963,N_1175,N_1304);
nor U3964 (N_3964,N_528,N_2177);
nand U3965 (N_3965,N_967,N_598);
xnor U3966 (N_3966,N_121,N_404);
or U3967 (N_3967,N_1810,N_733);
nor U3968 (N_3968,N_2021,N_46);
nand U3969 (N_3969,N_562,N_888);
nand U3970 (N_3970,N_576,N_479);
nand U3971 (N_3971,N_239,N_395);
and U3972 (N_3972,N_1203,N_1748);
and U3973 (N_3973,N_862,N_142);
and U3974 (N_3974,N_2469,N_2361);
or U3975 (N_3975,N_1624,N_282);
or U3976 (N_3976,N_621,N_1994);
xnor U3977 (N_3977,N_1178,N_1991);
nor U3978 (N_3978,N_1995,N_1513);
nand U3979 (N_3979,N_1151,N_1842);
and U3980 (N_3980,N_1237,N_86);
or U3981 (N_3981,N_1971,N_247);
or U3982 (N_3982,N_286,N_1611);
nand U3983 (N_3983,N_1140,N_2373);
or U3984 (N_3984,N_642,N_49);
or U3985 (N_3985,N_398,N_1794);
or U3986 (N_3986,N_2035,N_1164);
xnor U3987 (N_3987,N_306,N_1709);
xor U3988 (N_3988,N_2171,N_700);
and U3989 (N_3989,N_1943,N_1865);
xor U3990 (N_3990,N_945,N_890);
xor U3991 (N_3991,N_913,N_789);
nor U3992 (N_3992,N_2435,N_340);
xnor U3993 (N_3993,N_1971,N_740);
xnor U3994 (N_3994,N_2211,N_1170);
xor U3995 (N_3995,N_213,N_2101);
or U3996 (N_3996,N_1178,N_1916);
or U3997 (N_3997,N_532,N_1561);
or U3998 (N_3998,N_575,N_1398);
nor U3999 (N_3999,N_511,N_1256);
nor U4000 (N_4000,N_1008,N_1990);
nor U4001 (N_4001,N_311,N_2363);
and U4002 (N_4002,N_1514,N_2353);
nand U4003 (N_4003,N_636,N_2325);
xnor U4004 (N_4004,N_1931,N_1569);
xor U4005 (N_4005,N_1398,N_1172);
nor U4006 (N_4006,N_1941,N_1397);
and U4007 (N_4007,N_1258,N_2061);
nand U4008 (N_4008,N_1611,N_150);
nor U4009 (N_4009,N_2137,N_1581);
xnor U4010 (N_4010,N_1882,N_877);
xor U4011 (N_4011,N_2116,N_867);
nor U4012 (N_4012,N_661,N_1446);
and U4013 (N_4013,N_2358,N_1935);
or U4014 (N_4014,N_1427,N_985);
nand U4015 (N_4015,N_1929,N_102);
nand U4016 (N_4016,N_1205,N_2164);
xor U4017 (N_4017,N_1516,N_1166);
nor U4018 (N_4018,N_2180,N_4);
and U4019 (N_4019,N_60,N_1011);
or U4020 (N_4020,N_2498,N_1416);
and U4021 (N_4021,N_757,N_2462);
and U4022 (N_4022,N_1551,N_2197);
nand U4023 (N_4023,N_1015,N_514);
nand U4024 (N_4024,N_795,N_1732);
nand U4025 (N_4025,N_2055,N_1274);
and U4026 (N_4026,N_1584,N_1636);
xor U4027 (N_4027,N_1186,N_1265);
xor U4028 (N_4028,N_30,N_1362);
nand U4029 (N_4029,N_719,N_1254);
or U4030 (N_4030,N_228,N_621);
nor U4031 (N_4031,N_961,N_2096);
and U4032 (N_4032,N_22,N_26);
xor U4033 (N_4033,N_1511,N_2225);
and U4034 (N_4034,N_2312,N_843);
or U4035 (N_4035,N_1268,N_984);
and U4036 (N_4036,N_1812,N_2166);
nand U4037 (N_4037,N_515,N_317);
nand U4038 (N_4038,N_1469,N_714);
nor U4039 (N_4039,N_1459,N_675);
and U4040 (N_4040,N_336,N_174);
or U4041 (N_4041,N_259,N_1754);
xor U4042 (N_4042,N_1669,N_831);
xnor U4043 (N_4043,N_1947,N_22);
nor U4044 (N_4044,N_2251,N_950);
xnor U4045 (N_4045,N_343,N_1121);
nor U4046 (N_4046,N_231,N_2378);
xnor U4047 (N_4047,N_912,N_437);
nor U4048 (N_4048,N_906,N_1329);
and U4049 (N_4049,N_1789,N_68);
and U4050 (N_4050,N_418,N_891);
nor U4051 (N_4051,N_1423,N_1624);
nand U4052 (N_4052,N_1236,N_2454);
xor U4053 (N_4053,N_247,N_1177);
and U4054 (N_4054,N_391,N_604);
and U4055 (N_4055,N_1664,N_1912);
nand U4056 (N_4056,N_1147,N_1236);
or U4057 (N_4057,N_56,N_1363);
nor U4058 (N_4058,N_350,N_2432);
or U4059 (N_4059,N_2184,N_597);
nand U4060 (N_4060,N_1424,N_2069);
nor U4061 (N_4061,N_649,N_966);
xnor U4062 (N_4062,N_1318,N_2056);
xnor U4063 (N_4063,N_1840,N_1924);
nor U4064 (N_4064,N_428,N_1251);
nor U4065 (N_4065,N_1328,N_310);
and U4066 (N_4066,N_2054,N_2094);
or U4067 (N_4067,N_1718,N_617);
xnor U4068 (N_4068,N_87,N_944);
and U4069 (N_4069,N_409,N_1541);
nand U4070 (N_4070,N_1352,N_645);
nor U4071 (N_4071,N_1816,N_227);
nor U4072 (N_4072,N_1040,N_113);
nor U4073 (N_4073,N_1449,N_420);
nor U4074 (N_4074,N_772,N_903);
nor U4075 (N_4075,N_2086,N_490);
nand U4076 (N_4076,N_1134,N_2080);
nand U4077 (N_4077,N_1196,N_77);
nand U4078 (N_4078,N_1422,N_2027);
xnor U4079 (N_4079,N_1808,N_2029);
nor U4080 (N_4080,N_1506,N_67);
xnor U4081 (N_4081,N_1034,N_1946);
nand U4082 (N_4082,N_1368,N_1651);
xor U4083 (N_4083,N_1124,N_809);
nor U4084 (N_4084,N_138,N_2006);
xnor U4085 (N_4085,N_1173,N_342);
nand U4086 (N_4086,N_439,N_2302);
and U4087 (N_4087,N_1796,N_471);
and U4088 (N_4088,N_62,N_1336);
and U4089 (N_4089,N_2050,N_411);
nand U4090 (N_4090,N_671,N_88);
xnor U4091 (N_4091,N_2493,N_1836);
xor U4092 (N_4092,N_1762,N_142);
or U4093 (N_4093,N_1544,N_527);
nor U4094 (N_4094,N_359,N_2430);
xor U4095 (N_4095,N_2279,N_149);
and U4096 (N_4096,N_1720,N_2335);
xor U4097 (N_4097,N_2347,N_644);
or U4098 (N_4098,N_812,N_313);
xnor U4099 (N_4099,N_1659,N_1047);
and U4100 (N_4100,N_540,N_428);
nand U4101 (N_4101,N_933,N_958);
nand U4102 (N_4102,N_1155,N_968);
and U4103 (N_4103,N_2319,N_1654);
or U4104 (N_4104,N_500,N_948);
or U4105 (N_4105,N_586,N_1810);
xor U4106 (N_4106,N_20,N_144);
or U4107 (N_4107,N_1528,N_1075);
nor U4108 (N_4108,N_144,N_1320);
nor U4109 (N_4109,N_2027,N_1337);
nand U4110 (N_4110,N_1272,N_638);
nand U4111 (N_4111,N_180,N_1262);
xnor U4112 (N_4112,N_1993,N_1693);
nor U4113 (N_4113,N_1565,N_1313);
and U4114 (N_4114,N_1053,N_632);
nand U4115 (N_4115,N_1971,N_1100);
or U4116 (N_4116,N_28,N_1427);
nor U4117 (N_4117,N_2183,N_720);
or U4118 (N_4118,N_1404,N_459);
xnor U4119 (N_4119,N_2367,N_1753);
nand U4120 (N_4120,N_1042,N_678);
and U4121 (N_4121,N_1634,N_1630);
or U4122 (N_4122,N_2388,N_2297);
nor U4123 (N_4123,N_1236,N_1028);
and U4124 (N_4124,N_2414,N_1251);
nor U4125 (N_4125,N_1180,N_2318);
nor U4126 (N_4126,N_2499,N_219);
xnor U4127 (N_4127,N_1590,N_2063);
and U4128 (N_4128,N_2036,N_105);
nor U4129 (N_4129,N_1044,N_324);
and U4130 (N_4130,N_2192,N_1564);
or U4131 (N_4131,N_695,N_400);
xnor U4132 (N_4132,N_2040,N_1254);
nand U4133 (N_4133,N_84,N_970);
xnor U4134 (N_4134,N_1442,N_675);
nand U4135 (N_4135,N_15,N_246);
and U4136 (N_4136,N_944,N_1119);
and U4137 (N_4137,N_1111,N_1203);
xor U4138 (N_4138,N_2399,N_1414);
xnor U4139 (N_4139,N_1216,N_1704);
and U4140 (N_4140,N_1696,N_1846);
and U4141 (N_4141,N_2492,N_732);
nor U4142 (N_4142,N_367,N_24);
and U4143 (N_4143,N_1972,N_1498);
nand U4144 (N_4144,N_2345,N_760);
nand U4145 (N_4145,N_1503,N_575);
or U4146 (N_4146,N_1617,N_102);
nor U4147 (N_4147,N_422,N_1782);
nand U4148 (N_4148,N_310,N_195);
xor U4149 (N_4149,N_1207,N_80);
nand U4150 (N_4150,N_1545,N_584);
nor U4151 (N_4151,N_18,N_906);
or U4152 (N_4152,N_2232,N_1699);
and U4153 (N_4153,N_104,N_2449);
and U4154 (N_4154,N_781,N_2353);
and U4155 (N_4155,N_712,N_722);
nor U4156 (N_4156,N_137,N_1901);
and U4157 (N_4157,N_615,N_1418);
nor U4158 (N_4158,N_538,N_1811);
and U4159 (N_4159,N_2301,N_841);
and U4160 (N_4160,N_1032,N_384);
and U4161 (N_4161,N_586,N_1137);
xor U4162 (N_4162,N_1737,N_856);
nand U4163 (N_4163,N_1656,N_788);
nand U4164 (N_4164,N_593,N_2123);
and U4165 (N_4165,N_44,N_1658);
xor U4166 (N_4166,N_1052,N_2290);
and U4167 (N_4167,N_1448,N_885);
nor U4168 (N_4168,N_954,N_1192);
xor U4169 (N_4169,N_1710,N_836);
nand U4170 (N_4170,N_631,N_1479);
nand U4171 (N_4171,N_267,N_194);
or U4172 (N_4172,N_101,N_282);
or U4173 (N_4173,N_2373,N_406);
nor U4174 (N_4174,N_1413,N_2033);
and U4175 (N_4175,N_2061,N_1575);
xnor U4176 (N_4176,N_1618,N_214);
or U4177 (N_4177,N_346,N_1671);
and U4178 (N_4178,N_1859,N_671);
xor U4179 (N_4179,N_796,N_1118);
xnor U4180 (N_4180,N_1428,N_89);
nor U4181 (N_4181,N_1017,N_968);
and U4182 (N_4182,N_2020,N_2462);
or U4183 (N_4183,N_978,N_1632);
xor U4184 (N_4184,N_2324,N_933);
xnor U4185 (N_4185,N_2140,N_1993);
and U4186 (N_4186,N_545,N_2333);
and U4187 (N_4187,N_650,N_651);
or U4188 (N_4188,N_1151,N_324);
xnor U4189 (N_4189,N_2265,N_1082);
xor U4190 (N_4190,N_388,N_443);
nand U4191 (N_4191,N_2399,N_641);
and U4192 (N_4192,N_1264,N_1551);
nand U4193 (N_4193,N_778,N_1966);
nand U4194 (N_4194,N_2442,N_1076);
nand U4195 (N_4195,N_0,N_1177);
and U4196 (N_4196,N_804,N_892);
nand U4197 (N_4197,N_638,N_1279);
nor U4198 (N_4198,N_2010,N_1132);
and U4199 (N_4199,N_898,N_2049);
and U4200 (N_4200,N_99,N_1711);
nor U4201 (N_4201,N_2383,N_2082);
nand U4202 (N_4202,N_277,N_1177);
and U4203 (N_4203,N_2154,N_569);
nor U4204 (N_4204,N_1978,N_1650);
nor U4205 (N_4205,N_812,N_59);
nand U4206 (N_4206,N_214,N_924);
nor U4207 (N_4207,N_2058,N_2436);
or U4208 (N_4208,N_505,N_1976);
nor U4209 (N_4209,N_570,N_498);
xor U4210 (N_4210,N_1028,N_1751);
nor U4211 (N_4211,N_2346,N_584);
and U4212 (N_4212,N_1919,N_647);
and U4213 (N_4213,N_2233,N_763);
nand U4214 (N_4214,N_2275,N_57);
nand U4215 (N_4215,N_1918,N_2305);
and U4216 (N_4216,N_1454,N_860);
nand U4217 (N_4217,N_1905,N_1686);
nor U4218 (N_4218,N_1056,N_1172);
or U4219 (N_4219,N_1939,N_390);
or U4220 (N_4220,N_1761,N_2154);
nand U4221 (N_4221,N_2255,N_1918);
nand U4222 (N_4222,N_1259,N_1192);
nor U4223 (N_4223,N_1375,N_1395);
or U4224 (N_4224,N_1002,N_1817);
xor U4225 (N_4225,N_1838,N_1313);
xnor U4226 (N_4226,N_761,N_1658);
nor U4227 (N_4227,N_1542,N_1736);
or U4228 (N_4228,N_1437,N_1280);
or U4229 (N_4229,N_1360,N_929);
and U4230 (N_4230,N_76,N_396);
nand U4231 (N_4231,N_1105,N_24);
nand U4232 (N_4232,N_880,N_786);
nor U4233 (N_4233,N_1573,N_2378);
nor U4234 (N_4234,N_2412,N_669);
and U4235 (N_4235,N_663,N_1144);
nor U4236 (N_4236,N_2229,N_1711);
and U4237 (N_4237,N_2031,N_1088);
nand U4238 (N_4238,N_672,N_827);
or U4239 (N_4239,N_830,N_1164);
or U4240 (N_4240,N_1502,N_2172);
nand U4241 (N_4241,N_733,N_1459);
and U4242 (N_4242,N_988,N_1211);
and U4243 (N_4243,N_856,N_555);
and U4244 (N_4244,N_326,N_628);
xor U4245 (N_4245,N_1367,N_191);
xor U4246 (N_4246,N_108,N_1374);
xnor U4247 (N_4247,N_1740,N_1311);
nand U4248 (N_4248,N_618,N_1211);
or U4249 (N_4249,N_1338,N_526);
and U4250 (N_4250,N_1078,N_2177);
or U4251 (N_4251,N_555,N_802);
nor U4252 (N_4252,N_2363,N_1602);
or U4253 (N_4253,N_1621,N_2094);
nor U4254 (N_4254,N_1933,N_2239);
nand U4255 (N_4255,N_959,N_1272);
or U4256 (N_4256,N_395,N_2477);
or U4257 (N_4257,N_527,N_566);
xnor U4258 (N_4258,N_1558,N_1536);
nor U4259 (N_4259,N_1008,N_1486);
xor U4260 (N_4260,N_635,N_1068);
nor U4261 (N_4261,N_994,N_289);
or U4262 (N_4262,N_1450,N_27);
or U4263 (N_4263,N_2473,N_241);
or U4264 (N_4264,N_2208,N_2387);
or U4265 (N_4265,N_860,N_581);
or U4266 (N_4266,N_2240,N_1837);
or U4267 (N_4267,N_510,N_229);
nor U4268 (N_4268,N_122,N_1265);
and U4269 (N_4269,N_1140,N_27);
or U4270 (N_4270,N_2221,N_37);
xor U4271 (N_4271,N_1385,N_2334);
and U4272 (N_4272,N_1509,N_1452);
nor U4273 (N_4273,N_420,N_1200);
or U4274 (N_4274,N_5,N_1150);
and U4275 (N_4275,N_648,N_1398);
or U4276 (N_4276,N_405,N_1111);
xor U4277 (N_4277,N_465,N_404);
or U4278 (N_4278,N_268,N_1042);
nand U4279 (N_4279,N_1650,N_1932);
and U4280 (N_4280,N_1663,N_878);
nor U4281 (N_4281,N_1786,N_1875);
xnor U4282 (N_4282,N_608,N_612);
xor U4283 (N_4283,N_2476,N_1062);
or U4284 (N_4284,N_7,N_1135);
xor U4285 (N_4285,N_2315,N_2159);
nor U4286 (N_4286,N_1389,N_971);
xnor U4287 (N_4287,N_1742,N_1510);
nor U4288 (N_4288,N_2311,N_1286);
nand U4289 (N_4289,N_1932,N_1955);
xnor U4290 (N_4290,N_347,N_1750);
xor U4291 (N_4291,N_1082,N_1742);
nor U4292 (N_4292,N_205,N_1882);
nand U4293 (N_4293,N_228,N_105);
nor U4294 (N_4294,N_101,N_415);
nor U4295 (N_4295,N_893,N_2098);
xnor U4296 (N_4296,N_729,N_1305);
xor U4297 (N_4297,N_1461,N_347);
or U4298 (N_4298,N_1769,N_2082);
nor U4299 (N_4299,N_386,N_1392);
xnor U4300 (N_4300,N_1565,N_2352);
nor U4301 (N_4301,N_190,N_400);
or U4302 (N_4302,N_2461,N_1111);
and U4303 (N_4303,N_106,N_504);
and U4304 (N_4304,N_544,N_281);
nor U4305 (N_4305,N_1143,N_315);
or U4306 (N_4306,N_2019,N_886);
nor U4307 (N_4307,N_1798,N_843);
nor U4308 (N_4308,N_1389,N_1699);
nand U4309 (N_4309,N_741,N_1496);
nand U4310 (N_4310,N_948,N_1764);
and U4311 (N_4311,N_1751,N_2200);
nor U4312 (N_4312,N_88,N_1765);
nand U4313 (N_4313,N_1602,N_978);
xor U4314 (N_4314,N_1291,N_55);
or U4315 (N_4315,N_2180,N_1272);
nor U4316 (N_4316,N_1596,N_2463);
and U4317 (N_4317,N_1141,N_1556);
xor U4318 (N_4318,N_1,N_1968);
and U4319 (N_4319,N_2350,N_2225);
and U4320 (N_4320,N_1647,N_1846);
nand U4321 (N_4321,N_726,N_397);
or U4322 (N_4322,N_899,N_1684);
and U4323 (N_4323,N_2156,N_1572);
and U4324 (N_4324,N_310,N_1489);
nand U4325 (N_4325,N_2022,N_23);
or U4326 (N_4326,N_710,N_452);
xor U4327 (N_4327,N_289,N_1271);
nor U4328 (N_4328,N_1320,N_152);
and U4329 (N_4329,N_474,N_1251);
xnor U4330 (N_4330,N_2075,N_1864);
nand U4331 (N_4331,N_1996,N_1438);
xor U4332 (N_4332,N_1044,N_2096);
nor U4333 (N_4333,N_865,N_1086);
xor U4334 (N_4334,N_1796,N_2154);
nand U4335 (N_4335,N_1661,N_2379);
nand U4336 (N_4336,N_866,N_1735);
xor U4337 (N_4337,N_275,N_2333);
or U4338 (N_4338,N_458,N_1985);
xnor U4339 (N_4339,N_1320,N_873);
nor U4340 (N_4340,N_574,N_1981);
nor U4341 (N_4341,N_584,N_780);
xor U4342 (N_4342,N_285,N_1041);
nor U4343 (N_4343,N_2135,N_1827);
nor U4344 (N_4344,N_617,N_1829);
xnor U4345 (N_4345,N_739,N_2015);
or U4346 (N_4346,N_2354,N_1980);
xnor U4347 (N_4347,N_1485,N_956);
or U4348 (N_4348,N_7,N_1752);
nor U4349 (N_4349,N_2119,N_1821);
nand U4350 (N_4350,N_2271,N_118);
nor U4351 (N_4351,N_664,N_1937);
nor U4352 (N_4352,N_2295,N_1934);
or U4353 (N_4353,N_2412,N_693);
or U4354 (N_4354,N_692,N_2374);
and U4355 (N_4355,N_34,N_1119);
nand U4356 (N_4356,N_2104,N_2378);
xnor U4357 (N_4357,N_1379,N_699);
or U4358 (N_4358,N_892,N_146);
nor U4359 (N_4359,N_2416,N_96);
and U4360 (N_4360,N_874,N_1162);
and U4361 (N_4361,N_2064,N_1511);
nor U4362 (N_4362,N_2358,N_927);
and U4363 (N_4363,N_2378,N_222);
and U4364 (N_4364,N_391,N_1120);
nor U4365 (N_4365,N_1149,N_1274);
or U4366 (N_4366,N_2486,N_1559);
nand U4367 (N_4367,N_1265,N_699);
nor U4368 (N_4368,N_913,N_1033);
and U4369 (N_4369,N_616,N_0);
xor U4370 (N_4370,N_2144,N_1690);
and U4371 (N_4371,N_1994,N_195);
nor U4372 (N_4372,N_1218,N_2338);
or U4373 (N_4373,N_2420,N_2301);
xor U4374 (N_4374,N_547,N_1507);
nand U4375 (N_4375,N_1561,N_2282);
or U4376 (N_4376,N_1897,N_738);
nand U4377 (N_4377,N_2269,N_2427);
nand U4378 (N_4378,N_433,N_1074);
nor U4379 (N_4379,N_2320,N_457);
xor U4380 (N_4380,N_112,N_1554);
nand U4381 (N_4381,N_451,N_2345);
and U4382 (N_4382,N_375,N_1874);
nor U4383 (N_4383,N_806,N_1133);
or U4384 (N_4384,N_432,N_411);
nand U4385 (N_4385,N_1025,N_877);
or U4386 (N_4386,N_1636,N_473);
xor U4387 (N_4387,N_188,N_1645);
xor U4388 (N_4388,N_121,N_1902);
or U4389 (N_4389,N_1121,N_1998);
nand U4390 (N_4390,N_1875,N_415);
and U4391 (N_4391,N_2239,N_1034);
xnor U4392 (N_4392,N_760,N_1378);
and U4393 (N_4393,N_360,N_697);
xor U4394 (N_4394,N_714,N_2317);
nor U4395 (N_4395,N_206,N_1717);
and U4396 (N_4396,N_801,N_1854);
xor U4397 (N_4397,N_1354,N_1268);
xor U4398 (N_4398,N_170,N_249);
or U4399 (N_4399,N_2210,N_1071);
nand U4400 (N_4400,N_1157,N_420);
and U4401 (N_4401,N_1886,N_797);
xor U4402 (N_4402,N_714,N_1474);
xnor U4403 (N_4403,N_283,N_1124);
or U4404 (N_4404,N_233,N_1870);
or U4405 (N_4405,N_1231,N_1292);
and U4406 (N_4406,N_1233,N_1545);
and U4407 (N_4407,N_2259,N_1775);
nor U4408 (N_4408,N_620,N_1688);
xor U4409 (N_4409,N_1592,N_1206);
and U4410 (N_4410,N_2045,N_2353);
nor U4411 (N_4411,N_1356,N_1511);
nand U4412 (N_4412,N_1185,N_1926);
xnor U4413 (N_4413,N_2356,N_547);
nand U4414 (N_4414,N_1275,N_1524);
nand U4415 (N_4415,N_1346,N_1647);
nand U4416 (N_4416,N_2478,N_756);
and U4417 (N_4417,N_391,N_394);
or U4418 (N_4418,N_973,N_2132);
nand U4419 (N_4419,N_180,N_1327);
xor U4420 (N_4420,N_1526,N_686);
nand U4421 (N_4421,N_455,N_1518);
xnor U4422 (N_4422,N_1557,N_1252);
and U4423 (N_4423,N_2423,N_1658);
xor U4424 (N_4424,N_78,N_825);
nand U4425 (N_4425,N_1561,N_206);
xor U4426 (N_4426,N_2071,N_2437);
xnor U4427 (N_4427,N_698,N_2298);
or U4428 (N_4428,N_353,N_1349);
and U4429 (N_4429,N_443,N_1153);
nor U4430 (N_4430,N_1028,N_1143);
xor U4431 (N_4431,N_1143,N_498);
and U4432 (N_4432,N_2402,N_1358);
nand U4433 (N_4433,N_1546,N_1072);
nor U4434 (N_4434,N_1477,N_2449);
xnor U4435 (N_4435,N_2376,N_494);
nand U4436 (N_4436,N_1834,N_1622);
nand U4437 (N_4437,N_2162,N_472);
and U4438 (N_4438,N_795,N_23);
xor U4439 (N_4439,N_744,N_1402);
xor U4440 (N_4440,N_1534,N_1552);
nand U4441 (N_4441,N_1594,N_1189);
nor U4442 (N_4442,N_789,N_1109);
xor U4443 (N_4443,N_1693,N_1617);
and U4444 (N_4444,N_1646,N_2244);
xor U4445 (N_4445,N_1534,N_2165);
and U4446 (N_4446,N_201,N_1613);
or U4447 (N_4447,N_1775,N_566);
nor U4448 (N_4448,N_2345,N_2236);
nand U4449 (N_4449,N_1136,N_1386);
xnor U4450 (N_4450,N_315,N_568);
xnor U4451 (N_4451,N_2496,N_558);
nand U4452 (N_4452,N_2380,N_1651);
or U4453 (N_4453,N_854,N_2115);
nand U4454 (N_4454,N_1011,N_636);
or U4455 (N_4455,N_1488,N_856);
or U4456 (N_4456,N_2395,N_373);
nand U4457 (N_4457,N_960,N_925);
nand U4458 (N_4458,N_1870,N_551);
or U4459 (N_4459,N_118,N_657);
nand U4460 (N_4460,N_1925,N_1672);
or U4461 (N_4461,N_1436,N_1622);
nand U4462 (N_4462,N_1459,N_1658);
nand U4463 (N_4463,N_294,N_1933);
or U4464 (N_4464,N_2342,N_1749);
nand U4465 (N_4465,N_1672,N_1623);
xor U4466 (N_4466,N_1035,N_151);
or U4467 (N_4467,N_46,N_183);
xor U4468 (N_4468,N_839,N_1486);
and U4469 (N_4469,N_2385,N_462);
nor U4470 (N_4470,N_2344,N_1794);
xor U4471 (N_4471,N_231,N_1203);
nor U4472 (N_4472,N_1939,N_2262);
and U4473 (N_4473,N_1385,N_1138);
nand U4474 (N_4474,N_1618,N_2202);
or U4475 (N_4475,N_599,N_1387);
xor U4476 (N_4476,N_1933,N_417);
nand U4477 (N_4477,N_2220,N_798);
or U4478 (N_4478,N_2004,N_2267);
nor U4479 (N_4479,N_2117,N_998);
or U4480 (N_4480,N_2364,N_1745);
nand U4481 (N_4481,N_1961,N_91);
or U4482 (N_4482,N_2072,N_1048);
or U4483 (N_4483,N_1084,N_1189);
and U4484 (N_4484,N_1452,N_880);
nor U4485 (N_4485,N_1436,N_1404);
nor U4486 (N_4486,N_1596,N_626);
or U4487 (N_4487,N_2128,N_1068);
and U4488 (N_4488,N_1534,N_768);
and U4489 (N_4489,N_2274,N_1588);
nor U4490 (N_4490,N_2410,N_73);
nor U4491 (N_4491,N_1005,N_2428);
and U4492 (N_4492,N_833,N_1070);
and U4493 (N_4493,N_789,N_619);
nand U4494 (N_4494,N_429,N_1216);
and U4495 (N_4495,N_2125,N_404);
nand U4496 (N_4496,N_242,N_489);
nor U4497 (N_4497,N_1760,N_2282);
xor U4498 (N_4498,N_1356,N_1062);
xnor U4499 (N_4499,N_709,N_890);
xnor U4500 (N_4500,N_893,N_603);
and U4501 (N_4501,N_511,N_1898);
xor U4502 (N_4502,N_2140,N_1043);
or U4503 (N_4503,N_1901,N_1704);
or U4504 (N_4504,N_1812,N_188);
or U4505 (N_4505,N_864,N_1275);
and U4506 (N_4506,N_1159,N_1083);
xor U4507 (N_4507,N_2090,N_2222);
and U4508 (N_4508,N_2088,N_1466);
and U4509 (N_4509,N_926,N_1849);
nand U4510 (N_4510,N_1943,N_2057);
nand U4511 (N_4511,N_2384,N_392);
and U4512 (N_4512,N_1487,N_1266);
and U4513 (N_4513,N_2086,N_1062);
xor U4514 (N_4514,N_741,N_226);
and U4515 (N_4515,N_749,N_1466);
nor U4516 (N_4516,N_920,N_583);
nand U4517 (N_4517,N_412,N_1834);
or U4518 (N_4518,N_1784,N_1412);
nor U4519 (N_4519,N_1949,N_352);
nor U4520 (N_4520,N_1665,N_715);
xor U4521 (N_4521,N_2407,N_2443);
nand U4522 (N_4522,N_2095,N_620);
or U4523 (N_4523,N_2289,N_1450);
or U4524 (N_4524,N_791,N_1301);
xnor U4525 (N_4525,N_861,N_837);
nor U4526 (N_4526,N_2129,N_2254);
nand U4527 (N_4527,N_1151,N_2245);
nand U4528 (N_4528,N_69,N_786);
and U4529 (N_4529,N_249,N_266);
or U4530 (N_4530,N_1146,N_1281);
or U4531 (N_4531,N_774,N_1305);
and U4532 (N_4532,N_2343,N_51);
nand U4533 (N_4533,N_14,N_1824);
nand U4534 (N_4534,N_1687,N_1073);
and U4535 (N_4535,N_2099,N_1972);
or U4536 (N_4536,N_130,N_434);
nor U4537 (N_4537,N_1657,N_1968);
or U4538 (N_4538,N_1731,N_220);
and U4539 (N_4539,N_1373,N_601);
nand U4540 (N_4540,N_804,N_336);
or U4541 (N_4541,N_2133,N_1680);
or U4542 (N_4542,N_1396,N_853);
nor U4543 (N_4543,N_1510,N_1722);
xor U4544 (N_4544,N_1771,N_74);
xnor U4545 (N_4545,N_1566,N_322);
nand U4546 (N_4546,N_2138,N_2055);
nor U4547 (N_4547,N_577,N_1980);
nor U4548 (N_4548,N_1944,N_1937);
or U4549 (N_4549,N_2273,N_1756);
and U4550 (N_4550,N_1521,N_194);
and U4551 (N_4551,N_311,N_1465);
nor U4552 (N_4552,N_714,N_772);
or U4553 (N_4553,N_33,N_1397);
nor U4554 (N_4554,N_1809,N_1208);
nand U4555 (N_4555,N_614,N_78);
xor U4556 (N_4556,N_1734,N_880);
xor U4557 (N_4557,N_131,N_2223);
nand U4558 (N_4558,N_1090,N_533);
nor U4559 (N_4559,N_426,N_85);
xor U4560 (N_4560,N_2440,N_2257);
nand U4561 (N_4561,N_254,N_1399);
xor U4562 (N_4562,N_1667,N_2196);
xor U4563 (N_4563,N_667,N_846);
or U4564 (N_4564,N_1249,N_1063);
xor U4565 (N_4565,N_2450,N_1281);
and U4566 (N_4566,N_1409,N_1590);
and U4567 (N_4567,N_2387,N_88);
xor U4568 (N_4568,N_725,N_1644);
or U4569 (N_4569,N_1540,N_1370);
or U4570 (N_4570,N_803,N_2087);
xor U4571 (N_4571,N_1680,N_958);
or U4572 (N_4572,N_1378,N_1270);
and U4573 (N_4573,N_1156,N_504);
nor U4574 (N_4574,N_603,N_2408);
nor U4575 (N_4575,N_2441,N_1259);
nor U4576 (N_4576,N_493,N_578);
and U4577 (N_4577,N_896,N_1929);
nand U4578 (N_4578,N_1023,N_1077);
xor U4579 (N_4579,N_1299,N_197);
or U4580 (N_4580,N_2485,N_629);
xor U4581 (N_4581,N_750,N_1459);
and U4582 (N_4582,N_1740,N_592);
or U4583 (N_4583,N_2299,N_1345);
or U4584 (N_4584,N_2168,N_2397);
or U4585 (N_4585,N_356,N_2348);
and U4586 (N_4586,N_987,N_1539);
nand U4587 (N_4587,N_21,N_79);
and U4588 (N_4588,N_2004,N_1136);
and U4589 (N_4589,N_692,N_1638);
or U4590 (N_4590,N_1383,N_483);
or U4591 (N_4591,N_1479,N_1732);
nand U4592 (N_4592,N_1022,N_459);
or U4593 (N_4593,N_2055,N_2307);
nor U4594 (N_4594,N_958,N_650);
and U4595 (N_4595,N_1907,N_2115);
or U4596 (N_4596,N_1696,N_588);
and U4597 (N_4597,N_2102,N_880);
or U4598 (N_4598,N_2047,N_2338);
nand U4599 (N_4599,N_1833,N_775);
and U4600 (N_4600,N_1304,N_1899);
or U4601 (N_4601,N_152,N_891);
xor U4602 (N_4602,N_1612,N_2103);
or U4603 (N_4603,N_1353,N_2185);
and U4604 (N_4604,N_1771,N_2257);
or U4605 (N_4605,N_1015,N_2347);
and U4606 (N_4606,N_847,N_1511);
nand U4607 (N_4607,N_771,N_184);
nor U4608 (N_4608,N_1607,N_781);
nor U4609 (N_4609,N_821,N_1876);
nand U4610 (N_4610,N_1732,N_1094);
nand U4611 (N_4611,N_33,N_906);
nand U4612 (N_4612,N_1865,N_1984);
nor U4613 (N_4613,N_2134,N_892);
xor U4614 (N_4614,N_263,N_2345);
xnor U4615 (N_4615,N_2402,N_465);
and U4616 (N_4616,N_1076,N_2108);
and U4617 (N_4617,N_499,N_690);
xnor U4618 (N_4618,N_648,N_1775);
or U4619 (N_4619,N_2367,N_2473);
and U4620 (N_4620,N_120,N_2478);
and U4621 (N_4621,N_1387,N_76);
nand U4622 (N_4622,N_1609,N_2269);
xor U4623 (N_4623,N_2396,N_2197);
nor U4624 (N_4624,N_2273,N_1741);
nand U4625 (N_4625,N_1075,N_2256);
nand U4626 (N_4626,N_1837,N_1883);
nand U4627 (N_4627,N_230,N_799);
and U4628 (N_4628,N_2117,N_578);
nor U4629 (N_4629,N_272,N_458);
nand U4630 (N_4630,N_142,N_1038);
xor U4631 (N_4631,N_1971,N_574);
and U4632 (N_4632,N_2455,N_1246);
nor U4633 (N_4633,N_1422,N_2068);
or U4634 (N_4634,N_1036,N_102);
or U4635 (N_4635,N_1531,N_799);
nand U4636 (N_4636,N_525,N_1118);
or U4637 (N_4637,N_725,N_913);
or U4638 (N_4638,N_2139,N_2035);
xor U4639 (N_4639,N_680,N_563);
nor U4640 (N_4640,N_410,N_1906);
nor U4641 (N_4641,N_460,N_271);
and U4642 (N_4642,N_1896,N_254);
and U4643 (N_4643,N_1932,N_1428);
nand U4644 (N_4644,N_786,N_304);
xor U4645 (N_4645,N_2201,N_594);
xnor U4646 (N_4646,N_616,N_112);
xor U4647 (N_4647,N_502,N_570);
nand U4648 (N_4648,N_2400,N_780);
xnor U4649 (N_4649,N_1023,N_797);
nand U4650 (N_4650,N_923,N_1962);
nor U4651 (N_4651,N_1560,N_1233);
and U4652 (N_4652,N_751,N_2236);
nand U4653 (N_4653,N_1292,N_1072);
or U4654 (N_4654,N_848,N_880);
nand U4655 (N_4655,N_1208,N_1148);
or U4656 (N_4656,N_732,N_785);
or U4657 (N_4657,N_2226,N_425);
nand U4658 (N_4658,N_1393,N_1990);
nand U4659 (N_4659,N_1639,N_1766);
nor U4660 (N_4660,N_7,N_1264);
and U4661 (N_4661,N_429,N_689);
and U4662 (N_4662,N_1906,N_875);
xnor U4663 (N_4663,N_1627,N_2359);
and U4664 (N_4664,N_1391,N_153);
or U4665 (N_4665,N_483,N_1236);
or U4666 (N_4666,N_932,N_1765);
or U4667 (N_4667,N_1293,N_823);
nor U4668 (N_4668,N_604,N_2256);
nand U4669 (N_4669,N_807,N_2406);
or U4670 (N_4670,N_481,N_1767);
or U4671 (N_4671,N_1852,N_1301);
nor U4672 (N_4672,N_1921,N_1822);
and U4673 (N_4673,N_2259,N_593);
xnor U4674 (N_4674,N_1863,N_173);
or U4675 (N_4675,N_1218,N_2172);
and U4676 (N_4676,N_2439,N_919);
nor U4677 (N_4677,N_753,N_803);
nand U4678 (N_4678,N_2212,N_1398);
and U4679 (N_4679,N_2434,N_1747);
nand U4680 (N_4680,N_1869,N_1167);
and U4681 (N_4681,N_36,N_391);
nor U4682 (N_4682,N_46,N_1963);
xnor U4683 (N_4683,N_1478,N_49);
nor U4684 (N_4684,N_1537,N_1622);
xor U4685 (N_4685,N_1423,N_607);
xor U4686 (N_4686,N_1058,N_1174);
nand U4687 (N_4687,N_1563,N_730);
nand U4688 (N_4688,N_331,N_410);
nor U4689 (N_4689,N_1599,N_904);
and U4690 (N_4690,N_1693,N_598);
and U4691 (N_4691,N_349,N_1555);
xor U4692 (N_4692,N_163,N_1040);
or U4693 (N_4693,N_1243,N_2241);
and U4694 (N_4694,N_735,N_363);
nand U4695 (N_4695,N_2377,N_675);
nand U4696 (N_4696,N_586,N_103);
and U4697 (N_4697,N_2484,N_975);
and U4698 (N_4698,N_322,N_2169);
or U4699 (N_4699,N_1016,N_2040);
xnor U4700 (N_4700,N_298,N_1720);
nand U4701 (N_4701,N_2331,N_386);
nand U4702 (N_4702,N_492,N_423);
and U4703 (N_4703,N_296,N_2072);
xor U4704 (N_4704,N_1206,N_2069);
or U4705 (N_4705,N_671,N_473);
or U4706 (N_4706,N_506,N_36);
and U4707 (N_4707,N_21,N_2302);
xnor U4708 (N_4708,N_312,N_348);
nor U4709 (N_4709,N_66,N_1026);
nor U4710 (N_4710,N_965,N_127);
nor U4711 (N_4711,N_926,N_2350);
xnor U4712 (N_4712,N_412,N_1286);
nand U4713 (N_4713,N_583,N_640);
or U4714 (N_4714,N_378,N_293);
nor U4715 (N_4715,N_2213,N_484);
xnor U4716 (N_4716,N_105,N_690);
or U4717 (N_4717,N_77,N_2253);
or U4718 (N_4718,N_1456,N_1214);
or U4719 (N_4719,N_833,N_1472);
or U4720 (N_4720,N_704,N_2054);
nand U4721 (N_4721,N_1443,N_264);
and U4722 (N_4722,N_2030,N_457);
nand U4723 (N_4723,N_887,N_1669);
nand U4724 (N_4724,N_143,N_427);
nand U4725 (N_4725,N_1985,N_1847);
or U4726 (N_4726,N_1380,N_1796);
nand U4727 (N_4727,N_1392,N_349);
nor U4728 (N_4728,N_1745,N_195);
nand U4729 (N_4729,N_103,N_566);
or U4730 (N_4730,N_2100,N_2456);
nand U4731 (N_4731,N_1431,N_1560);
and U4732 (N_4732,N_1920,N_2045);
nand U4733 (N_4733,N_517,N_45);
nor U4734 (N_4734,N_226,N_2469);
xnor U4735 (N_4735,N_2171,N_858);
nor U4736 (N_4736,N_1785,N_2314);
nand U4737 (N_4737,N_2322,N_1842);
xor U4738 (N_4738,N_2212,N_671);
nand U4739 (N_4739,N_420,N_221);
xnor U4740 (N_4740,N_2133,N_339);
or U4741 (N_4741,N_2039,N_439);
and U4742 (N_4742,N_923,N_972);
or U4743 (N_4743,N_2435,N_1931);
and U4744 (N_4744,N_2233,N_2028);
or U4745 (N_4745,N_1656,N_1919);
xor U4746 (N_4746,N_139,N_2431);
and U4747 (N_4747,N_122,N_1687);
or U4748 (N_4748,N_2048,N_934);
or U4749 (N_4749,N_1417,N_2016);
and U4750 (N_4750,N_296,N_90);
nor U4751 (N_4751,N_645,N_2387);
xnor U4752 (N_4752,N_2421,N_698);
xnor U4753 (N_4753,N_1682,N_668);
xor U4754 (N_4754,N_1707,N_1202);
nand U4755 (N_4755,N_35,N_980);
or U4756 (N_4756,N_793,N_607);
xor U4757 (N_4757,N_2261,N_1003);
nor U4758 (N_4758,N_1927,N_962);
xor U4759 (N_4759,N_1298,N_1482);
nor U4760 (N_4760,N_2138,N_1855);
and U4761 (N_4761,N_1133,N_1764);
nor U4762 (N_4762,N_625,N_2384);
xor U4763 (N_4763,N_1870,N_1961);
nand U4764 (N_4764,N_364,N_1904);
or U4765 (N_4765,N_1259,N_1195);
nor U4766 (N_4766,N_1499,N_903);
nand U4767 (N_4767,N_1948,N_1969);
nor U4768 (N_4768,N_1147,N_678);
nand U4769 (N_4769,N_1584,N_168);
xor U4770 (N_4770,N_2374,N_593);
and U4771 (N_4771,N_2296,N_514);
nor U4772 (N_4772,N_2446,N_541);
xnor U4773 (N_4773,N_1844,N_1839);
and U4774 (N_4774,N_620,N_1029);
xnor U4775 (N_4775,N_1624,N_2328);
nand U4776 (N_4776,N_1101,N_538);
nand U4777 (N_4777,N_38,N_469);
or U4778 (N_4778,N_1379,N_199);
or U4779 (N_4779,N_1167,N_2005);
nor U4780 (N_4780,N_1628,N_1335);
nor U4781 (N_4781,N_1397,N_365);
or U4782 (N_4782,N_1308,N_1085);
and U4783 (N_4783,N_1586,N_1035);
and U4784 (N_4784,N_2145,N_318);
or U4785 (N_4785,N_426,N_520);
nor U4786 (N_4786,N_1995,N_56);
nor U4787 (N_4787,N_2291,N_1873);
nor U4788 (N_4788,N_1240,N_492);
xnor U4789 (N_4789,N_2400,N_130);
and U4790 (N_4790,N_778,N_2479);
and U4791 (N_4791,N_1424,N_1111);
and U4792 (N_4792,N_1333,N_1276);
nand U4793 (N_4793,N_322,N_1769);
xnor U4794 (N_4794,N_122,N_822);
nor U4795 (N_4795,N_2289,N_1579);
and U4796 (N_4796,N_495,N_364);
nand U4797 (N_4797,N_708,N_1461);
nand U4798 (N_4798,N_517,N_1342);
nor U4799 (N_4799,N_2276,N_2002);
xor U4800 (N_4800,N_452,N_2361);
and U4801 (N_4801,N_2173,N_1034);
nand U4802 (N_4802,N_1805,N_413);
xor U4803 (N_4803,N_2109,N_1349);
or U4804 (N_4804,N_1860,N_2450);
nand U4805 (N_4805,N_858,N_2360);
nand U4806 (N_4806,N_41,N_1113);
and U4807 (N_4807,N_447,N_2057);
or U4808 (N_4808,N_118,N_1778);
nand U4809 (N_4809,N_1883,N_1833);
or U4810 (N_4810,N_2398,N_469);
xnor U4811 (N_4811,N_111,N_1251);
or U4812 (N_4812,N_1788,N_1144);
and U4813 (N_4813,N_976,N_802);
or U4814 (N_4814,N_317,N_853);
and U4815 (N_4815,N_1579,N_440);
nand U4816 (N_4816,N_95,N_1551);
or U4817 (N_4817,N_439,N_1348);
nand U4818 (N_4818,N_863,N_2291);
and U4819 (N_4819,N_1150,N_868);
nor U4820 (N_4820,N_817,N_2375);
xor U4821 (N_4821,N_1505,N_661);
nand U4822 (N_4822,N_1291,N_2476);
and U4823 (N_4823,N_1483,N_120);
and U4824 (N_4824,N_1525,N_488);
nor U4825 (N_4825,N_719,N_318);
nor U4826 (N_4826,N_725,N_2003);
nand U4827 (N_4827,N_1035,N_404);
nand U4828 (N_4828,N_1949,N_2368);
or U4829 (N_4829,N_761,N_1599);
and U4830 (N_4830,N_489,N_828);
and U4831 (N_4831,N_1926,N_1202);
nand U4832 (N_4832,N_699,N_445);
nand U4833 (N_4833,N_955,N_1047);
or U4834 (N_4834,N_550,N_1690);
xor U4835 (N_4835,N_1333,N_2325);
or U4836 (N_4836,N_516,N_1881);
and U4837 (N_4837,N_80,N_2417);
or U4838 (N_4838,N_1701,N_505);
or U4839 (N_4839,N_602,N_1707);
nand U4840 (N_4840,N_1623,N_574);
and U4841 (N_4841,N_2017,N_2051);
nand U4842 (N_4842,N_2411,N_555);
or U4843 (N_4843,N_1943,N_1263);
or U4844 (N_4844,N_1997,N_1923);
nand U4845 (N_4845,N_1051,N_2104);
nor U4846 (N_4846,N_254,N_1964);
and U4847 (N_4847,N_420,N_817);
or U4848 (N_4848,N_2084,N_537);
nor U4849 (N_4849,N_1928,N_341);
nand U4850 (N_4850,N_1188,N_1967);
nor U4851 (N_4851,N_706,N_988);
and U4852 (N_4852,N_1295,N_10);
xnor U4853 (N_4853,N_682,N_1292);
or U4854 (N_4854,N_1064,N_1845);
nand U4855 (N_4855,N_1323,N_1195);
and U4856 (N_4856,N_1768,N_1331);
nand U4857 (N_4857,N_1455,N_779);
and U4858 (N_4858,N_2236,N_590);
and U4859 (N_4859,N_1652,N_855);
xor U4860 (N_4860,N_1772,N_70);
xnor U4861 (N_4861,N_504,N_1170);
nand U4862 (N_4862,N_2074,N_1975);
nand U4863 (N_4863,N_1640,N_698);
and U4864 (N_4864,N_1486,N_353);
and U4865 (N_4865,N_194,N_1885);
nand U4866 (N_4866,N_404,N_2098);
and U4867 (N_4867,N_1133,N_2217);
or U4868 (N_4868,N_2112,N_1202);
xor U4869 (N_4869,N_2048,N_289);
xnor U4870 (N_4870,N_606,N_320);
xor U4871 (N_4871,N_2196,N_901);
nor U4872 (N_4872,N_1981,N_669);
or U4873 (N_4873,N_1644,N_481);
or U4874 (N_4874,N_1777,N_751);
nand U4875 (N_4875,N_327,N_773);
and U4876 (N_4876,N_1931,N_9);
nor U4877 (N_4877,N_376,N_2208);
xor U4878 (N_4878,N_1931,N_169);
or U4879 (N_4879,N_1193,N_1470);
xnor U4880 (N_4880,N_2389,N_1050);
or U4881 (N_4881,N_700,N_1473);
or U4882 (N_4882,N_2032,N_900);
xor U4883 (N_4883,N_1713,N_983);
xnor U4884 (N_4884,N_2183,N_1737);
or U4885 (N_4885,N_1909,N_17);
and U4886 (N_4886,N_1938,N_1001);
or U4887 (N_4887,N_2077,N_1563);
or U4888 (N_4888,N_1855,N_322);
xor U4889 (N_4889,N_1577,N_1845);
and U4890 (N_4890,N_1489,N_1638);
nand U4891 (N_4891,N_257,N_174);
and U4892 (N_4892,N_1688,N_1493);
xnor U4893 (N_4893,N_370,N_74);
nand U4894 (N_4894,N_221,N_726);
nor U4895 (N_4895,N_2096,N_1011);
and U4896 (N_4896,N_2352,N_1397);
nand U4897 (N_4897,N_1003,N_1860);
nor U4898 (N_4898,N_1703,N_510);
or U4899 (N_4899,N_5,N_2428);
and U4900 (N_4900,N_2033,N_991);
nor U4901 (N_4901,N_1219,N_231);
nand U4902 (N_4902,N_109,N_777);
nand U4903 (N_4903,N_272,N_725);
xnor U4904 (N_4904,N_773,N_2164);
nor U4905 (N_4905,N_1494,N_1377);
xnor U4906 (N_4906,N_693,N_628);
or U4907 (N_4907,N_484,N_968);
nand U4908 (N_4908,N_293,N_1678);
nand U4909 (N_4909,N_2484,N_613);
and U4910 (N_4910,N_1862,N_1047);
and U4911 (N_4911,N_249,N_1912);
nor U4912 (N_4912,N_122,N_1317);
nor U4913 (N_4913,N_1024,N_1933);
nand U4914 (N_4914,N_1965,N_1031);
xnor U4915 (N_4915,N_545,N_691);
nand U4916 (N_4916,N_2482,N_21);
nor U4917 (N_4917,N_2069,N_1139);
nand U4918 (N_4918,N_415,N_626);
nor U4919 (N_4919,N_573,N_1131);
and U4920 (N_4920,N_1151,N_260);
nor U4921 (N_4921,N_1422,N_1317);
nor U4922 (N_4922,N_599,N_1862);
or U4923 (N_4923,N_1811,N_448);
and U4924 (N_4924,N_1737,N_729);
xnor U4925 (N_4925,N_1755,N_2235);
xor U4926 (N_4926,N_1387,N_249);
nor U4927 (N_4927,N_542,N_1483);
nand U4928 (N_4928,N_2476,N_1352);
or U4929 (N_4929,N_226,N_773);
and U4930 (N_4930,N_277,N_910);
nor U4931 (N_4931,N_395,N_2177);
or U4932 (N_4932,N_377,N_2349);
nor U4933 (N_4933,N_2152,N_484);
nor U4934 (N_4934,N_1071,N_2233);
nand U4935 (N_4935,N_290,N_2127);
nand U4936 (N_4936,N_98,N_57);
nor U4937 (N_4937,N_1300,N_434);
nand U4938 (N_4938,N_334,N_2422);
nor U4939 (N_4939,N_1033,N_986);
xnor U4940 (N_4940,N_173,N_1720);
nand U4941 (N_4941,N_593,N_1878);
or U4942 (N_4942,N_844,N_1669);
and U4943 (N_4943,N_1571,N_2427);
or U4944 (N_4944,N_1347,N_1501);
xnor U4945 (N_4945,N_1876,N_613);
or U4946 (N_4946,N_283,N_1657);
nor U4947 (N_4947,N_2034,N_1478);
and U4948 (N_4948,N_2378,N_2201);
nor U4949 (N_4949,N_243,N_1065);
nand U4950 (N_4950,N_1986,N_802);
nand U4951 (N_4951,N_1823,N_545);
nand U4952 (N_4952,N_1676,N_1727);
and U4953 (N_4953,N_434,N_976);
and U4954 (N_4954,N_1049,N_53);
nand U4955 (N_4955,N_920,N_1967);
or U4956 (N_4956,N_1097,N_892);
and U4957 (N_4957,N_1658,N_468);
or U4958 (N_4958,N_1326,N_2490);
nor U4959 (N_4959,N_1787,N_236);
nand U4960 (N_4960,N_500,N_1404);
and U4961 (N_4961,N_1557,N_1570);
nor U4962 (N_4962,N_2325,N_1204);
nor U4963 (N_4963,N_473,N_1786);
xor U4964 (N_4964,N_837,N_295);
xor U4965 (N_4965,N_367,N_1675);
nor U4966 (N_4966,N_2480,N_174);
nor U4967 (N_4967,N_694,N_1953);
nand U4968 (N_4968,N_1439,N_2199);
nand U4969 (N_4969,N_652,N_214);
xnor U4970 (N_4970,N_990,N_805);
nand U4971 (N_4971,N_750,N_2077);
nor U4972 (N_4972,N_1600,N_528);
and U4973 (N_4973,N_644,N_1741);
xnor U4974 (N_4974,N_792,N_1837);
nor U4975 (N_4975,N_1271,N_875);
nor U4976 (N_4976,N_1035,N_451);
nor U4977 (N_4977,N_1068,N_1195);
nor U4978 (N_4978,N_1360,N_510);
nand U4979 (N_4979,N_564,N_1731);
or U4980 (N_4980,N_95,N_1075);
xor U4981 (N_4981,N_207,N_1375);
xor U4982 (N_4982,N_212,N_1801);
or U4983 (N_4983,N_1517,N_344);
nand U4984 (N_4984,N_1802,N_1113);
xnor U4985 (N_4985,N_814,N_2054);
or U4986 (N_4986,N_1647,N_1708);
xor U4987 (N_4987,N_854,N_958);
nand U4988 (N_4988,N_1800,N_2100);
or U4989 (N_4989,N_2380,N_1764);
nor U4990 (N_4990,N_1024,N_137);
nor U4991 (N_4991,N_228,N_106);
and U4992 (N_4992,N_1985,N_1429);
nor U4993 (N_4993,N_867,N_1469);
and U4994 (N_4994,N_2412,N_148);
nand U4995 (N_4995,N_1067,N_1834);
and U4996 (N_4996,N_97,N_553);
and U4997 (N_4997,N_1239,N_1044);
nand U4998 (N_4998,N_1919,N_1782);
nand U4999 (N_4999,N_388,N_1371);
nand U5000 (N_5000,N_3810,N_4979);
nand U5001 (N_5001,N_3831,N_2677);
nand U5002 (N_5002,N_4025,N_3243);
xor U5003 (N_5003,N_4807,N_4969);
or U5004 (N_5004,N_4966,N_4331);
xnor U5005 (N_5005,N_2887,N_2557);
and U5006 (N_5006,N_3836,N_4198);
nand U5007 (N_5007,N_2848,N_3753);
nand U5008 (N_5008,N_3085,N_2732);
nand U5009 (N_5009,N_4061,N_2869);
xor U5010 (N_5010,N_2582,N_4813);
nor U5011 (N_5011,N_3435,N_3083);
nand U5012 (N_5012,N_4836,N_4497);
xor U5013 (N_5013,N_4475,N_3001);
xor U5014 (N_5014,N_4476,N_4839);
nor U5015 (N_5015,N_4482,N_3593);
nor U5016 (N_5016,N_3691,N_4354);
and U5017 (N_5017,N_2516,N_4717);
and U5018 (N_5018,N_2881,N_3550);
nand U5019 (N_5019,N_2715,N_4699);
and U5020 (N_5020,N_3141,N_4631);
and U5021 (N_5021,N_3358,N_3467);
and U5022 (N_5022,N_4693,N_3636);
and U5023 (N_5023,N_4275,N_2822);
xnor U5024 (N_5024,N_3166,N_4703);
nor U5025 (N_5025,N_2933,N_2700);
or U5026 (N_5026,N_3168,N_3882);
nor U5027 (N_5027,N_4056,N_4570);
xnor U5028 (N_5028,N_2517,N_4307);
and U5029 (N_5029,N_3616,N_3665);
nand U5030 (N_5030,N_3104,N_3486);
nor U5031 (N_5031,N_3761,N_2581);
and U5032 (N_5032,N_3638,N_3458);
and U5033 (N_5033,N_3605,N_2753);
or U5034 (N_5034,N_3056,N_4060);
or U5035 (N_5035,N_4862,N_3337);
nand U5036 (N_5036,N_2878,N_4353);
or U5037 (N_5037,N_4943,N_2917);
or U5038 (N_5038,N_2653,N_2718);
nand U5039 (N_5039,N_2756,N_3024);
nor U5040 (N_5040,N_4594,N_4081);
and U5041 (N_5041,N_2730,N_4287);
xor U5042 (N_5042,N_3362,N_4547);
xor U5043 (N_5043,N_3228,N_3971);
xor U5044 (N_5044,N_3142,N_3652);
and U5045 (N_5045,N_3967,N_3203);
nor U5046 (N_5046,N_4471,N_4278);
and U5047 (N_5047,N_4762,N_3409);
xor U5048 (N_5048,N_4940,N_2793);
nor U5049 (N_5049,N_3021,N_3192);
and U5050 (N_5050,N_4560,N_3277);
nand U5051 (N_5051,N_3783,N_2851);
nand U5052 (N_5052,N_2791,N_2725);
nor U5053 (N_5053,N_3892,N_4310);
nor U5054 (N_5054,N_3596,N_4024);
and U5055 (N_5055,N_2622,N_4067);
nand U5056 (N_5056,N_4069,N_4652);
xor U5057 (N_5057,N_4835,N_2987);
nor U5058 (N_5058,N_2561,N_4998);
nand U5059 (N_5059,N_4246,N_3426);
nand U5060 (N_5060,N_2646,N_3822);
nand U5061 (N_5061,N_4696,N_4820);
nor U5062 (N_5062,N_4956,N_2785);
or U5063 (N_5063,N_3842,N_2775);
and U5064 (N_5064,N_3431,N_4096);
or U5065 (N_5065,N_4898,N_4826);
and U5066 (N_5066,N_4445,N_3380);
xnor U5067 (N_5067,N_4095,N_3457);
or U5068 (N_5068,N_3630,N_4959);
and U5069 (N_5069,N_3093,N_4506);
nor U5070 (N_5070,N_3786,N_4416);
xor U5071 (N_5071,N_3960,N_3938);
nand U5072 (N_5072,N_4641,N_4350);
nand U5073 (N_5073,N_3549,N_3007);
xnor U5074 (N_5074,N_3449,N_3555);
and U5075 (N_5075,N_4563,N_4662);
and U5076 (N_5076,N_3463,N_3535);
nor U5077 (N_5077,N_4156,N_4248);
xor U5078 (N_5078,N_2918,N_3931);
nand U5079 (N_5079,N_3330,N_3412);
nand U5080 (N_5080,N_3137,N_3666);
or U5081 (N_5081,N_4910,N_2584);
nand U5082 (N_5082,N_3875,N_3559);
and U5083 (N_5083,N_4617,N_3706);
or U5084 (N_5084,N_4455,N_3461);
nand U5085 (N_5085,N_3052,N_3454);
xnor U5086 (N_5086,N_3191,N_3382);
or U5087 (N_5087,N_2518,N_4403);
nand U5088 (N_5088,N_3282,N_4197);
nor U5089 (N_5089,N_2911,N_3333);
or U5090 (N_5090,N_3547,N_4660);
or U5091 (N_5091,N_2832,N_4963);
or U5092 (N_5092,N_2662,N_2663);
xor U5093 (N_5093,N_4494,N_2945);
or U5094 (N_5094,N_4972,N_3769);
nand U5095 (N_5095,N_3235,N_3516);
nand U5096 (N_5096,N_4390,N_3470);
or U5097 (N_5097,N_4742,N_2652);
nor U5098 (N_5098,N_3254,N_4185);
and U5099 (N_5099,N_4167,N_4632);
nor U5100 (N_5100,N_2932,N_3447);
or U5101 (N_5101,N_4099,N_4834);
or U5102 (N_5102,N_4000,N_3906);
and U5103 (N_5103,N_4859,N_2991);
xor U5104 (N_5104,N_2706,N_4170);
nand U5105 (N_5105,N_3640,N_3830);
and U5106 (N_5106,N_2684,N_3301);
nor U5107 (N_5107,N_3058,N_2858);
nand U5108 (N_5108,N_3629,N_3552);
or U5109 (N_5109,N_4319,N_3494);
nor U5110 (N_5110,N_4753,N_2555);
and U5111 (N_5111,N_3854,N_4544);
nand U5112 (N_5112,N_4785,N_4819);
nand U5113 (N_5113,N_4871,N_4485);
xor U5114 (N_5114,N_4378,N_4181);
and U5115 (N_5115,N_4573,N_3386);
xnor U5116 (N_5116,N_4578,N_4131);
xnor U5117 (N_5117,N_3713,N_3539);
and U5118 (N_5118,N_3534,N_4811);
nand U5119 (N_5119,N_3818,N_4326);
nand U5120 (N_5120,N_4894,N_3963);
nor U5121 (N_5121,N_3866,N_2538);
nor U5122 (N_5122,N_2537,N_3434);
xor U5123 (N_5123,N_3112,N_4486);
or U5124 (N_5124,N_4759,N_4428);
nor U5125 (N_5125,N_4419,N_2890);
xor U5126 (N_5126,N_4335,N_4001);
or U5127 (N_5127,N_3576,N_4384);
or U5128 (N_5128,N_2977,N_3273);
and U5129 (N_5129,N_4603,N_2692);
and U5130 (N_5130,N_3639,N_4640);
nor U5131 (N_5131,N_4234,N_4997);
and U5132 (N_5132,N_2701,N_2962);
nand U5133 (N_5133,N_4680,N_3921);
nor U5134 (N_5134,N_4418,N_3482);
nand U5135 (N_5135,N_4540,N_2636);
xnor U5136 (N_5136,N_4609,N_2560);
and U5137 (N_5137,N_3767,N_3694);
nor U5138 (N_5138,N_3149,N_4723);
and U5139 (N_5139,N_4174,N_4017);
or U5140 (N_5140,N_4949,N_3765);
nand U5141 (N_5141,N_4417,N_4621);
xnor U5142 (N_5142,N_3130,N_4187);
xnor U5143 (N_5143,N_4232,N_4851);
nand U5144 (N_5144,N_4736,N_3060);
and U5145 (N_5145,N_4802,N_3451);
nor U5146 (N_5146,N_3909,N_4284);
nand U5147 (N_5147,N_3088,N_3441);
xor U5148 (N_5148,N_4464,N_3226);
and U5149 (N_5149,N_4944,N_3263);
nor U5150 (N_5150,N_3844,N_4683);
nand U5151 (N_5151,N_4149,N_4108);
and U5152 (N_5152,N_2596,N_3951);
nor U5153 (N_5153,N_2912,N_4302);
or U5154 (N_5154,N_4987,N_3527);
xnor U5155 (N_5155,N_2824,N_3568);
and U5156 (N_5156,N_4760,N_4144);
nor U5157 (N_5157,N_4143,N_2861);
or U5158 (N_5158,N_4827,N_4064);
nand U5159 (N_5159,N_2673,N_2626);
nand U5160 (N_5160,N_4038,N_2674);
nor U5161 (N_5161,N_4946,N_4450);
nand U5162 (N_5162,N_2639,N_4814);
and U5163 (N_5163,N_3813,N_3400);
or U5164 (N_5164,N_2751,N_2857);
and U5165 (N_5165,N_2812,N_4868);
xnor U5166 (N_5166,N_3657,N_4713);
or U5167 (N_5167,N_3891,N_2925);
or U5168 (N_5168,N_4176,N_3538);
and U5169 (N_5169,N_3712,N_4664);
or U5170 (N_5170,N_4155,N_3178);
xnor U5171 (N_5171,N_3816,N_4950);
xnor U5172 (N_5172,N_3331,N_3513);
or U5173 (N_5173,N_4113,N_3075);
nand U5174 (N_5174,N_3986,N_3393);
and U5175 (N_5175,N_2585,N_2610);
xor U5176 (N_5176,N_2600,N_3013);
or U5177 (N_5177,N_4220,N_4247);
and U5178 (N_5178,N_4294,N_4301);
xor U5179 (N_5179,N_3889,N_4519);
or U5180 (N_5180,N_4414,N_4424);
nand U5181 (N_5181,N_4899,N_2580);
xnor U5182 (N_5182,N_2532,N_4077);
nand U5183 (N_5183,N_3834,N_2839);
xnor U5184 (N_5184,N_3850,N_4228);
xnor U5185 (N_5185,N_4022,N_3586);
nor U5186 (N_5186,N_4120,N_4342);
xnor U5187 (N_5187,N_4180,N_2886);
or U5188 (N_5188,N_4537,N_4973);
and U5189 (N_5189,N_2528,N_4379);
nor U5190 (N_5190,N_3190,N_4088);
and U5191 (N_5191,N_3325,N_3182);
and U5192 (N_5192,N_4748,N_3053);
xnor U5193 (N_5193,N_4205,N_3741);
or U5194 (N_5194,N_2823,N_4195);
xor U5195 (N_5195,N_3624,N_4504);
and U5196 (N_5196,N_2989,N_3027);
nor U5197 (N_5197,N_4720,N_3840);
xnor U5198 (N_5198,N_4984,N_3020);
xor U5199 (N_5199,N_4731,N_4928);
and U5200 (N_5200,N_4566,N_3558);
nand U5201 (N_5201,N_3914,N_2844);
nand U5202 (N_5202,N_2860,N_3432);
nor U5203 (N_5203,N_3096,N_3643);
xnor U5204 (N_5204,N_4536,N_4732);
or U5205 (N_5205,N_4581,N_3403);
nand U5206 (N_5206,N_3355,N_3528);
and U5207 (N_5207,N_4217,N_2770);
and U5208 (N_5208,N_4021,N_4675);
and U5209 (N_5209,N_4382,N_3312);
xnor U5210 (N_5210,N_4087,N_2882);
nor U5211 (N_5211,N_3120,N_3949);
xnor U5212 (N_5212,N_3496,N_4325);
nand U5213 (N_5213,N_4716,N_3587);
xnor U5214 (N_5214,N_4211,N_4858);
nand U5215 (N_5215,N_4793,N_3530);
or U5216 (N_5216,N_4635,N_3995);
xnor U5217 (N_5217,N_3398,N_3578);
xor U5218 (N_5218,N_3029,N_4863);
and U5219 (N_5219,N_4479,N_3920);
xor U5220 (N_5220,N_3114,N_2536);
nor U5221 (N_5221,N_3123,N_3016);
xnor U5222 (N_5222,N_3611,N_3134);
nor U5223 (N_5223,N_3579,N_3208);
nor U5224 (N_5224,N_4459,N_3543);
xnor U5225 (N_5225,N_3401,N_4602);
and U5226 (N_5226,N_3430,N_3523);
and U5227 (N_5227,N_2985,N_2510);
nor U5228 (N_5228,N_4535,N_4468);
nand U5229 (N_5229,N_4656,N_4206);
xor U5230 (N_5230,N_3988,N_2849);
and U5231 (N_5231,N_3746,N_4221);
or U5232 (N_5232,N_2810,N_4242);
xnor U5233 (N_5233,N_3233,N_4089);
and U5234 (N_5234,N_4100,N_3040);
nand U5235 (N_5235,N_3385,N_3781);
nand U5236 (N_5236,N_3855,N_2603);
or U5237 (N_5237,N_3933,N_3899);
and U5238 (N_5238,N_4068,N_4867);
xor U5239 (N_5239,N_4639,N_4572);
xor U5240 (N_5240,N_3803,N_4323);
and U5241 (N_5241,N_3390,N_2968);
nand U5242 (N_5242,N_3151,N_3551);
xor U5243 (N_5243,N_4329,N_3727);
nor U5244 (N_5244,N_3147,N_3344);
and U5245 (N_5245,N_2734,N_4596);
nand U5246 (N_5246,N_4229,N_4383);
or U5247 (N_5247,N_2619,N_4129);
or U5248 (N_5248,N_4360,N_2893);
and U5249 (N_5249,N_3728,N_3491);
xor U5250 (N_5250,N_4746,N_3760);
nor U5251 (N_5251,N_3250,N_3747);
xnor U5252 (N_5252,N_3062,N_3105);
xor U5253 (N_5253,N_2675,N_3623);
and U5254 (N_5254,N_4942,N_3853);
xnor U5255 (N_5255,N_3846,N_4125);
and U5256 (N_5256,N_4882,N_4258);
nor U5257 (N_5257,N_3796,N_2661);
nor U5258 (N_5258,N_3809,N_2820);
nor U5259 (N_5259,N_2787,N_4999);
xor U5260 (N_5260,N_3485,N_4072);
nor U5261 (N_5261,N_3257,N_4209);
or U5262 (N_5262,N_4559,N_3992);
xnor U5263 (N_5263,N_4238,N_3363);
xnor U5264 (N_5264,N_4592,N_3987);
nor U5265 (N_5265,N_3455,N_4550);
nor U5266 (N_5266,N_3265,N_2884);
xor U5267 (N_5267,N_4279,N_4633);
or U5268 (N_5268,N_4150,N_4083);
or U5269 (N_5269,N_2888,N_2742);
nor U5270 (N_5270,N_4672,N_3678);
and U5271 (N_5271,N_3165,N_4488);
xnor U5272 (N_5272,N_2963,N_2697);
nor U5273 (N_5273,N_4786,N_4381);
xor U5274 (N_5274,N_2616,N_3492);
or U5275 (N_5275,N_3059,N_4066);
and U5276 (N_5276,N_4637,N_4577);
nand U5277 (N_5277,N_3839,N_4904);
or U5278 (N_5278,N_4292,N_3205);
or U5279 (N_5279,N_4140,N_2815);
or U5280 (N_5280,N_4196,N_2634);
or U5281 (N_5281,N_4816,N_3041);
nand U5282 (N_5282,N_3934,N_3940);
nor U5283 (N_5283,N_3019,N_2923);
xnor U5284 (N_5284,N_4044,N_4583);
xnor U5285 (N_5285,N_4362,N_4757);
or U5286 (N_5286,N_3782,N_3696);
or U5287 (N_5287,N_3102,N_3659);
and U5288 (N_5288,N_2608,N_3805);
nand U5289 (N_5289,N_4796,N_3708);
nor U5290 (N_5290,N_2960,N_4257);
or U5291 (N_5291,N_4576,N_3011);
nor U5292 (N_5292,N_4124,N_4626);
xnor U5293 (N_5293,N_4955,N_3873);
xnor U5294 (N_5294,N_3500,N_3111);
and U5295 (N_5295,N_2744,N_3721);
or U5296 (N_5296,N_3172,N_2948);
and U5297 (N_5297,N_2651,N_4800);
nand U5298 (N_5298,N_3081,N_2588);
nand U5299 (N_5299,N_4415,N_3258);
xor U5300 (N_5300,N_3739,N_4348);
xnor U5301 (N_5301,N_2831,N_2828);
and U5302 (N_5302,N_4924,N_3685);
and U5303 (N_5303,N_3662,N_3907);
nand U5304 (N_5304,N_4495,N_4437);
nand U5305 (N_5305,N_4616,N_2638);
nor U5306 (N_5306,N_3507,N_3961);
nand U5307 (N_5307,N_3904,N_3702);
nor U5308 (N_5308,N_3542,N_2698);
nor U5309 (N_5309,N_4297,N_3010);
or U5310 (N_5310,N_3724,N_4273);
and U5311 (N_5311,N_2975,N_3768);
and U5312 (N_5312,N_4651,N_2628);
nor U5313 (N_5313,N_2830,N_2906);
and U5314 (N_5314,N_4507,N_4063);
nor U5315 (N_5315,N_3043,N_3893);
nor U5316 (N_5316,N_3827,N_2723);
nand U5317 (N_5317,N_3188,N_4788);
or U5318 (N_5318,N_4630,N_4968);
nor U5319 (N_5319,N_4891,N_4778);
xor U5320 (N_5320,N_2821,N_3663);
nor U5321 (N_5321,N_4715,N_2826);
or U5322 (N_5322,N_4094,N_2834);
nand U5323 (N_5323,N_3022,N_4308);
nor U5324 (N_5324,N_4106,N_3865);
xnor U5325 (N_5325,N_3994,N_3080);
or U5326 (N_5326,N_2577,N_3135);
nor U5327 (N_5327,N_3119,N_3717);
nand U5328 (N_5328,N_3778,N_3249);
nand U5329 (N_5329,N_4905,N_4490);
nor U5330 (N_5330,N_3672,N_4521);
or U5331 (N_5331,N_2798,N_3144);
xor U5332 (N_5332,N_2609,N_3477);
or U5333 (N_5333,N_2615,N_3162);
xnor U5334 (N_5334,N_3614,N_3674);
and U5335 (N_5335,N_4877,N_3206);
and U5336 (N_5336,N_2789,N_2569);
or U5337 (N_5337,N_3991,N_4643);
xor U5338 (N_5338,N_3255,N_4971);
and U5339 (N_5339,N_4875,N_4389);
or U5340 (N_5340,N_2784,N_2944);
nand U5341 (N_5341,N_2618,N_4380);
xor U5342 (N_5342,N_4556,N_3957);
nand U5343 (N_5343,N_3063,N_4932);
nor U5344 (N_5344,N_4900,N_3481);
or U5345 (N_5345,N_4937,N_3014);
xnor U5346 (N_5346,N_3773,N_3997);
xor U5347 (N_5347,N_3795,N_3679);
nand U5348 (N_5348,N_4116,N_3095);
and U5349 (N_5349,N_3086,N_4613);
or U5350 (N_5350,N_3384,N_4747);
or U5351 (N_5351,N_3718,N_3342);
nor U5352 (N_5352,N_4227,N_4373);
nor U5353 (N_5353,N_3368,N_4841);
xnor U5354 (N_5354,N_2909,N_4030);
or U5355 (N_5355,N_3396,N_3688);
nor U5356 (N_5356,N_3026,N_4281);
and U5357 (N_5357,N_4398,N_2591);
nand U5358 (N_5358,N_2599,N_4545);
xnor U5359 (N_5359,N_4431,N_4579);
nand U5360 (N_5360,N_3510,N_4339);
or U5361 (N_5361,N_2875,N_3219);
or U5362 (N_5362,N_2867,N_2795);
xnor U5363 (N_5363,N_4792,N_4316);
nor U5364 (N_5364,N_4172,N_4915);
or U5365 (N_5365,N_4073,N_4138);
and U5366 (N_5366,N_2589,N_4502);
xor U5367 (N_5367,N_3881,N_2563);
nand U5368 (N_5368,N_4791,N_4847);
nor U5369 (N_5369,N_4309,N_2980);
and U5370 (N_5370,N_3811,N_4260);
or U5371 (N_5371,N_3560,N_3154);
or U5372 (N_5372,N_2666,N_2621);
and U5373 (N_5373,N_3048,N_3388);
nand U5374 (N_5374,N_2773,N_3962);
or U5375 (N_5375,N_3556,N_3828);
nand U5376 (N_5376,N_4085,N_3935);
or U5377 (N_5377,N_2930,N_4480);
and U5378 (N_5378,N_3240,N_2606);
or U5379 (N_5379,N_3750,N_3554);
nand U5380 (N_5380,N_3139,N_2656);
or U5381 (N_5381,N_4817,N_4013);
xnor U5382 (N_5382,N_3886,N_3730);
nor U5383 (N_5383,N_3705,N_3199);
and U5384 (N_5384,N_2546,N_2722);
or U5385 (N_5385,N_2919,N_3927);
and U5386 (N_5386,N_4520,N_3448);
xnor U5387 (N_5387,N_3184,N_3136);
or U5388 (N_5388,N_4527,N_2691);
nor U5389 (N_5389,N_4684,N_2951);
nand U5390 (N_5390,N_2748,N_4710);
and U5391 (N_5391,N_4688,N_4427);
nand U5392 (N_5392,N_2935,N_3101);
nor U5393 (N_5393,N_2984,N_2576);
nand U5394 (N_5394,N_3719,N_4148);
nand U5395 (N_5395,N_4860,N_4371);
and U5396 (N_5396,N_3793,N_2859);
nand U5397 (N_5397,N_2524,N_4745);
nand U5398 (N_5398,N_4023,N_4744);
and U5399 (N_5399,N_3817,N_3701);
xor U5400 (N_5400,N_2625,N_3784);
nand U5401 (N_5401,N_4532,N_2614);
nor U5402 (N_5402,N_2871,N_4884);
xnor U5403 (N_5403,N_3797,N_3890);
xor U5404 (N_5404,N_4727,N_3099);
nor U5405 (N_5405,N_3852,N_2708);
nand U5406 (N_5406,N_3641,N_4533);
nor U5407 (N_5407,N_2665,N_3653);
nand U5408 (N_5408,N_3771,N_3505);
xor U5409 (N_5409,N_3220,N_3469);
nand U5410 (N_5410,N_4250,N_4780);
or U5411 (N_5411,N_3518,N_2529);
nor U5412 (N_5412,N_3667,N_4794);
nor U5413 (N_5413,N_3731,N_4756);
xnor U5414 (N_5414,N_2946,N_3353);
or U5415 (N_5415,N_4305,N_4920);
and U5416 (N_5416,N_2549,N_2680);
nand U5417 (N_5417,N_4663,N_4674);
xnor U5418 (N_5418,N_4477,N_4879);
nand U5419 (N_5419,N_3474,N_2833);
nand U5420 (N_5420,N_4190,N_4991);
nand U5421 (N_5421,N_4874,N_2559);
or U5422 (N_5422,N_4948,N_2901);
xor U5423 (N_5423,N_3015,N_3117);
and U5424 (N_5424,N_3580,N_2696);
nand U5425 (N_5425,N_2737,N_2921);
nand U5426 (N_5426,N_4926,N_3187);
nor U5427 (N_5427,N_4127,N_4470);
nand U5428 (N_5428,N_2897,N_3131);
nand U5429 (N_5429,N_2883,N_3752);
xnor U5430 (N_5430,N_4412,N_3323);
nor U5431 (N_5431,N_3174,N_4356);
or U5432 (N_5432,N_4123,N_2741);
xor U5433 (N_5433,N_3375,N_3310);
nor U5434 (N_5434,N_3217,N_4327);
xor U5435 (N_5435,N_4865,N_3664);
or U5436 (N_5436,N_4912,N_4518);
and U5437 (N_5437,N_3573,N_4838);
nor U5438 (N_5438,N_4837,N_3153);
xnor U5439 (N_5439,N_2894,N_2876);
xor U5440 (N_5440,N_2633,N_2586);
xnor U5441 (N_5441,N_4829,N_3068);
or U5442 (N_5442,N_3395,N_2892);
xor U5443 (N_5443,N_3456,N_3429);
nand U5444 (N_5444,N_3391,N_4296);
and U5445 (N_5445,N_3300,N_3600);
and U5446 (N_5446,N_3862,N_4117);
or U5447 (N_5447,N_4918,N_3266);
xnor U5448 (N_5448,N_4509,N_3861);
nand U5449 (N_5449,N_3009,N_2966);
nor U5450 (N_5450,N_3780,N_4885);
or U5451 (N_5451,N_4618,N_4552);
or U5452 (N_5452,N_3480,N_3097);
nand U5453 (N_5453,N_4469,N_4266);
nor U5454 (N_5454,N_4806,N_3291);
xor U5455 (N_5455,N_3700,N_2659);
xor U5456 (N_5456,N_3416,N_2854);
xnor U5457 (N_5457,N_4958,N_4553);
or U5458 (N_5458,N_3606,N_2829);
and U5459 (N_5459,N_3309,N_4009);
nand U5460 (N_5460,N_4065,N_4401);
nand U5461 (N_5461,N_4989,N_3589);
xor U5462 (N_5462,N_2624,N_4890);
and U5463 (N_5463,N_3107,N_4110);
or U5464 (N_5464,N_3113,N_3436);
xor U5465 (N_5465,N_4259,N_3078);
nor U5466 (N_5466,N_4739,N_4330);
and U5467 (N_5467,N_2566,N_3847);
nor U5468 (N_5468,N_4845,N_4611);
nor U5469 (N_5469,N_2678,N_3180);
nand U5470 (N_5470,N_2551,N_4769);
nor U5471 (N_5471,N_4848,N_3159);
xnor U5472 (N_5472,N_4027,N_3379);
nor U5473 (N_5473,N_2969,N_3681);
xnor U5474 (N_5474,N_4893,N_3617);
or U5475 (N_5475,N_2686,N_4755);
and U5476 (N_5476,N_3037,N_4317);
or U5477 (N_5477,N_4191,N_3532);
or U5478 (N_5478,N_4036,N_3733);
or U5479 (N_5479,N_3374,N_3036);
nand U5480 (N_5480,N_2736,N_2738);
nand U5481 (N_5481,N_4134,N_4019);
and U5482 (N_5482,N_4584,N_3756);
nand U5483 (N_5483,N_4601,N_4654);
or U5484 (N_5484,N_4749,N_2643);
or U5485 (N_5485,N_3794,N_4233);
or U5486 (N_5486,N_2632,N_3253);
nand U5487 (N_5487,N_2740,N_2745);
nor U5488 (N_5488,N_3156,N_3256);
nor U5489 (N_5489,N_2762,N_3128);
nor U5490 (N_5490,N_2855,N_3157);
or U5491 (N_5491,N_3109,N_3517);
nand U5492 (N_5492,N_4164,N_3929);
nand U5493 (N_5493,N_3164,N_4016);
and U5494 (N_5494,N_4184,N_4192);
and U5495 (N_5495,N_2533,N_4557);
nand U5496 (N_5496,N_2952,N_3369);
xor U5497 (N_5497,N_4054,N_4719);
or U5498 (N_5498,N_3976,N_3592);
and U5499 (N_5499,N_4457,N_3615);
nand U5500 (N_5500,N_4312,N_4620);
xor U5501 (N_5501,N_4118,N_2801);
and U5502 (N_5502,N_4619,N_3295);
nand U5503 (N_5503,N_3069,N_3194);
or U5504 (N_5504,N_4567,N_4290);
and U5505 (N_5505,N_4853,N_2645);
nor U5506 (N_5506,N_3945,N_3487);
nand U5507 (N_5507,N_3757,N_2605);
and U5508 (N_5508,N_3418,N_4015);
nand U5509 (N_5509,N_4346,N_3092);
nor U5510 (N_5510,N_3497,N_2534);
and U5511 (N_5511,N_3654,N_3524);
and U5512 (N_5512,N_4681,N_4690);
xnor U5513 (N_5513,N_2814,N_2993);
nor U5514 (N_5514,N_4698,N_3346);
nor U5515 (N_5515,N_4650,N_2670);
nor U5516 (N_5516,N_3901,N_2950);
nor U5517 (N_5517,N_2955,N_4995);
or U5518 (N_5518,N_4236,N_4411);
and U5519 (N_5519,N_4409,N_4673);
nand U5520 (N_5520,N_4033,N_3584);
or U5521 (N_5521,N_4400,N_4208);
xor U5522 (N_5522,N_4996,N_3582);
xnor U5523 (N_5523,N_2712,N_4008);
or U5524 (N_5524,N_2852,N_4523);
nor U5525 (N_5525,N_4004,N_2819);
xor U5526 (N_5526,N_3227,N_4644);
nand U5527 (N_5527,N_2913,N_4886);
or U5528 (N_5528,N_3321,N_3898);
or U5529 (N_5529,N_3874,N_3407);
nor U5530 (N_5530,N_3484,N_4869);
or U5531 (N_5531,N_4162,N_4394);
and U5532 (N_5532,N_4665,N_3236);
nor U5533 (N_5533,N_4598,N_3627);
xnor U5534 (N_5534,N_3999,N_3671);
or U5535 (N_5535,N_3686,N_3122);
or U5536 (N_5536,N_3464,N_4318);
nand U5537 (N_5537,N_4677,N_3417);
nand U5538 (N_5538,N_4659,N_4333);
xor U5539 (N_5539,N_3952,N_4256);
nand U5540 (N_5540,N_3888,N_3821);
or U5541 (N_5541,N_3975,N_4372);
or U5542 (N_5542,N_4645,N_3758);
xnor U5543 (N_5543,N_3424,N_2922);
xnor U5544 (N_5544,N_4515,N_3919);
nor U5545 (N_5545,N_4976,N_4337);
and U5546 (N_5546,N_4965,N_3722);
nor U5547 (N_5547,N_3536,N_3361);
nand U5548 (N_5548,N_4655,N_4773);
or U5549 (N_5549,N_4104,N_3322);
and U5550 (N_5550,N_2799,N_2761);
xnor U5551 (N_5551,N_4005,N_2902);
nand U5552 (N_5552,N_2807,N_3110);
and U5553 (N_5553,N_3735,N_3108);
and U5554 (N_5554,N_3138,N_3711);
nand U5555 (N_5555,N_3443,N_3851);
nor U5556 (N_5556,N_4147,N_3977);
xor U5557 (N_5557,N_2936,N_2630);
nor U5558 (N_5558,N_4101,N_3057);
xor U5559 (N_5559,N_3471,N_3204);
nand U5560 (N_5560,N_2982,N_4889);
or U5561 (N_5561,N_3742,N_3425);
and U5562 (N_5562,N_2601,N_4831);
xnor U5563 (N_5563,N_3651,N_2514);
nor U5564 (N_5564,N_3476,N_4241);
nand U5565 (N_5565,N_4355,N_4718);
and U5566 (N_5566,N_4365,N_3089);
nand U5567 (N_5567,N_2726,N_3675);
or U5568 (N_5568,N_2777,N_3175);
xor U5569 (N_5569,N_2521,N_4797);
xnor U5570 (N_5570,N_4303,N_3006);
xor U5571 (N_5571,N_3948,N_2681);
and U5572 (N_5572,N_4990,N_4994);
nand U5573 (N_5573,N_3468,N_2842);
nor U5574 (N_5574,N_3790,N_3381);
and U5575 (N_5575,N_4421,N_4115);
and U5576 (N_5576,N_3612,N_4954);
nand U5577 (N_5577,N_2898,N_2573);
nor U5578 (N_5578,N_3302,N_4237);
nand U5579 (N_5579,N_3533,N_4695);
and U5580 (N_5580,N_4014,N_3317);
nor U5581 (N_5581,N_4048,N_3034);
and U5582 (N_5582,N_4870,N_4152);
xor U5583 (N_5583,N_4850,N_3947);
or U5584 (N_5584,N_3079,N_2664);
xnor U5585 (N_5585,N_4031,N_2598);
nor U5586 (N_5586,N_4391,N_4909);
xnor U5587 (N_5587,N_2927,N_4689);
nand U5588 (N_5588,N_2940,N_3293);
and U5589 (N_5589,N_4906,N_3376);
nand U5590 (N_5590,N_2978,N_4808);
nand U5591 (N_5591,N_4512,N_4255);
nor U5592 (N_5592,N_3460,N_3268);
nand U5593 (N_5593,N_4105,N_4440);
and U5594 (N_5594,N_4628,N_4453);
or U5595 (N_5595,N_4565,N_2719);
nor U5596 (N_5596,N_4590,N_3050);
or U5597 (N_5597,N_3347,N_2511);
nand U5598 (N_5598,N_2702,N_3699);
xnor U5599 (N_5599,N_3503,N_3423);
nand U5600 (N_5600,N_2905,N_3937);
nand U5601 (N_5601,N_3506,N_3121);
xor U5602 (N_5602,N_3224,N_3913);
or U5603 (N_5603,N_4002,N_2836);
and U5604 (N_5604,N_3276,N_4824);
nor U5605 (N_5605,N_3126,N_4981);
and U5606 (N_5606,N_4513,N_4474);
and U5607 (N_5607,N_4707,N_4936);
nor U5608 (N_5608,N_4114,N_3360);
and U5609 (N_5609,N_2850,N_3779);
nor U5610 (N_5610,N_3124,N_4055);
xor U5611 (N_5611,N_3304,N_3863);
xor U5612 (N_5612,N_2781,N_3242);
xnor U5613 (N_5613,N_2853,N_2938);
xor U5614 (N_5614,N_4254,N_2682);
xor U5615 (N_5615,N_4914,N_3002);
xnor U5616 (N_5616,N_2676,N_3032);
nand U5617 (N_5617,N_3303,N_4697);
and U5618 (N_5618,N_4210,N_3341);
nor U5619 (N_5619,N_4528,N_3896);
nand U5620 (N_5620,N_2800,N_2690);
nand U5621 (N_5621,N_2746,N_3023);
xnor U5622 (N_5622,N_3189,N_3176);
and U5623 (N_5623,N_4057,N_3008);
nor U5624 (N_5624,N_3098,N_2575);
nand U5625 (N_5625,N_2542,N_4447);
xnor U5626 (N_5626,N_4151,N_3859);
nand U5627 (N_5627,N_2788,N_4978);
nand U5628 (N_5628,N_2520,N_4933);
nand U5629 (N_5629,N_3285,N_3878);
or U5630 (N_5630,N_4574,N_3478);
and U5631 (N_5631,N_4084,N_3439);
or U5632 (N_5632,N_3815,N_3479);
nand U5633 (N_5633,N_2629,N_4102);
or U5634 (N_5634,N_2779,N_4974);
or U5635 (N_5635,N_2870,N_3966);
nand U5636 (N_5636,N_4046,N_2964);
or U5637 (N_5637,N_3290,N_3748);
or U5638 (N_5638,N_3213,N_3905);
nand U5639 (N_5639,N_3649,N_3613);
and U5640 (N_5640,N_2776,N_3049);
nand U5641 (N_5641,N_3444,N_4530);
nand U5642 (N_5642,N_4261,N_3197);
xnor U5643 (N_5643,N_2817,N_2749);
xor U5644 (N_5644,N_4472,N_4338);
nand U5645 (N_5645,N_3656,N_3956);
and U5646 (N_5646,N_2525,N_4153);
nand U5647 (N_5647,N_4171,N_4052);
nand U5648 (N_5648,N_4587,N_4525);
nor U5649 (N_5649,N_3405,N_4934);
nand U5650 (N_5650,N_3450,N_2843);
or U5651 (N_5651,N_4280,N_2772);
xnor U5652 (N_5652,N_3248,N_3218);
and U5653 (N_5653,N_4569,N_3996);
or U5654 (N_5654,N_4895,N_4435);
nand U5655 (N_5655,N_2556,N_4568);
nand U5656 (N_5656,N_3260,N_3209);
or U5657 (N_5657,N_3915,N_4709);
nand U5658 (N_5658,N_2545,N_3690);
nand U5659 (N_5659,N_4451,N_4923);
nor U5660 (N_5660,N_2729,N_4299);
or U5661 (N_5661,N_4803,N_4623);
or U5662 (N_5662,N_2595,N_3676);
nand U5663 (N_5663,N_3215,N_3682);
and U5664 (N_5664,N_3047,N_3259);
xnor U5665 (N_5665,N_2818,N_4582);
xnor U5666 (N_5666,N_3352,N_3744);
nand U5667 (N_5667,N_4789,N_2607);
and U5668 (N_5668,N_4142,N_2974);
xnor U5669 (N_5669,N_4441,N_4661);
or U5670 (N_5670,N_4770,N_4517);
nor U5671 (N_5671,N_3799,N_3601);
xor U5672 (N_5672,N_2825,N_3541);
or U5673 (N_5673,N_4952,N_4189);
or U5674 (N_5674,N_4341,N_4006);
nor U5675 (N_5675,N_3787,N_4622);
and U5676 (N_5676,N_4202,N_3709);
or U5677 (N_5677,N_2937,N_4591);
and U5678 (N_5678,N_2910,N_4289);
nand U5679 (N_5679,N_4436,N_3392);
and U5680 (N_5680,N_3211,N_4627);
nand U5681 (N_5681,N_4712,N_2868);
nor U5682 (N_5682,N_3521,N_3894);
and U5683 (N_5683,N_4636,N_3677);
and U5684 (N_5684,N_3658,N_2769);
or U5685 (N_5685,N_3288,N_2939);
nand U5686 (N_5686,N_4321,N_2505);
xnor U5687 (N_5687,N_2641,N_4043);
nand U5688 (N_5688,N_2597,N_3774);
or U5689 (N_5689,N_4489,N_4941);
xnor U5690 (N_5690,N_3504,N_2847);
and U5691 (N_5691,N_2637,N_4407);
or U5692 (N_5692,N_2866,N_3177);
nand U5693 (N_5693,N_4224,N_3459);
xor U5694 (N_5694,N_4496,N_4249);
xnor U5695 (N_5695,N_4666,N_3872);
and U5696 (N_5696,N_4975,N_3529);
nor U5697 (N_5697,N_2763,N_4078);
xnor U5698 (N_5698,N_3697,N_2757);
nand U5699 (N_5699,N_2928,N_3522);
and U5700 (N_5700,N_4200,N_4178);
nand U5701 (N_5701,N_2727,N_3626);
and U5702 (N_5702,N_2967,N_3824);
and U5703 (N_5703,N_4861,N_4678);
nor U5704 (N_5704,N_3628,N_3483);
nor U5705 (N_5705,N_4825,N_4215);
or U5706 (N_5706,N_4892,N_2703);
nor U5707 (N_5707,N_3725,N_3223);
and U5708 (N_5708,N_4163,N_4763);
nor U5709 (N_5709,N_3359,N_2895);
nor U5710 (N_5710,N_3028,N_4599);
and U5711 (N_5711,N_4432,N_3267);
xor U5712 (N_5712,N_3406,N_3350);
and U5713 (N_5713,N_4076,N_3158);
xor U5714 (N_5714,N_3094,N_2976);
xor U5715 (N_5715,N_3129,N_3585);
and U5716 (N_5716,N_4080,N_4776);
nor U5717 (N_5717,N_4774,N_3241);
nand U5718 (N_5718,N_2506,N_4487);
xor U5719 (N_5719,N_3619,N_2889);
and U5720 (N_5720,N_4951,N_4269);
nor U5721 (N_5721,N_2709,N_4529);
and U5722 (N_5722,N_3885,N_4543);
or U5723 (N_5723,N_3715,N_4691);
nand U5724 (N_5724,N_4810,N_4854);
nor U5725 (N_5725,N_4589,N_4324);
and U5726 (N_5726,N_4953,N_4268);
nor U5727 (N_5727,N_3823,N_3936);
xor U5728 (N_5728,N_3941,N_3160);
nand U5729 (N_5729,N_4881,N_4919);
or U5730 (N_5730,N_3005,N_2627);
xor U5731 (N_5731,N_4434,N_3819);
nand U5732 (N_5732,N_3087,N_3335);
and U5733 (N_5733,N_2669,N_2707);
nor U5734 (N_5734,N_3070,N_3514);
xor U5735 (N_5735,N_4728,N_2717);
nor U5736 (N_5736,N_4186,N_4604);
nand U5737 (N_5737,N_4272,N_4751);
nor U5738 (N_5738,N_3732,N_2885);
and U5739 (N_5739,N_4145,N_2640);
and U5740 (N_5740,N_2970,N_4558);
xor U5741 (N_5741,N_4705,N_3389);
xor U5742 (N_5742,N_4929,N_3595);
and U5743 (N_5743,N_2655,N_3442);
nand U5744 (N_5744,N_2949,N_3283);
or U5745 (N_5745,N_3917,N_4571);
xor U5746 (N_5746,N_3140,N_3314);
xor U5747 (N_5747,N_4107,N_3225);
nor U5748 (N_5748,N_4028,N_3729);
xor U5749 (N_5749,N_4740,N_4833);
and U5750 (N_5750,N_4286,N_4872);
nand U5751 (N_5751,N_3264,N_4642);
xor U5752 (N_5752,N_2837,N_2879);
and U5753 (N_5753,N_4916,N_2981);
and U5754 (N_5754,N_4037,N_3707);
xor U5755 (N_5755,N_2713,N_2594);
xnor U5756 (N_5756,N_3978,N_4597);
nor U5757 (N_5757,N_3912,N_4396);
nor U5758 (N_5758,N_4026,N_3884);
nand U5759 (N_5759,N_3411,N_3332);
nand U5760 (N_5760,N_2806,N_4798);
and U5761 (N_5761,N_2782,N_4805);
or U5762 (N_5762,N_3055,N_3804);
nor U5763 (N_5763,N_4694,N_4734);
nand U5764 (N_5764,N_3445,N_3438);
or U5765 (N_5765,N_3736,N_4729);
and U5766 (N_5766,N_3054,N_3902);
or U5767 (N_5767,N_3132,N_4423);
nand U5768 (N_5768,N_2531,N_4767);
xor U5769 (N_5769,N_3785,N_3631);
nor U5770 (N_5770,N_3887,N_3680);
xnor U5771 (N_5771,N_4032,N_3546);
xnor U5772 (N_5772,N_3324,N_3634);
nor U5773 (N_5773,N_3738,N_3196);
and U5774 (N_5774,N_3670,N_4313);
and U5775 (N_5775,N_4970,N_3645);
nand U5776 (N_5776,N_3367,N_2552);
nand U5777 (N_5777,N_4374,N_2931);
nor U5778 (N_5778,N_3848,N_4315);
nor U5779 (N_5779,N_3230,N_4347);
nand U5780 (N_5780,N_3798,N_3308);
nand U5781 (N_5781,N_2947,N_3714);
nand U5782 (N_5782,N_3849,N_2767);
or U5783 (N_5783,N_4930,N_3574);
and U5784 (N_5784,N_2693,N_4157);
xnor U5785 (N_5785,N_4982,N_3959);
and U5786 (N_5786,N_3012,N_3106);
and U5787 (N_5787,N_3826,N_2694);
nor U5788 (N_5788,N_4908,N_3064);
and U5789 (N_5789,N_3766,N_4961);
or U5790 (N_5790,N_3326,N_2695);
and U5791 (N_5791,N_4704,N_4967);
or U5792 (N_5792,N_3356,N_2720);
and U5793 (N_5793,N_2926,N_4377);
nor U5794 (N_5794,N_2813,N_3462);
xnor U5795 (N_5795,N_3646,N_4243);
nor U5796 (N_5796,N_4430,N_3939);
xnor U5797 (N_5797,N_3943,N_3755);
nand U5798 (N_5798,N_4300,N_2513);
nor U5799 (N_5799,N_2796,N_3954);
and U5800 (N_5800,N_3590,N_2808);
xnor U5801 (N_5801,N_3970,N_3599);
nand U5802 (N_5802,N_3833,N_3588);
nand U5803 (N_5803,N_4361,N_4925);
nor U5804 (N_5804,N_4843,N_2803);
nor U5805 (N_5805,N_4039,N_4173);
or U5806 (N_5806,N_3942,N_4752);
xnor U5807 (N_5807,N_3155,N_4600);
and U5808 (N_5808,N_4047,N_3270);
or U5809 (N_5809,N_3150,N_2735);
xor U5810 (N_5810,N_4011,N_4132);
or U5811 (N_5811,N_3399,N_3788);
and U5812 (N_5812,N_4711,N_2685);
or U5813 (N_5813,N_3704,N_3625);
and U5814 (N_5814,N_3868,N_3775);
nor U5815 (N_5815,N_4059,N_4448);
and U5816 (N_5816,N_3229,N_2809);
xor U5817 (N_5817,N_3378,N_4334);
xnor U5818 (N_5818,N_2530,N_3982);
and U5819 (N_5819,N_3565,N_3419);
or U5820 (N_5820,N_2986,N_4075);
nor U5821 (N_5821,N_3922,N_3620);
and U5822 (N_5822,N_4282,N_3046);
and U5823 (N_5823,N_2509,N_3608);
or U5824 (N_5824,N_3493,N_3591);
and U5825 (N_5825,N_3319,N_3918);
or U5826 (N_5826,N_4179,N_2631);
and U5827 (N_5827,N_3740,N_2650);
nand U5828 (N_5828,N_2574,N_3090);
and U5829 (N_5829,N_4399,N_2804);
nor U5830 (N_5830,N_2846,N_3415);
xnor U5831 (N_5831,N_4158,N_3537);
xor U5832 (N_5832,N_3743,N_3557);
nand U5833 (N_5833,N_4126,N_2774);
or U5834 (N_5834,N_3067,N_4830);
nand U5835 (N_5835,N_4082,N_3508);
and U5836 (N_5836,N_3373,N_3287);
nor U5837 (N_5837,N_4768,N_3495);
or U5838 (N_5838,N_4779,N_4702);
nor U5839 (N_5839,N_3869,N_4074);
nand U5840 (N_5840,N_2983,N_4093);
xnor U5841 (N_5841,N_4931,N_3575);
nand U5842 (N_5842,N_4491,N_4071);
nor U5843 (N_5843,N_4866,N_3511);
xnor U5844 (N_5844,N_3038,N_3812);
and U5845 (N_5845,N_2994,N_4306);
and U5846 (N_5846,N_3051,N_4692);
or U5847 (N_5847,N_2896,N_2766);
xnor U5848 (N_5848,N_3562,N_4203);
nand U5849 (N_5849,N_2864,N_2500);
and U5850 (N_5850,N_3076,N_4050);
and U5851 (N_5851,N_4864,N_3669);
nor U5852 (N_5852,N_4079,N_2965);
nand U5853 (N_5853,N_4492,N_3895);
and U5854 (N_5854,N_2759,N_4304);
xor U5855 (N_5855,N_3789,N_3509);
xnor U5856 (N_5856,N_3408,N_4135);
and U5857 (N_5857,N_3983,N_3465);
and U5858 (N_5858,N_2667,N_4385);
or U5859 (N_5859,N_2523,N_4741);
nand U5860 (N_5860,N_3602,N_3271);
nor U5861 (N_5861,N_3103,N_4730);
or U5862 (N_5862,N_2764,N_4765);
xnor U5863 (N_5863,N_4947,N_3566);
xor U5864 (N_5864,N_3955,N_3163);
xnor U5865 (N_5865,N_3564,N_4873);
and U5866 (N_5866,N_3762,N_4795);
nand U5867 (N_5867,N_3179,N_3035);
nand U5868 (N_5868,N_2721,N_3598);
nand U5869 (N_5869,N_4370,N_4562);
or U5870 (N_5870,N_3660,N_3161);
nor U5871 (N_5871,N_3985,N_3452);
nor U5872 (N_5872,N_3900,N_4460);
and U5873 (N_5873,N_4701,N_3025);
and U5874 (N_5874,N_4510,N_3239);
nor U5875 (N_5875,N_3622,N_3252);
nor U5876 (N_5876,N_2862,N_2512);
and U5877 (N_5877,N_4413,N_4034);
or U5878 (N_5878,N_3974,N_2593);
nand U5879 (N_5879,N_3148,N_3519);
and U5880 (N_5880,N_4183,N_4443);
and U5881 (N_5881,N_3498,N_3512);
xor U5882 (N_5882,N_4393,N_4531);
nor U5883 (N_5883,N_2841,N_3000);
and U5884 (N_5884,N_4405,N_3232);
nor U5885 (N_5885,N_4498,N_2877);
and U5886 (N_5886,N_3198,N_4288);
nand U5887 (N_5887,N_3349,N_2644);
and U5888 (N_5888,N_4700,N_3860);
or U5889 (N_5889,N_3916,N_3170);
xnor U5890 (N_5890,N_3410,N_3501);
nand U5891 (N_5891,N_4340,N_3281);
nor U5892 (N_5892,N_4901,N_4575);
and U5893 (N_5893,N_3490,N_4465);
or U5894 (N_5894,N_4667,N_3820);
and U5895 (N_5895,N_4388,N_3597);
nand U5896 (N_5896,N_3200,N_3567);
and U5897 (N_5897,N_3515,N_4625);
nor U5898 (N_5898,N_3647,N_4896);
or U5899 (N_5899,N_4986,N_4722);
and U5900 (N_5900,N_2654,N_4624);
and U5901 (N_5901,N_3387,N_2920);
nor U5902 (N_5902,N_3127,N_4426);
and U5903 (N_5903,N_2613,N_4526);
xnor U5904 (N_5904,N_2671,N_2535);
xor U5905 (N_5905,N_4669,N_2567);
nand U5906 (N_5906,N_4721,N_3306);
xor U5907 (N_5907,N_2527,N_3207);
and U5908 (N_5908,N_3698,N_4336);
and U5909 (N_5909,N_2579,N_3313);
nand U5910 (N_5910,N_4214,N_4781);
or U5911 (N_5911,N_3169,N_4349);
nor U5912 (N_5912,N_2750,N_3637);
or U5913 (N_5913,N_4483,N_3973);
nor U5914 (N_5914,N_2731,N_4070);
nand U5915 (N_5915,N_2973,N_4086);
or U5916 (N_5916,N_4514,N_2522);
or U5917 (N_5917,N_2908,N_3298);
and U5918 (N_5918,N_3668,N_3299);
or U5919 (N_5919,N_3100,N_2572);
and U5920 (N_5920,N_4395,N_2953);
or U5921 (N_5921,N_3466,N_3222);
and U5922 (N_5922,N_3751,N_2797);
nor U5923 (N_5923,N_2562,N_4392);
xor U5924 (N_5924,N_3320,N_3609);
nor U5925 (N_5925,N_2647,N_3338);
or U5926 (N_5926,N_3993,N_3212);
and U5927 (N_5927,N_2783,N_4442);
nand U5928 (N_5928,N_3689,N_3737);
xor U5929 (N_5929,N_4939,N_3329);
and U5930 (N_5930,N_4685,N_4818);
nor U5931 (N_5931,N_4375,N_2526);
nor U5932 (N_5932,N_2956,N_4109);
xnor U5933 (N_5933,N_4408,N_3570);
and U5934 (N_5934,N_3540,N_3234);
nand U5935 (N_5935,N_4463,N_2942);
and U5936 (N_5936,N_3437,N_4444);
xor U5937 (N_5937,N_4352,N_3923);
xor U5938 (N_5938,N_3402,N_3475);
and U5939 (N_5939,N_2957,N_4649);
nor U5940 (N_5940,N_4883,N_3801);
nor U5941 (N_5941,N_2780,N_3371);
or U5942 (N_5942,N_4429,N_4449);
nand U5943 (N_5943,N_4277,N_4985);
nor U5944 (N_5944,N_3604,N_3932);
nand U5945 (N_5945,N_3274,N_3814);
and U5946 (N_5946,N_3577,N_4917);
nand U5947 (N_5947,N_2865,N_4128);
nor U5948 (N_5948,N_4511,N_4962);
and U5949 (N_5949,N_3296,N_3764);
xnor U5950 (N_5950,N_4458,N_4772);
xnor U5951 (N_5951,N_3262,N_3366);
and U5952 (N_5952,N_3428,N_4516);
xnor U5953 (N_5953,N_3339,N_4840);
nor U5954 (N_5954,N_4832,N_4588);
and U5955 (N_5955,N_4686,N_4274);
nor U5956 (N_5956,N_3334,N_4397);
xnor U5957 (N_5957,N_4657,N_3928);
nor U5958 (N_5958,N_3871,N_3980);
nand U5959 (N_5959,N_2683,N_4119);
nand U5960 (N_5960,N_3754,N_3173);
and U5961 (N_5961,N_2874,N_4585);
or U5962 (N_5962,N_2873,N_4549);
xor U5963 (N_5963,N_3286,N_2548);
nand U5964 (N_5964,N_2604,N_3650);
nand U5965 (N_5965,N_3989,N_4708);
nand U5966 (N_5966,N_3867,N_3427);
nor U5967 (N_5967,N_3116,N_4098);
and U5968 (N_5968,N_4446,N_3214);
xnor U5969 (N_5969,N_2838,N_4606);
xor U5970 (N_5970,N_3687,N_3311);
nand U5971 (N_5971,N_4771,N_4366);
nor U5972 (N_5972,N_2743,N_4225);
nor U5973 (N_5973,N_4823,N_4314);
nand U5974 (N_5974,N_2635,N_3003);
or U5975 (N_5975,N_2711,N_3018);
nor U5976 (N_5976,N_3316,N_2689);
and U5977 (N_5977,N_3433,N_4505);
nand U5978 (N_5978,N_4668,N_3031);
and U5979 (N_5979,N_3171,N_4035);
nor U5980 (N_5980,N_4546,N_4658);
xnor U5981 (N_5981,N_2515,N_3440);
and U5982 (N_5982,N_3044,N_2688);
and U5983 (N_5983,N_3348,N_4878);
and U5984 (N_5984,N_3231,N_3684);
or U5985 (N_5985,N_4983,N_3548);
xor U5986 (N_5986,N_2672,N_3969);
nand U5987 (N_5987,N_4849,N_2805);
xor U5988 (N_5988,N_3186,N_4593);
and U5989 (N_5989,N_4239,N_3525);
nor U5990 (N_5990,N_4103,N_3526);
or U5991 (N_5991,N_2996,N_3261);
xnor U5992 (N_5992,N_4357,N_4524);
or U5993 (N_5993,N_4204,N_4647);
nor U5994 (N_5994,N_4844,N_3883);
xor U5995 (N_5995,N_2845,N_4508);
xnor U5996 (N_5996,N_2997,N_4363);
or U5997 (N_5997,N_4235,N_4466);
or U5998 (N_5998,N_2508,N_4218);
and U5999 (N_5999,N_3473,N_4332);
nor U6000 (N_6000,N_3284,N_4012);
xor U6001 (N_6001,N_3297,N_2739);
and U6002 (N_6002,N_3792,N_3964);
nand U6003 (N_6003,N_3777,N_4605);
xor U6004 (N_6004,N_4737,N_3074);
nand U6005 (N_6005,N_3910,N_4422);
or U6006 (N_6006,N_4761,N_4777);
nor U6007 (N_6007,N_3563,N_3772);
and U6008 (N_6008,N_3569,N_2943);
nor U6009 (N_6009,N_3143,N_3802);
or U6010 (N_6010,N_4168,N_4262);
nand U6011 (N_6011,N_4481,N_2929);
and U6012 (N_6012,N_2587,N_3825);
or U6013 (N_6013,N_3251,N_3835);
nor U6014 (N_6014,N_4907,N_4298);
and U6015 (N_6015,N_4358,N_4534);
or U6016 (N_6016,N_4935,N_2880);
or U6017 (N_6017,N_4433,N_4058);
or U6018 (N_6018,N_4738,N_3897);
nand U6019 (N_6019,N_4240,N_4045);
xnor U6020 (N_6020,N_3354,N_3413);
nand U6021 (N_6021,N_3520,N_4783);
xnor U6022 (N_6022,N_3201,N_4452);
nor U6023 (N_6023,N_3953,N_3181);
nand U6024 (N_6024,N_2915,N_2728);
xor U6025 (N_6025,N_4580,N_2540);
nor U6026 (N_6026,N_4226,N_3857);
nor U6027 (N_6027,N_3336,N_3603);
or U6028 (N_6028,N_3195,N_3091);
nor U6029 (N_6029,N_3618,N_4406);
and U6030 (N_6030,N_4213,N_3327);
xnor U6031 (N_6031,N_3998,N_3305);
and U6032 (N_6032,N_2752,N_3193);
xnor U6033 (N_6033,N_2771,N_3377);
and U6034 (N_6034,N_2995,N_3221);
or U6035 (N_6035,N_3238,N_4706);
and U6036 (N_6036,N_4439,N_3318);
nor U6037 (N_6037,N_2768,N_3042);
xnor U6038 (N_6038,N_2502,N_3502);
and U6039 (N_6039,N_2705,N_3745);
or U6040 (N_6040,N_4960,N_3280);
or U6041 (N_6041,N_3066,N_2754);
nor U6042 (N_6042,N_3061,N_3880);
and U6043 (N_6043,N_2827,N_3545);
nand U6044 (N_6044,N_4244,N_3693);
xor U6045 (N_6045,N_3245,N_4880);
or U6046 (N_6046,N_2916,N_2899);
nor U6047 (N_6047,N_3633,N_4161);
nand U6048 (N_6048,N_4499,N_4897);
nand U6049 (N_6049,N_4041,N_4367);
and U6050 (N_6050,N_3958,N_4784);
or U6051 (N_6051,N_4344,N_3404);
or U6052 (N_6052,N_4799,N_4276);
or U6053 (N_6053,N_3829,N_4283);
nand U6054 (N_6054,N_4219,N_3944);
nand U6055 (N_6055,N_4608,N_3837);
xor U6056 (N_6056,N_3125,N_4137);
nor U6057 (N_6057,N_2704,N_3370);
or U6058 (N_6058,N_4522,N_4787);
nand U6059 (N_6059,N_4473,N_3118);
and U6060 (N_6060,N_4188,N_3365);
or U6061 (N_6061,N_2924,N_4438);
nor U6062 (N_6062,N_4676,N_2872);
and U6063 (N_6063,N_4493,N_3673);
xor U6064 (N_6064,N_4501,N_4993);
xor U6065 (N_6065,N_3908,N_3272);
or U6066 (N_6066,N_3571,N_4222);
nor U6067 (N_6067,N_4539,N_2990);
nor U6068 (N_6068,N_3642,N_3357);
and U6069 (N_6069,N_4790,N_2519);
nor U6070 (N_6070,N_4852,N_3661);
and U6071 (N_6071,N_4538,N_3082);
or U6072 (N_6072,N_4913,N_4542);
xnor U6073 (N_6073,N_3216,N_4311);
or U6074 (N_6074,N_4177,N_4467);
and U6075 (N_6075,N_3372,N_4121);
xor U6076 (N_6076,N_3621,N_4040);
or U6077 (N_6077,N_3343,N_3692);
nand U6078 (N_6078,N_2570,N_4136);
xnor U6079 (N_6079,N_4945,N_3870);
nor U6080 (N_6080,N_3644,N_3553);
nor U6081 (N_6081,N_3152,N_4345);
and U6082 (N_6082,N_4212,N_3030);
xor U6083 (N_6083,N_3446,N_4018);
xnor U6084 (N_6084,N_4615,N_3420);
xor U6085 (N_6085,N_4634,N_2934);
nor U6086 (N_6086,N_4402,N_3328);
nand U6087 (N_6087,N_4648,N_4735);
or U6088 (N_6088,N_2903,N_4750);
and U6089 (N_6089,N_4146,N_4160);
or U6090 (N_6090,N_3632,N_2794);
nand U6091 (N_6091,N_3364,N_4815);
xor U6092 (N_6092,N_3581,N_4293);
and U6093 (N_6093,N_2554,N_4724);
nand U6094 (N_6094,N_3084,N_2623);
or U6095 (N_6095,N_4638,N_2558);
and U6096 (N_6096,N_4166,N_3307);
and U6097 (N_6097,N_2816,N_2611);
nand U6098 (N_6098,N_4051,N_3397);
nand U6099 (N_6099,N_4270,N_3864);
and U6100 (N_6100,N_3572,N_3315);
nand U6101 (N_6101,N_4733,N_2565);
nand U6102 (N_6102,N_2998,N_4291);
xor U6103 (N_6103,N_4462,N_2792);
nor U6104 (N_6104,N_4193,N_4484);
nand U6105 (N_6105,N_3499,N_3903);
xor U6106 (N_6106,N_2972,N_2811);
nor U6107 (N_6107,N_4285,N_4725);
and U6108 (N_6108,N_4130,N_3635);
nor U6109 (N_6109,N_2988,N_4822);
and U6110 (N_6110,N_4503,N_4614);
xnor U6111 (N_6111,N_4376,N_3710);
nor U6112 (N_6112,N_4387,N_2602);
nand U6113 (N_6113,N_2592,N_4320);
and U6114 (N_6114,N_2961,N_2724);
nor U6115 (N_6115,N_3017,N_3791);
nand U6116 (N_6116,N_3806,N_3726);
nor U6117 (N_6117,N_4454,N_2658);
xnor U6118 (N_6118,N_3594,N_4245);
or U6119 (N_6119,N_4343,N_3723);
xnor U6120 (N_6120,N_4159,N_4368);
xnor U6121 (N_6121,N_4754,N_3292);
nand U6122 (N_6122,N_2550,N_2891);
and U6123 (N_6123,N_4564,N_4223);
and U6124 (N_6124,N_2765,N_4782);
nand U6125 (N_6125,N_3289,N_3695);
and U6126 (N_6126,N_3246,N_4165);
nor U6127 (N_6127,N_3965,N_3683);
or U6128 (N_6128,N_3489,N_4964);
or U6129 (N_6129,N_2620,N_2590);
nor U6130 (N_6130,N_4322,N_3269);
xnor U6131 (N_6131,N_4062,N_2747);
xor U6132 (N_6132,N_4876,N_3039);
and U6133 (N_6133,N_4231,N_3984);
nand U6134 (N_6134,N_3946,N_4679);
nand U6135 (N_6135,N_2840,N_4646);
and U6136 (N_6136,N_4992,N_2979);
and U6137 (N_6137,N_3610,N_4812);
nand U6138 (N_6138,N_4364,N_4175);
xnor U6139 (N_6139,N_2660,N_3703);
and U6140 (N_6140,N_3279,N_3926);
xor U6141 (N_6141,N_4500,N_2583);
nor U6142 (N_6142,N_4263,N_4856);
nor U6143 (N_6143,N_4049,N_2571);
or U6144 (N_6144,N_4169,N_4980);
and U6145 (N_6145,N_3071,N_2941);
or U6146 (N_6146,N_3544,N_4828);
and U6147 (N_6147,N_3843,N_2786);
xnor U6148 (N_6148,N_4855,N_4133);
or U6149 (N_6149,N_3278,N_2760);
and U6150 (N_6150,N_2612,N_3950);
nor U6151 (N_6151,N_2863,N_4478);
nor U6152 (N_6152,N_4194,N_4957);
nand U6153 (N_6153,N_4612,N_2790);
nand U6154 (N_6154,N_4555,N_4141);
nand U6155 (N_6155,N_3979,N_4764);
xnor U6156 (N_6156,N_3734,N_4671);
nand U6157 (N_6157,N_4207,N_2657);
nor U6158 (N_6158,N_4267,N_4554);
and U6159 (N_6159,N_3237,N_4010);
or U6160 (N_6160,N_4386,N_4097);
nand U6161 (N_6161,N_3531,N_4846);
and U6162 (N_6162,N_3763,N_2568);
and U6163 (N_6163,N_4053,N_3838);
or U6164 (N_6164,N_2959,N_3421);
or U6165 (N_6165,N_3807,N_3472);
nand U6166 (N_6166,N_4216,N_2544);
or U6167 (N_6167,N_4887,N_2668);
xnor U6168 (N_6168,N_4911,N_2642);
and U6169 (N_6169,N_4295,N_4682);
or U6170 (N_6170,N_4842,N_4977);
xnor U6171 (N_6171,N_2733,N_4687);
or U6172 (N_6172,N_2835,N_3202);
nor U6173 (N_6173,N_3607,N_4586);
nand U6174 (N_6174,N_4351,N_4020);
or U6175 (N_6175,N_4090,N_3879);
nand U6176 (N_6176,N_4541,N_4548);
xor U6177 (N_6177,N_2649,N_2999);
nor U6178 (N_6178,N_3972,N_4801);
xnor U6179 (N_6179,N_3749,N_3183);
nand U6180 (N_6180,N_3776,N_4369);
nand U6181 (N_6181,N_2539,N_4007);
xnor U6182 (N_6182,N_2617,N_4922);
or U6183 (N_6183,N_2687,N_2755);
and U6184 (N_6184,N_2564,N_4265);
or U6185 (N_6185,N_3422,N_2758);
nor U6186 (N_6186,N_3340,N_2958);
and U6187 (N_6187,N_3925,N_4903);
and U6188 (N_6188,N_4595,N_3648);
nand U6189 (N_6189,N_4610,N_3167);
or U6190 (N_6190,N_3808,N_4888);
or U6191 (N_6191,N_4252,N_2541);
nand U6192 (N_6192,N_3294,N_4264);
or U6193 (N_6193,N_4139,N_3924);
and U6194 (N_6194,N_3145,N_4726);
nand U6195 (N_6195,N_3990,N_3210);
nor U6196 (N_6196,N_2802,N_4456);
or U6197 (N_6197,N_4230,N_3394);
and U6198 (N_6198,N_4607,N_3453);
nor U6199 (N_6199,N_3911,N_2778);
or U6200 (N_6200,N_3383,N_4271);
nand U6201 (N_6201,N_4199,N_4988);
or U6202 (N_6202,N_2856,N_2501);
nand U6203 (N_6203,N_2578,N_3561);
and U6204 (N_6204,N_4092,N_3414);
and U6205 (N_6205,N_3876,N_2543);
xnor U6206 (N_6206,N_3275,N_4743);
nor U6207 (N_6207,N_2503,N_3004);
and U6208 (N_6208,N_4804,N_3832);
nand U6209 (N_6209,N_4629,N_4927);
nand U6210 (N_6210,N_3077,N_2954);
and U6211 (N_6211,N_4766,N_3800);
or U6212 (N_6212,N_2547,N_4714);
nand U6213 (N_6213,N_3583,N_3115);
nor U6214 (N_6214,N_4653,N_3247);
and U6215 (N_6215,N_2553,N_2907);
nand U6216 (N_6216,N_3351,N_3981);
or U6217 (N_6217,N_4112,N_4921);
xnor U6218 (N_6218,N_2904,N_3072);
or U6219 (N_6219,N_4251,N_4182);
xor U6220 (N_6220,N_2900,N_4461);
or U6221 (N_6221,N_4359,N_4201);
nor U6222 (N_6222,N_3968,N_4042);
or U6223 (N_6223,N_3244,N_4821);
and U6224 (N_6224,N_4551,N_3858);
and U6225 (N_6225,N_3073,N_4111);
nor U6226 (N_6226,N_4154,N_3345);
and U6227 (N_6227,N_4029,N_2971);
nor U6228 (N_6228,N_3841,N_4420);
nand U6229 (N_6229,N_3877,N_4561);
or U6230 (N_6230,N_2992,N_3759);
nand U6231 (N_6231,N_4253,N_3488);
nor U6232 (N_6232,N_4328,N_4410);
xnor U6233 (N_6233,N_2679,N_3033);
or U6234 (N_6234,N_4404,N_2714);
xnor U6235 (N_6235,N_4670,N_4003);
nand U6236 (N_6236,N_2716,N_3856);
nor U6237 (N_6237,N_4857,N_4775);
or U6238 (N_6238,N_3845,N_2648);
or U6239 (N_6239,N_3065,N_4122);
and U6240 (N_6240,N_4758,N_3716);
xnor U6241 (N_6241,N_2710,N_4809);
xnor U6242 (N_6242,N_4902,N_3770);
nor U6243 (N_6243,N_3146,N_2507);
nand U6244 (N_6244,N_2914,N_3655);
nor U6245 (N_6245,N_4425,N_4091);
xnor U6246 (N_6246,N_2504,N_3930);
nor U6247 (N_6247,N_2699,N_4938);
xnor U6248 (N_6248,N_3720,N_3185);
nand U6249 (N_6249,N_3133,N_3045);
nor U6250 (N_6250,N_2907,N_2631);
nor U6251 (N_6251,N_4703,N_4682);
or U6252 (N_6252,N_4554,N_3141);
nand U6253 (N_6253,N_3285,N_3573);
xnor U6254 (N_6254,N_4925,N_3224);
xor U6255 (N_6255,N_2887,N_2773);
nand U6256 (N_6256,N_3756,N_4654);
nor U6257 (N_6257,N_4636,N_4474);
nor U6258 (N_6258,N_3869,N_3872);
and U6259 (N_6259,N_2615,N_4059);
and U6260 (N_6260,N_2759,N_3718);
and U6261 (N_6261,N_4209,N_3520);
and U6262 (N_6262,N_2996,N_3237);
or U6263 (N_6263,N_3008,N_4249);
or U6264 (N_6264,N_2866,N_3562);
or U6265 (N_6265,N_4753,N_3351);
or U6266 (N_6266,N_4815,N_3253);
nand U6267 (N_6267,N_3498,N_3573);
xor U6268 (N_6268,N_3007,N_2741);
xor U6269 (N_6269,N_3910,N_4126);
nor U6270 (N_6270,N_2848,N_4282);
or U6271 (N_6271,N_2967,N_4578);
or U6272 (N_6272,N_2909,N_4443);
nor U6273 (N_6273,N_3175,N_4624);
nor U6274 (N_6274,N_2967,N_4235);
xnor U6275 (N_6275,N_4184,N_4072);
and U6276 (N_6276,N_4405,N_4097);
or U6277 (N_6277,N_3390,N_4192);
xor U6278 (N_6278,N_3211,N_3841);
or U6279 (N_6279,N_3897,N_2935);
or U6280 (N_6280,N_4215,N_4709);
nand U6281 (N_6281,N_3654,N_4009);
and U6282 (N_6282,N_3066,N_3227);
or U6283 (N_6283,N_3004,N_2932);
nor U6284 (N_6284,N_3678,N_4027);
nand U6285 (N_6285,N_4818,N_4186);
or U6286 (N_6286,N_3157,N_3557);
nor U6287 (N_6287,N_3823,N_4196);
xor U6288 (N_6288,N_4427,N_4013);
nor U6289 (N_6289,N_4747,N_3349);
nor U6290 (N_6290,N_2649,N_3167);
and U6291 (N_6291,N_3185,N_4444);
nand U6292 (N_6292,N_4673,N_3621);
and U6293 (N_6293,N_3824,N_2814);
nand U6294 (N_6294,N_3962,N_2545);
nor U6295 (N_6295,N_2795,N_3026);
nor U6296 (N_6296,N_4431,N_3354);
nand U6297 (N_6297,N_4117,N_4912);
nor U6298 (N_6298,N_4633,N_4280);
xnor U6299 (N_6299,N_4079,N_3911);
or U6300 (N_6300,N_4520,N_3713);
nor U6301 (N_6301,N_4120,N_3912);
nor U6302 (N_6302,N_3943,N_2767);
nor U6303 (N_6303,N_4133,N_4558);
nand U6304 (N_6304,N_3395,N_2678);
and U6305 (N_6305,N_2853,N_3795);
or U6306 (N_6306,N_3427,N_3522);
or U6307 (N_6307,N_3851,N_4549);
xor U6308 (N_6308,N_4279,N_2933);
nand U6309 (N_6309,N_3195,N_3178);
xnor U6310 (N_6310,N_4405,N_4494);
and U6311 (N_6311,N_4553,N_3022);
nand U6312 (N_6312,N_4919,N_2676);
nor U6313 (N_6313,N_3012,N_2819);
and U6314 (N_6314,N_3707,N_2535);
and U6315 (N_6315,N_4544,N_4401);
nor U6316 (N_6316,N_2595,N_3824);
xor U6317 (N_6317,N_4516,N_4281);
xnor U6318 (N_6318,N_4535,N_4074);
nor U6319 (N_6319,N_4130,N_2618);
xor U6320 (N_6320,N_4205,N_4606);
nand U6321 (N_6321,N_2608,N_4429);
nand U6322 (N_6322,N_4984,N_2930);
nand U6323 (N_6323,N_3877,N_3347);
xor U6324 (N_6324,N_4417,N_3714);
and U6325 (N_6325,N_3455,N_4223);
and U6326 (N_6326,N_2916,N_4804);
nor U6327 (N_6327,N_2617,N_3186);
nor U6328 (N_6328,N_4368,N_4245);
or U6329 (N_6329,N_3498,N_3121);
nor U6330 (N_6330,N_2891,N_4925);
xnor U6331 (N_6331,N_4757,N_4358);
nor U6332 (N_6332,N_3031,N_2741);
nand U6333 (N_6333,N_4323,N_3943);
or U6334 (N_6334,N_3192,N_2573);
nor U6335 (N_6335,N_2616,N_3448);
or U6336 (N_6336,N_3237,N_2774);
nor U6337 (N_6337,N_4850,N_4348);
nand U6338 (N_6338,N_4331,N_3674);
and U6339 (N_6339,N_3214,N_4511);
nand U6340 (N_6340,N_2813,N_3131);
nor U6341 (N_6341,N_4542,N_4789);
nor U6342 (N_6342,N_2691,N_3872);
and U6343 (N_6343,N_3034,N_3145);
and U6344 (N_6344,N_4683,N_4068);
and U6345 (N_6345,N_4325,N_4326);
and U6346 (N_6346,N_2543,N_3806);
xor U6347 (N_6347,N_4676,N_4403);
and U6348 (N_6348,N_2827,N_4719);
nand U6349 (N_6349,N_3778,N_4043);
nor U6350 (N_6350,N_2548,N_2953);
or U6351 (N_6351,N_4957,N_4621);
xnor U6352 (N_6352,N_4218,N_3015);
nand U6353 (N_6353,N_2912,N_3353);
nor U6354 (N_6354,N_4820,N_3614);
or U6355 (N_6355,N_4503,N_4327);
and U6356 (N_6356,N_4027,N_4175);
nand U6357 (N_6357,N_4056,N_3331);
nor U6358 (N_6358,N_4813,N_4525);
and U6359 (N_6359,N_3926,N_2865);
xor U6360 (N_6360,N_3868,N_4093);
xor U6361 (N_6361,N_3431,N_4219);
or U6362 (N_6362,N_3839,N_3957);
nor U6363 (N_6363,N_3918,N_2740);
or U6364 (N_6364,N_4164,N_3570);
nand U6365 (N_6365,N_2864,N_2947);
and U6366 (N_6366,N_4145,N_4038);
nand U6367 (N_6367,N_3663,N_2521);
and U6368 (N_6368,N_2739,N_2540);
or U6369 (N_6369,N_4150,N_3424);
xor U6370 (N_6370,N_3028,N_3899);
nand U6371 (N_6371,N_4842,N_2947);
and U6372 (N_6372,N_3509,N_4709);
nand U6373 (N_6373,N_3029,N_4319);
or U6374 (N_6374,N_4412,N_4012);
or U6375 (N_6375,N_3047,N_3429);
or U6376 (N_6376,N_4978,N_3812);
nand U6377 (N_6377,N_3722,N_4410);
or U6378 (N_6378,N_3030,N_3762);
xor U6379 (N_6379,N_4462,N_3695);
and U6380 (N_6380,N_4583,N_4702);
xor U6381 (N_6381,N_3807,N_4571);
xnor U6382 (N_6382,N_3294,N_2904);
nand U6383 (N_6383,N_4130,N_4112);
nor U6384 (N_6384,N_3014,N_3264);
or U6385 (N_6385,N_2643,N_4721);
or U6386 (N_6386,N_4815,N_4947);
nand U6387 (N_6387,N_2662,N_3652);
nor U6388 (N_6388,N_4999,N_3614);
nand U6389 (N_6389,N_3344,N_2900);
xor U6390 (N_6390,N_3258,N_2993);
nand U6391 (N_6391,N_4224,N_3819);
and U6392 (N_6392,N_3910,N_4698);
xor U6393 (N_6393,N_3190,N_4606);
and U6394 (N_6394,N_2512,N_4693);
nor U6395 (N_6395,N_4038,N_4690);
or U6396 (N_6396,N_3864,N_2558);
and U6397 (N_6397,N_3176,N_3503);
xor U6398 (N_6398,N_3062,N_4738);
nand U6399 (N_6399,N_3177,N_2845);
and U6400 (N_6400,N_4522,N_3122);
and U6401 (N_6401,N_4614,N_4262);
nor U6402 (N_6402,N_4759,N_2608);
and U6403 (N_6403,N_3702,N_4493);
xor U6404 (N_6404,N_3731,N_3844);
nor U6405 (N_6405,N_3837,N_3280);
nand U6406 (N_6406,N_4647,N_3228);
and U6407 (N_6407,N_4989,N_2870);
and U6408 (N_6408,N_2904,N_3403);
and U6409 (N_6409,N_4632,N_3421);
xnor U6410 (N_6410,N_3769,N_4118);
nand U6411 (N_6411,N_3916,N_2982);
nor U6412 (N_6412,N_3593,N_2648);
and U6413 (N_6413,N_4136,N_3228);
nand U6414 (N_6414,N_2763,N_4891);
nor U6415 (N_6415,N_4085,N_4339);
and U6416 (N_6416,N_3059,N_4879);
xor U6417 (N_6417,N_4448,N_3480);
nand U6418 (N_6418,N_3785,N_3817);
or U6419 (N_6419,N_4905,N_3900);
and U6420 (N_6420,N_3557,N_3668);
xnor U6421 (N_6421,N_4833,N_4989);
nand U6422 (N_6422,N_4589,N_3082);
or U6423 (N_6423,N_2874,N_3481);
nor U6424 (N_6424,N_4449,N_4734);
nor U6425 (N_6425,N_3740,N_4422);
nand U6426 (N_6426,N_3303,N_2630);
and U6427 (N_6427,N_3977,N_4083);
or U6428 (N_6428,N_3651,N_4434);
nor U6429 (N_6429,N_2795,N_4718);
nor U6430 (N_6430,N_3066,N_4003);
nor U6431 (N_6431,N_3034,N_3153);
and U6432 (N_6432,N_3604,N_4035);
and U6433 (N_6433,N_4891,N_3547);
or U6434 (N_6434,N_4299,N_4053);
nor U6435 (N_6435,N_2972,N_3092);
nor U6436 (N_6436,N_2940,N_3756);
nand U6437 (N_6437,N_4694,N_4530);
nand U6438 (N_6438,N_2566,N_3384);
and U6439 (N_6439,N_3853,N_4644);
xor U6440 (N_6440,N_3219,N_4764);
or U6441 (N_6441,N_3847,N_3799);
or U6442 (N_6442,N_2827,N_3514);
nand U6443 (N_6443,N_4303,N_4360);
or U6444 (N_6444,N_3367,N_2950);
nor U6445 (N_6445,N_4586,N_3810);
nand U6446 (N_6446,N_2881,N_4468);
xnor U6447 (N_6447,N_4232,N_4222);
and U6448 (N_6448,N_3439,N_2575);
xor U6449 (N_6449,N_3166,N_2967);
nor U6450 (N_6450,N_4004,N_3555);
nor U6451 (N_6451,N_4681,N_3829);
xor U6452 (N_6452,N_4596,N_4483);
nor U6453 (N_6453,N_3583,N_4609);
and U6454 (N_6454,N_2986,N_3417);
nand U6455 (N_6455,N_4989,N_3047);
and U6456 (N_6456,N_4419,N_3025);
xor U6457 (N_6457,N_4799,N_2861);
nor U6458 (N_6458,N_3379,N_3277);
and U6459 (N_6459,N_3024,N_2654);
nor U6460 (N_6460,N_3680,N_4865);
nand U6461 (N_6461,N_2577,N_3627);
or U6462 (N_6462,N_2685,N_3299);
nor U6463 (N_6463,N_3815,N_3057);
and U6464 (N_6464,N_3318,N_3273);
nand U6465 (N_6465,N_3026,N_4786);
nand U6466 (N_6466,N_3834,N_4002);
xnor U6467 (N_6467,N_4437,N_4824);
xnor U6468 (N_6468,N_3504,N_3649);
nor U6469 (N_6469,N_4968,N_3081);
nor U6470 (N_6470,N_2843,N_2913);
xnor U6471 (N_6471,N_4861,N_2729);
and U6472 (N_6472,N_4406,N_3409);
or U6473 (N_6473,N_2813,N_4069);
and U6474 (N_6474,N_2531,N_4194);
nor U6475 (N_6475,N_4493,N_3907);
nand U6476 (N_6476,N_2639,N_2844);
nor U6477 (N_6477,N_4919,N_4887);
or U6478 (N_6478,N_3720,N_2818);
and U6479 (N_6479,N_2535,N_2717);
xnor U6480 (N_6480,N_4101,N_2674);
or U6481 (N_6481,N_2612,N_3392);
or U6482 (N_6482,N_4837,N_3924);
nor U6483 (N_6483,N_4478,N_4911);
or U6484 (N_6484,N_4680,N_3488);
nand U6485 (N_6485,N_4386,N_3093);
nand U6486 (N_6486,N_3034,N_3795);
nand U6487 (N_6487,N_3374,N_3378);
nor U6488 (N_6488,N_4372,N_3714);
or U6489 (N_6489,N_2806,N_3971);
and U6490 (N_6490,N_2900,N_3228);
and U6491 (N_6491,N_3425,N_3444);
xnor U6492 (N_6492,N_2969,N_2717);
and U6493 (N_6493,N_3074,N_2676);
or U6494 (N_6494,N_4066,N_4190);
or U6495 (N_6495,N_2993,N_3230);
and U6496 (N_6496,N_4103,N_3318);
nor U6497 (N_6497,N_3266,N_2503);
nor U6498 (N_6498,N_3366,N_4256);
and U6499 (N_6499,N_4214,N_3535);
nand U6500 (N_6500,N_4464,N_3490);
nand U6501 (N_6501,N_3392,N_2985);
and U6502 (N_6502,N_3411,N_2750);
nand U6503 (N_6503,N_4458,N_3426);
or U6504 (N_6504,N_4090,N_2650);
nand U6505 (N_6505,N_3422,N_4412);
nand U6506 (N_6506,N_4542,N_2967);
or U6507 (N_6507,N_4215,N_4077);
and U6508 (N_6508,N_4399,N_2865);
xor U6509 (N_6509,N_3274,N_3765);
nand U6510 (N_6510,N_4659,N_4253);
and U6511 (N_6511,N_4657,N_3954);
xnor U6512 (N_6512,N_2954,N_3157);
or U6513 (N_6513,N_3782,N_2511);
and U6514 (N_6514,N_2685,N_2516);
nor U6515 (N_6515,N_3248,N_3176);
xnor U6516 (N_6516,N_4638,N_4949);
nand U6517 (N_6517,N_3980,N_3892);
or U6518 (N_6518,N_2649,N_4536);
nand U6519 (N_6519,N_3721,N_4631);
nand U6520 (N_6520,N_4818,N_4037);
and U6521 (N_6521,N_4284,N_3176);
nor U6522 (N_6522,N_3045,N_2585);
and U6523 (N_6523,N_4710,N_4611);
and U6524 (N_6524,N_4483,N_4634);
and U6525 (N_6525,N_3217,N_3013);
nor U6526 (N_6526,N_2851,N_3996);
xor U6527 (N_6527,N_4664,N_4962);
or U6528 (N_6528,N_4263,N_4763);
nor U6529 (N_6529,N_3231,N_3346);
nand U6530 (N_6530,N_4866,N_3804);
and U6531 (N_6531,N_4678,N_3384);
nand U6532 (N_6532,N_2697,N_2900);
nand U6533 (N_6533,N_4109,N_4558);
xor U6534 (N_6534,N_4377,N_3784);
and U6535 (N_6535,N_3788,N_4949);
or U6536 (N_6536,N_2671,N_3622);
nor U6537 (N_6537,N_4316,N_4223);
or U6538 (N_6538,N_3289,N_4641);
nor U6539 (N_6539,N_2785,N_3673);
and U6540 (N_6540,N_4449,N_4937);
nand U6541 (N_6541,N_2959,N_4040);
and U6542 (N_6542,N_2855,N_3586);
or U6543 (N_6543,N_2749,N_2714);
and U6544 (N_6544,N_4886,N_4629);
nand U6545 (N_6545,N_4384,N_4644);
nor U6546 (N_6546,N_3968,N_2828);
and U6547 (N_6547,N_3494,N_2933);
or U6548 (N_6548,N_2903,N_3356);
xor U6549 (N_6549,N_4565,N_4344);
xor U6550 (N_6550,N_4704,N_4432);
and U6551 (N_6551,N_2886,N_3008);
or U6552 (N_6552,N_4232,N_3495);
xor U6553 (N_6553,N_4767,N_3385);
or U6554 (N_6554,N_4674,N_4978);
and U6555 (N_6555,N_3004,N_4181);
nor U6556 (N_6556,N_3033,N_2510);
and U6557 (N_6557,N_4759,N_2601);
nor U6558 (N_6558,N_2600,N_4185);
nand U6559 (N_6559,N_3912,N_4898);
nor U6560 (N_6560,N_3629,N_4733);
nand U6561 (N_6561,N_3436,N_2742);
and U6562 (N_6562,N_4455,N_3438);
nand U6563 (N_6563,N_3908,N_4598);
and U6564 (N_6564,N_4914,N_4356);
and U6565 (N_6565,N_3790,N_2750);
nor U6566 (N_6566,N_4459,N_4538);
xnor U6567 (N_6567,N_2871,N_3834);
or U6568 (N_6568,N_3832,N_4266);
nor U6569 (N_6569,N_3105,N_3005);
nand U6570 (N_6570,N_4805,N_4169);
and U6571 (N_6571,N_3740,N_3520);
nand U6572 (N_6572,N_3917,N_3568);
nor U6573 (N_6573,N_4136,N_3957);
nand U6574 (N_6574,N_4876,N_3437);
and U6575 (N_6575,N_2865,N_3284);
nand U6576 (N_6576,N_2872,N_3368);
and U6577 (N_6577,N_4291,N_2809);
nor U6578 (N_6578,N_2780,N_3762);
nand U6579 (N_6579,N_3633,N_4422);
nor U6580 (N_6580,N_4534,N_3013);
xnor U6581 (N_6581,N_2503,N_3145);
or U6582 (N_6582,N_4987,N_2845);
and U6583 (N_6583,N_2838,N_3853);
and U6584 (N_6584,N_3713,N_3717);
or U6585 (N_6585,N_2689,N_2545);
and U6586 (N_6586,N_4840,N_3824);
and U6587 (N_6587,N_4335,N_2760);
xnor U6588 (N_6588,N_4789,N_2515);
and U6589 (N_6589,N_3273,N_4797);
nor U6590 (N_6590,N_4516,N_4667);
and U6591 (N_6591,N_3905,N_3368);
nor U6592 (N_6592,N_4738,N_3240);
or U6593 (N_6593,N_2728,N_3549);
xor U6594 (N_6594,N_4211,N_3054);
xnor U6595 (N_6595,N_3875,N_4833);
and U6596 (N_6596,N_2767,N_3070);
nor U6597 (N_6597,N_2996,N_3812);
nand U6598 (N_6598,N_2993,N_4855);
nand U6599 (N_6599,N_3098,N_2957);
and U6600 (N_6600,N_3818,N_3271);
and U6601 (N_6601,N_4447,N_2892);
nor U6602 (N_6602,N_3742,N_3306);
xor U6603 (N_6603,N_4400,N_4276);
nand U6604 (N_6604,N_4401,N_4214);
and U6605 (N_6605,N_4246,N_2888);
and U6606 (N_6606,N_4331,N_3621);
nor U6607 (N_6607,N_2550,N_4338);
nor U6608 (N_6608,N_4523,N_4337);
xor U6609 (N_6609,N_3654,N_4480);
or U6610 (N_6610,N_4027,N_3863);
or U6611 (N_6611,N_2819,N_4549);
nand U6612 (N_6612,N_3964,N_3745);
nor U6613 (N_6613,N_3294,N_4817);
and U6614 (N_6614,N_3759,N_3290);
xor U6615 (N_6615,N_3264,N_4437);
xnor U6616 (N_6616,N_2504,N_4624);
or U6617 (N_6617,N_3947,N_2755);
or U6618 (N_6618,N_3626,N_4811);
xnor U6619 (N_6619,N_4428,N_4107);
or U6620 (N_6620,N_2620,N_4695);
and U6621 (N_6621,N_3213,N_4394);
and U6622 (N_6622,N_3884,N_4943);
nor U6623 (N_6623,N_4114,N_4014);
nor U6624 (N_6624,N_3609,N_2679);
nor U6625 (N_6625,N_3816,N_4068);
xor U6626 (N_6626,N_3547,N_3670);
nand U6627 (N_6627,N_3253,N_4785);
nand U6628 (N_6628,N_4829,N_2927);
nor U6629 (N_6629,N_2576,N_4346);
or U6630 (N_6630,N_4932,N_4986);
nand U6631 (N_6631,N_4622,N_2656);
xnor U6632 (N_6632,N_3014,N_3805);
and U6633 (N_6633,N_2597,N_4777);
or U6634 (N_6634,N_4729,N_2943);
xor U6635 (N_6635,N_2724,N_3266);
and U6636 (N_6636,N_3220,N_2989);
or U6637 (N_6637,N_2799,N_3223);
xnor U6638 (N_6638,N_2963,N_2549);
nor U6639 (N_6639,N_3000,N_2972);
nand U6640 (N_6640,N_3662,N_3403);
nor U6641 (N_6641,N_4009,N_3108);
nand U6642 (N_6642,N_3829,N_3893);
or U6643 (N_6643,N_2984,N_3639);
or U6644 (N_6644,N_4366,N_4780);
and U6645 (N_6645,N_2973,N_4019);
nor U6646 (N_6646,N_3238,N_3089);
and U6647 (N_6647,N_4510,N_3149);
nand U6648 (N_6648,N_3394,N_4478);
nor U6649 (N_6649,N_4124,N_2564);
nand U6650 (N_6650,N_4961,N_4739);
xnor U6651 (N_6651,N_3368,N_3774);
xnor U6652 (N_6652,N_2555,N_4774);
xnor U6653 (N_6653,N_3747,N_4743);
nor U6654 (N_6654,N_4468,N_4970);
nor U6655 (N_6655,N_4898,N_2721);
and U6656 (N_6656,N_4505,N_3562);
or U6657 (N_6657,N_2591,N_3311);
nor U6658 (N_6658,N_2778,N_2793);
and U6659 (N_6659,N_4207,N_4164);
nand U6660 (N_6660,N_3064,N_3257);
and U6661 (N_6661,N_3286,N_3247);
nor U6662 (N_6662,N_2835,N_4994);
xor U6663 (N_6663,N_2674,N_3130);
nor U6664 (N_6664,N_3817,N_3201);
or U6665 (N_6665,N_2583,N_4116);
and U6666 (N_6666,N_2959,N_4213);
nand U6667 (N_6667,N_3949,N_4074);
xnor U6668 (N_6668,N_3148,N_2934);
or U6669 (N_6669,N_3371,N_2614);
nor U6670 (N_6670,N_3435,N_4080);
or U6671 (N_6671,N_3309,N_3224);
nor U6672 (N_6672,N_3639,N_3641);
nand U6673 (N_6673,N_3627,N_4902);
xor U6674 (N_6674,N_3366,N_2694);
xor U6675 (N_6675,N_4127,N_4054);
and U6676 (N_6676,N_2798,N_3752);
nand U6677 (N_6677,N_3494,N_3084);
xor U6678 (N_6678,N_4002,N_2512);
xnor U6679 (N_6679,N_4028,N_4447);
or U6680 (N_6680,N_3764,N_2852);
or U6681 (N_6681,N_2590,N_3977);
or U6682 (N_6682,N_4725,N_4119);
xnor U6683 (N_6683,N_4771,N_2672);
xnor U6684 (N_6684,N_3890,N_2926);
nand U6685 (N_6685,N_4480,N_4662);
nor U6686 (N_6686,N_4324,N_3706);
nor U6687 (N_6687,N_3095,N_2510);
nand U6688 (N_6688,N_4942,N_4015);
xor U6689 (N_6689,N_3201,N_2946);
xor U6690 (N_6690,N_4008,N_4407);
xnor U6691 (N_6691,N_3951,N_2736);
xnor U6692 (N_6692,N_3205,N_4854);
or U6693 (N_6693,N_3718,N_3613);
xor U6694 (N_6694,N_2718,N_4056);
xnor U6695 (N_6695,N_2659,N_4003);
xnor U6696 (N_6696,N_4916,N_3453);
xor U6697 (N_6697,N_2893,N_4423);
and U6698 (N_6698,N_3660,N_2608);
nand U6699 (N_6699,N_3815,N_3318);
nor U6700 (N_6700,N_4638,N_3658);
nor U6701 (N_6701,N_4283,N_3745);
and U6702 (N_6702,N_4274,N_4933);
xnor U6703 (N_6703,N_4796,N_4452);
and U6704 (N_6704,N_2716,N_3509);
or U6705 (N_6705,N_2501,N_2557);
or U6706 (N_6706,N_4859,N_3203);
or U6707 (N_6707,N_4585,N_4502);
nand U6708 (N_6708,N_3069,N_4696);
and U6709 (N_6709,N_3048,N_3738);
nor U6710 (N_6710,N_3775,N_2933);
xor U6711 (N_6711,N_2833,N_3368);
and U6712 (N_6712,N_3614,N_2907);
nand U6713 (N_6713,N_2928,N_2549);
xor U6714 (N_6714,N_2556,N_3968);
nor U6715 (N_6715,N_2526,N_3006);
or U6716 (N_6716,N_4990,N_2743);
nor U6717 (N_6717,N_2997,N_4225);
nand U6718 (N_6718,N_2664,N_2726);
nand U6719 (N_6719,N_4062,N_3647);
nor U6720 (N_6720,N_3676,N_3581);
nand U6721 (N_6721,N_4304,N_3853);
and U6722 (N_6722,N_3508,N_3600);
nand U6723 (N_6723,N_4430,N_3000);
nor U6724 (N_6724,N_3946,N_2915);
nand U6725 (N_6725,N_3106,N_4101);
xnor U6726 (N_6726,N_3001,N_2741);
nand U6727 (N_6727,N_4648,N_4966);
nor U6728 (N_6728,N_4879,N_3291);
and U6729 (N_6729,N_4373,N_4274);
and U6730 (N_6730,N_3551,N_3018);
nor U6731 (N_6731,N_2662,N_3491);
nand U6732 (N_6732,N_3383,N_3686);
nor U6733 (N_6733,N_4779,N_2524);
or U6734 (N_6734,N_3625,N_2624);
nor U6735 (N_6735,N_3800,N_3946);
or U6736 (N_6736,N_4140,N_3005);
nand U6737 (N_6737,N_3793,N_3024);
nand U6738 (N_6738,N_4081,N_4104);
nor U6739 (N_6739,N_4218,N_4184);
nor U6740 (N_6740,N_3670,N_3018);
nor U6741 (N_6741,N_4250,N_4835);
nand U6742 (N_6742,N_4620,N_4860);
xor U6743 (N_6743,N_3175,N_3061);
nand U6744 (N_6744,N_4436,N_2668);
nand U6745 (N_6745,N_3460,N_3928);
and U6746 (N_6746,N_2972,N_4767);
nand U6747 (N_6747,N_2509,N_3569);
and U6748 (N_6748,N_3033,N_3383);
xnor U6749 (N_6749,N_2919,N_2823);
or U6750 (N_6750,N_4888,N_4159);
or U6751 (N_6751,N_2641,N_4511);
xnor U6752 (N_6752,N_2979,N_4039);
or U6753 (N_6753,N_3643,N_4486);
or U6754 (N_6754,N_3768,N_3895);
nor U6755 (N_6755,N_4216,N_2548);
xor U6756 (N_6756,N_3308,N_3671);
nor U6757 (N_6757,N_2513,N_4520);
nor U6758 (N_6758,N_2817,N_3560);
xnor U6759 (N_6759,N_2715,N_4681);
or U6760 (N_6760,N_4087,N_3380);
nor U6761 (N_6761,N_4167,N_3580);
nand U6762 (N_6762,N_4189,N_3737);
and U6763 (N_6763,N_4857,N_3234);
nand U6764 (N_6764,N_4436,N_3722);
and U6765 (N_6765,N_4235,N_4242);
or U6766 (N_6766,N_2789,N_4654);
and U6767 (N_6767,N_4192,N_4028);
xor U6768 (N_6768,N_3872,N_3773);
nor U6769 (N_6769,N_4273,N_4539);
xnor U6770 (N_6770,N_3431,N_3412);
xnor U6771 (N_6771,N_3441,N_3457);
or U6772 (N_6772,N_3091,N_2704);
nand U6773 (N_6773,N_2982,N_4929);
or U6774 (N_6774,N_4234,N_4639);
nand U6775 (N_6775,N_3381,N_3105);
or U6776 (N_6776,N_2713,N_2821);
nand U6777 (N_6777,N_4257,N_4302);
xnor U6778 (N_6778,N_3816,N_4565);
nor U6779 (N_6779,N_3417,N_2800);
and U6780 (N_6780,N_3422,N_4589);
nand U6781 (N_6781,N_4960,N_2691);
nand U6782 (N_6782,N_4722,N_2979);
nor U6783 (N_6783,N_2735,N_4382);
xor U6784 (N_6784,N_2974,N_3638);
or U6785 (N_6785,N_3856,N_4723);
nand U6786 (N_6786,N_4165,N_4162);
and U6787 (N_6787,N_4386,N_3507);
or U6788 (N_6788,N_2796,N_4957);
and U6789 (N_6789,N_4094,N_4189);
nand U6790 (N_6790,N_4910,N_2812);
nand U6791 (N_6791,N_2686,N_4910);
or U6792 (N_6792,N_4971,N_4243);
nand U6793 (N_6793,N_3227,N_3762);
nand U6794 (N_6794,N_2848,N_4241);
nor U6795 (N_6795,N_3082,N_2951);
or U6796 (N_6796,N_3610,N_3857);
or U6797 (N_6797,N_4543,N_2683);
xnor U6798 (N_6798,N_4654,N_4480);
and U6799 (N_6799,N_3551,N_3324);
or U6800 (N_6800,N_3122,N_4758);
or U6801 (N_6801,N_4290,N_3208);
nand U6802 (N_6802,N_4921,N_3485);
nor U6803 (N_6803,N_4228,N_3053);
nand U6804 (N_6804,N_2546,N_2670);
xor U6805 (N_6805,N_4061,N_3089);
and U6806 (N_6806,N_4662,N_3115);
nor U6807 (N_6807,N_2879,N_3976);
and U6808 (N_6808,N_4689,N_4156);
nor U6809 (N_6809,N_4899,N_2683);
nand U6810 (N_6810,N_4275,N_3236);
and U6811 (N_6811,N_2522,N_4825);
nand U6812 (N_6812,N_2933,N_2657);
or U6813 (N_6813,N_4013,N_3196);
xnor U6814 (N_6814,N_3404,N_3340);
nand U6815 (N_6815,N_3530,N_4411);
and U6816 (N_6816,N_3641,N_3528);
or U6817 (N_6817,N_3753,N_2798);
nand U6818 (N_6818,N_3259,N_3501);
nor U6819 (N_6819,N_4164,N_3659);
xor U6820 (N_6820,N_4502,N_3620);
or U6821 (N_6821,N_4400,N_4971);
and U6822 (N_6822,N_2751,N_4951);
or U6823 (N_6823,N_2990,N_2739);
or U6824 (N_6824,N_3678,N_3388);
xor U6825 (N_6825,N_3316,N_3999);
nor U6826 (N_6826,N_4836,N_2919);
or U6827 (N_6827,N_2898,N_4373);
nor U6828 (N_6828,N_4039,N_4207);
nand U6829 (N_6829,N_4794,N_3150);
nand U6830 (N_6830,N_3474,N_3659);
and U6831 (N_6831,N_3637,N_3380);
or U6832 (N_6832,N_3174,N_3850);
nand U6833 (N_6833,N_4500,N_2585);
xor U6834 (N_6834,N_2871,N_4788);
and U6835 (N_6835,N_3618,N_4476);
nand U6836 (N_6836,N_3295,N_2915);
nor U6837 (N_6837,N_3841,N_4354);
and U6838 (N_6838,N_3406,N_4391);
nor U6839 (N_6839,N_4304,N_4210);
xnor U6840 (N_6840,N_3637,N_3961);
and U6841 (N_6841,N_3022,N_3854);
nand U6842 (N_6842,N_3813,N_4650);
xnor U6843 (N_6843,N_2884,N_4585);
nand U6844 (N_6844,N_2896,N_3540);
and U6845 (N_6845,N_4972,N_2606);
xnor U6846 (N_6846,N_3853,N_3388);
xnor U6847 (N_6847,N_4955,N_2716);
or U6848 (N_6848,N_3509,N_2629);
or U6849 (N_6849,N_4605,N_3622);
and U6850 (N_6850,N_3508,N_4255);
nor U6851 (N_6851,N_4124,N_3981);
and U6852 (N_6852,N_3914,N_2601);
nand U6853 (N_6853,N_4141,N_4910);
or U6854 (N_6854,N_3512,N_4929);
or U6855 (N_6855,N_3931,N_4145);
and U6856 (N_6856,N_3591,N_3774);
xor U6857 (N_6857,N_3273,N_3868);
nand U6858 (N_6858,N_3668,N_3746);
xnor U6859 (N_6859,N_4283,N_4195);
and U6860 (N_6860,N_3495,N_2523);
nor U6861 (N_6861,N_4584,N_4238);
nand U6862 (N_6862,N_3526,N_4580);
xnor U6863 (N_6863,N_3640,N_4105);
nor U6864 (N_6864,N_3763,N_4674);
or U6865 (N_6865,N_2597,N_3965);
and U6866 (N_6866,N_2523,N_2841);
and U6867 (N_6867,N_3211,N_3933);
or U6868 (N_6868,N_3586,N_3756);
and U6869 (N_6869,N_2702,N_4476);
xnor U6870 (N_6870,N_2559,N_4083);
and U6871 (N_6871,N_4218,N_3096);
xnor U6872 (N_6872,N_3751,N_4308);
nand U6873 (N_6873,N_3243,N_2989);
xnor U6874 (N_6874,N_3726,N_3756);
xnor U6875 (N_6875,N_4554,N_3321);
nand U6876 (N_6876,N_4276,N_3180);
xor U6877 (N_6877,N_2672,N_3683);
or U6878 (N_6878,N_4980,N_3123);
nand U6879 (N_6879,N_2885,N_4627);
nand U6880 (N_6880,N_3777,N_2706);
nand U6881 (N_6881,N_3308,N_3504);
nand U6882 (N_6882,N_3434,N_4784);
nand U6883 (N_6883,N_3314,N_4725);
nor U6884 (N_6884,N_3064,N_2524);
xnor U6885 (N_6885,N_3957,N_4966);
and U6886 (N_6886,N_3331,N_2640);
nor U6887 (N_6887,N_3941,N_3069);
nor U6888 (N_6888,N_3530,N_4987);
nor U6889 (N_6889,N_4557,N_3098);
and U6890 (N_6890,N_4629,N_4192);
xor U6891 (N_6891,N_3024,N_3619);
xnor U6892 (N_6892,N_4193,N_3154);
and U6893 (N_6893,N_3347,N_4108);
nand U6894 (N_6894,N_4957,N_3621);
nand U6895 (N_6895,N_2612,N_4406);
and U6896 (N_6896,N_4249,N_2825);
and U6897 (N_6897,N_4035,N_2625);
nand U6898 (N_6898,N_4884,N_2708);
nand U6899 (N_6899,N_4733,N_3589);
and U6900 (N_6900,N_4111,N_3410);
nand U6901 (N_6901,N_4274,N_3237);
or U6902 (N_6902,N_3532,N_4609);
and U6903 (N_6903,N_3309,N_3105);
and U6904 (N_6904,N_4093,N_2764);
xnor U6905 (N_6905,N_2713,N_4943);
xor U6906 (N_6906,N_4975,N_3481);
or U6907 (N_6907,N_2842,N_4600);
and U6908 (N_6908,N_4486,N_3357);
nand U6909 (N_6909,N_3155,N_3921);
and U6910 (N_6910,N_4889,N_3342);
and U6911 (N_6911,N_2546,N_3096);
or U6912 (N_6912,N_4970,N_3594);
nor U6913 (N_6913,N_4496,N_2733);
nor U6914 (N_6914,N_2735,N_4481);
and U6915 (N_6915,N_3485,N_3666);
or U6916 (N_6916,N_2931,N_4455);
or U6917 (N_6917,N_4427,N_3804);
nor U6918 (N_6918,N_3453,N_3553);
or U6919 (N_6919,N_4280,N_4423);
xor U6920 (N_6920,N_4763,N_3851);
nor U6921 (N_6921,N_3700,N_4451);
and U6922 (N_6922,N_4915,N_3600);
nand U6923 (N_6923,N_4904,N_2944);
xnor U6924 (N_6924,N_4930,N_3506);
and U6925 (N_6925,N_4410,N_2668);
xnor U6926 (N_6926,N_4416,N_2585);
and U6927 (N_6927,N_3320,N_3214);
or U6928 (N_6928,N_4311,N_2799);
and U6929 (N_6929,N_4315,N_4384);
or U6930 (N_6930,N_4930,N_3494);
nand U6931 (N_6931,N_4057,N_3217);
xnor U6932 (N_6932,N_2908,N_3191);
and U6933 (N_6933,N_4656,N_4716);
or U6934 (N_6934,N_2774,N_4806);
nand U6935 (N_6935,N_2657,N_2647);
nor U6936 (N_6936,N_4588,N_3668);
and U6937 (N_6937,N_3875,N_3735);
nor U6938 (N_6938,N_4380,N_4113);
and U6939 (N_6939,N_4304,N_2942);
or U6940 (N_6940,N_3144,N_4756);
nand U6941 (N_6941,N_2816,N_4586);
xnor U6942 (N_6942,N_4344,N_3309);
nand U6943 (N_6943,N_3412,N_4456);
xor U6944 (N_6944,N_3664,N_4044);
xnor U6945 (N_6945,N_4412,N_3864);
and U6946 (N_6946,N_3283,N_3589);
xnor U6947 (N_6947,N_3552,N_3683);
and U6948 (N_6948,N_4572,N_4924);
or U6949 (N_6949,N_2560,N_3439);
and U6950 (N_6950,N_4073,N_4268);
xnor U6951 (N_6951,N_3679,N_3779);
nand U6952 (N_6952,N_2951,N_2966);
or U6953 (N_6953,N_4164,N_4959);
or U6954 (N_6954,N_3991,N_3027);
xnor U6955 (N_6955,N_4914,N_3111);
or U6956 (N_6956,N_3707,N_3115);
or U6957 (N_6957,N_4244,N_3301);
xor U6958 (N_6958,N_3977,N_3703);
xor U6959 (N_6959,N_4786,N_3453);
nor U6960 (N_6960,N_4481,N_2828);
nand U6961 (N_6961,N_4781,N_2764);
and U6962 (N_6962,N_2874,N_4381);
nor U6963 (N_6963,N_4527,N_4014);
nor U6964 (N_6964,N_4600,N_2705);
and U6965 (N_6965,N_3760,N_2601);
xor U6966 (N_6966,N_4042,N_3327);
or U6967 (N_6967,N_3592,N_3714);
xor U6968 (N_6968,N_4797,N_2942);
and U6969 (N_6969,N_2688,N_3838);
nand U6970 (N_6970,N_4101,N_3460);
nor U6971 (N_6971,N_4590,N_4348);
or U6972 (N_6972,N_3004,N_3454);
xnor U6973 (N_6973,N_2959,N_3924);
nand U6974 (N_6974,N_4825,N_3542);
nand U6975 (N_6975,N_4232,N_4522);
and U6976 (N_6976,N_3755,N_3084);
xnor U6977 (N_6977,N_4111,N_4854);
xnor U6978 (N_6978,N_3402,N_2548);
xnor U6979 (N_6979,N_3563,N_4343);
nand U6980 (N_6980,N_3839,N_4311);
or U6981 (N_6981,N_3838,N_3439);
xnor U6982 (N_6982,N_3072,N_3375);
nor U6983 (N_6983,N_4473,N_2658);
nand U6984 (N_6984,N_2689,N_3219);
nand U6985 (N_6985,N_3168,N_4606);
nand U6986 (N_6986,N_4984,N_3040);
nor U6987 (N_6987,N_3614,N_4394);
xor U6988 (N_6988,N_4242,N_4806);
xnor U6989 (N_6989,N_4843,N_4882);
and U6990 (N_6990,N_4859,N_3907);
and U6991 (N_6991,N_4380,N_4846);
xnor U6992 (N_6992,N_3044,N_3529);
or U6993 (N_6993,N_4511,N_4402);
xnor U6994 (N_6994,N_3816,N_4081);
xor U6995 (N_6995,N_4900,N_2996);
xor U6996 (N_6996,N_4411,N_4955);
nor U6997 (N_6997,N_2903,N_3580);
nor U6998 (N_6998,N_4881,N_3651);
and U6999 (N_6999,N_2661,N_4112);
nor U7000 (N_7000,N_4337,N_4922);
or U7001 (N_7001,N_4120,N_2619);
nor U7002 (N_7002,N_3997,N_3751);
and U7003 (N_7003,N_3386,N_4261);
or U7004 (N_7004,N_3469,N_4529);
and U7005 (N_7005,N_3314,N_3624);
xnor U7006 (N_7006,N_3990,N_3906);
or U7007 (N_7007,N_2969,N_3385);
or U7008 (N_7008,N_4812,N_3551);
or U7009 (N_7009,N_4140,N_4771);
xor U7010 (N_7010,N_3085,N_2986);
or U7011 (N_7011,N_4267,N_3674);
nor U7012 (N_7012,N_4114,N_2612);
xnor U7013 (N_7013,N_4188,N_4830);
and U7014 (N_7014,N_2949,N_4106);
or U7015 (N_7015,N_3038,N_4924);
nand U7016 (N_7016,N_2928,N_4816);
xor U7017 (N_7017,N_4340,N_3493);
nand U7018 (N_7018,N_4575,N_2714);
or U7019 (N_7019,N_4274,N_3974);
or U7020 (N_7020,N_3995,N_4239);
and U7021 (N_7021,N_4420,N_4809);
xnor U7022 (N_7022,N_2520,N_4550);
and U7023 (N_7023,N_3221,N_3700);
or U7024 (N_7024,N_4665,N_3047);
nor U7025 (N_7025,N_4095,N_3775);
or U7026 (N_7026,N_4336,N_3094);
xnor U7027 (N_7027,N_3987,N_3352);
or U7028 (N_7028,N_3254,N_3286);
and U7029 (N_7029,N_3719,N_4400);
xnor U7030 (N_7030,N_3928,N_4623);
or U7031 (N_7031,N_3656,N_3205);
nor U7032 (N_7032,N_2597,N_4514);
nor U7033 (N_7033,N_4541,N_2717);
nor U7034 (N_7034,N_3910,N_3029);
and U7035 (N_7035,N_4259,N_4812);
and U7036 (N_7036,N_3632,N_4613);
or U7037 (N_7037,N_3987,N_3174);
xnor U7038 (N_7038,N_4946,N_3961);
xnor U7039 (N_7039,N_2615,N_3206);
or U7040 (N_7040,N_3464,N_4809);
and U7041 (N_7041,N_3889,N_2898);
or U7042 (N_7042,N_2785,N_3795);
xor U7043 (N_7043,N_3668,N_4614);
nand U7044 (N_7044,N_3067,N_3531);
nand U7045 (N_7045,N_3322,N_3166);
and U7046 (N_7046,N_4549,N_3820);
and U7047 (N_7047,N_3130,N_3564);
or U7048 (N_7048,N_2652,N_4484);
nand U7049 (N_7049,N_4891,N_4387);
nor U7050 (N_7050,N_4692,N_3478);
nor U7051 (N_7051,N_3870,N_3301);
and U7052 (N_7052,N_4949,N_3147);
nand U7053 (N_7053,N_3992,N_3183);
nand U7054 (N_7054,N_3570,N_2897);
nor U7055 (N_7055,N_3673,N_3687);
nand U7056 (N_7056,N_3859,N_3851);
and U7057 (N_7057,N_4207,N_4092);
xnor U7058 (N_7058,N_4070,N_3352);
or U7059 (N_7059,N_4801,N_3663);
and U7060 (N_7060,N_3744,N_4542);
or U7061 (N_7061,N_2742,N_3940);
and U7062 (N_7062,N_4116,N_3055);
nand U7063 (N_7063,N_2595,N_4597);
xnor U7064 (N_7064,N_4877,N_4876);
and U7065 (N_7065,N_3569,N_3139);
nand U7066 (N_7066,N_3893,N_3832);
xor U7067 (N_7067,N_3495,N_4995);
nand U7068 (N_7068,N_2676,N_3210);
or U7069 (N_7069,N_4530,N_3547);
or U7070 (N_7070,N_3661,N_4481);
and U7071 (N_7071,N_3527,N_4718);
nand U7072 (N_7072,N_3769,N_4003);
xnor U7073 (N_7073,N_3740,N_4421);
or U7074 (N_7074,N_2616,N_3033);
or U7075 (N_7075,N_4739,N_2570);
or U7076 (N_7076,N_4974,N_2770);
nand U7077 (N_7077,N_3671,N_3154);
xor U7078 (N_7078,N_3620,N_4232);
xnor U7079 (N_7079,N_3590,N_3426);
or U7080 (N_7080,N_4094,N_3612);
and U7081 (N_7081,N_3513,N_3185);
nor U7082 (N_7082,N_2883,N_3505);
or U7083 (N_7083,N_3066,N_3777);
and U7084 (N_7084,N_3736,N_3463);
xnor U7085 (N_7085,N_4754,N_4001);
and U7086 (N_7086,N_4164,N_3387);
nor U7087 (N_7087,N_3480,N_3611);
nand U7088 (N_7088,N_4539,N_3265);
nor U7089 (N_7089,N_4355,N_4082);
or U7090 (N_7090,N_3017,N_4496);
xor U7091 (N_7091,N_4502,N_4912);
xnor U7092 (N_7092,N_3365,N_4644);
nor U7093 (N_7093,N_2706,N_2850);
nand U7094 (N_7094,N_3967,N_4517);
or U7095 (N_7095,N_3746,N_3082);
xnor U7096 (N_7096,N_3820,N_4088);
nor U7097 (N_7097,N_2779,N_2548);
nand U7098 (N_7098,N_2892,N_3485);
xnor U7099 (N_7099,N_3168,N_3509);
or U7100 (N_7100,N_4988,N_4894);
and U7101 (N_7101,N_2527,N_2855);
nand U7102 (N_7102,N_3071,N_4818);
xnor U7103 (N_7103,N_4576,N_3105);
xor U7104 (N_7104,N_2845,N_3050);
xnor U7105 (N_7105,N_3299,N_2576);
xor U7106 (N_7106,N_4003,N_3314);
xnor U7107 (N_7107,N_4637,N_4893);
and U7108 (N_7108,N_3994,N_3844);
and U7109 (N_7109,N_3447,N_2933);
or U7110 (N_7110,N_2545,N_3388);
nor U7111 (N_7111,N_4302,N_4925);
and U7112 (N_7112,N_3580,N_4424);
or U7113 (N_7113,N_3662,N_4364);
nand U7114 (N_7114,N_3889,N_4271);
nand U7115 (N_7115,N_4245,N_3803);
and U7116 (N_7116,N_3514,N_2659);
nand U7117 (N_7117,N_4352,N_3115);
xnor U7118 (N_7118,N_4443,N_4194);
nand U7119 (N_7119,N_3544,N_4501);
or U7120 (N_7120,N_4399,N_3642);
and U7121 (N_7121,N_3464,N_4769);
xor U7122 (N_7122,N_4080,N_2858);
or U7123 (N_7123,N_3097,N_3061);
or U7124 (N_7124,N_3175,N_3579);
xnor U7125 (N_7125,N_3041,N_2529);
xnor U7126 (N_7126,N_4172,N_3617);
xor U7127 (N_7127,N_4992,N_2584);
xor U7128 (N_7128,N_2953,N_4377);
nor U7129 (N_7129,N_2571,N_3024);
nor U7130 (N_7130,N_3476,N_4913);
xor U7131 (N_7131,N_3039,N_2997);
nor U7132 (N_7132,N_2513,N_3174);
nor U7133 (N_7133,N_4453,N_4647);
nand U7134 (N_7134,N_3863,N_4458);
or U7135 (N_7135,N_3086,N_2888);
or U7136 (N_7136,N_4811,N_3831);
and U7137 (N_7137,N_3012,N_2720);
xor U7138 (N_7138,N_3799,N_3538);
and U7139 (N_7139,N_3113,N_2570);
nor U7140 (N_7140,N_3796,N_4929);
and U7141 (N_7141,N_3901,N_2873);
and U7142 (N_7142,N_4634,N_2502);
nor U7143 (N_7143,N_4737,N_4653);
xor U7144 (N_7144,N_4598,N_4706);
nor U7145 (N_7145,N_4442,N_3072);
or U7146 (N_7146,N_4781,N_4008);
xor U7147 (N_7147,N_2868,N_4137);
and U7148 (N_7148,N_3870,N_2969);
nand U7149 (N_7149,N_2913,N_2994);
nor U7150 (N_7150,N_3994,N_4718);
xnor U7151 (N_7151,N_4552,N_4398);
or U7152 (N_7152,N_3630,N_2744);
nand U7153 (N_7153,N_4806,N_4816);
nand U7154 (N_7154,N_2965,N_4777);
nand U7155 (N_7155,N_4183,N_4919);
and U7156 (N_7156,N_4958,N_4947);
and U7157 (N_7157,N_3336,N_4928);
or U7158 (N_7158,N_4686,N_3636);
or U7159 (N_7159,N_3310,N_4787);
nand U7160 (N_7160,N_4103,N_2577);
and U7161 (N_7161,N_3010,N_4686);
and U7162 (N_7162,N_4630,N_4423);
nor U7163 (N_7163,N_3739,N_3190);
or U7164 (N_7164,N_4480,N_4499);
xor U7165 (N_7165,N_2654,N_4161);
and U7166 (N_7166,N_3472,N_4036);
and U7167 (N_7167,N_3275,N_2798);
nor U7168 (N_7168,N_3696,N_4815);
and U7169 (N_7169,N_4697,N_4589);
and U7170 (N_7170,N_3495,N_2894);
and U7171 (N_7171,N_2810,N_4795);
xor U7172 (N_7172,N_4588,N_3337);
or U7173 (N_7173,N_3077,N_3708);
nand U7174 (N_7174,N_3270,N_3694);
nand U7175 (N_7175,N_3072,N_4600);
or U7176 (N_7176,N_2842,N_4553);
xor U7177 (N_7177,N_4142,N_4446);
nand U7178 (N_7178,N_3668,N_3774);
nand U7179 (N_7179,N_3381,N_4034);
nor U7180 (N_7180,N_3543,N_3700);
xnor U7181 (N_7181,N_2830,N_3180);
and U7182 (N_7182,N_4325,N_3642);
nor U7183 (N_7183,N_3773,N_3260);
and U7184 (N_7184,N_2769,N_3976);
xor U7185 (N_7185,N_3940,N_4890);
and U7186 (N_7186,N_2958,N_3096);
xnor U7187 (N_7187,N_4384,N_3023);
nand U7188 (N_7188,N_4668,N_3430);
xnor U7189 (N_7189,N_3088,N_2620);
nor U7190 (N_7190,N_3345,N_3103);
and U7191 (N_7191,N_3809,N_4546);
and U7192 (N_7192,N_2587,N_4003);
nand U7193 (N_7193,N_4599,N_2974);
xor U7194 (N_7194,N_3982,N_4948);
xor U7195 (N_7195,N_4694,N_4760);
nor U7196 (N_7196,N_4046,N_4011);
or U7197 (N_7197,N_3631,N_3889);
xnor U7198 (N_7198,N_3927,N_3047);
and U7199 (N_7199,N_3334,N_3430);
and U7200 (N_7200,N_4589,N_3351);
nor U7201 (N_7201,N_4370,N_4899);
xnor U7202 (N_7202,N_3477,N_4715);
or U7203 (N_7203,N_3211,N_3846);
xnor U7204 (N_7204,N_3156,N_3944);
or U7205 (N_7205,N_3334,N_3067);
or U7206 (N_7206,N_4735,N_4974);
and U7207 (N_7207,N_4608,N_3391);
nor U7208 (N_7208,N_3921,N_3471);
xnor U7209 (N_7209,N_3061,N_4226);
and U7210 (N_7210,N_3829,N_3820);
nor U7211 (N_7211,N_3062,N_4886);
xnor U7212 (N_7212,N_2632,N_4758);
nor U7213 (N_7213,N_2714,N_3114);
and U7214 (N_7214,N_4273,N_2927);
nor U7215 (N_7215,N_3108,N_2648);
or U7216 (N_7216,N_2612,N_4753);
nand U7217 (N_7217,N_3138,N_3452);
or U7218 (N_7218,N_4290,N_4586);
nand U7219 (N_7219,N_3243,N_3298);
nor U7220 (N_7220,N_3837,N_4579);
xor U7221 (N_7221,N_3336,N_2552);
nor U7222 (N_7222,N_4475,N_4127);
nand U7223 (N_7223,N_4072,N_3066);
nand U7224 (N_7224,N_4540,N_3798);
nand U7225 (N_7225,N_2765,N_3787);
nand U7226 (N_7226,N_4238,N_4653);
nand U7227 (N_7227,N_2746,N_4378);
nor U7228 (N_7228,N_3811,N_2604);
xnor U7229 (N_7229,N_2973,N_3580);
nor U7230 (N_7230,N_3698,N_4811);
nor U7231 (N_7231,N_3713,N_4411);
nor U7232 (N_7232,N_3682,N_2983);
nand U7233 (N_7233,N_3773,N_3790);
and U7234 (N_7234,N_3578,N_4445);
xnor U7235 (N_7235,N_2766,N_4438);
or U7236 (N_7236,N_4410,N_3871);
nor U7237 (N_7237,N_3120,N_4059);
or U7238 (N_7238,N_3652,N_3884);
and U7239 (N_7239,N_2711,N_4822);
or U7240 (N_7240,N_4848,N_3818);
nor U7241 (N_7241,N_4991,N_3407);
nand U7242 (N_7242,N_4660,N_3581);
nor U7243 (N_7243,N_3932,N_3696);
nand U7244 (N_7244,N_4348,N_3751);
or U7245 (N_7245,N_2959,N_2663);
nor U7246 (N_7246,N_3963,N_3536);
nand U7247 (N_7247,N_3349,N_2865);
or U7248 (N_7248,N_3916,N_2646);
nand U7249 (N_7249,N_3245,N_4049);
and U7250 (N_7250,N_4896,N_4237);
and U7251 (N_7251,N_3838,N_4102);
xor U7252 (N_7252,N_4696,N_4959);
nor U7253 (N_7253,N_3438,N_4436);
nand U7254 (N_7254,N_4663,N_3846);
or U7255 (N_7255,N_4981,N_3362);
xnor U7256 (N_7256,N_2527,N_3086);
nor U7257 (N_7257,N_4585,N_3819);
nand U7258 (N_7258,N_3899,N_2574);
or U7259 (N_7259,N_2897,N_3995);
nor U7260 (N_7260,N_3025,N_3474);
nand U7261 (N_7261,N_4857,N_4804);
nand U7262 (N_7262,N_2729,N_4105);
nor U7263 (N_7263,N_4103,N_2838);
or U7264 (N_7264,N_3949,N_4846);
xor U7265 (N_7265,N_4894,N_4842);
or U7266 (N_7266,N_3592,N_2610);
xor U7267 (N_7267,N_4392,N_4931);
or U7268 (N_7268,N_3078,N_4926);
or U7269 (N_7269,N_2959,N_4197);
nand U7270 (N_7270,N_4827,N_4072);
nor U7271 (N_7271,N_2724,N_4380);
xor U7272 (N_7272,N_3663,N_4392);
xor U7273 (N_7273,N_3026,N_4534);
nor U7274 (N_7274,N_4488,N_3442);
nand U7275 (N_7275,N_3502,N_2540);
and U7276 (N_7276,N_4709,N_4707);
nand U7277 (N_7277,N_3842,N_3149);
xnor U7278 (N_7278,N_4028,N_4751);
or U7279 (N_7279,N_2908,N_3602);
or U7280 (N_7280,N_4764,N_2971);
xnor U7281 (N_7281,N_2554,N_2547);
xnor U7282 (N_7282,N_3029,N_2707);
or U7283 (N_7283,N_2939,N_4592);
nand U7284 (N_7284,N_4761,N_3370);
xnor U7285 (N_7285,N_4938,N_3939);
and U7286 (N_7286,N_4916,N_3009);
and U7287 (N_7287,N_4946,N_4657);
and U7288 (N_7288,N_4876,N_3051);
xnor U7289 (N_7289,N_2682,N_4121);
or U7290 (N_7290,N_3211,N_3347);
xor U7291 (N_7291,N_2908,N_3660);
or U7292 (N_7292,N_2815,N_2637);
nor U7293 (N_7293,N_4738,N_3971);
nand U7294 (N_7294,N_3794,N_3289);
nor U7295 (N_7295,N_4563,N_3818);
nor U7296 (N_7296,N_4978,N_3805);
nor U7297 (N_7297,N_2649,N_4701);
nor U7298 (N_7298,N_4032,N_4743);
or U7299 (N_7299,N_3872,N_4194);
or U7300 (N_7300,N_3228,N_3987);
nor U7301 (N_7301,N_2999,N_4780);
or U7302 (N_7302,N_3025,N_4416);
or U7303 (N_7303,N_4985,N_2773);
nor U7304 (N_7304,N_2880,N_3524);
xnor U7305 (N_7305,N_3815,N_4605);
nand U7306 (N_7306,N_3687,N_2970);
and U7307 (N_7307,N_4512,N_4020);
nor U7308 (N_7308,N_4428,N_2799);
or U7309 (N_7309,N_2513,N_3955);
or U7310 (N_7310,N_3396,N_4590);
nor U7311 (N_7311,N_4166,N_4974);
nand U7312 (N_7312,N_4894,N_4965);
and U7313 (N_7313,N_4546,N_4160);
nand U7314 (N_7314,N_3480,N_4214);
nand U7315 (N_7315,N_3753,N_4026);
xor U7316 (N_7316,N_3084,N_2860);
and U7317 (N_7317,N_3388,N_4231);
or U7318 (N_7318,N_3006,N_4829);
and U7319 (N_7319,N_2948,N_2743);
xor U7320 (N_7320,N_2674,N_4854);
xnor U7321 (N_7321,N_4889,N_2807);
or U7322 (N_7322,N_4714,N_3183);
or U7323 (N_7323,N_4308,N_4935);
xnor U7324 (N_7324,N_2932,N_4287);
or U7325 (N_7325,N_3233,N_3345);
nor U7326 (N_7326,N_4874,N_3824);
xnor U7327 (N_7327,N_2624,N_3507);
xor U7328 (N_7328,N_3857,N_3574);
xnor U7329 (N_7329,N_2865,N_4598);
or U7330 (N_7330,N_3244,N_2909);
and U7331 (N_7331,N_3574,N_4813);
nand U7332 (N_7332,N_3802,N_4479);
or U7333 (N_7333,N_4412,N_4638);
xnor U7334 (N_7334,N_3643,N_3095);
and U7335 (N_7335,N_4017,N_3949);
or U7336 (N_7336,N_3205,N_3385);
xnor U7337 (N_7337,N_4225,N_3558);
or U7338 (N_7338,N_4655,N_3862);
or U7339 (N_7339,N_3741,N_2798);
nand U7340 (N_7340,N_4149,N_3763);
and U7341 (N_7341,N_3833,N_3931);
xnor U7342 (N_7342,N_4510,N_4287);
xor U7343 (N_7343,N_4688,N_2500);
and U7344 (N_7344,N_3348,N_4688);
or U7345 (N_7345,N_4856,N_4366);
and U7346 (N_7346,N_2609,N_2530);
nor U7347 (N_7347,N_3438,N_3560);
xnor U7348 (N_7348,N_4103,N_4437);
nand U7349 (N_7349,N_2563,N_2660);
or U7350 (N_7350,N_2971,N_4975);
or U7351 (N_7351,N_3601,N_4984);
nor U7352 (N_7352,N_2950,N_3453);
and U7353 (N_7353,N_3293,N_4261);
and U7354 (N_7354,N_4137,N_4623);
or U7355 (N_7355,N_3565,N_4750);
and U7356 (N_7356,N_2727,N_4334);
or U7357 (N_7357,N_2768,N_2871);
nand U7358 (N_7358,N_3822,N_4359);
or U7359 (N_7359,N_4861,N_3400);
and U7360 (N_7360,N_2713,N_3578);
nor U7361 (N_7361,N_2792,N_3746);
xnor U7362 (N_7362,N_3224,N_4849);
nand U7363 (N_7363,N_4112,N_4004);
and U7364 (N_7364,N_3453,N_3955);
and U7365 (N_7365,N_3305,N_4822);
xnor U7366 (N_7366,N_3682,N_3292);
nor U7367 (N_7367,N_2505,N_2570);
or U7368 (N_7368,N_4403,N_4840);
xnor U7369 (N_7369,N_3863,N_2839);
nor U7370 (N_7370,N_2930,N_2663);
nor U7371 (N_7371,N_4569,N_2509);
nand U7372 (N_7372,N_3947,N_4121);
or U7373 (N_7373,N_4551,N_4818);
and U7374 (N_7374,N_3032,N_4823);
and U7375 (N_7375,N_3092,N_3550);
or U7376 (N_7376,N_2870,N_3424);
or U7377 (N_7377,N_2578,N_3405);
and U7378 (N_7378,N_3344,N_4928);
nand U7379 (N_7379,N_4138,N_4203);
and U7380 (N_7380,N_4895,N_4684);
nor U7381 (N_7381,N_4217,N_2565);
or U7382 (N_7382,N_3823,N_4649);
or U7383 (N_7383,N_3840,N_4531);
xnor U7384 (N_7384,N_4635,N_4221);
and U7385 (N_7385,N_3471,N_3852);
nand U7386 (N_7386,N_3024,N_4535);
xor U7387 (N_7387,N_4987,N_4389);
nand U7388 (N_7388,N_3931,N_3706);
nand U7389 (N_7389,N_4114,N_3484);
and U7390 (N_7390,N_2997,N_3197);
nand U7391 (N_7391,N_3234,N_3086);
nor U7392 (N_7392,N_3781,N_4189);
nand U7393 (N_7393,N_4481,N_4204);
xor U7394 (N_7394,N_3583,N_2602);
xor U7395 (N_7395,N_3544,N_3789);
and U7396 (N_7396,N_3261,N_4271);
or U7397 (N_7397,N_2895,N_3731);
xnor U7398 (N_7398,N_4477,N_3477);
or U7399 (N_7399,N_3658,N_2603);
and U7400 (N_7400,N_2852,N_3339);
and U7401 (N_7401,N_2586,N_3991);
and U7402 (N_7402,N_4327,N_4022);
nand U7403 (N_7403,N_4177,N_3298);
nor U7404 (N_7404,N_4291,N_2723);
nor U7405 (N_7405,N_4640,N_3379);
nand U7406 (N_7406,N_2890,N_3087);
xnor U7407 (N_7407,N_3420,N_4411);
nand U7408 (N_7408,N_4609,N_3526);
or U7409 (N_7409,N_3673,N_2872);
xor U7410 (N_7410,N_3063,N_3301);
and U7411 (N_7411,N_4393,N_3541);
and U7412 (N_7412,N_4416,N_3426);
nand U7413 (N_7413,N_3215,N_3846);
xor U7414 (N_7414,N_4582,N_4938);
nor U7415 (N_7415,N_3034,N_4006);
or U7416 (N_7416,N_3347,N_4211);
xor U7417 (N_7417,N_3748,N_4461);
and U7418 (N_7418,N_3735,N_4510);
xnor U7419 (N_7419,N_4378,N_3447);
and U7420 (N_7420,N_4383,N_4424);
nor U7421 (N_7421,N_3367,N_3090);
or U7422 (N_7422,N_4641,N_2572);
nor U7423 (N_7423,N_3785,N_3334);
and U7424 (N_7424,N_4071,N_3316);
nor U7425 (N_7425,N_3327,N_3445);
or U7426 (N_7426,N_2611,N_4038);
or U7427 (N_7427,N_4787,N_4674);
nand U7428 (N_7428,N_4281,N_4108);
or U7429 (N_7429,N_4858,N_2813);
xnor U7430 (N_7430,N_4570,N_4330);
or U7431 (N_7431,N_4975,N_3609);
nor U7432 (N_7432,N_2847,N_4476);
nor U7433 (N_7433,N_3551,N_3553);
nor U7434 (N_7434,N_4722,N_3769);
nor U7435 (N_7435,N_3157,N_2643);
xnor U7436 (N_7436,N_3327,N_4606);
or U7437 (N_7437,N_2966,N_3461);
nor U7438 (N_7438,N_4140,N_4295);
and U7439 (N_7439,N_4442,N_3798);
and U7440 (N_7440,N_3720,N_4090);
nand U7441 (N_7441,N_2922,N_3084);
nand U7442 (N_7442,N_2942,N_4638);
or U7443 (N_7443,N_4519,N_3003);
xor U7444 (N_7444,N_3031,N_4763);
and U7445 (N_7445,N_4102,N_4991);
nand U7446 (N_7446,N_4977,N_4094);
and U7447 (N_7447,N_3527,N_3931);
nand U7448 (N_7448,N_4718,N_3946);
or U7449 (N_7449,N_4200,N_3705);
xnor U7450 (N_7450,N_4881,N_4992);
xor U7451 (N_7451,N_3107,N_3688);
nor U7452 (N_7452,N_4998,N_2868);
and U7453 (N_7453,N_2944,N_4440);
nand U7454 (N_7454,N_3384,N_3033);
nor U7455 (N_7455,N_4243,N_3695);
xnor U7456 (N_7456,N_3609,N_3133);
xor U7457 (N_7457,N_3350,N_2890);
or U7458 (N_7458,N_3607,N_3711);
nor U7459 (N_7459,N_4213,N_3836);
or U7460 (N_7460,N_2507,N_2891);
nand U7461 (N_7461,N_3164,N_2715);
nand U7462 (N_7462,N_4218,N_2902);
nor U7463 (N_7463,N_2818,N_3512);
and U7464 (N_7464,N_4670,N_4972);
nor U7465 (N_7465,N_3987,N_4950);
nand U7466 (N_7466,N_4615,N_2660);
nor U7467 (N_7467,N_2888,N_4552);
nor U7468 (N_7468,N_4491,N_2833);
or U7469 (N_7469,N_3451,N_2656);
and U7470 (N_7470,N_4333,N_4886);
nand U7471 (N_7471,N_3283,N_4608);
and U7472 (N_7472,N_4465,N_4637);
nor U7473 (N_7473,N_3039,N_3680);
or U7474 (N_7474,N_3950,N_3605);
or U7475 (N_7475,N_3016,N_4480);
or U7476 (N_7476,N_3038,N_4586);
xor U7477 (N_7477,N_4861,N_3797);
or U7478 (N_7478,N_4651,N_4804);
or U7479 (N_7479,N_4710,N_3738);
nor U7480 (N_7480,N_3289,N_3775);
nand U7481 (N_7481,N_4384,N_2755);
xor U7482 (N_7482,N_2876,N_3677);
and U7483 (N_7483,N_3447,N_4227);
xor U7484 (N_7484,N_2880,N_3067);
nor U7485 (N_7485,N_4846,N_2986);
nand U7486 (N_7486,N_4805,N_3074);
nand U7487 (N_7487,N_3419,N_4534);
xnor U7488 (N_7488,N_4196,N_3194);
or U7489 (N_7489,N_3772,N_4797);
xnor U7490 (N_7490,N_3381,N_4351);
and U7491 (N_7491,N_4619,N_3228);
nor U7492 (N_7492,N_3310,N_3510);
xor U7493 (N_7493,N_3212,N_4085);
and U7494 (N_7494,N_4071,N_4348);
or U7495 (N_7495,N_3411,N_2680);
and U7496 (N_7496,N_4441,N_2514);
or U7497 (N_7497,N_3299,N_3823);
nor U7498 (N_7498,N_2580,N_4614);
nor U7499 (N_7499,N_4932,N_4943);
xnor U7500 (N_7500,N_5460,N_7469);
and U7501 (N_7501,N_6760,N_7242);
and U7502 (N_7502,N_6906,N_5500);
or U7503 (N_7503,N_7028,N_7002);
nand U7504 (N_7504,N_6502,N_5731);
xor U7505 (N_7505,N_6320,N_7425);
xor U7506 (N_7506,N_5171,N_7300);
or U7507 (N_7507,N_7333,N_5117);
xnor U7508 (N_7508,N_7004,N_5102);
or U7509 (N_7509,N_6232,N_7016);
nor U7510 (N_7510,N_5188,N_5626);
nand U7511 (N_7511,N_6148,N_6490);
xor U7512 (N_7512,N_6503,N_5431);
or U7513 (N_7513,N_6084,N_5657);
xor U7514 (N_7514,N_6060,N_6671);
xor U7515 (N_7515,N_5800,N_7225);
or U7516 (N_7516,N_7387,N_5282);
xnor U7517 (N_7517,N_6007,N_5200);
and U7518 (N_7518,N_5549,N_6939);
and U7519 (N_7519,N_6241,N_5374);
and U7520 (N_7520,N_6545,N_7116);
or U7521 (N_7521,N_7495,N_6116);
nor U7522 (N_7522,N_6147,N_6220);
or U7523 (N_7523,N_5107,N_6223);
nand U7524 (N_7524,N_5133,N_6643);
nor U7525 (N_7525,N_6819,N_7172);
nand U7526 (N_7526,N_5695,N_6588);
and U7527 (N_7527,N_5059,N_5675);
xor U7528 (N_7528,N_5994,N_6036);
or U7529 (N_7529,N_5013,N_6401);
and U7530 (N_7530,N_5357,N_5017);
nand U7531 (N_7531,N_6156,N_6962);
or U7532 (N_7532,N_6552,N_6211);
nor U7533 (N_7533,N_6488,N_5104);
or U7534 (N_7534,N_5796,N_5077);
nand U7535 (N_7535,N_5398,N_7201);
nor U7536 (N_7536,N_6646,N_6308);
nand U7537 (N_7537,N_6780,N_6064);
and U7538 (N_7538,N_5339,N_5973);
or U7539 (N_7539,N_5176,N_6542);
nor U7540 (N_7540,N_7184,N_6628);
xor U7541 (N_7541,N_5049,N_5518);
xor U7542 (N_7542,N_6208,N_5365);
and U7543 (N_7543,N_5141,N_6394);
nor U7544 (N_7544,N_6594,N_7293);
nand U7545 (N_7545,N_7091,N_6432);
nor U7546 (N_7546,N_7388,N_5445);
xnor U7547 (N_7547,N_5429,N_6992);
and U7548 (N_7548,N_7243,N_7200);
or U7549 (N_7549,N_7284,N_5438);
or U7550 (N_7550,N_5498,N_6586);
and U7551 (N_7551,N_6321,N_5856);
nand U7552 (N_7552,N_5301,N_6080);
or U7553 (N_7553,N_6100,N_5385);
nand U7554 (N_7554,N_6904,N_5825);
xnor U7555 (N_7555,N_5725,N_6551);
or U7556 (N_7556,N_5435,N_6338);
nand U7557 (N_7557,N_7251,N_7268);
xnor U7558 (N_7558,N_6374,N_6250);
nand U7559 (N_7559,N_5162,N_6442);
nor U7560 (N_7560,N_5192,N_7176);
xnor U7561 (N_7561,N_6027,N_5560);
or U7562 (N_7562,N_5862,N_7338);
or U7563 (N_7563,N_7072,N_6290);
or U7564 (N_7564,N_6342,N_5978);
nand U7565 (N_7565,N_6969,N_6294);
or U7566 (N_7566,N_6896,N_5260);
nor U7567 (N_7567,N_5961,N_5410);
nor U7568 (N_7568,N_6828,N_5934);
nor U7569 (N_7569,N_5362,N_6443);
nand U7570 (N_7570,N_7205,N_5240);
or U7571 (N_7571,N_6960,N_5408);
and U7572 (N_7572,N_6304,N_5003);
and U7573 (N_7573,N_7000,N_6310);
nor U7574 (N_7574,N_7427,N_6203);
or U7575 (N_7575,N_5783,N_5343);
nand U7576 (N_7576,N_5330,N_6331);
and U7577 (N_7577,N_5633,N_5294);
nand U7578 (N_7578,N_5517,N_7165);
and U7579 (N_7579,N_5782,N_5131);
and U7580 (N_7580,N_6804,N_6648);
nor U7581 (N_7581,N_6987,N_6596);
nand U7582 (N_7582,N_6165,N_5291);
nor U7583 (N_7583,N_6664,N_6576);
or U7584 (N_7584,N_5839,N_5119);
or U7585 (N_7585,N_6172,N_5000);
xnor U7586 (N_7586,N_7210,N_7109);
xnor U7587 (N_7587,N_6766,N_6273);
or U7588 (N_7588,N_6425,N_5273);
and U7589 (N_7589,N_6974,N_6091);
and U7590 (N_7590,N_6189,N_7066);
nand U7591 (N_7591,N_7032,N_5110);
nand U7592 (N_7592,N_5641,N_7168);
xnor U7593 (N_7593,N_7438,N_5457);
xnor U7594 (N_7594,N_7418,N_6621);
xor U7595 (N_7595,N_5718,N_6427);
nand U7596 (N_7596,N_6641,N_6805);
and U7597 (N_7597,N_5160,N_6219);
nand U7598 (N_7598,N_6402,N_7270);
nand U7599 (N_7599,N_5363,N_6185);
xnor U7600 (N_7600,N_5703,N_7453);
nor U7601 (N_7601,N_6270,N_6692);
and U7602 (N_7602,N_5661,N_5381);
xor U7603 (N_7603,N_7164,N_6434);
nor U7604 (N_7604,N_7173,N_5074);
or U7605 (N_7605,N_7157,N_6650);
xor U7606 (N_7606,N_6891,N_7351);
xor U7607 (N_7607,N_7045,N_5719);
nor U7608 (N_7608,N_5653,N_5752);
xor U7609 (N_7609,N_5341,N_6476);
or U7610 (N_7610,N_6030,N_6920);
nand U7611 (N_7611,N_5004,N_7189);
nand U7612 (N_7612,N_5267,N_5544);
xnor U7613 (N_7613,N_6843,N_6979);
nand U7614 (N_7614,N_7101,N_7250);
or U7615 (N_7615,N_7148,N_5832);
or U7616 (N_7616,N_6395,N_5726);
nand U7617 (N_7617,N_7328,N_5737);
and U7618 (N_7618,N_6753,N_6759);
xor U7619 (N_7619,N_5925,N_5182);
nand U7620 (N_7620,N_7127,N_6140);
nor U7621 (N_7621,N_6360,N_7070);
nand U7622 (N_7622,N_5336,N_7337);
and U7623 (N_7623,N_7299,N_5519);
nor U7624 (N_7624,N_5993,N_6302);
and U7625 (N_7625,N_6940,N_7140);
nand U7626 (N_7626,N_7391,N_6106);
nor U7627 (N_7627,N_5103,N_5067);
or U7628 (N_7628,N_7206,N_6396);
and U7629 (N_7629,N_6644,N_6584);
nor U7630 (N_7630,N_7353,N_5366);
xor U7631 (N_7631,N_5837,N_5411);
and U7632 (N_7632,N_6484,N_5802);
xnor U7633 (N_7633,N_7138,N_7443);
nand U7634 (N_7634,N_6371,N_5161);
xnor U7635 (N_7635,N_6066,N_5210);
or U7636 (N_7636,N_5450,N_5114);
xor U7637 (N_7637,N_5801,N_6417);
nand U7638 (N_7638,N_5533,N_5577);
nand U7639 (N_7639,N_5579,N_5252);
nand U7640 (N_7640,N_5520,N_6405);
xnor U7641 (N_7641,N_7130,N_5685);
nor U7642 (N_7642,N_6052,N_6235);
nor U7643 (N_7643,N_5478,N_6566);
nor U7644 (N_7644,N_5100,N_6034);
and U7645 (N_7645,N_5525,N_5673);
and U7646 (N_7646,N_6251,N_7497);
and U7647 (N_7647,N_7113,N_5574);
xor U7648 (N_7648,N_5591,N_6433);
nand U7649 (N_7649,N_6178,N_6240);
or U7650 (N_7650,N_7098,N_6000);
nand U7651 (N_7651,N_6244,N_6101);
xor U7652 (N_7652,N_6806,N_6718);
xor U7653 (N_7653,N_6212,N_7074);
or U7654 (N_7654,N_6218,N_6154);
nor U7655 (N_7655,N_6568,N_6480);
or U7656 (N_7656,N_6821,N_5654);
xor U7657 (N_7657,N_6949,N_7218);
and U7658 (N_7658,N_6537,N_5687);
or U7659 (N_7659,N_6726,N_5486);
or U7660 (N_7660,N_5937,N_6793);
and U7661 (N_7661,N_5553,N_5600);
nand U7662 (N_7662,N_5557,N_6337);
or U7663 (N_7663,N_7481,N_5268);
nand U7664 (N_7664,N_6961,N_5762);
or U7665 (N_7665,N_7463,N_6051);
nand U7666 (N_7666,N_5543,N_7194);
and U7667 (N_7667,N_6067,N_7363);
xor U7668 (N_7668,N_6851,N_5281);
or U7669 (N_7669,N_6550,N_5694);
nand U7670 (N_7670,N_6216,N_5873);
or U7671 (N_7671,N_7022,N_5901);
xnor U7672 (N_7672,N_7137,N_7464);
xnor U7673 (N_7673,N_5037,N_6840);
nor U7674 (N_7674,N_5691,N_7457);
xnor U7675 (N_7675,N_5639,N_7343);
or U7676 (N_7676,N_6820,N_7383);
and U7677 (N_7677,N_5382,N_7372);
nand U7678 (N_7678,N_7232,N_5417);
xor U7679 (N_7679,N_6543,N_7245);
nor U7680 (N_7680,N_7327,N_7001);
nor U7681 (N_7681,N_6248,N_5091);
xnor U7682 (N_7682,N_5640,N_5045);
and U7683 (N_7683,N_6177,N_5667);
or U7684 (N_7684,N_6951,N_5052);
or U7685 (N_7685,N_5092,N_5872);
xnor U7686 (N_7686,N_5088,N_5256);
and U7687 (N_7687,N_5581,N_7269);
nand U7688 (N_7688,N_7038,N_6050);
or U7689 (N_7689,N_6298,N_7491);
xor U7690 (N_7690,N_6553,N_6815);
and U7691 (N_7691,N_5396,N_5170);
xnor U7692 (N_7692,N_6312,N_5356);
nor U7693 (N_7693,N_5936,N_7399);
xor U7694 (N_7694,N_7365,N_6869);
nand U7695 (N_7695,N_7234,N_7472);
or U7696 (N_7696,N_6514,N_6998);
nand U7697 (N_7697,N_6778,N_6271);
nand U7698 (N_7698,N_6303,N_5916);
nand U7699 (N_7699,N_6547,N_6860);
nand U7700 (N_7700,N_6075,N_6842);
and U7701 (N_7701,N_5881,N_5477);
or U7702 (N_7702,N_5875,N_6506);
or U7703 (N_7703,N_6015,N_6365);
xnor U7704 (N_7704,N_7429,N_7092);
and U7705 (N_7705,N_6830,N_5361);
nor U7706 (N_7706,N_5242,N_6682);
xor U7707 (N_7707,N_7492,N_6744);
nor U7708 (N_7708,N_7371,N_5137);
nor U7709 (N_7709,N_6014,N_6288);
or U7710 (N_7710,N_6202,N_5124);
and U7711 (N_7711,N_5423,N_5788);
nor U7712 (N_7712,N_5157,N_6436);
and U7713 (N_7713,N_7292,N_5266);
nor U7714 (N_7714,N_5746,N_7442);
or U7715 (N_7715,N_5727,N_6237);
nor U7716 (N_7716,N_5205,N_5546);
xnor U7717 (N_7717,N_5809,N_6572);
or U7718 (N_7718,N_7424,N_6756);
nand U7719 (N_7719,N_5563,N_5007);
and U7720 (N_7720,N_6149,N_6755);
nand U7721 (N_7721,N_5020,N_5305);
and U7722 (N_7722,N_6781,N_5771);
nor U7723 (N_7723,N_6006,N_7440);
nor U7724 (N_7724,N_7095,N_7008);
nand U7725 (N_7725,N_5204,N_5975);
or U7726 (N_7726,N_5008,N_6640);
or U7727 (N_7727,N_7480,N_7123);
nand U7728 (N_7728,N_5774,N_6309);
xor U7729 (N_7729,N_5097,N_6113);
or U7730 (N_7730,N_5548,N_7026);
xnor U7731 (N_7731,N_5314,N_5140);
xnor U7732 (N_7732,N_6608,N_7386);
xor U7733 (N_7733,N_7256,N_6965);
nor U7734 (N_7734,N_6261,N_6582);
nand U7735 (N_7735,N_5526,N_5624);
nor U7736 (N_7736,N_5216,N_7308);
nand U7737 (N_7737,N_5354,N_7125);
xor U7738 (N_7738,N_7190,N_6257);
or U7739 (N_7739,N_6012,N_7483);
nand U7740 (N_7740,N_6859,N_6844);
nor U7741 (N_7741,N_5985,N_7192);
and U7742 (N_7742,N_5813,N_5159);
nand U7743 (N_7743,N_6131,N_7393);
and U7744 (N_7744,N_5995,N_7494);
or U7745 (N_7745,N_6872,N_6201);
xnor U7746 (N_7746,N_6354,N_5912);
nand U7747 (N_7747,N_5595,N_7407);
nand U7748 (N_7748,N_6526,N_5803);
xor U7749 (N_7749,N_5387,N_6653);
and U7750 (N_7750,N_7482,N_7454);
nor U7751 (N_7751,N_7163,N_5467);
nor U7752 (N_7752,N_5741,N_7275);
xnor U7753 (N_7753,N_5482,N_5288);
nand U7754 (N_7754,N_5617,N_6814);
nand U7755 (N_7755,N_5014,N_7410);
nor U7756 (N_7756,N_6573,N_7191);
or U7757 (N_7757,N_6004,N_5596);
and U7758 (N_7758,N_7277,N_6236);
nor U7759 (N_7759,N_6347,N_6512);
nand U7760 (N_7760,N_6757,N_7342);
xnor U7761 (N_7761,N_6112,N_5938);
xor U7762 (N_7762,N_6262,N_6867);
xor U7763 (N_7763,N_5243,N_6481);
or U7764 (N_7764,N_5605,N_5223);
nand U7765 (N_7765,N_5906,N_5972);
xnor U7766 (N_7766,N_5736,N_7226);
nor U7767 (N_7767,N_5849,N_6467);
xnor U7768 (N_7768,N_6746,N_5487);
nand U7769 (N_7769,N_6922,N_7392);
or U7770 (N_7770,N_5735,N_6192);
or U7771 (N_7771,N_5218,N_6794);
or U7772 (N_7772,N_7015,N_5147);
nor U7773 (N_7773,N_5742,N_7291);
nor U7774 (N_7774,N_6964,N_6912);
nand U7775 (N_7775,N_5129,N_5241);
and U7776 (N_7776,N_7063,N_5384);
or U7777 (N_7777,N_6109,N_6021);
and U7778 (N_7778,N_6372,N_6721);
nor U7779 (N_7779,N_7025,N_5466);
xnor U7780 (N_7780,N_7334,N_5461);
xor U7781 (N_7781,N_5247,N_5175);
or U7782 (N_7782,N_6130,N_5528);
and U7783 (N_7783,N_6611,N_6703);
or U7784 (N_7784,N_6665,N_5127);
nor U7785 (N_7785,N_5493,N_6779);
xor U7786 (N_7786,N_5503,N_7068);
nand U7787 (N_7787,N_6833,N_5649);
nand U7788 (N_7788,N_7118,N_6413);
and U7789 (N_7789,N_6120,N_6351);
nand U7790 (N_7790,N_6022,N_6194);
xnor U7791 (N_7791,N_5132,N_7126);
nand U7792 (N_7792,N_5815,N_7255);
and U7793 (N_7793,N_6631,N_5660);
or U7794 (N_7794,N_5767,N_5785);
or U7795 (N_7795,N_5619,N_6018);
and U7796 (N_7796,N_7145,N_6745);
xor U7797 (N_7797,N_6437,N_5562);
nand U7798 (N_7798,N_7428,N_5709);
and U7799 (N_7799,N_5510,N_6375);
and U7800 (N_7800,N_7107,N_6911);
or U7801 (N_7801,N_7366,N_5778);
nor U7802 (N_7802,N_6296,N_6564);
or U7803 (N_7803,N_7433,N_6069);
or U7804 (N_7804,N_7448,N_6187);
or U7805 (N_7805,N_5250,N_6930);
nor U7806 (N_7806,N_5035,N_6901);
xnor U7807 (N_7807,N_6412,N_6186);
nor U7808 (N_7808,N_5075,N_6724);
xnor U7809 (N_7809,N_6485,N_5748);
and U7810 (N_7810,N_5342,N_7005);
and U7811 (N_7811,N_6300,N_6556);
or U7812 (N_7812,N_5958,N_6517);
xnor U7813 (N_7813,N_5884,N_5733);
or U7814 (N_7814,N_5468,N_6945);
nor U7815 (N_7815,N_5113,N_5949);
nor U7816 (N_7816,N_6438,N_5062);
and U7817 (N_7817,N_6111,N_7430);
nand U7818 (N_7818,N_7304,N_6875);
or U7819 (N_7819,N_6801,N_7043);
or U7820 (N_7820,N_6649,N_5126);
xor U7821 (N_7821,N_5812,N_6970);
or U7822 (N_7822,N_5854,N_6093);
and U7823 (N_7823,N_7082,N_5959);
xor U7824 (N_7824,N_6157,N_5195);
nand U7825 (N_7825,N_5980,N_6175);
nand U7826 (N_7826,N_5261,N_5723);
nand U7827 (N_7827,N_5564,N_6155);
xor U7828 (N_7828,N_5257,N_6426);
nor U7829 (N_7829,N_6439,N_7394);
nor U7830 (N_7830,N_5756,N_6441);
and U7831 (N_7831,N_6733,N_6910);
nand U7832 (N_7832,N_6670,N_6297);
nor U7833 (N_7833,N_6368,N_7489);
nor U7834 (N_7834,N_6180,N_6095);
nand U7835 (N_7835,N_5939,N_6919);
nor U7836 (N_7836,N_5621,N_6638);
nand U7837 (N_7837,N_5300,N_6902);
xor U7838 (N_7838,N_5966,N_6651);
xor U7839 (N_7839,N_5632,N_5513);
and U7840 (N_7840,N_7094,N_6104);
or U7841 (N_7841,N_6316,N_6719);
nand U7842 (N_7842,N_6404,N_7061);
nor U7843 (N_7843,N_6062,N_7437);
nand U7844 (N_7844,N_7326,N_6834);
xor U7845 (N_7845,N_5227,N_6619);
nand U7846 (N_7846,N_5848,N_6739);
or U7847 (N_7847,N_6010,N_6336);
and U7848 (N_7848,N_5146,N_7170);
nor U7849 (N_7849,N_5860,N_6415);
or U7850 (N_7850,N_5514,N_7247);
or U7851 (N_7851,N_7104,N_5747);
and U7852 (N_7852,N_5616,N_6934);
nor U7853 (N_7853,N_6943,N_6418);
and U7854 (N_7854,N_7455,N_6306);
nor U7855 (N_7855,N_5547,N_7236);
xnor U7856 (N_7856,N_5618,N_5597);
or U7857 (N_7857,N_5473,N_6457);
or U7858 (N_7858,N_5427,N_6046);
nand U7859 (N_7859,N_5350,N_5297);
or U7860 (N_7860,N_5886,N_5692);
and U7861 (N_7861,N_7133,N_5263);
nor U7862 (N_7862,N_6174,N_5941);
nand U7863 (N_7863,N_7035,N_5515);
xor U7864 (N_7864,N_5507,N_6164);
and U7865 (N_7865,N_5644,N_7354);
nor U7866 (N_7866,N_6121,N_6520);
xor U7867 (N_7867,N_5932,N_7271);
nand U7868 (N_7868,N_6725,N_7166);
xnor U7869 (N_7869,N_6575,N_5948);
nor U7870 (N_7870,N_7389,N_6055);
or U7871 (N_7871,N_7196,N_7136);
or U7872 (N_7872,N_7128,N_6836);
and U7873 (N_7873,N_6269,N_6074);
nor U7874 (N_7874,N_5522,N_6039);
and U7875 (N_7875,N_5040,N_6266);
nand U7876 (N_7876,N_5693,N_6222);
or U7877 (N_7877,N_6953,N_5531);
and U7878 (N_7878,N_7278,N_6926);
and U7879 (N_7879,N_5338,N_7306);
xor U7880 (N_7880,N_6089,N_6880);
nand U7881 (N_7881,N_7317,N_6571);
and U7882 (N_7882,N_5602,N_5303);
and U7883 (N_7883,N_5454,N_6486);
and U7884 (N_7884,N_7416,N_6678);
nor U7885 (N_7885,N_6361,N_7030);
nand U7886 (N_7886,N_6785,N_6795);
nand U7887 (N_7887,N_5590,N_6802);
nor U7888 (N_7888,N_6838,N_6455);
xor U7889 (N_7889,N_6874,N_5720);
or U7890 (N_7890,N_5572,N_5318);
and U7891 (N_7891,N_6217,N_6882);
xor U7892 (N_7892,N_6097,N_6330);
nand U7893 (N_7893,N_6344,N_5850);
nand U7894 (N_7894,N_5877,N_6715);
and U7895 (N_7895,N_5090,N_5455);
nand U7896 (N_7896,N_7285,N_6740);
xor U7897 (N_7897,N_6799,N_7311);
or U7898 (N_7898,N_5630,N_5348);
or U7899 (N_7899,N_6346,N_7010);
nand U7900 (N_7900,N_7488,N_6213);
nor U7901 (N_7901,N_7009,N_6808);
nand U7902 (N_7902,N_6042,N_5857);
nand U7903 (N_7903,N_6508,N_5781);
nand U7904 (N_7904,N_5430,N_5697);
xnor U7905 (N_7905,N_5797,N_5952);
nor U7906 (N_7906,N_6702,N_7402);
and U7907 (N_7907,N_5744,N_7182);
nor U7908 (N_7908,N_5983,N_7048);
xnor U7909 (N_7909,N_6536,N_5858);
and U7910 (N_7910,N_5022,N_7207);
xnor U7911 (N_7911,N_7409,N_6655);
nor U7912 (N_7912,N_5681,N_5570);
and U7913 (N_7913,N_7151,N_6141);
xnor U7914 (N_7914,N_7090,N_6958);
nand U7915 (N_7915,N_6792,N_6377);
nor U7916 (N_7916,N_5221,N_6458);
or U7917 (N_7917,N_5036,N_5496);
or U7918 (N_7918,N_6658,N_6966);
or U7919 (N_7919,N_6105,N_5108);
or U7920 (N_7920,N_5831,N_6139);
and U7921 (N_7921,N_6258,N_6431);
nor U7922 (N_7922,N_6166,N_7057);
nand U7923 (N_7923,N_5764,N_5909);
and U7924 (N_7924,N_7290,N_5180);
xnor U7925 (N_7925,N_6334,N_6414);
or U7926 (N_7926,N_6138,N_5766);
nor U7927 (N_7927,N_6676,N_6761);
nand U7928 (N_7928,N_5665,N_5163);
nor U7929 (N_7929,N_5947,N_6690);
nor U7930 (N_7930,N_6590,N_6352);
nor U7931 (N_7931,N_7310,N_5298);
and U7932 (N_7932,N_6424,N_6108);
xnor U7933 (N_7933,N_6706,N_7466);
or U7934 (N_7934,N_6398,N_7117);
or U7935 (N_7935,N_5270,N_6276);
nand U7936 (N_7936,N_7423,N_5229);
nand U7937 (N_7937,N_5392,N_5915);
and U7938 (N_7938,N_6391,N_7077);
and U7939 (N_7939,N_5824,N_6350);
nand U7940 (N_7940,N_7186,N_5592);
or U7941 (N_7941,N_5842,N_6256);
xor U7942 (N_7942,N_7422,N_6152);
nand U7943 (N_7943,N_6409,N_7315);
xnor U7944 (N_7944,N_7047,N_6662);
nand U7945 (N_7945,N_7021,N_7325);
or U7946 (N_7946,N_5255,N_6846);
xnor U7947 (N_7947,N_6206,N_5076);
nor U7948 (N_7948,N_5511,N_5235);
nor U7949 (N_7949,N_6950,N_5643);
or U7950 (N_7950,N_6086,N_5754);
and U7951 (N_7951,N_5502,N_5760);
nand U7952 (N_7952,N_7162,N_5441);
xnor U7953 (N_7953,N_5529,N_7451);
and U7954 (N_7954,N_6511,N_5679);
nand U7955 (N_7955,N_5072,N_6159);
nor U7956 (N_7956,N_5155,N_7356);
nor U7957 (N_7957,N_5743,N_7396);
or U7958 (N_7958,N_5729,N_5304);
nand U7959 (N_7959,N_5488,N_6666);
and U7960 (N_7960,N_7431,N_5678);
nand U7961 (N_7961,N_6873,N_5702);
nand U7962 (N_7962,N_6126,N_7320);
nand U7963 (N_7963,N_5080,N_5717);
xnor U7964 (N_7964,N_7312,N_5279);
or U7965 (N_7965,N_7141,N_6031);
xnor U7966 (N_7966,N_6981,N_6868);
or U7967 (N_7967,N_6143,N_6973);
nand U7968 (N_7968,N_7281,N_6025);
nand U7969 (N_7969,N_6047,N_5228);
xor U7970 (N_7970,N_7297,N_7198);
or U7971 (N_7971,N_6593,N_5295);
and U7972 (N_7972,N_5931,N_5686);
or U7973 (N_7973,N_5763,N_6366);
or U7974 (N_7974,N_5780,N_5607);
xor U7975 (N_7975,N_5979,N_5704);
or U7976 (N_7976,N_5835,N_5047);
xor U7977 (N_7977,N_5765,N_6599);
nand U7978 (N_7978,N_5044,N_7213);
or U7979 (N_7979,N_6995,N_6931);
nand U7980 (N_7980,N_7377,N_5405);
nor U7981 (N_7981,N_7199,N_6393);
nand U7982 (N_7982,N_5453,N_6362);
nand U7983 (N_7983,N_7093,N_7274);
xor U7984 (N_7984,N_6672,N_6249);
and U7985 (N_7985,N_6913,N_6278);
nor U7986 (N_7986,N_6777,N_5506);
or U7987 (N_7987,N_5933,N_5475);
and U7988 (N_7988,N_5566,N_5096);
or U7989 (N_7989,N_5805,N_7359);
nand U7990 (N_7990,N_6311,N_6035);
nor U7991 (N_7991,N_5086,N_7462);
and U7992 (N_7992,N_5734,N_5919);
nand U7993 (N_7993,N_6574,N_6900);
and U7994 (N_7994,N_5606,N_5373);
and U7995 (N_7995,N_7011,N_6983);
and U7996 (N_7996,N_6559,N_5761);
nor U7997 (N_7997,N_6661,N_7003);
and U7998 (N_7998,N_5728,N_6659);
nor U7999 (N_7999,N_5016,N_5990);
and U8000 (N_8000,N_6818,N_6209);
nor U8001 (N_8001,N_7335,N_6054);
or U8002 (N_8002,N_6698,N_6153);
nand U8003 (N_8003,N_5779,N_7111);
nand U8004 (N_8004,N_6783,N_5474);
nand U8005 (N_8005,N_6348,N_5191);
or U8006 (N_8006,N_6464,N_5057);
and U8007 (N_8007,N_6102,N_6247);
nor U8008 (N_8008,N_6689,N_5005);
and U8009 (N_8009,N_5817,N_6207);
nand U8010 (N_8010,N_5612,N_6171);
xnor U8011 (N_8011,N_6460,N_6612);
xor U8012 (N_8012,N_7339,N_6299);
nand U8013 (N_8013,N_5462,N_5174);
xnor U8014 (N_8014,N_6978,N_6115);
xor U8015 (N_8015,N_6195,N_6623);
or U8016 (N_8016,N_7239,N_6103);
nand U8017 (N_8017,N_6829,N_5890);
xnor U8018 (N_8018,N_5436,N_5065);
and U8019 (N_8019,N_6685,N_6639);
or U8020 (N_8020,N_6977,N_7079);
nor U8021 (N_8021,N_5355,N_5420);
nor U8022 (N_8022,N_7134,N_7373);
and U8023 (N_8023,N_6758,N_5629);
and U8024 (N_8024,N_6549,N_7102);
and U8025 (N_8025,N_5225,N_6267);
and U8026 (N_8026,N_7360,N_5287);
nor U8027 (N_8027,N_6866,N_7295);
and U8028 (N_8028,N_5541,N_6997);
xor U8029 (N_8029,N_7479,N_5627);
and U8030 (N_8030,N_6494,N_5311);
or U8031 (N_8031,N_7209,N_6136);
or U8032 (N_8032,N_7042,N_7108);
xor U8033 (N_8033,N_6204,N_5969);
or U8034 (N_8034,N_7078,N_6327);
nor U8035 (N_8035,N_6478,N_5212);
and U8036 (N_8036,N_7355,N_7318);
nand U8037 (N_8037,N_7340,N_5964);
and U8038 (N_8038,N_6863,N_5121);
xnor U8039 (N_8039,N_6011,N_6636);
nor U8040 (N_8040,N_5187,N_6667);
xor U8041 (N_8041,N_6092,N_7178);
nor U8042 (N_8042,N_5153,N_5677);
or U8043 (N_8043,N_6772,N_7050);
or U8044 (N_8044,N_5289,N_5816);
nor U8045 (N_8045,N_6620,N_6546);
and U8046 (N_8046,N_6720,N_6989);
xor U8047 (N_8047,N_5053,N_6170);
nand U8048 (N_8048,N_7379,N_7217);
and U8049 (N_8049,N_6061,N_6482);
and U8050 (N_8050,N_6317,N_5009);
and U8051 (N_8051,N_7253,N_6363);
nor U8052 (N_8052,N_5164,N_6696);
and U8053 (N_8053,N_5613,N_6775);
xnor U8054 (N_8054,N_5700,N_6190);
nand U8055 (N_8055,N_7062,N_5545);
or U8056 (N_8056,N_6079,N_5340);
and U8057 (N_8057,N_5565,N_5950);
nand U8058 (N_8058,N_5142,N_5390);
xor U8059 (N_8059,N_5069,N_6076);
and U8060 (N_8060,N_5209,N_5991);
nor U8061 (N_8061,N_5594,N_6504);
nor U8062 (N_8062,N_5177,N_6797);
xor U8063 (N_8063,N_5484,N_6854);
nand U8064 (N_8064,N_5573,N_7231);
and U8065 (N_8065,N_6253,N_5715);
and U8066 (N_8066,N_5231,N_5208);
nor U8067 (N_8067,N_7033,N_5151);
nor U8068 (N_8068,N_5470,N_6403);
nor U8069 (N_8069,N_6524,N_6447);
xnor U8070 (N_8070,N_6697,N_5489);
nand U8071 (N_8071,N_5651,N_6453);
or U8072 (N_8072,N_7073,N_6070);
or U8073 (N_8073,N_5409,N_6026);
nand U8074 (N_8074,N_7046,N_6008);
and U8075 (N_8075,N_7493,N_6370);
and U8076 (N_8076,N_5039,N_5603);
nand U8077 (N_8077,N_5904,N_5285);
nand U8078 (N_8078,N_5926,N_5636);
or U8079 (N_8079,N_6565,N_6229);
and U8080 (N_8080,N_6226,N_5672);
nor U8081 (N_8081,N_7100,N_5112);
nor U8082 (N_8082,N_7435,N_5066);
and U8083 (N_8083,N_5061,N_7237);
nor U8084 (N_8084,N_7263,N_5957);
xor U8085 (N_8085,N_6392,N_6287);
and U8086 (N_8086,N_5395,N_5928);
nor U8087 (N_8087,N_5122,N_5609);
and U8088 (N_8088,N_6373,N_5918);
xnor U8089 (N_8089,N_5232,N_6845);
nand U8090 (N_8090,N_5149,N_7056);
or U8091 (N_8091,N_6059,N_5965);
and U8092 (N_8092,N_5433,N_6522);
nand U8093 (N_8093,N_5988,N_5101);
and U8094 (N_8094,N_6876,N_7276);
or U8095 (N_8095,N_5823,N_5945);
nor U8096 (N_8096,N_6088,N_5943);
nand U8097 (N_8097,N_5404,N_5169);
and U8098 (N_8098,N_5173,N_5997);
nor U8099 (N_8099,N_5683,N_6385);
xnor U8100 (N_8100,N_7307,N_6787);
or U8101 (N_8101,N_5087,N_5874);
xor U8102 (N_8102,N_5758,N_6625);
nor U8103 (N_8103,N_5202,N_6376);
and U8104 (N_8104,N_5682,N_5811);
nand U8105 (N_8105,N_6461,N_6410);
nand U8106 (N_8106,N_5194,N_7378);
nor U8107 (N_8107,N_7283,N_6605);
and U8108 (N_8108,N_7401,N_6325);
nand U8109 (N_8109,N_7461,N_5593);
or U8110 (N_8110,N_5292,N_5418);
or U8111 (N_8111,N_5716,N_6734);
nand U8112 (N_8112,N_6768,N_6452);
nor U8113 (N_8113,N_5516,N_5532);
nor U8114 (N_8114,N_5063,N_5415);
xor U8115 (N_8115,N_7459,N_7309);
and U8116 (N_8116,N_6683,N_6822);
nand U8117 (N_8117,N_6839,N_6633);
nor U8118 (N_8118,N_6917,N_5434);
and U8119 (N_8119,N_5334,N_5822);
nor U8120 (N_8120,N_5237,N_5668);
xnor U8121 (N_8121,N_6474,N_5028);
xor U8122 (N_8122,N_7280,N_5903);
or U8123 (N_8123,N_6764,N_6789);
nor U8124 (N_8124,N_6918,N_7303);
xnor U8125 (N_8125,N_6005,N_5986);
or U8126 (N_8126,N_5711,N_6731);
nor U8127 (N_8127,N_6577,N_5830);
and U8128 (N_8128,N_6798,N_6519);
nor U8129 (N_8129,N_5601,N_7110);
and U8130 (N_8130,N_5587,N_7227);
or U8131 (N_8131,N_5054,N_7161);
xor U8132 (N_8132,N_7014,N_5808);
xor U8133 (N_8133,N_5472,N_6811);
or U8134 (N_8134,N_5923,N_5944);
nand U8135 (N_8135,N_7081,N_6462);
nor U8136 (N_8136,N_6708,N_6823);
or U8137 (N_8137,N_5469,N_6579);
nand U8138 (N_8138,N_5910,N_6637);
or U8139 (N_8139,N_6645,N_5259);
or U8140 (N_8140,N_5233,N_6073);
xor U8141 (N_8141,N_5451,N_5154);
or U8142 (N_8142,N_6946,N_6428);
and U8143 (N_8143,N_5222,N_6479);
nand U8144 (N_8144,N_6384,N_7272);
nand U8145 (N_8145,N_6349,N_5777);
xnor U8146 (N_8146,N_6832,N_7319);
nor U8147 (N_8147,N_6032,N_6448);
nor U8148 (N_8148,N_5265,N_5981);
nand U8149 (N_8149,N_7254,N_5306);
or U8150 (N_8150,N_5970,N_7132);
nor U8151 (N_8151,N_5887,N_5327);
or U8152 (N_8152,N_5650,N_6252);
and U8153 (N_8153,N_5960,N_5847);
nor U8154 (N_8154,N_5144,N_6784);
and U8155 (N_8155,N_5971,N_5414);
nand U8156 (N_8156,N_5530,N_5642);
and U8157 (N_8157,N_7332,N_5838);
and U8158 (N_8158,N_6603,N_5280);
or U8159 (N_8159,N_6591,N_7368);
or U8160 (N_8160,N_5393,N_7223);
and U8161 (N_8161,N_7499,N_7490);
nand U8162 (N_8162,N_6824,N_6686);
nand U8163 (N_8163,N_5775,N_5714);
xnor U8164 (N_8164,N_6435,N_6763);
xnor U8165 (N_8165,N_5332,N_6957);
and U8166 (N_8166,N_5422,N_5658);
and U8167 (N_8167,N_5073,N_7013);
nor U8168 (N_8168,N_7397,N_5662);
nand U8169 (N_8169,N_5328,N_7018);
xor U8170 (N_8170,N_5118,N_5999);
nor U8171 (N_8171,N_6386,N_5319);
or U8172 (N_8172,N_6680,N_5085);
nand U8173 (N_8173,N_6728,N_6314);
nand U8174 (N_8174,N_6956,N_5001);
nor U8175 (N_8175,N_5504,N_5810);
nor U8176 (N_8176,N_5599,N_5021);
nand U8177 (N_8177,N_5792,N_6057);
or U8178 (N_8178,N_6286,N_7144);
nand U8179 (N_8179,N_6118,N_5738);
xor U8180 (N_8180,N_6145,N_5956);
nand U8181 (N_8181,N_5614,N_5620);
or U8182 (N_8182,N_5019,N_6466);
nand U8183 (N_8183,N_5967,N_7204);
xnor U8184 (N_8184,N_6916,N_6602);
xor U8185 (N_8185,N_5820,N_6897);
or U8186 (N_8186,N_7211,N_7323);
nand U8187 (N_8187,N_6001,N_7169);
and U8188 (N_8188,N_5604,N_6492);
nand U8189 (N_8189,N_6390,N_5867);
nand U8190 (N_8190,N_6117,N_6016);
or U8191 (N_8191,N_5670,N_5056);
xor U8192 (N_8192,N_5798,N_5776);
and U8193 (N_8193,N_7121,N_6284);
and U8194 (N_8194,N_5753,N_7432);
or U8195 (N_8195,N_6694,N_5179);
or U8196 (N_8196,N_5556,N_5196);
and U8197 (N_8197,N_6183,N_7058);
nand U8198 (N_8198,N_6285,N_6040);
nor U8199 (N_8199,N_5406,N_7385);
xor U8200 (N_8200,N_6329,N_5929);
nand U8201 (N_8201,N_5413,N_7449);
nand U8202 (N_8202,N_7258,N_5026);
nand U8203 (N_8203,N_7471,N_5631);
xnor U8204 (N_8204,N_7087,N_7348);
xnor U8205 (N_8205,N_5308,N_6144);
xor U8206 (N_8206,N_5561,N_6500);
nor U8207 (N_8207,N_5251,N_5951);
nor U8208 (N_8208,N_5552,N_7224);
nand U8209 (N_8209,N_6529,N_7390);
xnor U8210 (N_8210,N_6137,N_6322);
and U8211 (N_8211,N_7498,N_5023);
or U8212 (N_8212,N_7436,N_5134);
nand U8213 (N_8213,N_6225,N_6233);
nand U8214 (N_8214,N_6289,N_7412);
and U8215 (N_8215,N_5181,N_6381);
and U8216 (N_8216,N_6971,N_7474);
nand U8217 (N_8217,N_7007,N_5819);
xor U8218 (N_8218,N_5859,N_5033);
xor U8219 (N_8219,N_6096,N_5568);
and U8220 (N_8220,N_6319,N_6701);
nor U8221 (N_8221,N_5902,N_7384);
xnor U8222 (N_8222,N_6292,N_5680);
xnor U8223 (N_8223,N_5197,N_5578);
and U8224 (N_8224,N_5322,N_6470);
and U8225 (N_8225,N_7065,N_7114);
xor U8226 (N_8226,N_6679,N_6954);
nor U8227 (N_8227,N_6497,N_5628);
or U8228 (N_8228,N_6020,N_7017);
and U8229 (N_8229,N_6214,N_6128);
nand U8230 (N_8230,N_7465,N_5239);
nand U8231 (N_8231,N_7006,N_6635);
xor U8232 (N_8232,N_5189,N_5998);
nor U8233 (N_8233,N_7414,N_5724);
and U8234 (N_8234,N_7467,N_5070);
xnor U8235 (N_8235,N_7187,N_5220);
or U8236 (N_8236,N_5081,N_5807);
or U8237 (N_8237,N_6463,N_6700);
xnor U8238 (N_8238,N_5920,N_5710);
nand U8239 (N_8239,N_6421,N_5900);
and U8240 (N_8240,N_6955,N_7341);
and U8241 (N_8241,N_5010,N_6525);
nand U8242 (N_8242,N_5437,N_6210);
nor U8243 (N_8243,N_6383,N_5655);
or U8244 (N_8244,N_7249,N_5921);
and U8245 (N_8245,N_7301,N_6454);
xor U8246 (N_8246,N_6864,N_6423);
nor U8247 (N_8247,N_5942,N_7456);
nand U8248 (N_8248,N_5246,N_6850);
or U8249 (N_8249,N_6999,N_6800);
nor U8250 (N_8250,N_5804,N_6752);
or U8251 (N_8251,N_5375,N_6400);
nor U8252 (N_8252,N_6947,N_5855);
xor U8253 (N_8253,N_5705,N_7103);
nor U8254 (N_8254,N_6558,N_7286);
or U8255 (N_8255,N_7324,N_7468);
xnor U8256 (N_8256,N_6127,N_5828);
or U8257 (N_8257,N_7413,N_7287);
or U8258 (N_8258,N_6509,N_7230);
or U8259 (N_8259,N_6446,N_6038);
and U8260 (N_8260,N_5321,N_5768);
nor U8261 (N_8261,N_6563,N_5345);
and U8262 (N_8262,N_5795,N_7150);
nor U8263 (N_8263,N_7040,N_7426);
or U8264 (N_8264,N_7034,N_5283);
nand U8265 (N_8265,N_5109,N_6307);
nand U8266 (N_8266,N_6493,N_5712);
nand U8267 (N_8267,N_5058,N_6388);
nor U8268 (N_8268,N_6132,N_5419);
nor U8269 (N_8269,N_5708,N_6293);
xnor U8270 (N_8270,N_5769,N_6730);
nand U8271 (N_8271,N_6626,N_5987);
nand U8272 (N_8272,N_6892,N_6107);
and U8273 (N_8273,N_5567,N_5550);
nand U8274 (N_8274,N_5786,N_5099);
nand U8275 (N_8275,N_5272,N_5523);
or U8276 (N_8276,N_6037,N_7404);
xor U8277 (N_8277,N_6150,N_5401);
xor U8278 (N_8278,N_5236,N_6673);
nand U8279 (N_8279,N_7475,N_5821);
xor U8280 (N_8280,N_6009,N_7485);
xor U8281 (N_8281,N_6885,N_5864);
and U8282 (N_8282,N_5868,N_5701);
nand U8283 (N_8283,N_7374,N_7235);
and U8284 (N_8284,N_5539,N_5082);
or U8285 (N_8285,N_6776,N_7195);
xor U8286 (N_8286,N_7403,N_5105);
nand U8287 (N_8287,N_6932,N_5845);
or U8288 (N_8288,N_6326,N_7444);
nand U8289 (N_8289,N_5184,N_6632);
and U8290 (N_8290,N_7302,N_6541);
nor U8291 (N_8291,N_5083,N_7159);
nor U8292 (N_8292,N_7458,N_6451);
nand U8293 (N_8293,N_6416,N_6615);
and U8294 (N_8294,N_7447,N_6765);
and U8295 (N_8295,N_5584,N_5465);
nand U8296 (N_8296,N_5588,N_6199);
or U8297 (N_8297,N_5172,N_6274);
and U8298 (N_8298,N_5030,N_5483);
nor U8299 (N_8299,N_7439,N_6907);
and U8300 (N_8300,N_7228,N_5827);
xnor U8301 (N_8301,N_6053,N_6855);
and U8302 (N_8302,N_7105,N_7273);
or U8303 (N_8303,N_5402,N_6749);
and U8304 (N_8304,N_7064,N_6968);
xor U8305 (N_8305,N_5015,N_5494);
xor U8306 (N_8306,N_5917,N_6515);
or U8307 (N_8307,N_7060,N_5492);
or U8308 (N_8308,N_6704,N_6903);
xnor U8309 (N_8309,N_7067,N_5271);
nor U8310 (N_8310,N_6616,N_5896);
and U8311 (N_8311,N_6975,N_5689);
nor U8312 (N_8312,N_7175,N_5869);
nand U8313 (N_8313,N_7445,N_7282);
xor U8314 (N_8314,N_6786,N_6245);
or U8315 (N_8315,N_5589,N_5011);
or U8316 (N_8316,N_6647,N_6119);
xnor U8317 (N_8317,N_6712,N_6856);
or U8318 (N_8318,N_5025,N_6905);
xnor U8319 (N_8319,N_5537,N_6369);
nand U8320 (N_8320,N_6886,N_5481);
or U8321 (N_8321,N_5051,N_6339);
xnor U8322 (N_8322,N_7106,N_6182);
or U8323 (N_8323,N_6928,N_6770);
or U8324 (N_8324,N_7219,N_7215);
or U8325 (N_8325,N_5183,N_5598);
and U8326 (N_8326,N_5722,N_6263);
or U8327 (N_8327,N_6420,N_6002);
and U8328 (N_8328,N_6343,N_5745);
nand U8329 (N_8329,N_5575,N_6122);
nor U8330 (N_8330,N_6695,N_6279);
xnor U8331 (N_8331,N_6264,N_6228);
nand U8332 (N_8332,N_7039,N_6281);
nor U8333 (N_8333,N_5358,N_5818);
and U8334 (N_8334,N_5757,N_7131);
nand U8335 (N_8335,N_6569,N_6341);
nor U8336 (N_8336,N_7313,N_6861);
xor U8337 (N_8337,N_5032,N_5098);
xnor U8338 (N_8338,N_6534,N_6959);
and U8339 (N_8339,N_5739,N_6847);
or U8340 (N_8340,N_7321,N_6355);
or U8341 (N_8341,N_6967,N_5352);
xor U8342 (N_8342,N_5645,N_5698);
nand U8343 (N_8343,N_7020,N_6389);
xor U8344 (N_8344,N_5249,N_6048);
xor U8345 (N_8345,N_6929,N_5571);
nor U8346 (N_8346,N_7305,N_6589);
nor U8347 (N_8347,N_6809,N_6523);
or U8348 (N_8348,N_5038,N_6738);
nor U8349 (N_8349,N_6936,N_5186);
and U8350 (N_8350,N_6193,N_6068);
nand U8351 (N_8351,N_5721,N_6767);
and U8352 (N_8352,N_6909,N_5789);
nor U8353 (N_8353,N_7152,N_6544);
nor U8354 (N_8354,N_6614,N_6056);
xnor U8355 (N_8355,N_6528,N_5888);
and U8356 (N_8356,N_5178,N_5094);
nand U8357 (N_8357,N_5120,N_7260);
nor U8358 (N_8358,N_6849,N_7369);
nor U8359 (N_8359,N_5006,N_7080);
or U8360 (N_8360,N_5707,N_6554);
nor U8361 (N_8361,N_6238,N_5138);
and U8362 (N_8362,N_5326,N_6246);
and U8363 (N_8363,N_7153,N_5898);
nor U8364 (N_8364,N_5012,N_7329);
nor U8365 (N_8365,N_6532,N_5889);
or U8366 (N_8366,N_5150,N_5002);
nand U8367 (N_8367,N_5652,N_5031);
xor U8368 (N_8368,N_6705,N_7460);
and U8369 (N_8369,N_7041,N_5397);
nand U8370 (N_8370,N_7470,N_6411);
xnor U8371 (N_8371,N_6991,N_6996);
nand U8372 (N_8372,N_5580,N_5214);
or U8373 (N_8373,N_5713,N_6471);
and U8374 (N_8374,N_5879,N_7298);
nand U8375 (N_8375,N_7171,N_5331);
or U8376 (N_8376,N_6578,N_6272);
nor U8377 (N_8377,N_6714,N_6883);
xor U8378 (N_8378,N_5479,N_5388);
or U8379 (N_8379,N_6677,N_5784);
nand U8380 (N_8380,N_5740,N_5863);
or U8381 (N_8381,N_6908,N_5145);
and U8382 (N_8382,N_5968,N_7174);
nand U8383 (N_8383,N_5277,N_7382);
or U8384 (N_8384,N_7099,N_6747);
and U8385 (N_8385,N_6058,N_5659);
nand U8386 (N_8386,N_5688,N_6162);
xor U8387 (N_8387,N_5190,N_5368);
nor U8388 (N_8388,N_5320,N_6260);
nand U8389 (N_8389,N_6606,N_5974);
or U8390 (N_8390,N_6835,N_6890);
xor U8391 (N_8391,N_7261,N_5834);
and U8392 (N_8392,N_7279,N_6642);
nand U8393 (N_8393,N_6518,N_6239);
xnor U8394 (N_8394,N_6587,N_7088);
nand U8395 (N_8395,N_6816,N_6711);
nor U8396 (N_8396,N_7346,N_6449);
xnor U8397 (N_8397,N_6445,N_6469);
nand U8398 (N_8398,N_5911,N_5215);
nand U8399 (N_8399,N_5111,N_6938);
xnor U8400 (N_8400,N_5432,N_6937);
nor U8401 (N_8401,N_6135,N_5199);
xnor U8402 (N_8402,N_5324,N_6444);
xor U8403 (N_8403,N_6168,N_6161);
nor U8404 (N_8404,N_6133,N_5851);
nor U8405 (N_8405,N_5316,N_6871);
nand U8406 (N_8406,N_5463,N_5610);
nor U8407 (N_8407,N_5307,N_7212);
and U8408 (N_8408,N_5646,N_5953);
or U8409 (N_8409,N_5464,N_6505);
nand U8410 (N_8410,N_5676,N_6429);
nor U8411 (N_8411,N_5622,N_7314);
xnor U8412 (N_8412,N_5213,N_6813);
nor U8413 (N_8413,N_6803,N_7364);
nand U8414 (N_8414,N_6110,N_7478);
xor U8415 (N_8415,N_7406,N_5490);
nor U8416 (N_8416,N_5095,N_7345);
nand U8417 (N_8417,N_5663,N_7135);
nand U8418 (N_8418,N_6142,N_6315);
or U8419 (N_8419,N_5412,N_6723);
nand U8420 (N_8420,N_6151,N_5372);
nand U8421 (N_8421,N_6530,N_5759);
nor U8422 (N_8422,N_5773,N_6762);
or U8423 (N_8423,N_5671,N_6041);
xor U8424 (N_8424,N_6681,N_6313);
or U8425 (N_8425,N_7119,N_5349);
nand U8426 (N_8426,N_5024,N_5637);
nand U8427 (N_8427,N_5424,N_5922);
or U8428 (N_8428,N_6387,N_5509);
nand U8429 (N_8429,N_5542,N_5491);
and U8430 (N_8430,N_6465,N_5442);
and U8431 (N_8431,N_5569,N_7370);
or U8432 (N_8432,N_6674,N_6215);
or U8433 (N_8433,N_5696,N_5317);
nor U8434 (N_8434,N_5286,N_5262);
xnor U8435 (N_8435,N_5399,N_5068);
nand U8436 (N_8436,N_6601,N_6812);
nand U8437 (N_8437,N_6627,N_6567);
nor U8438 (N_8438,N_6675,N_6406);
nand U8439 (N_8439,N_5930,N_5583);
or U8440 (N_8440,N_6827,N_5136);
or U8441 (N_8441,N_7051,N_5871);
nor U8442 (N_8442,N_6163,N_6345);
nor U8443 (N_8443,N_7044,N_6167);
nand U8444 (N_8444,N_5559,N_6751);
and U8445 (N_8445,N_5684,N_5623);
or U8446 (N_8446,N_6609,N_5895);
xnor U8447 (N_8447,N_6687,N_6501);
xnor U8448 (N_8448,N_5690,N_6538);
xnor U8449 (N_8449,N_7197,N_7244);
nand U8450 (N_8450,N_5244,N_5383);
nand U8451 (N_8451,N_5278,N_6607);
and U8452 (N_8452,N_7452,N_6098);
and U8453 (N_8453,N_5329,N_6858);
nand U8454 (N_8454,N_7264,N_6540);
nor U8455 (N_8455,N_5106,N_6948);
and U8456 (N_8456,N_5907,N_7139);
and U8457 (N_8457,N_7420,N_5264);
nand U8458 (N_8458,N_6742,N_5814);
nand U8459 (N_8459,N_5647,N_5505);
nand U8460 (N_8460,N_5485,N_5400);
and U8461 (N_8461,N_5524,N_5143);
or U8462 (N_8462,N_7052,N_5501);
nand U8463 (N_8463,N_5377,N_7421);
nor U8464 (N_8464,N_6807,N_5123);
and U8465 (N_8465,N_7362,N_7142);
or U8466 (N_8466,N_6732,N_5290);
xor U8467 (N_8467,N_6862,N_5656);
or U8468 (N_8468,N_6181,N_5315);
xor U8469 (N_8469,N_5551,N_5034);
xor U8470 (N_8470,N_7122,N_5078);
nor U8471 (N_8471,N_5421,N_5165);
nand U8472 (N_8472,N_5125,N_6817);
or U8473 (N_8473,N_5276,N_6899);
or U8474 (N_8474,N_7233,N_5829);
and U8475 (N_8475,N_5224,N_5585);
nor U8476 (N_8476,N_5876,N_7259);
and U8477 (N_8477,N_7203,N_6081);
nor U8478 (N_8478,N_7395,N_5924);
nor U8479 (N_8479,N_5093,N_5060);
nor U8480 (N_8480,N_6017,N_5166);
or U8481 (N_8481,N_7336,N_5428);
xor U8482 (N_8482,N_6585,N_6472);
or U8483 (N_8483,N_6291,N_5055);
and U8484 (N_8484,N_5908,N_6750);
nor U8485 (N_8485,N_7375,N_6114);
or U8486 (N_8486,N_6280,N_5364);
nor U8487 (N_8487,N_5128,N_5206);
xnor U8488 (N_8488,N_5732,N_6124);
or U8489 (N_8489,N_6788,N_7083);
xor U8490 (N_8490,N_7248,N_6184);
and U8491 (N_8491,N_6399,N_7049);
and U8492 (N_8492,N_5772,N_5203);
nand U8493 (N_8493,N_6895,N_6707);
nand U8494 (N_8494,N_7089,N_6255);
xnor U8495 (N_8495,N_7450,N_6933);
nor U8496 (N_8496,N_7361,N_7358);
nand U8497 (N_8497,N_6710,N_5156);
nor U8498 (N_8498,N_5234,N_5913);
nand U8499 (N_8499,N_5346,N_5258);
or U8500 (N_8500,N_5448,N_5211);
xor U8501 (N_8501,N_5148,N_7154);
and U8502 (N_8502,N_6521,N_5927);
or U8503 (N_8503,N_6033,N_6487);
or U8504 (N_8504,N_6942,N_6555);
and U8505 (N_8505,N_6191,N_7193);
or U8506 (N_8506,N_5538,N_7069);
xor U8507 (N_8507,N_6924,N_6358);
xnor U8508 (N_8508,N_5495,N_6197);
xnor U8509 (N_8509,N_5443,N_7408);
xor U8510 (N_8510,N_7434,N_5755);
or U8511 (N_8511,N_5378,N_7214);
nand U8512 (N_8512,N_6129,N_6889);
nand U8513 (N_8513,N_6630,N_5416);
and U8514 (N_8514,N_7055,N_5440);
xor U8515 (N_8515,N_7129,N_5296);
nand U8516 (N_8516,N_6848,N_7216);
nor U8517 (N_8517,N_7027,N_6160);
nor U8518 (N_8518,N_5826,N_6134);
xnor U8519 (N_8519,N_5230,N_6531);
nand U8520 (N_8520,N_6513,N_5870);
nor U8521 (N_8521,N_6560,N_6691);
nand U8522 (N_8522,N_5840,N_6982);
nor U8523 (N_8523,N_5335,N_6468);
or U8524 (N_8524,N_6925,N_6254);
and U8525 (N_8525,N_7183,N_6548);
nor U8526 (N_8526,N_7288,N_7096);
nor U8527 (N_8527,N_6944,N_7350);
nand U8528 (N_8528,N_6618,N_6176);
nor U8529 (N_8529,N_6921,N_6450);
nor U8530 (N_8530,N_6243,N_7036);
or U8531 (N_8531,N_5476,N_5674);
nand U8532 (N_8532,N_6408,N_6332);
nor U8533 (N_8533,N_6976,N_5892);
nor U8534 (N_8534,N_5730,N_7221);
nand U8535 (N_8535,N_5426,N_5167);
and U8536 (N_8536,N_5310,N_5615);
nand U8537 (N_8537,N_6972,N_5852);
xnor U8538 (N_8538,N_5293,N_6242);
nor U8539 (N_8539,N_6234,N_5846);
xnor U8540 (N_8540,N_6072,N_6810);
nor U8541 (N_8541,N_5861,N_6562);
or U8542 (N_8542,N_5323,N_5706);
and U8543 (N_8543,N_6382,N_6333);
xor U8544 (N_8544,N_6188,N_5955);
and U8545 (N_8545,N_7347,N_6065);
nand U8546 (N_8546,N_5446,N_6475);
nor U8547 (N_8547,N_6570,N_5369);
nand U8548 (N_8548,N_7146,N_5992);
nand U8549 (N_8549,N_5806,N_5843);
and U8550 (N_8550,N_5299,N_7240);
or U8551 (N_8551,N_5333,N_6044);
or U8552 (N_8552,N_6877,N_5508);
xor U8553 (N_8553,N_6613,N_7059);
and U8554 (N_8554,N_5638,N_7156);
xnor U8555 (N_8555,N_6729,N_6622);
nand U8556 (N_8556,N_6028,N_5071);
xnor U8557 (N_8557,N_5989,N_6496);
xor U8558 (N_8558,N_7084,N_7266);
nand U8559 (N_8559,N_6099,N_5751);
nand U8560 (N_8560,N_5787,N_7405);
or U8561 (N_8561,N_5139,N_5344);
nand U8562 (N_8562,N_7181,N_6598);
nand U8563 (N_8563,N_6324,N_5459);
or U8564 (N_8564,N_6790,N_5791);
xnor U8565 (N_8565,N_5555,N_5894);
nor U8566 (N_8566,N_6557,N_6527);
nor U8567 (N_8567,N_6748,N_7202);
nor U8568 (N_8568,N_6654,N_6782);
and U8569 (N_8569,N_6507,N_6884);
nor U8570 (N_8570,N_6898,N_6397);
nor U8571 (N_8571,N_7188,N_6796);
nor U8572 (N_8572,N_5790,N_6231);
xnor U8573 (N_8573,N_7400,N_6927);
xnor U8574 (N_8574,N_6259,N_7229);
nand U8575 (N_8575,N_6456,N_6179);
xor U8576 (N_8576,N_6736,N_5582);
or U8577 (N_8577,N_5880,N_6024);
nor U8578 (N_8578,N_6268,N_7265);
nor U8579 (N_8579,N_6592,N_6985);
nand U8580 (N_8580,N_5274,N_6318);
nor U8581 (N_8581,N_5558,N_5380);
or U8582 (N_8582,N_5158,N_5043);
nand U8583 (N_8583,N_5946,N_5193);
nand U8584 (N_8584,N_6914,N_6357);
and U8585 (N_8585,N_5853,N_6894);
nand U8586 (N_8586,N_6709,N_7262);
nor U8587 (N_8587,N_7180,N_7417);
nor U8588 (N_8588,N_5394,N_7177);
xnor U8589 (N_8589,N_6743,N_6125);
and U8590 (N_8590,N_7097,N_7380);
nor U8591 (N_8591,N_5914,N_5370);
or U8592 (N_8592,N_6087,N_5219);
and U8593 (N_8593,N_5029,N_5245);
nor U8594 (N_8594,N_6600,N_5079);
or U8595 (N_8595,N_5882,N_6986);
and U8596 (N_8596,N_5084,N_7075);
nand U8597 (N_8597,N_5449,N_5866);
nand U8598 (N_8598,N_6200,N_5976);
or U8599 (N_8599,N_5954,N_6652);
xnor U8600 (N_8600,N_5447,N_6561);
nor U8601 (N_8601,N_6669,N_6735);
or U8602 (N_8602,N_7246,N_5883);
and U8603 (N_8603,N_5608,N_6498);
xnor U8604 (N_8604,N_7357,N_7484);
xnor U8605 (N_8605,N_5353,N_5201);
xnor U8606 (N_8606,N_5371,N_6221);
and U8607 (N_8607,N_6230,N_5749);
nor U8608 (N_8608,N_6510,N_7053);
nand U8609 (N_8609,N_6083,N_5379);
and U8610 (N_8610,N_6380,N_6003);
or U8611 (N_8611,N_5891,N_6629);
and U8612 (N_8612,N_6158,N_6077);
and U8613 (N_8613,N_7071,N_7349);
and U8614 (N_8614,N_5027,N_6323);
nand U8615 (N_8615,N_5226,N_6473);
nand U8616 (N_8616,N_5050,N_5089);
nor U8617 (N_8617,N_7149,N_5064);
or U8618 (N_8618,N_6993,N_6227);
nor U8619 (N_8619,N_6275,N_6878);
xor U8620 (N_8620,N_5407,N_5521);
nor U8621 (N_8621,N_7220,N_6353);
nor U8622 (N_8622,N_6668,N_5799);
xnor U8623 (N_8623,N_6980,N_5878);
nor U8624 (N_8624,N_6581,N_6716);
xor U8625 (N_8625,N_6663,N_7381);
and U8626 (N_8626,N_5275,N_7419);
and U8627 (N_8627,N_5625,N_5135);
nand U8628 (N_8628,N_5770,N_5238);
or U8629 (N_8629,N_6430,N_6941);
nand U8630 (N_8630,N_5635,N_5750);
xor U8631 (N_8631,N_5389,N_7031);
xnor U8632 (N_8632,N_5905,N_7257);
nor U8633 (N_8633,N_7179,N_7398);
xor U8634 (N_8634,N_6379,N_6043);
and U8635 (N_8635,N_6422,N_6301);
or U8636 (N_8636,N_5248,N_7241);
nand U8637 (N_8637,N_6094,N_6173);
nand U8638 (N_8638,N_6923,N_6356);
or U8639 (N_8639,N_5471,N_6773);
and U8640 (N_8640,N_5940,N_5403);
nand U8641 (N_8641,N_7155,N_7143);
nor U8642 (N_8642,N_6359,N_6440);
or U8643 (N_8643,N_6045,N_5367);
or U8644 (N_8644,N_5217,N_6597);
xor U8645 (N_8645,N_5284,N_6754);
xor U8646 (N_8646,N_5984,N_6367);
xor U8647 (N_8647,N_5185,N_6771);
xnor U8648 (N_8648,N_6499,N_5425);
or U8649 (N_8649,N_7185,N_6196);
nor U8650 (N_8650,N_7331,N_6624);
nand U8651 (N_8651,N_6224,N_5048);
and U8652 (N_8652,N_6013,N_5444);
nand U8653 (N_8653,N_6841,N_6198);
nand U8654 (N_8654,N_5347,N_6090);
nand U8655 (N_8655,N_6722,N_5359);
nand U8656 (N_8656,N_5046,N_5337);
or U8657 (N_8657,N_5480,N_5836);
or U8658 (N_8658,N_7120,N_5439);
nor U8659 (N_8659,N_7367,N_6693);
and U8660 (N_8660,N_6023,N_7124);
xnor U8661 (N_8661,N_6984,N_6535);
xor U8662 (N_8662,N_5198,N_5351);
nor U8663 (N_8663,N_5269,N_5699);
or U8664 (N_8664,N_7024,N_5935);
nor U8665 (N_8665,N_7496,N_6881);
xor U8666 (N_8666,N_7076,N_7112);
nor U8667 (N_8667,N_6419,N_7029);
nand U8668 (N_8668,N_5885,N_6516);
nand U8669 (N_8669,N_6283,N_5309);
or U8670 (N_8670,N_5897,N_7477);
or U8671 (N_8671,N_7415,N_6295);
nor U8672 (N_8672,N_5313,N_5253);
and U8673 (N_8673,N_6887,N_6205);
or U8674 (N_8674,N_5152,N_6769);
nand U8675 (N_8675,N_6459,N_6604);
nand U8676 (N_8676,N_6265,N_5386);
nor U8677 (N_8677,N_7267,N_6071);
nor U8678 (N_8678,N_7222,N_6364);
or U8679 (N_8679,N_7115,N_6893);
xnor U8680 (N_8680,N_5115,N_7208);
and U8681 (N_8681,N_6727,N_7238);
and U8682 (N_8682,N_7012,N_6713);
xor U8683 (N_8683,N_6305,N_5536);
nor U8684 (N_8684,N_7486,N_5512);
nor U8685 (N_8685,N_6583,N_5325);
nand U8686 (N_8686,N_6491,N_5963);
nand U8687 (N_8687,N_7473,N_5586);
nand U8688 (N_8688,N_7376,N_5996);
nand U8689 (N_8689,N_5534,N_6340);
nand U8690 (N_8690,N_7085,N_6610);
xor U8691 (N_8691,N_7344,N_7446);
nor U8692 (N_8692,N_6852,N_6169);
xor U8693 (N_8693,N_7023,N_5962);
nand U8694 (N_8694,N_6988,N_5168);
or U8695 (N_8695,N_6282,N_7316);
and U8696 (N_8696,N_5116,N_5899);
or U8697 (N_8697,N_6539,N_7037);
or U8698 (N_8698,N_6837,N_6870);
or U8699 (N_8699,N_7322,N_6888);
nor U8700 (N_8700,N_5554,N_5977);
nand U8701 (N_8701,N_6580,N_5865);
nor U8702 (N_8702,N_7252,N_6853);
xor U8703 (N_8703,N_7487,N_6963);
nor U8704 (N_8704,N_5844,N_6477);
nand U8705 (N_8705,N_5793,N_6085);
and U8706 (N_8706,N_6990,N_7054);
xor U8707 (N_8707,N_6019,N_7167);
or U8708 (N_8708,N_5376,N_6994);
nand U8709 (N_8709,N_5540,N_7289);
or U8710 (N_8710,N_7147,N_5041);
nand U8711 (N_8711,N_5611,N_6831);
nor U8712 (N_8712,N_5018,N_6146);
or U8713 (N_8713,N_5456,N_5794);
nor U8714 (N_8714,N_5833,N_6082);
xor U8715 (N_8715,N_7296,N_6774);
and U8716 (N_8716,N_5391,N_6656);
or U8717 (N_8717,N_5452,N_5527);
xor U8718 (N_8718,N_5666,N_5254);
and U8719 (N_8719,N_5648,N_5634);
and U8720 (N_8720,N_7019,N_6029);
nand U8721 (N_8721,N_7294,N_6634);
or U8722 (N_8722,N_6826,N_6495);
or U8723 (N_8723,N_6857,N_6049);
nand U8724 (N_8724,N_6489,N_6078);
xor U8725 (N_8725,N_7330,N_6879);
and U8726 (N_8726,N_6407,N_6717);
or U8727 (N_8727,N_6915,N_7086);
and U8728 (N_8728,N_6328,N_6378);
and U8729 (N_8729,N_6123,N_5360);
xnor U8730 (N_8730,N_6935,N_5664);
nor U8731 (N_8731,N_6483,N_6741);
xor U8732 (N_8732,N_7352,N_6865);
nor U8733 (N_8733,N_5535,N_6825);
or U8734 (N_8734,N_5499,N_6791);
nand U8735 (N_8735,N_7160,N_5982);
xor U8736 (N_8736,N_5841,N_6737);
xnor U8737 (N_8737,N_5669,N_6660);
or U8738 (N_8738,N_6688,N_6699);
and U8739 (N_8739,N_6595,N_6277);
and U8740 (N_8740,N_5312,N_5042);
xnor U8741 (N_8741,N_5497,N_6684);
or U8742 (N_8742,N_5207,N_7411);
nor U8743 (N_8743,N_5302,N_7158);
nand U8744 (N_8744,N_5130,N_7476);
nor U8745 (N_8745,N_6533,N_6335);
nor U8746 (N_8746,N_5458,N_6063);
nor U8747 (N_8747,N_6952,N_6617);
or U8748 (N_8748,N_7441,N_5893);
nand U8749 (N_8749,N_6657,N_5576);
or U8750 (N_8750,N_5600,N_5242);
nand U8751 (N_8751,N_6065,N_6895);
xor U8752 (N_8752,N_5392,N_6939);
nor U8753 (N_8753,N_5721,N_5518);
nand U8754 (N_8754,N_5945,N_6468);
xnor U8755 (N_8755,N_5451,N_6784);
nand U8756 (N_8756,N_6282,N_5005);
nand U8757 (N_8757,N_5654,N_6663);
xor U8758 (N_8758,N_5883,N_7202);
xnor U8759 (N_8759,N_6730,N_6792);
nor U8760 (N_8760,N_5613,N_7229);
xor U8761 (N_8761,N_6411,N_6975);
or U8762 (N_8762,N_5265,N_6381);
nand U8763 (N_8763,N_6995,N_5108);
and U8764 (N_8764,N_5957,N_6019);
nor U8765 (N_8765,N_6634,N_6401);
and U8766 (N_8766,N_6860,N_5198);
xnor U8767 (N_8767,N_7250,N_5714);
or U8768 (N_8768,N_6853,N_5324);
or U8769 (N_8769,N_6062,N_5094);
or U8770 (N_8770,N_6748,N_5146);
xor U8771 (N_8771,N_5430,N_5464);
xor U8772 (N_8772,N_6198,N_5678);
and U8773 (N_8773,N_7357,N_5644);
or U8774 (N_8774,N_7066,N_5573);
nor U8775 (N_8775,N_7163,N_6427);
or U8776 (N_8776,N_7349,N_5357);
nand U8777 (N_8777,N_7062,N_7228);
nor U8778 (N_8778,N_5492,N_6271);
nand U8779 (N_8779,N_6632,N_6707);
nand U8780 (N_8780,N_7023,N_5359);
and U8781 (N_8781,N_6796,N_5632);
xnor U8782 (N_8782,N_7210,N_5996);
nor U8783 (N_8783,N_6259,N_5990);
nand U8784 (N_8784,N_5405,N_6837);
and U8785 (N_8785,N_5428,N_6479);
nand U8786 (N_8786,N_5075,N_6275);
xor U8787 (N_8787,N_6046,N_5550);
nand U8788 (N_8788,N_6960,N_5969);
nand U8789 (N_8789,N_6890,N_7244);
or U8790 (N_8790,N_6192,N_6126);
nor U8791 (N_8791,N_5705,N_5637);
and U8792 (N_8792,N_7032,N_5437);
or U8793 (N_8793,N_5707,N_6020);
nand U8794 (N_8794,N_5802,N_6425);
xnor U8795 (N_8795,N_5860,N_5148);
xor U8796 (N_8796,N_7483,N_6445);
xor U8797 (N_8797,N_5717,N_6470);
nand U8798 (N_8798,N_7424,N_6271);
xnor U8799 (N_8799,N_6900,N_7237);
nand U8800 (N_8800,N_6547,N_6823);
and U8801 (N_8801,N_6517,N_5606);
nand U8802 (N_8802,N_7311,N_6967);
xnor U8803 (N_8803,N_5041,N_6307);
nor U8804 (N_8804,N_6209,N_7456);
or U8805 (N_8805,N_5532,N_5385);
nand U8806 (N_8806,N_6635,N_5765);
nand U8807 (N_8807,N_6929,N_5154);
nand U8808 (N_8808,N_5480,N_5068);
or U8809 (N_8809,N_6267,N_7472);
or U8810 (N_8810,N_5579,N_6269);
nor U8811 (N_8811,N_6485,N_6501);
xnor U8812 (N_8812,N_5879,N_5410);
and U8813 (N_8813,N_6740,N_6379);
nor U8814 (N_8814,N_5058,N_6342);
nand U8815 (N_8815,N_6975,N_5825);
nor U8816 (N_8816,N_5650,N_6402);
nor U8817 (N_8817,N_6686,N_5108);
xnor U8818 (N_8818,N_6092,N_7209);
nor U8819 (N_8819,N_7228,N_6321);
and U8820 (N_8820,N_6227,N_5386);
nand U8821 (N_8821,N_6244,N_7484);
or U8822 (N_8822,N_5742,N_6398);
nand U8823 (N_8823,N_5425,N_7297);
and U8824 (N_8824,N_6365,N_6065);
and U8825 (N_8825,N_6014,N_5769);
nor U8826 (N_8826,N_5786,N_5485);
or U8827 (N_8827,N_6933,N_6416);
nand U8828 (N_8828,N_6751,N_7357);
and U8829 (N_8829,N_6692,N_6224);
and U8830 (N_8830,N_7388,N_6859);
nand U8831 (N_8831,N_6243,N_5483);
nand U8832 (N_8832,N_6578,N_6083);
nor U8833 (N_8833,N_6234,N_7421);
nor U8834 (N_8834,N_5419,N_6525);
or U8835 (N_8835,N_6315,N_5758);
and U8836 (N_8836,N_5728,N_5881);
nand U8837 (N_8837,N_5260,N_6364);
nor U8838 (N_8838,N_7227,N_6877);
nor U8839 (N_8839,N_6886,N_5384);
nor U8840 (N_8840,N_5326,N_5510);
and U8841 (N_8841,N_5539,N_5749);
and U8842 (N_8842,N_5862,N_5429);
or U8843 (N_8843,N_6724,N_6793);
nand U8844 (N_8844,N_5410,N_7019);
nor U8845 (N_8845,N_5406,N_6780);
or U8846 (N_8846,N_7179,N_5342);
nor U8847 (N_8847,N_6964,N_5816);
nand U8848 (N_8848,N_5629,N_6183);
xor U8849 (N_8849,N_6112,N_6432);
and U8850 (N_8850,N_6142,N_5203);
or U8851 (N_8851,N_5539,N_7283);
nor U8852 (N_8852,N_5256,N_7019);
nand U8853 (N_8853,N_6074,N_6000);
or U8854 (N_8854,N_5384,N_6800);
nor U8855 (N_8855,N_5857,N_7191);
nor U8856 (N_8856,N_6988,N_5296);
and U8857 (N_8857,N_5457,N_6356);
nor U8858 (N_8858,N_7234,N_6195);
and U8859 (N_8859,N_6874,N_5079);
and U8860 (N_8860,N_6422,N_5817);
and U8861 (N_8861,N_5247,N_5069);
xor U8862 (N_8862,N_6283,N_6501);
and U8863 (N_8863,N_5460,N_5321);
nor U8864 (N_8864,N_7193,N_6624);
nor U8865 (N_8865,N_7076,N_5060);
and U8866 (N_8866,N_6159,N_5641);
xnor U8867 (N_8867,N_5510,N_5515);
and U8868 (N_8868,N_5675,N_5442);
or U8869 (N_8869,N_6180,N_7434);
or U8870 (N_8870,N_6400,N_6344);
nand U8871 (N_8871,N_7048,N_7300);
or U8872 (N_8872,N_5868,N_6890);
or U8873 (N_8873,N_7424,N_5603);
nand U8874 (N_8874,N_7340,N_5200);
or U8875 (N_8875,N_6655,N_6770);
and U8876 (N_8876,N_6071,N_5023);
xnor U8877 (N_8877,N_6726,N_6193);
or U8878 (N_8878,N_6224,N_6952);
and U8879 (N_8879,N_6278,N_5371);
nor U8880 (N_8880,N_6941,N_5179);
or U8881 (N_8881,N_6003,N_6632);
and U8882 (N_8882,N_6762,N_5759);
xor U8883 (N_8883,N_7295,N_7131);
nor U8884 (N_8884,N_6785,N_5215);
and U8885 (N_8885,N_5027,N_7498);
nor U8886 (N_8886,N_5176,N_5885);
nor U8887 (N_8887,N_6660,N_5711);
and U8888 (N_8888,N_5180,N_6096);
or U8889 (N_8889,N_7138,N_6415);
and U8890 (N_8890,N_5012,N_6413);
and U8891 (N_8891,N_5470,N_5405);
and U8892 (N_8892,N_5398,N_6494);
xor U8893 (N_8893,N_5739,N_6931);
or U8894 (N_8894,N_5614,N_6764);
and U8895 (N_8895,N_7201,N_6153);
nand U8896 (N_8896,N_6232,N_5216);
or U8897 (N_8897,N_7006,N_6827);
nand U8898 (N_8898,N_6938,N_5861);
or U8899 (N_8899,N_7288,N_5394);
and U8900 (N_8900,N_7324,N_6018);
xnor U8901 (N_8901,N_6832,N_6144);
xor U8902 (N_8902,N_5470,N_6768);
and U8903 (N_8903,N_6435,N_6694);
or U8904 (N_8904,N_7163,N_7499);
xor U8905 (N_8905,N_6821,N_6922);
xor U8906 (N_8906,N_6850,N_5657);
or U8907 (N_8907,N_6680,N_7218);
nand U8908 (N_8908,N_7252,N_6522);
or U8909 (N_8909,N_5640,N_7000);
and U8910 (N_8910,N_6423,N_5924);
nand U8911 (N_8911,N_5697,N_7305);
nor U8912 (N_8912,N_5308,N_6384);
and U8913 (N_8913,N_6268,N_7045);
nand U8914 (N_8914,N_6893,N_6389);
or U8915 (N_8915,N_6295,N_6982);
xor U8916 (N_8916,N_7284,N_5567);
xnor U8917 (N_8917,N_5738,N_6988);
nor U8918 (N_8918,N_7251,N_6111);
or U8919 (N_8919,N_5846,N_6391);
xor U8920 (N_8920,N_5816,N_5874);
or U8921 (N_8921,N_6248,N_5963);
nor U8922 (N_8922,N_6411,N_6657);
and U8923 (N_8923,N_6021,N_6995);
xnor U8924 (N_8924,N_6272,N_7054);
nor U8925 (N_8925,N_5564,N_6026);
nor U8926 (N_8926,N_6507,N_7112);
nand U8927 (N_8927,N_5338,N_5208);
xnor U8928 (N_8928,N_6304,N_5982);
or U8929 (N_8929,N_5928,N_7443);
or U8930 (N_8930,N_6056,N_7401);
and U8931 (N_8931,N_5130,N_5056);
and U8932 (N_8932,N_7482,N_5030);
xnor U8933 (N_8933,N_7012,N_6293);
xnor U8934 (N_8934,N_5235,N_6815);
and U8935 (N_8935,N_6731,N_6756);
xnor U8936 (N_8936,N_5918,N_5495);
xnor U8937 (N_8937,N_6856,N_6694);
or U8938 (N_8938,N_5218,N_6803);
nand U8939 (N_8939,N_7138,N_7132);
and U8940 (N_8940,N_6713,N_5152);
and U8941 (N_8941,N_5841,N_7252);
or U8942 (N_8942,N_7199,N_5446);
nand U8943 (N_8943,N_5792,N_6970);
xor U8944 (N_8944,N_5749,N_5689);
nor U8945 (N_8945,N_6624,N_5932);
xnor U8946 (N_8946,N_6363,N_7184);
and U8947 (N_8947,N_7286,N_5955);
xor U8948 (N_8948,N_5334,N_6385);
xor U8949 (N_8949,N_5539,N_7329);
and U8950 (N_8950,N_6364,N_6189);
nand U8951 (N_8951,N_5690,N_6712);
nor U8952 (N_8952,N_6553,N_6414);
nand U8953 (N_8953,N_5208,N_5040);
and U8954 (N_8954,N_5659,N_6470);
or U8955 (N_8955,N_5260,N_5057);
nand U8956 (N_8956,N_5879,N_5808);
nand U8957 (N_8957,N_6071,N_7252);
xnor U8958 (N_8958,N_6396,N_6179);
nor U8959 (N_8959,N_7085,N_5768);
nor U8960 (N_8960,N_6900,N_7241);
or U8961 (N_8961,N_7285,N_6831);
nor U8962 (N_8962,N_5309,N_6974);
nand U8963 (N_8963,N_5218,N_6970);
nand U8964 (N_8964,N_6827,N_6121);
nand U8965 (N_8965,N_6175,N_6824);
or U8966 (N_8966,N_7302,N_5596);
or U8967 (N_8967,N_5529,N_6491);
or U8968 (N_8968,N_7332,N_5120);
nand U8969 (N_8969,N_5859,N_7396);
nor U8970 (N_8970,N_6823,N_5875);
nand U8971 (N_8971,N_5426,N_7464);
xnor U8972 (N_8972,N_7477,N_6512);
and U8973 (N_8973,N_5600,N_7005);
nor U8974 (N_8974,N_5752,N_5346);
and U8975 (N_8975,N_5448,N_7448);
and U8976 (N_8976,N_6274,N_6930);
and U8977 (N_8977,N_5249,N_5566);
xnor U8978 (N_8978,N_7021,N_6521);
xor U8979 (N_8979,N_5901,N_7425);
nand U8980 (N_8980,N_6298,N_5099);
nor U8981 (N_8981,N_6081,N_5926);
xor U8982 (N_8982,N_7328,N_5114);
and U8983 (N_8983,N_5738,N_6937);
or U8984 (N_8984,N_6929,N_7190);
and U8985 (N_8985,N_6754,N_6623);
or U8986 (N_8986,N_6314,N_6832);
or U8987 (N_8987,N_6076,N_6817);
and U8988 (N_8988,N_5430,N_7374);
xor U8989 (N_8989,N_6176,N_5152);
or U8990 (N_8990,N_5951,N_6676);
or U8991 (N_8991,N_6563,N_6529);
and U8992 (N_8992,N_6140,N_6693);
nor U8993 (N_8993,N_5880,N_7346);
and U8994 (N_8994,N_6349,N_7365);
and U8995 (N_8995,N_5509,N_5850);
xnor U8996 (N_8996,N_6120,N_6703);
and U8997 (N_8997,N_6917,N_6632);
nor U8998 (N_8998,N_5513,N_7001);
nor U8999 (N_8999,N_6201,N_7071);
and U9000 (N_9000,N_7359,N_5005);
nand U9001 (N_9001,N_6471,N_6060);
nand U9002 (N_9002,N_7283,N_5725);
or U9003 (N_9003,N_7182,N_6010);
and U9004 (N_9004,N_7013,N_5581);
xor U9005 (N_9005,N_5687,N_5959);
nand U9006 (N_9006,N_5433,N_6503);
nor U9007 (N_9007,N_7496,N_7049);
xor U9008 (N_9008,N_5013,N_6671);
nor U9009 (N_9009,N_5539,N_5376);
or U9010 (N_9010,N_6592,N_6997);
nand U9011 (N_9011,N_7413,N_6695);
and U9012 (N_9012,N_6322,N_6416);
and U9013 (N_9013,N_6305,N_5421);
nor U9014 (N_9014,N_5459,N_5148);
and U9015 (N_9015,N_5162,N_6433);
xnor U9016 (N_9016,N_5037,N_7127);
nor U9017 (N_9017,N_6066,N_5320);
xor U9018 (N_9018,N_5578,N_5336);
or U9019 (N_9019,N_5246,N_5533);
nand U9020 (N_9020,N_7378,N_6738);
or U9021 (N_9021,N_5010,N_5219);
nand U9022 (N_9022,N_6448,N_6170);
and U9023 (N_9023,N_5749,N_5861);
or U9024 (N_9024,N_6197,N_6942);
nand U9025 (N_9025,N_7473,N_5167);
or U9026 (N_9026,N_7437,N_7423);
nor U9027 (N_9027,N_6622,N_7377);
and U9028 (N_9028,N_5876,N_5772);
and U9029 (N_9029,N_5376,N_6848);
or U9030 (N_9030,N_5065,N_5914);
and U9031 (N_9031,N_6592,N_5734);
nor U9032 (N_9032,N_6441,N_5269);
or U9033 (N_9033,N_6860,N_5250);
xnor U9034 (N_9034,N_7121,N_5680);
and U9035 (N_9035,N_6604,N_6154);
or U9036 (N_9036,N_5482,N_6031);
and U9037 (N_9037,N_5717,N_5231);
nand U9038 (N_9038,N_6396,N_5732);
or U9039 (N_9039,N_5617,N_5414);
xnor U9040 (N_9040,N_6794,N_6418);
or U9041 (N_9041,N_5225,N_5889);
and U9042 (N_9042,N_6904,N_6798);
and U9043 (N_9043,N_7082,N_6728);
nor U9044 (N_9044,N_7268,N_6420);
nor U9045 (N_9045,N_5163,N_7468);
and U9046 (N_9046,N_5744,N_6230);
or U9047 (N_9047,N_5177,N_6871);
nor U9048 (N_9048,N_5595,N_5113);
nor U9049 (N_9049,N_6307,N_6638);
and U9050 (N_9050,N_5542,N_6748);
nor U9051 (N_9051,N_5841,N_7426);
or U9052 (N_9052,N_7006,N_6807);
nor U9053 (N_9053,N_5845,N_7280);
and U9054 (N_9054,N_5874,N_6692);
xor U9055 (N_9055,N_6548,N_5577);
nand U9056 (N_9056,N_6137,N_6044);
or U9057 (N_9057,N_6453,N_5204);
and U9058 (N_9058,N_7197,N_5245);
nor U9059 (N_9059,N_5434,N_5090);
nand U9060 (N_9060,N_5727,N_7461);
xor U9061 (N_9061,N_5921,N_5409);
and U9062 (N_9062,N_5449,N_6880);
and U9063 (N_9063,N_5663,N_5798);
xnor U9064 (N_9064,N_5110,N_5709);
nand U9065 (N_9065,N_6419,N_5077);
and U9066 (N_9066,N_5831,N_5815);
or U9067 (N_9067,N_7336,N_5775);
nor U9068 (N_9068,N_5580,N_6249);
nor U9069 (N_9069,N_5855,N_7431);
nor U9070 (N_9070,N_5007,N_5224);
or U9071 (N_9071,N_5299,N_6174);
or U9072 (N_9072,N_7265,N_7332);
nand U9073 (N_9073,N_5585,N_5659);
nand U9074 (N_9074,N_5096,N_6617);
or U9075 (N_9075,N_5908,N_7279);
nand U9076 (N_9076,N_6689,N_7497);
nor U9077 (N_9077,N_6954,N_5948);
nor U9078 (N_9078,N_5879,N_5089);
and U9079 (N_9079,N_6412,N_6756);
nor U9080 (N_9080,N_5558,N_6333);
xnor U9081 (N_9081,N_5578,N_6498);
xnor U9082 (N_9082,N_5770,N_7284);
nor U9083 (N_9083,N_7000,N_6356);
nor U9084 (N_9084,N_6720,N_5452);
or U9085 (N_9085,N_5081,N_5241);
xor U9086 (N_9086,N_5487,N_6401);
xnor U9087 (N_9087,N_7108,N_5103);
nand U9088 (N_9088,N_6006,N_5051);
or U9089 (N_9089,N_5733,N_6761);
nand U9090 (N_9090,N_6827,N_6211);
xor U9091 (N_9091,N_6675,N_7363);
nor U9092 (N_9092,N_5099,N_5671);
xor U9093 (N_9093,N_6643,N_6487);
or U9094 (N_9094,N_7455,N_6642);
or U9095 (N_9095,N_5745,N_5119);
nand U9096 (N_9096,N_6466,N_7377);
or U9097 (N_9097,N_6491,N_5195);
nor U9098 (N_9098,N_5030,N_7475);
and U9099 (N_9099,N_7105,N_5616);
nand U9100 (N_9100,N_6234,N_6851);
or U9101 (N_9101,N_5812,N_7093);
or U9102 (N_9102,N_6588,N_6718);
or U9103 (N_9103,N_6434,N_5896);
or U9104 (N_9104,N_5154,N_5183);
and U9105 (N_9105,N_7234,N_5564);
and U9106 (N_9106,N_5172,N_7233);
or U9107 (N_9107,N_6457,N_6108);
xor U9108 (N_9108,N_5250,N_7352);
nor U9109 (N_9109,N_7217,N_7232);
and U9110 (N_9110,N_7459,N_5841);
nand U9111 (N_9111,N_6101,N_6693);
xor U9112 (N_9112,N_6522,N_5229);
xor U9113 (N_9113,N_5328,N_5329);
or U9114 (N_9114,N_5349,N_6267);
nor U9115 (N_9115,N_6450,N_6093);
and U9116 (N_9116,N_6809,N_6386);
and U9117 (N_9117,N_5842,N_7477);
or U9118 (N_9118,N_7477,N_7419);
nand U9119 (N_9119,N_5529,N_6627);
xor U9120 (N_9120,N_6695,N_6139);
or U9121 (N_9121,N_7129,N_5247);
nor U9122 (N_9122,N_5089,N_6711);
nor U9123 (N_9123,N_6686,N_6772);
xnor U9124 (N_9124,N_5613,N_5294);
and U9125 (N_9125,N_5878,N_5704);
nand U9126 (N_9126,N_5092,N_5235);
and U9127 (N_9127,N_7183,N_7393);
or U9128 (N_9128,N_6765,N_6909);
nand U9129 (N_9129,N_6756,N_5951);
nand U9130 (N_9130,N_5714,N_6459);
nand U9131 (N_9131,N_6089,N_7417);
nor U9132 (N_9132,N_7111,N_6660);
nor U9133 (N_9133,N_5925,N_5384);
xor U9134 (N_9134,N_5953,N_6232);
xor U9135 (N_9135,N_6857,N_5645);
nor U9136 (N_9136,N_6220,N_7253);
xor U9137 (N_9137,N_5048,N_5902);
and U9138 (N_9138,N_5662,N_7071);
nand U9139 (N_9139,N_5287,N_6840);
nand U9140 (N_9140,N_6533,N_5786);
nor U9141 (N_9141,N_7256,N_6681);
nand U9142 (N_9142,N_5476,N_7477);
and U9143 (N_9143,N_7457,N_6458);
nor U9144 (N_9144,N_5416,N_6795);
and U9145 (N_9145,N_5932,N_6750);
xor U9146 (N_9146,N_6511,N_5776);
nor U9147 (N_9147,N_6139,N_5316);
xnor U9148 (N_9148,N_6945,N_7259);
or U9149 (N_9149,N_5840,N_6995);
nor U9150 (N_9150,N_6743,N_7237);
nor U9151 (N_9151,N_5034,N_5115);
nor U9152 (N_9152,N_6631,N_5651);
nor U9153 (N_9153,N_6569,N_7373);
or U9154 (N_9154,N_5877,N_6485);
nor U9155 (N_9155,N_7174,N_7291);
or U9156 (N_9156,N_6658,N_7470);
and U9157 (N_9157,N_7359,N_5804);
nor U9158 (N_9158,N_5565,N_7201);
nand U9159 (N_9159,N_5358,N_6834);
or U9160 (N_9160,N_7140,N_5121);
or U9161 (N_9161,N_5206,N_6326);
nor U9162 (N_9162,N_5535,N_6323);
nor U9163 (N_9163,N_6055,N_7446);
nor U9164 (N_9164,N_6745,N_7116);
nor U9165 (N_9165,N_6991,N_7250);
or U9166 (N_9166,N_6488,N_7067);
or U9167 (N_9167,N_6880,N_5057);
and U9168 (N_9168,N_6590,N_6572);
and U9169 (N_9169,N_5395,N_6751);
and U9170 (N_9170,N_5209,N_5806);
or U9171 (N_9171,N_5281,N_6353);
or U9172 (N_9172,N_5345,N_5497);
and U9173 (N_9173,N_6505,N_6875);
xnor U9174 (N_9174,N_5714,N_5718);
nand U9175 (N_9175,N_7211,N_5513);
or U9176 (N_9176,N_7489,N_5412);
and U9177 (N_9177,N_6858,N_5849);
and U9178 (N_9178,N_5878,N_7413);
and U9179 (N_9179,N_5560,N_5675);
and U9180 (N_9180,N_6927,N_7179);
xnor U9181 (N_9181,N_5406,N_5493);
nand U9182 (N_9182,N_6550,N_6116);
and U9183 (N_9183,N_6241,N_5220);
nand U9184 (N_9184,N_6421,N_7470);
and U9185 (N_9185,N_6812,N_6895);
and U9186 (N_9186,N_7297,N_5711);
and U9187 (N_9187,N_6979,N_6071);
xor U9188 (N_9188,N_6981,N_6628);
nand U9189 (N_9189,N_6317,N_6421);
and U9190 (N_9190,N_7191,N_6886);
nor U9191 (N_9191,N_7008,N_6328);
or U9192 (N_9192,N_5039,N_6979);
or U9193 (N_9193,N_6642,N_6622);
or U9194 (N_9194,N_7210,N_7002);
and U9195 (N_9195,N_6432,N_5805);
or U9196 (N_9196,N_5946,N_6853);
nand U9197 (N_9197,N_7350,N_5571);
or U9198 (N_9198,N_6899,N_6695);
and U9199 (N_9199,N_7114,N_7250);
or U9200 (N_9200,N_6488,N_6476);
xnor U9201 (N_9201,N_6392,N_6985);
or U9202 (N_9202,N_6455,N_7487);
xnor U9203 (N_9203,N_7475,N_7173);
nor U9204 (N_9204,N_6690,N_5537);
xnor U9205 (N_9205,N_7399,N_6936);
and U9206 (N_9206,N_7486,N_5597);
xnor U9207 (N_9207,N_5084,N_6657);
nor U9208 (N_9208,N_5195,N_5892);
or U9209 (N_9209,N_6959,N_6140);
and U9210 (N_9210,N_5202,N_5058);
xnor U9211 (N_9211,N_7215,N_5598);
or U9212 (N_9212,N_6438,N_6274);
or U9213 (N_9213,N_7477,N_6775);
nand U9214 (N_9214,N_6867,N_5204);
xor U9215 (N_9215,N_6164,N_5453);
nand U9216 (N_9216,N_6520,N_6226);
nor U9217 (N_9217,N_6695,N_5645);
nand U9218 (N_9218,N_7418,N_5685);
or U9219 (N_9219,N_7310,N_5948);
nor U9220 (N_9220,N_7074,N_5883);
and U9221 (N_9221,N_7177,N_6247);
nand U9222 (N_9222,N_5715,N_5634);
or U9223 (N_9223,N_7021,N_6128);
and U9224 (N_9224,N_6423,N_6334);
nand U9225 (N_9225,N_7179,N_5097);
nand U9226 (N_9226,N_6519,N_6932);
and U9227 (N_9227,N_5219,N_5006);
nand U9228 (N_9228,N_6124,N_6212);
nor U9229 (N_9229,N_6632,N_5785);
nor U9230 (N_9230,N_6670,N_6932);
nand U9231 (N_9231,N_6733,N_7191);
or U9232 (N_9232,N_6184,N_5975);
xnor U9233 (N_9233,N_5065,N_5493);
or U9234 (N_9234,N_7441,N_7181);
and U9235 (N_9235,N_7272,N_6743);
or U9236 (N_9236,N_7369,N_5982);
nand U9237 (N_9237,N_5756,N_5915);
nor U9238 (N_9238,N_5304,N_5018);
xor U9239 (N_9239,N_6189,N_7369);
or U9240 (N_9240,N_6510,N_5298);
or U9241 (N_9241,N_5392,N_6654);
nor U9242 (N_9242,N_7211,N_6891);
xor U9243 (N_9243,N_6167,N_7371);
or U9244 (N_9244,N_6315,N_6855);
xnor U9245 (N_9245,N_5575,N_5073);
nor U9246 (N_9246,N_7442,N_5668);
nor U9247 (N_9247,N_5435,N_5501);
xor U9248 (N_9248,N_5580,N_5067);
nand U9249 (N_9249,N_6444,N_5949);
nor U9250 (N_9250,N_6848,N_7147);
nor U9251 (N_9251,N_7077,N_7321);
nor U9252 (N_9252,N_7407,N_5846);
and U9253 (N_9253,N_6897,N_5232);
nor U9254 (N_9254,N_6195,N_5872);
and U9255 (N_9255,N_6546,N_5386);
nor U9256 (N_9256,N_6809,N_6017);
nand U9257 (N_9257,N_7047,N_5454);
and U9258 (N_9258,N_5133,N_6118);
nor U9259 (N_9259,N_7204,N_5797);
nand U9260 (N_9260,N_7154,N_7238);
nor U9261 (N_9261,N_7477,N_7227);
nand U9262 (N_9262,N_6341,N_5660);
nand U9263 (N_9263,N_5988,N_7276);
xor U9264 (N_9264,N_6898,N_5653);
and U9265 (N_9265,N_6446,N_5204);
xnor U9266 (N_9266,N_5165,N_7076);
nor U9267 (N_9267,N_5760,N_6204);
xnor U9268 (N_9268,N_6293,N_6648);
nor U9269 (N_9269,N_5293,N_7268);
or U9270 (N_9270,N_6491,N_5109);
and U9271 (N_9271,N_5154,N_6405);
nor U9272 (N_9272,N_6830,N_5869);
and U9273 (N_9273,N_5448,N_5358);
nand U9274 (N_9274,N_7483,N_5241);
nor U9275 (N_9275,N_6330,N_5638);
or U9276 (N_9276,N_7077,N_6070);
nor U9277 (N_9277,N_5568,N_6951);
xor U9278 (N_9278,N_6467,N_5090);
or U9279 (N_9279,N_7296,N_5802);
xor U9280 (N_9280,N_7396,N_5186);
xor U9281 (N_9281,N_7327,N_6866);
and U9282 (N_9282,N_7371,N_7294);
nor U9283 (N_9283,N_6186,N_6585);
nor U9284 (N_9284,N_6813,N_5768);
nand U9285 (N_9285,N_6599,N_7105);
and U9286 (N_9286,N_5455,N_6690);
xnor U9287 (N_9287,N_6859,N_5044);
xnor U9288 (N_9288,N_5324,N_6768);
xor U9289 (N_9289,N_6488,N_7283);
and U9290 (N_9290,N_5295,N_7262);
and U9291 (N_9291,N_5350,N_6068);
or U9292 (N_9292,N_7373,N_6915);
and U9293 (N_9293,N_6852,N_6847);
xor U9294 (N_9294,N_6906,N_6328);
or U9295 (N_9295,N_7401,N_6497);
or U9296 (N_9296,N_5929,N_7008);
xnor U9297 (N_9297,N_7207,N_6083);
nand U9298 (N_9298,N_6949,N_7008);
nand U9299 (N_9299,N_5936,N_6910);
xor U9300 (N_9300,N_6554,N_7348);
nand U9301 (N_9301,N_6603,N_5400);
or U9302 (N_9302,N_5592,N_6709);
xor U9303 (N_9303,N_5124,N_6893);
nand U9304 (N_9304,N_6974,N_7211);
xor U9305 (N_9305,N_5822,N_6379);
and U9306 (N_9306,N_5161,N_6908);
nand U9307 (N_9307,N_6580,N_7090);
and U9308 (N_9308,N_5933,N_6934);
nand U9309 (N_9309,N_6005,N_5026);
nand U9310 (N_9310,N_5915,N_5396);
xnor U9311 (N_9311,N_6273,N_6042);
nor U9312 (N_9312,N_7309,N_7255);
nand U9313 (N_9313,N_5428,N_6164);
and U9314 (N_9314,N_6282,N_5817);
nand U9315 (N_9315,N_5544,N_5117);
nand U9316 (N_9316,N_6972,N_5463);
nand U9317 (N_9317,N_5596,N_6721);
and U9318 (N_9318,N_5497,N_7460);
nor U9319 (N_9319,N_7321,N_5278);
nand U9320 (N_9320,N_5468,N_5242);
and U9321 (N_9321,N_6569,N_5309);
nor U9322 (N_9322,N_6973,N_6495);
xor U9323 (N_9323,N_6843,N_7078);
and U9324 (N_9324,N_6642,N_7211);
nor U9325 (N_9325,N_5725,N_7179);
xor U9326 (N_9326,N_7472,N_6818);
and U9327 (N_9327,N_6475,N_5853);
or U9328 (N_9328,N_6187,N_7346);
or U9329 (N_9329,N_6800,N_7254);
xnor U9330 (N_9330,N_6939,N_6226);
and U9331 (N_9331,N_6976,N_5890);
nor U9332 (N_9332,N_5830,N_7148);
nor U9333 (N_9333,N_7028,N_7247);
nand U9334 (N_9334,N_5118,N_7340);
xor U9335 (N_9335,N_5256,N_7212);
or U9336 (N_9336,N_5218,N_6059);
or U9337 (N_9337,N_5942,N_6784);
nand U9338 (N_9338,N_6379,N_6796);
xor U9339 (N_9339,N_5658,N_6701);
and U9340 (N_9340,N_5369,N_5732);
or U9341 (N_9341,N_5505,N_6948);
nand U9342 (N_9342,N_6152,N_6133);
nor U9343 (N_9343,N_6716,N_5911);
or U9344 (N_9344,N_6050,N_5713);
and U9345 (N_9345,N_5416,N_6060);
nor U9346 (N_9346,N_5739,N_5370);
xnor U9347 (N_9347,N_6479,N_5429);
nand U9348 (N_9348,N_5498,N_5016);
nand U9349 (N_9349,N_5018,N_5971);
nand U9350 (N_9350,N_5766,N_7353);
nand U9351 (N_9351,N_6695,N_7331);
xnor U9352 (N_9352,N_6237,N_6949);
nand U9353 (N_9353,N_6326,N_6358);
nor U9354 (N_9354,N_5848,N_6653);
and U9355 (N_9355,N_6852,N_5133);
or U9356 (N_9356,N_6044,N_7434);
and U9357 (N_9357,N_5176,N_6295);
or U9358 (N_9358,N_7078,N_5795);
xor U9359 (N_9359,N_5701,N_5398);
xor U9360 (N_9360,N_6959,N_6746);
nor U9361 (N_9361,N_6573,N_7011);
nor U9362 (N_9362,N_5235,N_5183);
or U9363 (N_9363,N_5640,N_7184);
and U9364 (N_9364,N_7274,N_6538);
nand U9365 (N_9365,N_6887,N_5289);
nand U9366 (N_9366,N_6531,N_5915);
nand U9367 (N_9367,N_7394,N_5133);
nand U9368 (N_9368,N_6706,N_6160);
nor U9369 (N_9369,N_7017,N_6619);
and U9370 (N_9370,N_6696,N_6319);
nand U9371 (N_9371,N_6182,N_5690);
nor U9372 (N_9372,N_6566,N_6941);
xor U9373 (N_9373,N_5798,N_5032);
and U9374 (N_9374,N_5277,N_6922);
nand U9375 (N_9375,N_6501,N_7240);
nand U9376 (N_9376,N_5539,N_6105);
and U9377 (N_9377,N_7063,N_6826);
and U9378 (N_9378,N_5261,N_5371);
or U9379 (N_9379,N_5290,N_5269);
and U9380 (N_9380,N_5226,N_7258);
nor U9381 (N_9381,N_5841,N_5822);
or U9382 (N_9382,N_5147,N_7397);
nor U9383 (N_9383,N_5926,N_7418);
or U9384 (N_9384,N_5329,N_6057);
and U9385 (N_9385,N_5660,N_5696);
and U9386 (N_9386,N_6249,N_6685);
or U9387 (N_9387,N_6282,N_6271);
or U9388 (N_9388,N_5590,N_5526);
xnor U9389 (N_9389,N_6487,N_6765);
nand U9390 (N_9390,N_5383,N_6788);
nand U9391 (N_9391,N_7396,N_6136);
and U9392 (N_9392,N_7271,N_5738);
xor U9393 (N_9393,N_6655,N_6749);
xnor U9394 (N_9394,N_5333,N_5558);
xnor U9395 (N_9395,N_7136,N_6781);
and U9396 (N_9396,N_6354,N_5165);
nand U9397 (N_9397,N_5382,N_5559);
nand U9398 (N_9398,N_7368,N_7048);
or U9399 (N_9399,N_5058,N_7215);
nor U9400 (N_9400,N_6813,N_6304);
nand U9401 (N_9401,N_5637,N_6369);
or U9402 (N_9402,N_7391,N_6921);
xnor U9403 (N_9403,N_7088,N_5271);
nor U9404 (N_9404,N_6222,N_6298);
or U9405 (N_9405,N_7468,N_7089);
nor U9406 (N_9406,N_5959,N_6286);
xor U9407 (N_9407,N_5048,N_7090);
or U9408 (N_9408,N_5901,N_7432);
xor U9409 (N_9409,N_5088,N_5620);
and U9410 (N_9410,N_5171,N_6452);
or U9411 (N_9411,N_7107,N_6370);
or U9412 (N_9412,N_5814,N_6776);
nor U9413 (N_9413,N_5827,N_5567);
or U9414 (N_9414,N_7277,N_7102);
nand U9415 (N_9415,N_6350,N_7469);
xnor U9416 (N_9416,N_7232,N_6809);
or U9417 (N_9417,N_6957,N_5247);
xor U9418 (N_9418,N_5801,N_5101);
nor U9419 (N_9419,N_5261,N_7263);
nor U9420 (N_9420,N_5402,N_6289);
xor U9421 (N_9421,N_6767,N_7037);
and U9422 (N_9422,N_5622,N_5807);
or U9423 (N_9423,N_6612,N_6683);
nand U9424 (N_9424,N_7082,N_7038);
and U9425 (N_9425,N_5919,N_5949);
xnor U9426 (N_9426,N_6611,N_5348);
xnor U9427 (N_9427,N_7236,N_5948);
xor U9428 (N_9428,N_5703,N_6540);
and U9429 (N_9429,N_6065,N_5501);
or U9430 (N_9430,N_5221,N_6599);
nand U9431 (N_9431,N_5444,N_7200);
nor U9432 (N_9432,N_5100,N_5993);
or U9433 (N_9433,N_6886,N_6796);
nand U9434 (N_9434,N_5342,N_5876);
and U9435 (N_9435,N_5339,N_6733);
nor U9436 (N_9436,N_7197,N_6306);
or U9437 (N_9437,N_5191,N_6680);
and U9438 (N_9438,N_6841,N_7275);
nor U9439 (N_9439,N_5550,N_7359);
and U9440 (N_9440,N_6939,N_6648);
xor U9441 (N_9441,N_6097,N_6814);
or U9442 (N_9442,N_7328,N_7050);
nand U9443 (N_9443,N_6662,N_6108);
xor U9444 (N_9444,N_6256,N_5677);
and U9445 (N_9445,N_5626,N_5075);
or U9446 (N_9446,N_5907,N_5615);
nand U9447 (N_9447,N_6603,N_5358);
nor U9448 (N_9448,N_6211,N_6605);
xor U9449 (N_9449,N_5079,N_5908);
nor U9450 (N_9450,N_6384,N_6967);
or U9451 (N_9451,N_5526,N_7021);
xor U9452 (N_9452,N_5154,N_6334);
xor U9453 (N_9453,N_5697,N_6382);
nand U9454 (N_9454,N_6380,N_6995);
or U9455 (N_9455,N_5259,N_6393);
nand U9456 (N_9456,N_6753,N_7256);
nor U9457 (N_9457,N_5832,N_5904);
xor U9458 (N_9458,N_7047,N_5565);
or U9459 (N_9459,N_5260,N_5000);
xor U9460 (N_9460,N_7389,N_5312);
nor U9461 (N_9461,N_5809,N_6010);
nor U9462 (N_9462,N_5776,N_6506);
nor U9463 (N_9463,N_7403,N_7119);
nand U9464 (N_9464,N_5023,N_6085);
and U9465 (N_9465,N_5443,N_6775);
or U9466 (N_9466,N_6641,N_5834);
or U9467 (N_9467,N_7034,N_6889);
xnor U9468 (N_9468,N_5763,N_5124);
nor U9469 (N_9469,N_6201,N_6775);
nor U9470 (N_9470,N_5930,N_7079);
nand U9471 (N_9471,N_7352,N_6886);
nor U9472 (N_9472,N_6916,N_5009);
nand U9473 (N_9473,N_5106,N_5023);
or U9474 (N_9474,N_5212,N_6659);
and U9475 (N_9475,N_7311,N_5535);
xnor U9476 (N_9476,N_5917,N_5696);
nor U9477 (N_9477,N_7461,N_5587);
xor U9478 (N_9478,N_6163,N_7438);
and U9479 (N_9479,N_7393,N_6339);
xnor U9480 (N_9480,N_5632,N_6033);
and U9481 (N_9481,N_5816,N_6485);
or U9482 (N_9482,N_5679,N_6218);
xnor U9483 (N_9483,N_6152,N_5889);
xor U9484 (N_9484,N_5281,N_5450);
or U9485 (N_9485,N_7183,N_5000);
or U9486 (N_9486,N_5793,N_6482);
nand U9487 (N_9487,N_6328,N_7090);
xnor U9488 (N_9488,N_5393,N_6593);
nand U9489 (N_9489,N_5834,N_5815);
or U9490 (N_9490,N_6105,N_6396);
and U9491 (N_9491,N_5129,N_7347);
nor U9492 (N_9492,N_7289,N_5330);
xor U9493 (N_9493,N_5743,N_6736);
nor U9494 (N_9494,N_5374,N_5302);
nand U9495 (N_9495,N_7075,N_6884);
and U9496 (N_9496,N_6160,N_7484);
xnor U9497 (N_9497,N_5056,N_6842);
xor U9498 (N_9498,N_6020,N_5817);
or U9499 (N_9499,N_7494,N_5951);
or U9500 (N_9500,N_6166,N_6433);
xor U9501 (N_9501,N_5932,N_7030);
and U9502 (N_9502,N_5043,N_5445);
nand U9503 (N_9503,N_6045,N_7195);
xnor U9504 (N_9504,N_5298,N_5374);
nand U9505 (N_9505,N_5969,N_6751);
nor U9506 (N_9506,N_6864,N_6854);
xor U9507 (N_9507,N_5765,N_5784);
and U9508 (N_9508,N_6591,N_7151);
nand U9509 (N_9509,N_6457,N_5202);
or U9510 (N_9510,N_5460,N_6428);
and U9511 (N_9511,N_5368,N_7443);
xnor U9512 (N_9512,N_6324,N_6466);
nor U9513 (N_9513,N_7374,N_6726);
nand U9514 (N_9514,N_6667,N_5785);
xnor U9515 (N_9515,N_6643,N_7460);
nand U9516 (N_9516,N_6466,N_6520);
or U9517 (N_9517,N_6756,N_6757);
and U9518 (N_9518,N_5416,N_5052);
nor U9519 (N_9519,N_7483,N_6018);
and U9520 (N_9520,N_6654,N_5428);
nor U9521 (N_9521,N_6431,N_6591);
xor U9522 (N_9522,N_7278,N_6146);
or U9523 (N_9523,N_6111,N_5511);
nor U9524 (N_9524,N_6078,N_6905);
nor U9525 (N_9525,N_6418,N_5212);
xnor U9526 (N_9526,N_6251,N_5451);
xnor U9527 (N_9527,N_5037,N_6935);
xnor U9528 (N_9528,N_7092,N_5038);
nor U9529 (N_9529,N_6689,N_6113);
nand U9530 (N_9530,N_7338,N_5834);
and U9531 (N_9531,N_5627,N_5184);
and U9532 (N_9532,N_5075,N_6044);
xnor U9533 (N_9533,N_5145,N_6835);
or U9534 (N_9534,N_7016,N_6349);
xor U9535 (N_9535,N_6667,N_6725);
and U9536 (N_9536,N_6066,N_5815);
xor U9537 (N_9537,N_5748,N_6516);
or U9538 (N_9538,N_6000,N_5384);
or U9539 (N_9539,N_6317,N_5747);
xnor U9540 (N_9540,N_5358,N_5824);
nand U9541 (N_9541,N_7187,N_6655);
and U9542 (N_9542,N_7209,N_6681);
or U9543 (N_9543,N_6044,N_6110);
or U9544 (N_9544,N_6231,N_5955);
and U9545 (N_9545,N_5410,N_6399);
and U9546 (N_9546,N_6428,N_5074);
and U9547 (N_9547,N_5407,N_5492);
nand U9548 (N_9548,N_7465,N_5554);
and U9549 (N_9549,N_5924,N_7221);
nand U9550 (N_9550,N_5801,N_5811);
xnor U9551 (N_9551,N_7362,N_6017);
nor U9552 (N_9552,N_6777,N_6444);
or U9553 (N_9553,N_6479,N_5764);
nor U9554 (N_9554,N_6862,N_5249);
and U9555 (N_9555,N_6632,N_6424);
xnor U9556 (N_9556,N_7417,N_6321);
xnor U9557 (N_9557,N_5801,N_5580);
and U9558 (N_9558,N_7315,N_5073);
and U9559 (N_9559,N_6905,N_7054);
nand U9560 (N_9560,N_6193,N_5773);
or U9561 (N_9561,N_7168,N_5771);
and U9562 (N_9562,N_5903,N_6974);
and U9563 (N_9563,N_6624,N_5611);
and U9564 (N_9564,N_5955,N_6566);
nand U9565 (N_9565,N_7331,N_7158);
and U9566 (N_9566,N_6930,N_5380);
nor U9567 (N_9567,N_6910,N_5491);
xnor U9568 (N_9568,N_5749,N_6041);
xnor U9569 (N_9569,N_5295,N_7119);
xnor U9570 (N_9570,N_5446,N_6686);
nand U9571 (N_9571,N_5066,N_5540);
xor U9572 (N_9572,N_6718,N_5310);
and U9573 (N_9573,N_7384,N_7034);
xor U9574 (N_9574,N_7296,N_5188);
xor U9575 (N_9575,N_7336,N_7432);
nand U9576 (N_9576,N_5942,N_5803);
xor U9577 (N_9577,N_6641,N_5700);
xor U9578 (N_9578,N_7260,N_6499);
or U9579 (N_9579,N_7265,N_7481);
nor U9580 (N_9580,N_6669,N_5962);
xnor U9581 (N_9581,N_7079,N_6165);
nand U9582 (N_9582,N_5229,N_5219);
nand U9583 (N_9583,N_5162,N_5493);
or U9584 (N_9584,N_5552,N_5594);
and U9585 (N_9585,N_6106,N_7461);
xor U9586 (N_9586,N_5765,N_7173);
xnor U9587 (N_9587,N_6852,N_5122);
and U9588 (N_9588,N_6066,N_5089);
nor U9589 (N_9589,N_5024,N_6952);
xor U9590 (N_9590,N_6506,N_7495);
xnor U9591 (N_9591,N_6273,N_5733);
and U9592 (N_9592,N_7391,N_6535);
and U9593 (N_9593,N_7479,N_5127);
or U9594 (N_9594,N_7468,N_6853);
xnor U9595 (N_9595,N_7391,N_6008);
nor U9596 (N_9596,N_6109,N_5392);
and U9597 (N_9597,N_6837,N_5882);
nor U9598 (N_9598,N_6012,N_5804);
xnor U9599 (N_9599,N_5047,N_6034);
xnor U9600 (N_9600,N_5705,N_6653);
or U9601 (N_9601,N_5820,N_5339);
and U9602 (N_9602,N_5686,N_7418);
xor U9603 (N_9603,N_6535,N_5280);
xnor U9604 (N_9604,N_7130,N_7470);
nand U9605 (N_9605,N_6407,N_6065);
or U9606 (N_9606,N_5026,N_7169);
nor U9607 (N_9607,N_6357,N_7198);
and U9608 (N_9608,N_5993,N_6564);
nand U9609 (N_9609,N_5364,N_5927);
and U9610 (N_9610,N_6051,N_5817);
nand U9611 (N_9611,N_6965,N_6379);
or U9612 (N_9612,N_7197,N_7209);
nor U9613 (N_9613,N_5714,N_6470);
or U9614 (N_9614,N_5840,N_7120);
or U9615 (N_9615,N_6938,N_5921);
and U9616 (N_9616,N_5561,N_6770);
nor U9617 (N_9617,N_6438,N_6208);
xor U9618 (N_9618,N_7068,N_6856);
nand U9619 (N_9619,N_7136,N_5335);
xnor U9620 (N_9620,N_7084,N_6605);
or U9621 (N_9621,N_5902,N_5539);
xor U9622 (N_9622,N_6905,N_5162);
and U9623 (N_9623,N_6891,N_7022);
or U9624 (N_9624,N_5341,N_6203);
and U9625 (N_9625,N_6560,N_5780);
xnor U9626 (N_9626,N_7165,N_5372);
nand U9627 (N_9627,N_5181,N_6395);
xnor U9628 (N_9628,N_6793,N_5084);
or U9629 (N_9629,N_5882,N_5343);
xor U9630 (N_9630,N_5142,N_6862);
nand U9631 (N_9631,N_5352,N_5430);
or U9632 (N_9632,N_5469,N_5643);
or U9633 (N_9633,N_5375,N_6186);
nand U9634 (N_9634,N_5929,N_5177);
or U9635 (N_9635,N_6952,N_5718);
or U9636 (N_9636,N_5737,N_5829);
nand U9637 (N_9637,N_5426,N_6629);
nand U9638 (N_9638,N_5820,N_6416);
and U9639 (N_9639,N_6041,N_5595);
or U9640 (N_9640,N_7492,N_5524);
nand U9641 (N_9641,N_5530,N_6802);
and U9642 (N_9642,N_7484,N_6606);
and U9643 (N_9643,N_5029,N_5415);
nor U9644 (N_9644,N_5189,N_5337);
nand U9645 (N_9645,N_7478,N_5810);
or U9646 (N_9646,N_7021,N_5533);
or U9647 (N_9647,N_5959,N_5783);
or U9648 (N_9648,N_5271,N_5910);
nor U9649 (N_9649,N_5181,N_6723);
nor U9650 (N_9650,N_7195,N_5899);
or U9651 (N_9651,N_5297,N_5616);
nand U9652 (N_9652,N_7331,N_5242);
or U9653 (N_9653,N_7341,N_7150);
nor U9654 (N_9654,N_6748,N_5700);
nor U9655 (N_9655,N_7086,N_6809);
nand U9656 (N_9656,N_6797,N_6410);
and U9657 (N_9657,N_5380,N_7465);
and U9658 (N_9658,N_5730,N_6750);
nand U9659 (N_9659,N_6058,N_5314);
xor U9660 (N_9660,N_5102,N_5471);
or U9661 (N_9661,N_6287,N_5264);
xnor U9662 (N_9662,N_6953,N_7447);
nand U9663 (N_9663,N_5160,N_6537);
xnor U9664 (N_9664,N_6248,N_6547);
nor U9665 (N_9665,N_5925,N_6084);
and U9666 (N_9666,N_5845,N_6911);
and U9667 (N_9667,N_5883,N_7363);
nor U9668 (N_9668,N_6840,N_5984);
nor U9669 (N_9669,N_5802,N_7493);
or U9670 (N_9670,N_6734,N_6071);
nand U9671 (N_9671,N_5763,N_6966);
xor U9672 (N_9672,N_6147,N_7236);
and U9673 (N_9673,N_5140,N_7106);
nand U9674 (N_9674,N_6734,N_5490);
nand U9675 (N_9675,N_7480,N_6641);
nand U9676 (N_9676,N_5663,N_5913);
and U9677 (N_9677,N_5968,N_6073);
nand U9678 (N_9678,N_6651,N_6378);
nor U9679 (N_9679,N_6720,N_5707);
or U9680 (N_9680,N_6421,N_6477);
xnor U9681 (N_9681,N_7151,N_6776);
or U9682 (N_9682,N_6608,N_7486);
nor U9683 (N_9683,N_5351,N_6419);
xor U9684 (N_9684,N_5933,N_5651);
or U9685 (N_9685,N_7307,N_7054);
and U9686 (N_9686,N_5829,N_7084);
nor U9687 (N_9687,N_5103,N_6899);
nand U9688 (N_9688,N_6225,N_6787);
nand U9689 (N_9689,N_7264,N_6983);
and U9690 (N_9690,N_6087,N_5059);
nor U9691 (N_9691,N_5555,N_6984);
nor U9692 (N_9692,N_6612,N_6959);
xor U9693 (N_9693,N_6402,N_6489);
xor U9694 (N_9694,N_5163,N_7305);
and U9695 (N_9695,N_5568,N_7053);
xor U9696 (N_9696,N_6468,N_5493);
xnor U9697 (N_9697,N_7148,N_6490);
nand U9698 (N_9698,N_5107,N_6565);
xor U9699 (N_9699,N_5786,N_6246);
or U9700 (N_9700,N_6359,N_7432);
nand U9701 (N_9701,N_5351,N_5098);
xnor U9702 (N_9702,N_5515,N_5478);
or U9703 (N_9703,N_5857,N_6438);
or U9704 (N_9704,N_7322,N_7078);
xnor U9705 (N_9705,N_5603,N_5894);
nor U9706 (N_9706,N_5983,N_7080);
and U9707 (N_9707,N_5431,N_5565);
or U9708 (N_9708,N_6371,N_6534);
and U9709 (N_9709,N_5887,N_6686);
or U9710 (N_9710,N_6954,N_7426);
nor U9711 (N_9711,N_6535,N_5872);
nand U9712 (N_9712,N_5296,N_6087);
or U9713 (N_9713,N_5609,N_5031);
nand U9714 (N_9714,N_7373,N_6941);
or U9715 (N_9715,N_5545,N_5379);
xor U9716 (N_9716,N_5008,N_7037);
or U9717 (N_9717,N_6169,N_6789);
or U9718 (N_9718,N_5067,N_7025);
nor U9719 (N_9719,N_6095,N_6314);
nor U9720 (N_9720,N_6188,N_5761);
or U9721 (N_9721,N_6138,N_5384);
nand U9722 (N_9722,N_6737,N_6753);
xnor U9723 (N_9723,N_5065,N_5126);
nand U9724 (N_9724,N_7300,N_6819);
xor U9725 (N_9725,N_7027,N_7065);
or U9726 (N_9726,N_6118,N_6932);
xor U9727 (N_9727,N_6403,N_7283);
nor U9728 (N_9728,N_5310,N_6162);
nor U9729 (N_9729,N_5134,N_5657);
xor U9730 (N_9730,N_6724,N_7333);
and U9731 (N_9731,N_6245,N_5465);
nor U9732 (N_9732,N_6168,N_6626);
nor U9733 (N_9733,N_6932,N_7304);
nand U9734 (N_9734,N_6431,N_7010);
and U9735 (N_9735,N_5624,N_6020);
nand U9736 (N_9736,N_6103,N_5232);
and U9737 (N_9737,N_6831,N_7277);
nor U9738 (N_9738,N_6115,N_5654);
or U9739 (N_9739,N_5628,N_5663);
nor U9740 (N_9740,N_7472,N_6455);
or U9741 (N_9741,N_6797,N_5104);
xnor U9742 (N_9742,N_7127,N_5006);
nor U9743 (N_9743,N_5546,N_7386);
nor U9744 (N_9744,N_6211,N_7404);
nand U9745 (N_9745,N_6643,N_7368);
nor U9746 (N_9746,N_7402,N_5787);
nor U9747 (N_9747,N_5899,N_6771);
nor U9748 (N_9748,N_6956,N_6263);
xor U9749 (N_9749,N_7398,N_6018);
xnor U9750 (N_9750,N_6516,N_5106);
nand U9751 (N_9751,N_6865,N_7167);
or U9752 (N_9752,N_5070,N_6814);
nor U9753 (N_9753,N_5548,N_5283);
nand U9754 (N_9754,N_6953,N_7184);
or U9755 (N_9755,N_6761,N_6416);
nor U9756 (N_9756,N_6989,N_6379);
xnor U9757 (N_9757,N_5274,N_5522);
nor U9758 (N_9758,N_5614,N_5771);
and U9759 (N_9759,N_7266,N_7206);
nor U9760 (N_9760,N_5805,N_5974);
nor U9761 (N_9761,N_6031,N_5591);
and U9762 (N_9762,N_5243,N_7434);
and U9763 (N_9763,N_6906,N_6277);
nor U9764 (N_9764,N_7403,N_6522);
xor U9765 (N_9765,N_6385,N_5230);
nand U9766 (N_9766,N_6067,N_5278);
nand U9767 (N_9767,N_6710,N_5314);
nor U9768 (N_9768,N_7453,N_6455);
xor U9769 (N_9769,N_6937,N_5297);
nor U9770 (N_9770,N_6849,N_5298);
xnor U9771 (N_9771,N_7231,N_6988);
xor U9772 (N_9772,N_6524,N_6920);
or U9773 (N_9773,N_6269,N_6444);
and U9774 (N_9774,N_5808,N_5233);
nand U9775 (N_9775,N_5107,N_6651);
and U9776 (N_9776,N_5820,N_6342);
xor U9777 (N_9777,N_5249,N_6463);
nor U9778 (N_9778,N_7248,N_7471);
xnor U9779 (N_9779,N_5745,N_5146);
nand U9780 (N_9780,N_6055,N_5483);
nor U9781 (N_9781,N_5654,N_6659);
nor U9782 (N_9782,N_5599,N_5511);
and U9783 (N_9783,N_5585,N_5296);
and U9784 (N_9784,N_7066,N_6476);
nand U9785 (N_9785,N_5424,N_6478);
or U9786 (N_9786,N_6956,N_5593);
nand U9787 (N_9787,N_5870,N_7121);
nand U9788 (N_9788,N_5094,N_5477);
nor U9789 (N_9789,N_7367,N_7052);
xnor U9790 (N_9790,N_7294,N_6892);
or U9791 (N_9791,N_7222,N_6326);
nor U9792 (N_9792,N_7114,N_6478);
and U9793 (N_9793,N_5508,N_6808);
or U9794 (N_9794,N_7056,N_6580);
xnor U9795 (N_9795,N_6196,N_6280);
or U9796 (N_9796,N_6118,N_7135);
nand U9797 (N_9797,N_5376,N_6750);
or U9798 (N_9798,N_7410,N_6006);
and U9799 (N_9799,N_5477,N_5026);
or U9800 (N_9800,N_6268,N_6290);
nor U9801 (N_9801,N_6751,N_6856);
xnor U9802 (N_9802,N_6415,N_6733);
or U9803 (N_9803,N_6647,N_6234);
or U9804 (N_9804,N_6281,N_6330);
nand U9805 (N_9805,N_5536,N_7239);
nand U9806 (N_9806,N_6628,N_6119);
nand U9807 (N_9807,N_5770,N_5879);
or U9808 (N_9808,N_5962,N_5455);
nand U9809 (N_9809,N_7218,N_5385);
xnor U9810 (N_9810,N_7369,N_5287);
nand U9811 (N_9811,N_6463,N_5154);
and U9812 (N_9812,N_6502,N_6545);
or U9813 (N_9813,N_7399,N_5315);
nand U9814 (N_9814,N_5271,N_7369);
nand U9815 (N_9815,N_5441,N_6530);
xnor U9816 (N_9816,N_6082,N_6936);
and U9817 (N_9817,N_5272,N_5520);
nor U9818 (N_9818,N_6746,N_6174);
or U9819 (N_9819,N_5246,N_6873);
or U9820 (N_9820,N_5292,N_5035);
nand U9821 (N_9821,N_7083,N_7310);
or U9822 (N_9822,N_6142,N_6395);
nor U9823 (N_9823,N_6569,N_5715);
and U9824 (N_9824,N_6779,N_5201);
xnor U9825 (N_9825,N_5143,N_7023);
xnor U9826 (N_9826,N_5186,N_6356);
and U9827 (N_9827,N_7376,N_7295);
nor U9828 (N_9828,N_7123,N_6653);
xnor U9829 (N_9829,N_6262,N_7172);
or U9830 (N_9830,N_7485,N_6331);
nor U9831 (N_9831,N_7377,N_5712);
or U9832 (N_9832,N_5423,N_6744);
or U9833 (N_9833,N_6827,N_5761);
nand U9834 (N_9834,N_6902,N_5028);
and U9835 (N_9835,N_7092,N_5861);
and U9836 (N_9836,N_6178,N_6693);
xnor U9837 (N_9837,N_6225,N_6937);
nand U9838 (N_9838,N_5451,N_6692);
xor U9839 (N_9839,N_7224,N_6699);
xnor U9840 (N_9840,N_5697,N_5039);
or U9841 (N_9841,N_6681,N_5038);
nor U9842 (N_9842,N_5876,N_5072);
and U9843 (N_9843,N_7433,N_7064);
xnor U9844 (N_9844,N_6753,N_6666);
nand U9845 (N_9845,N_5656,N_5077);
or U9846 (N_9846,N_6824,N_5249);
nand U9847 (N_9847,N_7071,N_7427);
xor U9848 (N_9848,N_6254,N_6873);
and U9849 (N_9849,N_5368,N_6261);
and U9850 (N_9850,N_7375,N_6968);
nor U9851 (N_9851,N_5873,N_6286);
or U9852 (N_9852,N_7359,N_5859);
or U9853 (N_9853,N_6451,N_6638);
nand U9854 (N_9854,N_7233,N_6050);
nor U9855 (N_9855,N_5016,N_5051);
xnor U9856 (N_9856,N_5780,N_5307);
nor U9857 (N_9857,N_5489,N_5424);
and U9858 (N_9858,N_6576,N_5600);
xnor U9859 (N_9859,N_5578,N_5949);
xnor U9860 (N_9860,N_6633,N_5402);
xnor U9861 (N_9861,N_5397,N_5360);
or U9862 (N_9862,N_6373,N_5114);
and U9863 (N_9863,N_5719,N_7233);
and U9864 (N_9864,N_5411,N_7009);
or U9865 (N_9865,N_5878,N_5797);
xnor U9866 (N_9866,N_5036,N_5669);
nand U9867 (N_9867,N_5973,N_5150);
nand U9868 (N_9868,N_5721,N_7145);
or U9869 (N_9869,N_6790,N_5295);
and U9870 (N_9870,N_5805,N_6877);
nand U9871 (N_9871,N_6599,N_5674);
nand U9872 (N_9872,N_6827,N_5874);
nand U9873 (N_9873,N_5304,N_6083);
and U9874 (N_9874,N_7085,N_5708);
and U9875 (N_9875,N_6307,N_6590);
or U9876 (N_9876,N_6203,N_6735);
and U9877 (N_9877,N_6616,N_5146);
nand U9878 (N_9878,N_5321,N_7248);
or U9879 (N_9879,N_6514,N_6224);
or U9880 (N_9880,N_5587,N_5989);
nand U9881 (N_9881,N_7337,N_6163);
or U9882 (N_9882,N_6620,N_6539);
and U9883 (N_9883,N_7249,N_5107);
nor U9884 (N_9884,N_6325,N_6957);
and U9885 (N_9885,N_5554,N_5205);
and U9886 (N_9886,N_6256,N_5148);
or U9887 (N_9887,N_7164,N_5576);
xor U9888 (N_9888,N_5215,N_6194);
and U9889 (N_9889,N_5321,N_7068);
nand U9890 (N_9890,N_6643,N_6891);
or U9891 (N_9891,N_6505,N_7347);
nand U9892 (N_9892,N_6290,N_6839);
xnor U9893 (N_9893,N_7023,N_5569);
nor U9894 (N_9894,N_5774,N_6959);
and U9895 (N_9895,N_7245,N_5536);
xor U9896 (N_9896,N_5407,N_6366);
and U9897 (N_9897,N_7036,N_6827);
and U9898 (N_9898,N_5326,N_5530);
nand U9899 (N_9899,N_6627,N_5661);
and U9900 (N_9900,N_7045,N_5290);
or U9901 (N_9901,N_5138,N_5743);
xor U9902 (N_9902,N_5661,N_6040);
and U9903 (N_9903,N_6320,N_5380);
and U9904 (N_9904,N_7264,N_5695);
xnor U9905 (N_9905,N_7344,N_5147);
xnor U9906 (N_9906,N_7375,N_6253);
nand U9907 (N_9907,N_6942,N_7268);
or U9908 (N_9908,N_6442,N_6832);
xnor U9909 (N_9909,N_6811,N_6930);
and U9910 (N_9910,N_7484,N_5069);
nor U9911 (N_9911,N_5139,N_6844);
nor U9912 (N_9912,N_6867,N_6522);
and U9913 (N_9913,N_6736,N_5772);
nand U9914 (N_9914,N_5951,N_6363);
xnor U9915 (N_9915,N_5788,N_7130);
and U9916 (N_9916,N_6235,N_6495);
xor U9917 (N_9917,N_5332,N_6886);
xnor U9918 (N_9918,N_5906,N_5961);
nor U9919 (N_9919,N_5799,N_7084);
nor U9920 (N_9920,N_6657,N_5406);
nand U9921 (N_9921,N_6533,N_6940);
nor U9922 (N_9922,N_5137,N_6600);
and U9923 (N_9923,N_6604,N_6240);
or U9924 (N_9924,N_6152,N_6050);
xor U9925 (N_9925,N_6193,N_6409);
nor U9926 (N_9926,N_6492,N_6718);
or U9927 (N_9927,N_5461,N_6312);
nor U9928 (N_9928,N_6499,N_5437);
xor U9929 (N_9929,N_5960,N_6150);
nor U9930 (N_9930,N_7364,N_5741);
xor U9931 (N_9931,N_5723,N_6280);
nand U9932 (N_9932,N_6517,N_6986);
or U9933 (N_9933,N_6327,N_5031);
xnor U9934 (N_9934,N_5074,N_7484);
nand U9935 (N_9935,N_5743,N_5382);
or U9936 (N_9936,N_5681,N_6986);
xnor U9937 (N_9937,N_7495,N_6184);
nor U9938 (N_9938,N_7434,N_6448);
nand U9939 (N_9939,N_7272,N_5115);
and U9940 (N_9940,N_5544,N_5854);
or U9941 (N_9941,N_6974,N_5991);
nand U9942 (N_9942,N_5865,N_6133);
or U9943 (N_9943,N_5304,N_5878);
nor U9944 (N_9944,N_6589,N_6108);
nand U9945 (N_9945,N_6367,N_6230);
nor U9946 (N_9946,N_5362,N_5404);
or U9947 (N_9947,N_7387,N_6069);
nor U9948 (N_9948,N_5347,N_7133);
or U9949 (N_9949,N_5544,N_6068);
nor U9950 (N_9950,N_5943,N_5476);
or U9951 (N_9951,N_6721,N_6184);
nor U9952 (N_9952,N_5193,N_6560);
or U9953 (N_9953,N_7057,N_6947);
nor U9954 (N_9954,N_6811,N_7152);
nor U9955 (N_9955,N_6665,N_6562);
and U9956 (N_9956,N_5311,N_5898);
nor U9957 (N_9957,N_5404,N_6399);
nand U9958 (N_9958,N_5702,N_5053);
nor U9959 (N_9959,N_7040,N_5230);
or U9960 (N_9960,N_6315,N_5681);
nor U9961 (N_9961,N_5500,N_7405);
nand U9962 (N_9962,N_5392,N_6208);
and U9963 (N_9963,N_6865,N_5592);
or U9964 (N_9964,N_6343,N_5832);
or U9965 (N_9965,N_5767,N_5157);
nand U9966 (N_9966,N_6884,N_7436);
nor U9967 (N_9967,N_6436,N_5633);
xnor U9968 (N_9968,N_5853,N_5704);
nor U9969 (N_9969,N_5732,N_5011);
nor U9970 (N_9970,N_7051,N_6778);
or U9971 (N_9971,N_5311,N_5285);
nor U9972 (N_9972,N_7061,N_6355);
nand U9973 (N_9973,N_5843,N_6574);
nand U9974 (N_9974,N_5621,N_6992);
xnor U9975 (N_9975,N_5321,N_7060);
xor U9976 (N_9976,N_6840,N_5362);
and U9977 (N_9977,N_5774,N_5771);
and U9978 (N_9978,N_6106,N_6551);
and U9979 (N_9979,N_6292,N_5438);
xnor U9980 (N_9980,N_5764,N_6296);
and U9981 (N_9981,N_6324,N_6618);
and U9982 (N_9982,N_6119,N_7079);
nor U9983 (N_9983,N_5657,N_7380);
and U9984 (N_9984,N_6603,N_5604);
xnor U9985 (N_9985,N_5533,N_5667);
or U9986 (N_9986,N_5409,N_5616);
or U9987 (N_9987,N_5792,N_7403);
nor U9988 (N_9988,N_6236,N_6137);
xnor U9989 (N_9989,N_7311,N_7472);
xnor U9990 (N_9990,N_6114,N_6777);
nand U9991 (N_9991,N_7091,N_6197);
nand U9992 (N_9992,N_7164,N_5409);
or U9993 (N_9993,N_5708,N_7030);
nor U9994 (N_9994,N_6490,N_5116);
or U9995 (N_9995,N_6693,N_6665);
or U9996 (N_9996,N_5540,N_7019);
nand U9997 (N_9997,N_6680,N_7171);
xor U9998 (N_9998,N_5491,N_5247);
and U9999 (N_9999,N_5592,N_7486);
and U10000 (N_10000,N_7669,N_9924);
or U10001 (N_10001,N_8061,N_8806);
and U10002 (N_10002,N_8274,N_7731);
nand U10003 (N_10003,N_7561,N_9834);
xnor U10004 (N_10004,N_8126,N_8426);
and U10005 (N_10005,N_8399,N_8889);
xnor U10006 (N_10006,N_8744,N_8090);
or U10007 (N_10007,N_9102,N_9179);
nand U10008 (N_10008,N_7687,N_8443);
or U10009 (N_10009,N_9851,N_9552);
nand U10010 (N_10010,N_8020,N_8284);
or U10011 (N_10011,N_9893,N_7694);
or U10012 (N_10012,N_9481,N_7945);
nand U10013 (N_10013,N_9634,N_8936);
and U10014 (N_10014,N_9566,N_8603);
xnor U10015 (N_10015,N_9994,N_9105);
nand U10016 (N_10016,N_7696,N_9604);
nand U10017 (N_10017,N_8533,N_9396);
or U10018 (N_10018,N_9943,N_8336);
or U10019 (N_10019,N_8411,N_9240);
and U10020 (N_10020,N_7540,N_8618);
or U10021 (N_10021,N_9072,N_9565);
or U10022 (N_10022,N_9232,N_8287);
or U10023 (N_10023,N_8129,N_8259);
nor U10024 (N_10024,N_8225,N_7647);
nor U10025 (N_10025,N_7937,N_8439);
xnor U10026 (N_10026,N_8140,N_9981);
and U10027 (N_10027,N_8491,N_8160);
or U10028 (N_10028,N_9767,N_8453);
xor U10029 (N_10029,N_9425,N_8428);
and U10030 (N_10030,N_9722,N_9287);
nand U10031 (N_10031,N_9795,N_9688);
and U10032 (N_10032,N_7651,N_9131);
and U10033 (N_10033,N_8264,N_7592);
xor U10034 (N_10034,N_9182,N_9781);
nor U10035 (N_10035,N_9282,N_9819);
nor U10036 (N_10036,N_9450,N_8986);
nor U10037 (N_10037,N_8239,N_7867);
xnor U10038 (N_10038,N_8574,N_8954);
or U10039 (N_10039,N_8783,N_9522);
or U10040 (N_10040,N_8698,N_8731);
and U10041 (N_10041,N_8250,N_8525);
or U10042 (N_10042,N_8372,N_8114);
xnor U10043 (N_10043,N_9147,N_7819);
xor U10044 (N_10044,N_9486,N_7512);
xor U10045 (N_10045,N_8504,N_8522);
nand U10046 (N_10046,N_9163,N_8254);
nand U10047 (N_10047,N_8243,N_8570);
nand U10048 (N_10048,N_8103,N_9739);
xor U10049 (N_10049,N_9961,N_8261);
and U10050 (N_10050,N_9153,N_8375);
or U10051 (N_10051,N_8024,N_9247);
or U10052 (N_10052,N_7681,N_8031);
and U10053 (N_10053,N_9161,N_9038);
nor U10054 (N_10054,N_9034,N_9580);
and U10055 (N_10055,N_9510,N_7785);
xnor U10056 (N_10056,N_9007,N_7641);
nor U10057 (N_10057,N_7514,N_9435);
nor U10058 (N_10058,N_8653,N_8076);
nand U10059 (N_10059,N_8005,N_8384);
nand U10060 (N_10060,N_9397,N_8791);
nor U10061 (N_10061,N_8959,N_8348);
xor U10062 (N_10062,N_9668,N_7500);
and U10063 (N_10063,N_7718,N_9611);
and U10064 (N_10064,N_8328,N_9143);
nor U10065 (N_10065,N_8787,N_7515);
nand U10066 (N_10066,N_8033,N_8645);
nand U10067 (N_10067,N_7725,N_8374);
and U10068 (N_10068,N_9125,N_8000);
or U10069 (N_10069,N_8325,N_8467);
nand U10070 (N_10070,N_9132,N_8838);
nor U10071 (N_10071,N_8086,N_9364);
nor U10072 (N_10072,N_8978,N_9355);
nor U10073 (N_10073,N_8650,N_7902);
nand U10074 (N_10074,N_7831,N_9896);
or U10075 (N_10075,N_7730,N_8640);
nor U10076 (N_10076,N_8178,N_9244);
nor U10077 (N_10077,N_8257,N_9075);
and U10078 (N_10078,N_7633,N_8560);
xnor U10079 (N_10079,N_8980,N_9964);
nor U10080 (N_10080,N_9277,N_9890);
and U10081 (N_10081,N_8686,N_7903);
xor U10082 (N_10082,N_9198,N_9097);
and U10083 (N_10083,N_8923,N_8052);
xor U10084 (N_10084,N_8371,N_7848);
and U10085 (N_10085,N_9049,N_8711);
nand U10086 (N_10086,N_8098,N_9770);
and U10087 (N_10087,N_9672,N_9360);
and U10088 (N_10088,N_8565,N_8855);
and U10089 (N_10089,N_8726,N_9561);
nand U10090 (N_10090,N_9539,N_8768);
nor U10091 (N_10091,N_9606,N_8356);
nand U10092 (N_10092,N_8095,N_8065);
nor U10093 (N_10093,N_8790,N_9638);
or U10094 (N_10094,N_9667,N_8846);
or U10095 (N_10095,N_8001,N_8048);
or U10096 (N_10096,N_8938,N_9550);
nand U10097 (N_10097,N_7728,N_7792);
nand U10098 (N_10098,N_8104,N_8083);
xnor U10099 (N_10099,N_7671,N_9839);
xor U10100 (N_10100,N_9267,N_7572);
nor U10101 (N_10101,N_8755,N_8868);
nand U10102 (N_10102,N_9117,N_7897);
and U10103 (N_10103,N_9520,N_7533);
or U10104 (N_10104,N_8702,N_8432);
xnor U10105 (N_10105,N_7830,N_9710);
nor U10106 (N_10106,N_8493,N_9177);
nand U10107 (N_10107,N_8420,N_9379);
nor U10108 (N_10108,N_9024,N_7801);
and U10109 (N_10109,N_9926,N_8499);
and U10110 (N_10110,N_7690,N_7553);
xor U10111 (N_10111,N_9256,N_9879);
xor U10112 (N_10112,N_9378,N_9808);
xor U10113 (N_10113,N_8530,N_9938);
xor U10114 (N_10114,N_8720,N_9204);
nand U10115 (N_10115,N_7768,N_9400);
xor U10116 (N_10116,N_8394,N_9316);
xor U10117 (N_10117,N_7784,N_9508);
or U10118 (N_10118,N_7838,N_8277);
or U10119 (N_10119,N_9241,N_8767);
nor U10120 (N_10120,N_8183,N_9393);
or U10121 (N_10121,N_8282,N_7611);
and U10122 (N_10122,N_8575,N_8827);
and U10123 (N_10123,N_7814,N_9181);
or U10124 (N_10124,N_9597,N_9029);
or U10125 (N_10125,N_8144,N_7535);
or U10126 (N_10126,N_8405,N_9152);
xnor U10127 (N_10127,N_9050,N_8200);
or U10128 (N_10128,N_8634,N_9262);
nor U10129 (N_10129,N_8182,N_8311);
xor U10130 (N_10130,N_8485,N_9016);
nand U10131 (N_10131,N_9327,N_8648);
and U10132 (N_10132,N_9637,N_8012);
nand U10133 (N_10133,N_9031,N_7780);
nand U10134 (N_10134,N_8041,N_9503);
xnor U10135 (N_10135,N_8666,N_9923);
xor U10136 (N_10136,N_9404,N_8637);
xor U10137 (N_10137,N_9293,N_8919);
xnor U10138 (N_10138,N_8409,N_9333);
and U10139 (N_10139,N_9226,N_7762);
or U10140 (N_10140,N_8018,N_9423);
and U10141 (N_10141,N_8699,N_9209);
xnor U10142 (N_10142,N_7721,N_8623);
and U10143 (N_10143,N_8749,N_8106);
and U10144 (N_10144,N_8970,N_9903);
xor U10145 (N_10145,N_8376,N_8177);
nand U10146 (N_10146,N_8722,N_8404);
or U10147 (N_10147,N_9046,N_8059);
xnor U10148 (N_10148,N_9382,N_9058);
or U10149 (N_10149,N_7988,N_8147);
and U10150 (N_10150,N_8882,N_8351);
nand U10151 (N_10151,N_8946,N_9140);
or U10152 (N_10152,N_7652,N_9060);
and U10153 (N_10153,N_9185,N_9831);
nand U10154 (N_10154,N_8927,N_9136);
or U10155 (N_10155,N_9974,N_9040);
xnor U10156 (N_10156,N_7623,N_7948);
nor U10157 (N_10157,N_8292,N_7583);
or U10158 (N_10158,N_8445,N_9366);
nand U10159 (N_10159,N_8867,N_8102);
and U10160 (N_10160,N_7776,N_8361);
xnor U10161 (N_10161,N_7552,N_8554);
xor U10162 (N_10162,N_9801,N_8382);
and U10163 (N_10163,N_8937,N_9946);
nand U10164 (N_10164,N_8812,N_9982);
nor U10165 (N_10165,N_8926,N_9763);
nand U10166 (N_10166,N_8547,N_9933);
nand U10167 (N_10167,N_9236,N_8281);
or U10168 (N_10168,N_9035,N_9600);
nor U10169 (N_10169,N_8381,N_7981);
nor U10170 (N_10170,N_9250,N_7850);
or U10171 (N_10171,N_8856,N_9854);
xor U10172 (N_10172,N_9973,N_9625);
nor U10173 (N_10173,N_9560,N_7812);
nand U10174 (N_10174,N_9548,N_9211);
nand U10175 (N_10175,N_9986,N_9484);
nand U10176 (N_10176,N_8230,N_7699);
nand U10177 (N_10177,N_7970,N_8778);
or U10178 (N_10178,N_9299,N_9555);
and U10179 (N_10179,N_7567,N_9434);
nand U10180 (N_10180,N_8466,N_9726);
and U10181 (N_10181,N_7823,N_9339);
xor U10182 (N_10182,N_9084,N_8777);
xor U10183 (N_10183,N_9453,N_8089);
nor U10184 (N_10184,N_8258,N_9892);
and U10185 (N_10185,N_7501,N_8473);
xor U10186 (N_10186,N_9138,N_8630);
nand U10187 (N_10187,N_9718,N_9305);
xnor U10188 (N_10188,N_7817,N_8481);
or U10189 (N_10189,N_8263,N_7807);
or U10190 (N_10190,N_9330,N_9797);
or U10191 (N_10191,N_9899,N_9458);
xor U10192 (N_10192,N_7983,N_8814);
xnor U10193 (N_10193,N_9095,N_8668);
xor U10194 (N_10194,N_8172,N_9012);
xor U10195 (N_10195,N_7639,N_9289);
nand U10196 (N_10196,N_8690,N_7524);
nor U10197 (N_10197,N_8136,N_9681);
nor U10198 (N_10198,N_9409,N_9536);
nand U10199 (N_10199,N_9092,N_8171);
xor U10200 (N_10200,N_7582,N_8229);
or U10201 (N_10201,N_7570,N_9081);
nand U10202 (N_10202,N_9912,N_9067);
xor U10203 (N_10203,N_9671,N_8290);
or U10204 (N_10204,N_7846,N_8507);
xor U10205 (N_10205,N_8810,N_9094);
nand U10206 (N_10206,N_8111,N_7634);
or U10207 (N_10207,N_8319,N_8782);
nand U10208 (N_10208,N_8543,N_8070);
nand U10209 (N_10209,N_9771,N_9275);
and U10210 (N_10210,N_8933,N_8826);
or U10211 (N_10211,N_8784,N_8380);
or U10212 (N_10212,N_9288,N_8951);
nand U10213 (N_10213,N_9459,N_8793);
nor U10214 (N_10214,N_8987,N_9817);
xor U10215 (N_10215,N_8246,N_8370);
nor U10216 (N_10216,N_8527,N_7859);
xnor U10217 (N_10217,N_8809,N_7542);
xnor U10218 (N_10218,N_9874,N_9215);
nor U10219 (N_10219,N_7824,N_8629);
and U10220 (N_10220,N_7861,N_9569);
nand U10221 (N_10221,N_8419,N_8515);
xor U10222 (N_10222,N_9314,N_8644);
or U10223 (N_10223,N_7832,N_8217);
xnor U10224 (N_10224,N_7788,N_8056);
and U10225 (N_10225,N_8393,N_7711);
xnor U10226 (N_10226,N_7982,N_9609);
or U10227 (N_10227,N_9533,N_8685);
nor U10228 (N_10228,N_8154,N_8053);
xnor U10229 (N_10229,N_8847,N_9922);
nand U10230 (N_10230,N_7714,N_9804);
and U10231 (N_10231,N_8143,N_8609);
and U10232 (N_10232,N_8684,N_9729);
or U10233 (N_10233,N_8683,N_7640);
or U10234 (N_10234,N_9989,N_9937);
nor U10235 (N_10235,N_9862,N_9587);
xnor U10236 (N_10236,N_9608,N_8181);
nor U10237 (N_10237,N_9649,N_8823);
nor U10238 (N_10238,N_8446,N_8843);
or U10239 (N_10239,N_8479,N_7560);
or U10240 (N_10240,N_7506,N_8478);
xnor U10241 (N_10241,N_8349,N_9723);
xnor U10242 (N_10242,N_7673,N_7769);
or U10243 (N_10243,N_8006,N_7607);
and U10244 (N_10244,N_8664,N_9821);
nand U10245 (N_10245,N_9412,N_8004);
and U10246 (N_10246,N_8624,N_9919);
nand U10247 (N_10247,N_8444,N_8423);
xnor U10248 (N_10248,N_8895,N_7949);
or U10249 (N_10249,N_8231,N_9605);
and U10250 (N_10250,N_7740,N_9054);
nor U10251 (N_10251,N_8400,N_8063);
or U10252 (N_10252,N_7763,N_8656);
and U10253 (N_10253,N_7891,N_8465);
nand U10254 (N_10254,N_8825,N_9384);
and U10255 (N_10255,N_9166,N_8576);
xor U10256 (N_10256,N_9374,N_9253);
xnor U10257 (N_10257,N_8861,N_8733);
xnor U10258 (N_10258,N_9653,N_8240);
nor U10259 (N_10259,N_7624,N_7794);
nor U10260 (N_10260,N_9074,N_7606);
xor U10261 (N_10261,N_7894,N_7736);
xor U10262 (N_10262,N_9523,N_9123);
nand U10263 (N_10263,N_8360,N_7680);
nand U10264 (N_10264,N_9853,N_7627);
nand U10265 (N_10265,N_7765,N_8730);
or U10266 (N_10266,N_8027,N_8416);
or U10267 (N_10267,N_8635,N_8128);
or U10268 (N_10268,N_7940,N_9659);
and U10269 (N_10269,N_9913,N_7907);
xor U10270 (N_10270,N_9113,N_8235);
xor U10271 (N_10271,N_9243,N_8222);
xor U10272 (N_10272,N_7944,N_9535);
nand U10273 (N_10273,N_8100,N_7756);
xor U10274 (N_10274,N_8321,N_7920);
or U10275 (N_10275,N_8367,N_7919);
nand U10276 (N_10276,N_7523,N_9342);
or U10277 (N_10277,N_9189,N_9370);
nand U10278 (N_10278,N_7688,N_9008);
nand U10279 (N_10279,N_7781,N_9942);
and U10280 (N_10280,N_8770,N_8109);
nor U10281 (N_10281,N_8494,N_9551);
or U10282 (N_10282,N_9660,N_8194);
or U10283 (N_10283,N_7929,N_8245);
nor U10284 (N_10284,N_9794,N_8511);
nand U10285 (N_10285,N_7893,N_7620);
or U10286 (N_10286,N_7536,N_9640);
nor U10287 (N_10287,N_9789,N_9106);
xnor U10288 (N_10288,N_9880,N_8304);
xnor U10289 (N_10289,N_9354,N_9515);
nand U10290 (N_10290,N_9971,N_9077);
nor U10291 (N_10291,N_9875,N_7899);
or U10292 (N_10292,N_8813,N_8836);
and U10293 (N_10293,N_8654,N_9583);
nand U10294 (N_10294,N_8537,N_7986);
nor U10295 (N_10295,N_9344,N_7521);
or U10296 (N_10296,N_8953,N_9297);
nand U10297 (N_10297,N_9571,N_9061);
xor U10298 (N_10298,N_9888,N_8971);
xor U10299 (N_10299,N_8617,N_9765);
xnor U10300 (N_10300,N_7643,N_8158);
nand U10301 (N_10301,N_7519,N_9741);
and U10302 (N_10302,N_8312,N_9784);
xnor U10303 (N_10303,N_9742,N_8622);
nand U10304 (N_10304,N_7742,N_9644);
and U10305 (N_10305,N_8452,N_8950);
nand U10306 (N_10306,N_7663,N_7974);
or U10307 (N_10307,N_8191,N_8584);
nand U10308 (N_10308,N_8687,N_8712);
or U10309 (N_10309,N_8262,N_7895);
nor U10310 (N_10310,N_8459,N_8119);
xor U10311 (N_10311,N_8205,N_8794);
nand U10312 (N_10312,N_8363,N_9184);
nor U10313 (N_10313,N_9151,N_9208);
nand U10314 (N_10314,N_8976,N_8669);
or U10315 (N_10315,N_8430,N_8947);
nand U10316 (N_10316,N_9513,N_9304);
and U10317 (N_10317,N_9005,N_7892);
nand U10318 (N_10318,N_9658,N_8665);
or U10319 (N_10319,N_9323,N_9957);
xnor U10320 (N_10320,N_9042,N_8280);
nor U10321 (N_10321,N_7616,N_8449);
or U10322 (N_10322,N_8115,N_8117);
or U10323 (N_10323,N_8567,N_9670);
nand U10324 (N_10324,N_7576,N_7682);
nand U10325 (N_10325,N_8204,N_9401);
xnor U10326 (N_10326,N_8773,N_7834);
and U10327 (N_10327,N_8188,N_9891);
nand U10328 (N_10328,N_9696,N_7588);
xor U10329 (N_10329,N_7855,N_7556);
and U10330 (N_10330,N_8415,N_7549);
nand U10331 (N_10331,N_8993,N_9415);
nand U10332 (N_10332,N_8237,N_8973);
and U10333 (N_10333,N_9750,N_9978);
nor U10334 (N_10334,N_9233,N_9646);
nor U10335 (N_10335,N_8030,N_9692);
nand U10336 (N_10336,N_9391,N_9712);
nor U10337 (N_10337,N_9227,N_8307);
nand U10338 (N_10338,N_8450,N_7558);
or U10339 (N_10339,N_9180,N_8228);
nand U10340 (N_10340,N_8022,N_8845);
or U10341 (N_10341,N_8910,N_8192);
nor U10342 (N_10342,N_9709,N_8285);
nor U10343 (N_10343,N_7888,N_9183);
or U10344 (N_10344,N_9258,N_9169);
xnor U10345 (N_10345,N_9492,N_8403);
nor U10346 (N_10346,N_7637,N_7666);
and U10347 (N_10347,N_7551,N_9932);
or U10348 (N_10348,N_8410,N_9736);
xnor U10349 (N_10349,N_8613,N_9114);
nand U10350 (N_10350,N_8969,N_7569);
nand U10351 (N_10351,N_9955,N_9015);
nor U10352 (N_10352,N_7766,N_8700);
and U10353 (N_10353,N_9628,N_9908);
nand U10354 (N_10354,N_7635,N_7581);
and U10355 (N_10355,N_9787,N_9811);
xor U10356 (N_10356,N_8967,N_8998);
nand U10357 (N_10357,N_9642,N_7918);
nor U10358 (N_10358,N_8692,N_9348);
nand U10359 (N_10359,N_9694,N_9822);
xor U10360 (N_10360,N_9099,N_9849);
and U10361 (N_10361,N_8462,N_9705);
and U10362 (N_10362,N_7962,N_8146);
or U10363 (N_10363,N_9501,N_8865);
and U10364 (N_10364,N_7923,N_8518);
nor U10365 (N_10365,N_7770,N_9438);
nand U10366 (N_10366,N_7702,N_8579);
nor U10367 (N_10367,N_9684,N_7909);
nand U10368 (N_10368,N_7978,N_9641);
xnor U10369 (N_10369,N_8344,N_8691);
nor U10370 (N_10370,N_8387,N_8124);
and U10371 (N_10371,N_8903,N_8358);
and U10372 (N_10372,N_7729,N_9969);
nand U10373 (N_10373,N_8600,N_7664);
xnor U10374 (N_10374,N_9915,N_7954);
nor U10375 (N_10375,N_8273,N_7516);
or U10376 (N_10376,N_7589,N_9086);
nand U10377 (N_10377,N_8091,N_8580);
nor U10378 (N_10378,N_8837,N_9776);
or U10379 (N_10379,N_9272,N_9477);
nor U10380 (N_10380,N_7648,N_9442);
and U10381 (N_10381,N_8614,N_9907);
and U10382 (N_10382,N_9619,N_7713);
nor U10383 (N_10383,N_7779,N_7939);
nor U10384 (N_10384,N_9349,N_9698);
nor U10385 (N_10385,N_8299,N_7672);
or U10386 (N_10386,N_9996,N_9499);
and U10387 (N_10387,N_8853,N_7719);
nand U10388 (N_10388,N_9708,N_9193);
nand U10389 (N_10389,N_9167,N_9753);
or U10390 (N_10390,N_9457,N_9863);
nor U10391 (N_10391,N_9351,N_7999);
nand U10392 (N_10392,N_9388,N_9329);
or U10393 (N_10393,N_7979,N_7550);
nand U10394 (N_10394,N_8226,N_9298);
or U10395 (N_10395,N_9900,N_7679);
nor U10396 (N_10396,N_9706,N_9895);
nor U10397 (N_10397,N_8113,N_8815);
or U10398 (N_10398,N_8835,N_8829);
nor U10399 (N_10399,N_8477,N_8539);
or U10400 (N_10400,N_8206,N_9228);
or U10401 (N_10401,N_9768,N_8101);
nor U10402 (N_10402,N_9021,N_7532);
nor U10403 (N_10403,N_9365,N_9413);
nor U10404 (N_10404,N_9371,N_9011);
or U10405 (N_10405,N_8558,N_8424);
or U10406 (N_10406,N_8197,N_7998);
or U10407 (N_10407,N_8379,N_9655);
or U10408 (N_10408,N_9968,N_8639);
nand U10409 (N_10409,N_9857,N_9856);
xnor U10410 (N_10410,N_8887,N_8215);
xor U10411 (N_10411,N_8710,N_9213);
nand U10412 (N_10412,N_9279,N_7615);
xnor U10413 (N_10413,N_7879,N_8286);
nor U10414 (N_10414,N_8077,N_9216);
and U10415 (N_10415,N_8460,N_9221);
nor U10416 (N_10416,N_8714,N_7659);
and U10417 (N_10417,N_9647,N_8786);
and U10418 (N_10418,N_9128,N_8725);
or U10419 (N_10419,N_9291,N_9278);
nor U10420 (N_10420,N_8981,N_8906);
xor U10421 (N_10421,N_8353,N_8159);
nand U10422 (N_10422,N_7543,N_9172);
xor U10423 (N_10423,N_8877,N_7836);
xnor U10424 (N_10424,N_9559,N_9576);
nor U10425 (N_10425,N_9737,N_9663);
or U10426 (N_10426,N_9301,N_9917);
nand U10427 (N_10427,N_8435,N_9991);
and U10428 (N_10428,N_9249,N_8412);
xor U10429 (N_10429,N_9069,N_8116);
nor U10430 (N_10430,N_8924,N_8441);
nor U10431 (N_10431,N_9855,N_7710);
nand U10432 (N_10432,N_9773,N_9290);
or U10433 (N_10433,N_9998,N_8604);
xor U10434 (N_10434,N_8072,N_9848);
nand U10435 (N_10435,N_8357,N_8572);
nor U10436 (N_10436,N_9420,N_8619);
or U10437 (N_10437,N_8081,N_9758);
nor U10438 (N_10438,N_8772,N_9427);
or U10439 (N_10439,N_7874,N_9487);
nor U10440 (N_10440,N_7808,N_8501);
nor U10441 (N_10441,N_9041,N_9721);
xor U10442 (N_10442,N_9341,N_7590);
and U10443 (N_10443,N_9951,N_9433);
xor U10444 (N_10444,N_8727,N_9695);
nor U10445 (N_10445,N_8766,N_8999);
nand U10446 (N_10446,N_8084,N_8017);
nand U10447 (N_10447,N_7605,N_8750);
nor U10448 (N_10448,N_8148,N_8442);
nor U10449 (N_10449,N_8509,N_9199);
or U10450 (N_10450,N_8152,N_8520);
xnor U10451 (N_10451,N_8538,N_9121);
xnor U10452 (N_10452,N_8037,N_8740);
xor U10453 (N_10453,N_8649,N_8628);
nand U10454 (N_10454,N_9877,N_8288);
nand U10455 (N_10455,N_7987,N_7946);
and U10456 (N_10456,N_8094,N_9636);
xor U10457 (N_10457,N_7693,N_7636);
and U10458 (N_10458,N_7802,N_8427);
nor U10459 (N_10459,N_7915,N_9633);
nand U10460 (N_10460,N_7594,N_9357);
nand U10461 (N_10461,N_9500,N_9159);
and U10462 (N_10462,N_8392,N_9219);
xnor U10463 (N_10463,N_8193,N_9246);
nand U10464 (N_10464,N_9562,N_8941);
or U10465 (N_10465,N_7700,N_8821);
xnor U10466 (N_10466,N_9144,N_8422);
and U10467 (N_10467,N_8289,N_9626);
and U10468 (N_10468,N_8737,N_9790);
xnor U10469 (N_10469,N_8536,N_7689);
nor U10470 (N_10470,N_9764,N_8220);
and U10471 (N_10471,N_9308,N_8717);
nor U10472 (N_10472,N_9346,N_9976);
nor U10473 (N_10473,N_7658,N_7804);
xor U10474 (N_10474,N_8035,N_9368);
and U10475 (N_10475,N_8896,N_7670);
or U10476 (N_10476,N_9174,N_9703);
and U10477 (N_10477,N_9156,N_9883);
xor U10478 (N_10478,N_7930,N_8524);
xor U10479 (N_10479,N_8820,N_9623);
xnor U10480 (N_10480,N_7657,N_8674);
xnor U10481 (N_10481,N_8383,N_8122);
xor U10482 (N_10482,N_7889,N_9292);
nor U10483 (N_10483,N_9700,N_8626);
or U10484 (N_10484,N_9683,N_9098);
xnor U10485 (N_10485,N_7691,N_9137);
or U10486 (N_10486,N_8093,N_9643);
xnor U10487 (N_10487,N_9904,N_9018);
or U10488 (N_10488,N_9124,N_7741);
xnor U10489 (N_10489,N_8042,N_9935);
nand U10490 (N_10490,N_9884,N_9043);
nor U10491 (N_10491,N_8345,N_7864);
or U10492 (N_10492,N_8928,N_8055);
or U10493 (N_10493,N_9345,N_9494);
nand U10494 (N_10494,N_8247,N_7996);
nor U10495 (N_10495,N_8503,N_7782);
nor U10496 (N_10496,N_9734,N_9940);
nor U10497 (N_10497,N_9352,N_8131);
nor U10498 (N_10498,N_7900,N_8211);
and U10499 (N_10499,N_7618,N_9443);
xnor U10500 (N_10500,N_8858,N_9101);
nand U10501 (N_10501,N_9088,N_8992);
and U10502 (N_10502,N_8899,N_8464);
nand U10503 (N_10503,N_8120,N_7863);
xnor U10504 (N_10504,N_8023,N_9203);
nor U10505 (N_10505,N_9025,N_9607);
or U10506 (N_10506,N_8064,N_8859);
nand U10507 (N_10507,N_9343,N_7809);
nand U10508 (N_10508,N_9390,N_9837);
nand U10509 (N_10509,N_7761,N_8003);
nand U10510 (N_10510,N_7504,N_9909);
and U10511 (N_10511,N_8590,N_8627);
nand U10512 (N_10512,N_9129,N_7667);
nor U10513 (N_10513,N_9373,N_7732);
xnor U10514 (N_10514,N_7904,N_9680);
and U10515 (N_10515,N_8327,N_9052);
xor U10516 (N_10516,N_7628,N_8917);
xnor U10517 (N_10517,N_8811,N_8661);
and U10518 (N_10518,N_7562,N_8354);
and U10519 (N_10519,N_7518,N_7822);
and U10520 (N_10520,N_7827,N_7966);
nand U10521 (N_10521,N_9516,N_9752);
xor U10522 (N_10522,N_9358,N_9630);
nor U10523 (N_10523,N_7580,N_9376);
and U10524 (N_10524,N_9687,N_8180);
xnor U10525 (N_10525,N_8918,N_9263);
or U10526 (N_10526,N_9059,N_9673);
or U10527 (N_10527,N_9595,N_8212);
nand U10528 (N_10528,N_7885,N_8689);
nor U10529 (N_10529,N_8632,N_8985);
and U10530 (N_10530,N_8242,N_7829);
nor U10531 (N_10531,N_9003,N_8173);
nor U10532 (N_10532,N_7701,N_8391);
nor U10533 (N_10533,N_8300,N_8021);
xnor U10534 (N_10534,N_9044,N_7748);
xor U10535 (N_10535,N_8474,N_9534);
xnor U10536 (N_10536,N_7798,N_9280);
and U10537 (N_10537,N_8943,N_9980);
and U10538 (N_10538,N_8955,N_7803);
xor U10539 (N_10539,N_8483,N_7810);
nand U10540 (N_10540,N_8703,N_9568);
xnor U10541 (N_10541,N_9104,N_9313);
xnor U10542 (N_10542,N_7957,N_7773);
or U10543 (N_10543,N_7811,N_8233);
nand U10544 (N_10544,N_9451,N_9732);
and U10545 (N_10545,N_8893,N_8581);
or U10546 (N_10546,N_8704,N_8870);
or U10547 (N_10547,N_8534,N_7815);
nand U10548 (N_10548,N_8886,N_9239);
xnor U10549 (N_10549,N_9230,N_9283);
or U10550 (N_10550,N_7676,N_8852);
nor U10551 (N_10551,N_7835,N_8911);
nand U10552 (N_10552,N_9586,N_9531);
and U10553 (N_10553,N_9234,N_8832);
and U10554 (N_10554,N_8014,N_8974);
xor U10555 (N_10555,N_8545,N_7557);
xor U10556 (N_10556,N_7598,N_9222);
xnor U10557 (N_10557,N_9497,N_9777);
or U10558 (N_10558,N_8002,N_8050);
and U10559 (N_10559,N_9887,N_8913);
nand U10560 (N_10560,N_8996,N_7744);
xnor U10561 (N_10561,N_9806,N_8655);
xor U10562 (N_10562,N_9835,N_7632);
nor U10563 (N_10563,N_9859,N_8802);
and U10564 (N_10564,N_9910,N_9463);
nand U10565 (N_10565,N_8139,N_9073);
nand U10566 (N_10566,N_8378,N_9334);
nand U10567 (N_10567,N_9507,N_8025);
or U10568 (N_10568,N_8834,N_9666);
and U10569 (N_10569,N_9885,N_9745);
or U10570 (N_10570,N_8972,N_8232);
and U10571 (N_10571,N_9432,N_9632);
xor U10572 (N_10572,N_9437,N_7953);
xnor U10573 (N_10573,N_9727,N_9911);
and U10574 (N_10574,N_9191,N_8688);
xnor U10575 (N_10575,N_9558,N_8385);
xnor U10576 (N_10576,N_9774,N_7901);
nor U10577 (N_10577,N_9861,N_8615);
xnor U10578 (N_10578,N_7602,N_8352);
or U10579 (N_10579,N_8330,N_7882);
and U10580 (N_10580,N_7505,N_8339);
or U10581 (N_10581,N_7674,N_8675);
nand U10582 (N_10582,N_9266,N_8302);
or U10583 (N_10583,N_8592,N_8716);
nor U10584 (N_10584,N_9554,N_9296);
or U10585 (N_10585,N_7712,N_8642);
nand U10586 (N_10586,N_8607,N_8071);
nor U10587 (N_10587,N_7530,N_7997);
and U10588 (N_10588,N_9631,N_9027);
and U10589 (N_10589,N_9078,N_9319);
nand U10590 (N_10590,N_9852,N_8407);
nand U10591 (N_10591,N_8301,N_7875);
or U10592 (N_10592,N_8347,N_7797);
and U10593 (N_10593,N_8774,N_7960);
and U10594 (N_10594,N_8482,N_9017);
xor U10595 (N_10595,N_9905,N_9820);
nor U10596 (N_10596,N_8082,N_8073);
or U10597 (N_10597,N_8492,N_8269);
and U10598 (N_10598,N_9573,N_9719);
nand U10599 (N_10599,N_8236,N_9830);
xnor U10600 (N_10600,N_8087,N_9422);
nand U10601 (N_10601,N_7963,N_8549);
or U10602 (N_10602,N_9402,N_8553);
nor U10603 (N_10603,N_8715,N_7717);
and U10604 (N_10604,N_8529,N_8792);
xor U10605 (N_10605,N_8564,N_8818);
and U10606 (N_10606,N_7968,N_9269);
and U10607 (N_10607,N_8315,N_7912);
xnor U10608 (N_10608,N_9112,N_7771);
nand U10609 (N_10609,N_9881,N_9563);
xnor U10610 (N_10610,N_8036,N_9010);
and U10611 (N_10611,N_9871,N_8841);
and U10612 (N_10612,N_8697,N_7967);
or U10613 (N_10613,N_9385,N_9004);
nand U10614 (N_10614,N_8454,N_9841);
nand U10615 (N_10615,N_8914,N_9452);
nor U10616 (N_10616,N_9134,N_9925);
xor U10617 (N_10617,N_9449,N_7760);
nor U10618 (N_10618,N_8966,N_7517);
or U10619 (N_10619,N_9530,N_9403);
nand U10620 (N_10620,N_9386,N_7943);
nor U10621 (N_10621,N_7853,N_9840);
xor U10622 (N_10622,N_8546,N_9307);
xnor U10623 (N_10623,N_9218,N_7621);
and U10624 (N_10624,N_8293,N_9429);
nand U10625 (N_10625,N_9541,N_8851);
xor U10626 (N_10626,N_8573,N_9603);
or U10627 (N_10627,N_7821,N_8643);
nand U10628 (N_10628,N_7653,N_9567);
or U10629 (N_10629,N_8272,N_7914);
and U10630 (N_10630,N_9627,N_8209);
nor U10631 (N_10631,N_9148,N_9679);
xnor U10632 (N_10632,N_7924,N_8673);
nor U10633 (N_10633,N_7753,N_9546);
nand U10634 (N_10634,N_8141,N_8164);
nor U10635 (N_10635,N_8541,N_8900);
nand U10636 (N_10636,N_8659,N_8413);
or U10637 (N_10637,N_8577,N_7527);
and U10638 (N_10638,N_9273,N_7984);
or U10639 (N_10639,N_8046,N_9738);
and U10640 (N_10640,N_8939,N_8857);
xor U10641 (N_10641,N_8198,N_7520);
and U10642 (N_10642,N_8747,N_9332);
nand U10643 (N_10643,N_8196,N_9941);
xor U10644 (N_10644,N_8651,N_7692);
xor U10645 (N_10645,N_7869,N_8185);
nor U10646 (N_10646,N_8170,N_7833);
nor U10647 (N_10647,N_9825,N_9171);
nor U10648 (N_10648,N_9898,N_8088);
nand U10649 (N_10649,N_7507,N_8085);
nor U10650 (N_10650,N_7843,N_9048);
and U10651 (N_10651,N_9190,N_8758);
nor U10652 (N_10652,N_7529,N_8862);
and U10653 (N_10653,N_9544,N_8963);
xnor U10654 (N_10654,N_9096,N_7825);
or U10655 (N_10655,N_8118,N_8601);
xor U10656 (N_10656,N_9460,N_9950);
nand U10657 (N_10657,N_8223,N_9972);
nor U10658 (N_10658,N_7548,N_8149);
nor U10659 (N_10659,N_8706,N_8952);
xor U10660 (N_10660,N_9066,N_8157);
nand U10661 (N_10661,N_8219,N_9707);
and U10662 (N_10662,N_9635,N_9116);
nor U10663 (N_10663,N_9802,N_9194);
and U10664 (N_10664,N_8105,N_9843);
or U10665 (N_10665,N_8038,N_8043);
nor U10666 (N_10666,N_7858,N_8256);
or U10667 (N_10667,N_7705,N_9410);
nand U10668 (N_10668,N_7965,N_7752);
xor U10669 (N_10669,N_8599,N_9495);
nor U10670 (N_10670,N_9699,N_7757);
nand U10671 (N_10671,N_8099,N_8935);
or U10672 (N_10672,N_9108,N_8934);
and U10673 (N_10673,N_9650,N_7655);
and U10674 (N_10674,N_9735,N_9109);
and U10675 (N_10675,N_7544,N_8161);
xnor U10676 (N_10676,N_7587,N_9214);
nand U10677 (N_10677,N_9200,N_9257);
and U10678 (N_10678,N_9051,N_9711);
nor U10679 (N_10679,N_7727,N_9949);
and U10680 (N_10680,N_7545,N_8238);
and U10681 (N_10681,N_8587,N_9873);
and U10682 (N_10682,N_8418,N_7707);
xor U10683 (N_10683,N_9255,N_8342);
xnor U10684 (N_10684,N_9844,N_9997);
and U10685 (N_10685,N_9062,N_7614);
nand U10686 (N_10686,N_9306,N_9829);
xor U10687 (N_10687,N_9947,N_8807);
nand U10688 (N_10688,N_9897,N_8519);
xor U10689 (N_10689,N_8047,N_7884);
xnor U10690 (N_10690,N_8265,N_7575);
xnor U10691 (N_10691,N_9115,N_8500);
nand U10692 (N_10692,N_7629,N_8854);
nor U10693 (N_10693,N_8092,N_8531);
or U10694 (N_10694,N_8625,N_9579);
or U10695 (N_10695,N_9085,N_8753);
nor U10696 (N_10696,N_8819,N_9009);
nor U10697 (N_10697,N_8029,N_8894);
nand U10698 (N_10698,N_9466,N_7783);
or U10699 (N_10699,N_9780,N_9574);
or U10700 (N_10700,N_8708,N_8267);
nor U10701 (N_10701,N_9845,N_9444);
and U10702 (N_10702,N_8723,N_9514);
and U10703 (N_10703,N_7816,N_7839);
or U10704 (N_10704,N_8804,N_8646);
or U10705 (N_10705,N_8742,N_9584);
nor U10706 (N_10706,N_7793,N_8436);
xor U10707 (N_10707,N_9419,N_9577);
and U10708 (N_10708,N_9894,N_8458);
nand U10709 (N_10709,N_9261,N_7746);
nor U10710 (N_10710,N_7820,N_7555);
nand U10711 (N_10711,N_7599,N_8165);
nand U10712 (N_10712,N_9248,N_9621);
nand U10713 (N_10713,N_9476,N_8563);
or U10714 (N_10714,N_7574,N_8308);
nand U10715 (N_10715,N_7739,N_7928);
xor U10716 (N_10716,N_9818,N_9175);
nand U10717 (N_10717,N_7715,N_9381);
xnor U10718 (N_10718,N_7980,N_7786);
nor U10719 (N_10719,N_8060,N_9921);
xnor U10720 (N_10720,N_8979,N_8881);
or U10721 (N_10721,N_8447,N_9446);
xor U10722 (N_10722,N_9599,N_9999);
and U10723 (N_10723,N_8875,N_9070);
nor U10724 (N_10724,N_8550,N_7539);
or U10725 (N_10725,N_9869,N_8902);
nand U10726 (N_10726,N_9268,N_9992);
xnor U10727 (N_10727,N_8658,N_7601);
xnor U10728 (N_10728,N_8752,N_9398);
nand U10729 (N_10729,N_9490,N_8251);
nor U10730 (N_10730,N_8879,N_8968);
and U10731 (N_10731,N_8130,N_8224);
nor U10732 (N_10732,N_9170,N_8808);
xor U10733 (N_10733,N_9164,N_8011);
and U10734 (N_10734,N_8457,N_8320);
and U10735 (N_10735,N_8561,N_8368);
and U10736 (N_10736,N_7644,N_7706);
nand U10737 (N_10737,N_8578,N_7564);
nand U10738 (N_10738,N_9053,N_9809);
xnor U10739 (N_10739,N_9733,N_8296);
and U10740 (N_10740,N_9591,N_9716);
or U10741 (N_10741,N_9033,N_7678);
nand U10742 (N_10742,N_9392,N_7951);
and U10743 (N_10743,N_8695,N_8125);
nor U10744 (N_10744,N_8512,N_9528);
xnor U10745 (N_10745,N_8366,N_9755);
xnor U10746 (N_10746,N_7865,N_8860);
or U10747 (N_10747,N_8513,N_9119);
or U10748 (N_10748,N_8514,N_7985);
nand U10749 (N_10749,N_8800,N_8638);
or U10750 (N_10750,N_9759,N_7724);
xnor U10751 (N_10751,N_8487,N_8169);
nor U10752 (N_10752,N_8738,N_9614);
and U10753 (N_10753,N_9440,N_8724);
nor U10754 (N_10754,N_8878,N_9945);
xor U10755 (N_10755,N_9271,N_9076);
or U10756 (N_10756,N_9265,N_8516);
xor U10757 (N_10757,N_8335,N_9928);
and U10758 (N_10758,N_9080,N_9697);
or U10759 (N_10759,N_8341,N_8540);
nand U10760 (N_10760,N_8278,N_8309);
xnor U10761 (N_10761,N_7660,N_7913);
nor U10762 (N_10762,N_7510,N_8765);
or U10763 (N_10763,N_8839,N_7931);
nand U10764 (N_10764,N_9701,N_8528);
or U10765 (N_10765,N_8605,N_9772);
or U10766 (N_10766,N_8521,N_7709);
xnor U10767 (N_10767,N_8762,N_8163);
xnor U10768 (N_10768,N_9657,N_8276);
nand U10769 (N_10769,N_7977,N_8798);
and U10770 (N_10770,N_8763,N_9447);
nor U10771 (N_10771,N_9782,N_9675);
xor U10772 (N_10772,N_7845,N_7847);
nand U10773 (N_10773,N_7778,N_8785);
and U10774 (N_10774,N_9740,N_8472);
xnor U10775 (N_10775,N_7935,N_8401);
xnor U10776 (N_10776,N_8156,N_7608);
or U10777 (N_10777,N_7840,N_8801);
nand U10778 (N_10778,N_9870,N_9962);
nand U10779 (N_10779,N_9220,N_7559);
or U10780 (N_10780,N_8880,N_8068);
nand U10781 (N_10781,N_7538,N_8075);
xor U10782 (N_10782,N_9865,N_7565);
nor U10783 (N_10783,N_9963,N_9967);
nor U10784 (N_10784,N_9496,N_9775);
nor U10785 (N_10785,N_7932,N_8833);
xor U10786 (N_10786,N_9610,N_8313);
or U10787 (N_10787,N_8015,N_7665);
nor U10788 (N_10788,N_7883,N_7563);
xor U10789 (N_10789,N_9532,N_9988);
nor U10790 (N_10790,N_8057,N_8523);
and U10791 (N_10791,N_8764,N_9578);
nor U10792 (N_10792,N_9842,N_7733);
nand U10793 (N_10793,N_8962,N_9464);
xnor U10794 (N_10794,N_7584,N_9353);
nor U10795 (N_10795,N_9019,N_8678);
nor U10796 (N_10796,N_8891,N_7767);
xor U10797 (N_10797,N_8396,N_9596);
nor U10798 (N_10798,N_7841,N_9006);
and U10799 (N_10799,N_8677,N_7697);
or U10800 (N_10800,N_7638,N_8476);
nand U10801 (N_10801,N_8316,N_8922);
xnor U10802 (N_10802,N_8034,N_7675);
or U10803 (N_10803,N_7787,N_8334);
and U10804 (N_10804,N_9110,N_8249);
or U10805 (N_10805,N_8597,N_8713);
or U10806 (N_10806,N_9788,N_8797);
nor U10807 (N_10807,N_9648,N_7654);
xnor U10808 (N_10808,N_7926,N_9762);
xor U10809 (N_10809,N_8636,N_9920);
and U10810 (N_10810,N_8298,N_9286);
and U10811 (N_10811,N_9549,N_7626);
nor U10812 (N_10812,N_8662,N_9876);
and U10813 (N_10813,N_9524,N_7683);
or U10814 (N_10814,N_9310,N_9757);
nand U10815 (N_10815,N_9622,N_8402);
nor U10816 (N_10816,N_8994,N_8754);
or U10817 (N_10817,N_8408,N_8871);
and U10818 (N_10818,N_8390,N_7645);
nand U10819 (N_10819,N_8097,N_9939);
or U10820 (N_10820,N_8932,N_9302);
and U10821 (N_10821,N_7578,N_9411);
nand U10822 (N_10822,N_9965,N_8145);
xnor U10823 (N_10823,N_7952,N_9540);
nand U10824 (N_10824,N_8051,N_8275);
and U10825 (N_10825,N_9320,N_8471);
xor U10826 (N_10826,N_9377,N_8925);
nor U10827 (N_10827,N_9426,N_8074);
nor U10828 (N_10828,N_8942,N_8045);
nand U10829 (N_10829,N_7958,N_8451);
xor U10830 (N_10830,N_8468,N_9761);
nand U10831 (N_10831,N_8369,N_7990);
xor U10832 (N_10832,N_7872,N_7513);
nor U10833 (N_10833,N_9186,N_8680);
nor U10834 (N_10834,N_9620,N_9954);
xnor U10835 (N_10835,N_9324,N_9037);
xor U10836 (N_10836,N_7772,N_8270);
and U10837 (N_10837,N_7596,N_9868);
nand U10838 (N_10838,N_9195,N_8732);
and U10839 (N_10839,N_8983,N_8912);
nor U10840 (N_10840,N_9087,N_8216);
nor U10841 (N_10841,N_7795,N_8965);
xnor U10842 (N_10842,N_9953,N_9285);
and U10843 (N_10843,N_8890,N_9704);
nand U10844 (N_10844,N_9485,N_9424);
nand U10845 (N_10845,N_9724,N_9483);
and U10846 (N_10846,N_7964,N_8647);
nor U10847 (N_10847,N_7973,N_9235);
nand U10848 (N_10848,N_9461,N_8679);
nand U10849 (N_10849,N_9303,N_8310);
nor U10850 (N_10850,N_9356,N_9975);
and U10851 (N_10851,N_9055,N_9807);
and U10852 (N_10852,N_8123,N_9001);
xor U10853 (N_10853,N_9064,N_8377);
and U10854 (N_10854,N_9126,N_8314);
and U10855 (N_10855,N_9545,N_8995);
and U10856 (N_10856,N_9375,N_9103);
nor U10857 (N_10857,N_7541,N_8438);
nand U10858 (N_10858,N_9803,N_9321);
or U10859 (N_10859,N_9677,N_9118);
nor U10860 (N_10860,N_7877,N_9431);
xor U10861 (N_10861,N_9047,N_7642);
nand U10862 (N_10862,N_9328,N_8593);
nor U10863 (N_10863,N_9335,N_7871);
and U10864 (N_10864,N_9512,N_7704);
nor U10865 (N_10865,N_8748,N_9960);
or U10866 (N_10866,N_8054,N_9827);
nand U10867 (N_10867,N_9509,N_9952);
or U10868 (N_10868,N_8032,N_9867);
or U10869 (N_10869,N_9956,N_9783);
nor U10870 (N_10870,N_8869,N_7503);
nand U10871 (N_10871,N_7622,N_9418);
nand U10872 (N_10872,N_8921,N_8517);
and U10873 (N_10873,N_9471,N_9178);
nor U10874 (N_10874,N_8333,N_8324);
or U10875 (N_10875,N_9714,N_8701);
and U10876 (N_10876,N_9785,N_8305);
xor U10877 (N_10877,N_9661,N_8343);
xnor U10878 (N_10878,N_9749,N_8283);
nand U10879 (N_10879,N_9395,N_8326);
and U10880 (N_10880,N_9479,N_7942);
nand U10881 (N_10881,N_8039,N_8417);
and U10882 (N_10882,N_8929,N_9192);
nand U10883 (N_10883,N_7837,N_7961);
or U10884 (N_10884,N_9654,N_9616);
and U10885 (N_10885,N_9406,N_9380);
and U10886 (N_10886,N_8026,N_8295);
xnor U10887 (N_10887,N_7571,N_7880);
nor U10888 (N_10888,N_9002,N_9020);
or U10889 (N_10889,N_8266,N_8872);
and U10890 (N_10890,N_9063,N_7908);
and U10891 (N_10891,N_9168,N_7790);
and U10892 (N_10892,N_7755,N_8150);
nor U10893 (N_10893,N_9810,N_8824);
xor U10894 (N_10894,N_8850,N_7870);
xor U10895 (N_10895,N_9205,N_9439);
and U10896 (N_10896,N_8741,N_9537);
xor U10897 (N_10897,N_7849,N_9363);
nor U10898 (N_10898,N_8218,N_8013);
nand U10899 (N_10899,N_8583,N_8621);
and U10900 (N_10900,N_9743,N_8956);
nand U10901 (N_10901,N_8350,N_8736);
and U10902 (N_10902,N_7844,N_7862);
and U10903 (N_10903,N_8332,N_8780);
nor U10904 (N_10904,N_7703,N_9542);
or U10905 (N_10905,N_9791,N_8803);
or U10906 (N_10906,N_8840,N_9556);
or U10907 (N_10907,N_8991,N_8108);
nand U10908 (N_10908,N_7854,N_7917);
xor U10909 (N_10909,N_9480,N_9237);
nand U10910 (N_10910,N_8557,N_9336);
nor U10911 (N_10911,N_8544,N_9196);
nand U10912 (N_10912,N_7934,N_8016);
nor U10913 (N_10913,N_9225,N_9948);
or U10914 (N_10914,N_9428,N_9135);
or U10915 (N_10915,N_9206,N_7758);
and U10916 (N_10916,N_9456,N_8365);
or U10917 (N_10917,N_8260,N_9274);
and U10918 (N_10918,N_8176,N_7649);
and U10919 (N_10919,N_8155,N_9068);
or U10920 (N_10920,N_7600,N_8582);
nand U10921 (N_10921,N_8162,N_9518);
and U10922 (N_10922,N_7941,N_9936);
or U10923 (N_10923,N_8957,N_9122);
and U10924 (N_10924,N_9778,N_8489);
nand U10925 (N_10925,N_7502,N_9931);
nor U10926 (N_10926,N_9421,N_7723);
and U10927 (N_10927,N_8398,N_8694);
nor U10928 (N_10928,N_8234,N_8663);
nor U10929 (N_10929,N_8010,N_8433);
nand U10930 (N_10930,N_9645,N_8268);
nand U10931 (N_10931,N_7851,N_8132);
xor U10932 (N_10932,N_8340,N_8496);
nor U10933 (N_10933,N_9294,N_7522);
or U10934 (N_10934,N_8598,N_8945);
nor U10935 (N_10935,N_7989,N_9730);
nor U10936 (N_10936,N_9526,N_8187);
and U10937 (N_10937,N_9590,N_9664);
xnor U10938 (N_10938,N_7936,N_9315);
nor U10939 (N_10939,N_9686,N_8975);
nor U10940 (N_10940,N_9519,N_7568);
and U10941 (N_10941,N_8961,N_9399);
and U10942 (N_10942,N_8789,N_8682);
nand U10943 (N_10943,N_9543,N_9521);
nor U10944 (N_10944,N_8189,N_7800);
or U10945 (N_10945,N_9914,N_8201);
xnor U10946 (N_10946,N_9141,N_7805);
xnor U10947 (N_10947,N_7818,N_8566);
or U10948 (N_10948,N_8406,N_9455);
and U10949 (N_10949,N_8127,N_7661);
or U10950 (N_10950,N_8864,N_8490);
nand U10951 (N_10951,N_9902,N_7950);
xnor U10952 (N_10952,N_8331,N_9593);
and U10953 (N_10953,N_7547,N_8153);
xor U10954 (N_10954,N_8138,N_8488);
nor U10955 (N_10955,N_9359,N_8508);
and U10956 (N_10956,N_7789,N_8885);
nor U10957 (N_10957,N_9618,N_9889);
nor U10958 (N_10958,N_9229,N_8728);
xor U10959 (N_10959,N_9799,N_9120);
nor U10960 (N_10960,N_9833,N_8588);
or U10961 (N_10961,N_7737,N_8739);
or U10962 (N_10962,N_7531,N_9207);
and U10963 (N_10963,N_9201,N_9416);
or U10964 (N_10964,N_8586,N_8337);
or U10965 (N_10965,N_8556,N_9629);
nand U10966 (N_10966,N_8480,N_8759);
xnor U10967 (N_10967,N_8568,N_8667);
or U10968 (N_10968,N_9473,N_8799);
or U10969 (N_10969,N_7751,N_9760);
nor U10970 (N_10970,N_8329,N_9405);
nand U10971 (N_10971,N_7708,N_8873);
or U10972 (N_10972,N_8776,N_9090);
nor U10973 (N_10973,N_8608,N_8977);
or U10974 (N_10974,N_8672,N_9553);
nand U10975 (N_10975,N_9491,N_9441);
nor U10976 (N_10976,N_9678,N_9139);
or U10977 (N_10977,N_8721,N_8338);
nand U10978 (N_10978,N_9570,N_7554);
nand U10979 (N_10979,N_8397,N_9505);
nor U10980 (N_10980,N_9281,N_8920);
nor U10981 (N_10981,N_8248,N_8502);
nor U10982 (N_10982,N_9517,N_7896);
or U10983 (N_10983,N_8134,N_8252);
or U10984 (N_10984,N_7750,N_9828);
xnor U10985 (N_10985,N_9860,N_7759);
xnor U10986 (N_10986,N_8734,N_9815);
nand U10987 (N_10987,N_9886,N_9079);
nand U10988 (N_10988,N_7972,N_8058);
xor U10989 (N_10989,N_9202,N_9387);
or U10990 (N_10990,N_8805,N_9462);
and U10991 (N_10991,N_9300,N_8552);
nor U10992 (N_10992,N_9082,N_8681);
nand U10993 (N_10993,N_9489,N_8830);
xor U10994 (N_10994,N_8190,N_7747);
nand U10995 (N_10995,N_7956,N_7630);
nand U10996 (N_10996,N_9731,N_9254);
and U10997 (N_10997,N_8729,N_8897);
nor U10998 (N_10998,N_7905,N_7610);
xor U10999 (N_10999,N_8195,N_8535);
and U11000 (N_11000,N_9538,N_8930);
or U11001 (N_11001,N_9934,N_9039);
nand U11002 (N_11002,N_9154,N_8633);
nor U11003 (N_11003,N_9504,N_8110);
and U11004 (N_11004,N_7726,N_9197);
nor U11005 (N_11005,N_9469,N_7662);
or U11006 (N_11006,N_8988,N_9944);
xnor U11007 (N_11007,N_9475,N_8486);
and U11008 (N_11008,N_8760,N_8414);
and U11009 (N_11009,N_9032,N_8007);
xor U11010 (N_11010,N_9317,N_7566);
nand U11011 (N_11011,N_7537,N_7650);
nand U11012 (N_11012,N_8842,N_8386);
nor U11013 (N_11013,N_8596,N_7866);
or U11014 (N_11014,N_7597,N_7860);
or U11015 (N_11015,N_9769,N_9045);
nand U11016 (N_11016,N_9506,N_9796);
nand U11017 (N_11017,N_7716,N_9000);
nor U11018 (N_11018,N_8044,N_8816);
nor U11019 (N_11019,N_8019,N_8166);
or U11020 (N_11020,N_7959,N_8373);
and U11021 (N_11021,N_8495,N_9057);
or U11022 (N_11022,N_8989,N_8940);
nor U11023 (N_11023,N_7916,N_8362);
nor U11024 (N_11024,N_9575,N_9445);
nor U11025 (N_11025,N_9468,N_7868);
xnor U11026 (N_11026,N_8469,N_9916);
nor U11027 (N_11027,N_7754,N_9984);
nand U11028 (N_11028,N_7722,N_7631);
nor U11029 (N_11029,N_8244,N_8949);
and U11030 (N_11030,N_8844,N_8795);
xor U11031 (N_11031,N_8049,N_8831);
and U11032 (N_11032,N_7876,N_8676);
nand U11033 (N_11033,N_9036,N_8510);
nand U11034 (N_11034,N_9685,N_7828);
nor U11035 (N_11035,N_9798,N_9318);
nand U11036 (N_11036,N_7720,N_8318);
and U11037 (N_11037,N_9188,N_7947);
and U11038 (N_11038,N_9754,N_7546);
or U11039 (N_11039,N_8696,N_8562);
xnor U11040 (N_11040,N_8997,N_8429);
nor U11041 (N_11041,N_7528,N_7898);
or U11042 (N_11042,N_8745,N_7646);
nand U11043 (N_11043,N_9093,N_9985);
xor U11044 (N_11044,N_9744,N_9836);
and U11045 (N_11045,N_9338,N_8822);
xor U11046 (N_11046,N_9766,N_8434);
and U11047 (N_11047,N_8107,N_9394);
or U11048 (N_11048,N_7612,N_7745);
or U11049 (N_11049,N_9547,N_8931);
or U11050 (N_11050,N_9071,N_7738);
xor U11051 (N_11051,N_7743,N_8828);
and U11052 (N_11052,N_8916,N_8388);
and U11053 (N_11053,N_8175,N_8364);
or U11054 (N_11054,N_8008,N_9100);
nor U11055 (N_11055,N_9467,N_9013);
or U11056 (N_11056,N_9160,N_8498);
and U11057 (N_11057,N_7799,N_8883);
xnor U11058 (N_11058,N_9858,N_8788);
nor U11059 (N_11059,N_8096,N_8660);
nor U11060 (N_11060,N_7625,N_9748);
or U11061 (N_11061,N_9866,N_8069);
xnor U11062 (N_11062,N_8079,N_7842);
xnor U11063 (N_11063,N_9624,N_9502);
and U11064 (N_11064,N_9901,N_9028);
and U11065 (N_11065,N_8719,N_7873);
nand U11066 (N_11066,N_7734,N_9158);
or U11067 (N_11067,N_7806,N_9824);
nand U11068 (N_11068,N_8892,N_8317);
and U11069 (N_11069,N_8184,N_8781);
nand U11070 (N_11070,N_7886,N_8761);
and U11071 (N_11071,N_8448,N_9276);
or U11072 (N_11072,N_8641,N_7922);
and U11073 (N_11073,N_9813,N_7586);
xor U11074 (N_11074,N_8743,N_8866);
and U11075 (N_11075,N_9812,N_9878);
nor U11076 (N_11076,N_8990,N_9823);
or U11077 (N_11077,N_8915,N_8542);
or U11078 (N_11078,N_9617,N_7911);
or U11079 (N_11079,N_8670,N_7991);
or U11080 (N_11080,N_9747,N_9414);
nand U11081 (N_11081,N_9850,N_9389);
or U11082 (N_11082,N_9150,N_8395);
nor U11083 (N_11083,N_8631,N_9525);
xnor U11084 (N_11084,N_9582,N_9430);
nand U11085 (N_11085,N_7525,N_8591);
nor U11086 (N_11086,N_9800,N_9311);
nor U11087 (N_11087,N_9728,N_9656);
nor U11088 (N_11088,N_9918,N_9793);
xor U11089 (N_11089,N_7796,N_8909);
nand U11090 (N_11090,N_9026,N_9493);
nand U11091 (N_11091,N_7509,N_8888);
nand U11092 (N_11092,N_9746,N_7585);
nor U11093 (N_11093,N_8849,N_7994);
xor U11094 (N_11094,N_7604,N_9407);
or U11095 (N_11095,N_8585,N_8532);
xor U11096 (N_11096,N_8905,N_9369);
and U11097 (N_11097,N_9022,N_9367);
and U11098 (N_11098,N_7976,N_8425);
and U11099 (N_11099,N_8705,N_9133);
nor U11100 (N_11100,N_7617,N_8214);
and U11101 (N_11101,N_9295,N_8904);
and U11102 (N_11102,N_9652,N_9805);
nor U11103 (N_11103,N_8589,N_9146);
and U11104 (N_11104,N_8594,N_9284);
xor U11105 (N_11105,N_9408,N_8611);
nand U11106 (N_11106,N_8040,N_8028);
or U11107 (N_11107,N_9792,N_8066);
and U11108 (N_11108,N_8569,N_8202);
or U11109 (N_11109,N_8657,N_8693);
nand U11110 (N_11110,N_9231,N_9260);
xnor U11111 (N_11111,N_9847,N_8227);
and U11112 (N_11112,N_9786,N_7508);
xor U11113 (N_11113,N_7955,N_9927);
nand U11114 (N_11114,N_9436,N_9979);
nand U11115 (N_11115,N_9270,N_9107);
nand U11116 (N_11116,N_9581,N_9245);
nor U11117 (N_11117,N_8848,N_7813);
and U11118 (N_11118,N_7969,N_9470);
nand U11119 (N_11119,N_8944,N_8559);
or U11120 (N_11120,N_8135,N_9210);
nand U11121 (N_11121,N_9482,N_9639);
nand U11122 (N_11122,N_8389,N_9983);
nor U11123 (N_11123,N_9155,N_8186);
nor U11124 (N_11124,N_9966,N_9340);
or U11125 (N_11125,N_9142,N_8322);
nand U11126 (N_11126,N_8437,N_8907);
or U11127 (N_11127,N_9662,N_8203);
or U11128 (N_11128,N_9224,N_9322);
and U11129 (N_11129,N_7975,N_7591);
or U11130 (N_11130,N_7992,N_8964);
xor U11131 (N_11131,N_9598,N_9252);
and U11132 (N_11132,N_8062,N_9362);
or U11133 (N_11133,N_8271,N_7938);
nand U11134 (N_11134,N_8142,N_8359);
nand U11135 (N_11135,N_8297,N_8255);
nor U11136 (N_11136,N_8796,N_8775);
nand U11137 (N_11137,N_9089,N_9223);
nor U11138 (N_11138,N_9682,N_7887);
nand U11139 (N_11139,N_9676,N_8506);
or U11140 (N_11140,N_8167,N_7826);
and U11141 (N_11141,N_9725,N_9238);
nand U11142 (N_11142,N_8484,N_9970);
nand U11143 (N_11143,N_8555,N_8080);
xnor U11144 (N_11144,N_9474,N_8610);
xor U11145 (N_11145,N_7685,N_7511);
xor U11146 (N_11146,N_9613,N_7910);
and U11147 (N_11147,N_8620,N_9990);
nand U11148 (N_11148,N_8960,N_7921);
and U11149 (N_11149,N_8463,N_8303);
nor U11150 (N_11150,N_9715,N_8526);
nand U11151 (N_11151,N_8876,N_8671);
xnor U11152 (N_11152,N_8505,N_9615);
nor U11153 (N_11153,N_7577,N_8757);
or U11154 (N_11154,N_9588,N_7993);
and U11155 (N_11155,N_8497,N_9111);
and U11156 (N_11156,N_8958,N_9173);
xor U11157 (N_11157,N_9511,N_8470);
and U11158 (N_11158,N_9987,N_9217);
and U11159 (N_11159,N_9846,N_8984);
xor U11160 (N_11160,N_9091,N_8863);
or U11161 (N_11161,N_9251,N_9779);
xnor U11162 (N_11162,N_9756,N_8908);
and U11163 (N_11163,N_8221,N_9527);
or U11164 (N_11164,N_7609,N_7890);
and U11165 (N_11165,N_7656,N_9145);
and U11166 (N_11166,N_8174,N_9693);
or U11167 (N_11167,N_9690,N_9601);
xor U11168 (N_11168,N_8709,N_8151);
or U11169 (N_11169,N_7777,N_8253);
or U11170 (N_11170,N_8078,N_7698);
or U11171 (N_11171,N_7593,N_9176);
or U11172 (N_11172,N_9065,N_7775);
nor U11173 (N_11173,N_9242,N_8718);
or U11174 (N_11174,N_8456,N_9977);
nor U11175 (N_11175,N_9691,N_9864);
xnor U11176 (N_11176,N_8771,N_9127);
xnor U11177 (N_11177,N_9383,N_8355);
and U11178 (N_11178,N_8121,N_8210);
and U11179 (N_11179,N_8455,N_9826);
or U11180 (N_11180,N_9751,N_8137);
and U11181 (N_11181,N_8294,N_9882);
or U11182 (N_11182,N_7906,N_8067);
and U11183 (N_11183,N_8769,N_8901);
or U11184 (N_11184,N_9651,N_9585);
or U11185 (N_11185,N_8421,N_8291);
or U11186 (N_11186,N_9720,N_9309);
xnor U11187 (N_11187,N_9056,N_8874);
nand U11188 (N_11188,N_9157,N_9713);
nor U11189 (N_11189,N_8595,N_9331);
xor U11190 (N_11190,N_9337,N_9589);
and U11191 (N_11191,N_8306,N_9030);
or U11192 (N_11192,N_8606,N_7695);
or U11193 (N_11193,N_7856,N_9594);
and U11194 (N_11194,N_9612,N_9361);
nor U11195 (N_11195,N_7534,N_9472);
or U11196 (N_11196,N_9212,N_7881);
and U11197 (N_11197,N_9529,N_8948);
or U11198 (N_11198,N_7668,N_9083);
xor U11199 (N_11199,N_9702,N_9162);
and U11200 (N_11200,N_7995,N_7603);
nand U11201 (N_11201,N_9014,N_8884);
xnor U11202 (N_11202,N_8207,N_9959);
xor U11203 (N_11203,N_8982,N_8112);
xor U11204 (N_11204,N_7764,N_8756);
or U11205 (N_11205,N_9478,N_9312);
or U11206 (N_11206,N_8548,N_9187);
and U11207 (N_11207,N_8213,N_7791);
and U11208 (N_11208,N_9557,N_8323);
and U11209 (N_11209,N_8652,N_9130);
xnor U11210 (N_11210,N_7735,N_9717);
and U11211 (N_11211,N_7526,N_9958);
xnor U11212 (N_11212,N_8735,N_8346);
or U11213 (N_11213,N_7573,N_8779);
or U11214 (N_11214,N_9872,N_9149);
and U11215 (N_11215,N_9325,N_9165);
and U11216 (N_11216,N_8612,N_7684);
xnor U11217 (N_11217,N_9326,N_9665);
or U11218 (N_11218,N_8133,N_8571);
nand U11219 (N_11219,N_8168,N_7933);
and U11220 (N_11220,N_9930,N_8279);
or U11221 (N_11221,N_7595,N_8208);
nand U11222 (N_11222,N_7878,N_7613);
xor U11223 (N_11223,N_9023,N_9488);
xor U11224 (N_11224,N_9448,N_7852);
nor U11225 (N_11225,N_7925,N_8009);
or U11226 (N_11226,N_8602,N_9689);
nor U11227 (N_11227,N_9465,N_9592);
nor U11228 (N_11228,N_7971,N_8475);
or U11229 (N_11229,N_9564,N_9498);
or U11230 (N_11230,N_9995,N_9264);
nand U11231 (N_11231,N_9816,N_9602);
or U11232 (N_11232,N_9814,N_8241);
nand U11233 (N_11233,N_7686,N_9906);
and U11234 (N_11234,N_9929,N_9347);
or U11235 (N_11235,N_9669,N_7927);
nor U11236 (N_11236,N_8817,N_8431);
nand U11237 (N_11237,N_9454,N_7579);
nand U11238 (N_11238,N_9259,N_7857);
nand U11239 (N_11239,N_9572,N_8461);
nand U11240 (N_11240,N_9832,N_8616);
nand U11241 (N_11241,N_8199,N_9350);
xnor U11242 (N_11242,N_8551,N_8898);
or U11243 (N_11243,N_8179,N_9417);
nor U11244 (N_11244,N_7774,N_9372);
nand U11245 (N_11245,N_7619,N_8440);
xnor U11246 (N_11246,N_8746,N_8751);
xor U11247 (N_11247,N_9674,N_9993);
and U11248 (N_11248,N_7677,N_8707);
xnor U11249 (N_11249,N_9838,N_7749);
nand U11250 (N_11250,N_9822,N_9608);
and U11251 (N_11251,N_8243,N_8136);
and U11252 (N_11252,N_9945,N_7938);
and U11253 (N_11253,N_7538,N_8842);
and U11254 (N_11254,N_7670,N_7797);
or U11255 (N_11255,N_9507,N_8265);
nand U11256 (N_11256,N_9063,N_8231);
and U11257 (N_11257,N_9008,N_8470);
xor U11258 (N_11258,N_7846,N_8304);
xnor U11259 (N_11259,N_8541,N_8577);
xnor U11260 (N_11260,N_9528,N_9361);
nand U11261 (N_11261,N_9087,N_8787);
or U11262 (N_11262,N_9088,N_9407);
or U11263 (N_11263,N_8960,N_9588);
xor U11264 (N_11264,N_8806,N_7691);
and U11265 (N_11265,N_7753,N_8583);
nand U11266 (N_11266,N_9307,N_7668);
nand U11267 (N_11267,N_8112,N_8797);
and U11268 (N_11268,N_7564,N_7965);
or U11269 (N_11269,N_7594,N_8324);
or U11270 (N_11270,N_9169,N_8025);
nand U11271 (N_11271,N_8938,N_9662);
xor U11272 (N_11272,N_9218,N_8686);
or U11273 (N_11273,N_7812,N_9640);
nand U11274 (N_11274,N_7657,N_9883);
or U11275 (N_11275,N_8207,N_8456);
nand U11276 (N_11276,N_8634,N_9178);
and U11277 (N_11277,N_7530,N_8355);
xnor U11278 (N_11278,N_9247,N_7903);
nor U11279 (N_11279,N_9332,N_9844);
and U11280 (N_11280,N_8133,N_8290);
and U11281 (N_11281,N_7520,N_7562);
or U11282 (N_11282,N_9195,N_7994);
or U11283 (N_11283,N_7527,N_7978);
or U11284 (N_11284,N_8400,N_7538);
and U11285 (N_11285,N_8147,N_9222);
or U11286 (N_11286,N_9025,N_7594);
nor U11287 (N_11287,N_8848,N_8598);
nor U11288 (N_11288,N_7745,N_9008);
and U11289 (N_11289,N_8949,N_7672);
or U11290 (N_11290,N_8762,N_8390);
and U11291 (N_11291,N_9827,N_8152);
xnor U11292 (N_11292,N_8999,N_7635);
nor U11293 (N_11293,N_8889,N_9831);
xor U11294 (N_11294,N_8026,N_9338);
or U11295 (N_11295,N_8226,N_9897);
nor U11296 (N_11296,N_8617,N_8819);
and U11297 (N_11297,N_9904,N_8505);
nand U11298 (N_11298,N_8556,N_9749);
nand U11299 (N_11299,N_8273,N_9837);
nor U11300 (N_11300,N_7503,N_9911);
or U11301 (N_11301,N_9677,N_9197);
and U11302 (N_11302,N_9505,N_8738);
nor U11303 (N_11303,N_8408,N_9973);
or U11304 (N_11304,N_9388,N_8739);
or U11305 (N_11305,N_7982,N_9699);
nor U11306 (N_11306,N_7989,N_7549);
and U11307 (N_11307,N_8521,N_8398);
xnor U11308 (N_11308,N_8289,N_9733);
xor U11309 (N_11309,N_8256,N_9956);
or U11310 (N_11310,N_9715,N_8070);
and U11311 (N_11311,N_9072,N_9499);
and U11312 (N_11312,N_8961,N_8002);
or U11313 (N_11313,N_9318,N_7639);
or U11314 (N_11314,N_7846,N_8091);
nor U11315 (N_11315,N_8387,N_9566);
xor U11316 (N_11316,N_8467,N_8994);
and U11317 (N_11317,N_9063,N_9867);
nor U11318 (N_11318,N_7868,N_9609);
or U11319 (N_11319,N_7994,N_8893);
and U11320 (N_11320,N_7713,N_9191);
or U11321 (N_11321,N_9322,N_8241);
or U11322 (N_11322,N_7746,N_8980);
and U11323 (N_11323,N_9571,N_8611);
or U11324 (N_11324,N_7766,N_9200);
nor U11325 (N_11325,N_7520,N_8481);
or U11326 (N_11326,N_8352,N_7914);
nand U11327 (N_11327,N_8580,N_9712);
and U11328 (N_11328,N_8901,N_7986);
and U11329 (N_11329,N_8399,N_8573);
nor U11330 (N_11330,N_9584,N_8116);
xor U11331 (N_11331,N_9893,N_8296);
and U11332 (N_11332,N_7661,N_7962);
xor U11333 (N_11333,N_9925,N_8664);
nand U11334 (N_11334,N_8489,N_9197);
and U11335 (N_11335,N_8240,N_9422);
nand U11336 (N_11336,N_8292,N_8676);
and U11337 (N_11337,N_9075,N_9789);
and U11338 (N_11338,N_9848,N_8243);
xnor U11339 (N_11339,N_9496,N_9097);
nor U11340 (N_11340,N_9794,N_8881);
and U11341 (N_11341,N_8409,N_7664);
nand U11342 (N_11342,N_9735,N_8086);
xnor U11343 (N_11343,N_9706,N_9399);
xnor U11344 (N_11344,N_8565,N_8722);
or U11345 (N_11345,N_9666,N_8042);
and U11346 (N_11346,N_9427,N_9123);
nand U11347 (N_11347,N_7909,N_9418);
xnor U11348 (N_11348,N_8059,N_7742);
nor U11349 (N_11349,N_9995,N_8680);
xor U11350 (N_11350,N_8050,N_9049);
nor U11351 (N_11351,N_7745,N_8259);
nand U11352 (N_11352,N_9133,N_9225);
nand U11353 (N_11353,N_9476,N_8321);
xor U11354 (N_11354,N_9645,N_7599);
or U11355 (N_11355,N_7914,N_8685);
and U11356 (N_11356,N_8754,N_8350);
nor U11357 (N_11357,N_7757,N_7996);
nand U11358 (N_11358,N_7970,N_9184);
nand U11359 (N_11359,N_9563,N_8064);
nand U11360 (N_11360,N_8462,N_9052);
or U11361 (N_11361,N_9813,N_7842);
and U11362 (N_11362,N_9670,N_8314);
and U11363 (N_11363,N_8831,N_9546);
or U11364 (N_11364,N_8018,N_9780);
nor U11365 (N_11365,N_8077,N_7572);
nor U11366 (N_11366,N_9756,N_9310);
xnor U11367 (N_11367,N_8702,N_7992);
or U11368 (N_11368,N_8702,N_9184);
and U11369 (N_11369,N_9678,N_8057);
and U11370 (N_11370,N_8357,N_9079);
or U11371 (N_11371,N_9947,N_9168);
nand U11372 (N_11372,N_8545,N_9430);
or U11373 (N_11373,N_9399,N_9370);
nand U11374 (N_11374,N_8503,N_8977);
or U11375 (N_11375,N_8646,N_8877);
nor U11376 (N_11376,N_9988,N_8487);
and U11377 (N_11377,N_8024,N_8481);
nand U11378 (N_11378,N_9948,N_9817);
nor U11379 (N_11379,N_9215,N_8531);
or U11380 (N_11380,N_9785,N_9862);
nor U11381 (N_11381,N_9806,N_8129);
and U11382 (N_11382,N_7911,N_7975);
xor U11383 (N_11383,N_7805,N_7687);
or U11384 (N_11384,N_8161,N_9814);
or U11385 (N_11385,N_8145,N_9479);
and U11386 (N_11386,N_8486,N_7588);
xor U11387 (N_11387,N_8739,N_7944);
nand U11388 (N_11388,N_8700,N_8514);
xnor U11389 (N_11389,N_8392,N_9923);
or U11390 (N_11390,N_9210,N_9546);
xnor U11391 (N_11391,N_7977,N_7737);
xor U11392 (N_11392,N_8845,N_8707);
nand U11393 (N_11393,N_9479,N_7720);
or U11394 (N_11394,N_8973,N_7822);
xnor U11395 (N_11395,N_8912,N_9484);
nand U11396 (N_11396,N_8876,N_8531);
or U11397 (N_11397,N_7945,N_7525);
nor U11398 (N_11398,N_8109,N_7515);
nand U11399 (N_11399,N_9786,N_8299);
nor U11400 (N_11400,N_9718,N_9924);
xnor U11401 (N_11401,N_8866,N_8827);
xor U11402 (N_11402,N_7717,N_8877);
and U11403 (N_11403,N_7891,N_9079);
or U11404 (N_11404,N_7561,N_9005);
nor U11405 (N_11405,N_8303,N_7648);
nand U11406 (N_11406,N_8548,N_8723);
and U11407 (N_11407,N_9492,N_8618);
or U11408 (N_11408,N_7728,N_8517);
xor U11409 (N_11409,N_8244,N_7869);
nor U11410 (N_11410,N_8189,N_9472);
and U11411 (N_11411,N_8312,N_9306);
nand U11412 (N_11412,N_7897,N_7765);
and U11413 (N_11413,N_8462,N_9228);
nor U11414 (N_11414,N_9961,N_8540);
xnor U11415 (N_11415,N_9637,N_9589);
xor U11416 (N_11416,N_9042,N_7614);
and U11417 (N_11417,N_9946,N_8212);
and U11418 (N_11418,N_8803,N_7891);
or U11419 (N_11419,N_9453,N_9685);
and U11420 (N_11420,N_9957,N_9417);
xnor U11421 (N_11421,N_8706,N_7827);
xnor U11422 (N_11422,N_8838,N_7809);
or U11423 (N_11423,N_9187,N_8996);
nand U11424 (N_11424,N_9782,N_9745);
nand U11425 (N_11425,N_7917,N_7927);
and U11426 (N_11426,N_8747,N_9687);
nor U11427 (N_11427,N_8116,N_7927);
nor U11428 (N_11428,N_7575,N_9875);
nor U11429 (N_11429,N_9528,N_8830);
and U11430 (N_11430,N_8115,N_8264);
nand U11431 (N_11431,N_8620,N_7730);
and U11432 (N_11432,N_7574,N_8368);
xnor U11433 (N_11433,N_8260,N_8291);
or U11434 (N_11434,N_9551,N_9323);
and U11435 (N_11435,N_9630,N_8294);
and U11436 (N_11436,N_8299,N_9062);
and U11437 (N_11437,N_9426,N_8336);
and U11438 (N_11438,N_8545,N_8669);
nor U11439 (N_11439,N_9161,N_9087);
and U11440 (N_11440,N_8351,N_9061);
xnor U11441 (N_11441,N_8577,N_8552);
or U11442 (N_11442,N_8492,N_8739);
nand U11443 (N_11443,N_7635,N_8291);
and U11444 (N_11444,N_7563,N_9572);
nand U11445 (N_11445,N_8626,N_8513);
xor U11446 (N_11446,N_9392,N_9044);
nor U11447 (N_11447,N_9096,N_7684);
nand U11448 (N_11448,N_9285,N_7916);
and U11449 (N_11449,N_9594,N_7557);
and U11450 (N_11450,N_7517,N_8606);
and U11451 (N_11451,N_8957,N_7520);
xnor U11452 (N_11452,N_9168,N_9679);
and U11453 (N_11453,N_7918,N_9241);
or U11454 (N_11454,N_9222,N_9149);
xor U11455 (N_11455,N_8256,N_7911);
and U11456 (N_11456,N_9912,N_9367);
nor U11457 (N_11457,N_7783,N_8142);
or U11458 (N_11458,N_7792,N_7982);
xor U11459 (N_11459,N_9800,N_7647);
or U11460 (N_11460,N_8478,N_9138);
nor U11461 (N_11461,N_9788,N_9806);
nor U11462 (N_11462,N_9405,N_7581);
and U11463 (N_11463,N_9985,N_9605);
and U11464 (N_11464,N_7548,N_8063);
xor U11465 (N_11465,N_9612,N_9831);
and U11466 (N_11466,N_7881,N_8253);
nand U11467 (N_11467,N_8938,N_9344);
nor U11468 (N_11468,N_9479,N_8228);
xor U11469 (N_11469,N_7683,N_9985);
xor U11470 (N_11470,N_7552,N_8526);
nor U11471 (N_11471,N_8857,N_8004);
or U11472 (N_11472,N_9553,N_9046);
nand U11473 (N_11473,N_7724,N_7957);
nor U11474 (N_11474,N_8392,N_8820);
and U11475 (N_11475,N_8661,N_8210);
xnor U11476 (N_11476,N_9012,N_9167);
nand U11477 (N_11477,N_8278,N_8938);
or U11478 (N_11478,N_8961,N_9094);
xor U11479 (N_11479,N_9162,N_9300);
or U11480 (N_11480,N_8380,N_9467);
and U11481 (N_11481,N_9036,N_9641);
xnor U11482 (N_11482,N_7539,N_9994);
xnor U11483 (N_11483,N_7687,N_8717);
xor U11484 (N_11484,N_7791,N_7717);
nor U11485 (N_11485,N_7849,N_9076);
nor U11486 (N_11486,N_9797,N_9204);
and U11487 (N_11487,N_8721,N_8283);
or U11488 (N_11488,N_9170,N_7800);
nor U11489 (N_11489,N_9792,N_8448);
nand U11490 (N_11490,N_9150,N_7783);
and U11491 (N_11491,N_7508,N_9317);
nand U11492 (N_11492,N_9852,N_7653);
and U11493 (N_11493,N_8734,N_7746);
and U11494 (N_11494,N_7900,N_7510);
nor U11495 (N_11495,N_7700,N_8744);
xnor U11496 (N_11496,N_9206,N_8309);
xor U11497 (N_11497,N_7999,N_9683);
or U11498 (N_11498,N_7613,N_9916);
nand U11499 (N_11499,N_9488,N_9656);
nand U11500 (N_11500,N_7678,N_9126);
xor U11501 (N_11501,N_8016,N_8404);
or U11502 (N_11502,N_9523,N_9080);
nand U11503 (N_11503,N_9381,N_9146);
nor U11504 (N_11504,N_8345,N_8204);
or U11505 (N_11505,N_7974,N_8335);
xor U11506 (N_11506,N_9902,N_9583);
and U11507 (N_11507,N_9234,N_9450);
nor U11508 (N_11508,N_9728,N_7794);
xor U11509 (N_11509,N_8774,N_8924);
xor U11510 (N_11510,N_9370,N_9710);
and U11511 (N_11511,N_8997,N_8043);
nand U11512 (N_11512,N_8792,N_8133);
xnor U11513 (N_11513,N_8057,N_9573);
nor U11514 (N_11514,N_7875,N_8051);
or U11515 (N_11515,N_7967,N_8197);
nand U11516 (N_11516,N_9025,N_7502);
xnor U11517 (N_11517,N_7589,N_9004);
and U11518 (N_11518,N_7999,N_7570);
or U11519 (N_11519,N_9401,N_8015);
nor U11520 (N_11520,N_7568,N_7984);
xor U11521 (N_11521,N_8988,N_9249);
and U11522 (N_11522,N_9004,N_7632);
or U11523 (N_11523,N_7984,N_8079);
nor U11524 (N_11524,N_8382,N_9388);
or U11525 (N_11525,N_9554,N_8070);
nor U11526 (N_11526,N_8706,N_9369);
xor U11527 (N_11527,N_7525,N_8588);
or U11528 (N_11528,N_7764,N_8071);
nor U11529 (N_11529,N_8748,N_9916);
xor U11530 (N_11530,N_9503,N_8918);
nor U11531 (N_11531,N_9922,N_9300);
and U11532 (N_11532,N_8271,N_7586);
xnor U11533 (N_11533,N_8125,N_7999);
or U11534 (N_11534,N_7561,N_7793);
nand U11535 (N_11535,N_9829,N_8098);
and U11536 (N_11536,N_7623,N_9349);
nand U11537 (N_11537,N_7625,N_8155);
and U11538 (N_11538,N_9381,N_8517);
nor U11539 (N_11539,N_8680,N_8889);
and U11540 (N_11540,N_9006,N_8687);
xnor U11541 (N_11541,N_8234,N_9575);
nand U11542 (N_11542,N_8605,N_8556);
xor U11543 (N_11543,N_8006,N_8063);
xor U11544 (N_11544,N_9481,N_8540);
xor U11545 (N_11545,N_9691,N_7673);
nor U11546 (N_11546,N_9106,N_8767);
nand U11547 (N_11547,N_8587,N_8969);
xor U11548 (N_11548,N_7774,N_7914);
xnor U11549 (N_11549,N_9052,N_8231);
or U11550 (N_11550,N_8066,N_8574);
xnor U11551 (N_11551,N_9082,N_8986);
nand U11552 (N_11552,N_8908,N_8544);
nand U11553 (N_11553,N_7510,N_7700);
or U11554 (N_11554,N_8964,N_7756);
or U11555 (N_11555,N_8934,N_8717);
and U11556 (N_11556,N_9577,N_8368);
and U11557 (N_11557,N_7847,N_8416);
xor U11558 (N_11558,N_8612,N_9925);
and U11559 (N_11559,N_8158,N_8875);
or U11560 (N_11560,N_8296,N_7968);
xnor U11561 (N_11561,N_9048,N_7727);
nor U11562 (N_11562,N_9436,N_7731);
nand U11563 (N_11563,N_9544,N_7531);
nor U11564 (N_11564,N_9128,N_7654);
nand U11565 (N_11565,N_9036,N_8699);
xnor U11566 (N_11566,N_9709,N_7549);
nand U11567 (N_11567,N_7590,N_9672);
or U11568 (N_11568,N_7673,N_9877);
nand U11569 (N_11569,N_8878,N_7721);
or U11570 (N_11570,N_8604,N_9652);
and U11571 (N_11571,N_9084,N_9053);
nor U11572 (N_11572,N_8093,N_9215);
xor U11573 (N_11573,N_9285,N_9957);
xor U11574 (N_11574,N_9247,N_9061);
nor U11575 (N_11575,N_7516,N_8303);
nand U11576 (N_11576,N_9860,N_9479);
xor U11577 (N_11577,N_7859,N_8568);
xor U11578 (N_11578,N_9863,N_9537);
and U11579 (N_11579,N_8104,N_7576);
xor U11580 (N_11580,N_8644,N_8010);
or U11581 (N_11581,N_9726,N_9877);
nor U11582 (N_11582,N_9473,N_8848);
or U11583 (N_11583,N_9750,N_8440);
nand U11584 (N_11584,N_8126,N_8907);
nor U11585 (N_11585,N_7630,N_9111);
xnor U11586 (N_11586,N_8863,N_7905);
nor U11587 (N_11587,N_8251,N_8930);
xnor U11588 (N_11588,N_8978,N_7773);
nor U11589 (N_11589,N_9255,N_7618);
nand U11590 (N_11590,N_8075,N_9071);
and U11591 (N_11591,N_8728,N_8975);
xor U11592 (N_11592,N_9226,N_9895);
and U11593 (N_11593,N_9420,N_7929);
nand U11594 (N_11594,N_9134,N_8780);
nor U11595 (N_11595,N_8229,N_9289);
and U11596 (N_11596,N_7650,N_8390);
or U11597 (N_11597,N_9098,N_8889);
and U11598 (N_11598,N_8733,N_7558);
and U11599 (N_11599,N_8757,N_8192);
nand U11600 (N_11600,N_7504,N_9887);
nand U11601 (N_11601,N_8549,N_7815);
or U11602 (N_11602,N_9369,N_9968);
or U11603 (N_11603,N_7858,N_7547);
nand U11604 (N_11604,N_8041,N_9597);
nor U11605 (N_11605,N_8030,N_7534);
and U11606 (N_11606,N_8826,N_9069);
or U11607 (N_11607,N_7597,N_9408);
nand U11608 (N_11608,N_7587,N_8901);
and U11609 (N_11609,N_9774,N_8569);
nor U11610 (N_11610,N_9518,N_8075);
nand U11611 (N_11611,N_9411,N_9472);
nor U11612 (N_11612,N_9114,N_9126);
and U11613 (N_11613,N_9907,N_9986);
nor U11614 (N_11614,N_8387,N_7612);
nand U11615 (N_11615,N_7719,N_9421);
xnor U11616 (N_11616,N_9846,N_9700);
xnor U11617 (N_11617,N_8885,N_7962);
or U11618 (N_11618,N_8292,N_9110);
nand U11619 (N_11619,N_7635,N_9666);
or U11620 (N_11620,N_8398,N_7893);
nand U11621 (N_11621,N_9820,N_9290);
nand U11622 (N_11622,N_7759,N_9069);
and U11623 (N_11623,N_9183,N_8233);
xnor U11624 (N_11624,N_9176,N_9975);
nand U11625 (N_11625,N_8257,N_8508);
or U11626 (N_11626,N_8754,N_7893);
nor U11627 (N_11627,N_8670,N_8354);
xnor U11628 (N_11628,N_9202,N_9592);
or U11629 (N_11629,N_8365,N_8578);
nand U11630 (N_11630,N_9433,N_8966);
nor U11631 (N_11631,N_9042,N_8289);
or U11632 (N_11632,N_9992,N_8521);
and U11633 (N_11633,N_9191,N_9394);
xnor U11634 (N_11634,N_9488,N_9332);
nor U11635 (N_11635,N_7633,N_9094);
nor U11636 (N_11636,N_8521,N_9463);
nand U11637 (N_11637,N_9857,N_8684);
nand U11638 (N_11638,N_7914,N_9403);
xnor U11639 (N_11639,N_8719,N_8823);
and U11640 (N_11640,N_8931,N_7825);
and U11641 (N_11641,N_8004,N_7899);
nor U11642 (N_11642,N_9829,N_9217);
nor U11643 (N_11643,N_8759,N_8733);
xor U11644 (N_11644,N_9745,N_9734);
xnor U11645 (N_11645,N_9233,N_9831);
xnor U11646 (N_11646,N_9746,N_9448);
or U11647 (N_11647,N_7717,N_8523);
xnor U11648 (N_11648,N_8579,N_8409);
or U11649 (N_11649,N_8279,N_8462);
or U11650 (N_11650,N_8264,N_7911);
nor U11651 (N_11651,N_8773,N_9080);
nor U11652 (N_11652,N_8524,N_9301);
and U11653 (N_11653,N_8180,N_9495);
nor U11654 (N_11654,N_8595,N_8325);
xnor U11655 (N_11655,N_9337,N_8114);
and U11656 (N_11656,N_8580,N_9269);
nand U11657 (N_11657,N_9832,N_9417);
or U11658 (N_11658,N_9103,N_9728);
and U11659 (N_11659,N_7633,N_8323);
nor U11660 (N_11660,N_9359,N_9487);
and U11661 (N_11661,N_9370,N_8574);
nor U11662 (N_11662,N_9294,N_7797);
or U11663 (N_11663,N_9584,N_8808);
nand U11664 (N_11664,N_9553,N_9356);
nand U11665 (N_11665,N_8079,N_9128);
and U11666 (N_11666,N_7790,N_9575);
nand U11667 (N_11667,N_8831,N_8106);
nor U11668 (N_11668,N_8538,N_9112);
and U11669 (N_11669,N_9591,N_8947);
or U11670 (N_11670,N_8012,N_8943);
xnor U11671 (N_11671,N_9062,N_9597);
xor U11672 (N_11672,N_8485,N_8068);
nand U11673 (N_11673,N_9709,N_8127);
and U11674 (N_11674,N_9676,N_9927);
or U11675 (N_11675,N_7779,N_9027);
and U11676 (N_11676,N_8195,N_8450);
nand U11677 (N_11677,N_7824,N_9809);
or U11678 (N_11678,N_9088,N_9331);
nand U11679 (N_11679,N_9170,N_8389);
nor U11680 (N_11680,N_8095,N_9593);
nand U11681 (N_11681,N_8153,N_9163);
and U11682 (N_11682,N_9717,N_9048);
nand U11683 (N_11683,N_8452,N_7692);
nor U11684 (N_11684,N_9216,N_8996);
nand U11685 (N_11685,N_8860,N_9468);
and U11686 (N_11686,N_9731,N_9305);
nand U11687 (N_11687,N_9766,N_8020);
and U11688 (N_11688,N_9114,N_9480);
nand U11689 (N_11689,N_8804,N_7858);
xnor U11690 (N_11690,N_8687,N_8929);
xor U11691 (N_11691,N_9921,N_8819);
xor U11692 (N_11692,N_8968,N_9360);
or U11693 (N_11693,N_8628,N_8723);
and U11694 (N_11694,N_9887,N_7558);
nor U11695 (N_11695,N_8066,N_8455);
nand U11696 (N_11696,N_8091,N_8942);
xnor U11697 (N_11697,N_9331,N_8680);
or U11698 (N_11698,N_8041,N_9658);
or U11699 (N_11699,N_9731,N_7918);
xor U11700 (N_11700,N_9030,N_8726);
nor U11701 (N_11701,N_8178,N_9871);
or U11702 (N_11702,N_9809,N_8576);
nand U11703 (N_11703,N_9793,N_9798);
and U11704 (N_11704,N_9387,N_8223);
nor U11705 (N_11705,N_9086,N_9731);
and U11706 (N_11706,N_7854,N_8023);
xnor U11707 (N_11707,N_9437,N_8285);
nand U11708 (N_11708,N_9784,N_9533);
nor U11709 (N_11709,N_8559,N_8808);
nand U11710 (N_11710,N_7803,N_8681);
nor U11711 (N_11711,N_8965,N_8132);
xnor U11712 (N_11712,N_8533,N_7654);
xor U11713 (N_11713,N_8158,N_8642);
and U11714 (N_11714,N_9429,N_7546);
and U11715 (N_11715,N_7501,N_8417);
xor U11716 (N_11716,N_9133,N_8579);
or U11717 (N_11717,N_8437,N_8281);
xor U11718 (N_11718,N_7740,N_9253);
xnor U11719 (N_11719,N_8363,N_9563);
nand U11720 (N_11720,N_8559,N_8590);
nor U11721 (N_11721,N_8754,N_8610);
and U11722 (N_11722,N_9573,N_9328);
or U11723 (N_11723,N_9278,N_9609);
nor U11724 (N_11724,N_8835,N_7827);
nor U11725 (N_11725,N_8105,N_9765);
or U11726 (N_11726,N_9121,N_8344);
xor U11727 (N_11727,N_9491,N_8440);
nor U11728 (N_11728,N_9101,N_8169);
nor U11729 (N_11729,N_8897,N_9667);
or U11730 (N_11730,N_8106,N_8094);
nor U11731 (N_11731,N_9843,N_9177);
or U11732 (N_11732,N_9562,N_9478);
or U11733 (N_11733,N_8154,N_7535);
and U11734 (N_11734,N_8907,N_9709);
nand U11735 (N_11735,N_9234,N_8248);
nor U11736 (N_11736,N_7629,N_7519);
or U11737 (N_11737,N_9578,N_7689);
and U11738 (N_11738,N_8419,N_8052);
nor U11739 (N_11739,N_8829,N_7780);
nand U11740 (N_11740,N_9740,N_7843);
or U11741 (N_11741,N_8106,N_9875);
and U11742 (N_11742,N_9630,N_8467);
or U11743 (N_11743,N_8899,N_9057);
xor U11744 (N_11744,N_9588,N_8731);
and U11745 (N_11745,N_8967,N_7503);
nor U11746 (N_11746,N_8696,N_7551);
or U11747 (N_11747,N_8643,N_8236);
and U11748 (N_11748,N_8375,N_7859);
and U11749 (N_11749,N_8494,N_9360);
xor U11750 (N_11750,N_8881,N_7837);
xnor U11751 (N_11751,N_9302,N_8861);
or U11752 (N_11752,N_9971,N_9865);
or U11753 (N_11753,N_9786,N_9522);
nor U11754 (N_11754,N_8400,N_8956);
nand U11755 (N_11755,N_9660,N_8844);
or U11756 (N_11756,N_7808,N_9933);
nor U11757 (N_11757,N_7720,N_8277);
and U11758 (N_11758,N_9730,N_9316);
and U11759 (N_11759,N_8586,N_9878);
or U11760 (N_11760,N_8455,N_8128);
nand U11761 (N_11761,N_7897,N_8958);
xor U11762 (N_11762,N_9353,N_8875);
or U11763 (N_11763,N_8474,N_7775);
xor U11764 (N_11764,N_7696,N_9280);
and U11765 (N_11765,N_7992,N_8229);
nand U11766 (N_11766,N_8672,N_7710);
nand U11767 (N_11767,N_9505,N_7500);
and U11768 (N_11768,N_7650,N_9411);
nand U11769 (N_11769,N_9275,N_9980);
and U11770 (N_11770,N_9059,N_9038);
and U11771 (N_11771,N_9674,N_8237);
nor U11772 (N_11772,N_9053,N_8127);
nor U11773 (N_11773,N_8702,N_7654);
nand U11774 (N_11774,N_9009,N_8872);
and U11775 (N_11775,N_8442,N_9958);
and U11776 (N_11776,N_9865,N_9177);
nand U11777 (N_11777,N_7888,N_7664);
xor U11778 (N_11778,N_7981,N_9441);
nor U11779 (N_11779,N_9695,N_9587);
nor U11780 (N_11780,N_8447,N_9727);
xor U11781 (N_11781,N_9081,N_9824);
xor U11782 (N_11782,N_9860,N_8282);
nor U11783 (N_11783,N_9831,N_8998);
or U11784 (N_11784,N_7875,N_9424);
nand U11785 (N_11785,N_8685,N_8028);
or U11786 (N_11786,N_9925,N_8376);
or U11787 (N_11787,N_8944,N_9924);
xnor U11788 (N_11788,N_9474,N_7939);
or U11789 (N_11789,N_9656,N_8642);
nand U11790 (N_11790,N_9546,N_8332);
nor U11791 (N_11791,N_9512,N_8373);
nand U11792 (N_11792,N_9680,N_8186);
or U11793 (N_11793,N_8527,N_7851);
xor U11794 (N_11794,N_9843,N_9784);
xor U11795 (N_11795,N_7670,N_8266);
nor U11796 (N_11796,N_7890,N_8625);
xnor U11797 (N_11797,N_8491,N_9862);
xnor U11798 (N_11798,N_7595,N_8999);
or U11799 (N_11799,N_9983,N_7774);
or U11800 (N_11800,N_9366,N_9835);
xnor U11801 (N_11801,N_8051,N_7884);
xor U11802 (N_11802,N_8462,N_8603);
nand U11803 (N_11803,N_9152,N_9504);
xor U11804 (N_11804,N_8698,N_8885);
nand U11805 (N_11805,N_7684,N_8354);
or U11806 (N_11806,N_8128,N_9048);
or U11807 (N_11807,N_9191,N_9879);
nor U11808 (N_11808,N_7640,N_8371);
nor U11809 (N_11809,N_9567,N_9184);
or U11810 (N_11810,N_8008,N_8382);
xnor U11811 (N_11811,N_9224,N_7789);
or U11812 (N_11812,N_9423,N_9880);
nand U11813 (N_11813,N_7579,N_8935);
xor U11814 (N_11814,N_8198,N_9567);
nor U11815 (N_11815,N_9061,N_8447);
nand U11816 (N_11816,N_9602,N_8673);
nand U11817 (N_11817,N_9344,N_9053);
nand U11818 (N_11818,N_8608,N_8670);
nand U11819 (N_11819,N_8386,N_8219);
xor U11820 (N_11820,N_8095,N_9987);
or U11821 (N_11821,N_7634,N_9141);
xnor U11822 (N_11822,N_8019,N_9293);
or U11823 (N_11823,N_8227,N_9078);
and U11824 (N_11824,N_7964,N_9347);
nor U11825 (N_11825,N_7575,N_8337);
or U11826 (N_11826,N_8000,N_9843);
xor U11827 (N_11827,N_8618,N_8311);
and U11828 (N_11828,N_8461,N_9272);
or U11829 (N_11829,N_9828,N_9226);
nor U11830 (N_11830,N_9737,N_7519);
or U11831 (N_11831,N_9727,N_8947);
xor U11832 (N_11832,N_8800,N_8504);
nand U11833 (N_11833,N_7504,N_9576);
and U11834 (N_11834,N_7955,N_8969);
and U11835 (N_11835,N_7923,N_8713);
or U11836 (N_11836,N_9636,N_8819);
xor U11837 (N_11837,N_9312,N_9019);
xnor U11838 (N_11838,N_7566,N_8112);
nor U11839 (N_11839,N_9648,N_8834);
or U11840 (N_11840,N_9417,N_9810);
nor U11841 (N_11841,N_7887,N_9227);
or U11842 (N_11842,N_9504,N_8257);
and U11843 (N_11843,N_8031,N_8641);
xor U11844 (N_11844,N_9942,N_8038);
nand U11845 (N_11845,N_8318,N_8731);
and U11846 (N_11846,N_8088,N_9071);
nor U11847 (N_11847,N_9209,N_9267);
or U11848 (N_11848,N_8892,N_8970);
or U11849 (N_11849,N_8845,N_9405);
xor U11850 (N_11850,N_7537,N_7514);
or U11851 (N_11851,N_9112,N_9781);
or U11852 (N_11852,N_7681,N_7937);
or U11853 (N_11853,N_9290,N_9104);
nor U11854 (N_11854,N_7503,N_7941);
nor U11855 (N_11855,N_7645,N_7662);
nor U11856 (N_11856,N_9042,N_8254);
or U11857 (N_11857,N_9846,N_8745);
nor U11858 (N_11858,N_7955,N_9109);
xnor U11859 (N_11859,N_7846,N_9073);
or U11860 (N_11860,N_9461,N_8852);
or U11861 (N_11861,N_8676,N_7849);
or U11862 (N_11862,N_9145,N_8797);
or U11863 (N_11863,N_9590,N_9588);
xor U11864 (N_11864,N_8563,N_8464);
nand U11865 (N_11865,N_8258,N_8698);
or U11866 (N_11866,N_9034,N_7617);
and U11867 (N_11867,N_7621,N_8026);
or U11868 (N_11868,N_7751,N_9044);
nand U11869 (N_11869,N_7629,N_9199);
or U11870 (N_11870,N_8080,N_9576);
nand U11871 (N_11871,N_8798,N_8649);
nor U11872 (N_11872,N_9983,N_8049);
nor U11873 (N_11873,N_7980,N_9636);
and U11874 (N_11874,N_7980,N_9082);
xor U11875 (N_11875,N_8929,N_7524);
xor U11876 (N_11876,N_8272,N_9093);
nand U11877 (N_11877,N_9492,N_9191);
nand U11878 (N_11878,N_9558,N_8856);
and U11879 (N_11879,N_8013,N_7824);
nand U11880 (N_11880,N_8882,N_8423);
nor U11881 (N_11881,N_7906,N_8474);
xor U11882 (N_11882,N_8027,N_8992);
xnor U11883 (N_11883,N_7553,N_8522);
xor U11884 (N_11884,N_7719,N_9506);
nand U11885 (N_11885,N_7508,N_8961);
xor U11886 (N_11886,N_9240,N_7879);
and U11887 (N_11887,N_8095,N_9935);
or U11888 (N_11888,N_8731,N_9546);
or U11889 (N_11889,N_9458,N_9389);
and U11890 (N_11890,N_8787,N_7686);
nand U11891 (N_11891,N_8209,N_9513);
nand U11892 (N_11892,N_9939,N_9203);
or U11893 (N_11893,N_9358,N_9448);
and U11894 (N_11894,N_9108,N_9691);
xor U11895 (N_11895,N_9328,N_9683);
xor U11896 (N_11896,N_9529,N_9244);
nor U11897 (N_11897,N_7894,N_8123);
xor U11898 (N_11898,N_9837,N_7538);
or U11899 (N_11899,N_8737,N_9616);
nand U11900 (N_11900,N_9123,N_9993);
nor U11901 (N_11901,N_9727,N_9487);
or U11902 (N_11902,N_7864,N_9988);
or U11903 (N_11903,N_9926,N_9095);
xor U11904 (N_11904,N_9109,N_9106);
and U11905 (N_11905,N_9127,N_9383);
or U11906 (N_11906,N_8936,N_8760);
xnor U11907 (N_11907,N_8563,N_8133);
nor U11908 (N_11908,N_9404,N_8537);
and U11909 (N_11909,N_7895,N_8774);
nor U11910 (N_11910,N_7838,N_8121);
or U11911 (N_11911,N_9357,N_9781);
xnor U11912 (N_11912,N_9121,N_8989);
or U11913 (N_11913,N_9905,N_9640);
or U11914 (N_11914,N_9802,N_8730);
nand U11915 (N_11915,N_9720,N_9090);
and U11916 (N_11916,N_8259,N_7832);
nor U11917 (N_11917,N_9954,N_8062);
and U11918 (N_11918,N_8488,N_8717);
xnor U11919 (N_11919,N_7801,N_8297);
nor U11920 (N_11920,N_9613,N_8838);
xor U11921 (N_11921,N_8957,N_9425);
or U11922 (N_11922,N_9801,N_9436);
and U11923 (N_11923,N_9740,N_7783);
nor U11924 (N_11924,N_9875,N_9697);
nor U11925 (N_11925,N_9277,N_7690);
nand U11926 (N_11926,N_8199,N_8135);
xnor U11927 (N_11927,N_8414,N_9945);
xnor U11928 (N_11928,N_7943,N_7754);
nor U11929 (N_11929,N_8073,N_8761);
xnor U11930 (N_11930,N_9679,N_8977);
xnor U11931 (N_11931,N_7997,N_8040);
nor U11932 (N_11932,N_8752,N_9515);
nand U11933 (N_11933,N_8694,N_9063);
and U11934 (N_11934,N_8790,N_8216);
or U11935 (N_11935,N_7751,N_8522);
nor U11936 (N_11936,N_8715,N_9814);
nand U11937 (N_11937,N_9863,N_8554);
nor U11938 (N_11938,N_8275,N_8894);
xor U11939 (N_11939,N_8198,N_8174);
or U11940 (N_11940,N_8410,N_8483);
and U11941 (N_11941,N_7541,N_7895);
or U11942 (N_11942,N_8189,N_8199);
or U11943 (N_11943,N_7568,N_7990);
nand U11944 (N_11944,N_8800,N_8191);
xor U11945 (N_11945,N_8593,N_8319);
xnor U11946 (N_11946,N_9927,N_8816);
and U11947 (N_11947,N_8541,N_9758);
and U11948 (N_11948,N_9087,N_9653);
nand U11949 (N_11949,N_9482,N_9035);
xor U11950 (N_11950,N_7870,N_8773);
nand U11951 (N_11951,N_8632,N_9826);
xnor U11952 (N_11952,N_9588,N_8230);
or U11953 (N_11953,N_7823,N_9084);
nand U11954 (N_11954,N_7823,N_9434);
and U11955 (N_11955,N_9313,N_9404);
or U11956 (N_11956,N_9618,N_9832);
nor U11957 (N_11957,N_9894,N_9248);
or U11958 (N_11958,N_8073,N_9254);
or U11959 (N_11959,N_7657,N_7790);
or U11960 (N_11960,N_9596,N_8500);
nand U11961 (N_11961,N_9158,N_7913);
or U11962 (N_11962,N_9734,N_7787);
xor U11963 (N_11963,N_8606,N_8148);
and U11964 (N_11964,N_7700,N_7995);
and U11965 (N_11965,N_8928,N_8083);
and U11966 (N_11966,N_8833,N_9947);
and U11967 (N_11967,N_7964,N_7927);
nand U11968 (N_11968,N_9101,N_8605);
nand U11969 (N_11969,N_8642,N_9940);
or U11970 (N_11970,N_8676,N_7631);
nand U11971 (N_11971,N_8472,N_8063);
xor U11972 (N_11972,N_8646,N_8531);
and U11973 (N_11973,N_8745,N_7865);
xnor U11974 (N_11974,N_9923,N_8743);
nand U11975 (N_11975,N_8152,N_9185);
nor U11976 (N_11976,N_8774,N_7838);
or U11977 (N_11977,N_9091,N_8120);
or U11978 (N_11978,N_9433,N_7670);
xor U11979 (N_11979,N_7754,N_8199);
xor U11980 (N_11980,N_8946,N_9652);
nand U11981 (N_11981,N_9315,N_7841);
xnor U11982 (N_11982,N_7886,N_8605);
xor U11983 (N_11983,N_8317,N_8117);
or U11984 (N_11984,N_7872,N_7987);
nand U11985 (N_11985,N_7845,N_9363);
nor U11986 (N_11986,N_8361,N_8419);
xor U11987 (N_11987,N_9304,N_9591);
nand U11988 (N_11988,N_8302,N_7880);
nand U11989 (N_11989,N_7687,N_8265);
nand U11990 (N_11990,N_9050,N_9790);
nor U11991 (N_11991,N_9625,N_7719);
xnor U11992 (N_11992,N_9002,N_8739);
and U11993 (N_11993,N_8288,N_7925);
and U11994 (N_11994,N_8889,N_8470);
or U11995 (N_11995,N_8213,N_9795);
nor U11996 (N_11996,N_7575,N_7686);
nor U11997 (N_11997,N_8272,N_9739);
nor U11998 (N_11998,N_8793,N_9514);
xor U11999 (N_11999,N_9500,N_8010);
nor U12000 (N_12000,N_7857,N_7988);
nor U12001 (N_12001,N_8561,N_9658);
nand U12002 (N_12002,N_9064,N_8403);
xor U12003 (N_12003,N_7845,N_8423);
xor U12004 (N_12004,N_9707,N_8400);
nand U12005 (N_12005,N_9813,N_9450);
and U12006 (N_12006,N_9157,N_7942);
nand U12007 (N_12007,N_9005,N_7568);
nor U12008 (N_12008,N_9381,N_7662);
xnor U12009 (N_12009,N_9397,N_7500);
and U12010 (N_12010,N_8684,N_7808);
or U12011 (N_12011,N_9893,N_8850);
or U12012 (N_12012,N_9766,N_9278);
and U12013 (N_12013,N_9335,N_9431);
nand U12014 (N_12014,N_9645,N_8791);
nor U12015 (N_12015,N_9578,N_9901);
or U12016 (N_12016,N_9706,N_9847);
nor U12017 (N_12017,N_7961,N_7880);
nor U12018 (N_12018,N_9282,N_9220);
nand U12019 (N_12019,N_9467,N_7714);
xnor U12020 (N_12020,N_7522,N_7871);
and U12021 (N_12021,N_8365,N_8897);
and U12022 (N_12022,N_8518,N_9599);
or U12023 (N_12023,N_9981,N_8412);
nor U12024 (N_12024,N_9207,N_7599);
nand U12025 (N_12025,N_7575,N_9443);
or U12026 (N_12026,N_7545,N_9549);
nand U12027 (N_12027,N_9736,N_8983);
nor U12028 (N_12028,N_9354,N_8294);
nand U12029 (N_12029,N_7730,N_7539);
or U12030 (N_12030,N_7654,N_7568);
and U12031 (N_12031,N_8005,N_7733);
and U12032 (N_12032,N_9927,N_7750);
or U12033 (N_12033,N_9474,N_8492);
nand U12034 (N_12034,N_8923,N_8795);
or U12035 (N_12035,N_8983,N_9106);
nor U12036 (N_12036,N_8057,N_8172);
xor U12037 (N_12037,N_8964,N_8306);
xnor U12038 (N_12038,N_9483,N_7966);
xnor U12039 (N_12039,N_8379,N_9102);
or U12040 (N_12040,N_7926,N_9747);
xnor U12041 (N_12041,N_7799,N_7649);
xnor U12042 (N_12042,N_9237,N_7681);
nand U12043 (N_12043,N_8841,N_8432);
or U12044 (N_12044,N_8347,N_9671);
nor U12045 (N_12045,N_9858,N_9077);
or U12046 (N_12046,N_9605,N_9113);
and U12047 (N_12047,N_8223,N_8342);
nor U12048 (N_12048,N_8920,N_8706);
nand U12049 (N_12049,N_7867,N_8055);
and U12050 (N_12050,N_9134,N_7681);
or U12051 (N_12051,N_8538,N_9970);
and U12052 (N_12052,N_8714,N_7991);
nand U12053 (N_12053,N_8720,N_7965);
and U12054 (N_12054,N_9123,N_9120);
xnor U12055 (N_12055,N_8919,N_8884);
nand U12056 (N_12056,N_7838,N_9572);
xor U12057 (N_12057,N_8682,N_9776);
and U12058 (N_12058,N_7653,N_8480);
and U12059 (N_12059,N_8548,N_8982);
nor U12060 (N_12060,N_8282,N_9364);
and U12061 (N_12061,N_9465,N_8410);
nor U12062 (N_12062,N_7604,N_9884);
xnor U12063 (N_12063,N_7691,N_8503);
or U12064 (N_12064,N_8307,N_9756);
xnor U12065 (N_12065,N_8881,N_8180);
or U12066 (N_12066,N_9691,N_7914);
nand U12067 (N_12067,N_7564,N_9977);
nor U12068 (N_12068,N_9417,N_7851);
xor U12069 (N_12069,N_8955,N_8253);
nor U12070 (N_12070,N_9878,N_8888);
xnor U12071 (N_12071,N_9138,N_9732);
or U12072 (N_12072,N_7889,N_8128);
and U12073 (N_12073,N_8348,N_7715);
xor U12074 (N_12074,N_8258,N_9512);
and U12075 (N_12075,N_9771,N_9226);
xnor U12076 (N_12076,N_7620,N_9255);
nand U12077 (N_12077,N_9645,N_8352);
nand U12078 (N_12078,N_8189,N_7985);
and U12079 (N_12079,N_8922,N_9467);
and U12080 (N_12080,N_9199,N_8380);
nand U12081 (N_12081,N_8027,N_7847);
or U12082 (N_12082,N_9204,N_8136);
nand U12083 (N_12083,N_9266,N_8009);
and U12084 (N_12084,N_9746,N_8713);
or U12085 (N_12085,N_9796,N_8075);
xor U12086 (N_12086,N_9251,N_9036);
and U12087 (N_12087,N_8867,N_8273);
nor U12088 (N_12088,N_9923,N_8856);
or U12089 (N_12089,N_8667,N_8030);
and U12090 (N_12090,N_9050,N_8319);
and U12091 (N_12091,N_9510,N_9221);
and U12092 (N_12092,N_8154,N_7673);
xnor U12093 (N_12093,N_9267,N_8937);
nor U12094 (N_12094,N_9247,N_8757);
or U12095 (N_12095,N_8160,N_8522);
or U12096 (N_12096,N_9084,N_9735);
nand U12097 (N_12097,N_7842,N_8120);
nand U12098 (N_12098,N_8819,N_9178);
or U12099 (N_12099,N_9533,N_7929);
nand U12100 (N_12100,N_8043,N_8089);
nor U12101 (N_12101,N_9398,N_9980);
xnor U12102 (N_12102,N_7692,N_8838);
nand U12103 (N_12103,N_9786,N_9447);
and U12104 (N_12104,N_7995,N_9511);
nand U12105 (N_12105,N_9995,N_8688);
or U12106 (N_12106,N_7551,N_9119);
and U12107 (N_12107,N_9665,N_9246);
nor U12108 (N_12108,N_9613,N_8525);
and U12109 (N_12109,N_9250,N_8762);
xnor U12110 (N_12110,N_8031,N_9224);
nor U12111 (N_12111,N_9562,N_8245);
and U12112 (N_12112,N_9013,N_7709);
xor U12113 (N_12113,N_8821,N_8759);
xnor U12114 (N_12114,N_8939,N_9110);
xnor U12115 (N_12115,N_9066,N_8241);
nor U12116 (N_12116,N_7861,N_8178);
nand U12117 (N_12117,N_8420,N_9457);
xor U12118 (N_12118,N_9246,N_8575);
and U12119 (N_12119,N_7698,N_8845);
nor U12120 (N_12120,N_9653,N_7542);
and U12121 (N_12121,N_8846,N_8958);
nand U12122 (N_12122,N_8755,N_9343);
xor U12123 (N_12123,N_8752,N_9339);
xnor U12124 (N_12124,N_8814,N_8994);
nor U12125 (N_12125,N_7663,N_9462);
xnor U12126 (N_12126,N_7578,N_9452);
or U12127 (N_12127,N_9361,N_8729);
nand U12128 (N_12128,N_8315,N_9091);
nor U12129 (N_12129,N_9578,N_9436);
nand U12130 (N_12130,N_8084,N_8152);
xor U12131 (N_12131,N_8423,N_8044);
nor U12132 (N_12132,N_7658,N_8353);
xnor U12133 (N_12133,N_8956,N_7786);
nand U12134 (N_12134,N_9044,N_7721);
xnor U12135 (N_12135,N_7833,N_8643);
nand U12136 (N_12136,N_7637,N_9266);
nand U12137 (N_12137,N_7937,N_9963);
nand U12138 (N_12138,N_7918,N_8414);
and U12139 (N_12139,N_7828,N_8708);
nor U12140 (N_12140,N_8807,N_9794);
xnor U12141 (N_12141,N_8044,N_8860);
xnor U12142 (N_12142,N_8944,N_8041);
or U12143 (N_12143,N_8592,N_9230);
nand U12144 (N_12144,N_7584,N_8544);
nor U12145 (N_12145,N_7604,N_8452);
and U12146 (N_12146,N_7952,N_8404);
or U12147 (N_12147,N_7885,N_8171);
nor U12148 (N_12148,N_7696,N_8815);
xor U12149 (N_12149,N_8751,N_9348);
xnor U12150 (N_12150,N_9965,N_9136);
and U12151 (N_12151,N_8087,N_7822);
and U12152 (N_12152,N_8275,N_8599);
nand U12153 (N_12153,N_9835,N_7755);
or U12154 (N_12154,N_7860,N_8723);
or U12155 (N_12155,N_7724,N_9373);
and U12156 (N_12156,N_8476,N_9491);
nand U12157 (N_12157,N_8945,N_8002);
nor U12158 (N_12158,N_8377,N_9029);
or U12159 (N_12159,N_7603,N_7772);
nand U12160 (N_12160,N_9558,N_8050);
or U12161 (N_12161,N_9396,N_7614);
nand U12162 (N_12162,N_7510,N_8473);
nor U12163 (N_12163,N_9921,N_7827);
or U12164 (N_12164,N_8788,N_8889);
and U12165 (N_12165,N_7950,N_7711);
or U12166 (N_12166,N_9942,N_9941);
nand U12167 (N_12167,N_8457,N_9515);
nor U12168 (N_12168,N_7894,N_9857);
nand U12169 (N_12169,N_9436,N_9529);
xor U12170 (N_12170,N_8476,N_8016);
xor U12171 (N_12171,N_9509,N_8130);
xor U12172 (N_12172,N_9106,N_7887);
nor U12173 (N_12173,N_9887,N_8385);
or U12174 (N_12174,N_8754,N_9760);
and U12175 (N_12175,N_9760,N_8726);
and U12176 (N_12176,N_8120,N_7627);
xor U12177 (N_12177,N_7744,N_9561);
and U12178 (N_12178,N_7562,N_7552);
xnor U12179 (N_12179,N_9376,N_9901);
nand U12180 (N_12180,N_8648,N_7541);
or U12181 (N_12181,N_8971,N_9973);
xor U12182 (N_12182,N_8642,N_8542);
nand U12183 (N_12183,N_8549,N_9107);
nor U12184 (N_12184,N_9907,N_8173);
and U12185 (N_12185,N_9997,N_9543);
xnor U12186 (N_12186,N_7803,N_8785);
and U12187 (N_12187,N_9801,N_9081);
or U12188 (N_12188,N_8698,N_7965);
xnor U12189 (N_12189,N_9051,N_8357);
or U12190 (N_12190,N_8776,N_8642);
and U12191 (N_12191,N_8225,N_9010);
nand U12192 (N_12192,N_9692,N_7914);
or U12193 (N_12193,N_8719,N_9323);
or U12194 (N_12194,N_8471,N_8940);
or U12195 (N_12195,N_8358,N_8709);
or U12196 (N_12196,N_9795,N_9807);
xor U12197 (N_12197,N_7565,N_9396);
or U12198 (N_12198,N_8203,N_9087);
nand U12199 (N_12199,N_9048,N_9747);
nor U12200 (N_12200,N_8191,N_7619);
nor U12201 (N_12201,N_9131,N_7996);
or U12202 (N_12202,N_9659,N_9313);
and U12203 (N_12203,N_8333,N_9925);
nor U12204 (N_12204,N_7990,N_9579);
xnor U12205 (N_12205,N_8848,N_9069);
nor U12206 (N_12206,N_8047,N_8068);
xor U12207 (N_12207,N_9984,N_8610);
xor U12208 (N_12208,N_8627,N_9767);
or U12209 (N_12209,N_8945,N_8949);
or U12210 (N_12210,N_8385,N_7846);
and U12211 (N_12211,N_9994,N_8702);
or U12212 (N_12212,N_9950,N_8145);
nor U12213 (N_12213,N_8981,N_8636);
nor U12214 (N_12214,N_8235,N_9399);
and U12215 (N_12215,N_9024,N_8707);
or U12216 (N_12216,N_9690,N_8421);
nand U12217 (N_12217,N_8738,N_7764);
xnor U12218 (N_12218,N_9369,N_8361);
nor U12219 (N_12219,N_9671,N_9983);
nor U12220 (N_12220,N_8224,N_8490);
nor U12221 (N_12221,N_9265,N_8989);
nor U12222 (N_12222,N_8861,N_7930);
nor U12223 (N_12223,N_8808,N_9455);
or U12224 (N_12224,N_9579,N_8240);
nor U12225 (N_12225,N_8030,N_7865);
xnor U12226 (N_12226,N_7557,N_7522);
and U12227 (N_12227,N_9138,N_7838);
and U12228 (N_12228,N_9418,N_9663);
and U12229 (N_12229,N_7937,N_8760);
nor U12230 (N_12230,N_8533,N_8816);
or U12231 (N_12231,N_8530,N_8397);
and U12232 (N_12232,N_9701,N_9589);
nand U12233 (N_12233,N_7712,N_7525);
nor U12234 (N_12234,N_9746,N_8711);
xor U12235 (N_12235,N_7883,N_9810);
or U12236 (N_12236,N_9557,N_8304);
xor U12237 (N_12237,N_9652,N_9862);
nor U12238 (N_12238,N_7827,N_9996);
nor U12239 (N_12239,N_7725,N_9611);
nor U12240 (N_12240,N_8202,N_9598);
or U12241 (N_12241,N_7568,N_8471);
nor U12242 (N_12242,N_7500,N_9462);
and U12243 (N_12243,N_8086,N_8211);
xor U12244 (N_12244,N_7650,N_7666);
xnor U12245 (N_12245,N_7548,N_7882);
nor U12246 (N_12246,N_9626,N_9422);
and U12247 (N_12247,N_8224,N_9258);
and U12248 (N_12248,N_8809,N_7950);
and U12249 (N_12249,N_8774,N_9632);
xor U12250 (N_12250,N_9589,N_9075);
or U12251 (N_12251,N_8480,N_9096);
and U12252 (N_12252,N_8593,N_9997);
nand U12253 (N_12253,N_9719,N_9514);
or U12254 (N_12254,N_8922,N_9478);
or U12255 (N_12255,N_8581,N_9534);
and U12256 (N_12256,N_7572,N_8768);
xor U12257 (N_12257,N_8491,N_9215);
xnor U12258 (N_12258,N_8234,N_9005);
xor U12259 (N_12259,N_8567,N_8979);
nand U12260 (N_12260,N_8235,N_8385);
nand U12261 (N_12261,N_9638,N_8028);
or U12262 (N_12262,N_9447,N_8281);
xor U12263 (N_12263,N_8260,N_9737);
xnor U12264 (N_12264,N_9178,N_9913);
and U12265 (N_12265,N_9897,N_8522);
nand U12266 (N_12266,N_8175,N_8163);
and U12267 (N_12267,N_7707,N_7889);
nor U12268 (N_12268,N_8871,N_8213);
or U12269 (N_12269,N_8448,N_8104);
nor U12270 (N_12270,N_8508,N_9321);
nand U12271 (N_12271,N_7744,N_9931);
xnor U12272 (N_12272,N_8459,N_9667);
or U12273 (N_12273,N_7804,N_8513);
and U12274 (N_12274,N_7885,N_9792);
nand U12275 (N_12275,N_9350,N_8118);
and U12276 (N_12276,N_9005,N_9957);
nor U12277 (N_12277,N_9966,N_7944);
or U12278 (N_12278,N_9816,N_9147);
nand U12279 (N_12279,N_8991,N_7578);
xnor U12280 (N_12280,N_8878,N_8880);
nor U12281 (N_12281,N_7688,N_9273);
or U12282 (N_12282,N_7564,N_8317);
xor U12283 (N_12283,N_8444,N_9468);
nor U12284 (N_12284,N_9369,N_9923);
or U12285 (N_12285,N_9977,N_9211);
xor U12286 (N_12286,N_9802,N_8016);
nand U12287 (N_12287,N_9931,N_9882);
nor U12288 (N_12288,N_7557,N_7809);
and U12289 (N_12289,N_8132,N_8861);
or U12290 (N_12290,N_9166,N_9405);
nand U12291 (N_12291,N_7865,N_8036);
nand U12292 (N_12292,N_8466,N_9630);
nand U12293 (N_12293,N_8695,N_9258);
xnor U12294 (N_12294,N_9198,N_8490);
xor U12295 (N_12295,N_7922,N_9126);
or U12296 (N_12296,N_9099,N_7616);
xor U12297 (N_12297,N_9590,N_7502);
nand U12298 (N_12298,N_8205,N_8250);
nor U12299 (N_12299,N_7866,N_8915);
xnor U12300 (N_12300,N_9881,N_7946);
and U12301 (N_12301,N_9911,N_7596);
nand U12302 (N_12302,N_7731,N_8975);
or U12303 (N_12303,N_9672,N_9947);
xor U12304 (N_12304,N_8229,N_7982);
xor U12305 (N_12305,N_8073,N_7740);
and U12306 (N_12306,N_8890,N_8407);
or U12307 (N_12307,N_7783,N_8800);
nand U12308 (N_12308,N_8058,N_9054);
nand U12309 (N_12309,N_9671,N_9751);
and U12310 (N_12310,N_8013,N_8820);
nand U12311 (N_12311,N_7897,N_7714);
and U12312 (N_12312,N_7702,N_7506);
and U12313 (N_12313,N_7555,N_9395);
and U12314 (N_12314,N_9208,N_9844);
nor U12315 (N_12315,N_8871,N_8953);
or U12316 (N_12316,N_8214,N_7724);
nor U12317 (N_12317,N_9373,N_8906);
or U12318 (N_12318,N_8288,N_9583);
nand U12319 (N_12319,N_9490,N_7731);
nor U12320 (N_12320,N_7981,N_7956);
or U12321 (N_12321,N_9715,N_9578);
xnor U12322 (N_12322,N_9283,N_9924);
nand U12323 (N_12323,N_8468,N_9572);
and U12324 (N_12324,N_8339,N_9967);
and U12325 (N_12325,N_9937,N_8014);
and U12326 (N_12326,N_7575,N_9803);
or U12327 (N_12327,N_7982,N_8676);
nor U12328 (N_12328,N_8774,N_9856);
nand U12329 (N_12329,N_9885,N_7876);
and U12330 (N_12330,N_8969,N_8423);
and U12331 (N_12331,N_9080,N_8471);
and U12332 (N_12332,N_8010,N_8141);
and U12333 (N_12333,N_7523,N_9802);
xnor U12334 (N_12334,N_8454,N_9027);
xor U12335 (N_12335,N_7997,N_8596);
nor U12336 (N_12336,N_7873,N_7767);
nor U12337 (N_12337,N_9028,N_8698);
or U12338 (N_12338,N_9441,N_7883);
and U12339 (N_12339,N_9808,N_7933);
or U12340 (N_12340,N_8267,N_7642);
xnor U12341 (N_12341,N_9152,N_8739);
and U12342 (N_12342,N_9880,N_8222);
nand U12343 (N_12343,N_8452,N_8397);
nand U12344 (N_12344,N_9996,N_9226);
or U12345 (N_12345,N_9508,N_8452);
xor U12346 (N_12346,N_8099,N_8254);
nand U12347 (N_12347,N_8859,N_9789);
nand U12348 (N_12348,N_9343,N_9522);
and U12349 (N_12349,N_8689,N_8760);
and U12350 (N_12350,N_9585,N_9795);
nand U12351 (N_12351,N_8496,N_8456);
nand U12352 (N_12352,N_8812,N_7500);
or U12353 (N_12353,N_8216,N_8340);
nand U12354 (N_12354,N_8905,N_9718);
and U12355 (N_12355,N_8204,N_9725);
nor U12356 (N_12356,N_9239,N_9226);
xnor U12357 (N_12357,N_7501,N_8343);
nand U12358 (N_12358,N_9301,N_7620);
or U12359 (N_12359,N_8051,N_8181);
or U12360 (N_12360,N_8164,N_9181);
xnor U12361 (N_12361,N_7914,N_8767);
nor U12362 (N_12362,N_8845,N_8100);
and U12363 (N_12363,N_9101,N_8248);
or U12364 (N_12364,N_9877,N_7678);
or U12365 (N_12365,N_9201,N_9856);
nor U12366 (N_12366,N_9785,N_9140);
and U12367 (N_12367,N_9900,N_8747);
xnor U12368 (N_12368,N_9261,N_8356);
nor U12369 (N_12369,N_9498,N_9967);
nor U12370 (N_12370,N_9599,N_7649);
nor U12371 (N_12371,N_8927,N_8158);
xnor U12372 (N_12372,N_9671,N_7735);
and U12373 (N_12373,N_9601,N_8848);
nand U12374 (N_12374,N_9897,N_8369);
xnor U12375 (N_12375,N_9185,N_9504);
nor U12376 (N_12376,N_8142,N_8400);
nand U12377 (N_12377,N_9823,N_8010);
and U12378 (N_12378,N_8962,N_9972);
or U12379 (N_12379,N_9177,N_9053);
nand U12380 (N_12380,N_8479,N_7658);
or U12381 (N_12381,N_9424,N_8266);
nand U12382 (N_12382,N_8830,N_7863);
nand U12383 (N_12383,N_9647,N_7502);
nor U12384 (N_12384,N_9479,N_8459);
xor U12385 (N_12385,N_8023,N_9998);
nor U12386 (N_12386,N_9820,N_9284);
nor U12387 (N_12387,N_9802,N_9912);
or U12388 (N_12388,N_9299,N_9742);
or U12389 (N_12389,N_9317,N_9271);
nand U12390 (N_12390,N_9798,N_7877);
or U12391 (N_12391,N_7806,N_7914);
and U12392 (N_12392,N_8479,N_8533);
nor U12393 (N_12393,N_7540,N_9333);
or U12394 (N_12394,N_9132,N_8733);
xnor U12395 (N_12395,N_9973,N_7745);
nand U12396 (N_12396,N_8023,N_8880);
nor U12397 (N_12397,N_7534,N_8016);
nor U12398 (N_12398,N_9284,N_9117);
and U12399 (N_12399,N_7899,N_8739);
xor U12400 (N_12400,N_7561,N_7706);
or U12401 (N_12401,N_9727,N_9327);
xnor U12402 (N_12402,N_8043,N_7620);
nand U12403 (N_12403,N_7606,N_9223);
or U12404 (N_12404,N_8706,N_8366);
nor U12405 (N_12405,N_8588,N_7840);
and U12406 (N_12406,N_9734,N_7508);
and U12407 (N_12407,N_8250,N_7674);
nor U12408 (N_12408,N_9012,N_7835);
or U12409 (N_12409,N_7558,N_9551);
and U12410 (N_12410,N_7530,N_7744);
xor U12411 (N_12411,N_9314,N_9381);
or U12412 (N_12412,N_7720,N_8469);
and U12413 (N_12413,N_8827,N_9789);
and U12414 (N_12414,N_9631,N_9804);
and U12415 (N_12415,N_9897,N_9813);
nand U12416 (N_12416,N_9928,N_9539);
nor U12417 (N_12417,N_9723,N_8108);
and U12418 (N_12418,N_7620,N_9268);
xor U12419 (N_12419,N_9754,N_8652);
and U12420 (N_12420,N_7513,N_9659);
nor U12421 (N_12421,N_7540,N_8529);
xnor U12422 (N_12422,N_7939,N_8880);
xor U12423 (N_12423,N_7554,N_8265);
nor U12424 (N_12424,N_8853,N_9364);
or U12425 (N_12425,N_9699,N_7773);
and U12426 (N_12426,N_9400,N_9746);
and U12427 (N_12427,N_8400,N_9094);
nand U12428 (N_12428,N_9697,N_8326);
or U12429 (N_12429,N_7909,N_9532);
nand U12430 (N_12430,N_8722,N_7769);
nor U12431 (N_12431,N_9948,N_9486);
and U12432 (N_12432,N_9462,N_8072);
nand U12433 (N_12433,N_9347,N_8304);
and U12434 (N_12434,N_9731,N_8400);
nand U12435 (N_12435,N_7792,N_7817);
xnor U12436 (N_12436,N_7602,N_9026);
and U12437 (N_12437,N_9232,N_9985);
xnor U12438 (N_12438,N_9730,N_8237);
xor U12439 (N_12439,N_9859,N_8685);
nor U12440 (N_12440,N_9160,N_9214);
or U12441 (N_12441,N_9223,N_8870);
xor U12442 (N_12442,N_9645,N_9676);
xor U12443 (N_12443,N_8745,N_7771);
or U12444 (N_12444,N_7826,N_8000);
and U12445 (N_12445,N_7522,N_8027);
xnor U12446 (N_12446,N_8989,N_9738);
and U12447 (N_12447,N_8833,N_7814);
or U12448 (N_12448,N_8717,N_9769);
xor U12449 (N_12449,N_9352,N_9092);
or U12450 (N_12450,N_8217,N_9884);
and U12451 (N_12451,N_8629,N_9417);
xor U12452 (N_12452,N_7913,N_7524);
nor U12453 (N_12453,N_8985,N_9727);
xor U12454 (N_12454,N_8140,N_7776);
nand U12455 (N_12455,N_7659,N_8625);
nor U12456 (N_12456,N_8395,N_8819);
nand U12457 (N_12457,N_8184,N_9753);
and U12458 (N_12458,N_7941,N_8464);
or U12459 (N_12459,N_9052,N_9786);
or U12460 (N_12460,N_9587,N_8108);
nor U12461 (N_12461,N_8420,N_9493);
nor U12462 (N_12462,N_8806,N_8448);
and U12463 (N_12463,N_7530,N_7822);
nor U12464 (N_12464,N_9693,N_8304);
xor U12465 (N_12465,N_9332,N_9501);
xor U12466 (N_12466,N_9889,N_9339);
or U12467 (N_12467,N_7921,N_8163);
xor U12468 (N_12468,N_8719,N_7535);
and U12469 (N_12469,N_9017,N_7803);
nand U12470 (N_12470,N_8687,N_7829);
and U12471 (N_12471,N_8595,N_9313);
and U12472 (N_12472,N_8953,N_9686);
or U12473 (N_12473,N_7979,N_9595);
and U12474 (N_12474,N_7634,N_8627);
xor U12475 (N_12475,N_9551,N_9967);
and U12476 (N_12476,N_9915,N_7565);
and U12477 (N_12477,N_9076,N_8473);
xor U12478 (N_12478,N_8642,N_9980);
nand U12479 (N_12479,N_9775,N_8321);
nor U12480 (N_12480,N_8141,N_8114);
xnor U12481 (N_12481,N_9758,N_8743);
xor U12482 (N_12482,N_8044,N_9596);
xnor U12483 (N_12483,N_8999,N_8953);
and U12484 (N_12484,N_8134,N_8327);
or U12485 (N_12485,N_7611,N_9767);
xnor U12486 (N_12486,N_9442,N_9640);
or U12487 (N_12487,N_8674,N_8454);
nor U12488 (N_12488,N_7980,N_7873);
or U12489 (N_12489,N_8329,N_8155);
xnor U12490 (N_12490,N_8667,N_9164);
or U12491 (N_12491,N_8080,N_8428);
nor U12492 (N_12492,N_9086,N_8751);
and U12493 (N_12493,N_7589,N_9349);
and U12494 (N_12494,N_9716,N_7777);
nand U12495 (N_12495,N_9306,N_9767);
and U12496 (N_12496,N_8629,N_9014);
xor U12497 (N_12497,N_9388,N_8094);
xnor U12498 (N_12498,N_9464,N_9476);
xnor U12499 (N_12499,N_8758,N_8134);
and U12500 (N_12500,N_12445,N_10296);
xnor U12501 (N_12501,N_10496,N_10716);
and U12502 (N_12502,N_10528,N_11722);
xnor U12503 (N_12503,N_10430,N_12102);
xor U12504 (N_12504,N_11465,N_10491);
nor U12505 (N_12505,N_11682,N_10271);
nand U12506 (N_12506,N_10860,N_12339);
or U12507 (N_12507,N_11270,N_11955);
and U12508 (N_12508,N_11740,N_11483);
xnor U12509 (N_12509,N_11837,N_11318);
nand U12510 (N_12510,N_11113,N_10704);
xor U12511 (N_12511,N_12136,N_10957);
or U12512 (N_12512,N_10295,N_12128);
xor U12513 (N_12513,N_11017,N_10299);
or U12514 (N_12514,N_11616,N_11251);
xnor U12515 (N_12515,N_11338,N_11329);
nor U12516 (N_12516,N_11103,N_11264);
and U12517 (N_12517,N_12322,N_12359);
nand U12518 (N_12518,N_12082,N_10002);
nor U12519 (N_12519,N_11424,N_11189);
or U12520 (N_12520,N_10055,N_10941);
or U12521 (N_12521,N_12204,N_10897);
or U12522 (N_12522,N_10687,N_11810);
or U12523 (N_12523,N_12378,N_11684);
xor U12524 (N_12524,N_12274,N_11351);
nor U12525 (N_12525,N_10390,N_10706);
and U12526 (N_12526,N_10555,N_10153);
or U12527 (N_12527,N_10066,N_11057);
or U12528 (N_12528,N_11414,N_10549);
nor U12529 (N_12529,N_11686,N_11354);
nor U12530 (N_12530,N_10877,N_11493);
or U12531 (N_12531,N_10473,N_12277);
nor U12532 (N_12532,N_11238,N_11924);
or U12533 (N_12533,N_11211,N_12326);
nand U12534 (N_12534,N_11223,N_11922);
and U12535 (N_12535,N_10566,N_10617);
and U12536 (N_12536,N_10280,N_10330);
nor U12537 (N_12537,N_12447,N_10070);
and U12538 (N_12538,N_10481,N_11903);
xnor U12539 (N_12539,N_11818,N_11366);
nor U12540 (N_12540,N_11869,N_11075);
xnor U12541 (N_12541,N_12116,N_11752);
xor U12542 (N_12542,N_12077,N_10080);
xor U12543 (N_12543,N_10712,N_10602);
or U12544 (N_12544,N_11213,N_11850);
or U12545 (N_12545,N_11167,N_10967);
nand U12546 (N_12546,N_11543,N_12216);
and U12547 (N_12547,N_12185,N_10592);
or U12548 (N_12548,N_11349,N_12047);
xnor U12549 (N_12549,N_11060,N_11120);
xor U12550 (N_12550,N_10419,N_11938);
nor U12551 (N_12551,N_11742,N_12352);
and U12552 (N_12552,N_12444,N_10908);
nand U12553 (N_12553,N_12475,N_10341);
or U12554 (N_12554,N_12081,N_12381);
or U12555 (N_12555,N_10527,N_12390);
or U12556 (N_12556,N_10583,N_11962);
nand U12557 (N_12557,N_11772,N_10115);
xor U12558 (N_12558,N_12417,N_11546);
and U12559 (N_12559,N_10287,N_10685);
xnor U12560 (N_12560,N_11111,N_12182);
nand U12561 (N_12561,N_10762,N_12002);
xnor U12562 (N_12562,N_11395,N_11530);
or U12563 (N_12563,N_11952,N_10626);
xnor U12564 (N_12564,N_11193,N_11510);
or U12565 (N_12565,N_11316,N_10820);
xor U12566 (N_12566,N_10771,N_11601);
xor U12567 (N_12567,N_11176,N_10684);
nand U12568 (N_12568,N_11524,N_11014);
nor U12569 (N_12569,N_11857,N_11032);
nand U12570 (N_12570,N_12334,N_10506);
and U12571 (N_12571,N_12060,N_11846);
or U12572 (N_12572,N_11638,N_12398);
nand U12573 (N_12573,N_12492,N_12178);
nand U12574 (N_12574,N_12411,N_11596);
and U12575 (N_12575,N_10093,N_12227);
and U12576 (N_12576,N_11816,N_10038);
and U12577 (N_12577,N_11241,N_11203);
nand U12578 (N_12578,N_12320,N_12246);
nor U12579 (N_12579,N_11308,N_11919);
xor U12580 (N_12580,N_11028,N_12033);
nand U12581 (N_12581,N_11458,N_11355);
and U12582 (N_12582,N_11324,N_10054);
xnor U12583 (N_12583,N_11501,N_12155);
or U12584 (N_12584,N_11487,N_10503);
or U12585 (N_12585,N_11352,N_11575);
and U12586 (N_12586,N_11831,N_11166);
or U12587 (N_12587,N_10278,N_10459);
and U12588 (N_12588,N_10558,N_11262);
nor U12589 (N_12589,N_10821,N_10560);
or U12590 (N_12590,N_10996,N_11974);
and U12591 (N_12591,N_11401,N_10791);
and U12592 (N_12592,N_10914,N_10199);
or U12593 (N_12593,N_10709,N_12016);
nand U12594 (N_12594,N_11147,N_12305);
and U12595 (N_12595,N_10323,N_11765);
or U12596 (N_12596,N_11893,N_10561);
and U12597 (N_12597,N_11978,N_12476);
nor U12598 (N_12598,N_11536,N_10983);
nor U12599 (N_12599,N_11729,N_11709);
nor U12600 (N_12600,N_10450,N_12197);
xnor U12601 (N_12601,N_11902,N_10067);
nor U12602 (N_12602,N_12371,N_10504);
and U12603 (N_12603,N_10679,N_10207);
nand U12604 (N_12604,N_10849,N_11997);
nand U12605 (N_12605,N_12027,N_12165);
nor U12606 (N_12606,N_12349,N_11126);
nor U12607 (N_12607,N_11931,N_10608);
xnor U12608 (N_12608,N_10866,N_10939);
and U12609 (N_12609,N_11710,N_10913);
or U12610 (N_12610,N_10845,N_10012);
and U12611 (N_12611,N_11631,N_11130);
and U12612 (N_12612,N_10343,N_10209);
nor U12613 (N_12613,N_12147,N_11158);
or U12614 (N_12614,N_11134,N_10895);
nand U12615 (N_12615,N_11376,N_12196);
xnor U12616 (N_12616,N_11399,N_12198);
and U12617 (N_12617,N_10361,N_10783);
or U12618 (N_12618,N_12361,N_12369);
or U12619 (N_12619,N_11894,N_11673);
nor U12620 (N_12620,N_12042,N_11610);
or U12621 (N_12621,N_12287,N_11252);
nand U12622 (N_12622,N_11625,N_10765);
nand U12623 (N_12623,N_10719,N_10382);
xnor U12624 (N_12624,N_10170,N_12223);
nor U12625 (N_12625,N_11975,N_11101);
and U12626 (N_12626,N_11909,N_10805);
and U12627 (N_12627,N_10814,N_11074);
nand U12628 (N_12628,N_12459,N_10963);
and U12629 (N_12629,N_10754,N_11467);
or U12630 (N_12630,N_11704,N_11331);
or U12631 (N_12631,N_12207,N_12259);
nor U12632 (N_12632,N_11152,N_10898);
nor U12633 (N_12633,N_12377,N_10412);
nor U12634 (N_12634,N_12154,N_10634);
nand U12635 (N_12635,N_11927,N_10136);
xnor U12636 (N_12636,N_12192,N_10091);
and U12637 (N_12637,N_10168,N_12142);
nand U12638 (N_12638,N_11701,N_12400);
and U12639 (N_12639,N_10391,N_11904);
and U12640 (N_12640,N_12222,N_10517);
xor U12641 (N_12641,N_10681,N_10014);
nand U12642 (N_12642,N_10127,N_11895);
and U12643 (N_12643,N_10578,N_10392);
nor U12644 (N_12644,N_11044,N_10605);
nor U12645 (N_12645,N_11164,N_12413);
or U12646 (N_12646,N_10722,N_11015);
and U12647 (N_12647,N_12432,N_11887);
or U12648 (N_12648,N_11808,N_11215);
nand U12649 (N_12649,N_11677,N_10970);
nor U12650 (N_12650,N_10004,N_12109);
or U12651 (N_12651,N_10497,N_11806);
xor U12652 (N_12652,N_12236,N_10520);
nand U12653 (N_12653,N_10863,N_11388);
or U12654 (N_12654,N_11052,N_11804);
nor U12655 (N_12655,N_12397,N_11650);
and U12656 (N_12656,N_10904,N_11774);
nor U12657 (N_12657,N_11732,N_11245);
xnor U12658 (N_12658,N_10058,N_11934);
xnor U12659 (N_12659,N_12433,N_10976);
nor U12660 (N_12660,N_10281,N_10173);
or U12661 (N_12661,N_10165,N_11754);
and U12662 (N_12662,N_12293,N_11538);
xor U12663 (N_12663,N_10793,N_11300);
and U12664 (N_12664,N_11606,N_11844);
nor U12665 (N_12665,N_10965,N_12212);
nand U12666 (N_12666,N_12086,N_11992);
nor U12667 (N_12667,N_11059,N_11009);
nor U12668 (N_12668,N_11498,N_12306);
nand U12669 (N_12669,N_12017,N_10064);
xor U12670 (N_12670,N_10697,N_12477);
xnor U12671 (N_12671,N_10163,N_12255);
xor U12672 (N_12672,N_10580,N_11186);
and U12673 (N_12673,N_12229,N_12497);
and U12674 (N_12674,N_10698,N_10922);
or U12675 (N_12675,N_10358,N_12450);
or U12676 (N_12676,N_10554,N_11875);
nand U12677 (N_12677,N_10891,N_11696);
xor U12678 (N_12678,N_10338,N_10594);
xor U12679 (N_12679,N_10662,N_10407);
or U12680 (N_12680,N_10905,N_10188);
nor U12681 (N_12681,N_12065,N_11348);
nand U12682 (N_12682,N_10625,N_10478);
nor U12683 (N_12683,N_10406,N_10943);
or U12684 (N_12684,N_12394,N_11259);
and U12685 (N_12685,N_12210,N_11076);
nand U12686 (N_12686,N_12262,N_12493);
xor U12687 (N_12687,N_10595,N_11666);
or U12688 (N_12688,N_12375,N_10256);
or U12689 (N_12689,N_10534,N_11121);
nand U12690 (N_12690,N_11471,N_10919);
or U12691 (N_12691,N_11634,N_10696);
nand U12692 (N_12692,N_11013,N_10337);
and U12693 (N_12693,N_12468,N_12125);
nand U12694 (N_12694,N_11146,N_11100);
nand U12695 (N_12695,N_11160,N_10183);
or U12696 (N_12696,N_10413,N_10312);
xnor U12697 (N_12697,N_11566,N_12064);
and U12698 (N_12698,N_11012,N_12130);
nor U12699 (N_12699,N_12135,N_12396);
or U12700 (N_12700,N_10158,N_11593);
or U12701 (N_12701,N_11550,N_10807);
and U12702 (N_12702,N_10861,N_12494);
nand U12703 (N_12703,N_10859,N_11107);
or U12704 (N_12704,N_10551,N_12333);
and U12705 (N_12705,N_10353,N_11700);
and U12706 (N_12706,N_11412,N_11557);
or U12707 (N_12707,N_11532,N_11626);
xnor U12708 (N_12708,N_10786,N_10345);
nor U12709 (N_12709,N_10034,N_10282);
or U12710 (N_12710,N_10700,N_10540);
xnor U12711 (N_12711,N_11861,N_11826);
nand U12712 (N_12712,N_11436,N_11144);
xnor U12713 (N_12713,N_12256,N_12111);
xor U12714 (N_12714,N_10801,N_11265);
and U12715 (N_12715,N_11481,N_11492);
nand U12716 (N_12716,N_12007,N_12195);
or U12717 (N_12717,N_11415,N_12465);
nand U12718 (N_12718,N_11637,N_11081);
nand U12719 (N_12719,N_10253,N_10446);
nor U12720 (N_12720,N_10451,N_11527);
and U12721 (N_12721,N_10693,N_12053);
xnor U12722 (N_12722,N_11583,N_11541);
xor U12723 (N_12723,N_12340,N_10324);
nand U12724 (N_12724,N_11764,N_12235);
nor U12725 (N_12725,N_12092,N_10006);
nor U12726 (N_12726,N_12491,N_11452);
nor U12727 (N_12727,N_11983,N_10699);
xor U12728 (N_12728,N_10105,N_10770);
or U12729 (N_12729,N_11592,N_10111);
nand U12730 (N_12730,N_11611,N_10665);
xnor U12731 (N_12731,N_11613,N_11460);
nor U12732 (N_12732,N_11562,N_11357);
and U12733 (N_12733,N_10039,N_10344);
nand U12734 (N_12734,N_11712,N_10180);
nand U12735 (N_12735,N_11309,N_12088);
xor U12736 (N_12736,N_11840,N_11942);
or U12737 (N_12737,N_10537,N_10829);
and U12738 (N_12738,N_12286,N_11208);
nand U12739 (N_12739,N_11283,N_10499);
and U12740 (N_12740,N_11254,N_10893);
xnor U12741 (N_12741,N_10531,N_12271);
or U12742 (N_12742,N_11038,N_10792);
nor U12743 (N_12743,N_10736,N_11271);
nand U12744 (N_12744,N_11248,N_11603);
nor U12745 (N_12745,N_11085,N_12302);
nand U12746 (N_12746,N_12159,N_11953);
and U12747 (N_12747,N_11797,N_10972);
or U12748 (N_12748,N_11434,N_10273);
nor U12749 (N_12749,N_10912,N_11124);
or U12750 (N_12750,N_10374,N_10755);
or U12751 (N_12751,N_10611,N_10760);
nor U12752 (N_12752,N_10899,N_10156);
and U12753 (N_12753,N_10892,N_10266);
or U12754 (N_12754,N_11499,N_12441);
xor U12755 (N_12755,N_10176,N_11125);
nand U12756 (N_12756,N_11668,N_11822);
nor U12757 (N_12757,N_12437,N_10936);
nor U12758 (N_12758,N_11128,N_12261);
nand U12759 (N_12759,N_11192,N_10572);
and U12760 (N_12760,N_11373,N_12211);
nand U12761 (N_12761,N_11217,N_11617);
xnor U12762 (N_12762,N_10140,N_10509);
nand U12763 (N_12763,N_11182,N_10663);
nor U12764 (N_12764,N_10079,N_11266);
xor U12765 (N_12765,N_10620,N_10095);
and U12766 (N_12766,N_12041,N_11896);
nand U12767 (N_12767,N_11190,N_11405);
and U12768 (N_12768,N_11106,N_12044);
nor U12769 (N_12769,N_12220,N_10053);
nand U12770 (N_12770,N_10251,N_12367);
xnor U12771 (N_12771,N_10813,N_10900);
nand U12772 (N_12772,N_12248,N_10515);
and U12773 (N_12773,N_10806,N_12480);
xor U12774 (N_12774,N_10394,N_11314);
or U12775 (N_12775,N_10688,N_11628);
nor U12776 (N_12776,N_11393,N_12453);
nor U12777 (N_12777,N_11917,N_12439);
and U12778 (N_12778,N_10667,N_11345);
nor U12779 (N_12779,N_11294,N_11762);
nor U12780 (N_12780,N_11222,N_11145);
and U12781 (N_12781,N_12416,N_11369);
or U12782 (N_12782,N_10514,N_11497);
and U12783 (N_12783,N_12119,N_10440);
xnor U12784 (N_12784,N_10599,N_10469);
and U12785 (N_12785,N_11132,N_11558);
nand U12786 (N_12786,N_11627,N_10160);
nand U12787 (N_12787,N_11973,N_12488);
and U12788 (N_12788,N_10935,N_12010);
nor U12789 (N_12789,N_10200,N_11289);
or U12790 (N_12790,N_11151,N_11127);
or U12791 (N_12791,N_11768,N_11018);
xnor U12792 (N_12792,N_11734,N_10449);
xnor U12793 (N_12793,N_11777,N_10128);
and U12794 (N_12794,N_11914,N_10521);
or U12795 (N_12795,N_10589,N_12311);
or U12796 (N_12796,N_11109,N_10529);
or U12797 (N_12797,N_10987,N_12085);
nand U12798 (N_12798,N_10735,N_10868);
xor U12799 (N_12799,N_10441,N_11240);
nor U12800 (N_12800,N_11398,N_11039);
xnor U12801 (N_12801,N_10564,N_11573);
nand U12802 (N_12802,N_10109,N_12057);
xnor U12803 (N_12803,N_11133,N_12383);
nand U12804 (N_12804,N_10366,N_12451);
nand U12805 (N_12805,N_10512,N_10896);
nand U12806 (N_12806,N_10037,N_10502);
or U12807 (N_12807,N_10099,N_11998);
xnor U12808 (N_12808,N_10991,N_10882);
nor U12809 (N_12809,N_12104,N_11430);
nand U12810 (N_12810,N_10981,N_11589);
nor U12811 (N_12811,N_10262,N_11739);
and U12812 (N_12812,N_10795,N_10225);
xnor U12813 (N_12813,N_10465,N_10257);
nand U12814 (N_12814,N_10742,N_11157);
or U12815 (N_12815,N_11711,N_10887);
nor U12816 (N_12816,N_11170,N_12455);
nand U12817 (N_12817,N_11091,N_11718);
and U12818 (N_12818,N_10516,N_11960);
xnor U12819 (N_12819,N_10297,N_11233);
or U12820 (N_12820,N_12244,N_10112);
and U12821 (N_12821,N_11612,N_10695);
and U12822 (N_12822,N_11343,N_11427);
or U12823 (N_12823,N_11814,N_10756);
or U12824 (N_12824,N_10216,N_11663);
nor U12825 (N_12825,N_11891,N_12279);
xor U12826 (N_12826,N_12382,N_11785);
or U12827 (N_12827,N_11702,N_10293);
xor U12828 (N_12828,N_11839,N_10428);
nand U12829 (N_12829,N_10781,N_11571);
xor U12830 (N_12830,N_12032,N_11544);
and U12831 (N_12831,N_12006,N_11420);
nor U12832 (N_12832,N_10751,N_12423);
or U12833 (N_12833,N_12001,N_12310);
nor U12834 (N_12834,N_11033,N_12422);
nor U12835 (N_12835,N_10445,N_10614);
or U12836 (N_12836,N_11521,N_11604);
or U12837 (N_12837,N_11695,N_10823);
and U12838 (N_12838,N_10576,N_11118);
nor U12839 (N_12839,N_10633,N_10997);
xnor U12840 (N_12840,N_11246,N_11476);
xnor U12841 (N_12841,N_10915,N_10321);
xor U12842 (N_12842,N_11915,N_11341);
nand U12843 (N_12843,N_11759,N_12031);
or U12844 (N_12844,N_10335,N_10232);
nand U12845 (N_12845,N_11923,N_12121);
and U12846 (N_12846,N_12122,N_10234);
nand U12847 (N_12847,N_12103,N_10371);
xnor U12848 (N_12848,N_11403,N_12307);
and U12849 (N_12849,N_10989,N_11561);
or U12850 (N_12850,N_12318,N_12113);
and U12851 (N_12851,N_10242,N_10498);
xnor U12852 (N_12852,N_10463,N_10717);
xor U12853 (N_12853,N_11746,N_10206);
xnor U12854 (N_12854,N_12008,N_11237);
and U12855 (N_12855,N_10068,N_11054);
xor U12856 (N_12856,N_11472,N_11559);
nand U12857 (N_12857,N_12025,N_11863);
and U12858 (N_12858,N_11332,N_11485);
or U12859 (N_12859,N_11438,N_11967);
xor U12860 (N_12860,N_10705,N_10618);
xor U12861 (N_12861,N_11825,N_10325);
nand U12862 (N_12862,N_10819,N_11657);
or U12863 (N_12863,N_11086,N_11884);
or U12864 (N_12864,N_11056,N_10089);
nor U12865 (N_12865,N_10869,N_10235);
xnor U12866 (N_12866,N_10584,N_10258);
nand U12867 (N_12867,N_10437,N_12139);
nor U12868 (N_12868,N_10279,N_10062);
nand U12869 (N_12869,N_11656,N_11336);
nand U12870 (N_12870,N_11016,N_12420);
nand U12871 (N_12871,N_10587,N_11003);
and U12872 (N_12872,N_11022,N_12172);
xnor U12873 (N_12873,N_12457,N_10581);
nand U12874 (N_12874,N_11225,N_10027);
and U12875 (N_12875,N_10149,N_10533);
nor U12876 (N_12876,N_11925,N_11776);
xor U12877 (N_12877,N_11433,N_12270);
nor U12878 (N_12878,N_10885,N_10992);
nor U12879 (N_12879,N_11936,N_10458);
xnor U12880 (N_12880,N_11569,N_12284);
xnor U12881 (N_12881,N_10910,N_11045);
xor U12882 (N_12882,N_10098,N_11916);
and U12883 (N_12883,N_12347,N_10732);
and U12884 (N_12884,N_10462,N_10776);
or U12885 (N_12885,N_11528,N_10721);
xor U12886 (N_12886,N_10818,N_11607);
nor U12887 (N_12887,N_10485,N_12335);
nand U12888 (N_12888,N_10400,N_11518);
xor U12889 (N_12889,N_11010,N_11047);
nor U12890 (N_12890,N_11907,N_11821);
and U12891 (N_12891,N_12254,N_10284);
or U12892 (N_12892,N_11214,N_11620);
or U12893 (N_12893,N_10134,N_11780);
and U12894 (N_12894,N_10249,N_11066);
and U12895 (N_12895,N_12215,N_11675);
and U12896 (N_12896,N_10927,N_10523);
xnor U12897 (N_12897,N_10045,N_10147);
nor U12898 (N_12898,N_12291,N_11690);
xnor U12899 (N_12899,N_11542,N_11939);
nor U12900 (N_12900,N_11970,N_12021);
xnor U12901 (N_12901,N_10017,N_12487);
and U12902 (N_12902,N_10303,N_12344);
nand U12903 (N_12903,N_10591,N_11775);
and U12904 (N_12904,N_10727,N_11568);
nor U12905 (N_12905,N_10162,N_10973);
nand U12906 (N_12906,N_12059,N_10233);
or U12907 (N_12907,N_10046,N_10703);
xor U12908 (N_12908,N_12043,N_11035);
nor U12909 (N_12909,N_10933,N_12187);
or U12910 (N_12910,N_10164,N_10944);
or U12911 (N_12911,N_11662,N_10610);
nor U12912 (N_12912,N_10956,N_11602);
xor U12913 (N_12913,N_12265,N_10375);
xor U12914 (N_12914,N_12110,N_11445);
xnor U12915 (N_12915,N_10978,N_11102);
and U12916 (N_12916,N_11212,N_10229);
nor U12917 (N_12917,N_12403,N_12167);
and U12918 (N_12918,N_11007,N_11930);
nor U12919 (N_12919,N_10192,N_11064);
nor U12920 (N_12920,N_11383,N_10385);
and U12921 (N_12921,N_10929,N_10415);
or U12922 (N_12922,N_11432,N_11790);
nand U12923 (N_12923,N_11954,N_11535);
xnor U12924 (N_12924,N_10141,N_11619);
nor U12925 (N_12925,N_11783,N_10539);
xor U12926 (N_12926,N_11577,N_11630);
xor U12927 (N_12927,N_10305,N_10026);
or U12928 (N_12928,N_10368,N_11811);
nor U12929 (N_12929,N_10713,N_10395);
and U12930 (N_12930,N_11387,N_10604);
xor U12931 (N_12931,N_11397,N_11050);
xnor U12932 (N_12932,N_10203,N_10668);
xnor U12933 (N_12933,N_10672,N_12175);
xor U12934 (N_12934,N_10318,N_10107);
and U12935 (N_12935,N_11115,N_11261);
nor U12936 (N_12936,N_10195,N_11719);
and U12937 (N_12937,N_10940,N_12332);
or U12938 (N_12938,N_11042,N_11046);
nor U12939 (N_12939,N_11714,N_10383);
nand U12940 (N_12940,N_10714,N_10548);
nand U12941 (N_12941,N_10349,N_11402);
or U12942 (N_12942,N_10986,N_11361);
or U12943 (N_12943,N_11880,N_12219);
nor U12944 (N_12944,N_10816,N_11323);
and U12945 (N_12945,N_10622,N_12199);
or U12946 (N_12946,N_12205,N_11671);
xnor U12947 (N_12947,N_10774,N_10950);
nand U12948 (N_12948,N_10525,N_12247);
nor U12949 (N_12949,N_10918,N_10047);
or U12950 (N_12950,N_10624,N_11736);
nand U12951 (N_12951,N_10669,N_10985);
xnor U12952 (N_12952,N_10488,N_10559);
nand U12953 (N_12953,N_11131,N_11478);
or U12954 (N_12954,N_11827,N_10686);
or U12955 (N_12955,N_12253,N_10865);
xnor U12956 (N_12956,N_11778,N_11726);
nor U12957 (N_12957,N_10088,N_11517);
and U12958 (N_12958,N_10676,N_10001);
nand U12959 (N_12959,N_12118,N_10308);
or U12960 (N_12960,N_10916,N_10352);
nor U12961 (N_12961,N_12145,N_11585);
nor U12962 (N_12962,N_10500,N_11933);
or U12963 (N_12963,N_11652,N_10186);
nand U12964 (N_12964,N_12000,N_10425);
or U12965 (N_12965,N_10511,N_10577);
or U12966 (N_12966,N_10600,N_10372);
xnor U12967 (N_12967,N_11644,N_10808);
or U12968 (N_12968,N_10606,N_10414);
nor U12969 (N_12969,N_12095,N_11812);
nand U12970 (N_12970,N_11587,N_12421);
xnor U12971 (N_12971,N_12232,N_12479);
nand U12972 (N_12972,N_10557,N_10590);
and U12973 (N_12973,N_12263,N_11892);
and U12974 (N_12974,N_12045,N_10175);
and U12975 (N_12975,N_12174,N_11554);
nor U12976 (N_12976,N_12233,N_10426);
and U12977 (N_12977,N_11024,N_10926);
nand U12978 (N_12978,N_11522,N_11859);
nand U12979 (N_12979,N_11371,N_11494);
xnor U12980 (N_12980,N_11748,N_10749);
and U12981 (N_12981,N_10272,N_12384);
nor U12982 (N_12982,N_10597,N_11841);
xnor U12983 (N_12983,N_10660,N_11443);
xor U12984 (N_12984,N_10680,N_11694);
and U12985 (N_12985,N_11731,N_11624);
xnor U12986 (N_12986,N_11871,N_10811);
or U12987 (N_12987,N_12496,N_11281);
nand U12988 (N_12988,N_11421,N_10048);
xor U12989 (N_12989,N_10184,N_11723);
xnor U12990 (N_12990,N_12298,N_12321);
nand U12991 (N_12991,N_11092,N_11717);
nor U12992 (N_12992,N_10009,N_12385);
or U12993 (N_12993,N_12485,N_10351);
nor U12994 (N_12994,N_11423,N_10778);
nor U12995 (N_12995,N_10775,N_11838);
and U12996 (N_12996,N_11474,N_11163);
and U12997 (N_12997,N_10870,N_11020);
xor U12998 (N_12998,N_12117,N_10457);
and U12999 (N_12999,N_11579,N_10975);
nand U13000 (N_13000,N_10326,N_11489);
and U13001 (N_13001,N_12267,N_10562);
xor U13002 (N_13002,N_10434,N_11834);
nor U13003 (N_13003,N_10355,N_11796);
nand U13004 (N_13004,N_11173,N_10020);
nor U13005 (N_13005,N_10876,N_11987);
nand U13006 (N_13006,N_10132,N_11114);
nor U13007 (N_13007,N_10448,N_12105);
and U13008 (N_13008,N_11547,N_11949);
or U13009 (N_13009,N_11755,N_12098);
xnor U13010 (N_13010,N_10433,N_11282);
nor U13011 (N_13011,N_12231,N_10479);
nand U13012 (N_13012,N_10619,N_11360);
nand U13013 (N_13013,N_12151,N_11647);
xor U13014 (N_13014,N_11805,N_11055);
xnor U13015 (N_13015,N_11991,N_10826);
nand U13016 (N_13016,N_12168,N_12304);
nor U13017 (N_13017,N_11330,N_11760);
or U13018 (N_13018,N_11287,N_12404);
or U13019 (N_13019,N_11431,N_12313);
xnor U13020 (N_13020,N_10103,N_11306);
xor U13021 (N_13021,N_10711,N_11094);
or U13022 (N_13022,N_11333,N_10844);
nor U13023 (N_13023,N_11951,N_12039);
nand U13024 (N_13024,N_11390,N_10911);
xor U13025 (N_13025,N_11231,N_12180);
or U13026 (N_13026,N_10924,N_11197);
or U13027 (N_13027,N_11006,N_11756);
xor U13028 (N_13028,N_10174,N_11781);
nand U13029 (N_13029,N_12337,N_10477);
nand U13030 (N_13030,N_10090,N_10274);
xnor U13031 (N_13031,N_10044,N_10131);
nor U13032 (N_13032,N_12426,N_10421);
nor U13033 (N_13033,N_12188,N_11272);
and U13034 (N_13034,N_11216,N_10708);
xor U13035 (N_13035,N_10389,N_10023);
nor U13036 (N_13036,N_10881,N_10431);
nor U13037 (N_13037,N_11082,N_10850);
and U13038 (N_13038,N_12079,N_11770);
nor U13039 (N_13039,N_12357,N_10336);
nand U13040 (N_13040,N_10211,N_10999);
and U13041 (N_13041,N_11315,N_10616);
nor U13042 (N_13042,N_12309,N_10227);
and U13043 (N_13043,N_11552,N_11110);
nand U13044 (N_13044,N_11364,N_11725);
nor U13045 (N_13045,N_11803,N_10628);
nor U13046 (N_13046,N_10052,N_12281);
nor U13047 (N_13047,N_10265,N_10471);
or U13048 (N_13048,N_10379,N_11757);
or U13049 (N_13049,N_10487,N_11477);
xor U13050 (N_13050,N_12250,N_10738);
nand U13051 (N_13051,N_11291,N_12170);
and U13052 (N_13052,N_12373,N_10642);
xnor U13053 (N_13053,N_12050,N_11910);
xor U13054 (N_13054,N_10946,N_11615);
and U13055 (N_13055,N_12124,N_12070);
and U13056 (N_13056,N_12327,N_10977);
or U13057 (N_13057,N_10061,N_10757);
nor U13058 (N_13058,N_10889,N_12202);
or U13059 (N_13059,N_11034,N_10853);
nand U13060 (N_13060,N_10042,N_11928);
xnor U13061 (N_13061,N_10315,N_10565);
nor U13062 (N_13062,N_10842,N_10930);
nor U13063 (N_13063,N_11404,N_11188);
xnor U13064 (N_13064,N_12186,N_11833);
nor U13065 (N_13065,N_11600,N_11672);
nor U13066 (N_13066,N_10033,N_11856);
xor U13067 (N_13067,N_10745,N_11174);
and U13068 (N_13068,N_12317,N_11932);
or U13069 (N_13069,N_12409,N_11011);
or U13070 (N_13070,N_10087,N_11002);
nand U13071 (N_13071,N_10726,N_10248);
and U13072 (N_13072,N_11649,N_12331);
xor U13073 (N_13073,N_11782,N_11267);
nand U13074 (N_13074,N_10051,N_10645);
or U13075 (N_13075,N_10028,N_11921);
and U13076 (N_13076,N_10144,N_10110);
xnor U13077 (N_13077,N_11288,N_11080);
xor U13078 (N_13078,N_12094,N_11870);
or U13079 (N_13079,N_11177,N_11758);
or U13080 (N_13080,N_11389,N_11986);
and U13081 (N_13081,N_10832,N_11835);
nand U13082 (N_13082,N_10219,N_11276);
or U13083 (N_13083,N_12481,N_11511);
and U13084 (N_13084,N_11463,N_11865);
xnor U13085 (N_13085,N_12075,N_12179);
or U13086 (N_13086,N_10678,N_12037);
nor U13087 (N_13087,N_11381,N_11202);
xor U13088 (N_13088,N_12464,N_11691);
and U13089 (N_13089,N_11848,N_10953);
xor U13090 (N_13090,N_10724,N_11000);
and U13091 (N_13091,N_10629,N_10650);
nor U13092 (N_13092,N_12431,N_12022);
xor U13093 (N_13093,N_10838,N_10541);
or U13094 (N_13094,N_11794,N_11971);
or U13095 (N_13095,N_10538,N_11486);
or U13096 (N_13096,N_11570,N_11353);
and U13097 (N_13097,N_10077,N_12312);
xnor U13098 (N_13098,N_11312,N_12091);
nand U13099 (N_13099,N_11643,N_11185);
nand U13100 (N_13100,N_12303,N_11621);
or U13101 (N_13101,N_12074,N_10436);
or U13102 (N_13102,N_10331,N_12407);
xor U13103 (N_13103,N_10884,N_10769);
nor U13104 (N_13104,N_10354,N_10015);
or U13105 (N_13105,N_11502,N_11849);
nor U13106 (N_13106,N_11908,N_12365);
or U13107 (N_13107,N_11290,N_11480);
and U13108 (N_13108,N_11860,N_11204);
nor U13109 (N_13109,N_12412,N_10875);
xor U13110 (N_13110,N_10785,N_11311);
and U13111 (N_13111,N_11560,N_10035);
and U13112 (N_13112,N_10960,N_10817);
nand U13113 (N_13113,N_11461,N_10171);
xnor U13114 (N_13114,N_10631,N_10029);
and U13115 (N_13115,N_10990,N_10187);
and U13116 (N_13116,N_10575,N_10456);
and U13117 (N_13117,N_10063,N_10964);
xor U13118 (N_13118,N_10571,N_12486);
nand U13119 (N_13119,N_10596,N_10729);
and U13120 (N_13120,N_11191,N_10720);
and U13121 (N_13121,N_10701,N_11221);
nor U13122 (N_13122,N_10137,N_12055);
xor U13123 (N_13123,N_11693,N_10317);
nand U13124 (N_13124,N_10984,N_12120);
or U13125 (N_13125,N_10022,N_10988);
xnor U13126 (N_13126,N_11031,N_11912);
nor U13127 (N_13127,N_12379,N_10942);
xnor U13128 (N_13128,N_10494,N_10150);
nand U13129 (N_13129,N_10261,N_11641);
nor U13130 (N_13130,N_11036,N_11779);
or U13131 (N_13131,N_10300,N_12443);
xnor U13132 (N_13132,N_11334,N_11374);
and U13133 (N_13133,N_11958,N_12366);
or U13134 (N_13134,N_11206,N_12458);
or U13135 (N_13135,N_10743,N_11491);
nand U13136 (N_13136,N_11515,N_12020);
and U13137 (N_13137,N_12346,N_10169);
xor U13138 (N_13138,N_11025,N_11703);
or U13139 (N_13139,N_10182,N_10734);
and U13140 (N_13140,N_10550,N_11873);
nor U13141 (N_13141,N_12015,N_11660);
xnor U13142 (N_13142,N_11139,N_11578);
or U13143 (N_13143,N_11407,N_11382);
and U13144 (N_13144,N_11843,N_11868);
nor U13145 (N_13145,N_11553,N_10032);
or U13146 (N_13146,N_11505,N_12434);
or U13147 (N_13147,N_11178,N_10526);
or U13148 (N_13148,N_10954,N_11588);
xnor U13149 (N_13149,N_10084,N_12097);
nand U13150 (N_13150,N_11500,N_11629);
nand U13151 (N_13151,N_11979,N_11256);
nor U13152 (N_13152,N_11898,N_12389);
xor U13153 (N_13153,N_11678,N_12438);
xor U13154 (N_13154,N_12153,N_11989);
and U13155 (N_13155,N_11852,N_11243);
and U13156 (N_13156,N_11302,N_11263);
and U13157 (N_13157,N_11400,N_11533);
and U13158 (N_13158,N_10210,N_10016);
xnor U13159 (N_13159,N_10513,N_11523);
and U13160 (N_13160,N_10447,N_11090);
and U13161 (N_13161,N_12030,N_10292);
nor U13162 (N_13162,N_12087,N_10283);
nand U13163 (N_13163,N_10191,N_11058);
or U13164 (N_13164,N_10789,N_10417);
and U13165 (N_13165,N_10056,N_12354);
nor U13166 (N_13166,N_10340,N_10423);
nand U13167 (N_13167,N_11980,N_10652);
nor U13168 (N_13168,N_10082,N_10205);
and U13169 (N_13169,N_12093,N_12414);
nand U13170 (N_13170,N_10364,N_11228);
or U13171 (N_13171,N_10834,N_11653);
or U13172 (N_13172,N_12014,N_10847);
and U13173 (N_13173,N_11450,N_11999);
xnor U13174 (N_13174,N_12213,N_11574);
nand U13175 (N_13175,N_11667,N_10563);
nand U13176 (N_13176,N_11129,N_12356);
nor U13177 (N_13177,N_12084,N_11688);
or U13178 (N_13178,N_11380,N_10490);
and U13179 (N_13179,N_11504,N_10097);
xor U13180 (N_13180,N_11292,N_10552);
and U13181 (N_13181,N_12046,N_10424);
and U13182 (N_13182,N_10830,N_12463);
nand U13183 (N_13183,N_12177,N_11944);
or U13184 (N_13184,N_11674,N_11854);
nor U13185 (N_13185,N_10118,N_11363);
nand U13186 (N_13186,N_11531,N_10856);
and U13187 (N_13187,N_10530,N_10078);
or U13188 (N_13188,N_11706,N_10670);
and U13189 (N_13189,N_11767,N_11162);
and U13190 (N_13190,N_11743,N_12063);
nor U13191 (N_13191,N_11088,N_12049);
and U13192 (N_13192,N_12169,N_10993);
xnor U13193 (N_13193,N_10615,N_10925);
or U13194 (N_13194,N_11008,N_11112);
nand U13195 (N_13195,N_11249,N_12068);
and U13196 (N_13196,N_11851,N_12252);
nand U13197 (N_13197,N_11963,N_11169);
nand U13198 (N_13198,N_12214,N_11707);
xnor U13199 (N_13199,N_11680,N_11614);
nand U13200 (N_13200,N_10694,N_10255);
xor U13201 (N_13201,N_11506,N_11829);
nor U13202 (N_13202,N_12143,N_11540);
or U13203 (N_13203,N_12360,N_11295);
xor U13204 (N_13204,N_11043,N_10360);
or U13205 (N_13205,N_10677,N_10827);
and U13206 (N_13206,N_11150,N_12058);
nand U13207 (N_13207,N_11298,N_10923);
nor U13208 (N_13208,N_12348,N_10784);
or U13209 (N_13209,N_10367,N_10193);
and U13210 (N_13210,N_10254,N_11026);
nor U13211 (N_13211,N_11137,N_11346);
and U13212 (N_13212,N_10259,N_11342);
xor U13213 (N_13213,N_10289,N_12080);
and U13214 (N_13214,N_12280,N_10130);
and U13215 (N_13215,N_11525,N_12370);
nor U13216 (N_13216,N_10648,N_10871);
xor U13217 (N_13217,N_11310,N_12200);
nor U13218 (N_13218,N_12221,N_10715);
nand U13219 (N_13219,N_11747,N_10763);
and U13220 (N_13220,N_12336,N_11180);
and U13221 (N_13221,N_10113,N_11823);
xnor U13222 (N_13222,N_10106,N_10654);
nand U13223 (N_13223,N_10172,N_11877);
and U13224 (N_13224,N_11096,N_10524);
xnor U13225 (N_13225,N_11943,N_11665);
or U13226 (N_13226,N_11609,N_10152);
or U13227 (N_13227,N_11099,N_10059);
and U13228 (N_13228,N_11595,N_11327);
or U13229 (N_13229,N_10947,N_10427);
xnor U13230 (N_13230,N_11409,N_11982);
nand U13231 (N_13231,N_10240,N_11156);
and U13232 (N_13232,N_12225,N_12374);
and U13233 (N_13233,N_11926,N_10815);
nand U13234 (N_13234,N_10673,N_12054);
or U13235 (N_13235,N_11049,N_10114);
and U13236 (N_13236,N_11095,N_11004);
nor U13237 (N_13237,N_11078,N_10021);
or U13238 (N_13238,N_12449,N_10075);
or U13239 (N_13239,N_11207,N_12242);
nor U13240 (N_13240,N_12183,N_12363);
nor U13241 (N_13241,N_10542,N_11209);
xor U13242 (N_13242,N_10000,N_10790);
xor U13243 (N_13243,N_10536,N_12460);
xnor U13244 (N_13244,N_12035,N_11422);
and U13245 (N_13245,N_10545,N_12206);
nand U13246 (N_13246,N_10104,N_10851);
or U13247 (N_13247,N_10903,N_10495);
and U13248 (N_13248,N_11449,N_11769);
and U13249 (N_13249,N_11027,N_11858);
nor U13250 (N_13250,N_12072,N_10069);
xor U13251 (N_13251,N_11813,N_10065);
and U13252 (N_13252,N_11800,N_11470);
and U13253 (N_13253,N_11705,N_12372);
nand U13254 (N_13254,N_12012,N_10702);
xor U13255 (N_13255,N_11845,N_10486);
or U13256 (N_13256,N_11572,N_12358);
nor U13257 (N_13257,N_12315,N_11123);
xnor U13258 (N_13258,N_12495,N_10854);
and U13259 (N_13259,N_11866,N_10072);
nor U13260 (N_13260,N_11179,N_10585);
xor U13261 (N_13261,N_12061,N_12162);
or U13262 (N_13262,N_11418,N_10613);
nand U13263 (N_13263,N_11040,N_10468);
xnor U13264 (N_13264,N_12160,N_11495);
nand U13265 (N_13265,N_10855,N_10547);
nand U13266 (N_13266,N_11881,N_10387);
nand U13267 (N_13267,N_12489,N_10181);
or U13268 (N_13268,N_12123,N_10085);
or U13269 (N_13269,N_10731,N_10142);
xnor U13270 (N_13270,N_10074,N_12440);
nand U13271 (N_13271,N_11766,N_10974);
xnor U13272 (N_13272,N_11229,N_12408);
or U13273 (N_13273,N_10812,N_11462);
and U13274 (N_13274,N_11855,N_12424);
and U13275 (N_13275,N_10398,N_10482);
xnor U13276 (N_13276,N_11253,N_11019);
or U13277 (N_13277,N_10612,N_11304);
or U13278 (N_13278,N_11842,N_11072);
xnor U13279 (N_13279,N_10196,N_12013);
nor U13280 (N_13280,N_11236,N_12323);
nand U13281 (N_13281,N_11715,N_10380);
and U13282 (N_13282,N_10011,N_10190);
nor U13283 (N_13283,N_10276,N_10476);
nand U13284 (N_13284,N_11689,N_10888);
nand U13285 (N_13285,N_10050,N_10707);
or U13286 (N_13286,N_10167,N_10399);
nand U13287 (N_13287,N_10040,N_11143);
or U13288 (N_13288,N_10836,N_10822);
nand U13289 (N_13289,N_12234,N_10733);
or U13290 (N_13290,N_10277,N_10108);
and U13291 (N_13291,N_12150,N_10568);
nand U13292 (N_13292,N_11172,N_10008);
or U13293 (N_13293,N_12478,N_10746);
or U13294 (N_13294,N_12456,N_12164);
or U13295 (N_13295,N_10094,N_11648);
or U13296 (N_13296,N_10133,N_10179);
or U13297 (N_13297,N_10119,N_11200);
or U13298 (N_13298,N_11444,N_12328);
and U13299 (N_13299,N_11230,N_12134);
nand U13300 (N_13300,N_10329,N_11738);
or U13301 (N_13301,N_10800,N_11285);
and U13302 (N_13302,N_10840,N_12268);
nor U13303 (N_13303,N_12282,N_10116);
nor U13304 (N_13304,N_12399,N_10857);
nor U13305 (N_13305,N_11716,N_12245);
or U13306 (N_13306,N_10553,N_11720);
or U13307 (N_13307,N_11632,N_12308);
xnor U13308 (N_13308,N_11836,N_10307);
or U13309 (N_13309,N_10226,N_11005);
xor U13310 (N_13310,N_11961,N_11940);
or U13311 (N_13311,N_10122,N_11874);
and U13312 (N_13312,N_12471,N_11001);
or U13313 (N_13313,N_12406,N_10799);
or U13314 (N_13314,N_11359,N_11062);
nand U13315 (N_13315,N_10643,N_11697);
and U13316 (N_13316,N_12101,N_12288);
xor U13317 (N_13317,N_10013,N_11784);
nor U13318 (N_13318,N_11069,N_10221);
xor U13319 (N_13319,N_10125,N_10388);
xnor U13320 (N_13320,N_10328,N_11937);
xnor U13321 (N_13321,N_11159,N_10998);
xnor U13322 (N_13322,N_11959,N_10788);
or U13323 (N_13323,N_11582,N_12226);
nor U13324 (N_13324,N_10835,N_11183);
xnor U13325 (N_13325,N_12392,N_12418);
xor U13326 (N_13326,N_10753,N_10138);
nor U13327 (N_13327,N_11293,N_11084);
nor U13328 (N_13328,N_12184,N_12131);
and U13329 (N_13329,N_11512,N_10522);
nand U13330 (N_13330,N_12386,N_11417);
and U13331 (N_13331,N_11370,N_12452);
and U13332 (N_13332,N_11957,N_12243);
xor U13333 (N_13333,N_11900,N_11148);
nor U13334 (N_13334,N_10378,N_12351);
nand U13335 (N_13335,N_12157,N_10766);
and U13336 (N_13336,N_12194,N_12038);
nand U13337 (N_13337,N_11659,N_10638);
nor U13338 (N_13338,N_11030,N_10270);
nor U13339 (N_13339,N_10260,N_10217);
xor U13340 (N_13340,N_11976,N_12144);
xor U13341 (N_13341,N_10228,N_10339);
nand U13342 (N_13342,N_10197,N_11503);
and U13343 (N_13343,N_11377,N_12051);
nor U13344 (N_13344,N_10041,N_10535);
or U13345 (N_13345,N_11750,N_10492);
xor U13346 (N_13346,N_12325,N_11149);
nor U13347 (N_13347,N_10573,N_10952);
nor U13348 (N_13348,N_11651,N_10664);
nor U13349 (N_13349,N_12129,N_11268);
nor U13350 (N_13350,N_12275,N_10828);
nor U13351 (N_13351,N_10401,N_10239);
or U13352 (N_13352,N_12166,N_10327);
xor U13353 (N_13353,N_11817,N_10402);
and U13354 (N_13354,N_10748,N_12342);
nor U13355 (N_13355,N_11367,N_11154);
xor U13356 (N_13356,N_10567,N_12089);
and U13357 (N_13357,N_11372,N_12158);
nor U13358 (N_13358,N_11721,N_12343);
and U13359 (N_13359,N_11795,N_10907);
or U13360 (N_13360,N_10031,N_10135);
nand U13361 (N_13361,N_10518,N_11442);
nand U13362 (N_13362,N_11640,N_10096);
or U13363 (N_13363,N_11104,N_11247);
xnor U13364 (N_13364,N_10655,N_12330);
and U13365 (N_13365,N_10178,N_11565);
xor U13366 (N_13366,N_11466,N_11279);
and U13367 (N_13367,N_12003,N_10018);
and U13368 (N_13368,N_10659,N_11220);
nor U13369 (N_13369,N_12338,N_12071);
and U13370 (N_13370,N_10920,N_11847);
nand U13371 (N_13371,N_11023,N_12228);
and U13372 (N_13372,N_11802,N_10843);
nor U13373 (N_13373,N_11475,N_10955);
xnor U13374 (N_13374,N_12100,N_11889);
xnor U13375 (N_13375,N_10802,N_10244);
xor U13376 (N_13376,N_12353,N_11735);
nand U13377 (N_13377,N_11277,N_11994);
nand U13378 (N_13378,N_12425,N_10208);
nor U13379 (N_13379,N_11325,N_10833);
and U13380 (N_13380,N_10747,N_11428);
and U13381 (N_13381,N_11138,N_11140);
or U13382 (N_13382,N_11622,N_11899);
or U13383 (N_13383,N_11224,N_11820);
or U13384 (N_13384,N_11319,N_12429);
and U13385 (N_13385,N_10304,N_10653);
or U13386 (N_13386,N_12273,N_11911);
xor U13387 (N_13387,N_11406,N_10365);
xor U13388 (N_13388,N_10081,N_11551);
xor U13389 (N_13389,N_11977,N_11328);
nor U13390 (N_13390,N_10831,N_11819);
nand U13391 (N_13391,N_11549,N_10237);
or U13392 (N_13392,N_11073,N_11520);
xor U13393 (N_13393,N_11386,N_12387);
and U13394 (N_13394,N_11670,N_10780);
nor U13395 (N_13395,N_11879,N_11168);
xnor U13396 (N_13396,N_10036,N_12258);
xor U13397 (N_13397,N_10603,N_11021);
and U13398 (N_13398,N_10268,N_10202);
or U13399 (N_13399,N_10454,N_11683);
nor U13400 (N_13400,N_11473,N_11175);
nand U13401 (N_13401,N_10357,N_12368);
xnor U13402 (N_13402,N_10464,N_11929);
nor U13403 (N_13403,N_12260,N_10761);
and U13404 (N_13404,N_11809,N_10723);
or U13405 (N_13405,N_12266,N_12290);
and U13406 (N_13406,N_10435,N_12436);
and U13407 (N_13407,N_11564,N_10246);
or U13408 (N_13408,N_12249,N_10100);
and U13409 (N_13409,N_11862,N_10740);
nor U13410 (N_13410,N_10231,N_10661);
xnor U13411 (N_13411,N_10264,N_12161);
nor U13412 (N_13412,N_10043,N_12314);
nor U13413 (N_13413,N_10852,N_12096);
or U13414 (N_13414,N_10864,N_10411);
nand U13415 (N_13415,N_10690,N_11165);
nand U13416 (N_13416,N_10647,N_10102);
xor U13417 (N_13417,N_11079,N_11067);
nor U13418 (N_13418,N_11322,N_11864);
and U13419 (N_13419,N_12251,N_11448);
or U13420 (N_13420,N_11853,N_10872);
xnor U13421 (N_13421,N_11744,N_11876);
xor U13422 (N_13422,N_11771,N_10263);
and U13423 (N_13423,N_12498,N_11068);
nand U13424 (N_13424,N_10286,N_10949);
and U13425 (N_13425,N_11984,N_12140);
or U13426 (N_13426,N_11633,N_12380);
nand U13427 (N_13427,N_10601,N_12193);
xor U13428 (N_13428,N_11872,N_11920);
or U13429 (N_13429,N_12300,N_11116);
and U13430 (N_13430,N_11798,N_10377);
nand U13431 (N_13431,N_10737,N_10569);
nand U13432 (N_13432,N_12428,N_11108);
nor U13433 (N_13433,N_10945,N_12350);
and U13434 (N_13434,N_10906,N_12239);
nand U13435 (N_13435,N_11687,N_11232);
or U13436 (N_13436,N_11642,N_11286);
nand U13437 (N_13437,N_11447,N_12141);
xnor U13438 (N_13438,N_10461,N_10928);
and U13439 (N_13439,N_10393,N_11227);
nor U13440 (N_13440,N_11250,N_10886);
xor U13441 (N_13441,N_10879,N_11469);
or U13442 (N_13442,N_11484,N_10909);
xor U13443 (N_13443,N_10958,N_11365);
and U13444 (N_13444,N_10294,N_10275);
nor U13445 (N_13445,N_11661,N_10267);
or U13446 (N_13446,N_11437,N_10384);
nor U13447 (N_13447,N_10145,N_12467);
or U13448 (N_13448,N_12152,N_11061);
and U13449 (N_13449,N_11882,N_11664);
nand U13450 (N_13450,N_10342,N_10129);
or U13451 (N_13451,N_10359,N_10373);
nand U13452 (N_13452,N_11394,N_12329);
or U13453 (N_13453,N_11459,N_12292);
or U13454 (N_13454,N_10376,N_12149);
and U13455 (N_13455,N_12364,N_11787);
nor U13456 (N_13456,N_11135,N_10510);
or U13457 (N_13457,N_10159,N_10593);
xnor U13458 (N_13458,N_10758,N_12107);
nand U13459 (N_13459,N_11317,N_11122);
xor U13460 (N_13460,N_12126,N_11883);
and U13461 (N_13461,N_12324,N_11098);
nor U13462 (N_13462,N_10319,N_12264);
xor U13463 (N_13463,N_12238,N_11464);
nand U13464 (N_13464,N_12106,N_11065);
or U13465 (N_13465,N_11187,N_12499);
xor U13466 (N_13466,N_12203,N_11763);
nand U13467 (N_13467,N_11435,N_10961);
xnor U13468 (N_13468,N_10410,N_10938);
xor U13469 (N_13469,N_11897,N_12237);
or U13470 (N_13470,N_12083,N_10636);
or U13471 (N_13471,N_10346,N_11303);
or U13472 (N_13472,N_10994,N_10146);
xnor U13473 (N_13473,N_10917,N_11210);
nor U13474 (N_13474,N_10030,N_11828);
or U13475 (N_13475,N_11995,N_11195);
xor U13476 (N_13476,N_10858,N_10290);
xnor U13477 (N_13477,N_12163,N_10810);
or U13478 (N_13478,N_10101,N_11635);
and U13479 (N_13479,N_10651,N_11597);
or U13480 (N_13480,N_12028,N_11792);
nor U13481 (N_13481,N_10452,N_10139);
or U13482 (N_13482,N_11416,N_10632);
nor U13483 (N_13483,N_12067,N_10543);
nor U13484 (N_13484,N_11117,N_11278);
nand U13485 (N_13485,N_12209,N_11456);
and U13486 (N_13486,N_11950,N_10322);
xnor U13487 (N_13487,N_12462,N_11141);
or U13488 (N_13488,N_10508,N_12240);
nand U13489 (N_13489,N_12296,N_10213);
nand U13490 (N_13490,N_11799,N_12036);
or U13491 (N_13491,N_10250,N_11886);
nor U13492 (N_13492,N_10637,N_12171);
and U13493 (N_13493,N_10121,N_10586);
nor U13494 (N_13494,N_10071,N_12011);
or U13495 (N_13495,N_11051,N_10621);
nor U13496 (N_13496,N_11545,N_10049);
and U13497 (N_13497,N_11425,N_11636);
or U13498 (N_13498,N_12026,N_11867);
and U13499 (N_13499,N_11618,N_12040);
or U13500 (N_13500,N_12395,N_10310);
and U13501 (N_13501,N_10467,N_11786);
or U13502 (N_13502,N_11815,N_11198);
nor U13503 (N_13503,N_12466,N_10348);
or U13504 (N_13504,N_12114,N_12257);
nand U13505 (N_13505,N_10880,N_10198);
or U13506 (N_13506,N_12217,N_10649);
or U13507 (N_13507,N_12289,N_10252);
and U13508 (N_13508,N_11580,N_11347);
or U13509 (N_13509,N_10683,N_10689);
nand U13510 (N_13510,N_11184,N_10505);
nand U13511 (N_13511,N_10767,N_12066);
nand U13512 (N_13512,N_11791,N_11089);
nand U13513 (N_13513,N_10460,N_11591);
or U13514 (N_13514,N_10777,N_10982);
nor U13515 (N_13515,N_12201,N_10218);
or U13516 (N_13516,N_10157,N_11083);
nand U13517 (N_13517,N_10640,N_11728);
nor U13518 (N_13518,N_11645,N_11988);
and U13519 (N_13519,N_12023,N_10222);
or U13520 (N_13520,N_11063,N_11362);
or U13521 (N_13521,N_12345,N_11273);
or U13522 (N_13522,N_10867,N_10501);
and U13523 (N_13523,N_10223,N_12230);
or U13524 (N_13524,N_11155,N_10470);
nor U13525 (N_13525,N_10837,N_11918);
xnor U13526 (N_13526,N_11878,N_10489);
nand U13527 (N_13527,N_10243,N_12469);
xnor U13528 (N_13528,N_11966,N_10422);
nor U13529 (N_13529,N_11457,N_10472);
and U13530 (N_13530,N_11301,N_10666);
xor U13531 (N_13531,N_10507,N_11375);
xor U13532 (N_13532,N_10641,N_10544);
nor U13533 (N_13533,N_10381,N_11384);
xor U13534 (N_13534,N_12285,N_11320);
xor U13535 (N_13535,N_11534,N_12189);
and U13536 (N_13536,N_11679,N_12148);
nand U13537 (N_13537,N_12176,N_10126);
or U13538 (N_13538,N_11196,N_10725);
or U13539 (N_13539,N_11789,N_11948);
xnor U13540 (N_13540,N_12283,N_11446);
xnor U13541 (N_13541,N_11257,N_10092);
and U13542 (N_13542,N_12132,N_11490);
nand U13543 (N_13543,N_11773,N_10313);
nand U13544 (N_13544,N_10532,N_11945);
nor U13545 (N_13545,N_11356,N_12391);
nor U13546 (N_13546,N_11548,N_11646);
nor U13547 (N_13547,N_10630,N_10220);
or U13548 (N_13548,N_11519,N_11514);
nand U13549 (N_13549,N_12490,N_12297);
xor U13550 (N_13550,N_11526,N_12078);
xor U13551 (N_13551,N_10073,N_11832);
or U13552 (N_13552,N_11454,N_12316);
nor U13553 (N_13553,N_12473,N_10846);
nand U13554 (N_13554,N_11479,N_10658);
and U13555 (N_13555,N_10466,N_10347);
or U13556 (N_13556,N_11161,N_10759);
xnor U13557 (N_13557,N_11194,N_10362);
nor U13558 (N_13558,N_11741,N_10301);
xor U13559 (N_13559,N_10124,N_10848);
and U13560 (N_13560,N_12269,N_11513);
xnor U13561 (N_13561,N_11529,N_10728);
nor U13562 (N_13562,N_10718,N_11905);
xor U13563 (N_13563,N_12062,N_11623);
xor U13564 (N_13564,N_12146,N_11260);
and U13565 (N_13565,N_10968,N_11901);
xor U13566 (N_13566,N_12484,N_11097);
nor U13567 (N_13567,N_10752,N_11153);
nand U13568 (N_13568,N_10579,N_10730);
nor U13569 (N_13569,N_11993,N_11946);
nand U13570 (N_13570,N_12018,N_10161);
or U13571 (N_13571,N_10741,N_11885);
nand U13572 (N_13572,N_11981,N_11234);
xnor U13573 (N_13573,N_11753,N_10003);
nor U13574 (N_13574,N_11598,N_10979);
nor U13575 (N_13575,N_12034,N_10750);
nand U13576 (N_13576,N_10332,N_10841);
xnor U13577 (N_13577,N_12435,N_10429);
nor U13578 (N_13578,N_10937,N_10883);
nor U13579 (N_13579,N_10475,N_10356);
xor U13580 (N_13580,N_10878,N_10809);
nand U13581 (N_13581,N_10675,N_10588);
xnor U13582 (N_13582,N_11284,N_10824);
nand U13583 (N_13583,N_11576,N_11077);
xor U13584 (N_13584,N_10969,N_12415);
or U13585 (N_13585,N_10291,N_12127);
nand U13586 (N_13586,N_11337,N_10405);
and U13587 (N_13587,N_11639,N_10627);
xnor U13588 (N_13588,N_11321,N_11171);
xor U13589 (N_13589,N_10873,N_11378);
nor U13590 (N_13590,N_10546,N_10117);
xor U13591 (N_13591,N_12362,N_10932);
or U13592 (N_13592,N_12454,N_11339);
nand U13593 (N_13593,N_12115,N_11801);
xor U13594 (N_13594,N_11581,N_11070);
or U13595 (N_13595,N_10794,N_11807);
or U13596 (N_13596,N_10123,N_11235);
or U13597 (N_13597,N_11654,N_11053);
nor U13598 (N_13598,N_10635,N_12190);
or U13599 (N_13599,N_10432,N_10418);
and U13600 (N_13600,N_11968,N_11087);
nand U13601 (N_13601,N_11708,N_10302);
nand U13602 (N_13602,N_12224,N_11242);
nor U13603 (N_13603,N_11201,N_12181);
xnor U13604 (N_13604,N_11516,N_11205);
and U13605 (N_13605,N_10306,N_10334);
xor U13606 (N_13606,N_10607,N_11996);
and U13607 (N_13607,N_11093,N_10519);
xor U13608 (N_13608,N_11392,N_10370);
or U13609 (N_13609,N_11749,N_10598);
and U13610 (N_13610,N_11439,N_10803);
or U13611 (N_13611,N_10298,N_10691);
nor U13612 (N_13612,N_11239,N_11586);
or U13613 (N_13613,N_11307,N_12272);
and U13614 (N_13614,N_10148,N_10143);
xor U13615 (N_13615,N_11419,N_12376);
nor U13616 (N_13616,N_12419,N_12410);
and U13617 (N_13617,N_10921,N_11737);
nand U13618 (N_13618,N_11244,N_12009);
nor U13619 (N_13619,N_11956,N_10236);
nand U13620 (N_13620,N_10995,N_10215);
and U13621 (N_13621,N_10060,N_10309);
nor U13622 (N_13622,N_12069,N_10798);
or U13623 (N_13623,N_10768,N_12461);
xnor U13624 (N_13624,N_11071,N_10019);
nor U13625 (N_13625,N_11713,N_11275);
nand U13626 (N_13626,N_10007,N_12004);
nand U13627 (N_13627,N_11413,N_10155);
or U13628 (N_13628,N_10120,N_11296);
or U13629 (N_13629,N_12024,N_12052);
or U13630 (N_13630,N_12341,N_11136);
nand U13631 (N_13631,N_12056,N_11037);
or U13632 (N_13632,N_10238,N_10189);
nand U13633 (N_13633,N_10772,N_11274);
or U13634 (N_13634,N_10744,N_12019);
or U13635 (N_13635,N_10397,N_10682);
and U13636 (N_13636,N_11692,N_10212);
or U13637 (N_13637,N_11830,N_10825);
or U13638 (N_13638,N_11730,N_10570);
nand U13639 (N_13639,N_11935,N_11411);
nand U13640 (N_13640,N_11280,N_12137);
or U13641 (N_13641,N_12442,N_11396);
nor U13642 (N_13642,N_10320,N_12112);
or U13643 (N_13643,N_12073,N_11488);
nand U13644 (N_13644,N_10874,N_12276);
or U13645 (N_13645,N_10201,N_10245);
xnor U13646 (N_13646,N_11556,N_12029);
or U13647 (N_13647,N_10350,N_10764);
or U13648 (N_13648,N_11453,N_11508);
nand U13649 (N_13649,N_12482,N_10438);
xnor U13650 (N_13650,N_11681,N_12173);
or U13651 (N_13651,N_10971,N_11941);
nor U13652 (N_13652,N_11658,N_10247);
or U13653 (N_13653,N_10657,N_11507);
or U13654 (N_13654,N_11305,N_10311);
and U13655 (N_13655,N_11655,N_10439);
nor U13656 (N_13656,N_12483,N_11733);
nor U13657 (N_13657,N_11496,N_12108);
xor U13658 (N_13658,N_12393,N_11340);
nand U13659 (N_13659,N_10314,N_11676);
nand U13660 (N_13660,N_12448,N_11385);
nor U13661 (N_13661,N_10839,N_11105);
nor U13662 (N_13662,N_10420,N_10493);
nor U13663 (N_13663,N_10484,N_12191);
nor U13664 (N_13664,N_11255,N_11368);
xor U13665 (N_13665,N_10214,N_10151);
xor U13666 (N_13666,N_10779,N_11426);
xor U13667 (N_13667,N_11297,N_10416);
xnor U13668 (N_13668,N_10453,N_12446);
or U13669 (N_13669,N_10656,N_10086);
and U13670 (N_13670,N_10154,N_11537);
xor U13671 (N_13671,N_12301,N_11724);
nor U13672 (N_13672,N_11906,N_10224);
xor U13673 (N_13673,N_10951,N_12299);
or U13674 (N_13674,N_11727,N_12208);
and U13675 (N_13675,N_10644,N_11344);
nor U13676 (N_13676,N_11299,N_10408);
nand U13677 (N_13677,N_11990,N_11669);
nand U13678 (N_13678,N_12090,N_11745);
or U13679 (N_13679,N_11509,N_10480);
nand U13680 (N_13680,N_12402,N_11890);
xnor U13681 (N_13681,N_10966,N_10269);
and U13682 (N_13682,N_12430,N_11788);
nor U13683 (N_13683,N_12048,N_11594);
and U13684 (N_13684,N_11410,N_12241);
nand U13685 (N_13685,N_11913,N_11379);
and U13686 (N_13686,N_11947,N_10025);
or U13687 (N_13687,N_10782,N_11041);
xor U13688 (N_13688,N_10443,N_11313);
xor U13689 (N_13689,N_10574,N_11391);
xnor U13690 (N_13690,N_11793,N_10288);
nor U13691 (N_13691,N_11350,N_11761);
xor U13692 (N_13692,N_12472,N_12401);
and U13693 (N_13693,N_12405,N_10787);
nand U13694 (N_13694,N_11599,N_10582);
xor U13695 (N_13695,N_12388,N_10894);
nor U13696 (N_13696,N_12294,N_10444);
nor U13697 (N_13697,N_12133,N_11539);
nor U13698 (N_13698,N_10369,N_10948);
nand U13699 (N_13699,N_12295,N_10083);
nor U13700 (N_13700,N_11181,N_11429);
or U13701 (N_13701,N_11965,N_11824);
or U13702 (N_13702,N_10902,N_12278);
nand U13703 (N_13703,N_10483,N_11563);
and U13704 (N_13704,N_12474,N_10005);
nand U13705 (N_13705,N_11608,N_10166);
nand U13706 (N_13706,N_10455,N_10710);
nor U13707 (N_13707,N_11482,N_10556);
or U13708 (N_13708,N_11326,N_10285);
or U13709 (N_13709,N_11455,N_10057);
nor U13710 (N_13710,N_11972,N_11584);
or U13711 (N_13711,N_11985,N_10931);
xor U13712 (N_13712,N_12099,N_10316);
nor U13713 (N_13713,N_10230,N_11605);
nor U13714 (N_13714,N_10796,N_11258);
xor U13715 (N_13715,N_12005,N_12138);
and U13716 (N_13716,N_12470,N_10671);
nand U13717 (N_13717,N_11358,N_10773);
or U13718 (N_13718,N_11269,N_12076);
or U13719 (N_13719,N_10442,N_10639);
xor U13720 (N_13720,N_10980,N_11451);
and U13721 (N_13721,N_10962,N_10890);
and U13722 (N_13722,N_11888,N_10363);
or U13723 (N_13723,N_10959,N_11567);
nor U13724 (N_13724,N_12355,N_10797);
xnor U13725 (N_13725,N_10386,N_11029);
or U13726 (N_13726,N_11698,N_11226);
nand U13727 (N_13727,N_10409,N_10901);
nor U13728 (N_13728,N_10204,N_11590);
or U13729 (N_13729,N_11218,N_11335);
nand U13730 (N_13730,N_10862,N_10404);
nor U13731 (N_13731,N_12218,N_11119);
nand U13732 (N_13732,N_11048,N_10241);
nand U13733 (N_13733,N_11408,N_11685);
nand U13734 (N_13734,N_10194,N_11219);
or U13735 (N_13735,N_12156,N_11969);
nor U13736 (N_13736,N_10739,N_11199);
or U13737 (N_13737,N_11751,N_12319);
nor U13738 (N_13738,N_10623,N_11468);
nand U13739 (N_13739,N_10396,N_10185);
xor U13740 (N_13740,N_11441,N_10474);
and U13741 (N_13741,N_10024,N_10934);
nand U13742 (N_13742,N_10403,N_10333);
xnor U13743 (N_13743,N_10692,N_11964);
nand U13744 (N_13744,N_10076,N_11142);
and U13745 (N_13745,N_10010,N_11699);
or U13746 (N_13746,N_10646,N_10177);
nand U13747 (N_13747,N_12427,N_10674);
and U13748 (N_13748,N_11555,N_10609);
nand U13749 (N_13749,N_11440,N_10804);
xor U13750 (N_13750,N_11054,N_11921);
or U13751 (N_13751,N_11524,N_11451);
nor U13752 (N_13752,N_11719,N_12326);
nand U13753 (N_13753,N_11846,N_10539);
nor U13754 (N_13754,N_11884,N_10870);
and U13755 (N_13755,N_11030,N_10376);
nor U13756 (N_13756,N_11687,N_10178);
xnor U13757 (N_13757,N_11144,N_12161);
xnor U13758 (N_13758,N_11247,N_10193);
xnor U13759 (N_13759,N_11754,N_10545);
nor U13760 (N_13760,N_11430,N_12107);
nand U13761 (N_13761,N_11498,N_12107);
or U13762 (N_13762,N_10394,N_11579);
nor U13763 (N_13763,N_11641,N_10985);
xnor U13764 (N_13764,N_10381,N_11310);
nand U13765 (N_13765,N_10041,N_12049);
xor U13766 (N_13766,N_11947,N_12244);
and U13767 (N_13767,N_10996,N_10079);
xor U13768 (N_13768,N_10944,N_12128);
and U13769 (N_13769,N_10271,N_12468);
or U13770 (N_13770,N_10260,N_12472);
xnor U13771 (N_13771,N_10345,N_12300);
nor U13772 (N_13772,N_10262,N_10104);
and U13773 (N_13773,N_11481,N_10285);
nand U13774 (N_13774,N_12088,N_10598);
xnor U13775 (N_13775,N_10772,N_10428);
nor U13776 (N_13776,N_11081,N_12298);
xor U13777 (N_13777,N_11919,N_12161);
or U13778 (N_13778,N_11542,N_11881);
or U13779 (N_13779,N_10289,N_10371);
xor U13780 (N_13780,N_11984,N_11734);
and U13781 (N_13781,N_10493,N_10231);
nor U13782 (N_13782,N_12293,N_10375);
nand U13783 (N_13783,N_10954,N_11741);
or U13784 (N_13784,N_11618,N_11127);
and U13785 (N_13785,N_11778,N_10621);
xor U13786 (N_13786,N_10180,N_10527);
xnor U13787 (N_13787,N_10639,N_10155);
nand U13788 (N_13788,N_11912,N_10262);
nand U13789 (N_13789,N_11362,N_11812);
nand U13790 (N_13790,N_10858,N_11340);
nand U13791 (N_13791,N_12439,N_11680);
nand U13792 (N_13792,N_10359,N_12128);
xnor U13793 (N_13793,N_11414,N_10543);
and U13794 (N_13794,N_11176,N_10140);
nor U13795 (N_13795,N_11022,N_10359);
or U13796 (N_13796,N_10303,N_11784);
xnor U13797 (N_13797,N_10725,N_11604);
xnor U13798 (N_13798,N_12419,N_10864);
xor U13799 (N_13799,N_10276,N_10312);
or U13800 (N_13800,N_12311,N_11419);
and U13801 (N_13801,N_10532,N_12359);
nor U13802 (N_13802,N_11748,N_11857);
nand U13803 (N_13803,N_12253,N_11363);
and U13804 (N_13804,N_12440,N_10948);
nor U13805 (N_13805,N_12451,N_10796);
or U13806 (N_13806,N_11812,N_10169);
nand U13807 (N_13807,N_11635,N_12039);
xor U13808 (N_13808,N_12171,N_11419);
nand U13809 (N_13809,N_11105,N_10480);
nor U13810 (N_13810,N_11446,N_11783);
nand U13811 (N_13811,N_10650,N_10947);
nand U13812 (N_13812,N_10062,N_11317);
xor U13813 (N_13813,N_11479,N_11187);
and U13814 (N_13814,N_10456,N_10900);
nand U13815 (N_13815,N_11659,N_11076);
nand U13816 (N_13816,N_11639,N_10036);
xor U13817 (N_13817,N_12096,N_11066);
xnor U13818 (N_13818,N_11777,N_11583);
nor U13819 (N_13819,N_10137,N_11676);
nand U13820 (N_13820,N_11124,N_12370);
nor U13821 (N_13821,N_10123,N_11980);
or U13822 (N_13822,N_12123,N_12073);
nor U13823 (N_13823,N_11702,N_11194);
or U13824 (N_13824,N_12025,N_12213);
and U13825 (N_13825,N_12212,N_11021);
or U13826 (N_13826,N_11371,N_11617);
nor U13827 (N_13827,N_11721,N_10969);
and U13828 (N_13828,N_11719,N_11088);
xor U13829 (N_13829,N_11353,N_10702);
nor U13830 (N_13830,N_11084,N_12486);
and U13831 (N_13831,N_11892,N_11153);
or U13832 (N_13832,N_11410,N_10401);
and U13833 (N_13833,N_11990,N_10813);
nand U13834 (N_13834,N_11692,N_10663);
or U13835 (N_13835,N_11551,N_11363);
nor U13836 (N_13836,N_11616,N_10278);
or U13837 (N_13837,N_10551,N_10685);
nor U13838 (N_13838,N_12191,N_10022);
nor U13839 (N_13839,N_10408,N_12061);
nor U13840 (N_13840,N_12224,N_10074);
xnor U13841 (N_13841,N_11473,N_11702);
or U13842 (N_13842,N_10891,N_11707);
or U13843 (N_13843,N_11604,N_10610);
nor U13844 (N_13844,N_11665,N_10905);
and U13845 (N_13845,N_10148,N_10300);
and U13846 (N_13846,N_11506,N_10536);
or U13847 (N_13847,N_10209,N_11629);
and U13848 (N_13848,N_10927,N_11207);
and U13849 (N_13849,N_10780,N_11474);
xnor U13850 (N_13850,N_11244,N_12368);
nor U13851 (N_13851,N_10062,N_11859);
and U13852 (N_13852,N_10560,N_10592);
and U13853 (N_13853,N_11685,N_10026);
nand U13854 (N_13854,N_10270,N_11633);
nand U13855 (N_13855,N_11308,N_11744);
xor U13856 (N_13856,N_11298,N_10010);
nand U13857 (N_13857,N_11834,N_12034);
and U13858 (N_13858,N_10896,N_10681);
nand U13859 (N_13859,N_11696,N_11318);
xor U13860 (N_13860,N_10462,N_12161);
nand U13861 (N_13861,N_11332,N_12026);
and U13862 (N_13862,N_11491,N_12330);
xnor U13863 (N_13863,N_11932,N_10908);
or U13864 (N_13864,N_11990,N_11726);
or U13865 (N_13865,N_11171,N_11874);
nand U13866 (N_13866,N_11025,N_10930);
xor U13867 (N_13867,N_10045,N_10677);
nor U13868 (N_13868,N_12058,N_11611);
nand U13869 (N_13869,N_10384,N_10778);
xor U13870 (N_13870,N_11656,N_11282);
and U13871 (N_13871,N_10224,N_11884);
nand U13872 (N_13872,N_11771,N_11969);
nor U13873 (N_13873,N_11476,N_10363);
or U13874 (N_13874,N_10966,N_10664);
nand U13875 (N_13875,N_11281,N_12100);
nor U13876 (N_13876,N_10961,N_10970);
xnor U13877 (N_13877,N_11067,N_11080);
or U13878 (N_13878,N_10869,N_12096);
xnor U13879 (N_13879,N_10836,N_11732);
xnor U13880 (N_13880,N_11036,N_11935);
xnor U13881 (N_13881,N_10986,N_11848);
or U13882 (N_13882,N_11671,N_11534);
xnor U13883 (N_13883,N_11688,N_10214);
nor U13884 (N_13884,N_11419,N_10980);
nand U13885 (N_13885,N_10255,N_10115);
or U13886 (N_13886,N_12190,N_11802);
and U13887 (N_13887,N_11621,N_11080);
and U13888 (N_13888,N_12393,N_10438);
or U13889 (N_13889,N_12145,N_10322);
or U13890 (N_13890,N_12140,N_11776);
or U13891 (N_13891,N_10325,N_10631);
nand U13892 (N_13892,N_11307,N_12248);
and U13893 (N_13893,N_10266,N_10666);
xor U13894 (N_13894,N_10934,N_11666);
or U13895 (N_13895,N_12131,N_10722);
nor U13896 (N_13896,N_10832,N_10287);
xnor U13897 (N_13897,N_11652,N_10933);
and U13898 (N_13898,N_11541,N_10687);
xnor U13899 (N_13899,N_12445,N_11936);
or U13900 (N_13900,N_10468,N_12450);
nor U13901 (N_13901,N_10521,N_10691);
or U13902 (N_13902,N_12070,N_10063);
nor U13903 (N_13903,N_11041,N_12336);
and U13904 (N_13904,N_11827,N_12120);
nor U13905 (N_13905,N_11005,N_10615);
nand U13906 (N_13906,N_10411,N_11401);
xor U13907 (N_13907,N_10516,N_10527);
nor U13908 (N_13908,N_10082,N_10259);
and U13909 (N_13909,N_12042,N_11075);
nand U13910 (N_13910,N_11480,N_11862);
nor U13911 (N_13911,N_11818,N_12324);
and U13912 (N_13912,N_11469,N_10839);
nor U13913 (N_13913,N_10528,N_10057);
or U13914 (N_13914,N_11293,N_10492);
and U13915 (N_13915,N_11792,N_10306);
nand U13916 (N_13916,N_11776,N_10027);
nor U13917 (N_13917,N_11608,N_11109);
and U13918 (N_13918,N_10200,N_11295);
and U13919 (N_13919,N_10326,N_10006);
nor U13920 (N_13920,N_10483,N_11946);
nor U13921 (N_13921,N_12195,N_10773);
nand U13922 (N_13922,N_10019,N_11783);
nor U13923 (N_13923,N_12392,N_11524);
and U13924 (N_13924,N_10385,N_11242);
or U13925 (N_13925,N_11196,N_11980);
xnor U13926 (N_13926,N_11260,N_11022);
xnor U13927 (N_13927,N_10014,N_10049);
xor U13928 (N_13928,N_11348,N_11221);
nor U13929 (N_13929,N_11764,N_10079);
or U13930 (N_13930,N_10610,N_10353);
or U13931 (N_13931,N_10906,N_11041);
and U13932 (N_13932,N_12338,N_11026);
and U13933 (N_13933,N_10387,N_11898);
nand U13934 (N_13934,N_12323,N_10477);
nor U13935 (N_13935,N_11415,N_10415);
xor U13936 (N_13936,N_11665,N_10099);
nand U13937 (N_13937,N_11821,N_12492);
and U13938 (N_13938,N_10425,N_10092);
or U13939 (N_13939,N_10036,N_11518);
xnor U13940 (N_13940,N_11815,N_11126);
and U13941 (N_13941,N_10895,N_11944);
or U13942 (N_13942,N_10136,N_10260);
or U13943 (N_13943,N_10943,N_10131);
nand U13944 (N_13944,N_10841,N_10545);
xnor U13945 (N_13945,N_11581,N_11201);
or U13946 (N_13946,N_10853,N_11611);
nand U13947 (N_13947,N_10005,N_11896);
xor U13948 (N_13948,N_10632,N_11437);
and U13949 (N_13949,N_10669,N_12170);
nor U13950 (N_13950,N_11459,N_10256);
xnor U13951 (N_13951,N_11379,N_10074);
nand U13952 (N_13952,N_10462,N_11084);
xor U13953 (N_13953,N_10109,N_10996);
or U13954 (N_13954,N_12017,N_10135);
nand U13955 (N_13955,N_12395,N_11707);
nor U13956 (N_13956,N_12413,N_10619);
nor U13957 (N_13957,N_12073,N_11374);
and U13958 (N_13958,N_11225,N_12092);
xor U13959 (N_13959,N_10575,N_10862);
or U13960 (N_13960,N_11724,N_11210);
xnor U13961 (N_13961,N_10973,N_11689);
or U13962 (N_13962,N_11713,N_12120);
xor U13963 (N_13963,N_10123,N_12213);
nand U13964 (N_13964,N_11249,N_11071);
and U13965 (N_13965,N_11179,N_11485);
nand U13966 (N_13966,N_12348,N_10506);
nor U13967 (N_13967,N_11130,N_12210);
or U13968 (N_13968,N_11158,N_11146);
or U13969 (N_13969,N_12086,N_12161);
xnor U13970 (N_13970,N_10149,N_11889);
nor U13971 (N_13971,N_12203,N_10130);
and U13972 (N_13972,N_11175,N_11152);
xor U13973 (N_13973,N_11773,N_12124);
and U13974 (N_13974,N_11846,N_11493);
nand U13975 (N_13975,N_11733,N_11439);
or U13976 (N_13976,N_11909,N_12138);
xor U13977 (N_13977,N_11633,N_10202);
nor U13978 (N_13978,N_10757,N_11478);
xor U13979 (N_13979,N_10263,N_11951);
nand U13980 (N_13980,N_10788,N_10634);
nand U13981 (N_13981,N_11137,N_11961);
nand U13982 (N_13982,N_11733,N_12151);
nand U13983 (N_13983,N_12228,N_12411);
and U13984 (N_13984,N_11735,N_10330);
or U13985 (N_13985,N_11307,N_11900);
xnor U13986 (N_13986,N_10062,N_10091);
xor U13987 (N_13987,N_11820,N_10825);
xor U13988 (N_13988,N_12434,N_12253);
nand U13989 (N_13989,N_11562,N_11812);
xor U13990 (N_13990,N_11624,N_12490);
xnor U13991 (N_13991,N_11703,N_10761);
nand U13992 (N_13992,N_11620,N_11978);
xor U13993 (N_13993,N_11926,N_10132);
or U13994 (N_13994,N_11140,N_10679);
and U13995 (N_13995,N_10084,N_10005);
xor U13996 (N_13996,N_11081,N_11414);
or U13997 (N_13997,N_11736,N_11301);
or U13998 (N_13998,N_12434,N_10388);
and U13999 (N_13999,N_10132,N_11381);
or U14000 (N_14000,N_10179,N_11597);
nand U14001 (N_14001,N_12264,N_12175);
and U14002 (N_14002,N_10151,N_11317);
xor U14003 (N_14003,N_11722,N_11920);
nor U14004 (N_14004,N_11648,N_10485);
xor U14005 (N_14005,N_11177,N_11763);
xor U14006 (N_14006,N_11668,N_10611);
and U14007 (N_14007,N_11499,N_11121);
or U14008 (N_14008,N_11037,N_12202);
nand U14009 (N_14009,N_10385,N_11800);
and U14010 (N_14010,N_12474,N_11732);
or U14011 (N_14011,N_10839,N_11583);
and U14012 (N_14012,N_10948,N_10763);
xor U14013 (N_14013,N_11362,N_11752);
nor U14014 (N_14014,N_11931,N_11243);
or U14015 (N_14015,N_10741,N_12328);
xor U14016 (N_14016,N_11931,N_10462);
nand U14017 (N_14017,N_11510,N_12201);
and U14018 (N_14018,N_10002,N_11442);
and U14019 (N_14019,N_11222,N_12249);
nand U14020 (N_14020,N_11140,N_11917);
nor U14021 (N_14021,N_10965,N_11056);
and U14022 (N_14022,N_10558,N_10268);
or U14023 (N_14023,N_11928,N_12320);
xor U14024 (N_14024,N_10050,N_11022);
and U14025 (N_14025,N_11093,N_11924);
nand U14026 (N_14026,N_10998,N_11733);
nand U14027 (N_14027,N_10278,N_11435);
xnor U14028 (N_14028,N_10472,N_12222);
nand U14029 (N_14029,N_11575,N_12121);
xor U14030 (N_14030,N_10207,N_11190);
or U14031 (N_14031,N_10834,N_11951);
nand U14032 (N_14032,N_10329,N_10402);
or U14033 (N_14033,N_11485,N_11631);
nor U14034 (N_14034,N_10629,N_10819);
xnor U14035 (N_14035,N_10112,N_10605);
or U14036 (N_14036,N_12020,N_11594);
nand U14037 (N_14037,N_10671,N_11234);
nor U14038 (N_14038,N_10162,N_10489);
and U14039 (N_14039,N_10860,N_10719);
xor U14040 (N_14040,N_12425,N_12020);
and U14041 (N_14041,N_10384,N_10078);
nand U14042 (N_14042,N_11935,N_10816);
xor U14043 (N_14043,N_11950,N_10038);
and U14044 (N_14044,N_11166,N_11003);
or U14045 (N_14045,N_12240,N_11617);
or U14046 (N_14046,N_11810,N_10863);
nand U14047 (N_14047,N_11279,N_10984);
nand U14048 (N_14048,N_11298,N_10448);
nand U14049 (N_14049,N_10791,N_11269);
and U14050 (N_14050,N_10909,N_10932);
xnor U14051 (N_14051,N_11329,N_10978);
nor U14052 (N_14052,N_11082,N_11972);
nand U14053 (N_14053,N_10062,N_12075);
xor U14054 (N_14054,N_11136,N_10926);
xnor U14055 (N_14055,N_12421,N_11981);
nor U14056 (N_14056,N_10726,N_11696);
nand U14057 (N_14057,N_10524,N_11251);
and U14058 (N_14058,N_11914,N_10639);
xor U14059 (N_14059,N_11599,N_10378);
nor U14060 (N_14060,N_12080,N_11443);
xnor U14061 (N_14061,N_10993,N_12485);
or U14062 (N_14062,N_10748,N_10293);
xor U14063 (N_14063,N_11148,N_10176);
xor U14064 (N_14064,N_12267,N_10940);
or U14065 (N_14065,N_12433,N_11044);
or U14066 (N_14066,N_11485,N_11194);
nor U14067 (N_14067,N_11091,N_10660);
xnor U14068 (N_14068,N_11838,N_12190);
and U14069 (N_14069,N_10975,N_11832);
or U14070 (N_14070,N_10674,N_10715);
or U14071 (N_14071,N_11858,N_11136);
or U14072 (N_14072,N_12326,N_10341);
nor U14073 (N_14073,N_11711,N_11540);
xnor U14074 (N_14074,N_11089,N_11110);
xnor U14075 (N_14075,N_11507,N_10728);
and U14076 (N_14076,N_11384,N_12443);
and U14077 (N_14077,N_10027,N_11764);
or U14078 (N_14078,N_11390,N_12002);
nand U14079 (N_14079,N_10061,N_10662);
xor U14080 (N_14080,N_10638,N_10363);
and U14081 (N_14081,N_11071,N_12498);
and U14082 (N_14082,N_12428,N_10533);
or U14083 (N_14083,N_11441,N_10133);
nor U14084 (N_14084,N_11589,N_10002);
nor U14085 (N_14085,N_12315,N_11177);
and U14086 (N_14086,N_12486,N_11352);
and U14087 (N_14087,N_10739,N_12198);
xnor U14088 (N_14088,N_11774,N_12370);
nand U14089 (N_14089,N_10020,N_11074);
nand U14090 (N_14090,N_11321,N_11375);
or U14091 (N_14091,N_11481,N_12478);
nor U14092 (N_14092,N_10359,N_10453);
and U14093 (N_14093,N_10038,N_11897);
nor U14094 (N_14094,N_10460,N_11362);
nor U14095 (N_14095,N_10847,N_10177);
nor U14096 (N_14096,N_10144,N_11610);
or U14097 (N_14097,N_11229,N_10823);
or U14098 (N_14098,N_10498,N_10715);
or U14099 (N_14099,N_11082,N_10690);
nand U14100 (N_14100,N_10827,N_11699);
and U14101 (N_14101,N_11790,N_10836);
nand U14102 (N_14102,N_11582,N_11167);
nand U14103 (N_14103,N_11973,N_10576);
xor U14104 (N_14104,N_11528,N_11749);
nor U14105 (N_14105,N_10914,N_10253);
and U14106 (N_14106,N_10729,N_10343);
or U14107 (N_14107,N_11403,N_12188);
xnor U14108 (N_14108,N_10865,N_11263);
or U14109 (N_14109,N_12483,N_11482);
or U14110 (N_14110,N_11566,N_12013);
xor U14111 (N_14111,N_12032,N_10825);
nand U14112 (N_14112,N_10958,N_11527);
xor U14113 (N_14113,N_11909,N_11232);
or U14114 (N_14114,N_12310,N_12494);
or U14115 (N_14115,N_12382,N_10092);
nor U14116 (N_14116,N_11332,N_10077);
xnor U14117 (N_14117,N_10269,N_12099);
nand U14118 (N_14118,N_11542,N_11648);
or U14119 (N_14119,N_11107,N_12167);
nand U14120 (N_14120,N_10434,N_11899);
and U14121 (N_14121,N_11323,N_10528);
or U14122 (N_14122,N_11363,N_10582);
xor U14123 (N_14123,N_12432,N_11678);
nand U14124 (N_14124,N_12293,N_10234);
xnor U14125 (N_14125,N_12466,N_10203);
and U14126 (N_14126,N_10458,N_12185);
and U14127 (N_14127,N_12417,N_12446);
or U14128 (N_14128,N_10296,N_11118);
or U14129 (N_14129,N_12078,N_11759);
nand U14130 (N_14130,N_10007,N_10296);
nor U14131 (N_14131,N_11271,N_10955);
xor U14132 (N_14132,N_11704,N_12433);
and U14133 (N_14133,N_10460,N_12200);
or U14134 (N_14134,N_10049,N_11548);
xor U14135 (N_14135,N_12298,N_10381);
nand U14136 (N_14136,N_10136,N_12340);
nor U14137 (N_14137,N_10222,N_10399);
or U14138 (N_14138,N_11624,N_11189);
xnor U14139 (N_14139,N_10598,N_11247);
nand U14140 (N_14140,N_11293,N_11192);
and U14141 (N_14141,N_10321,N_10815);
xor U14142 (N_14142,N_12306,N_10298);
nor U14143 (N_14143,N_11776,N_11019);
xnor U14144 (N_14144,N_11905,N_10353);
xnor U14145 (N_14145,N_10564,N_10151);
nor U14146 (N_14146,N_11874,N_10081);
and U14147 (N_14147,N_11675,N_12159);
and U14148 (N_14148,N_12296,N_10322);
or U14149 (N_14149,N_11592,N_12492);
nor U14150 (N_14150,N_11542,N_10450);
nand U14151 (N_14151,N_10034,N_10808);
or U14152 (N_14152,N_10473,N_12085);
xor U14153 (N_14153,N_12125,N_10769);
and U14154 (N_14154,N_11192,N_12188);
and U14155 (N_14155,N_11573,N_10207);
nand U14156 (N_14156,N_10553,N_12008);
xor U14157 (N_14157,N_10076,N_10317);
or U14158 (N_14158,N_11271,N_12437);
nor U14159 (N_14159,N_12227,N_12329);
nand U14160 (N_14160,N_11372,N_10459);
or U14161 (N_14161,N_11860,N_11609);
nand U14162 (N_14162,N_11057,N_11842);
nor U14163 (N_14163,N_12152,N_12218);
nor U14164 (N_14164,N_12312,N_10932);
or U14165 (N_14165,N_11567,N_12055);
nor U14166 (N_14166,N_12100,N_12006);
or U14167 (N_14167,N_11078,N_10728);
and U14168 (N_14168,N_11499,N_11685);
and U14169 (N_14169,N_11646,N_12233);
or U14170 (N_14170,N_10332,N_11914);
nand U14171 (N_14171,N_10109,N_12389);
or U14172 (N_14172,N_12195,N_10240);
or U14173 (N_14173,N_11808,N_11216);
and U14174 (N_14174,N_10901,N_10113);
or U14175 (N_14175,N_12126,N_11544);
nor U14176 (N_14176,N_11195,N_11775);
nor U14177 (N_14177,N_11739,N_11042);
nor U14178 (N_14178,N_10891,N_11230);
and U14179 (N_14179,N_11457,N_11637);
and U14180 (N_14180,N_10772,N_11805);
nor U14181 (N_14181,N_11567,N_10730);
xor U14182 (N_14182,N_11908,N_11175);
nand U14183 (N_14183,N_12254,N_12285);
nand U14184 (N_14184,N_11656,N_10818);
or U14185 (N_14185,N_12459,N_11006);
and U14186 (N_14186,N_12099,N_10400);
and U14187 (N_14187,N_12054,N_10976);
nor U14188 (N_14188,N_10896,N_11389);
or U14189 (N_14189,N_10933,N_10353);
or U14190 (N_14190,N_10031,N_11324);
nand U14191 (N_14191,N_10647,N_12085);
xor U14192 (N_14192,N_10929,N_11059);
nand U14193 (N_14193,N_10806,N_11781);
or U14194 (N_14194,N_10460,N_11308);
and U14195 (N_14195,N_10212,N_10353);
nand U14196 (N_14196,N_10477,N_11078);
and U14197 (N_14197,N_10832,N_12324);
and U14198 (N_14198,N_10664,N_10289);
nand U14199 (N_14199,N_11051,N_11075);
and U14200 (N_14200,N_11085,N_10635);
and U14201 (N_14201,N_10211,N_10875);
and U14202 (N_14202,N_11383,N_11859);
xor U14203 (N_14203,N_10466,N_10915);
xnor U14204 (N_14204,N_11953,N_11165);
and U14205 (N_14205,N_10594,N_11902);
xor U14206 (N_14206,N_11715,N_12344);
xnor U14207 (N_14207,N_10792,N_11786);
and U14208 (N_14208,N_11111,N_10217);
nor U14209 (N_14209,N_10186,N_11137);
or U14210 (N_14210,N_11493,N_11717);
xnor U14211 (N_14211,N_11844,N_10077);
nand U14212 (N_14212,N_11509,N_10820);
or U14213 (N_14213,N_10517,N_10185);
and U14214 (N_14214,N_11554,N_10043);
xnor U14215 (N_14215,N_11569,N_10085);
or U14216 (N_14216,N_11905,N_11712);
xor U14217 (N_14217,N_10296,N_11242);
or U14218 (N_14218,N_10595,N_10713);
xnor U14219 (N_14219,N_10103,N_11507);
nor U14220 (N_14220,N_12356,N_10032);
and U14221 (N_14221,N_11721,N_11020);
nor U14222 (N_14222,N_11526,N_10432);
nand U14223 (N_14223,N_12455,N_11773);
nor U14224 (N_14224,N_11596,N_10922);
nand U14225 (N_14225,N_11856,N_11757);
and U14226 (N_14226,N_11654,N_11271);
xnor U14227 (N_14227,N_11583,N_10804);
nor U14228 (N_14228,N_11659,N_10904);
and U14229 (N_14229,N_12052,N_11680);
xnor U14230 (N_14230,N_10664,N_11396);
or U14231 (N_14231,N_11053,N_10122);
and U14232 (N_14232,N_10615,N_10447);
and U14233 (N_14233,N_10534,N_10493);
nor U14234 (N_14234,N_11055,N_10120);
and U14235 (N_14235,N_12252,N_10479);
and U14236 (N_14236,N_11634,N_10914);
nor U14237 (N_14237,N_11146,N_10476);
nor U14238 (N_14238,N_11145,N_12199);
nor U14239 (N_14239,N_12107,N_12430);
and U14240 (N_14240,N_10434,N_12163);
nand U14241 (N_14241,N_11799,N_10138);
or U14242 (N_14242,N_12390,N_10992);
or U14243 (N_14243,N_10384,N_10245);
nor U14244 (N_14244,N_10291,N_10116);
nor U14245 (N_14245,N_11657,N_12111);
nand U14246 (N_14246,N_11323,N_12334);
nand U14247 (N_14247,N_11163,N_11830);
nand U14248 (N_14248,N_10095,N_11544);
and U14249 (N_14249,N_12244,N_10840);
and U14250 (N_14250,N_11469,N_12083);
xnor U14251 (N_14251,N_11171,N_11099);
nand U14252 (N_14252,N_10329,N_12448);
or U14253 (N_14253,N_10810,N_10520);
xnor U14254 (N_14254,N_11361,N_11199);
nor U14255 (N_14255,N_12185,N_12129);
nor U14256 (N_14256,N_11504,N_12220);
and U14257 (N_14257,N_10753,N_11101);
and U14258 (N_14258,N_11557,N_10462);
nor U14259 (N_14259,N_10753,N_11703);
or U14260 (N_14260,N_12272,N_11176);
or U14261 (N_14261,N_11234,N_10973);
xnor U14262 (N_14262,N_10616,N_12202);
nor U14263 (N_14263,N_11790,N_11136);
nor U14264 (N_14264,N_11850,N_11549);
nor U14265 (N_14265,N_12280,N_11425);
nor U14266 (N_14266,N_12070,N_11729);
xor U14267 (N_14267,N_10760,N_11744);
or U14268 (N_14268,N_11471,N_10865);
or U14269 (N_14269,N_11498,N_11251);
nor U14270 (N_14270,N_11692,N_11830);
or U14271 (N_14271,N_10398,N_11088);
nand U14272 (N_14272,N_10728,N_10447);
nand U14273 (N_14273,N_10489,N_10949);
nand U14274 (N_14274,N_10855,N_11684);
xnor U14275 (N_14275,N_11652,N_10545);
and U14276 (N_14276,N_12372,N_10160);
and U14277 (N_14277,N_10222,N_11870);
or U14278 (N_14278,N_12169,N_11663);
xnor U14279 (N_14279,N_11152,N_10483);
and U14280 (N_14280,N_11849,N_10316);
and U14281 (N_14281,N_12037,N_11306);
nand U14282 (N_14282,N_12251,N_11211);
xor U14283 (N_14283,N_12275,N_11189);
nor U14284 (N_14284,N_10710,N_10922);
and U14285 (N_14285,N_10633,N_10866);
and U14286 (N_14286,N_10706,N_12159);
and U14287 (N_14287,N_11894,N_12226);
or U14288 (N_14288,N_11336,N_10024);
nand U14289 (N_14289,N_10661,N_10897);
nand U14290 (N_14290,N_10657,N_11932);
and U14291 (N_14291,N_10968,N_11908);
or U14292 (N_14292,N_12041,N_10561);
nand U14293 (N_14293,N_12373,N_10474);
and U14294 (N_14294,N_10855,N_10399);
nand U14295 (N_14295,N_11773,N_11804);
xor U14296 (N_14296,N_10496,N_12023);
nand U14297 (N_14297,N_10561,N_11691);
nor U14298 (N_14298,N_12324,N_11553);
and U14299 (N_14299,N_10731,N_10525);
nand U14300 (N_14300,N_11355,N_10187);
xor U14301 (N_14301,N_11097,N_12214);
or U14302 (N_14302,N_10931,N_11796);
nor U14303 (N_14303,N_10185,N_11663);
nand U14304 (N_14304,N_11132,N_10850);
nand U14305 (N_14305,N_12082,N_12351);
nand U14306 (N_14306,N_11335,N_10013);
xnor U14307 (N_14307,N_12230,N_10340);
or U14308 (N_14308,N_12109,N_12273);
xor U14309 (N_14309,N_10798,N_10147);
or U14310 (N_14310,N_10557,N_11163);
or U14311 (N_14311,N_10993,N_10480);
or U14312 (N_14312,N_11294,N_10436);
or U14313 (N_14313,N_11304,N_11289);
and U14314 (N_14314,N_10581,N_11238);
nand U14315 (N_14315,N_10304,N_12055);
nand U14316 (N_14316,N_10585,N_11233);
and U14317 (N_14317,N_10948,N_10041);
and U14318 (N_14318,N_12202,N_10569);
and U14319 (N_14319,N_10822,N_10381);
xnor U14320 (N_14320,N_12247,N_10393);
and U14321 (N_14321,N_10394,N_10756);
nand U14322 (N_14322,N_12304,N_10075);
or U14323 (N_14323,N_10751,N_12387);
or U14324 (N_14324,N_11879,N_10344);
or U14325 (N_14325,N_10271,N_10833);
nand U14326 (N_14326,N_10201,N_10539);
xnor U14327 (N_14327,N_11774,N_10862);
nor U14328 (N_14328,N_11052,N_12015);
or U14329 (N_14329,N_12072,N_12366);
and U14330 (N_14330,N_10180,N_12147);
or U14331 (N_14331,N_10450,N_10990);
and U14332 (N_14332,N_10912,N_10713);
and U14333 (N_14333,N_11071,N_12354);
nor U14334 (N_14334,N_12323,N_10933);
nand U14335 (N_14335,N_10046,N_12439);
and U14336 (N_14336,N_10555,N_11398);
or U14337 (N_14337,N_11632,N_10686);
nor U14338 (N_14338,N_10804,N_10667);
and U14339 (N_14339,N_11797,N_10182);
nor U14340 (N_14340,N_11386,N_10554);
and U14341 (N_14341,N_12230,N_11746);
nor U14342 (N_14342,N_10444,N_10416);
xnor U14343 (N_14343,N_10600,N_11543);
and U14344 (N_14344,N_10362,N_10263);
xor U14345 (N_14345,N_11420,N_11924);
and U14346 (N_14346,N_12191,N_12096);
nand U14347 (N_14347,N_10695,N_11208);
and U14348 (N_14348,N_10969,N_11468);
and U14349 (N_14349,N_11628,N_11604);
nand U14350 (N_14350,N_11718,N_10439);
nand U14351 (N_14351,N_11176,N_10594);
or U14352 (N_14352,N_10433,N_11166);
or U14353 (N_14353,N_10416,N_11874);
or U14354 (N_14354,N_11223,N_11109);
nor U14355 (N_14355,N_10268,N_11662);
nand U14356 (N_14356,N_11447,N_10178);
nand U14357 (N_14357,N_11310,N_10498);
nand U14358 (N_14358,N_10769,N_11022);
nand U14359 (N_14359,N_10193,N_11640);
nand U14360 (N_14360,N_11574,N_11359);
nor U14361 (N_14361,N_10353,N_11060);
nor U14362 (N_14362,N_12245,N_11145);
and U14363 (N_14363,N_11856,N_12252);
or U14364 (N_14364,N_11059,N_10588);
and U14365 (N_14365,N_10658,N_11164);
nor U14366 (N_14366,N_10807,N_11473);
and U14367 (N_14367,N_10581,N_11075);
and U14368 (N_14368,N_10444,N_10114);
and U14369 (N_14369,N_10961,N_12300);
or U14370 (N_14370,N_12083,N_12001);
nand U14371 (N_14371,N_12339,N_12050);
and U14372 (N_14372,N_11436,N_10600);
nor U14373 (N_14373,N_10405,N_11396);
nor U14374 (N_14374,N_11379,N_12237);
and U14375 (N_14375,N_10727,N_11087);
nor U14376 (N_14376,N_12217,N_12085);
nand U14377 (N_14377,N_11975,N_11618);
nand U14378 (N_14378,N_12089,N_10665);
nor U14379 (N_14379,N_10920,N_10808);
or U14380 (N_14380,N_11757,N_11748);
xor U14381 (N_14381,N_11827,N_10649);
nor U14382 (N_14382,N_12038,N_12477);
or U14383 (N_14383,N_10923,N_11070);
and U14384 (N_14384,N_10136,N_10625);
and U14385 (N_14385,N_10960,N_11664);
nand U14386 (N_14386,N_12277,N_10497);
nand U14387 (N_14387,N_10943,N_11650);
and U14388 (N_14388,N_10236,N_10947);
nor U14389 (N_14389,N_12427,N_10741);
nand U14390 (N_14390,N_12392,N_11357);
nor U14391 (N_14391,N_12019,N_10856);
or U14392 (N_14392,N_11480,N_11295);
nor U14393 (N_14393,N_10403,N_12256);
xnor U14394 (N_14394,N_11718,N_10155);
or U14395 (N_14395,N_10549,N_11601);
or U14396 (N_14396,N_11294,N_12234);
and U14397 (N_14397,N_10869,N_10321);
nand U14398 (N_14398,N_11248,N_12206);
and U14399 (N_14399,N_12092,N_11005);
nand U14400 (N_14400,N_10128,N_10658);
nand U14401 (N_14401,N_11584,N_11796);
nor U14402 (N_14402,N_10166,N_11126);
and U14403 (N_14403,N_12391,N_11644);
nor U14404 (N_14404,N_12320,N_10141);
xor U14405 (N_14405,N_10422,N_10590);
nor U14406 (N_14406,N_11783,N_12103);
nor U14407 (N_14407,N_11309,N_11546);
nor U14408 (N_14408,N_11422,N_12414);
or U14409 (N_14409,N_12102,N_11382);
nand U14410 (N_14410,N_10592,N_10300);
nor U14411 (N_14411,N_12054,N_10624);
xor U14412 (N_14412,N_10498,N_11348);
nor U14413 (N_14413,N_12328,N_10445);
nand U14414 (N_14414,N_11124,N_10349);
xor U14415 (N_14415,N_10996,N_12263);
xor U14416 (N_14416,N_10335,N_11012);
or U14417 (N_14417,N_10632,N_12315);
xnor U14418 (N_14418,N_10797,N_10251);
nor U14419 (N_14419,N_10093,N_11825);
nor U14420 (N_14420,N_11032,N_12114);
or U14421 (N_14421,N_10788,N_10503);
nor U14422 (N_14422,N_11646,N_11808);
xor U14423 (N_14423,N_11850,N_11431);
and U14424 (N_14424,N_10163,N_10863);
nand U14425 (N_14425,N_11574,N_12208);
nor U14426 (N_14426,N_11693,N_12461);
nor U14427 (N_14427,N_12360,N_10053);
nand U14428 (N_14428,N_11692,N_10201);
nand U14429 (N_14429,N_11291,N_10620);
nand U14430 (N_14430,N_11632,N_12495);
nor U14431 (N_14431,N_11313,N_10600);
and U14432 (N_14432,N_10958,N_11280);
and U14433 (N_14433,N_12283,N_11326);
xor U14434 (N_14434,N_10383,N_10985);
nor U14435 (N_14435,N_11670,N_12053);
nand U14436 (N_14436,N_12256,N_10665);
xor U14437 (N_14437,N_10890,N_10235);
nor U14438 (N_14438,N_11774,N_12473);
and U14439 (N_14439,N_10676,N_12020);
or U14440 (N_14440,N_10949,N_11054);
nor U14441 (N_14441,N_11162,N_10718);
xor U14442 (N_14442,N_10151,N_11202);
or U14443 (N_14443,N_10992,N_12140);
xnor U14444 (N_14444,N_10766,N_12006);
or U14445 (N_14445,N_12318,N_11342);
and U14446 (N_14446,N_11627,N_11369);
nand U14447 (N_14447,N_10021,N_10508);
or U14448 (N_14448,N_11585,N_12059);
nor U14449 (N_14449,N_11454,N_12157);
or U14450 (N_14450,N_12165,N_11294);
or U14451 (N_14451,N_10060,N_10414);
and U14452 (N_14452,N_10613,N_11685);
and U14453 (N_14453,N_11886,N_10307);
and U14454 (N_14454,N_11696,N_12064);
nand U14455 (N_14455,N_11900,N_11227);
nand U14456 (N_14456,N_12056,N_10371);
nor U14457 (N_14457,N_12336,N_10665);
nor U14458 (N_14458,N_11844,N_10674);
xnor U14459 (N_14459,N_10324,N_11407);
xnor U14460 (N_14460,N_10098,N_10419);
nor U14461 (N_14461,N_10476,N_11372);
xor U14462 (N_14462,N_10089,N_10383);
nand U14463 (N_14463,N_11008,N_11678);
xnor U14464 (N_14464,N_12130,N_10361);
nand U14465 (N_14465,N_11499,N_12026);
or U14466 (N_14466,N_11429,N_11841);
xor U14467 (N_14467,N_10753,N_10538);
or U14468 (N_14468,N_10396,N_10377);
and U14469 (N_14469,N_10694,N_10241);
or U14470 (N_14470,N_10347,N_10586);
or U14471 (N_14471,N_10495,N_11950);
nor U14472 (N_14472,N_12393,N_12250);
xor U14473 (N_14473,N_10941,N_11286);
nand U14474 (N_14474,N_11736,N_11037);
xor U14475 (N_14475,N_11951,N_10926);
nand U14476 (N_14476,N_10484,N_10440);
or U14477 (N_14477,N_10132,N_12001);
nor U14478 (N_14478,N_10693,N_10315);
nor U14479 (N_14479,N_10177,N_11526);
nand U14480 (N_14480,N_11345,N_11932);
or U14481 (N_14481,N_12060,N_11759);
nand U14482 (N_14482,N_10849,N_10086);
and U14483 (N_14483,N_11121,N_11777);
nand U14484 (N_14484,N_12172,N_11291);
nand U14485 (N_14485,N_11867,N_11768);
and U14486 (N_14486,N_10894,N_11521);
xor U14487 (N_14487,N_11845,N_12167);
xnor U14488 (N_14488,N_10133,N_11882);
nand U14489 (N_14489,N_10048,N_10696);
nor U14490 (N_14490,N_10674,N_12442);
or U14491 (N_14491,N_10741,N_10800);
nor U14492 (N_14492,N_10695,N_10744);
xor U14493 (N_14493,N_11025,N_11264);
xor U14494 (N_14494,N_11726,N_11168);
xnor U14495 (N_14495,N_12236,N_11936);
xor U14496 (N_14496,N_10567,N_12497);
xor U14497 (N_14497,N_12451,N_11847);
nand U14498 (N_14498,N_11586,N_11856);
nor U14499 (N_14499,N_10459,N_10195);
xnor U14500 (N_14500,N_10816,N_10072);
or U14501 (N_14501,N_11197,N_12076);
nor U14502 (N_14502,N_10192,N_11209);
nand U14503 (N_14503,N_10207,N_12322);
nor U14504 (N_14504,N_12132,N_11902);
xor U14505 (N_14505,N_12022,N_10732);
or U14506 (N_14506,N_12297,N_10569);
nand U14507 (N_14507,N_12437,N_11392);
or U14508 (N_14508,N_12003,N_11420);
or U14509 (N_14509,N_11205,N_10756);
xor U14510 (N_14510,N_11765,N_10618);
nor U14511 (N_14511,N_11834,N_12436);
nor U14512 (N_14512,N_10121,N_11437);
or U14513 (N_14513,N_10352,N_12264);
nor U14514 (N_14514,N_12128,N_10254);
or U14515 (N_14515,N_10728,N_10343);
nor U14516 (N_14516,N_10498,N_10806);
or U14517 (N_14517,N_12008,N_10424);
or U14518 (N_14518,N_10409,N_12223);
xor U14519 (N_14519,N_12039,N_10341);
nand U14520 (N_14520,N_10224,N_11557);
nor U14521 (N_14521,N_11449,N_11458);
nor U14522 (N_14522,N_10916,N_12214);
nor U14523 (N_14523,N_11483,N_10449);
or U14524 (N_14524,N_11212,N_12025);
nor U14525 (N_14525,N_11710,N_11488);
or U14526 (N_14526,N_10505,N_10426);
nand U14527 (N_14527,N_11085,N_10715);
xor U14528 (N_14528,N_10995,N_11407);
xor U14529 (N_14529,N_11518,N_11399);
xor U14530 (N_14530,N_11587,N_11630);
and U14531 (N_14531,N_12481,N_10612);
or U14532 (N_14532,N_12490,N_11943);
and U14533 (N_14533,N_11087,N_11136);
nand U14534 (N_14534,N_10161,N_10446);
or U14535 (N_14535,N_10467,N_11270);
xnor U14536 (N_14536,N_11604,N_11551);
nor U14537 (N_14537,N_10559,N_12146);
or U14538 (N_14538,N_10120,N_11135);
and U14539 (N_14539,N_11301,N_12233);
nor U14540 (N_14540,N_10523,N_10464);
and U14541 (N_14541,N_11991,N_10759);
or U14542 (N_14542,N_11101,N_11992);
nor U14543 (N_14543,N_10598,N_12335);
and U14544 (N_14544,N_11850,N_10454);
nor U14545 (N_14545,N_10822,N_10492);
and U14546 (N_14546,N_12117,N_10774);
and U14547 (N_14547,N_12264,N_11500);
or U14548 (N_14548,N_12232,N_11799);
nand U14549 (N_14549,N_11589,N_11134);
nor U14550 (N_14550,N_11662,N_10982);
xor U14551 (N_14551,N_12376,N_10372);
or U14552 (N_14552,N_10772,N_10994);
xor U14553 (N_14553,N_10739,N_10979);
nor U14554 (N_14554,N_11709,N_11876);
nand U14555 (N_14555,N_10813,N_10787);
nand U14556 (N_14556,N_10551,N_11337);
and U14557 (N_14557,N_12033,N_11957);
xor U14558 (N_14558,N_12417,N_12257);
nor U14559 (N_14559,N_10341,N_12490);
xnor U14560 (N_14560,N_10067,N_10129);
and U14561 (N_14561,N_11394,N_11059);
xnor U14562 (N_14562,N_11959,N_12490);
or U14563 (N_14563,N_12110,N_11193);
nand U14564 (N_14564,N_11012,N_11159);
nand U14565 (N_14565,N_11957,N_11634);
nand U14566 (N_14566,N_12085,N_11764);
nor U14567 (N_14567,N_10074,N_11860);
nand U14568 (N_14568,N_11301,N_12077);
nand U14569 (N_14569,N_10363,N_10136);
nor U14570 (N_14570,N_12083,N_11612);
xor U14571 (N_14571,N_10030,N_11873);
nor U14572 (N_14572,N_10041,N_10737);
nor U14573 (N_14573,N_12118,N_11512);
xor U14574 (N_14574,N_12202,N_11874);
nand U14575 (N_14575,N_11734,N_12122);
and U14576 (N_14576,N_10656,N_12202);
and U14577 (N_14577,N_11080,N_12222);
nand U14578 (N_14578,N_12430,N_11600);
and U14579 (N_14579,N_11752,N_11295);
and U14580 (N_14580,N_11920,N_10731);
or U14581 (N_14581,N_10334,N_11583);
xnor U14582 (N_14582,N_10273,N_12446);
nor U14583 (N_14583,N_11380,N_11729);
xor U14584 (N_14584,N_11397,N_12167);
nand U14585 (N_14585,N_10693,N_11763);
nand U14586 (N_14586,N_11878,N_11638);
nor U14587 (N_14587,N_11738,N_11521);
nor U14588 (N_14588,N_12481,N_12093);
nor U14589 (N_14589,N_11680,N_10210);
xnor U14590 (N_14590,N_12035,N_12170);
and U14591 (N_14591,N_11412,N_10865);
and U14592 (N_14592,N_10193,N_10901);
and U14593 (N_14593,N_12145,N_10782);
xnor U14594 (N_14594,N_12496,N_11460);
nor U14595 (N_14595,N_11679,N_11198);
or U14596 (N_14596,N_11373,N_12480);
and U14597 (N_14597,N_10084,N_11031);
nand U14598 (N_14598,N_11435,N_10052);
or U14599 (N_14599,N_11633,N_11339);
and U14600 (N_14600,N_11096,N_11161);
or U14601 (N_14601,N_10428,N_12155);
nor U14602 (N_14602,N_10757,N_12066);
nand U14603 (N_14603,N_12241,N_10272);
nor U14604 (N_14604,N_11511,N_10585);
nand U14605 (N_14605,N_11843,N_12166);
nand U14606 (N_14606,N_11099,N_10798);
nor U14607 (N_14607,N_12478,N_12073);
or U14608 (N_14608,N_10731,N_12447);
or U14609 (N_14609,N_11665,N_11149);
xor U14610 (N_14610,N_10102,N_10148);
nor U14611 (N_14611,N_11444,N_11816);
nand U14612 (N_14612,N_12116,N_11034);
or U14613 (N_14613,N_10972,N_11775);
xnor U14614 (N_14614,N_10771,N_12433);
nand U14615 (N_14615,N_10020,N_10336);
xor U14616 (N_14616,N_10566,N_12101);
xnor U14617 (N_14617,N_10882,N_12473);
and U14618 (N_14618,N_11463,N_11456);
or U14619 (N_14619,N_11845,N_10094);
xnor U14620 (N_14620,N_10464,N_11918);
or U14621 (N_14621,N_10214,N_11731);
nor U14622 (N_14622,N_10276,N_11899);
xnor U14623 (N_14623,N_12296,N_11147);
xor U14624 (N_14624,N_11178,N_10264);
or U14625 (N_14625,N_11345,N_10699);
xor U14626 (N_14626,N_11835,N_10555);
xnor U14627 (N_14627,N_12029,N_10589);
xnor U14628 (N_14628,N_11987,N_10572);
nor U14629 (N_14629,N_11330,N_10403);
or U14630 (N_14630,N_10819,N_10977);
nor U14631 (N_14631,N_11223,N_11893);
and U14632 (N_14632,N_11100,N_11806);
nand U14633 (N_14633,N_10644,N_11491);
and U14634 (N_14634,N_10002,N_11818);
xor U14635 (N_14635,N_10847,N_10949);
or U14636 (N_14636,N_10817,N_11250);
nand U14637 (N_14637,N_12477,N_12324);
nor U14638 (N_14638,N_11896,N_11826);
xnor U14639 (N_14639,N_10224,N_12252);
xor U14640 (N_14640,N_11415,N_11047);
nor U14641 (N_14641,N_11544,N_12493);
nand U14642 (N_14642,N_11215,N_12453);
xnor U14643 (N_14643,N_10785,N_10021);
nor U14644 (N_14644,N_12082,N_11380);
xnor U14645 (N_14645,N_10088,N_12161);
and U14646 (N_14646,N_10724,N_10602);
nor U14647 (N_14647,N_11639,N_10456);
or U14648 (N_14648,N_11493,N_11725);
nor U14649 (N_14649,N_11683,N_11569);
nor U14650 (N_14650,N_10270,N_12013);
nand U14651 (N_14651,N_10801,N_10849);
or U14652 (N_14652,N_11369,N_12406);
xor U14653 (N_14653,N_10331,N_10944);
xnor U14654 (N_14654,N_11626,N_10659);
nor U14655 (N_14655,N_11623,N_11683);
or U14656 (N_14656,N_10688,N_11054);
nand U14657 (N_14657,N_11604,N_11832);
nor U14658 (N_14658,N_11909,N_10944);
xor U14659 (N_14659,N_10704,N_10902);
nand U14660 (N_14660,N_11438,N_11232);
xnor U14661 (N_14661,N_10758,N_12203);
and U14662 (N_14662,N_12343,N_11522);
nand U14663 (N_14663,N_11865,N_11134);
xnor U14664 (N_14664,N_11860,N_10469);
nand U14665 (N_14665,N_12127,N_10278);
or U14666 (N_14666,N_10041,N_11011);
and U14667 (N_14667,N_11106,N_12271);
nor U14668 (N_14668,N_10390,N_10506);
xnor U14669 (N_14669,N_11687,N_10106);
xnor U14670 (N_14670,N_10839,N_11165);
and U14671 (N_14671,N_10763,N_10224);
xnor U14672 (N_14672,N_11127,N_11776);
and U14673 (N_14673,N_12317,N_11218);
and U14674 (N_14674,N_11262,N_10560);
or U14675 (N_14675,N_12016,N_12340);
and U14676 (N_14676,N_12205,N_10621);
and U14677 (N_14677,N_12009,N_10288);
nand U14678 (N_14678,N_11739,N_11806);
nor U14679 (N_14679,N_10834,N_10888);
xnor U14680 (N_14680,N_11609,N_12380);
or U14681 (N_14681,N_10157,N_11829);
or U14682 (N_14682,N_10883,N_11341);
or U14683 (N_14683,N_10286,N_12126);
xor U14684 (N_14684,N_12004,N_11688);
nor U14685 (N_14685,N_11881,N_11275);
or U14686 (N_14686,N_10927,N_10144);
nor U14687 (N_14687,N_10009,N_10578);
nor U14688 (N_14688,N_11097,N_11930);
nor U14689 (N_14689,N_10436,N_10184);
nand U14690 (N_14690,N_11973,N_11957);
or U14691 (N_14691,N_11315,N_11693);
and U14692 (N_14692,N_10800,N_10131);
nor U14693 (N_14693,N_10528,N_12253);
nor U14694 (N_14694,N_10940,N_10317);
xor U14695 (N_14695,N_10985,N_11864);
nand U14696 (N_14696,N_12050,N_10101);
or U14697 (N_14697,N_11273,N_10679);
and U14698 (N_14698,N_10994,N_11132);
nand U14699 (N_14699,N_11201,N_10797);
nor U14700 (N_14700,N_10344,N_10511);
or U14701 (N_14701,N_10730,N_10177);
or U14702 (N_14702,N_10325,N_10587);
nor U14703 (N_14703,N_10883,N_10936);
nor U14704 (N_14704,N_10912,N_11138);
or U14705 (N_14705,N_11713,N_10366);
and U14706 (N_14706,N_10493,N_11511);
nor U14707 (N_14707,N_10394,N_11127);
or U14708 (N_14708,N_10927,N_11161);
nand U14709 (N_14709,N_10968,N_12164);
nor U14710 (N_14710,N_11529,N_10109);
and U14711 (N_14711,N_12208,N_10984);
or U14712 (N_14712,N_12052,N_11750);
nor U14713 (N_14713,N_10631,N_10339);
nor U14714 (N_14714,N_11445,N_11957);
nor U14715 (N_14715,N_10162,N_11628);
nor U14716 (N_14716,N_11397,N_10255);
nor U14717 (N_14717,N_11989,N_12453);
or U14718 (N_14718,N_11482,N_12354);
and U14719 (N_14719,N_12124,N_11254);
or U14720 (N_14720,N_11612,N_10511);
and U14721 (N_14721,N_10871,N_12306);
nand U14722 (N_14722,N_12491,N_11794);
nor U14723 (N_14723,N_11374,N_10235);
nand U14724 (N_14724,N_10121,N_10381);
and U14725 (N_14725,N_10846,N_11683);
nor U14726 (N_14726,N_10317,N_10575);
nor U14727 (N_14727,N_11003,N_10607);
or U14728 (N_14728,N_10637,N_10842);
nand U14729 (N_14729,N_10957,N_11106);
or U14730 (N_14730,N_11946,N_10324);
or U14731 (N_14731,N_12227,N_10965);
xor U14732 (N_14732,N_11533,N_12131);
xnor U14733 (N_14733,N_11361,N_10246);
xor U14734 (N_14734,N_10140,N_12292);
and U14735 (N_14735,N_10013,N_11749);
nor U14736 (N_14736,N_12392,N_11493);
nand U14737 (N_14737,N_10715,N_12097);
xnor U14738 (N_14738,N_11201,N_11160);
nand U14739 (N_14739,N_11618,N_12277);
xnor U14740 (N_14740,N_10296,N_10375);
nor U14741 (N_14741,N_10653,N_11567);
and U14742 (N_14742,N_10306,N_10010);
or U14743 (N_14743,N_11304,N_11998);
nand U14744 (N_14744,N_10492,N_11262);
nand U14745 (N_14745,N_11181,N_12170);
nand U14746 (N_14746,N_12280,N_11032);
xor U14747 (N_14747,N_10326,N_11263);
or U14748 (N_14748,N_12367,N_11296);
xnor U14749 (N_14749,N_10276,N_10008);
nor U14750 (N_14750,N_11817,N_10475);
and U14751 (N_14751,N_12017,N_11293);
and U14752 (N_14752,N_10991,N_11656);
xnor U14753 (N_14753,N_11180,N_10590);
or U14754 (N_14754,N_10904,N_11653);
nor U14755 (N_14755,N_10509,N_12177);
or U14756 (N_14756,N_10370,N_11988);
nand U14757 (N_14757,N_10846,N_10009);
and U14758 (N_14758,N_12399,N_10003);
xor U14759 (N_14759,N_10059,N_11113);
xor U14760 (N_14760,N_10406,N_11630);
or U14761 (N_14761,N_10680,N_11241);
nand U14762 (N_14762,N_11397,N_12409);
nand U14763 (N_14763,N_10737,N_12324);
or U14764 (N_14764,N_11331,N_12374);
and U14765 (N_14765,N_10300,N_10338);
or U14766 (N_14766,N_12120,N_10390);
xnor U14767 (N_14767,N_12181,N_11479);
and U14768 (N_14768,N_11447,N_10342);
or U14769 (N_14769,N_11016,N_11411);
nand U14770 (N_14770,N_11701,N_10595);
or U14771 (N_14771,N_11500,N_11455);
and U14772 (N_14772,N_12005,N_12113);
and U14773 (N_14773,N_11585,N_11114);
xnor U14774 (N_14774,N_10453,N_10610);
and U14775 (N_14775,N_11237,N_11949);
or U14776 (N_14776,N_11373,N_12472);
nand U14777 (N_14777,N_12203,N_11924);
nor U14778 (N_14778,N_11865,N_11226);
nand U14779 (N_14779,N_11974,N_12115);
nor U14780 (N_14780,N_10449,N_11452);
xor U14781 (N_14781,N_10133,N_10516);
or U14782 (N_14782,N_10732,N_11601);
nor U14783 (N_14783,N_11549,N_10341);
nor U14784 (N_14784,N_10427,N_10792);
nor U14785 (N_14785,N_11564,N_10859);
nor U14786 (N_14786,N_10239,N_12155);
xnor U14787 (N_14787,N_10120,N_11732);
nor U14788 (N_14788,N_11020,N_11181);
and U14789 (N_14789,N_10155,N_10003);
xor U14790 (N_14790,N_12266,N_10207);
xor U14791 (N_14791,N_10170,N_10158);
nor U14792 (N_14792,N_10102,N_11560);
and U14793 (N_14793,N_10920,N_10788);
and U14794 (N_14794,N_11663,N_11112);
xnor U14795 (N_14795,N_11731,N_12028);
or U14796 (N_14796,N_11081,N_10613);
nor U14797 (N_14797,N_12458,N_10530);
nand U14798 (N_14798,N_10955,N_12442);
and U14799 (N_14799,N_10723,N_10270);
or U14800 (N_14800,N_11401,N_10558);
xnor U14801 (N_14801,N_11981,N_11491);
or U14802 (N_14802,N_11577,N_11112);
nand U14803 (N_14803,N_11532,N_10102);
nand U14804 (N_14804,N_10426,N_10203);
nor U14805 (N_14805,N_10540,N_11626);
and U14806 (N_14806,N_10220,N_11103);
nor U14807 (N_14807,N_12058,N_10226);
xnor U14808 (N_14808,N_10660,N_10819);
nand U14809 (N_14809,N_11705,N_11701);
nand U14810 (N_14810,N_11449,N_11819);
or U14811 (N_14811,N_11639,N_10354);
and U14812 (N_14812,N_10794,N_12244);
nand U14813 (N_14813,N_10673,N_10684);
and U14814 (N_14814,N_11723,N_10716);
nor U14815 (N_14815,N_10047,N_10525);
or U14816 (N_14816,N_12272,N_10504);
or U14817 (N_14817,N_12088,N_11649);
nand U14818 (N_14818,N_12014,N_11991);
and U14819 (N_14819,N_11164,N_11460);
xnor U14820 (N_14820,N_10944,N_12466);
or U14821 (N_14821,N_11676,N_11828);
or U14822 (N_14822,N_11482,N_12187);
nand U14823 (N_14823,N_10579,N_10781);
or U14824 (N_14824,N_11002,N_11668);
and U14825 (N_14825,N_12114,N_11052);
nand U14826 (N_14826,N_11419,N_10052);
xor U14827 (N_14827,N_10272,N_11774);
and U14828 (N_14828,N_10784,N_10132);
nor U14829 (N_14829,N_12322,N_10799);
xor U14830 (N_14830,N_12236,N_10876);
nand U14831 (N_14831,N_11854,N_12146);
or U14832 (N_14832,N_11886,N_10876);
or U14833 (N_14833,N_10094,N_10794);
nand U14834 (N_14834,N_12407,N_11606);
nor U14835 (N_14835,N_10957,N_11849);
and U14836 (N_14836,N_11207,N_10538);
nor U14837 (N_14837,N_11713,N_11792);
nor U14838 (N_14838,N_12285,N_11031);
and U14839 (N_14839,N_12341,N_10986);
nor U14840 (N_14840,N_12289,N_12040);
nand U14841 (N_14841,N_12450,N_11245);
xnor U14842 (N_14842,N_10317,N_11420);
and U14843 (N_14843,N_10091,N_10084);
nor U14844 (N_14844,N_11689,N_11538);
nand U14845 (N_14845,N_11007,N_10426);
and U14846 (N_14846,N_10476,N_12435);
and U14847 (N_14847,N_11774,N_10552);
or U14848 (N_14848,N_11649,N_10131);
xor U14849 (N_14849,N_10889,N_10025);
nand U14850 (N_14850,N_11465,N_11991);
and U14851 (N_14851,N_11448,N_12389);
and U14852 (N_14852,N_10606,N_10464);
and U14853 (N_14853,N_11948,N_11380);
xor U14854 (N_14854,N_11882,N_10322);
nand U14855 (N_14855,N_11497,N_11692);
nand U14856 (N_14856,N_12163,N_10937);
nand U14857 (N_14857,N_10082,N_12268);
nor U14858 (N_14858,N_12305,N_11462);
nand U14859 (N_14859,N_12391,N_12498);
xor U14860 (N_14860,N_10919,N_11253);
and U14861 (N_14861,N_11890,N_11797);
nand U14862 (N_14862,N_11999,N_11415);
and U14863 (N_14863,N_12093,N_10590);
nand U14864 (N_14864,N_11478,N_10896);
or U14865 (N_14865,N_11948,N_11111);
xor U14866 (N_14866,N_11306,N_10640);
nand U14867 (N_14867,N_11132,N_11913);
nor U14868 (N_14868,N_12273,N_11730);
or U14869 (N_14869,N_11202,N_11579);
and U14870 (N_14870,N_10869,N_11131);
xor U14871 (N_14871,N_10726,N_12274);
nand U14872 (N_14872,N_11889,N_11245);
or U14873 (N_14873,N_11159,N_11672);
xnor U14874 (N_14874,N_12235,N_11598);
nand U14875 (N_14875,N_12449,N_10536);
and U14876 (N_14876,N_10747,N_12431);
and U14877 (N_14877,N_10452,N_12059);
xor U14878 (N_14878,N_10626,N_11561);
nor U14879 (N_14879,N_11804,N_11016);
nand U14880 (N_14880,N_11184,N_11679);
nand U14881 (N_14881,N_11286,N_11280);
nor U14882 (N_14882,N_11895,N_10417);
and U14883 (N_14883,N_11211,N_10593);
or U14884 (N_14884,N_10774,N_11024);
nor U14885 (N_14885,N_11792,N_10080);
xnor U14886 (N_14886,N_10680,N_10936);
and U14887 (N_14887,N_11440,N_12193);
or U14888 (N_14888,N_12158,N_11112);
nor U14889 (N_14889,N_12436,N_10039);
and U14890 (N_14890,N_11693,N_11935);
nand U14891 (N_14891,N_12157,N_10867);
nor U14892 (N_14892,N_12183,N_11350);
or U14893 (N_14893,N_11757,N_11881);
xor U14894 (N_14894,N_12363,N_12092);
and U14895 (N_14895,N_11438,N_11785);
nor U14896 (N_14896,N_10690,N_11432);
or U14897 (N_14897,N_11605,N_11460);
and U14898 (N_14898,N_11840,N_11696);
and U14899 (N_14899,N_11587,N_11035);
xor U14900 (N_14900,N_11730,N_10899);
xor U14901 (N_14901,N_11986,N_10573);
and U14902 (N_14902,N_10227,N_11089);
xnor U14903 (N_14903,N_10390,N_10325);
or U14904 (N_14904,N_10081,N_10012);
xnor U14905 (N_14905,N_12445,N_10043);
or U14906 (N_14906,N_11306,N_11114);
nand U14907 (N_14907,N_10702,N_11833);
and U14908 (N_14908,N_10055,N_11277);
xnor U14909 (N_14909,N_11453,N_12215);
xnor U14910 (N_14910,N_11917,N_10095);
and U14911 (N_14911,N_10589,N_10362);
xnor U14912 (N_14912,N_10662,N_12125);
xor U14913 (N_14913,N_12116,N_10836);
xnor U14914 (N_14914,N_11502,N_11246);
or U14915 (N_14915,N_10426,N_11598);
nand U14916 (N_14916,N_11066,N_12498);
and U14917 (N_14917,N_10505,N_10794);
or U14918 (N_14918,N_10818,N_11046);
or U14919 (N_14919,N_12136,N_10929);
nor U14920 (N_14920,N_10681,N_11683);
or U14921 (N_14921,N_12462,N_10364);
and U14922 (N_14922,N_11811,N_10286);
nand U14923 (N_14923,N_11945,N_10769);
and U14924 (N_14924,N_11967,N_11254);
nand U14925 (N_14925,N_12383,N_10568);
and U14926 (N_14926,N_10781,N_10553);
xnor U14927 (N_14927,N_11700,N_11918);
nor U14928 (N_14928,N_11307,N_10825);
and U14929 (N_14929,N_10121,N_10154);
xnor U14930 (N_14930,N_12110,N_11199);
xnor U14931 (N_14931,N_12476,N_10712);
xor U14932 (N_14932,N_12113,N_10663);
or U14933 (N_14933,N_10032,N_10079);
and U14934 (N_14934,N_10882,N_11252);
and U14935 (N_14935,N_11284,N_10918);
or U14936 (N_14936,N_12401,N_11140);
or U14937 (N_14937,N_11455,N_11350);
nand U14938 (N_14938,N_11778,N_11776);
nand U14939 (N_14939,N_10110,N_10353);
xnor U14940 (N_14940,N_10869,N_11172);
or U14941 (N_14941,N_11295,N_11963);
nor U14942 (N_14942,N_10483,N_11098);
xor U14943 (N_14943,N_11806,N_10918);
nor U14944 (N_14944,N_11332,N_12174);
nand U14945 (N_14945,N_11525,N_10362);
xnor U14946 (N_14946,N_12222,N_11599);
or U14947 (N_14947,N_10817,N_11297);
nand U14948 (N_14948,N_10221,N_12097);
nor U14949 (N_14949,N_11768,N_11436);
nand U14950 (N_14950,N_11215,N_11715);
or U14951 (N_14951,N_10237,N_12389);
and U14952 (N_14952,N_12171,N_11328);
xor U14953 (N_14953,N_10958,N_11877);
or U14954 (N_14954,N_10782,N_10837);
nand U14955 (N_14955,N_12236,N_10675);
nand U14956 (N_14956,N_10508,N_12188);
or U14957 (N_14957,N_11871,N_10947);
or U14958 (N_14958,N_10668,N_10743);
nand U14959 (N_14959,N_11902,N_12419);
nor U14960 (N_14960,N_11150,N_11895);
nor U14961 (N_14961,N_11944,N_10030);
and U14962 (N_14962,N_11975,N_11015);
nand U14963 (N_14963,N_10720,N_10908);
nand U14964 (N_14964,N_11264,N_10932);
nor U14965 (N_14965,N_11916,N_11968);
nor U14966 (N_14966,N_10856,N_10944);
xor U14967 (N_14967,N_11863,N_10426);
xor U14968 (N_14968,N_11367,N_10720);
and U14969 (N_14969,N_10519,N_10715);
nand U14970 (N_14970,N_10687,N_10126);
nor U14971 (N_14971,N_11959,N_10902);
nand U14972 (N_14972,N_10025,N_10088);
and U14973 (N_14973,N_11694,N_10580);
or U14974 (N_14974,N_11621,N_11511);
or U14975 (N_14975,N_12130,N_12481);
nor U14976 (N_14976,N_10037,N_11864);
nand U14977 (N_14977,N_10845,N_12032);
and U14978 (N_14978,N_12186,N_11531);
or U14979 (N_14979,N_10408,N_10039);
or U14980 (N_14980,N_11414,N_12246);
xor U14981 (N_14981,N_10133,N_12290);
and U14982 (N_14982,N_10545,N_10921);
or U14983 (N_14983,N_12403,N_10389);
xor U14984 (N_14984,N_11239,N_11978);
nand U14985 (N_14985,N_11246,N_10028);
or U14986 (N_14986,N_11483,N_10968);
nand U14987 (N_14987,N_11968,N_10334);
and U14988 (N_14988,N_10748,N_10637);
and U14989 (N_14989,N_11980,N_10662);
nand U14990 (N_14990,N_12069,N_11044);
or U14991 (N_14991,N_11355,N_11270);
nand U14992 (N_14992,N_11942,N_10351);
nand U14993 (N_14993,N_12411,N_11245);
or U14994 (N_14994,N_12171,N_11172);
nor U14995 (N_14995,N_11939,N_12033);
and U14996 (N_14996,N_10691,N_11929);
xnor U14997 (N_14997,N_12394,N_12484);
nand U14998 (N_14998,N_10523,N_10815);
xor U14999 (N_14999,N_10352,N_11108);
nor U15000 (N_15000,N_14758,N_14711);
nor U15001 (N_15001,N_13190,N_13950);
or U15002 (N_15002,N_14968,N_14942);
nand U15003 (N_15003,N_14755,N_13500);
nand U15004 (N_15004,N_14715,N_14527);
and U15005 (N_15005,N_13936,N_13405);
nand U15006 (N_15006,N_12522,N_12952);
or U15007 (N_15007,N_12515,N_12629);
or U15008 (N_15008,N_14111,N_14677);
or U15009 (N_15009,N_13513,N_13856);
nor U15010 (N_15010,N_14145,N_14375);
and U15011 (N_15011,N_14702,N_12760);
or U15012 (N_15012,N_14869,N_13421);
or U15013 (N_15013,N_12525,N_14509);
or U15014 (N_15014,N_14587,N_13084);
or U15015 (N_15015,N_13613,N_14633);
nand U15016 (N_15016,N_13952,N_13282);
and U15017 (N_15017,N_14689,N_13733);
and U15018 (N_15018,N_13690,N_14867);
nor U15019 (N_15019,N_14381,N_13675);
nor U15020 (N_15020,N_13018,N_13932);
nand U15021 (N_15021,N_14638,N_13959);
or U15022 (N_15022,N_14893,N_12813);
nor U15023 (N_15023,N_13633,N_14811);
nand U15024 (N_15024,N_12891,N_12580);
nor U15025 (N_15025,N_13810,N_13904);
nor U15026 (N_15026,N_12610,N_13585);
or U15027 (N_15027,N_13641,N_14520);
and U15028 (N_15028,N_13830,N_12634);
xor U15029 (N_15029,N_13109,N_14993);
nand U15030 (N_15030,N_14778,N_13747);
nand U15031 (N_15031,N_14861,N_12696);
xor U15032 (N_15032,N_13409,N_14110);
nor U15033 (N_15033,N_13578,N_14733);
nor U15034 (N_15034,N_12500,N_13668);
nor U15035 (N_15035,N_13478,N_12518);
and U15036 (N_15036,N_13678,N_13411);
or U15037 (N_15037,N_14316,N_13499);
nand U15038 (N_15038,N_13744,N_13473);
and U15039 (N_15039,N_14529,N_14089);
and U15040 (N_15040,N_13078,N_13134);
nor U15041 (N_15041,N_12882,N_13883);
nor U15042 (N_15042,N_14822,N_13593);
xnor U15043 (N_15043,N_14370,N_13820);
nor U15044 (N_15044,N_13958,N_14078);
nand U15045 (N_15045,N_13099,N_14443);
nand U15046 (N_15046,N_13406,N_13779);
and U15047 (N_15047,N_12674,N_13325);
xor U15048 (N_15048,N_14799,N_13617);
or U15049 (N_15049,N_13376,N_13843);
nor U15050 (N_15050,N_13080,N_13535);
and U15051 (N_15051,N_12709,N_14308);
or U15052 (N_15052,N_13941,N_12627);
and U15053 (N_15053,N_12785,N_14567);
nor U15054 (N_15054,N_14232,N_13789);
xor U15055 (N_15055,N_14432,N_14069);
nand U15056 (N_15056,N_12700,N_12579);
xnor U15057 (N_15057,N_12663,N_12915);
and U15058 (N_15058,N_13981,N_12756);
nand U15059 (N_15059,N_13157,N_12927);
or U15060 (N_15060,N_14900,N_14137);
nand U15061 (N_15061,N_14810,N_13693);
or U15062 (N_15062,N_14598,N_12514);
nor U15063 (N_15063,N_14533,N_14314);
nand U15064 (N_15064,N_14318,N_13854);
nand U15065 (N_15065,N_13168,N_13603);
xor U15066 (N_15066,N_13644,N_14305);
nor U15067 (N_15067,N_13247,N_13284);
and U15068 (N_15068,N_12949,N_14401);
and U15069 (N_15069,N_13555,N_14100);
or U15070 (N_15070,N_13433,N_12805);
nor U15071 (N_15071,N_13306,N_12622);
or U15072 (N_15072,N_14769,N_13703);
or U15073 (N_15073,N_13447,N_14120);
nor U15074 (N_15074,N_14940,N_14597);
xor U15075 (N_15075,N_14061,N_12816);
or U15076 (N_15076,N_14131,N_13750);
nand U15077 (N_15077,N_12963,N_13751);
xnor U15078 (N_15078,N_13058,N_13017);
xor U15079 (N_15079,N_13766,N_13414);
and U15080 (N_15080,N_14717,N_14691);
xnor U15081 (N_15081,N_12631,N_14267);
and U15082 (N_15082,N_14295,N_13313);
nand U15083 (N_15083,N_12691,N_14133);
and U15084 (N_15084,N_13418,N_12746);
or U15085 (N_15085,N_13492,N_13087);
and U15086 (N_15086,N_13467,N_14122);
nor U15087 (N_15087,N_14282,N_12985);
and U15088 (N_15088,N_14704,N_12635);
or U15089 (N_15089,N_14135,N_13713);
nand U15090 (N_15090,N_12716,N_12777);
xor U15091 (N_15091,N_14724,N_12980);
or U15092 (N_15092,N_12779,N_13209);
nand U15093 (N_15093,N_14080,N_12831);
and U15094 (N_15094,N_14038,N_12844);
nor U15095 (N_15095,N_13665,N_13090);
nand U15096 (N_15096,N_14088,N_14035);
or U15097 (N_15097,N_14218,N_12786);
nor U15098 (N_15098,N_12718,N_14700);
and U15099 (N_15099,N_12841,N_13022);
xor U15100 (N_15100,N_12724,N_12898);
and U15101 (N_15101,N_14323,N_14837);
and U15102 (N_15102,N_12600,N_14436);
or U15103 (N_15103,N_14410,N_12834);
or U15104 (N_15104,N_13587,N_13841);
nand U15105 (N_15105,N_12537,N_14846);
xnor U15106 (N_15106,N_14913,N_14173);
and U15107 (N_15107,N_13494,N_13538);
and U15108 (N_15108,N_14430,N_14506);
nor U15109 (N_15109,N_12945,N_13000);
nand U15110 (N_15110,N_13649,N_14586);
nor U15111 (N_15111,N_14224,N_14979);
xor U15112 (N_15112,N_13217,N_14439);
or U15113 (N_15113,N_14771,N_14682);
and U15114 (N_15114,N_13749,N_13575);
nand U15115 (N_15115,N_14376,N_14756);
and U15116 (N_15116,N_13752,N_14823);
nand U15117 (N_15117,N_13549,N_13577);
nand U15118 (N_15118,N_12860,N_13455);
nand U15119 (N_15119,N_13480,N_14132);
nand U15120 (N_15120,N_12658,N_13975);
xnor U15121 (N_15121,N_14334,N_12902);
nand U15122 (N_15122,N_13586,N_12955);
xor U15123 (N_15123,N_14855,N_14413);
nand U15124 (N_15124,N_14337,N_14492);
and U15125 (N_15125,N_12884,N_13025);
nor U15126 (N_15126,N_14783,N_14141);
and U15127 (N_15127,N_13312,N_13427);
nand U15128 (N_15128,N_13785,N_14876);
or U15129 (N_15129,N_13802,N_13239);
nand U15130 (N_15130,N_14419,N_13914);
and U15131 (N_15131,N_13263,N_13510);
nand U15132 (N_15132,N_13694,N_14858);
or U15133 (N_15133,N_13702,N_14695);
xnor U15134 (N_15134,N_12912,N_12977);
nand U15135 (N_15135,N_13194,N_13234);
or U15136 (N_15136,N_14409,N_14726);
or U15137 (N_15137,N_12685,N_14243);
and U15138 (N_15138,N_13884,N_13011);
nor U15139 (N_15139,N_14641,N_12857);
and U15140 (N_15140,N_14657,N_14910);
nor U15141 (N_15141,N_12976,N_14891);
xnor U15142 (N_15142,N_12588,N_13536);
nor U15143 (N_15143,N_13149,N_14997);
or U15144 (N_15144,N_14971,N_13051);
or U15145 (N_15145,N_13572,N_13591);
nand U15146 (N_15146,N_14601,N_13021);
nand U15147 (N_15147,N_14222,N_13137);
and U15148 (N_15148,N_12798,N_13470);
and U15149 (N_15149,N_14546,N_13272);
xnor U15150 (N_15150,N_13806,N_13348);
xor U15151 (N_15151,N_13908,N_13684);
nor U15152 (N_15152,N_13122,N_14919);
nand U15153 (N_15153,N_13285,N_12584);
nand U15154 (N_15154,N_13446,N_14906);
or U15155 (N_15155,N_14216,N_14670);
nor U15156 (N_15156,N_13745,N_13291);
and U15157 (N_15157,N_13023,N_13488);
or U15158 (N_15158,N_13029,N_14459);
xor U15159 (N_15159,N_13125,N_14552);
and U15160 (N_15160,N_14285,N_12863);
and U15161 (N_15161,N_14404,N_12865);
and U15162 (N_15162,N_14373,N_13777);
nor U15163 (N_15163,N_14757,N_14904);
and U15164 (N_15164,N_14475,N_14693);
and U15165 (N_15165,N_13191,N_13174);
or U15166 (N_15166,N_14836,N_14315);
nand U15167 (N_15167,N_12747,N_12710);
or U15168 (N_15168,N_13660,N_14452);
xnor U15169 (N_15169,N_14607,N_12640);
nor U15170 (N_15170,N_13482,N_13337);
or U15171 (N_15171,N_13623,N_14444);
nand U15172 (N_15172,N_13120,N_13842);
nand U15173 (N_15173,N_13160,N_13228);
nor U15174 (N_15174,N_12883,N_14818);
and U15175 (N_15175,N_14467,N_14049);
nand U15176 (N_15176,N_13179,N_14253);
xnor U15177 (N_15177,N_12571,N_14191);
nand U15178 (N_15178,N_12984,N_14204);
nand U15179 (N_15179,N_12970,N_14562);
xnor U15180 (N_15180,N_14515,N_13972);
nand U15181 (N_15181,N_12767,N_14147);
nor U15182 (N_15182,N_13844,N_13701);
xor U15183 (N_15183,N_12827,N_12543);
xnor U15184 (N_15184,N_14923,N_14931);
nand U15185 (N_15185,N_14990,N_12505);
xor U15186 (N_15186,N_13044,N_14096);
and U15187 (N_15187,N_13268,N_13154);
nor U15188 (N_15188,N_12694,N_13771);
or U15189 (N_15189,N_14938,N_14000);
nor U15190 (N_15190,N_12601,N_14539);
xor U15191 (N_15191,N_14849,N_14604);
nor U15192 (N_15192,N_14551,N_14673);
nor U15193 (N_15193,N_14434,N_13569);
nand U15194 (N_15194,N_13260,N_13719);
and U15195 (N_15195,N_13740,N_13273);
and U15196 (N_15196,N_12665,N_14431);
or U15197 (N_15197,N_14076,N_14197);
and U15198 (N_15198,N_14384,N_14781);
xor U15199 (N_15199,N_13695,N_14297);
nor U15200 (N_15200,N_13930,N_14885);
nand U15201 (N_15201,N_14887,N_14543);
and U15202 (N_15202,N_14895,N_12699);
nand U15203 (N_15203,N_14268,N_13115);
nor U15204 (N_15204,N_14104,N_12837);
and U15205 (N_15205,N_14421,N_14064);
nand U15206 (N_15206,N_14366,N_14044);
or U15207 (N_15207,N_13159,N_12649);
nor U15208 (N_15208,N_12692,N_12679);
xnor U15209 (N_15209,N_14451,N_14616);
xor U15210 (N_15210,N_12973,N_13636);
xor U15211 (N_15211,N_14981,N_14725);
and U15212 (N_15212,N_13146,N_14889);
xnor U15213 (N_15213,N_14896,N_14025);
xnor U15214 (N_15214,N_13040,N_14720);
or U15215 (N_15215,N_14200,N_13919);
nand U15216 (N_15216,N_14456,N_14507);
and U15217 (N_15217,N_13170,N_14531);
and U15218 (N_15218,N_13755,N_14738);
nor U15219 (N_15219,N_14184,N_12639);
nor U15220 (N_15220,N_14019,N_14559);
and U15221 (N_15221,N_14140,N_13805);
and U15222 (N_15222,N_14462,N_14407);
xor U15223 (N_15223,N_14261,N_13869);
xor U15224 (N_15224,N_12757,N_14329);
and U15225 (N_15225,N_12962,N_14223);
xor U15226 (N_15226,N_14010,N_14399);
and U15227 (N_15227,N_13836,N_14206);
xnor U15228 (N_15228,N_14944,N_14103);
and U15229 (N_15229,N_14390,N_14231);
xor U15230 (N_15230,N_13033,N_14678);
and U15231 (N_15231,N_13429,N_12565);
nor U15232 (N_15232,N_13768,N_14927);
nor U15233 (N_15233,N_13294,N_14383);
xnor U15234 (N_15234,N_12881,N_13308);
nand U15235 (N_15235,N_14335,N_13722);
or U15236 (N_15236,N_12540,N_14554);
xor U15237 (N_15237,N_14987,N_12788);
nand U15238 (N_15238,N_14663,N_14012);
or U15239 (N_15239,N_14826,N_14360);
xor U15240 (N_15240,N_12596,N_13725);
or U15241 (N_15241,N_14631,N_13351);
or U15242 (N_15242,N_13232,N_12890);
nor U15243 (N_15243,N_14408,N_12676);
nand U15244 (N_15244,N_14379,N_13413);
nor U15245 (N_15245,N_14589,N_14542);
and U15246 (N_15246,N_13412,N_14377);
xor U15247 (N_15247,N_13968,N_13692);
nor U15248 (N_15248,N_14310,N_13399);
nor U15249 (N_15249,N_12784,N_14468);
xnor U15250 (N_15250,N_14221,N_14264);
or U15251 (N_15251,N_12521,N_13622);
or U15252 (N_15252,N_14962,N_13092);
nand U15253 (N_15253,N_13946,N_13295);
nor U15254 (N_15254,N_13354,N_13542);
or U15255 (N_15255,N_14872,N_13948);
nand U15256 (N_15256,N_12545,N_12670);
or U15257 (N_15257,N_13073,N_13629);
nand U15258 (N_15258,N_13394,N_14945);
nand U15259 (N_15259,N_14692,N_13435);
or U15260 (N_15260,N_13821,N_13502);
and U15261 (N_15261,N_14512,N_12651);
nand U15262 (N_15262,N_13231,N_13955);
or U15263 (N_15263,N_13543,N_14679);
and U15264 (N_15264,N_13721,N_13216);
nand U15265 (N_15265,N_13043,N_13072);
xor U15266 (N_15266,N_14281,N_13226);
xor U15267 (N_15267,N_12808,N_13366);
and U15268 (N_15268,N_12939,N_14924);
nand U15269 (N_15269,N_13873,N_12541);
nor U15270 (N_15270,N_13527,N_13900);
xor U15271 (N_15271,N_13458,N_13550);
nor U15272 (N_15272,N_14814,N_14302);
or U15273 (N_15273,N_13410,N_12763);
nor U15274 (N_15274,N_14101,N_13403);
xor U15275 (N_15275,N_14193,N_12833);
nor U15276 (N_15276,N_13519,N_14414);
xor U15277 (N_15277,N_12899,N_14583);
xnor U15278 (N_15278,N_12737,N_12536);
and U15279 (N_15279,N_12698,N_14138);
and U15280 (N_15280,N_14721,N_13474);
xnor U15281 (N_15281,N_14211,N_14894);
or U15282 (N_15282,N_12971,N_13521);
xor U15283 (N_15283,N_13985,N_14652);
and U15284 (N_15284,N_14851,N_14286);
and U15285 (N_15285,N_13118,N_13734);
and U15286 (N_15286,N_14392,N_14819);
nor U15287 (N_15287,N_13392,N_14681);
nor U15288 (N_15288,N_13352,N_13003);
or U15289 (N_15289,N_13082,N_13404);
xnor U15290 (N_15290,N_13065,N_14006);
nor U15291 (N_15291,N_14427,N_13487);
and U15292 (N_15292,N_13143,N_14066);
nor U15293 (N_15293,N_14402,N_13726);
and U15294 (N_15294,N_12690,N_14943);
nor U15295 (N_15295,N_14621,N_13124);
and U15296 (N_15296,N_14859,N_14686);
nor U15297 (N_15297,N_14839,N_14510);
xor U15298 (N_15298,N_14807,N_13626);
nor U15299 (N_15299,N_12531,N_13566);
nand U15300 (N_15300,N_14538,N_14065);
xnor U15301 (N_15301,N_14608,N_13490);
and U15302 (N_15302,N_13992,N_14808);
and U15303 (N_15303,N_13200,N_13336);
or U15304 (N_15304,N_13012,N_13928);
and U15305 (N_15305,N_14087,N_13420);
xor U15306 (N_15306,N_14654,N_14151);
or U15307 (N_15307,N_14701,N_13748);
nor U15308 (N_15308,N_13653,N_13185);
nor U15309 (N_15309,N_13046,N_13434);
nor U15310 (N_15310,N_13286,N_14564);
nand U15311 (N_15311,N_13905,N_13901);
nor U15312 (N_15312,N_14494,N_14612);
or U15313 (N_15313,N_13288,N_12609);
and U15314 (N_15314,N_14320,N_13102);
nand U15315 (N_15315,N_14425,N_13620);
nand U15316 (N_15316,N_12678,N_13384);
nor U15317 (N_15317,N_14136,N_14134);
xnor U15318 (N_15318,N_14159,N_13552);
nor U15319 (N_15319,N_12569,N_14342);
and U15320 (N_15320,N_12815,N_13400);
nor U15321 (N_15321,N_13131,N_13982);
or U15322 (N_15322,N_12769,N_14916);
nand U15323 (N_15323,N_13426,N_12671);
xor U15324 (N_15324,N_14580,N_13172);
nand U15325 (N_15325,N_14610,N_14992);
or U15326 (N_15326,N_13350,N_12546);
xor U15327 (N_15327,N_14751,N_12607);
or U15328 (N_15328,N_13192,N_12944);
nand U15329 (N_15329,N_13370,N_14571);
and U15330 (N_15330,N_14759,N_12851);
and U15331 (N_15331,N_12697,N_13320);
or U15332 (N_15332,N_13704,N_13648);
nand U15333 (N_15333,N_14606,N_14176);
nor U15334 (N_15334,N_13775,N_12799);
nand U15335 (N_15335,N_13994,N_13706);
nor U15336 (N_15336,N_13442,N_13781);
xor U15337 (N_15337,N_13880,N_13503);
nand U15338 (N_15338,N_14745,N_13758);
nand U15339 (N_15339,N_12814,N_14048);
nor U15340 (N_15340,N_14125,N_13800);
nor U15341 (N_15341,N_12744,N_13515);
nand U15342 (N_15342,N_13189,N_12894);
nand U15343 (N_15343,N_13323,N_12858);
or U15344 (N_15344,N_14395,N_13865);
or U15345 (N_15345,N_14023,N_14675);
nor U15346 (N_15346,N_13452,N_14464);
nand U15347 (N_15347,N_14442,N_13221);
xor U15348 (N_15348,N_14278,N_13013);
nor U15349 (N_15349,N_14789,N_13266);
or U15350 (N_15350,N_12774,N_13047);
nand U15351 (N_15351,N_14473,N_12802);
or U15352 (N_15352,N_12503,N_12800);
xnor U15353 (N_15353,N_13727,N_14828);
nand U15354 (N_15354,N_14983,N_13643);
xnor U15355 (N_15355,N_12562,N_13275);
and U15356 (N_15356,N_13911,N_14341);
xor U15357 (N_15357,N_13604,N_14417);
xnor U15358 (N_15358,N_13113,N_13608);
nand U15359 (N_15359,N_14537,N_13846);
xnor U15360 (N_15360,N_13395,N_14747);
nand U15361 (N_15361,N_12720,N_13056);
nor U15362 (N_15362,N_12938,N_13639);
nor U15363 (N_15363,N_14142,N_13888);
and U15364 (N_15364,N_13035,N_13529);
and U15365 (N_15365,N_14574,N_12783);
nand U15366 (N_15366,N_12553,N_13477);
and U15367 (N_15367,N_13416,N_12590);
nand U15368 (N_15368,N_12714,N_13679);
or U15369 (N_15369,N_14393,N_13178);
nor U15370 (N_15370,N_14478,N_13222);
nor U15371 (N_15371,N_13193,N_14929);
nor U15372 (N_15372,N_13516,N_14592);
and U15373 (N_15373,N_13879,N_12706);
and U15374 (N_15374,N_14732,N_12563);
nand U15375 (N_15375,N_14975,N_14832);
xnor U15376 (N_15376,N_14791,N_12761);
xor U15377 (N_15377,N_14293,N_13823);
nand U15378 (N_15378,N_14016,N_12673);
or U15379 (N_15379,N_12787,N_12793);
nand U15380 (N_15380,N_12603,N_14215);
or U15381 (N_15381,N_12990,N_13307);
or U15382 (N_15382,N_14058,N_14219);
or U15383 (N_15383,N_12869,N_13920);
nor U15384 (N_15384,N_13004,N_12758);
nand U15385 (N_15385,N_12872,N_13229);
or U15386 (N_15386,N_13737,N_12740);
xnor U15387 (N_15387,N_14042,N_13728);
or U15388 (N_15388,N_14426,N_13672);
and U15389 (N_15389,N_12701,N_13619);
or U15390 (N_15390,N_13832,N_12991);
xnor U15391 (N_15391,N_13889,N_13450);
nor U15392 (N_15392,N_14183,N_14797);
xnor U15393 (N_15393,N_14787,N_12958);
nor U15394 (N_15394,N_12886,N_14713);
and U15395 (N_15395,N_14594,N_12731);
nor U15396 (N_15396,N_14483,N_14180);
xnor U15397 (N_15397,N_12585,N_13738);
nand U15398 (N_15398,N_12832,N_13364);
nand U15399 (N_15399,N_14912,N_13206);
xnor U15400 (N_15400,N_12824,N_13026);
xor U15401 (N_15401,N_12549,N_13197);
nor U15402 (N_15402,N_13481,N_12910);
xor U15403 (N_15403,N_12994,N_12840);
xnor U15404 (N_15404,N_13436,N_14306);
nand U15405 (N_15405,N_14388,N_13390);
nor U15406 (N_15406,N_12736,N_14965);
or U15407 (N_15407,N_13997,N_14474);
or U15408 (N_15408,N_13696,N_13038);
xor U15409 (N_15409,N_14844,N_12982);
nand U15410 (N_15410,N_13973,N_14175);
and U15411 (N_15411,N_14071,N_13428);
or U15412 (N_15412,N_13098,N_14820);
and U15413 (N_15413,N_14767,N_14046);
or U15414 (N_15414,N_14578,N_13872);
and U15415 (N_15415,N_13592,N_14952);
nor U15416 (N_15416,N_12820,N_13015);
xor U15417 (N_15417,N_14772,N_13373);
nor U15418 (N_15418,N_12703,N_13505);
nand U15419 (N_15419,N_12809,N_12729);
and U15420 (N_15420,N_13934,N_13265);
nor U15421 (N_15421,N_13152,N_12797);
nand U15422 (N_15422,N_13990,N_12542);
or U15423 (N_15423,N_14057,N_14655);
or U15424 (N_15424,N_14047,N_14217);
and U15425 (N_15425,N_12589,N_14569);
xnor U15426 (N_15426,N_13215,N_12683);
and U15427 (N_15427,N_13573,N_13584);
xnor U15428 (N_15428,N_13835,N_14613);
and U15429 (N_15429,N_12501,N_13864);
and U15430 (N_15430,N_13321,N_14866);
xnor U15431 (N_15431,N_13735,N_13951);
and U15432 (N_15432,N_14547,N_13169);
nand U15433 (N_15433,N_13237,N_14291);
or U15434 (N_15434,N_13465,N_14174);
and U15435 (N_15435,N_13681,N_13594);
and U15436 (N_15436,N_12926,N_12509);
xnor U15437 (N_15437,N_14036,N_14073);
nand U15438 (N_15438,N_14031,N_12913);
nand U15439 (N_15439,N_12504,N_13117);
and U15440 (N_15440,N_12957,N_14922);
nor U15441 (N_15441,N_13016,N_14697);
nor U15442 (N_15442,N_14918,N_13059);
or U15443 (N_15443,N_13741,N_12707);
xnor U15444 (N_15444,N_14950,N_13655);
nand U15445 (N_15445,N_13518,N_13671);
nor U15446 (N_15446,N_14500,N_14167);
nand U15447 (N_15447,N_13548,N_13523);
or U15448 (N_15448,N_13258,N_14195);
nor U15449 (N_15449,N_12989,N_12901);
xnor U15450 (N_15450,N_13381,N_12878);
nand U15451 (N_15451,N_12550,N_13252);
xor U15452 (N_15452,N_14699,N_13890);
or U15453 (N_15453,N_14760,N_14123);
nand U15454 (N_15454,N_13441,N_12527);
or U15455 (N_15455,N_14244,N_12742);
and U15456 (N_15456,N_14269,N_13974);
and U15457 (N_15457,N_14661,N_13760);
and U15458 (N_15458,N_12682,N_14403);
nand U15459 (N_15459,N_13977,N_12659);
nor U15460 (N_15460,N_13184,N_13007);
or U15461 (N_15461,N_12893,N_13245);
nor U15462 (N_15462,N_13219,N_13097);
and U15463 (N_15463,N_13689,N_14157);
or U15464 (N_15464,N_13297,N_12576);
nand U15465 (N_15465,N_14476,N_12780);
nand U15466 (N_15466,N_14972,N_12932);
xor U15467 (N_15467,N_14158,N_14688);
and U15468 (N_15468,N_13534,N_12508);
nor U15469 (N_15469,N_13605,N_12992);
nor U15470 (N_15470,N_14513,N_13255);
xor U15471 (N_15471,N_14115,N_14982);
nand U15472 (N_15472,N_13627,N_14091);
nand U15473 (N_15473,N_12606,N_14812);
or U15474 (N_15474,N_14013,N_12595);
nand U15475 (N_15475,N_14234,N_14511);
nand U15476 (N_15476,N_14907,N_12561);
and U15477 (N_15477,N_13868,N_14346);
xor U15478 (N_15478,N_12544,N_13826);
and U15479 (N_15479,N_13368,N_14186);
or U15480 (N_15480,N_14275,N_14497);
xor U15481 (N_15481,N_14097,N_13378);
or U15482 (N_15482,N_14685,N_14203);
nand U15483 (N_15483,N_13698,N_13769);
and U15484 (N_15484,N_14094,N_12759);
and U15485 (N_15485,N_12904,N_14148);
nor U15486 (N_15486,N_13765,N_14082);
xor U15487 (N_15487,N_13181,N_13031);
nand U15488 (N_15488,N_13114,N_12829);
nor U15489 (N_15489,N_13171,N_12846);
xnor U15490 (N_15490,N_14365,N_14189);
xnor U15491 (N_15491,N_14072,N_13443);
or U15492 (N_15492,N_13077,N_14603);
and U15493 (N_15493,N_13156,N_14873);
or U15494 (N_15494,N_14909,N_13345);
or U15495 (N_15495,N_14027,N_13874);
nor U15496 (N_15496,N_13032,N_14934);
nor U15497 (N_15497,N_14116,N_13661);
nand U15498 (N_15498,N_14045,N_12885);
nand U15499 (N_15499,N_12920,N_14199);
or U15500 (N_15500,N_14448,N_13828);
xor U15501 (N_15501,N_13922,N_13054);
nor U15502 (N_15502,N_13819,N_13783);
nor U15503 (N_15503,N_12650,N_13281);
nand U15504 (N_15504,N_14770,N_12775);
xnor U15505 (N_15505,N_13961,N_12772);
xnor U15506 (N_15506,N_12613,N_14458);
xnor U15507 (N_15507,N_12727,N_14722);
and U15508 (N_15508,N_14878,N_13576);
xor U15509 (N_15509,N_14300,N_12717);
xnor U15510 (N_15510,N_12965,N_13532);
xor U15511 (N_15511,N_13243,N_13799);
nor U15512 (N_15512,N_12507,N_13896);
and U15513 (N_15513,N_14272,N_14821);
xnor U15514 (N_15514,N_14795,N_13244);
and U15515 (N_15515,N_12776,N_13290);
nand U15516 (N_15516,N_13978,N_13316);
or U15517 (N_15517,N_14398,N_12765);
and U15518 (N_15518,N_13496,N_13002);
and U15519 (N_15519,N_14505,N_13372);
and U15520 (N_15520,N_12535,N_12933);
xnor U15521 (N_15521,N_12752,N_14153);
xor U15522 (N_15522,N_12506,N_14773);
and U15523 (N_15523,N_13293,N_14668);
xor U15524 (N_15524,N_14532,N_13508);
nor U15525 (N_15525,N_13456,N_14709);
nand U15526 (N_15526,N_14486,N_14623);
xnor U15527 (N_15527,N_14394,N_13396);
nor U15528 (N_15528,N_13935,N_14347);
or U15529 (N_15529,N_14524,N_13062);
or U15530 (N_15530,N_14892,N_14017);
or U15531 (N_15531,N_14660,N_14544);
and U15532 (N_15532,N_13132,N_14170);
xnor U15533 (N_15533,N_13203,N_13697);
nand U15534 (N_15534,N_12621,N_14187);
xnor U15535 (N_15535,N_14259,N_12722);
nor U15536 (N_15536,N_12633,N_13283);
or U15537 (N_15537,N_13332,N_13756);
and U15538 (N_15538,N_12875,N_14650);
and U15539 (N_15539,N_13790,N_12892);
or U15540 (N_15540,N_13898,N_14405);
nand U15541 (N_15541,N_13929,N_14570);
nand U15542 (N_15542,N_14958,N_14237);
nor U15543 (N_15543,N_14645,N_14591);
and U15544 (N_15544,N_13398,N_12654);
and U15545 (N_15545,N_13402,N_12964);
and U15546 (N_15546,N_14937,N_14238);
nor U15547 (N_15547,N_12810,N_13866);
and U15548 (N_15548,N_14847,N_13567);
nand U15549 (N_15549,N_14396,N_13196);
nor U15550 (N_15550,N_14880,N_14694);
and U15551 (N_15551,N_13401,N_12861);
or U15552 (N_15552,N_14932,N_14565);
and U15553 (N_15553,N_14882,N_14835);
nand U15554 (N_15554,N_14672,N_13770);
nand U15555 (N_15555,N_14782,N_13123);
and U15556 (N_15556,N_14241,N_14790);
or U15557 (N_15557,N_14470,N_12986);
nor U15558 (N_15558,N_14617,N_14067);
xnor U15559 (N_15559,N_13207,N_13645);
nand U15560 (N_15560,N_14437,N_13609);
or U15561 (N_15561,N_13367,N_14784);
and U15562 (N_15562,N_14647,N_13071);
xnor U15563 (N_15563,N_14372,N_13705);
nor U15564 (N_15564,N_13257,N_14643);
nor U15565 (N_15565,N_12728,N_14424);
or U15566 (N_15566,N_14941,N_13646);
nand U15567 (N_15567,N_13024,N_13631);
nand U15568 (N_15568,N_12708,N_14412);
nor U15569 (N_15569,N_13669,N_13772);
and U15570 (N_15570,N_14626,N_13612);
nor U15571 (N_15571,N_14463,N_14102);
and U15572 (N_15572,N_14420,N_12907);
and U15573 (N_15573,N_12764,N_13829);
nand U15574 (N_15574,N_14716,N_13101);
nand U15575 (N_15575,N_14126,N_13986);
nand U15576 (N_15576,N_12972,N_13069);
nand U15577 (N_15577,N_14461,N_13867);
nor U15578 (N_15578,N_14349,N_14504);
xnor U15579 (N_15579,N_13822,N_12523);
xnor U15580 (N_15580,N_14684,N_14914);
and U15581 (N_15581,N_14150,N_14946);
nor U15582 (N_15582,N_14680,N_12790);
nand U15583 (N_15583,N_14333,N_13471);
xor U15584 (N_15584,N_12732,N_12626);
xnor U15585 (N_15585,N_12620,N_14356);
nand U15586 (N_15586,N_14350,N_14605);
nor U15587 (N_15587,N_14753,N_13938);
and U15588 (N_15588,N_14179,N_12637);
or U15589 (N_15589,N_14317,N_12871);
or U15590 (N_15590,N_14595,N_14030);
and U15591 (N_15591,N_14834,N_14113);
nand U15592 (N_15592,N_14928,N_12520);
or U15593 (N_15593,N_14936,N_13019);
or U15594 (N_15594,N_12773,N_14744);
nor U15595 (N_15595,N_13878,N_14522);
or U15596 (N_15596,N_14739,N_13991);
nand U15597 (N_15597,N_13088,N_13673);
nand U15598 (N_15598,N_13556,N_14803);
nand U15599 (N_15599,N_12750,N_13859);
and U15600 (N_15600,N_14710,N_13659);
and U15601 (N_15601,N_13682,N_14870);
nor U15602 (N_15602,N_13128,N_14659);
and U15603 (N_15603,N_13177,N_13061);
xnor U15604 (N_15604,N_14780,N_12835);
xnor U15605 (N_15605,N_14618,N_13300);
nor U15606 (N_15606,N_13774,N_14263);
nand U15607 (N_15607,N_12655,N_13224);
xor U15608 (N_15608,N_12792,N_13831);
and U15609 (N_15609,N_13723,N_13795);
nand U15610 (N_15610,N_13230,N_12979);
nor U15611 (N_15611,N_12539,N_14277);
nand U15612 (N_15612,N_12615,N_14619);
nor U15613 (N_15613,N_13292,N_13979);
xor U15614 (N_15614,N_12547,N_14905);
nor U15615 (N_15615,N_14146,N_14387);
or U15616 (N_15616,N_12966,N_13957);
nand U15617 (N_15617,N_14575,N_13921);
or U15618 (N_15618,N_12560,N_13564);
nor U15619 (N_15619,N_12581,N_14611);
nor U15620 (N_15620,N_13495,N_14364);
xnor U15621 (N_15621,N_14809,N_14995);
and U15622 (N_15622,N_12770,N_13915);
nor U15623 (N_15623,N_14960,N_14001);
nor U15624 (N_15624,N_13993,N_14788);
xor U15625 (N_15625,N_13939,N_13792);
nand U15626 (N_15626,N_14632,N_14325);
and U15627 (N_15627,N_13151,N_13870);
and U15628 (N_15628,N_14785,N_14566);
or U15629 (N_15629,N_14228,N_12667);
nor U15630 (N_15630,N_14955,N_13107);
or U15631 (N_15631,N_12873,N_12723);
nand U15632 (N_15632,N_13355,N_14752);
xnor U15633 (N_15633,N_13305,N_14706);
or U15634 (N_15634,N_14117,N_12574);
nand U15635 (N_15635,N_13964,N_14921);
and U15636 (N_15636,N_13163,N_13611);
nand U15637 (N_15637,N_12811,N_12956);
nor U15638 (N_15638,N_13754,N_13034);
nand U15639 (N_15639,N_14041,N_13311);
nor U15640 (N_15640,N_13597,N_13246);
and U15641 (N_15641,N_14888,N_13530);
or U15642 (N_15642,N_14266,N_13079);
or U15643 (N_15643,N_14020,N_14852);
or U15644 (N_15644,N_13596,N_13111);
nand U15645 (N_15645,N_12602,N_14428);
and U15646 (N_15646,N_14954,N_13136);
xnor U15647 (N_15647,N_13233,N_13916);
nor U15648 (N_15648,N_14902,N_14005);
nand U15649 (N_15649,N_14056,N_13528);
and U15650 (N_15650,N_14062,N_12839);
nand U15651 (N_15651,N_13882,N_14026);
xnor U15652 (N_15652,N_14092,N_14074);
nor U15653 (N_15653,N_12781,N_13998);
and U15654 (N_15654,N_13423,N_14037);
and U15655 (N_15655,N_14590,N_14344);
nand U15656 (N_15656,N_12895,N_14884);
or U15657 (N_15657,N_12738,N_14994);
or U15658 (N_15658,N_12695,N_13526);
nand U15659 (N_15659,N_14099,N_14774);
or U15660 (N_15660,N_13155,N_12821);
nor U15661 (N_15661,N_14545,N_12914);
xor U15662 (N_15662,N_14637,N_12909);
nor U15663 (N_15663,N_13562,N_14925);
xnor U15664 (N_15664,N_14098,N_14600);
nand U15665 (N_15665,N_13485,N_14374);
xor U15666 (N_15666,N_13590,N_13853);
or U15667 (N_15667,N_12572,N_13342);
and U15668 (N_15668,N_13580,N_14168);
or U15669 (N_15669,N_14226,N_13814);
nand U15670 (N_15670,N_13987,N_14429);
nand U15671 (N_15671,N_14805,N_14897);
xor U15672 (N_15672,N_13718,N_13444);
or U15673 (N_15673,N_14304,N_13881);
nand U15674 (N_15674,N_13287,N_14558);
xor U15675 (N_15675,N_13801,N_12739);
and U15676 (N_15676,N_13074,N_14177);
and U15677 (N_15677,N_13302,N_12573);
and U15678 (N_15678,N_13338,N_14740);
xnor U15679 (N_15679,N_12903,N_14523);
or U15680 (N_15680,N_12870,N_14112);
nand U15681 (N_15681,N_13039,N_13663);
and U15682 (N_15682,N_14201,N_14625);
nor U15683 (N_15683,N_14161,N_14028);
nor U15684 (N_15684,N_14114,N_14319);
and U15685 (N_15685,N_13009,N_14213);
nand U15686 (N_15686,N_14786,N_13913);
nand U15687 (N_15687,N_14139,N_12604);
xnor U15688 (N_15688,N_14917,N_13897);
and U15689 (N_15689,N_14690,N_13383);
and U15690 (N_15690,N_13001,N_14864);
or U15691 (N_15691,N_13892,N_13212);
nand U15692 (N_15692,N_14576,N_13647);
nand U15693 (N_15693,N_14251,N_13717);
or U15694 (N_15694,N_14908,N_13895);
or U15695 (N_15695,N_13130,N_12993);
and U15696 (N_15696,N_13945,N_12591);
or U15697 (N_15697,N_14741,N_13885);
and U15698 (N_15698,N_14255,N_14230);
xor U15699 (N_15699,N_14879,N_14620);
or U15700 (N_15700,N_12513,N_14683);
or U15701 (N_15701,N_13037,N_14021);
xor U15702 (N_15702,N_13762,N_13753);
nor U15703 (N_15703,N_13280,N_12978);
nor U15704 (N_15704,N_14901,N_13960);
xor U15705 (N_15705,N_12940,N_14508);
and U15706 (N_15706,N_13318,N_13886);
and U15707 (N_15707,N_14453,N_13374);
or U15708 (N_15708,N_13780,N_13764);
nand U15709 (N_15709,N_14481,N_13028);
nor U15710 (N_15710,N_13610,N_14622);
xnor U15711 (N_15711,N_14166,N_14008);
nor U15712 (N_15712,N_13850,N_12753);
nand U15713 (N_15713,N_13797,N_14718);
and U15714 (N_15714,N_13857,N_13546);
and U15715 (N_15715,N_14129,N_13541);
or U15716 (N_15716,N_12931,N_13104);
or U15717 (N_15717,N_12859,N_13736);
and U15718 (N_15718,N_14324,N_12556);
nor U15719 (N_15719,N_13327,N_14980);
nor U15720 (N_15720,N_13010,N_14728);
nand U15721 (N_15721,N_14289,N_12877);
nor U15722 (N_15722,N_13763,N_14128);
or U15723 (N_15723,N_13511,N_13359);
nand U15724 (N_15724,N_14236,N_12608);
xor U15725 (N_15725,N_13432,N_13006);
or U15726 (N_15726,N_14843,N_13533);
and U15727 (N_15727,N_14060,N_13008);
or U15728 (N_15728,N_14160,N_14765);
nor U15729 (N_15729,N_12983,N_14838);
xor U15730 (N_15730,N_13439,N_13254);
xor U15731 (N_15731,N_14039,N_14764);
or U15732 (N_15732,N_13818,N_13808);
nand U15733 (N_15733,N_14214,N_12687);
or U15734 (N_15734,N_14415,N_14768);
nand U15735 (N_15735,N_13020,N_14351);
nor U15736 (N_15736,N_13066,N_14816);
or U15737 (N_15737,N_14883,N_14947);
and U15738 (N_15738,N_14252,N_14011);
nor U15739 (N_15739,N_13218,N_14313);
or U15740 (N_15740,N_14283,N_12641);
nor U15741 (N_15741,N_13264,N_13851);
nor U15742 (N_15742,N_14457,N_14903);
or U15743 (N_15743,N_13664,N_13827);
nor U15744 (N_15744,N_14178,N_12660);
and U15745 (N_15745,N_13005,N_14653);
or U15746 (N_15746,N_12817,N_13448);
xnor U15747 (N_15747,N_12713,N_12624);
nand U15748 (N_15748,N_12618,N_14106);
xor U15749 (N_15749,N_13761,N_12880);
nand U15750 (N_15750,N_13369,N_13570);
xor U15751 (N_15751,N_13537,N_13545);
or U15752 (N_15752,N_14518,N_13937);
or U15753 (N_15753,N_14671,N_12823);
nand U15754 (N_15754,N_14423,N_13145);
nor U15755 (N_15755,N_14144,N_14378);
nand U15756 (N_15756,N_13486,N_13927);
and U15757 (N_15757,N_13804,N_14970);
and U15758 (N_15758,N_14386,N_13942);
nand U15759 (N_15759,N_14119,N_13199);
xor U15760 (N_15760,N_14309,N_14326);
xnor U15761 (N_15761,N_14220,N_13309);
xor U15762 (N_15762,N_12825,N_13666);
nand U15763 (N_15763,N_13438,N_14288);
nor U15764 (N_15764,N_14354,N_13063);
and U15765 (N_15765,N_14053,N_14499);
and U15766 (N_15766,N_12652,N_13742);
nor U15767 (N_15767,N_14149,N_14548);
nand U15768 (N_15768,N_13809,N_13833);
nor U15769 (N_15769,N_14208,N_14059);
nand U15770 (N_15770,N_12593,N_13164);
xor U15771 (N_15771,N_14974,N_13340);
xor U15772 (N_15772,N_13158,N_14541);
or U15773 (N_15773,N_13720,N_12961);
xor U15774 (N_15774,N_13956,N_12856);
and U15775 (N_15775,N_14070,N_13504);
and U15776 (N_15776,N_13262,N_12975);
nor U15777 (N_15777,N_14235,N_13595);
or U15778 (N_15778,N_14705,N_13091);
xor U15779 (N_15779,N_14233,N_14959);
nand U15780 (N_15780,N_13525,N_12712);
xor U15781 (N_15781,N_14658,N_14748);
or U15782 (N_15782,N_13241,N_14163);
nand U15783 (N_15783,N_14939,N_14775);
nor U15784 (N_15784,N_12951,N_13589);
xor U15785 (N_15785,N_12843,N_13253);
nor U15786 (N_15786,N_13085,N_14493);
xnor U15787 (N_15787,N_12668,N_14182);
and U15788 (N_15788,N_12928,N_13324);
nor U15789 (N_15789,N_13425,N_14827);
nand U15790 (N_15790,N_13601,N_14963);
and U15791 (N_15791,N_12755,N_12919);
or U15792 (N_15792,N_13147,N_13096);
xor U15793 (N_15793,N_14517,N_14192);
nor U15794 (N_15794,N_13127,N_13568);
xor U15795 (N_15795,N_14081,N_14549);
xor U15796 (N_15796,N_12617,N_14095);
xor U15797 (N_15797,N_12852,N_14455);
nor U15798 (N_15798,N_14850,N_12996);
nor U15799 (N_15799,N_13807,N_13628);
nand U15800 (N_15800,N_14077,N_14860);
and U15801 (N_15801,N_14841,N_14991);
xor U15802 (N_15802,N_12930,N_13341);
and U15803 (N_15803,N_14957,N_13544);
nor U15804 (N_15804,N_13700,N_13947);
or U15805 (N_15805,N_14521,N_14435);
nor U15806 (N_15806,N_13094,N_14599);
nor U15807 (N_15807,N_14164,N_13296);
xor U15808 (N_15808,N_14806,N_12557);
nor U15809 (N_15809,N_14561,N_13784);
and U15810 (N_15810,N_12693,N_12664);
and U15811 (N_15811,N_14829,N_14815);
nor U15812 (N_15812,N_12564,N_14162);
or U15813 (N_15813,N_13662,N_13468);
xnor U15814 (N_15814,N_13965,N_13912);
or U15815 (N_15815,N_13457,N_14328);
nor U15816 (N_15816,N_14553,N_14385);
or U15817 (N_15817,N_13995,N_13574);
xnor U15818 (N_15818,N_13180,N_13052);
or U15819 (N_15819,N_12876,N_12552);
and U15820 (N_15820,N_13211,N_14881);
or U15821 (N_15821,N_14156,N_14582);
and U15822 (N_15822,N_14257,N_13161);
or U15823 (N_15823,N_13524,N_14015);
or U15824 (N_15824,N_13667,N_13289);
xnor U15825 (N_15825,N_14009,N_14557);
and U15826 (N_15826,N_14519,N_14502);
and U15827 (N_15827,N_12917,N_13497);
xor U15828 (N_15828,N_14746,N_12768);
and U15829 (N_15829,N_14920,N_12936);
and U15830 (N_15830,N_13279,N_13459);
nor U15831 (N_15831,N_13907,N_14043);
nor U15832 (N_15832,N_13274,N_14194);
xnor U15833 (N_15833,N_14440,N_13687);
nand U15834 (N_15834,N_13248,N_14794);
and U15835 (N_15835,N_14155,N_14400);
nor U15836 (N_15836,N_14465,N_13606);
nand U15837 (N_15837,N_12791,N_14276);
and U15838 (N_15838,N_14391,N_13520);
and U15839 (N_15839,N_14270,N_14363);
nor U15840 (N_15840,N_13724,N_13501);
and U15841 (N_15841,N_13558,N_13798);
or U15842 (N_15842,N_12526,N_14207);
nor U15843 (N_15843,N_12623,N_14629);
and U15844 (N_15844,N_12657,N_14628);
and U15845 (N_15845,N_14875,N_13531);
xnor U15846 (N_15846,N_14842,N_13277);
xnor U15847 (N_15847,N_14966,N_12959);
nor U15848 (N_15848,N_13250,N_13855);
or U15849 (N_15849,N_12897,N_13984);
and U15850 (N_15850,N_12551,N_13050);
nor U15851 (N_15851,N_13871,N_13583);
xnor U15852 (N_15852,N_14068,N_13793);
or U15853 (N_15853,N_13767,N_13845);
or U15854 (N_15854,N_13188,N_14615);
and U15855 (N_15855,N_12868,N_14051);
or U15856 (N_15856,N_14536,N_14406);
and U15857 (N_15857,N_13329,N_14798);
or U15858 (N_15858,N_14093,N_14886);
or U15859 (N_15859,N_14890,N_13377);
or U15860 (N_15860,N_13407,N_14246);
or U15861 (N_15861,N_14915,N_12998);
and U15862 (N_15862,N_14258,N_14169);
xnor U15863 (N_15863,N_14279,N_14022);
xor U15864 (N_15864,N_14079,N_13498);
nor U15865 (N_15865,N_13943,N_14534);
and U15866 (N_15866,N_14121,N_14825);
xnor U15867 (N_15867,N_14301,N_13553);
and U15868 (N_15868,N_14503,N_12950);
nand U15869 (N_15869,N_14857,N_12995);
nand U15870 (N_15870,N_13852,N_14948);
or U15871 (N_15871,N_13759,N_13182);
nor U15872 (N_15872,N_13811,N_13335);
or U15873 (N_15873,N_13632,N_12935);
xnor U15874 (N_15874,N_13953,N_13236);
or U15875 (N_15875,N_12688,N_14382);
nor U15876 (N_15876,N_13235,N_14256);
and U15877 (N_15877,N_14181,N_12796);
and U15878 (N_15878,N_13430,N_13242);
xnor U15879 (N_15879,N_12517,N_14292);
and U15880 (N_15880,N_13635,N_13256);
or U15881 (N_15881,N_14340,N_14550);
and U15882 (N_15882,N_12889,N_13086);
or U15883 (N_15883,N_12943,N_13624);
nand U15884 (N_15884,N_13787,N_13891);
or U15885 (N_15885,N_13899,N_13067);
nand U15886 (N_15886,N_13812,N_13676);
and U15887 (N_15887,N_12946,N_14714);
nand U15888 (N_15888,N_13688,N_12646);
xor U15889 (N_15889,N_14737,N_13112);
nand U15890 (N_15890,N_14813,N_13630);
and U15891 (N_15891,N_13382,N_13708);
nand U15892 (N_15892,N_12559,N_12900);
xor U15893 (N_15893,N_12818,N_14817);
xor U15894 (N_15894,N_13269,N_14501);
and U15895 (N_15895,N_14063,N_13141);
or U15896 (N_15896,N_14262,N_14322);
xor U15897 (N_15897,N_14801,N_13996);
and U15898 (N_15898,N_14988,N_13509);
nor U15899 (N_15899,N_13060,N_14416);
xnor U15900 (N_15900,N_14484,N_13339);
nor U15901 (N_15901,N_12534,N_12771);
and U15902 (N_15902,N_14648,N_14274);
and U15903 (N_15903,N_13862,N_12896);
xnor U15904 (N_15904,N_13213,N_12570);
and U15905 (N_15905,N_14212,N_14052);
or U15906 (N_15906,N_12830,N_14327);
xor U15907 (N_15907,N_13475,N_14472);
nand U15908 (N_15908,N_13554,N_14730);
or U15909 (N_15909,N_12879,N_13691);
xnor U15910 (N_15910,N_14792,N_13220);
nand U15911 (N_15911,N_12614,N_14642);
xnor U15912 (N_15912,N_13310,N_13514);
nor U15913 (N_15913,N_14649,N_13175);
or U15914 (N_15914,N_14107,N_14766);
nor U15915 (N_15915,N_13625,N_12529);
xor U15916 (N_15916,N_14824,N_12749);
xor U15917 (N_15917,N_13989,N_14754);
nor U15918 (N_15918,N_14338,N_12511);
or U15919 (N_15919,N_14245,N_14853);
nand U15920 (N_15920,N_14307,N_13731);
nand U15921 (N_15921,N_14339,N_14634);
or U15922 (N_15922,N_13931,N_13983);
and U15923 (N_15923,N_13198,N_13909);
nor U15924 (N_15924,N_14321,N_12681);
nor U15925 (N_15925,N_13963,N_12677);
nor U15926 (N_15926,N_13326,N_13121);
xnor U15927 (N_15927,N_13464,N_13729);
nand U15928 (N_15928,N_13615,N_13834);
or U15929 (N_15929,N_14964,N_13173);
or U15930 (N_15930,N_13607,N_13214);
or U15931 (N_15931,N_14874,N_12906);
nand U15932 (N_15932,N_12828,N_13358);
nor U15933 (N_15933,N_14397,N_13707);
or U15934 (N_15934,N_12847,N_14674);
nor U15935 (N_15935,N_12625,N_14007);
or U15936 (N_15936,N_13328,N_12619);
nand U15937 (N_15937,N_14188,N_13153);
or U15938 (N_15938,N_13424,N_12730);
nand U15939 (N_15939,N_13361,N_12554);
xor U15940 (N_15940,N_14999,N_13782);
nand U15941 (N_15941,N_14249,N_14225);
and U15942 (N_15942,N_12653,N_13148);
and U15943 (N_15943,N_14831,N_13906);
nor U15944 (N_15944,N_13138,N_14556);
xnor U15945 (N_15945,N_13600,N_13223);
xor U15946 (N_15946,N_13417,N_12838);
or U15947 (N_15947,N_14863,N_13375);
nand U15948 (N_15948,N_13651,N_12795);
xor U15949 (N_15949,N_13380,N_14185);
xor U15950 (N_15950,N_14004,N_13453);
or U15951 (N_15951,N_14312,N_14332);
and U15952 (N_15952,N_14703,N_12987);
or U15953 (N_15953,N_13142,N_14840);
nor U15954 (N_15954,N_14460,N_12662);
nor U15955 (N_15955,N_14800,N_14862);
or U15956 (N_15956,N_14389,N_14926);
xnor U15957 (N_15957,N_14086,N_12988);
nand U15958 (N_15958,N_13512,N_14240);
and U15959 (N_15959,N_14729,N_14345);
nor U15960 (N_15960,N_13971,N_12806);
and U15961 (N_15961,N_13652,N_13712);
and U15962 (N_15962,N_13877,N_12532);
xnor U15963 (N_15963,N_13999,N_14712);
xnor U15964 (N_15964,N_13362,N_14152);
or U15965 (N_15965,N_13208,N_13388);
xor U15966 (N_15966,N_13677,N_13278);
nand U15967 (N_15967,N_12855,N_14596);
nand U15968 (N_15968,N_12578,N_14528);
xor U15969 (N_15969,N_14254,N_13240);
and U15970 (N_15970,N_13637,N_14630);
nand U15971 (N_15971,N_13251,N_13582);
nand U15972 (N_15972,N_12845,N_13746);
nand U15973 (N_15973,N_14050,N_13144);
xor U15974 (N_15974,N_14573,N_13347);
xor U15975 (N_15975,N_14445,N_14563);
xnor U15976 (N_15976,N_13923,N_12558);
and U15977 (N_15977,N_13270,N_14949);
and U15978 (N_15978,N_12669,N_14449);
nand U15979 (N_15979,N_12643,N_13621);
nand U15980 (N_15980,N_12866,N_14090);
and U15981 (N_15981,N_13317,N_12555);
or U15982 (N_15982,N_13356,N_12524);
and U15983 (N_15983,N_12647,N_14804);
nand U15984 (N_15984,N_12862,N_12577);
or U15985 (N_15985,N_14935,N_14454);
nand U15986 (N_15986,N_12968,N_13803);
nand U15987 (N_15987,N_12848,N_13166);
and U15988 (N_15988,N_14568,N_13462);
or U15989 (N_15989,N_13949,N_14761);
or U15990 (N_15990,N_14284,N_14239);
nand U15991 (N_15991,N_13408,N_13944);
nor U15992 (N_15992,N_14369,N_12592);
xnor U15993 (N_15993,N_14743,N_12850);
or U15994 (N_15994,N_12566,N_13379);
xnor U15995 (N_15995,N_12734,N_12803);
nor U15996 (N_15996,N_14362,N_12754);
nor U15997 (N_15997,N_13133,N_14593);
xor U15998 (N_15998,N_14247,N_13757);
nor U15999 (N_15999,N_14124,N_13539);
and U16000 (N_16000,N_13540,N_14742);
or U16001 (N_16001,N_13918,N_13385);
xnor U16002 (N_16002,N_13840,N_13670);
nor U16003 (N_16003,N_14480,N_12711);
nor U16004 (N_16004,N_12942,N_12782);
nor U16005 (N_16005,N_12819,N_13560);
or U16006 (N_16006,N_14535,N_14330);
nand U16007 (N_16007,N_13353,N_13824);
nor U16008 (N_16008,N_14489,N_13933);
xnor U16009 (N_16009,N_14336,N_12548);
and U16010 (N_16010,N_13187,N_14248);
nor U16011 (N_16011,N_14933,N_14762);
and U16012 (N_16012,N_14495,N_13049);
or U16013 (N_16013,N_14355,N_12804);
xor U16014 (N_16014,N_13967,N_12675);
and U16015 (N_16015,N_12644,N_12586);
and U16016 (N_16016,N_14579,N_13105);
nand U16017 (N_16017,N_14118,N_13249);
xnor U16018 (N_16018,N_14165,N_12921);
nand U16019 (N_16019,N_14736,N_13848);
nand U16020 (N_16020,N_14749,N_13201);
nand U16021 (N_16021,N_14466,N_12567);
and U16022 (N_16022,N_13360,N_14584);
or U16023 (N_16023,N_12937,N_14986);
xnor U16024 (N_16024,N_12867,N_12922);
xnor U16025 (N_16025,N_13259,N_12974);
xnor U16026 (N_16026,N_14977,N_13349);
or U16027 (N_16027,N_12916,N_14664);
nand U16028 (N_16028,N_12680,N_13716);
nor U16029 (N_16029,N_13129,N_13903);
xor U16030 (N_16030,N_13027,N_12854);
nand U16031 (N_16031,N_13422,N_14976);
nand U16032 (N_16032,N_13469,N_13183);
xnor U16033 (N_16033,N_13186,N_13940);
and U16034 (N_16034,N_13969,N_14640);
and U16035 (N_16035,N_12969,N_13303);
xnor U16036 (N_16036,N_12751,N_12594);
and U16037 (N_16037,N_14985,N_13715);
xor U16038 (N_16038,N_14368,N_14560);
or U16039 (N_16039,N_13894,N_12719);
nand U16040 (N_16040,N_14930,N_13334);
or U16041 (N_16041,N_13506,N_12864);
xor U16042 (N_16042,N_13816,N_12648);
xnor U16043 (N_16043,N_13838,N_13616);
nand U16044 (N_16044,N_14488,N_13030);
xnor U16045 (N_16045,N_14075,N_12807);
or U16046 (N_16046,N_14656,N_13014);
nor U16047 (N_16047,N_14014,N_12502);
or U16048 (N_16048,N_12715,N_14540);
and U16049 (N_16049,N_13371,N_12516);
nor U16050 (N_16050,N_12887,N_13195);
nor U16051 (N_16051,N_13267,N_13786);
nand U16052 (N_16052,N_13656,N_13466);
nand U16053 (N_16053,N_12923,N_14639);
xor U16054 (N_16054,N_14777,N_12853);
nor U16055 (N_16055,N_12575,N_14635);
nand U16056 (N_16056,N_14418,N_13674);
or U16057 (N_16057,N_14998,N_12705);
nand U16058 (N_16058,N_13119,N_13135);
nand U16059 (N_16059,N_13489,N_13581);
or U16060 (N_16060,N_14154,N_12533);
nor U16061 (N_16061,N_12960,N_12597);
and U16062 (N_16062,N_14353,N_13791);
or U16063 (N_16063,N_13522,N_13064);
and U16064 (N_16064,N_14865,N_14109);
or U16065 (N_16065,N_12726,N_13070);
nand U16066 (N_16066,N_12743,N_13640);
nor U16067 (N_16067,N_14105,N_12530);
xor U16068 (N_16068,N_12582,N_12630);
xor U16069 (N_16069,N_12689,N_13565);
or U16070 (N_16070,N_14609,N_12616);
and U16071 (N_16071,N_14585,N_12733);
xnor U16072 (N_16072,N_12778,N_12826);
or U16073 (N_16073,N_14735,N_14845);
nor U16074 (N_16074,N_13089,N_13298);
and U16075 (N_16075,N_13463,N_14750);
and U16076 (N_16076,N_13730,N_14651);
xnor U16077 (N_16077,N_13075,N_13680);
nand U16078 (N_16078,N_13699,N_13966);
xnor U16079 (N_16079,N_13314,N_13926);
and U16080 (N_16080,N_12934,N_14898);
or U16081 (N_16081,N_13108,N_14727);
nor U16082 (N_16082,N_14491,N_12702);
and U16083 (N_16083,N_13271,N_13387);
and U16084 (N_16084,N_14229,N_13093);
nor U16085 (N_16085,N_13962,N_14085);
nor U16086 (N_16086,N_14171,N_14433);
or U16087 (N_16087,N_14854,N_12745);
nand U16088 (N_16088,N_14496,N_14498);
nor U16089 (N_16089,N_13773,N_13330);
xor U16090 (N_16090,N_13839,N_14273);
xor U16091 (N_16091,N_12812,N_13053);
or U16092 (N_16092,N_14032,N_14450);
nand U16093 (N_16093,N_13449,N_13598);
nand U16094 (N_16094,N_12766,N_14190);
xor U16095 (N_16095,N_14040,N_14877);
nor U16096 (N_16096,N_14973,N_14477);
and U16097 (N_16097,N_14514,N_12661);
nor U16098 (N_16098,N_13460,N_14485);
xnor U16099 (N_16099,N_12735,N_14367);
or U16100 (N_16100,N_12953,N_13357);
or U16101 (N_16101,N_12981,N_14446);
or U16102 (N_16102,N_14666,N_13686);
and U16103 (N_16103,N_14018,N_13391);
nor U16104 (N_16104,N_12512,N_14698);
or U16105 (N_16105,N_14447,N_14127);
nand U16106 (N_16106,N_13076,N_13634);
nand U16107 (N_16107,N_13988,N_12519);
and U16108 (N_16108,N_12789,N_13849);
and U16109 (N_16109,N_13068,N_14723);
nor U16110 (N_16110,N_12510,N_12836);
nor U16111 (N_16111,N_13484,N_14250);
nor U16112 (N_16112,N_13714,N_12704);
nor U16113 (N_16113,N_13363,N_13445);
nand U16114 (N_16114,N_14172,N_14487);
xnor U16115 (N_16115,N_13454,N_12794);
nand U16116 (N_16116,N_13204,N_12721);
and U16117 (N_16117,N_13602,N_14969);
nand U16118 (N_16118,N_14687,N_14024);
nand U16119 (N_16119,N_13711,N_14003);
xor U16120 (N_16120,N_13299,N_13210);
or U16121 (N_16121,N_12587,N_12636);
nand U16122 (N_16122,N_13893,N_12967);
nor U16123 (N_16123,N_14978,N_14380);
and U16124 (N_16124,N_13547,N_14776);
nor U16125 (N_16125,N_14669,N_13333);
xor U16126 (N_16126,N_13860,N_13483);
xor U16127 (N_16127,N_14602,N_14624);
or U16128 (N_16128,N_14636,N_14856);
and U16129 (N_16129,N_13389,N_14719);
xnor U16130 (N_16130,N_13917,N_13103);
nand U16131 (N_16131,N_13658,N_12725);
xor U16132 (N_16132,N_13167,N_13559);
xnor U16133 (N_16133,N_14830,N_13861);
and U16134 (N_16134,N_14296,N_14471);
nor U16135 (N_16135,N_14298,N_13150);
nand U16136 (N_16136,N_13551,N_12997);
and U16137 (N_16137,N_13654,N_13042);
or U16138 (N_16138,N_13386,N_12762);
or U16139 (N_16139,N_14644,N_12929);
nand U16140 (N_16140,N_14294,N_14763);
nand U16141 (N_16141,N_13910,N_14731);
and U16142 (N_16142,N_12686,N_14482);
nand U16143 (N_16143,N_13709,N_14371);
xnor U16144 (N_16144,N_13863,N_14242);
nor U16145 (N_16145,N_13925,N_13710);
and U16146 (N_16146,N_12583,N_12924);
and U16147 (N_16147,N_13319,N_12645);
xnor U16148 (N_16148,N_14260,N_13205);
nand U16149 (N_16149,N_14411,N_14953);
xnor U16150 (N_16150,N_12598,N_12638);
or U16151 (N_16151,N_14951,N_13739);
and U16152 (N_16152,N_13045,N_13365);
nor U16153 (N_16153,N_14196,N_13517);
nor U16154 (N_16154,N_14525,N_13140);
nand U16155 (N_16155,N_12941,N_14054);
nand U16156 (N_16156,N_14303,N_14209);
or U16157 (N_16157,N_12599,N_14438);
nor U16158 (N_16158,N_13683,N_13561);
or U16159 (N_16159,N_14833,N_14555);
xor U16160 (N_16160,N_14227,N_14989);
and U16161 (N_16161,N_12748,N_13479);
nor U16162 (N_16162,N_12918,N_13599);
nor U16163 (N_16163,N_14280,N_12908);
or U16164 (N_16164,N_13343,N_14299);
nand U16165 (N_16165,N_13301,N_13227);
nor U16166 (N_16166,N_14899,N_14614);
xor U16167 (N_16167,N_14002,N_14490);
xnor U16168 (N_16168,N_13618,N_13162);
and U16169 (N_16169,N_12925,N_14646);
xnor U16170 (N_16170,N_14033,N_12528);
nand U16171 (N_16171,N_13315,N_13858);
xnor U16172 (N_16172,N_13876,N_13588);
xor U16173 (N_16173,N_14343,N_12672);
or U16174 (N_16174,N_13794,N_13110);
nor U16175 (N_16175,N_14577,N_13976);
or U16176 (N_16176,N_14696,N_14707);
nand U16177 (N_16177,N_13083,N_13788);
xnor U16178 (N_16178,N_13304,N_14627);
nor U16179 (N_16179,N_14984,N_14083);
or U16180 (N_16180,N_14108,N_13847);
nor U16181 (N_16181,N_14290,N_12741);
nor U16182 (N_16182,N_14516,N_14422);
nand U16183 (N_16183,N_12801,N_13875);
xnor U16184 (N_16184,N_14848,N_14441);
or U16185 (N_16185,N_14287,N_13650);
nand U16186 (N_16186,N_14034,N_13331);
nor U16187 (N_16187,N_13980,N_14996);
or U16188 (N_16188,N_13642,N_13657);
nand U16189 (N_16189,N_14793,N_13165);
nand U16190 (N_16190,N_12947,N_14961);
and U16191 (N_16191,N_13036,N_13415);
and U16192 (N_16192,N_13954,N_13887);
nand U16193 (N_16193,N_12888,N_13778);
xor U16194 (N_16194,N_14802,N_13813);
and U16195 (N_16195,N_12628,N_12948);
nor U16196 (N_16196,N_13116,N_12632);
and U16197 (N_16197,N_14265,N_13055);
and U16198 (N_16198,N_13106,N_13970);
and U16199 (N_16199,N_12849,N_13095);
xnor U16200 (N_16200,N_13344,N_13176);
and U16201 (N_16201,N_12642,N_12822);
nor U16202 (N_16202,N_13743,N_13041);
xor U16203 (N_16203,N_13322,N_14202);
nand U16204 (N_16204,N_13817,N_12538);
and U16205 (N_16205,N_14348,N_13451);
nand U16206 (N_16206,N_13057,N_13437);
and U16207 (N_16207,N_14331,N_14359);
and U16208 (N_16208,N_13557,N_14871);
nor U16209 (N_16209,N_14779,N_14130);
and U16210 (N_16210,N_13614,N_13126);
nand U16211 (N_16211,N_14572,N_14911);
nand U16212 (N_16212,N_12911,N_13431);
nand U16213 (N_16213,N_14311,N_14526);
xor U16214 (N_16214,N_13825,N_14358);
nor U16215 (N_16215,N_12842,N_13100);
nand U16216 (N_16216,N_13924,N_12905);
xnor U16217 (N_16217,N_13491,N_13139);
xnor U16218 (N_16218,N_14956,N_13902);
xor U16219 (N_16219,N_14210,N_13048);
xnor U16220 (N_16220,N_13507,N_14667);
or U16221 (N_16221,N_14271,N_14530);
or U16222 (N_16222,N_14796,N_13440);
or U16223 (N_16223,N_14198,N_12568);
or U16224 (N_16224,N_14469,N_13563);
nand U16225 (N_16225,N_14581,N_14479);
or U16226 (N_16226,N_14352,N_13202);
and U16227 (N_16227,N_14588,N_14868);
xor U16228 (N_16228,N_12954,N_13476);
nand U16229 (N_16229,N_12874,N_13571);
and U16230 (N_16230,N_13796,N_12656);
nand U16231 (N_16231,N_13346,N_14662);
and U16232 (N_16232,N_13732,N_13393);
nor U16233 (N_16233,N_14357,N_13081);
and U16234 (N_16234,N_13461,N_14029);
xnor U16235 (N_16235,N_12611,N_14734);
xor U16236 (N_16236,N_14676,N_13276);
and U16237 (N_16237,N_13815,N_12612);
or U16238 (N_16238,N_14205,N_12999);
and U16239 (N_16239,N_13225,N_13579);
and U16240 (N_16240,N_14967,N_13261);
and U16241 (N_16241,N_12684,N_13472);
nor U16242 (N_16242,N_13238,N_13776);
xnor U16243 (N_16243,N_14084,N_13837);
and U16244 (N_16244,N_14361,N_13419);
and U16245 (N_16245,N_13397,N_14143);
and U16246 (N_16246,N_14708,N_12666);
nor U16247 (N_16247,N_14055,N_13685);
nand U16248 (N_16248,N_12605,N_13493);
and U16249 (N_16249,N_13638,N_14665);
and U16250 (N_16250,N_14491,N_13808);
nand U16251 (N_16251,N_14767,N_14061);
and U16252 (N_16252,N_13471,N_13535);
nor U16253 (N_16253,N_14424,N_14759);
or U16254 (N_16254,N_14642,N_12805);
and U16255 (N_16255,N_14280,N_12640);
and U16256 (N_16256,N_13657,N_14780);
nand U16257 (N_16257,N_13832,N_13560);
nand U16258 (N_16258,N_14296,N_13669);
and U16259 (N_16259,N_13961,N_13734);
or U16260 (N_16260,N_13613,N_13143);
and U16261 (N_16261,N_14762,N_12979);
nor U16262 (N_16262,N_13461,N_13293);
nand U16263 (N_16263,N_14089,N_13127);
nor U16264 (N_16264,N_13461,N_13757);
xor U16265 (N_16265,N_14519,N_13821);
nand U16266 (N_16266,N_13101,N_14011);
nand U16267 (N_16267,N_14492,N_13308);
or U16268 (N_16268,N_13369,N_14014);
nand U16269 (N_16269,N_13230,N_14045);
nand U16270 (N_16270,N_12712,N_14194);
nor U16271 (N_16271,N_14002,N_14766);
nor U16272 (N_16272,N_12804,N_14264);
xnor U16273 (N_16273,N_13808,N_13415);
nor U16274 (N_16274,N_13331,N_13183);
xor U16275 (N_16275,N_14868,N_12558);
nor U16276 (N_16276,N_14344,N_14606);
xor U16277 (N_16277,N_12861,N_14571);
nor U16278 (N_16278,N_14572,N_13463);
or U16279 (N_16279,N_14959,N_13598);
nand U16280 (N_16280,N_13221,N_12566);
xnor U16281 (N_16281,N_14074,N_14099);
nand U16282 (N_16282,N_13361,N_14331);
and U16283 (N_16283,N_12742,N_14893);
nand U16284 (N_16284,N_14137,N_13668);
xor U16285 (N_16285,N_13232,N_13535);
or U16286 (N_16286,N_14833,N_12525);
xnor U16287 (N_16287,N_12986,N_12901);
nor U16288 (N_16288,N_12890,N_14820);
and U16289 (N_16289,N_14723,N_13597);
and U16290 (N_16290,N_13438,N_13873);
nand U16291 (N_16291,N_14188,N_13326);
nor U16292 (N_16292,N_12914,N_13561);
nor U16293 (N_16293,N_14629,N_14719);
xor U16294 (N_16294,N_14079,N_12895);
and U16295 (N_16295,N_14017,N_13093);
nor U16296 (N_16296,N_13897,N_13092);
nand U16297 (N_16297,N_12872,N_14331);
and U16298 (N_16298,N_12963,N_12611);
xor U16299 (N_16299,N_13225,N_14644);
nand U16300 (N_16300,N_14373,N_12941);
or U16301 (N_16301,N_14824,N_13040);
or U16302 (N_16302,N_14539,N_13114);
xnor U16303 (N_16303,N_13387,N_14373);
and U16304 (N_16304,N_12930,N_13974);
nand U16305 (N_16305,N_14200,N_13473);
and U16306 (N_16306,N_14950,N_14829);
and U16307 (N_16307,N_12514,N_12572);
xnor U16308 (N_16308,N_14802,N_14828);
xor U16309 (N_16309,N_14914,N_14121);
and U16310 (N_16310,N_13904,N_12534);
or U16311 (N_16311,N_13429,N_14105);
and U16312 (N_16312,N_13986,N_13938);
and U16313 (N_16313,N_12965,N_14970);
or U16314 (N_16314,N_14544,N_14060);
nand U16315 (N_16315,N_13408,N_13048);
nand U16316 (N_16316,N_13849,N_13386);
nor U16317 (N_16317,N_13681,N_14909);
or U16318 (N_16318,N_14100,N_14824);
nand U16319 (N_16319,N_13843,N_13062);
and U16320 (N_16320,N_13912,N_14875);
or U16321 (N_16321,N_14596,N_14184);
nor U16322 (N_16322,N_14920,N_14702);
and U16323 (N_16323,N_13411,N_13094);
xnor U16324 (N_16324,N_12767,N_13818);
and U16325 (N_16325,N_14431,N_14293);
xnor U16326 (N_16326,N_12997,N_12910);
nand U16327 (N_16327,N_12833,N_13334);
and U16328 (N_16328,N_13986,N_12986);
and U16329 (N_16329,N_13629,N_13446);
or U16330 (N_16330,N_13189,N_14297);
nor U16331 (N_16331,N_12953,N_14195);
and U16332 (N_16332,N_14539,N_13073);
and U16333 (N_16333,N_13184,N_13529);
xnor U16334 (N_16334,N_13821,N_13565);
nand U16335 (N_16335,N_14659,N_13946);
nor U16336 (N_16336,N_14110,N_12600);
nand U16337 (N_16337,N_13182,N_13385);
or U16338 (N_16338,N_14670,N_12847);
xnor U16339 (N_16339,N_12845,N_13315);
and U16340 (N_16340,N_14827,N_12614);
nor U16341 (N_16341,N_12881,N_13855);
and U16342 (N_16342,N_13246,N_14354);
nand U16343 (N_16343,N_12958,N_14257);
xnor U16344 (N_16344,N_13851,N_14892);
xnor U16345 (N_16345,N_13871,N_13163);
and U16346 (N_16346,N_12886,N_14596);
nor U16347 (N_16347,N_14545,N_13124);
or U16348 (N_16348,N_13095,N_14925);
or U16349 (N_16349,N_12868,N_13042);
xor U16350 (N_16350,N_13174,N_13516);
xor U16351 (N_16351,N_12763,N_14623);
and U16352 (N_16352,N_13769,N_13272);
or U16353 (N_16353,N_13730,N_14275);
nor U16354 (N_16354,N_14652,N_13324);
and U16355 (N_16355,N_13177,N_13203);
xor U16356 (N_16356,N_14267,N_13082);
and U16357 (N_16357,N_14911,N_12521);
xnor U16358 (N_16358,N_14604,N_13821);
or U16359 (N_16359,N_12948,N_14429);
nor U16360 (N_16360,N_14689,N_14025);
or U16361 (N_16361,N_14066,N_13685);
nor U16362 (N_16362,N_14319,N_13532);
xor U16363 (N_16363,N_14719,N_13078);
nand U16364 (N_16364,N_14302,N_14663);
or U16365 (N_16365,N_14885,N_12816);
or U16366 (N_16366,N_14942,N_14264);
and U16367 (N_16367,N_14470,N_13138);
xor U16368 (N_16368,N_14205,N_14463);
or U16369 (N_16369,N_14622,N_13277);
nand U16370 (N_16370,N_12952,N_12682);
xor U16371 (N_16371,N_12577,N_12747);
or U16372 (N_16372,N_13609,N_12887);
and U16373 (N_16373,N_14422,N_12848);
and U16374 (N_16374,N_14644,N_12731);
or U16375 (N_16375,N_14697,N_13255);
and U16376 (N_16376,N_13749,N_14030);
or U16377 (N_16377,N_12823,N_12646);
and U16378 (N_16378,N_14269,N_13683);
nor U16379 (N_16379,N_14063,N_13912);
xnor U16380 (N_16380,N_12961,N_12829);
and U16381 (N_16381,N_13331,N_14487);
nand U16382 (N_16382,N_13266,N_14457);
and U16383 (N_16383,N_12863,N_13673);
and U16384 (N_16384,N_13035,N_12622);
nor U16385 (N_16385,N_13411,N_12853);
or U16386 (N_16386,N_14139,N_13814);
nand U16387 (N_16387,N_12796,N_13172);
or U16388 (N_16388,N_14267,N_13220);
and U16389 (N_16389,N_12947,N_14036);
and U16390 (N_16390,N_13763,N_14613);
or U16391 (N_16391,N_13013,N_13192);
nand U16392 (N_16392,N_14521,N_12606);
xnor U16393 (N_16393,N_13459,N_14846);
xnor U16394 (N_16394,N_12986,N_14878);
or U16395 (N_16395,N_14824,N_12600);
or U16396 (N_16396,N_13100,N_12545);
nor U16397 (N_16397,N_13945,N_14653);
nand U16398 (N_16398,N_13689,N_12610);
or U16399 (N_16399,N_14253,N_13541);
or U16400 (N_16400,N_14743,N_14635);
and U16401 (N_16401,N_14088,N_12737);
nor U16402 (N_16402,N_12823,N_14539);
and U16403 (N_16403,N_14037,N_14795);
nand U16404 (N_16404,N_13887,N_13102);
xnor U16405 (N_16405,N_13721,N_14808);
nand U16406 (N_16406,N_13978,N_13498);
nand U16407 (N_16407,N_13379,N_14597);
nor U16408 (N_16408,N_13567,N_12533);
or U16409 (N_16409,N_12939,N_13155);
and U16410 (N_16410,N_14096,N_14836);
xor U16411 (N_16411,N_13987,N_14920);
or U16412 (N_16412,N_13107,N_12847);
xnor U16413 (N_16413,N_14285,N_13694);
and U16414 (N_16414,N_14206,N_14188);
and U16415 (N_16415,N_14609,N_14215);
nand U16416 (N_16416,N_14320,N_13190);
nor U16417 (N_16417,N_13317,N_13573);
nor U16418 (N_16418,N_12888,N_14176);
xnor U16419 (N_16419,N_14770,N_13344);
or U16420 (N_16420,N_14118,N_13587);
xnor U16421 (N_16421,N_14270,N_13228);
nand U16422 (N_16422,N_12606,N_14736);
or U16423 (N_16423,N_13536,N_12507);
or U16424 (N_16424,N_12784,N_12884);
xor U16425 (N_16425,N_12800,N_13847);
or U16426 (N_16426,N_13858,N_13620);
and U16427 (N_16427,N_14589,N_14095);
and U16428 (N_16428,N_14292,N_14883);
nand U16429 (N_16429,N_13766,N_13987);
xnor U16430 (N_16430,N_13162,N_13041);
xnor U16431 (N_16431,N_14642,N_13679);
nand U16432 (N_16432,N_13552,N_13289);
xor U16433 (N_16433,N_14113,N_14614);
nand U16434 (N_16434,N_14175,N_12587);
or U16435 (N_16435,N_14657,N_13677);
nand U16436 (N_16436,N_12546,N_13278);
or U16437 (N_16437,N_14850,N_14836);
or U16438 (N_16438,N_12957,N_12868);
or U16439 (N_16439,N_13552,N_14092);
or U16440 (N_16440,N_14954,N_14799);
nor U16441 (N_16441,N_13923,N_14404);
or U16442 (N_16442,N_13388,N_14043);
and U16443 (N_16443,N_13738,N_14331);
or U16444 (N_16444,N_13075,N_14614);
and U16445 (N_16445,N_13704,N_12984);
nor U16446 (N_16446,N_13879,N_12872);
or U16447 (N_16447,N_12658,N_12929);
or U16448 (N_16448,N_12688,N_14560);
nand U16449 (N_16449,N_12650,N_14708);
nor U16450 (N_16450,N_13918,N_13044);
nand U16451 (N_16451,N_14602,N_14361);
nor U16452 (N_16452,N_13677,N_13140);
xnor U16453 (N_16453,N_14556,N_13908);
xor U16454 (N_16454,N_13319,N_12556);
xor U16455 (N_16455,N_14415,N_12718);
and U16456 (N_16456,N_12974,N_14944);
nor U16457 (N_16457,N_14363,N_12815);
or U16458 (N_16458,N_14308,N_14880);
nor U16459 (N_16459,N_13786,N_12580);
or U16460 (N_16460,N_12663,N_12751);
nor U16461 (N_16461,N_13663,N_14325);
nand U16462 (N_16462,N_14133,N_14843);
or U16463 (N_16463,N_12665,N_14399);
nand U16464 (N_16464,N_12942,N_14466);
nor U16465 (N_16465,N_13992,N_13237);
nand U16466 (N_16466,N_13664,N_14084);
and U16467 (N_16467,N_14724,N_14760);
or U16468 (N_16468,N_13697,N_14921);
nor U16469 (N_16469,N_13164,N_14852);
and U16470 (N_16470,N_13102,N_13343);
nand U16471 (N_16471,N_13692,N_13619);
nand U16472 (N_16472,N_12581,N_14694);
xor U16473 (N_16473,N_14230,N_14669);
or U16474 (N_16474,N_13993,N_14437);
nand U16475 (N_16475,N_14393,N_12802);
and U16476 (N_16476,N_13694,N_13572);
xnor U16477 (N_16477,N_12662,N_14120);
and U16478 (N_16478,N_12889,N_14051);
nand U16479 (N_16479,N_13224,N_14596);
xnor U16480 (N_16480,N_13534,N_13930);
xor U16481 (N_16481,N_14521,N_13268);
xnor U16482 (N_16482,N_13027,N_14229);
nand U16483 (N_16483,N_13071,N_14666);
nor U16484 (N_16484,N_14986,N_14171);
or U16485 (N_16485,N_14491,N_13358);
or U16486 (N_16486,N_14884,N_13634);
nor U16487 (N_16487,N_13393,N_12778);
and U16488 (N_16488,N_12953,N_12519);
or U16489 (N_16489,N_12964,N_12638);
xnor U16490 (N_16490,N_14445,N_13790);
nand U16491 (N_16491,N_14669,N_12582);
xor U16492 (N_16492,N_13183,N_14385);
xnor U16493 (N_16493,N_13095,N_13651);
or U16494 (N_16494,N_13053,N_14856);
nor U16495 (N_16495,N_14387,N_14800);
nand U16496 (N_16496,N_12759,N_14543);
or U16497 (N_16497,N_14630,N_14404);
nor U16498 (N_16498,N_14987,N_12731);
and U16499 (N_16499,N_13926,N_13927);
or U16500 (N_16500,N_14007,N_12586);
nor U16501 (N_16501,N_14047,N_14623);
and U16502 (N_16502,N_13604,N_14963);
xnor U16503 (N_16503,N_13661,N_13261);
and U16504 (N_16504,N_14786,N_14928);
nand U16505 (N_16505,N_14740,N_12928);
nand U16506 (N_16506,N_13616,N_13151);
nand U16507 (N_16507,N_13686,N_14109);
xnor U16508 (N_16508,N_14198,N_13663);
nand U16509 (N_16509,N_14175,N_13613);
and U16510 (N_16510,N_13743,N_14383);
xnor U16511 (N_16511,N_14265,N_14073);
or U16512 (N_16512,N_13169,N_13522);
nand U16513 (N_16513,N_14424,N_13665);
xor U16514 (N_16514,N_13712,N_14661);
nand U16515 (N_16515,N_13176,N_13997);
or U16516 (N_16516,N_14826,N_14929);
or U16517 (N_16517,N_13263,N_14194);
or U16518 (N_16518,N_13430,N_12957);
nand U16519 (N_16519,N_13427,N_13253);
nand U16520 (N_16520,N_13066,N_13626);
xnor U16521 (N_16521,N_12673,N_13269);
nand U16522 (N_16522,N_12730,N_13149);
xnor U16523 (N_16523,N_12849,N_13330);
or U16524 (N_16524,N_13852,N_14449);
nor U16525 (N_16525,N_13021,N_13547);
nand U16526 (N_16526,N_14755,N_13532);
or U16527 (N_16527,N_13526,N_12789);
or U16528 (N_16528,N_13879,N_14646);
nor U16529 (N_16529,N_13130,N_13325);
xnor U16530 (N_16530,N_14095,N_12828);
xnor U16531 (N_16531,N_14717,N_14327);
and U16532 (N_16532,N_13708,N_13350);
xor U16533 (N_16533,N_13759,N_14421);
and U16534 (N_16534,N_14684,N_13275);
and U16535 (N_16535,N_14333,N_13743);
xnor U16536 (N_16536,N_13806,N_14771);
and U16537 (N_16537,N_12970,N_13363);
nor U16538 (N_16538,N_14128,N_14985);
nor U16539 (N_16539,N_12936,N_13682);
and U16540 (N_16540,N_13035,N_14151);
and U16541 (N_16541,N_12587,N_14008);
or U16542 (N_16542,N_13556,N_12764);
and U16543 (N_16543,N_13959,N_14423);
xnor U16544 (N_16544,N_12909,N_14237);
or U16545 (N_16545,N_14321,N_13341);
nor U16546 (N_16546,N_13583,N_12584);
or U16547 (N_16547,N_14203,N_14501);
or U16548 (N_16548,N_13314,N_13752);
or U16549 (N_16549,N_12981,N_12597);
or U16550 (N_16550,N_13156,N_14778);
nor U16551 (N_16551,N_14584,N_13198);
and U16552 (N_16552,N_13775,N_14170);
and U16553 (N_16553,N_14654,N_13275);
xnor U16554 (N_16554,N_12947,N_12700);
and U16555 (N_16555,N_14190,N_13928);
xnor U16556 (N_16556,N_14248,N_13047);
xnor U16557 (N_16557,N_13834,N_14599);
nor U16558 (N_16558,N_14046,N_13588);
nor U16559 (N_16559,N_14360,N_14371);
or U16560 (N_16560,N_12755,N_14101);
xnor U16561 (N_16561,N_14801,N_12886);
xor U16562 (N_16562,N_14567,N_12820);
xor U16563 (N_16563,N_14720,N_13271);
xnor U16564 (N_16564,N_12623,N_13982);
xnor U16565 (N_16565,N_14514,N_13556);
and U16566 (N_16566,N_13752,N_14897);
xor U16567 (N_16567,N_13785,N_14341);
and U16568 (N_16568,N_13429,N_14803);
nor U16569 (N_16569,N_14430,N_12617);
nor U16570 (N_16570,N_13505,N_14118);
or U16571 (N_16571,N_13997,N_12780);
nand U16572 (N_16572,N_12639,N_14630);
or U16573 (N_16573,N_14316,N_13589);
and U16574 (N_16574,N_14565,N_14717);
and U16575 (N_16575,N_13486,N_14285);
nand U16576 (N_16576,N_14167,N_12810);
nor U16577 (N_16577,N_14857,N_12571);
nand U16578 (N_16578,N_14544,N_14715);
xor U16579 (N_16579,N_13513,N_13097);
and U16580 (N_16580,N_14671,N_13683);
nand U16581 (N_16581,N_14616,N_13165);
nor U16582 (N_16582,N_14260,N_12628);
nor U16583 (N_16583,N_14962,N_14995);
and U16584 (N_16584,N_13357,N_12957);
xor U16585 (N_16585,N_13794,N_14327);
and U16586 (N_16586,N_14985,N_12718);
and U16587 (N_16587,N_14996,N_13945);
xnor U16588 (N_16588,N_12935,N_12905);
or U16589 (N_16589,N_14783,N_14810);
xnor U16590 (N_16590,N_13997,N_13036);
nand U16591 (N_16591,N_14180,N_12911);
and U16592 (N_16592,N_14120,N_14200);
xor U16593 (N_16593,N_14601,N_14559);
xnor U16594 (N_16594,N_14900,N_13261);
xnor U16595 (N_16595,N_14900,N_13467);
nand U16596 (N_16596,N_14261,N_12718);
xor U16597 (N_16597,N_13077,N_14253);
nor U16598 (N_16598,N_14063,N_14465);
or U16599 (N_16599,N_13632,N_13413);
xnor U16600 (N_16600,N_13896,N_14931);
nand U16601 (N_16601,N_13479,N_13206);
xor U16602 (N_16602,N_13051,N_14598);
xnor U16603 (N_16603,N_12995,N_14232);
and U16604 (N_16604,N_14158,N_12892);
and U16605 (N_16605,N_13338,N_14140);
and U16606 (N_16606,N_14325,N_14317);
and U16607 (N_16607,N_12876,N_12694);
nand U16608 (N_16608,N_14847,N_14348);
xnor U16609 (N_16609,N_14969,N_12771);
or U16610 (N_16610,N_14194,N_14993);
nand U16611 (N_16611,N_13707,N_14412);
xor U16612 (N_16612,N_13081,N_13517);
or U16613 (N_16613,N_13624,N_14636);
or U16614 (N_16614,N_13209,N_13156);
xor U16615 (N_16615,N_12755,N_13851);
xnor U16616 (N_16616,N_13199,N_14278);
or U16617 (N_16617,N_12600,N_13988);
or U16618 (N_16618,N_12523,N_12526);
and U16619 (N_16619,N_13862,N_14535);
nor U16620 (N_16620,N_13061,N_13564);
and U16621 (N_16621,N_14977,N_14149);
nor U16622 (N_16622,N_13039,N_12694);
xnor U16623 (N_16623,N_13437,N_14236);
nor U16624 (N_16624,N_13163,N_13425);
and U16625 (N_16625,N_13723,N_13419);
nand U16626 (N_16626,N_14311,N_13599);
xnor U16627 (N_16627,N_12757,N_14155);
nand U16628 (N_16628,N_13089,N_13810);
or U16629 (N_16629,N_12695,N_13872);
nor U16630 (N_16630,N_14526,N_12752);
nor U16631 (N_16631,N_13477,N_13289);
nand U16632 (N_16632,N_13409,N_13963);
and U16633 (N_16633,N_14242,N_13440);
xnor U16634 (N_16634,N_14767,N_13545);
xnor U16635 (N_16635,N_14842,N_14986);
nand U16636 (N_16636,N_14983,N_13685);
nand U16637 (N_16637,N_13030,N_13975);
nand U16638 (N_16638,N_14276,N_14692);
xnor U16639 (N_16639,N_13613,N_14012);
and U16640 (N_16640,N_12592,N_14632);
xnor U16641 (N_16641,N_14112,N_14453);
and U16642 (N_16642,N_12632,N_14070);
nor U16643 (N_16643,N_14066,N_14346);
and U16644 (N_16644,N_14990,N_13439);
or U16645 (N_16645,N_14803,N_13213);
xor U16646 (N_16646,N_14737,N_13617);
or U16647 (N_16647,N_13690,N_14435);
nand U16648 (N_16648,N_14616,N_13040);
and U16649 (N_16649,N_13112,N_14495);
and U16650 (N_16650,N_13239,N_14272);
or U16651 (N_16651,N_12807,N_14896);
or U16652 (N_16652,N_13506,N_14740);
nor U16653 (N_16653,N_13480,N_13515);
xnor U16654 (N_16654,N_14449,N_14871);
and U16655 (N_16655,N_14848,N_14415);
xor U16656 (N_16656,N_13285,N_14279);
nor U16657 (N_16657,N_12870,N_12558);
and U16658 (N_16658,N_13136,N_13814);
and U16659 (N_16659,N_13801,N_12603);
or U16660 (N_16660,N_13435,N_13514);
nor U16661 (N_16661,N_14143,N_14952);
xnor U16662 (N_16662,N_13651,N_12657);
xnor U16663 (N_16663,N_13075,N_14064);
nand U16664 (N_16664,N_13878,N_13439);
nor U16665 (N_16665,N_13607,N_13879);
or U16666 (N_16666,N_14535,N_13851);
nand U16667 (N_16667,N_14311,N_13701);
and U16668 (N_16668,N_13375,N_14117);
or U16669 (N_16669,N_14457,N_13854);
nor U16670 (N_16670,N_14847,N_13423);
nand U16671 (N_16671,N_14978,N_14661);
or U16672 (N_16672,N_12563,N_13655);
xor U16673 (N_16673,N_14624,N_14186);
nor U16674 (N_16674,N_14442,N_12813);
nor U16675 (N_16675,N_12656,N_14858);
and U16676 (N_16676,N_12777,N_14277);
or U16677 (N_16677,N_14838,N_14381);
and U16678 (N_16678,N_14823,N_13254);
xor U16679 (N_16679,N_13838,N_13144);
xor U16680 (N_16680,N_12886,N_13309);
nand U16681 (N_16681,N_13194,N_14820);
xnor U16682 (N_16682,N_14359,N_14697);
nand U16683 (N_16683,N_14474,N_14712);
xnor U16684 (N_16684,N_14152,N_12629);
and U16685 (N_16685,N_13754,N_13626);
nor U16686 (N_16686,N_14255,N_14654);
xor U16687 (N_16687,N_12700,N_14539);
or U16688 (N_16688,N_13343,N_13301);
nor U16689 (N_16689,N_14897,N_13402);
nor U16690 (N_16690,N_13266,N_14294);
nor U16691 (N_16691,N_12882,N_14192);
xor U16692 (N_16692,N_14695,N_14715);
nor U16693 (N_16693,N_13625,N_13518);
nor U16694 (N_16694,N_12505,N_13960);
and U16695 (N_16695,N_13821,N_13730);
nor U16696 (N_16696,N_12547,N_13976);
nand U16697 (N_16697,N_14010,N_13777);
xor U16698 (N_16698,N_12587,N_12770);
xnor U16699 (N_16699,N_13204,N_12901);
nand U16700 (N_16700,N_13502,N_12860);
and U16701 (N_16701,N_13510,N_13303);
or U16702 (N_16702,N_14892,N_13859);
nand U16703 (N_16703,N_13668,N_13165);
nor U16704 (N_16704,N_13412,N_13673);
xnor U16705 (N_16705,N_13696,N_14037);
xor U16706 (N_16706,N_13090,N_13206);
or U16707 (N_16707,N_13433,N_12903);
nand U16708 (N_16708,N_12556,N_14736);
xor U16709 (N_16709,N_14235,N_13705);
nand U16710 (N_16710,N_13563,N_12877);
nand U16711 (N_16711,N_14579,N_13820);
and U16712 (N_16712,N_13339,N_13454);
xnor U16713 (N_16713,N_12840,N_14649);
nor U16714 (N_16714,N_14733,N_12652);
xor U16715 (N_16715,N_13942,N_13520);
nor U16716 (N_16716,N_13460,N_14883);
or U16717 (N_16717,N_14855,N_13204);
or U16718 (N_16718,N_13967,N_14225);
or U16719 (N_16719,N_14417,N_14821);
nand U16720 (N_16720,N_13495,N_14173);
nor U16721 (N_16721,N_13031,N_12577);
xor U16722 (N_16722,N_12541,N_13124);
and U16723 (N_16723,N_14827,N_13982);
and U16724 (N_16724,N_13416,N_14083);
nand U16725 (N_16725,N_13300,N_14806);
nor U16726 (N_16726,N_12949,N_13329);
nor U16727 (N_16727,N_13278,N_13653);
xnor U16728 (N_16728,N_12776,N_14382);
xnor U16729 (N_16729,N_13757,N_12561);
nor U16730 (N_16730,N_12922,N_13293);
nand U16731 (N_16731,N_14392,N_12553);
and U16732 (N_16732,N_14105,N_13482);
nand U16733 (N_16733,N_14614,N_12741);
nor U16734 (N_16734,N_14293,N_13957);
nor U16735 (N_16735,N_12956,N_14112);
nor U16736 (N_16736,N_13917,N_14843);
xor U16737 (N_16737,N_13201,N_13032);
nor U16738 (N_16738,N_14680,N_13885);
or U16739 (N_16739,N_13675,N_13904);
xor U16740 (N_16740,N_14986,N_13232);
or U16741 (N_16741,N_13936,N_13102);
xnor U16742 (N_16742,N_13896,N_13228);
nand U16743 (N_16743,N_14552,N_14985);
nand U16744 (N_16744,N_14007,N_13477);
or U16745 (N_16745,N_14591,N_14686);
xor U16746 (N_16746,N_12771,N_13152);
nor U16747 (N_16747,N_12764,N_13528);
nand U16748 (N_16748,N_12682,N_13236);
or U16749 (N_16749,N_14110,N_13047);
nand U16750 (N_16750,N_13745,N_14295);
nor U16751 (N_16751,N_13191,N_14123);
nor U16752 (N_16752,N_14958,N_13484);
or U16753 (N_16753,N_14698,N_13900);
and U16754 (N_16754,N_13441,N_13788);
nor U16755 (N_16755,N_12744,N_12742);
and U16756 (N_16756,N_14567,N_13224);
nor U16757 (N_16757,N_13163,N_13224);
and U16758 (N_16758,N_13951,N_12959);
nor U16759 (N_16759,N_12759,N_14933);
or U16760 (N_16760,N_13103,N_13225);
xnor U16761 (N_16761,N_14665,N_13227);
nand U16762 (N_16762,N_14589,N_13551);
and U16763 (N_16763,N_14925,N_13092);
xor U16764 (N_16764,N_13211,N_14788);
nor U16765 (N_16765,N_14265,N_14147);
nand U16766 (N_16766,N_13898,N_13156);
xor U16767 (N_16767,N_13560,N_14642);
xnor U16768 (N_16768,N_14293,N_13024);
nor U16769 (N_16769,N_14319,N_12724);
nor U16770 (N_16770,N_14287,N_14443);
xnor U16771 (N_16771,N_12567,N_14463);
nand U16772 (N_16772,N_14113,N_13702);
nand U16773 (N_16773,N_14451,N_12532);
or U16774 (N_16774,N_14251,N_12993);
nor U16775 (N_16775,N_14889,N_13867);
or U16776 (N_16776,N_14690,N_12715);
nand U16777 (N_16777,N_12934,N_13459);
xor U16778 (N_16778,N_14636,N_12536);
nand U16779 (N_16779,N_13630,N_13324);
and U16780 (N_16780,N_13837,N_14649);
nand U16781 (N_16781,N_13903,N_14483);
nor U16782 (N_16782,N_12692,N_14753);
and U16783 (N_16783,N_12663,N_12962);
nor U16784 (N_16784,N_12638,N_13080);
nand U16785 (N_16785,N_12656,N_14843);
and U16786 (N_16786,N_12957,N_12912);
and U16787 (N_16787,N_14288,N_14377);
xnor U16788 (N_16788,N_14104,N_13697);
xor U16789 (N_16789,N_14547,N_14400);
nor U16790 (N_16790,N_14227,N_13455);
nand U16791 (N_16791,N_14135,N_14567);
xor U16792 (N_16792,N_13677,N_13289);
nor U16793 (N_16793,N_14592,N_13049);
xnor U16794 (N_16794,N_12516,N_13090);
nor U16795 (N_16795,N_12552,N_13312);
nand U16796 (N_16796,N_13779,N_14648);
or U16797 (N_16797,N_13258,N_14793);
nand U16798 (N_16798,N_12567,N_13370);
and U16799 (N_16799,N_14679,N_13547);
or U16800 (N_16800,N_14596,N_14765);
xor U16801 (N_16801,N_13248,N_13445);
or U16802 (N_16802,N_14517,N_12535);
nor U16803 (N_16803,N_13415,N_13716);
nand U16804 (N_16804,N_14756,N_13039);
xor U16805 (N_16805,N_13175,N_13029);
or U16806 (N_16806,N_14027,N_14898);
nor U16807 (N_16807,N_14483,N_14737);
or U16808 (N_16808,N_12957,N_14292);
xor U16809 (N_16809,N_14997,N_13609);
nand U16810 (N_16810,N_13237,N_14832);
and U16811 (N_16811,N_13938,N_12786);
nand U16812 (N_16812,N_13877,N_14714);
xnor U16813 (N_16813,N_13866,N_12880);
xor U16814 (N_16814,N_13006,N_14129);
nor U16815 (N_16815,N_14936,N_14954);
nand U16816 (N_16816,N_14055,N_14393);
or U16817 (N_16817,N_14266,N_14531);
nand U16818 (N_16818,N_14814,N_12905);
xnor U16819 (N_16819,N_14840,N_14545);
and U16820 (N_16820,N_14109,N_12760);
xor U16821 (N_16821,N_14517,N_14147);
xor U16822 (N_16822,N_12547,N_12705);
and U16823 (N_16823,N_12626,N_13651);
nor U16824 (N_16824,N_14538,N_12686);
nor U16825 (N_16825,N_13732,N_13298);
or U16826 (N_16826,N_14880,N_13993);
xnor U16827 (N_16827,N_14604,N_14569);
and U16828 (N_16828,N_14992,N_14911);
nor U16829 (N_16829,N_14764,N_14087);
or U16830 (N_16830,N_13699,N_14393);
or U16831 (N_16831,N_14791,N_14480);
xnor U16832 (N_16832,N_14379,N_14829);
xor U16833 (N_16833,N_13520,N_13667);
or U16834 (N_16834,N_14819,N_14235);
or U16835 (N_16835,N_13369,N_14419);
nand U16836 (N_16836,N_12766,N_14044);
and U16837 (N_16837,N_14626,N_14485);
and U16838 (N_16838,N_13580,N_14890);
nor U16839 (N_16839,N_12625,N_12938);
nor U16840 (N_16840,N_13039,N_13520);
or U16841 (N_16841,N_14587,N_14965);
nor U16842 (N_16842,N_12870,N_14078);
and U16843 (N_16843,N_13374,N_14959);
nand U16844 (N_16844,N_14478,N_14419);
nor U16845 (N_16845,N_12798,N_13792);
or U16846 (N_16846,N_13544,N_14905);
or U16847 (N_16847,N_13513,N_14293);
xnor U16848 (N_16848,N_13013,N_14518);
or U16849 (N_16849,N_13295,N_14307);
xor U16850 (N_16850,N_14310,N_14039);
nor U16851 (N_16851,N_14966,N_14390);
xnor U16852 (N_16852,N_13921,N_14182);
nand U16853 (N_16853,N_14265,N_12592);
nor U16854 (N_16854,N_12624,N_13519);
and U16855 (N_16855,N_14437,N_14304);
xnor U16856 (N_16856,N_13700,N_13628);
nor U16857 (N_16857,N_14095,N_14731);
and U16858 (N_16858,N_14237,N_14844);
nand U16859 (N_16859,N_13675,N_14366);
nor U16860 (N_16860,N_13670,N_12861);
nand U16861 (N_16861,N_14464,N_13788);
or U16862 (N_16862,N_14024,N_14562);
nor U16863 (N_16863,N_14819,N_14048);
or U16864 (N_16864,N_14779,N_13217);
xnor U16865 (N_16865,N_13510,N_14844);
nand U16866 (N_16866,N_13113,N_12674);
or U16867 (N_16867,N_14000,N_13134);
xnor U16868 (N_16868,N_14208,N_13663);
nor U16869 (N_16869,N_14120,N_14825);
xnor U16870 (N_16870,N_12739,N_14485);
or U16871 (N_16871,N_12592,N_13996);
nand U16872 (N_16872,N_14281,N_13178);
nand U16873 (N_16873,N_13523,N_13674);
and U16874 (N_16874,N_12504,N_14208);
and U16875 (N_16875,N_13175,N_13877);
nor U16876 (N_16876,N_14976,N_13240);
nor U16877 (N_16877,N_14036,N_13358);
xnor U16878 (N_16878,N_12978,N_14075);
and U16879 (N_16879,N_13226,N_13659);
nor U16880 (N_16880,N_13122,N_12682);
nor U16881 (N_16881,N_14877,N_14484);
nor U16882 (N_16882,N_14892,N_14635);
xor U16883 (N_16883,N_14079,N_13226);
and U16884 (N_16884,N_14655,N_13411);
xnor U16885 (N_16885,N_12788,N_14084);
or U16886 (N_16886,N_14228,N_13720);
and U16887 (N_16887,N_14701,N_14179);
xor U16888 (N_16888,N_14015,N_13217);
and U16889 (N_16889,N_12601,N_12875);
nand U16890 (N_16890,N_14126,N_13800);
nor U16891 (N_16891,N_13186,N_14044);
and U16892 (N_16892,N_12887,N_13168);
nor U16893 (N_16893,N_13597,N_13110);
or U16894 (N_16894,N_14488,N_14641);
and U16895 (N_16895,N_13179,N_14868);
and U16896 (N_16896,N_14120,N_14289);
or U16897 (N_16897,N_12803,N_13935);
nor U16898 (N_16898,N_14290,N_14225);
and U16899 (N_16899,N_13206,N_13249);
and U16900 (N_16900,N_13124,N_13911);
nand U16901 (N_16901,N_13282,N_13508);
nor U16902 (N_16902,N_13637,N_13831);
nand U16903 (N_16903,N_14117,N_14841);
nand U16904 (N_16904,N_14977,N_12835);
nand U16905 (N_16905,N_13432,N_13673);
and U16906 (N_16906,N_12547,N_14500);
nor U16907 (N_16907,N_13978,N_14778);
nand U16908 (N_16908,N_13089,N_14849);
xor U16909 (N_16909,N_13325,N_14381);
nor U16910 (N_16910,N_14767,N_12827);
nand U16911 (N_16911,N_13547,N_14286);
nand U16912 (N_16912,N_14101,N_13602);
or U16913 (N_16913,N_13878,N_12708);
or U16914 (N_16914,N_14737,N_13428);
or U16915 (N_16915,N_14702,N_13132);
nand U16916 (N_16916,N_13163,N_14353);
or U16917 (N_16917,N_14686,N_14679);
nor U16918 (N_16918,N_14974,N_13628);
or U16919 (N_16919,N_14843,N_13659);
and U16920 (N_16920,N_13239,N_14550);
and U16921 (N_16921,N_14289,N_14957);
nor U16922 (N_16922,N_13179,N_13123);
and U16923 (N_16923,N_14306,N_13095);
or U16924 (N_16924,N_14082,N_13303);
nand U16925 (N_16925,N_14559,N_12935);
or U16926 (N_16926,N_13005,N_12868);
and U16927 (N_16927,N_13501,N_12966);
nor U16928 (N_16928,N_14384,N_14610);
and U16929 (N_16929,N_14606,N_12806);
and U16930 (N_16930,N_13849,N_13787);
nor U16931 (N_16931,N_13912,N_13751);
or U16932 (N_16932,N_14535,N_13904);
xnor U16933 (N_16933,N_13551,N_13542);
and U16934 (N_16934,N_13451,N_12551);
nor U16935 (N_16935,N_13236,N_12530);
and U16936 (N_16936,N_13191,N_13693);
nand U16937 (N_16937,N_13692,N_14417);
nor U16938 (N_16938,N_13299,N_13698);
xnor U16939 (N_16939,N_14329,N_14390);
and U16940 (N_16940,N_13165,N_14103);
or U16941 (N_16941,N_14234,N_13871);
nand U16942 (N_16942,N_13611,N_14358);
nand U16943 (N_16943,N_14532,N_14095);
or U16944 (N_16944,N_13835,N_14999);
and U16945 (N_16945,N_13874,N_13581);
xnor U16946 (N_16946,N_13969,N_14056);
nor U16947 (N_16947,N_14428,N_12645);
or U16948 (N_16948,N_13239,N_12978);
or U16949 (N_16949,N_14795,N_12700);
xnor U16950 (N_16950,N_13717,N_12588);
or U16951 (N_16951,N_13137,N_14177);
or U16952 (N_16952,N_13223,N_13556);
nand U16953 (N_16953,N_14264,N_14831);
or U16954 (N_16954,N_13110,N_13503);
nor U16955 (N_16955,N_14203,N_14491);
xor U16956 (N_16956,N_13119,N_12713);
xnor U16957 (N_16957,N_13324,N_14482);
nand U16958 (N_16958,N_13465,N_14544);
nor U16959 (N_16959,N_12863,N_14312);
nor U16960 (N_16960,N_12888,N_12882);
nand U16961 (N_16961,N_13956,N_14211);
and U16962 (N_16962,N_13230,N_13276);
nand U16963 (N_16963,N_14651,N_13648);
nor U16964 (N_16964,N_14571,N_13725);
or U16965 (N_16965,N_14447,N_12676);
nor U16966 (N_16966,N_12754,N_13000);
or U16967 (N_16967,N_13426,N_14774);
nor U16968 (N_16968,N_13788,N_14287);
xor U16969 (N_16969,N_12761,N_13020);
nor U16970 (N_16970,N_12550,N_13843);
xor U16971 (N_16971,N_14848,N_13020);
xnor U16972 (N_16972,N_12628,N_14769);
nand U16973 (N_16973,N_12705,N_13527);
nor U16974 (N_16974,N_12625,N_14392);
nand U16975 (N_16975,N_13918,N_14670);
or U16976 (N_16976,N_12716,N_14085);
and U16977 (N_16977,N_12593,N_14500);
nor U16978 (N_16978,N_12982,N_14723);
and U16979 (N_16979,N_13268,N_14130);
nand U16980 (N_16980,N_13432,N_13924);
nor U16981 (N_16981,N_12951,N_13728);
nand U16982 (N_16982,N_13179,N_14369);
nor U16983 (N_16983,N_12911,N_12950);
nand U16984 (N_16984,N_14876,N_12535);
or U16985 (N_16985,N_14064,N_12534);
nand U16986 (N_16986,N_14264,N_12911);
and U16987 (N_16987,N_14454,N_12565);
xnor U16988 (N_16988,N_14750,N_12724);
or U16989 (N_16989,N_12575,N_14192);
xnor U16990 (N_16990,N_12747,N_13593);
or U16991 (N_16991,N_13166,N_12802);
and U16992 (N_16992,N_13264,N_14243);
or U16993 (N_16993,N_14060,N_13689);
nor U16994 (N_16994,N_13957,N_14702);
xnor U16995 (N_16995,N_14949,N_12917);
nand U16996 (N_16996,N_12721,N_14185);
nand U16997 (N_16997,N_14419,N_13985);
and U16998 (N_16998,N_14013,N_13521);
or U16999 (N_16999,N_12535,N_13328);
nand U17000 (N_17000,N_14323,N_13813);
or U17001 (N_17001,N_14799,N_13188);
or U17002 (N_17002,N_12509,N_14123);
nor U17003 (N_17003,N_12749,N_13306);
nor U17004 (N_17004,N_14973,N_13031);
nor U17005 (N_17005,N_14059,N_13609);
nand U17006 (N_17006,N_12556,N_12820);
and U17007 (N_17007,N_12981,N_13227);
nand U17008 (N_17008,N_14041,N_13789);
and U17009 (N_17009,N_14644,N_14720);
nand U17010 (N_17010,N_14289,N_14664);
nor U17011 (N_17011,N_13397,N_14723);
nor U17012 (N_17012,N_12767,N_14847);
xor U17013 (N_17013,N_13710,N_12937);
and U17014 (N_17014,N_12957,N_14989);
nor U17015 (N_17015,N_12816,N_13826);
nor U17016 (N_17016,N_12963,N_13656);
nor U17017 (N_17017,N_13880,N_14228);
nor U17018 (N_17018,N_13148,N_14453);
xor U17019 (N_17019,N_12870,N_14236);
xor U17020 (N_17020,N_14409,N_12731);
xor U17021 (N_17021,N_14346,N_14488);
or U17022 (N_17022,N_13379,N_12890);
nand U17023 (N_17023,N_12915,N_12851);
nand U17024 (N_17024,N_14509,N_14612);
and U17025 (N_17025,N_13206,N_12619);
nand U17026 (N_17026,N_12719,N_13821);
or U17027 (N_17027,N_13648,N_13064);
nor U17028 (N_17028,N_13566,N_13919);
or U17029 (N_17029,N_14843,N_12844);
nand U17030 (N_17030,N_14412,N_13117);
or U17031 (N_17031,N_12531,N_13294);
or U17032 (N_17032,N_13603,N_12576);
and U17033 (N_17033,N_13999,N_14182);
nand U17034 (N_17034,N_14554,N_14388);
xor U17035 (N_17035,N_13460,N_14650);
xnor U17036 (N_17036,N_14069,N_14817);
and U17037 (N_17037,N_13375,N_13655);
or U17038 (N_17038,N_13265,N_14105);
nor U17039 (N_17039,N_13442,N_12795);
xnor U17040 (N_17040,N_13085,N_13785);
nand U17041 (N_17041,N_14939,N_13192);
nand U17042 (N_17042,N_13370,N_13841);
nor U17043 (N_17043,N_13477,N_14768);
nand U17044 (N_17044,N_14559,N_13417);
nor U17045 (N_17045,N_14680,N_12970);
nor U17046 (N_17046,N_14738,N_14165);
nand U17047 (N_17047,N_13567,N_14938);
or U17048 (N_17048,N_12510,N_14256);
or U17049 (N_17049,N_13888,N_12800);
xor U17050 (N_17050,N_13766,N_13543);
or U17051 (N_17051,N_14095,N_14157);
nand U17052 (N_17052,N_13488,N_13071);
and U17053 (N_17053,N_14297,N_14800);
and U17054 (N_17054,N_12843,N_12749);
nand U17055 (N_17055,N_13704,N_12615);
xor U17056 (N_17056,N_14675,N_13246);
nor U17057 (N_17057,N_12615,N_13541);
xnor U17058 (N_17058,N_13450,N_14459);
and U17059 (N_17059,N_12734,N_14258);
nand U17060 (N_17060,N_13073,N_14524);
or U17061 (N_17061,N_14283,N_14166);
nand U17062 (N_17062,N_14817,N_13945);
nor U17063 (N_17063,N_13233,N_12955);
and U17064 (N_17064,N_13793,N_13624);
and U17065 (N_17065,N_12749,N_14040);
nor U17066 (N_17066,N_14135,N_13958);
xnor U17067 (N_17067,N_13776,N_14347);
nor U17068 (N_17068,N_13510,N_14614);
xnor U17069 (N_17069,N_12838,N_12668);
or U17070 (N_17070,N_14341,N_13461);
nand U17071 (N_17071,N_12781,N_13497);
and U17072 (N_17072,N_12848,N_13320);
xnor U17073 (N_17073,N_13568,N_14727);
xnor U17074 (N_17074,N_13221,N_13721);
xnor U17075 (N_17075,N_13228,N_12633);
and U17076 (N_17076,N_14905,N_13554);
nand U17077 (N_17077,N_14075,N_13424);
nand U17078 (N_17078,N_14025,N_14162);
and U17079 (N_17079,N_14129,N_14144);
or U17080 (N_17080,N_14737,N_14247);
nand U17081 (N_17081,N_13987,N_14524);
nand U17082 (N_17082,N_14397,N_13507);
nor U17083 (N_17083,N_13322,N_14447);
or U17084 (N_17084,N_13520,N_13223);
nor U17085 (N_17085,N_14552,N_13499);
nor U17086 (N_17086,N_12570,N_14972);
or U17087 (N_17087,N_13301,N_14555);
or U17088 (N_17088,N_14195,N_14286);
or U17089 (N_17089,N_14268,N_13409);
or U17090 (N_17090,N_13537,N_13749);
or U17091 (N_17091,N_14292,N_13952);
or U17092 (N_17092,N_13853,N_13739);
or U17093 (N_17093,N_14452,N_13697);
xor U17094 (N_17094,N_13712,N_13127);
xor U17095 (N_17095,N_13333,N_14318);
nand U17096 (N_17096,N_13260,N_13725);
xnor U17097 (N_17097,N_12841,N_14270);
nor U17098 (N_17098,N_13812,N_13195);
or U17099 (N_17099,N_14624,N_14945);
and U17100 (N_17100,N_12948,N_14930);
xor U17101 (N_17101,N_12571,N_14300);
or U17102 (N_17102,N_13875,N_14115);
nand U17103 (N_17103,N_14105,N_12524);
nor U17104 (N_17104,N_13571,N_14823);
nor U17105 (N_17105,N_13899,N_12817);
nor U17106 (N_17106,N_12868,N_13851);
nor U17107 (N_17107,N_14658,N_12720);
or U17108 (N_17108,N_13236,N_14105);
xor U17109 (N_17109,N_13489,N_14532);
nand U17110 (N_17110,N_14041,N_13702);
nand U17111 (N_17111,N_14721,N_13277);
or U17112 (N_17112,N_14475,N_13637);
or U17113 (N_17113,N_14758,N_13732);
xnor U17114 (N_17114,N_14704,N_13047);
xor U17115 (N_17115,N_12782,N_13153);
xnor U17116 (N_17116,N_14835,N_14054);
and U17117 (N_17117,N_14001,N_12676);
nand U17118 (N_17118,N_13002,N_13947);
nor U17119 (N_17119,N_13910,N_12524);
or U17120 (N_17120,N_13767,N_14430);
or U17121 (N_17121,N_14369,N_13332);
nand U17122 (N_17122,N_14621,N_14642);
and U17123 (N_17123,N_13229,N_14231);
xor U17124 (N_17124,N_13598,N_14517);
or U17125 (N_17125,N_13944,N_14243);
and U17126 (N_17126,N_14724,N_14334);
and U17127 (N_17127,N_13976,N_12983);
nor U17128 (N_17128,N_13527,N_13321);
or U17129 (N_17129,N_13715,N_13001);
and U17130 (N_17130,N_13572,N_13252);
and U17131 (N_17131,N_12975,N_14576);
nand U17132 (N_17132,N_12637,N_13554);
or U17133 (N_17133,N_13381,N_14122);
nor U17134 (N_17134,N_14931,N_13484);
nor U17135 (N_17135,N_14400,N_13874);
and U17136 (N_17136,N_14265,N_13004);
and U17137 (N_17137,N_14370,N_13811);
or U17138 (N_17138,N_13606,N_14300);
and U17139 (N_17139,N_12658,N_13187);
nor U17140 (N_17140,N_12825,N_14691);
nor U17141 (N_17141,N_13523,N_13343);
or U17142 (N_17142,N_13777,N_14571);
and U17143 (N_17143,N_12650,N_14104);
xor U17144 (N_17144,N_12659,N_13954);
and U17145 (N_17145,N_12691,N_13880);
nor U17146 (N_17146,N_14002,N_12738);
nor U17147 (N_17147,N_14682,N_12992);
and U17148 (N_17148,N_12711,N_14110);
nor U17149 (N_17149,N_13601,N_13588);
xnor U17150 (N_17150,N_12885,N_13590);
and U17151 (N_17151,N_12831,N_13062);
nor U17152 (N_17152,N_14861,N_12962);
nand U17153 (N_17153,N_12502,N_13654);
and U17154 (N_17154,N_14849,N_14551);
nand U17155 (N_17155,N_14916,N_14479);
nor U17156 (N_17156,N_13990,N_14627);
and U17157 (N_17157,N_12647,N_14418);
nor U17158 (N_17158,N_13264,N_12708);
or U17159 (N_17159,N_12983,N_12626);
or U17160 (N_17160,N_14117,N_13238);
and U17161 (N_17161,N_13845,N_13806);
nor U17162 (N_17162,N_12821,N_13753);
and U17163 (N_17163,N_14076,N_14113);
or U17164 (N_17164,N_14176,N_13031);
or U17165 (N_17165,N_13399,N_13686);
nor U17166 (N_17166,N_14793,N_12810);
and U17167 (N_17167,N_13211,N_12827);
xnor U17168 (N_17168,N_13179,N_13575);
nor U17169 (N_17169,N_13771,N_14207);
or U17170 (N_17170,N_13534,N_13822);
and U17171 (N_17171,N_14477,N_12845);
and U17172 (N_17172,N_13667,N_12630);
xor U17173 (N_17173,N_14309,N_13834);
nor U17174 (N_17174,N_14821,N_13780);
nand U17175 (N_17175,N_13725,N_14369);
nand U17176 (N_17176,N_13387,N_12520);
nor U17177 (N_17177,N_14297,N_14438);
nand U17178 (N_17178,N_12895,N_12976);
and U17179 (N_17179,N_12665,N_12731);
xor U17180 (N_17180,N_14950,N_13899);
or U17181 (N_17181,N_13216,N_14087);
and U17182 (N_17182,N_13636,N_13258);
or U17183 (N_17183,N_12543,N_12667);
nand U17184 (N_17184,N_13400,N_13563);
xor U17185 (N_17185,N_14529,N_13325);
and U17186 (N_17186,N_14196,N_13921);
nand U17187 (N_17187,N_12659,N_14500);
and U17188 (N_17188,N_14811,N_12596);
or U17189 (N_17189,N_14301,N_12809);
nor U17190 (N_17190,N_13897,N_13678);
nand U17191 (N_17191,N_13726,N_12713);
xnor U17192 (N_17192,N_13550,N_14312);
and U17193 (N_17193,N_13753,N_14899);
xnor U17194 (N_17194,N_12937,N_13026);
or U17195 (N_17195,N_13216,N_13117);
nand U17196 (N_17196,N_14241,N_14843);
xnor U17197 (N_17197,N_14492,N_12568);
xnor U17198 (N_17198,N_13378,N_14930);
xnor U17199 (N_17199,N_12794,N_14650);
nand U17200 (N_17200,N_14622,N_14463);
xor U17201 (N_17201,N_13300,N_12514);
nor U17202 (N_17202,N_12575,N_13904);
nor U17203 (N_17203,N_14879,N_13573);
or U17204 (N_17204,N_13426,N_12884);
and U17205 (N_17205,N_13033,N_14423);
xnor U17206 (N_17206,N_14842,N_14946);
nand U17207 (N_17207,N_13561,N_12500);
and U17208 (N_17208,N_13553,N_13386);
nand U17209 (N_17209,N_12866,N_13845);
xnor U17210 (N_17210,N_13601,N_14447);
or U17211 (N_17211,N_14328,N_13169);
nor U17212 (N_17212,N_13954,N_13754);
or U17213 (N_17213,N_13479,N_13473);
nor U17214 (N_17214,N_14768,N_14573);
nand U17215 (N_17215,N_14340,N_13751);
or U17216 (N_17216,N_14438,N_14851);
xnor U17217 (N_17217,N_13755,N_14644);
nor U17218 (N_17218,N_13871,N_14707);
xnor U17219 (N_17219,N_13395,N_14946);
xor U17220 (N_17220,N_13196,N_14097);
and U17221 (N_17221,N_13318,N_12653);
or U17222 (N_17222,N_12610,N_12977);
and U17223 (N_17223,N_12870,N_14071);
nand U17224 (N_17224,N_14412,N_14352);
xor U17225 (N_17225,N_14059,N_12691);
and U17226 (N_17226,N_13046,N_12836);
nand U17227 (N_17227,N_14615,N_12941);
and U17228 (N_17228,N_14296,N_14123);
nand U17229 (N_17229,N_14461,N_14707);
xnor U17230 (N_17230,N_14303,N_14238);
xor U17231 (N_17231,N_13890,N_13602);
and U17232 (N_17232,N_13199,N_12552);
and U17233 (N_17233,N_13110,N_14333);
or U17234 (N_17234,N_12638,N_14688);
and U17235 (N_17235,N_12686,N_13318);
or U17236 (N_17236,N_14782,N_13797);
xnor U17237 (N_17237,N_13681,N_12755);
or U17238 (N_17238,N_12641,N_14533);
nand U17239 (N_17239,N_13817,N_14550);
xnor U17240 (N_17240,N_12733,N_12536);
or U17241 (N_17241,N_14072,N_13620);
or U17242 (N_17242,N_14984,N_12934);
nand U17243 (N_17243,N_14813,N_12985);
or U17244 (N_17244,N_13018,N_13733);
nand U17245 (N_17245,N_13944,N_14882);
or U17246 (N_17246,N_13057,N_12501);
nand U17247 (N_17247,N_13983,N_14697);
xor U17248 (N_17248,N_13082,N_12770);
nand U17249 (N_17249,N_12627,N_14107);
or U17250 (N_17250,N_13387,N_14972);
nor U17251 (N_17251,N_14955,N_13825);
nand U17252 (N_17252,N_13308,N_13551);
and U17253 (N_17253,N_13302,N_13870);
and U17254 (N_17254,N_12610,N_14343);
and U17255 (N_17255,N_13507,N_14117);
nor U17256 (N_17256,N_13153,N_14626);
xnor U17257 (N_17257,N_13899,N_14336);
and U17258 (N_17258,N_14102,N_13869);
nor U17259 (N_17259,N_14622,N_12715);
xnor U17260 (N_17260,N_13397,N_12552);
and U17261 (N_17261,N_12696,N_14865);
or U17262 (N_17262,N_13127,N_13021);
nand U17263 (N_17263,N_14820,N_13410);
nand U17264 (N_17264,N_14752,N_14811);
xor U17265 (N_17265,N_12811,N_13657);
xnor U17266 (N_17266,N_13128,N_12924);
and U17267 (N_17267,N_13285,N_13060);
xor U17268 (N_17268,N_14058,N_14826);
nand U17269 (N_17269,N_13979,N_14013);
nor U17270 (N_17270,N_12810,N_14978);
nand U17271 (N_17271,N_14781,N_14035);
nand U17272 (N_17272,N_14460,N_14228);
nand U17273 (N_17273,N_14282,N_14503);
or U17274 (N_17274,N_14346,N_14075);
or U17275 (N_17275,N_13297,N_13316);
nand U17276 (N_17276,N_13492,N_14248);
nand U17277 (N_17277,N_14873,N_14957);
nor U17278 (N_17278,N_13557,N_12552);
or U17279 (N_17279,N_13471,N_14545);
nor U17280 (N_17280,N_13378,N_13058);
xnor U17281 (N_17281,N_13664,N_14664);
or U17282 (N_17282,N_12813,N_13110);
nor U17283 (N_17283,N_13449,N_12943);
or U17284 (N_17284,N_14773,N_13836);
xnor U17285 (N_17285,N_13903,N_13834);
nor U17286 (N_17286,N_12682,N_14394);
and U17287 (N_17287,N_13159,N_13930);
or U17288 (N_17288,N_12541,N_14261);
nand U17289 (N_17289,N_13278,N_13287);
xnor U17290 (N_17290,N_13873,N_14275);
and U17291 (N_17291,N_14986,N_13139);
xnor U17292 (N_17292,N_14978,N_13864);
xnor U17293 (N_17293,N_14973,N_13608);
and U17294 (N_17294,N_13179,N_12624);
nor U17295 (N_17295,N_13483,N_14906);
nor U17296 (N_17296,N_13611,N_13572);
nand U17297 (N_17297,N_14870,N_13102);
xor U17298 (N_17298,N_13450,N_13865);
and U17299 (N_17299,N_13046,N_13192);
xor U17300 (N_17300,N_13130,N_14485);
xnor U17301 (N_17301,N_14937,N_14344);
and U17302 (N_17302,N_14944,N_14395);
xor U17303 (N_17303,N_13704,N_14235);
and U17304 (N_17304,N_14799,N_14434);
and U17305 (N_17305,N_12965,N_14915);
or U17306 (N_17306,N_14114,N_12625);
or U17307 (N_17307,N_14208,N_12874);
nand U17308 (N_17308,N_14477,N_13842);
nand U17309 (N_17309,N_13435,N_14678);
or U17310 (N_17310,N_14320,N_14272);
or U17311 (N_17311,N_13813,N_14006);
xnor U17312 (N_17312,N_13045,N_12866);
xor U17313 (N_17313,N_13545,N_13350);
or U17314 (N_17314,N_14449,N_13506);
xnor U17315 (N_17315,N_13377,N_14169);
xor U17316 (N_17316,N_13659,N_12613);
or U17317 (N_17317,N_14238,N_14767);
xor U17318 (N_17318,N_13063,N_13834);
xnor U17319 (N_17319,N_14361,N_14617);
nand U17320 (N_17320,N_14992,N_12855);
nand U17321 (N_17321,N_13872,N_13906);
nor U17322 (N_17322,N_14916,N_12995);
or U17323 (N_17323,N_13315,N_12588);
nand U17324 (N_17324,N_14670,N_13125);
and U17325 (N_17325,N_14823,N_13417);
nand U17326 (N_17326,N_13675,N_13943);
and U17327 (N_17327,N_13143,N_14636);
nand U17328 (N_17328,N_14026,N_13336);
nand U17329 (N_17329,N_14208,N_12873);
nand U17330 (N_17330,N_14555,N_14316);
nand U17331 (N_17331,N_13639,N_12725);
nand U17332 (N_17332,N_13760,N_12677);
and U17333 (N_17333,N_13539,N_13741);
and U17334 (N_17334,N_13119,N_13365);
nor U17335 (N_17335,N_13974,N_14281);
xor U17336 (N_17336,N_13798,N_13407);
and U17337 (N_17337,N_14559,N_13389);
xor U17338 (N_17338,N_14057,N_12683);
and U17339 (N_17339,N_13095,N_14847);
and U17340 (N_17340,N_13009,N_13182);
nor U17341 (N_17341,N_12501,N_14315);
xor U17342 (N_17342,N_14011,N_13277);
or U17343 (N_17343,N_13658,N_14612);
nor U17344 (N_17344,N_14324,N_14958);
xor U17345 (N_17345,N_14242,N_14334);
or U17346 (N_17346,N_13901,N_12568);
nor U17347 (N_17347,N_13340,N_14942);
and U17348 (N_17348,N_14031,N_14939);
or U17349 (N_17349,N_13366,N_13194);
nand U17350 (N_17350,N_12801,N_14700);
or U17351 (N_17351,N_13383,N_14705);
nor U17352 (N_17352,N_12547,N_14634);
xor U17353 (N_17353,N_13522,N_12984);
nand U17354 (N_17354,N_13298,N_13911);
or U17355 (N_17355,N_14939,N_14695);
nand U17356 (N_17356,N_14918,N_13559);
or U17357 (N_17357,N_13211,N_13880);
nand U17358 (N_17358,N_12875,N_13035);
and U17359 (N_17359,N_14457,N_14510);
or U17360 (N_17360,N_13443,N_13244);
xnor U17361 (N_17361,N_14675,N_13403);
nand U17362 (N_17362,N_12926,N_13666);
nor U17363 (N_17363,N_12632,N_13087);
nand U17364 (N_17364,N_13915,N_14065);
or U17365 (N_17365,N_12882,N_13822);
and U17366 (N_17366,N_13453,N_12585);
and U17367 (N_17367,N_14010,N_14066);
nand U17368 (N_17368,N_14989,N_13357);
and U17369 (N_17369,N_14550,N_14121);
or U17370 (N_17370,N_14314,N_13082);
xor U17371 (N_17371,N_14339,N_13918);
nor U17372 (N_17372,N_14861,N_12841);
and U17373 (N_17373,N_13871,N_12642);
nor U17374 (N_17374,N_13909,N_14491);
nand U17375 (N_17375,N_12577,N_13412);
or U17376 (N_17376,N_12839,N_14567);
or U17377 (N_17377,N_13516,N_13002);
nor U17378 (N_17378,N_14659,N_13129);
and U17379 (N_17379,N_13604,N_14227);
or U17380 (N_17380,N_14161,N_14569);
and U17381 (N_17381,N_13445,N_14132);
nor U17382 (N_17382,N_14538,N_14916);
nor U17383 (N_17383,N_14245,N_12876);
nand U17384 (N_17384,N_12540,N_12739);
nand U17385 (N_17385,N_12801,N_13080);
and U17386 (N_17386,N_12650,N_12523);
nand U17387 (N_17387,N_13531,N_13963);
nor U17388 (N_17388,N_13977,N_14706);
xor U17389 (N_17389,N_12755,N_13476);
nor U17390 (N_17390,N_13850,N_13615);
xor U17391 (N_17391,N_14742,N_13653);
nand U17392 (N_17392,N_13583,N_13437);
or U17393 (N_17393,N_14946,N_13553);
xnor U17394 (N_17394,N_14912,N_13457);
and U17395 (N_17395,N_12600,N_14138);
xnor U17396 (N_17396,N_14452,N_13287);
or U17397 (N_17397,N_14208,N_14038);
or U17398 (N_17398,N_12509,N_14759);
nor U17399 (N_17399,N_12982,N_14057);
or U17400 (N_17400,N_12643,N_13938);
or U17401 (N_17401,N_13558,N_12723);
xor U17402 (N_17402,N_14369,N_14254);
and U17403 (N_17403,N_13471,N_14599);
or U17404 (N_17404,N_12670,N_14058);
nor U17405 (N_17405,N_13616,N_14893);
and U17406 (N_17406,N_12986,N_13556);
nor U17407 (N_17407,N_14999,N_13644);
nand U17408 (N_17408,N_13123,N_14563);
or U17409 (N_17409,N_13197,N_14722);
nor U17410 (N_17410,N_14564,N_14204);
and U17411 (N_17411,N_12502,N_14134);
nand U17412 (N_17412,N_14563,N_12642);
or U17413 (N_17413,N_13481,N_12742);
xor U17414 (N_17414,N_14369,N_14766);
nand U17415 (N_17415,N_14174,N_12796);
nand U17416 (N_17416,N_13728,N_13008);
nand U17417 (N_17417,N_14444,N_14700);
or U17418 (N_17418,N_14310,N_12876);
nand U17419 (N_17419,N_13195,N_13332);
nor U17420 (N_17420,N_13524,N_13140);
xnor U17421 (N_17421,N_12669,N_14879);
or U17422 (N_17422,N_14283,N_12964);
nand U17423 (N_17423,N_14525,N_14286);
nand U17424 (N_17424,N_14120,N_14236);
nor U17425 (N_17425,N_13395,N_14609);
nor U17426 (N_17426,N_13590,N_12799);
nand U17427 (N_17427,N_13179,N_14881);
or U17428 (N_17428,N_13642,N_14011);
nand U17429 (N_17429,N_12903,N_14021);
or U17430 (N_17430,N_13992,N_13734);
xnor U17431 (N_17431,N_13649,N_12644);
or U17432 (N_17432,N_12886,N_14773);
nor U17433 (N_17433,N_13115,N_14723);
and U17434 (N_17434,N_13980,N_13928);
nor U17435 (N_17435,N_13868,N_13313);
xnor U17436 (N_17436,N_13581,N_13627);
nor U17437 (N_17437,N_13315,N_14159);
nand U17438 (N_17438,N_12564,N_13797);
nor U17439 (N_17439,N_13608,N_13491);
nand U17440 (N_17440,N_14600,N_13336);
nor U17441 (N_17441,N_14180,N_12780);
nor U17442 (N_17442,N_14884,N_14867);
xnor U17443 (N_17443,N_14874,N_13758);
xor U17444 (N_17444,N_13602,N_13343);
nand U17445 (N_17445,N_14703,N_12894);
nand U17446 (N_17446,N_12716,N_12952);
nand U17447 (N_17447,N_14179,N_13077);
and U17448 (N_17448,N_13463,N_14772);
nand U17449 (N_17449,N_12590,N_12683);
xnor U17450 (N_17450,N_12772,N_12626);
xor U17451 (N_17451,N_13117,N_12665);
xnor U17452 (N_17452,N_13663,N_14337);
or U17453 (N_17453,N_13020,N_13136);
or U17454 (N_17454,N_14128,N_12705);
xnor U17455 (N_17455,N_13788,N_13619);
nor U17456 (N_17456,N_14755,N_12869);
nand U17457 (N_17457,N_13314,N_13055);
or U17458 (N_17458,N_13609,N_12954);
and U17459 (N_17459,N_14336,N_14167);
and U17460 (N_17460,N_12794,N_13945);
or U17461 (N_17461,N_12951,N_12784);
or U17462 (N_17462,N_14671,N_13285);
or U17463 (N_17463,N_12606,N_13923);
nor U17464 (N_17464,N_13025,N_13426);
xor U17465 (N_17465,N_13004,N_12766);
xor U17466 (N_17466,N_13742,N_14913);
nor U17467 (N_17467,N_14614,N_13989);
xor U17468 (N_17468,N_13256,N_13649);
nor U17469 (N_17469,N_14571,N_14096);
and U17470 (N_17470,N_13845,N_14857);
xnor U17471 (N_17471,N_12668,N_14110);
nor U17472 (N_17472,N_12643,N_12538);
and U17473 (N_17473,N_14360,N_14044);
nor U17474 (N_17474,N_13118,N_12716);
or U17475 (N_17475,N_14576,N_12969);
nand U17476 (N_17476,N_13118,N_14482);
or U17477 (N_17477,N_14263,N_14041);
nor U17478 (N_17478,N_12595,N_13176);
or U17479 (N_17479,N_13546,N_14830);
or U17480 (N_17480,N_13556,N_14588);
nand U17481 (N_17481,N_13554,N_14758);
nor U17482 (N_17482,N_14118,N_14306);
or U17483 (N_17483,N_13312,N_14881);
or U17484 (N_17484,N_12708,N_14894);
nor U17485 (N_17485,N_14389,N_13543);
nand U17486 (N_17486,N_13333,N_13293);
xnor U17487 (N_17487,N_13876,N_13244);
and U17488 (N_17488,N_12846,N_14104);
nand U17489 (N_17489,N_13462,N_14453);
xnor U17490 (N_17490,N_14350,N_13925);
nand U17491 (N_17491,N_13191,N_13902);
and U17492 (N_17492,N_14449,N_14901);
and U17493 (N_17493,N_12951,N_14079);
and U17494 (N_17494,N_13627,N_12552);
and U17495 (N_17495,N_14033,N_14223);
nand U17496 (N_17496,N_14340,N_14654);
or U17497 (N_17497,N_14602,N_13098);
or U17498 (N_17498,N_14583,N_14152);
nand U17499 (N_17499,N_13158,N_13203);
xnor U17500 (N_17500,N_16403,N_15469);
nor U17501 (N_17501,N_17334,N_16652);
xor U17502 (N_17502,N_15705,N_15527);
nand U17503 (N_17503,N_15007,N_15140);
and U17504 (N_17504,N_17027,N_15202);
or U17505 (N_17505,N_15882,N_15937);
nor U17506 (N_17506,N_15994,N_15358);
xnor U17507 (N_17507,N_17168,N_17443);
xnor U17508 (N_17508,N_17242,N_17088);
or U17509 (N_17509,N_16214,N_15460);
xor U17510 (N_17510,N_15100,N_16309);
nor U17511 (N_17511,N_16137,N_16932);
and U17512 (N_17512,N_16730,N_17348);
nor U17513 (N_17513,N_17497,N_15655);
or U17514 (N_17514,N_15539,N_17092);
nand U17515 (N_17515,N_15292,N_17437);
nand U17516 (N_17516,N_16078,N_15636);
xor U17517 (N_17517,N_16820,N_17248);
nand U17518 (N_17518,N_15331,N_15870);
nand U17519 (N_17519,N_16866,N_15454);
xor U17520 (N_17520,N_17152,N_16639);
and U17521 (N_17521,N_16228,N_15429);
or U17522 (N_17522,N_17150,N_17204);
and U17523 (N_17523,N_16509,N_16842);
and U17524 (N_17524,N_15001,N_16011);
nand U17525 (N_17525,N_15376,N_15608);
nor U17526 (N_17526,N_16346,N_15055);
nor U17527 (N_17527,N_17199,N_15000);
xnor U17528 (N_17528,N_15375,N_15715);
xnor U17529 (N_17529,N_15592,N_17421);
or U17530 (N_17530,N_15488,N_16105);
or U17531 (N_17531,N_15582,N_15317);
and U17532 (N_17532,N_15296,N_15524);
and U17533 (N_17533,N_15258,N_16267);
nor U17534 (N_17534,N_15408,N_16771);
and U17535 (N_17535,N_16325,N_16609);
and U17536 (N_17536,N_15840,N_15673);
and U17537 (N_17537,N_16476,N_17144);
xnor U17538 (N_17538,N_15239,N_16173);
nand U17539 (N_17539,N_16254,N_16665);
and U17540 (N_17540,N_16411,N_15401);
nor U17541 (N_17541,N_16717,N_17285);
or U17542 (N_17542,N_17366,N_16538);
nor U17543 (N_17543,N_15976,N_15152);
xnor U17544 (N_17544,N_16149,N_16565);
nand U17545 (N_17545,N_15530,N_16017);
and U17546 (N_17546,N_15738,N_16582);
or U17547 (N_17547,N_16375,N_16579);
nand U17548 (N_17548,N_15628,N_16682);
nand U17549 (N_17549,N_16751,N_17457);
xnor U17550 (N_17550,N_17143,N_15122);
and U17551 (N_17551,N_15023,N_15145);
or U17552 (N_17552,N_16535,N_17371);
and U17553 (N_17553,N_16216,N_15692);
nor U17554 (N_17554,N_17394,N_15506);
nor U17555 (N_17555,N_15158,N_16742);
nor U17556 (N_17556,N_16797,N_15691);
nand U17557 (N_17557,N_15947,N_15323);
xnor U17558 (N_17558,N_17013,N_15373);
and U17559 (N_17559,N_16496,N_15679);
xor U17560 (N_17560,N_16289,N_15371);
xor U17561 (N_17561,N_16436,N_16780);
xnor U17562 (N_17562,N_17139,N_17173);
nor U17563 (N_17563,N_16077,N_16136);
nor U17564 (N_17564,N_15246,N_15726);
nor U17565 (N_17565,N_16855,N_17320);
nand U17566 (N_17566,N_15604,N_15484);
and U17567 (N_17567,N_16186,N_16131);
and U17568 (N_17568,N_16201,N_17131);
xor U17569 (N_17569,N_16259,N_16525);
nand U17570 (N_17570,N_16001,N_15987);
and U17571 (N_17571,N_15393,N_16208);
or U17572 (N_17572,N_15359,N_17191);
nor U17573 (N_17573,N_16757,N_17225);
nand U17574 (N_17574,N_17175,N_15154);
or U17575 (N_17575,N_16659,N_16548);
xnor U17576 (N_17576,N_17309,N_17222);
or U17577 (N_17577,N_16341,N_16898);
and U17578 (N_17578,N_17339,N_15717);
and U17579 (N_17579,N_17435,N_15379);
nor U17580 (N_17580,N_15347,N_16635);
or U17581 (N_17581,N_16069,N_15340);
and U17582 (N_17582,N_15443,N_16809);
nor U17583 (N_17583,N_16927,N_15553);
or U17584 (N_17584,N_16664,N_15517);
or U17585 (N_17585,N_17493,N_16728);
or U17586 (N_17586,N_17432,N_15273);
or U17587 (N_17587,N_15566,N_15234);
or U17588 (N_17588,N_17201,N_15412);
xnor U17589 (N_17589,N_16986,N_15218);
nor U17590 (N_17590,N_16108,N_15805);
and U17591 (N_17591,N_17134,N_15591);
nor U17592 (N_17592,N_17442,N_16115);
nand U17593 (N_17593,N_15561,N_16237);
or U17594 (N_17594,N_15541,N_16860);
nand U17595 (N_17595,N_17369,N_16291);
and U17596 (N_17596,N_15615,N_17426);
or U17597 (N_17597,N_15839,N_16911);
and U17598 (N_17598,N_17261,N_16401);
xor U17599 (N_17599,N_16057,N_16785);
and U17600 (N_17600,N_15330,N_17218);
or U17601 (N_17601,N_15046,N_15851);
or U17602 (N_17602,N_15792,N_17096);
nor U17603 (N_17603,N_15417,N_16451);
nor U17604 (N_17604,N_17087,N_16490);
nand U17605 (N_17605,N_17446,N_17350);
or U17606 (N_17606,N_15776,N_15384);
xnor U17607 (N_17607,N_16389,N_17321);
and U17608 (N_17608,N_16124,N_17060);
or U17609 (N_17609,N_16358,N_16220);
xor U17610 (N_17610,N_15645,N_16592);
nand U17611 (N_17611,N_15303,N_15857);
xor U17612 (N_17612,N_15021,N_15261);
or U17613 (N_17613,N_15377,N_16409);
and U17614 (N_17614,N_17488,N_16891);
xnor U17615 (N_17615,N_15310,N_16487);
xor U17616 (N_17616,N_17280,N_15755);
or U17617 (N_17617,N_16362,N_16079);
xor U17618 (N_17618,N_15022,N_15828);
xnor U17619 (N_17619,N_16407,N_16831);
or U17620 (N_17620,N_16713,N_16394);
nand U17621 (N_17621,N_15821,N_16980);
or U17622 (N_17622,N_15897,N_15436);
nor U17623 (N_17623,N_17351,N_17067);
or U17624 (N_17624,N_15868,N_16942);
or U17625 (N_17625,N_15033,N_15575);
nand U17626 (N_17626,N_16021,N_16469);
and U17627 (N_17627,N_16740,N_16619);
or U17628 (N_17628,N_16307,N_16262);
xor U17629 (N_17629,N_17465,N_17423);
xnor U17630 (N_17630,N_16647,N_15255);
nor U17631 (N_17631,N_15009,N_15298);
nor U17632 (N_17632,N_16963,N_15499);
xnor U17633 (N_17633,N_15954,N_17279);
nor U17634 (N_17634,N_16873,N_17378);
xnor U17635 (N_17635,N_16095,N_16611);
or U17636 (N_17636,N_15067,N_15071);
nor U17637 (N_17637,N_17240,N_17485);
nand U17638 (N_17638,N_17180,N_17386);
xor U17639 (N_17639,N_15574,N_16398);
and U17640 (N_17640,N_16955,N_15518);
and U17641 (N_17641,N_17315,N_17329);
nand U17642 (N_17642,N_15670,N_16002);
nand U17643 (N_17643,N_17030,N_17243);
xnor U17644 (N_17644,N_16848,N_15043);
xor U17645 (N_17645,N_15632,N_16627);
and U17646 (N_17646,N_15779,N_15667);
xor U17647 (N_17647,N_16392,N_16199);
nand U17648 (N_17648,N_17146,N_16205);
and U17649 (N_17649,N_16531,N_16890);
nor U17650 (N_17650,N_15943,N_16143);
xor U17651 (N_17651,N_16031,N_16504);
or U17652 (N_17652,N_15867,N_15559);
and U17653 (N_17653,N_16331,N_16892);
xnor U17654 (N_17654,N_17103,N_16112);
or U17655 (N_17655,N_17238,N_16298);
nand U17656 (N_17656,N_17151,N_16657);
or U17657 (N_17657,N_17031,N_16632);
nor U17658 (N_17658,N_16920,N_17254);
xor U17659 (N_17659,N_16372,N_17129);
xnor U17660 (N_17660,N_17049,N_16580);
and U17661 (N_17661,N_16861,N_15005);
nor U17662 (N_17662,N_16818,N_15528);
nor U17663 (N_17663,N_15849,N_16087);
or U17664 (N_17664,N_16448,N_16871);
nor U17665 (N_17665,N_15453,N_17498);
nand U17666 (N_17666,N_16655,N_15661);
nor U17667 (N_17667,N_17294,N_16889);
nand U17668 (N_17668,N_15911,N_16093);
and U17669 (N_17669,N_17221,N_15537);
and U17670 (N_17670,N_15769,N_16858);
xor U17671 (N_17671,N_16651,N_16577);
or U17672 (N_17672,N_16759,N_15590);
and U17673 (N_17673,N_16200,N_17020);
nand U17674 (N_17674,N_16134,N_15880);
or U17675 (N_17675,N_15759,N_15664);
and U17676 (N_17676,N_16122,N_16425);
or U17677 (N_17677,N_16284,N_16774);
xnor U17678 (N_17678,N_17335,N_15176);
nand U17679 (N_17679,N_16661,N_15611);
xor U17680 (N_17680,N_15569,N_16918);
nand U17681 (N_17681,N_16038,N_16806);
or U17682 (N_17682,N_16943,N_15380);
and U17683 (N_17683,N_16601,N_15749);
or U17684 (N_17684,N_16312,N_17099);
xnor U17685 (N_17685,N_16499,N_16456);
and U17686 (N_17686,N_15707,N_16669);
nor U17687 (N_17687,N_16534,N_16494);
xor U17688 (N_17688,N_15150,N_15980);
or U17689 (N_17689,N_16452,N_15984);
or U17690 (N_17690,N_16917,N_17215);
nor U17691 (N_17691,N_15964,N_16568);
or U17692 (N_17692,N_17082,N_17052);
and U17693 (N_17693,N_17115,N_15985);
and U17694 (N_17694,N_16258,N_15845);
xor U17695 (N_17695,N_15681,N_17272);
and U17696 (N_17696,N_16616,N_16765);
xnor U17697 (N_17697,N_16053,N_17063);
xor U17698 (N_17698,N_16128,N_15822);
and U17699 (N_17699,N_16054,N_15497);
nand U17700 (N_17700,N_15265,N_15638);
xor U17701 (N_17701,N_17072,N_16503);
or U17702 (N_17702,N_16825,N_15625);
and U17703 (N_17703,N_16792,N_17281);
and U17704 (N_17704,N_15061,N_15772);
nand U17705 (N_17705,N_16418,N_16670);
and U17706 (N_17706,N_17035,N_16354);
and U17707 (N_17707,N_15286,N_16060);
xnor U17708 (N_17708,N_16424,N_16996);
and U17709 (N_17709,N_16316,N_16347);
nor U17710 (N_17710,N_15956,N_16731);
and U17711 (N_17711,N_15748,N_16753);
xnor U17712 (N_17712,N_16822,N_15761);
nor U17713 (N_17713,N_17352,N_16073);
nor U17714 (N_17714,N_15040,N_16040);
or U17715 (N_17715,N_17444,N_15864);
xor U17716 (N_17716,N_17205,N_15272);
and U17717 (N_17717,N_15739,N_15220);
and U17718 (N_17718,N_16326,N_15813);
nor U17719 (N_17719,N_15355,N_15235);
nand U17720 (N_17720,N_15902,N_15231);
nand U17721 (N_17721,N_15648,N_15958);
xor U17722 (N_17722,N_15951,N_16790);
xnor U17723 (N_17723,N_17200,N_15843);
nor U17724 (N_17724,N_15971,N_15056);
nor U17725 (N_17725,N_17057,N_16266);
or U17726 (N_17726,N_15421,N_16754);
xor U17727 (N_17727,N_17015,N_17289);
nor U17728 (N_17728,N_16058,N_17210);
xor U17729 (N_17729,N_17490,N_17475);
and U17730 (N_17730,N_15297,N_15419);
xor U17731 (N_17731,N_16546,N_16747);
xor U17732 (N_17732,N_16319,N_15594);
and U17733 (N_17733,N_17086,N_15115);
and U17734 (N_17734,N_16399,N_16877);
nor U17735 (N_17735,N_15847,N_15778);
or U17736 (N_17736,N_15302,N_15498);
or U17737 (N_17737,N_16197,N_15568);
or U17738 (N_17738,N_15439,N_17417);
nor U17739 (N_17739,N_16042,N_16453);
nand U17740 (N_17740,N_15165,N_17036);
and U17741 (N_17741,N_15058,N_16374);
or U17742 (N_17742,N_17085,N_17479);
nand U17743 (N_17743,N_15836,N_16438);
xnor U17744 (N_17744,N_15117,N_16250);
nor U17745 (N_17745,N_15932,N_16636);
or U17746 (N_17746,N_16193,N_16246);
and U17747 (N_17747,N_16683,N_16332);
nor U17748 (N_17748,N_15136,N_15685);
nand U17749 (N_17749,N_15642,N_16221);
xor U17750 (N_17750,N_15113,N_17398);
or U17751 (N_17751,N_15182,N_16239);
nor U17752 (N_17752,N_15363,N_15786);
or U17753 (N_17753,N_15700,N_17239);
nor U17754 (N_17754,N_15844,N_16648);
and U17755 (N_17755,N_15941,N_15307);
nor U17756 (N_17756,N_17392,N_16823);
and U17757 (N_17757,N_16151,N_15088);
nor U17758 (N_17758,N_15074,N_15390);
xnor U17759 (N_17759,N_16204,N_17109);
or U17760 (N_17760,N_16559,N_17381);
xnor U17761 (N_17761,N_16182,N_17356);
xor U17762 (N_17762,N_15394,N_16313);
or U17763 (N_17763,N_15752,N_16213);
nand U17764 (N_17764,N_16646,N_16096);
or U17765 (N_17765,N_17193,N_16793);
and U17766 (N_17766,N_16882,N_15585);
nand U17767 (N_17767,N_15381,N_16899);
nand U17768 (N_17768,N_16853,N_17445);
or U17769 (N_17769,N_15190,N_17301);
nor U17770 (N_17770,N_15827,N_16830);
nand U17771 (N_17771,N_16714,N_16879);
or U17772 (N_17772,N_16119,N_17171);
nand U17773 (N_17773,N_15669,N_16689);
nand U17774 (N_17774,N_16166,N_16457);
nor U17775 (N_17775,N_16643,N_16048);
nor U17776 (N_17776,N_15597,N_15181);
and U17777 (N_17777,N_17383,N_15523);
or U17778 (N_17778,N_17219,N_16344);
xnor U17779 (N_17779,N_16970,N_15038);
xnor U17780 (N_17780,N_16441,N_16737);
xnor U17781 (N_17781,N_15892,N_16290);
nor U17782 (N_17782,N_16365,N_16941);
nand U17783 (N_17783,N_16716,N_15386);
xor U17784 (N_17784,N_15596,N_17075);
and U17785 (N_17785,N_15883,N_16706);
nor U17786 (N_17786,N_16743,N_15874);
xor U17787 (N_17787,N_15565,N_16323);
nand U17788 (N_17788,N_17018,N_15651);
nand U17789 (N_17789,N_16522,N_15988);
or U17790 (N_17790,N_17166,N_15912);
nand U17791 (N_17791,N_16395,N_16090);
and U17792 (N_17792,N_16008,N_15736);
nand U17793 (N_17793,N_16308,N_16019);
or U17794 (N_17794,N_15922,N_17303);
xnor U17795 (N_17795,N_16749,N_15513);
xnor U17796 (N_17796,N_15644,N_16868);
nor U17797 (N_17797,N_16964,N_15192);
nor U17798 (N_17798,N_15720,N_15407);
nand U17799 (N_17799,N_15535,N_17252);
xor U17800 (N_17800,N_17101,N_15175);
nor U17801 (N_17801,N_16458,N_15250);
nand U17802 (N_17802,N_15034,N_15825);
nand U17803 (N_17803,N_17212,N_15699);
or U17804 (N_17804,N_16972,N_16127);
nor U17805 (N_17805,N_17464,N_17042);
or U17806 (N_17806,N_16296,N_16931);
and U17807 (N_17807,N_16520,N_15948);
nor U17808 (N_17808,N_17438,N_16333);
or U17809 (N_17809,N_15169,N_16462);
or U17810 (N_17810,N_16680,N_15831);
and U17811 (N_17811,N_15881,N_16569);
nor U17812 (N_17812,N_16025,N_15756);
xor U17813 (N_17813,N_16514,N_17121);
xnor U17814 (N_17814,N_16612,N_17255);
nor U17815 (N_17815,N_17051,N_16360);
or U17816 (N_17816,N_16814,N_15395);
and U17817 (N_17817,N_16599,N_16243);
xnor U17818 (N_17818,N_15830,N_17056);
nand U17819 (N_17819,N_15826,N_15742);
and U17820 (N_17820,N_15149,N_16653);
nor U17821 (N_17821,N_15975,N_15962);
and U17822 (N_17822,N_15589,N_16832);
or U17823 (N_17823,N_16450,N_17170);
or U17824 (N_17824,N_16234,N_15352);
xnor U17825 (N_17825,N_17288,N_15986);
xnor U17826 (N_17826,N_16413,N_16685);
nor U17827 (N_17827,N_15556,N_15914);
xnor U17828 (N_17828,N_16356,N_16283);
and U17829 (N_17829,N_16808,N_16746);
xnor U17830 (N_17830,N_16106,N_15799);
nor U17831 (N_17831,N_16795,N_16431);
xnor U17832 (N_17832,N_16739,N_15509);
or U17833 (N_17833,N_16480,N_15650);
and U17834 (N_17834,N_16965,N_17265);
nand U17835 (N_17835,N_16063,N_15318);
nand U17836 (N_17836,N_16410,N_16439);
and U17837 (N_17837,N_17141,N_15946);
and U17838 (N_17838,N_15133,N_15570);
nor U17839 (N_17839,N_17062,N_15078);
nor U17840 (N_17840,N_16187,N_15745);
and U17841 (N_17841,N_16997,N_16429);
xor U17842 (N_17842,N_17157,N_17275);
nand U17843 (N_17843,N_15913,N_15425);
nor U17844 (N_17844,N_15048,N_16961);
and U17845 (N_17845,N_16082,N_15753);
xor U17846 (N_17846,N_15853,N_15172);
nand U17847 (N_17847,N_17068,N_17244);
nand U17848 (N_17848,N_16172,N_15276);
and U17849 (N_17849,N_15496,N_15368);
or U17850 (N_17850,N_17034,N_15508);
xor U17851 (N_17851,N_17307,N_16257);
xor U17852 (N_17852,N_16519,N_16400);
and U17853 (N_17853,N_15702,N_16727);
nand U17854 (N_17854,N_15737,N_15251);
nor U17855 (N_17855,N_15468,N_16273);
and U17856 (N_17856,N_16282,N_16036);
nor U17857 (N_17857,N_15901,N_16687);
xor U17858 (N_17858,N_15979,N_16287);
or U17859 (N_17859,N_17379,N_16238);
nand U17860 (N_17860,N_15014,N_15919);
xnor U17861 (N_17861,N_16386,N_15734);
and U17862 (N_17862,N_16440,N_16009);
and U17863 (N_17863,N_15112,N_17404);
nor U17864 (N_17864,N_15928,N_16274);
nor U17865 (N_17865,N_15185,N_15798);
xnor U17866 (N_17866,N_15435,N_15969);
nor U17867 (N_17867,N_16378,N_15059);
or U17868 (N_17868,N_15199,N_16966);
or U17869 (N_17869,N_15442,N_17290);
xnor U17870 (N_17870,N_16894,N_16623);
nand U17871 (N_17871,N_15540,N_15131);
or U17872 (N_17872,N_15212,N_16366);
and U17873 (N_17873,N_16761,N_17026);
or U17874 (N_17874,N_16851,N_17226);
and U17875 (N_17875,N_15787,N_17196);
xnor U17876 (N_17876,N_17153,N_15624);
nand U17877 (N_17877,N_16248,N_16596);
nand U17878 (N_17878,N_15557,N_16232);
or U17879 (N_17879,N_17232,N_16255);
xor U17880 (N_17880,N_16581,N_16428);
and U17881 (N_17881,N_16024,N_17282);
nor U17882 (N_17882,N_16505,N_17111);
or U17883 (N_17883,N_17078,N_16773);
and U17884 (N_17884,N_15507,N_15832);
or U17885 (N_17885,N_15316,N_15221);
and U17886 (N_17886,N_15094,N_16799);
nand U17887 (N_17887,N_16244,N_15188);
and U17888 (N_17888,N_16045,N_16098);
or U17889 (N_17889,N_15909,N_17390);
or U17890 (N_17890,N_16062,N_15287);
nand U17891 (N_17891,N_16498,N_15025);
and U17892 (N_17892,N_16107,N_16071);
xnor U17893 (N_17893,N_15965,N_17331);
and U17894 (N_17894,N_16829,N_15135);
and U17895 (N_17895,N_16992,N_16593);
xnor U17896 (N_17896,N_16828,N_15719);
xnor U17897 (N_17897,N_15977,N_16926);
nand U17898 (N_17898,N_16159,N_16555);
nor U17899 (N_17899,N_16276,N_15629);
nand U17900 (N_17900,N_16776,N_15503);
and U17901 (N_17901,N_16702,N_16109);
nor U17902 (N_17902,N_15917,N_15634);
nand U17903 (N_17903,N_16195,N_16461);
and U17904 (N_17904,N_17364,N_16603);
nor U17905 (N_17905,N_16583,N_15938);
nand U17906 (N_17906,N_16959,N_15333);
xor U17907 (N_17907,N_15328,N_15440);
xor U17908 (N_17908,N_16174,N_17066);
nor U17909 (N_17909,N_15906,N_17208);
and U17910 (N_17910,N_15254,N_15348);
xor U17911 (N_17911,N_15536,N_15019);
or U17912 (N_17912,N_16065,N_16876);
or U17913 (N_17913,N_17337,N_16999);
and U17914 (N_17914,N_15249,N_15065);
nor U17915 (N_17915,N_16540,N_16263);
and U17916 (N_17916,N_15583,N_16321);
xor U17917 (N_17917,N_16377,N_17106);
nor U17918 (N_17918,N_16495,N_16536);
xnor U17919 (N_17919,N_15259,N_15993);
xnor U17920 (N_17920,N_15683,N_15186);
nor U17921 (N_17921,N_17287,N_17105);
xor U17922 (N_17922,N_15751,N_16382);
or U17923 (N_17923,N_17164,N_16181);
xor U17924 (N_17924,N_16541,N_15807);
xor U17925 (N_17925,N_15674,N_17041);
or U17926 (N_17926,N_17341,N_15433);
or U17927 (N_17927,N_15837,N_16268);
or U17928 (N_17928,N_15978,N_15070);
xor U17929 (N_17929,N_16473,N_15162);
and U17930 (N_17930,N_17418,N_15099);
or U17931 (N_17931,N_17305,N_15184);
nand U17932 (N_17932,N_15411,N_16950);
nor U17933 (N_17933,N_15613,N_17167);
nand U17934 (N_17934,N_16352,N_15918);
xor U17935 (N_17935,N_15052,N_17274);
nand U17936 (N_17936,N_15290,N_16976);
xnor U17937 (N_17937,N_16253,N_15427);
or U17938 (N_17938,N_16606,N_16421);
or U17939 (N_17939,N_16769,N_17393);
xnor U17940 (N_17940,N_17100,N_16013);
and U17941 (N_17941,N_16081,N_15444);
and U17942 (N_17942,N_17223,N_15179);
or U17943 (N_17943,N_16697,N_17207);
nor U17944 (N_17944,N_16113,N_15542);
or U17945 (N_17945,N_16838,N_17028);
xor U17946 (N_17946,N_15723,N_15081);
nand U17947 (N_17947,N_16711,N_16154);
and U17948 (N_17948,N_16722,N_17293);
or U17949 (N_17949,N_16417,N_16190);
and U17950 (N_17950,N_15612,N_15775);
xor U17951 (N_17951,N_16383,N_16217);
and U17952 (N_17952,N_15223,N_15266);
or U17953 (N_17953,N_15662,N_17420);
nor U17954 (N_17954,N_15126,N_17247);
and U17955 (N_17955,N_16138,N_16049);
and U17956 (N_17956,N_16130,N_17388);
and U17957 (N_17957,N_16833,N_15972);
nor U17958 (N_17958,N_15233,N_17108);
nand U17959 (N_17959,N_17433,N_15973);
xor U17960 (N_17960,N_15332,N_17136);
and U17961 (N_17961,N_15168,N_15877);
xor U17962 (N_17962,N_15195,N_15130);
and U17963 (N_17963,N_16223,N_16218);
xnor U17964 (N_17964,N_17396,N_16416);
and U17965 (N_17965,N_15129,N_17298);
nor U17966 (N_17966,N_16967,N_15087);
and U17967 (N_17967,N_16988,N_15031);
nor U17968 (N_17968,N_15326,N_16721);
or U17969 (N_17969,N_16072,N_16311);
or U17970 (N_17970,N_16618,N_16317);
nor U17971 (N_17971,N_16293,N_16068);
and U17972 (N_17972,N_16445,N_17271);
or U17973 (N_17973,N_15462,N_16849);
xor U17974 (N_17974,N_16844,N_16630);
and U17975 (N_17975,N_15716,N_15047);
nand U17976 (N_17976,N_15207,N_16471);
or U17977 (N_17977,N_17332,N_16245);
and U17978 (N_17978,N_16951,N_16092);
or U17979 (N_17979,N_16513,N_15698);
nor U17980 (N_17980,N_15114,N_15802);
nand U17981 (N_17981,N_16598,N_16867);
and U17982 (N_17982,N_15603,N_15029);
xnor U17983 (N_17983,N_16962,N_15529);
xor U17984 (N_17984,N_16314,N_16361);
nand U17985 (N_17985,N_15438,N_16207);
nand U17986 (N_17986,N_16376,N_15500);
nand U17987 (N_17987,N_15456,N_15110);
or U17988 (N_17988,N_15105,N_16933);
and U17989 (N_17989,N_16497,N_17165);
or U17990 (N_17990,N_16168,N_17033);
nand U17991 (N_17991,N_17128,N_16800);
or U17992 (N_17992,N_15708,N_15607);
nor U17993 (N_17993,N_16121,N_15295);
and U17994 (N_17994,N_16016,N_15713);
xnor U17995 (N_17995,N_17074,N_17330);
xor U17996 (N_17996,N_15405,N_15731);
or U17997 (N_17997,N_17029,N_16297);
or U17998 (N_17998,N_16415,N_16954);
xor U17999 (N_17999,N_15610,N_15278);
nor U18000 (N_18000,N_17159,N_16805);
nor U18001 (N_18001,N_16788,N_16123);
nand U18002 (N_18002,N_15855,N_17227);
nor U18003 (N_18003,N_16798,N_16945);
xnor U18004 (N_18004,N_16444,N_15640);
or U18005 (N_18005,N_15658,N_16865);
nor U18006 (N_18006,N_16949,N_15534);
xor U18007 (N_18007,N_15346,N_16100);
or U18008 (N_18008,N_17185,N_16704);
nor U18009 (N_18009,N_15092,N_17094);
nor U18010 (N_18010,N_17220,N_17300);
or U18011 (N_18011,N_16171,N_16883);
and U18012 (N_18012,N_17499,N_16625);
nand U18013 (N_18013,N_16481,N_16396);
xor U18014 (N_18014,N_16156,N_15997);
or U18015 (N_18015,N_16897,N_17048);
and U18016 (N_18016,N_15201,N_16059);
or U18017 (N_18017,N_16247,N_16139);
nor U18018 (N_18018,N_15525,N_15865);
nand U18019 (N_18019,N_15230,N_16940);
and U18020 (N_18020,N_16050,N_17478);
or U18021 (N_18021,N_16703,N_15577);
xor U18022 (N_18022,N_17081,N_17452);
nand U18023 (N_18023,N_15372,N_15784);
or U18024 (N_18024,N_15863,N_15350);
nor U18025 (N_18025,N_15817,N_15064);
nand U18026 (N_18026,N_17380,N_17473);
nand U18027 (N_18027,N_15336,N_15815);
or U18028 (N_18028,N_15725,N_17477);
nand U18029 (N_18029,N_16745,N_15367);
and U18030 (N_18030,N_17043,N_16786);
nor U18031 (N_18031,N_15121,N_16299);
and U18032 (N_18032,N_16720,N_15974);
xor U18033 (N_18033,N_16908,N_15665);
and U18034 (N_18034,N_16506,N_16552);
nand U18035 (N_18035,N_17245,N_15396);
or U18036 (N_18036,N_17310,N_17313);
and U18037 (N_18037,N_15887,N_15319);
nor U18038 (N_18038,N_16169,N_15875);
and U18039 (N_18039,N_16930,N_15531);
nor U18040 (N_18040,N_15485,N_16859);
and U18041 (N_18041,N_15229,N_16000);
nand U18042 (N_18042,N_15079,N_15649);
nor U18043 (N_18043,N_16750,N_15512);
or U18044 (N_18044,N_17342,N_16732);
and U18045 (N_18045,N_15489,N_16455);
nor U18046 (N_18046,N_15155,N_15942);
nand U18047 (N_18047,N_16815,N_17323);
nand U18048 (N_18048,N_16944,N_15818);
nor U18049 (N_18049,N_16590,N_15406);
xnor U18050 (N_18050,N_16188,N_15890);
nor U18051 (N_18051,N_16391,N_16523);
nor U18052 (N_18052,N_17419,N_16226);
nor U18053 (N_18053,N_16155,N_16957);
and U18054 (N_18054,N_15795,N_17229);
or U18055 (N_18055,N_16281,N_15285);
nor U18056 (N_18056,N_15174,N_17104);
xor U18057 (N_18057,N_16304,N_17353);
nor U18058 (N_18058,N_17489,N_16663);
nor U18059 (N_18059,N_17314,N_15567);
and U18060 (N_18060,N_17070,N_17431);
or U18061 (N_18061,N_16435,N_16694);
nor U18062 (N_18062,N_16758,N_15511);
nor U18063 (N_18063,N_15089,N_15491);
nor U18064 (N_18064,N_16210,N_15322);
or U18065 (N_18065,N_16938,N_17156);
nand U18066 (N_18066,N_15687,N_16474);
nand U18067 (N_18067,N_17284,N_17080);
or U18068 (N_18068,N_16693,N_15486);
or U18069 (N_18069,N_16686,N_16576);
or U18070 (N_18070,N_16554,N_16175);
or U18071 (N_18071,N_17359,N_16483);
nand U18072 (N_18072,N_15467,N_16550);
or U18073 (N_18073,N_15659,N_16690);
or U18074 (N_18074,N_16044,N_16709);
xor U18075 (N_18075,N_16126,N_17237);
or U18076 (N_18076,N_15116,N_15247);
xnor U18077 (N_18077,N_15730,N_15492);
nor U18078 (N_18078,N_16251,N_15431);
nand U18079 (N_18079,N_16629,N_16432);
and U18080 (N_18080,N_16227,N_15086);
and U18081 (N_18081,N_17148,N_16684);
xor U18082 (N_18082,N_16637,N_15324);
or U18083 (N_18083,N_15045,N_16230);
or U18084 (N_18084,N_17361,N_17058);
nor U18085 (N_18085,N_16140,N_15068);
nand U18086 (N_18086,N_15360,N_16787);
nor U18087 (N_18087,N_15312,N_15620);
nor U18088 (N_18088,N_15950,N_16604);
nor U18089 (N_18089,N_15036,N_15013);
nor U18090 (N_18090,N_15671,N_17095);
nor U18091 (N_18091,N_15037,N_16286);
or U18092 (N_18092,N_16982,N_16236);
nand U18093 (N_18093,N_16922,N_15676);
or U18094 (N_18094,N_17069,N_16192);
or U18095 (N_18095,N_17194,N_16114);
xnor U18096 (N_18096,N_15107,N_16974);
xor U18097 (N_18097,N_16152,N_17198);
nand U18098 (N_18098,N_17482,N_17117);
xor U18099 (N_18099,N_17114,N_15501);
or U18100 (N_18100,N_16734,N_15688);
xor U18101 (N_18101,N_16544,N_17195);
xnor U18102 (N_18102,N_16085,N_16766);
or U18103 (N_18103,N_17188,N_16224);
or U18104 (N_18104,N_15672,N_16367);
nand U18105 (N_18105,N_15128,N_17411);
and U18106 (N_18106,N_16671,N_16390);
or U18107 (N_18107,N_15160,N_15504);
xnor U18108 (N_18108,N_15378,N_15595);
and U18109 (N_18109,N_15284,N_16640);
and U18110 (N_18110,N_17257,N_16330);
and U18111 (N_18111,N_15224,N_16755);
or U18112 (N_18112,N_16222,N_15441);
nand U18113 (N_18113,N_15183,N_17453);
or U18114 (N_18114,N_15757,N_16198);
and U18115 (N_18115,N_15876,N_15794);
and U18116 (N_18116,N_16952,N_16294);
nand U18117 (N_18117,N_16909,N_15095);
and U18118 (N_18118,N_16558,N_15908);
nor U18119 (N_18119,N_15647,N_17365);
or U18120 (N_18120,N_16161,N_16512);
xor U18121 (N_18121,N_16878,N_15552);
and U18122 (N_18122,N_16574,N_17316);
nand U18123 (N_18123,N_15690,N_16280);
nor U18124 (N_18124,N_15006,N_16666);
xor U18125 (N_18125,N_16705,N_16212);
nand U18126 (N_18126,N_15850,N_16995);
or U18127 (N_18127,N_15189,N_16929);
nor U18128 (N_18128,N_16783,N_16179);
xnor U18129 (N_18129,N_15814,N_16014);
and U18130 (N_18130,N_15364,N_16427);
xnor U18131 (N_18131,N_15008,N_15341);
and U18132 (N_18132,N_16695,N_15983);
nor U18133 (N_18133,N_16470,N_17064);
xnor U18134 (N_18134,N_17250,N_16960);
nand U18135 (N_18135,N_16782,N_16948);
xnor U18136 (N_18136,N_15245,N_16673);
nor U18137 (N_18137,N_16412,N_15996);
nor U18138 (N_18138,N_16784,N_15637);
or U18139 (N_18139,N_17079,N_15098);
or U18140 (N_18140,N_17262,N_15762);
xor U18141 (N_18141,N_15859,N_16338);
nand U18142 (N_18142,N_15093,N_17090);
nor U18143 (N_18143,N_15766,N_17328);
and U18144 (N_18144,N_16925,N_16772);
or U18145 (N_18145,N_16379,N_16340);
nand U18146 (N_18146,N_16863,N_17135);
and U18147 (N_18147,N_15196,N_16339);
nand U18148 (N_18148,N_16353,N_15617);
and U18149 (N_18149,N_15907,N_16994);
and U18150 (N_18150,N_16030,N_15473);
or U18151 (N_18151,N_15694,N_16562);
or U18152 (N_18152,N_15895,N_16501);
xnor U18153 (N_18153,N_15633,N_17358);
nor U18154 (N_18154,N_16370,N_15487);
xor U18155 (N_18155,N_15306,N_15082);
and U18156 (N_18156,N_15641,N_17091);
or U18157 (N_18157,N_15198,N_15414);
xnor U18158 (N_18158,N_16420,N_16384);
or U18159 (N_18159,N_15933,N_16895);
xor U18160 (N_18160,N_16888,N_16385);
xor U18161 (N_18161,N_17344,N_16012);
and U18162 (N_18162,N_15146,N_15402);
nand U18163 (N_18163,N_15173,N_15810);
and U18164 (N_18164,N_17256,N_16368);
nand U18165 (N_18165,N_16404,N_16811);
xor U18166 (N_18166,N_16479,N_15271);
and U18167 (N_18167,N_17206,N_17133);
and U18168 (N_18168,N_16572,N_16147);
and U18169 (N_18169,N_15957,N_16229);
nand U18170 (N_18170,N_15780,N_16668);
xnor U18171 (N_18171,N_15765,N_16781);
nand U18172 (N_18172,N_15243,N_16373);
and U18173 (N_18173,N_16594,N_15461);
xor U18174 (N_18174,N_16904,N_16906);
or U18175 (N_18175,N_15714,N_16145);
xnor U18176 (N_18176,N_16560,N_16464);
or U18177 (N_18177,N_15516,N_15208);
nand U18178 (N_18178,N_17299,N_15558);
xnor U18179 (N_18179,N_16348,N_16981);
xor U18180 (N_18180,N_17406,N_16408);
or U18181 (N_18181,N_17161,N_17055);
and U18182 (N_18182,N_16277,N_16973);
nor U18183 (N_18183,N_17044,N_15383);
xor U18184 (N_18184,N_16857,N_15598);
and U18185 (N_18185,N_15833,N_17140);
xnor U18186 (N_18186,N_16887,N_15927);
nand U18187 (N_18187,N_15820,N_17495);
nand U18188 (N_18188,N_16342,N_16153);
or U18189 (N_18189,N_17414,N_17428);
xor U18190 (N_18190,N_15652,N_16029);
xor U18191 (N_18191,N_17410,N_16422);
and U18192 (N_18192,N_17116,N_17228);
nand U18193 (N_18193,N_17107,N_15788);
and U18194 (N_18194,N_15361,N_17021);
nor U18195 (N_18195,N_16946,N_15018);
and U18196 (N_18196,N_15063,N_16320);
xor U18197 (N_18197,N_15522,N_16443);
nor U18198 (N_18198,N_16032,N_15370);
or U18199 (N_18199,N_16055,N_16023);
or U18200 (N_18200,N_16423,N_15343);
or U18201 (N_18201,N_15657,N_16380);
nand U18202 (N_18202,N_16148,N_15538);
xor U18203 (N_18203,N_15357,N_16595);
and U18204 (N_18204,N_16511,N_16300);
nand U18205 (N_18205,N_15413,N_15123);
or U18206 (N_18206,N_17130,N_15959);
nand U18207 (N_18207,N_15619,N_17311);
or U18208 (N_18208,N_15228,N_16936);
or U18209 (N_18209,N_16700,N_15900);
and U18210 (N_18210,N_16900,N_15623);
nand U18211 (N_18211,N_17496,N_17373);
nand U18212 (N_18212,N_17259,N_15746);
and U18213 (N_18213,N_15300,N_16066);
or U18214 (N_18214,N_16588,N_16834);
and U18215 (N_18215,N_15365,N_15869);
or U18216 (N_18216,N_16419,N_15403);
nand U18217 (N_18217,N_15069,N_16270);
xor U18218 (N_18218,N_15995,N_15311);
xnor U18219 (N_18219,N_16209,N_17125);
nor U18220 (N_18220,N_16261,N_15423);
and U18221 (N_18221,N_16760,N_16135);
and U18222 (N_18222,N_16807,N_16035);
and U18223 (N_18223,N_16821,N_15621);
nand U18224 (N_18224,N_17407,N_17137);
nand U18225 (N_18225,N_17241,N_16968);
xnor U18226 (N_18226,N_16295,N_17395);
nor U18227 (N_18227,N_16144,N_16796);
xnor U18228 (N_18228,N_16364,N_16841);
and U18229 (N_18229,N_16624,N_16020);
xnor U18230 (N_18230,N_15464,N_16816);
and U18231 (N_18231,N_16658,N_15819);
nor U18232 (N_18232,N_15680,N_15695);
nor U18233 (N_18233,N_17450,N_15533);
or U18234 (N_18234,N_17336,N_15515);
nand U18235 (N_18235,N_16846,N_15675);
nand U18236 (N_18236,N_15432,N_15342);
or U18237 (N_18237,N_17469,N_15187);
and U18238 (N_18238,N_15144,N_15521);
xor U18239 (N_18239,N_16542,N_15770);
and U18240 (N_18240,N_16978,N_15242);
nor U18241 (N_18241,N_15686,N_15550);
nor U18242 (N_18242,N_15967,N_15280);
or U18243 (N_18243,N_15344,N_17382);
and U18244 (N_18244,N_16870,N_15472);
and U18245 (N_18245,N_15451,N_16862);
xnor U18246 (N_18246,N_16827,N_15106);
or U18247 (N_18247,N_16465,N_17391);
xor U18248 (N_18248,N_17375,N_16285);
xnor U18249 (N_18249,N_16791,N_15796);
nor U18250 (N_18250,N_16028,N_16589);
xor U18251 (N_18251,N_15510,N_15580);
nand U18252 (N_18252,N_17354,N_15862);
nor U18253 (N_18253,N_16345,N_16489);
or U18254 (N_18254,N_15711,N_17397);
xor U18255 (N_18255,N_16724,N_17474);
or U18256 (N_18256,N_17054,N_15109);
and U18257 (N_18257,N_16163,N_16613);
or U18258 (N_18258,N_15899,N_15614);
xor U18259 (N_18259,N_16905,N_16094);
nand U18260 (N_18260,N_16076,N_16916);
nor U18261 (N_18261,N_16708,N_16667);
xnor U18262 (N_18262,N_15744,N_15777);
xnor U18263 (N_18263,N_17374,N_16676);
xnor U18264 (N_18264,N_17076,N_15945);
xor U18265 (N_18265,N_16363,N_17045);
nor U18266 (N_18266,N_16305,N_17278);
and U18267 (N_18267,N_15709,N_16493);
nand U18268 (N_18268,N_15459,N_16710);
xnor U18269 (N_18269,N_15041,N_17008);
nand U18270 (N_18270,N_17363,N_15156);
xor U18271 (N_18271,N_17186,N_16587);
or U18272 (N_18272,N_15422,N_16203);
and U18273 (N_18273,N_17447,N_15502);
nand U18274 (N_18274,N_16650,N_16913);
nor U18275 (N_18275,N_16041,N_15313);
xor U18276 (N_18276,N_15545,N_15931);
or U18277 (N_18277,N_16748,N_17126);
nor U18278 (N_18278,N_15345,N_15269);
xor U18279 (N_18279,N_15547,N_17047);
nand U18280 (N_18280,N_17470,N_15118);
or U18281 (N_18281,N_17142,N_16924);
and U18282 (N_18282,N_15327,N_15238);
xnor U18283 (N_18283,N_15076,N_16712);
or U18284 (N_18284,N_17038,N_17440);
and U18285 (N_18285,N_17408,N_15463);
nor U18286 (N_18286,N_16269,N_15111);
nand U18287 (N_18287,N_15856,N_17462);
nor U18288 (N_18288,N_15428,N_17160);
and U18289 (N_18289,N_15147,N_16585);
nor U18290 (N_18290,N_17183,N_17273);
nor U18291 (N_18291,N_17295,N_16884);
nand U18292 (N_18292,N_17024,N_16804);
xnor U18293 (N_18293,N_16459,N_15584);
xor U18294 (N_18294,N_17184,N_16477);
nor U18295 (N_18295,N_15213,N_15693);
and U18296 (N_18296,N_15119,N_15834);
nand U18297 (N_18297,N_15434,N_16817);
or U18298 (N_18298,N_15476,N_16051);
nor U18299 (N_18299,N_16919,N_17177);
or U18300 (N_18300,N_17327,N_15314);
xor U18301 (N_18301,N_16303,N_15733);
or U18302 (N_18302,N_16064,N_15409);
nand U18303 (N_18303,N_16117,N_17399);
or U18304 (N_18304,N_16767,N_16644);
nand U18305 (N_18305,N_16993,N_15003);
nor U18306 (N_18306,N_17025,N_15102);
nand U18307 (N_18307,N_15399,N_15325);
or U18308 (N_18308,N_17124,N_15410);
nor U18309 (N_18309,N_16132,N_15823);
and U18310 (N_18310,N_16046,N_16843);
or U18311 (N_18311,N_15493,N_17120);
nand U18312 (N_18312,N_17268,N_15703);
or U18313 (N_18313,N_16775,N_15354);
and U18314 (N_18314,N_15470,N_16160);
nor U18315 (N_18315,N_17347,N_17384);
and U18316 (N_18316,N_16634,N_15562);
and U18317 (N_18317,N_15563,N_16158);
nor U18318 (N_18318,N_17197,N_16414);
nor U18319 (N_18319,N_15809,N_16921);
nor U18320 (N_18320,N_15701,N_16545);
and U18321 (N_18321,N_15137,N_17234);
xnor U18322 (N_18322,N_16633,N_16642);
xor U18323 (N_18323,N_16164,N_15054);
nor U18324 (N_18324,N_17235,N_16812);
nand U18325 (N_18325,N_17097,N_17118);
nor U18326 (N_18326,N_15177,N_16901);
and U18327 (N_18327,N_15012,N_17004);
nor U18328 (N_18328,N_17270,N_16875);
and U18329 (N_18329,N_15952,N_15631);
nor U18330 (N_18330,N_15543,N_15315);
nand U18331 (N_18331,N_17266,N_17325);
nand U18332 (N_18332,N_17296,N_15712);
nor U18333 (N_18333,N_15334,N_15635);
xnor U18334 (N_18334,N_16492,N_16983);
and U18335 (N_18335,N_17376,N_16947);
and U18336 (N_18336,N_15935,N_15279);
xnor U18337 (N_18337,N_16764,N_16406);
xor U18338 (N_18338,N_17413,N_15389);
and U18339 (N_18339,N_16524,N_16770);
nand U18340 (N_18340,N_16165,N_15781);
nor U18341 (N_18341,N_16310,N_15727);
xor U18342 (N_18342,N_16327,N_16662);
nand U18343 (N_18343,N_16869,N_17224);
xnor U18344 (N_18344,N_17147,N_16537);
xor U18345 (N_18345,N_17217,N_17145);
xor U18346 (N_18346,N_15760,N_17277);
nor U18347 (N_18347,N_16824,N_16631);
and U18348 (N_18348,N_15171,N_16488);
nand U18349 (N_18349,N_16211,N_16252);
and U18350 (N_18350,N_15127,N_15894);
and U18351 (N_18351,N_15573,N_15896);
nor U18352 (N_18352,N_16910,N_16956);
nor U18353 (N_18353,N_15066,N_15939);
nor U18354 (N_18354,N_17324,N_17010);
nand U18355 (N_18355,N_15926,N_16975);
nor U18356 (N_18356,N_17154,N_15609);
or U18357 (N_18357,N_16672,N_16037);
and U18358 (N_18358,N_17061,N_15010);
nor U18359 (N_18359,N_15773,N_16102);
or U18360 (N_18360,N_17326,N_15288);
xnor U18361 (N_18361,N_15458,N_16191);
and U18362 (N_18362,N_16070,N_15206);
and U18363 (N_18363,N_15758,N_16442);
and U18364 (N_18364,N_16756,N_15049);
xnor U18365 (N_18365,N_17456,N_16675);
and U18366 (N_18366,N_16741,N_15846);
nand U18367 (N_18367,N_17037,N_17360);
and U18368 (N_18368,N_17089,N_17040);
or U18369 (N_18369,N_16736,N_16953);
or U18370 (N_18370,N_16231,N_15885);
nor U18371 (N_18371,N_15077,N_16515);
xor U18372 (N_18372,N_17211,N_15743);
nor U18373 (N_18373,N_16826,N_17182);
and U18374 (N_18374,N_16696,N_15858);
and U18375 (N_18375,N_16454,N_15588);
nor U18376 (N_18376,N_16052,N_15252);
or U18377 (N_18377,N_15546,N_15949);
or U18378 (N_18378,N_17163,N_16608);
or U18379 (N_18379,N_15167,N_16185);
nor U18380 (N_18380,N_16005,N_16349);
nand U18381 (N_18381,N_16485,N_15889);
and U18382 (N_18382,N_15741,N_16864);
and U18383 (N_18383,N_17346,N_17427);
nand U18384 (N_18384,N_16516,N_16854);
nand U18385 (N_18385,N_16845,N_16621);
nand U18386 (N_18386,N_15134,N_16835);
nor U18387 (N_18387,N_15481,N_16729);
nand U18388 (N_18388,N_15554,N_15002);
xor U18389 (N_18389,N_16083,N_16551);
nand U18390 (N_18390,N_15842,N_15921);
or U18391 (N_18391,N_16170,N_15981);
xnor U18392 (N_18392,N_15886,N_16111);
or U18393 (N_18393,N_15936,N_17127);
nand U18394 (N_18394,N_15578,N_15191);
nand U18395 (N_18395,N_16116,N_17377);
or U18396 (N_18396,N_15905,N_16810);
or U18397 (N_18397,N_16004,N_15268);
and U18398 (N_18398,N_15480,N_15852);
or U18399 (N_18399,N_15477,N_16486);
or U18400 (N_18400,N_15955,N_17001);
and U18401 (N_18401,N_16564,N_15349);
nand U18402 (N_18402,N_17138,N_15044);
and U18403 (N_18403,N_15989,N_15968);
and U18404 (N_18404,N_17455,N_16433);
xor U18405 (N_18405,N_15204,N_15970);
or U18406 (N_18406,N_16977,N_15020);
xor U18407 (N_18407,N_15482,N_15599);
xnor U18408 (N_18408,N_16369,N_15446);
nand U18409 (N_18409,N_16539,N_17005);
xor U18410 (N_18410,N_15240,N_15763);
nor U18411 (N_18411,N_16874,N_15264);
nand U18412 (N_18412,N_15353,N_15581);
nor U18413 (N_18413,N_15024,N_15448);
nand U18414 (N_18414,N_15387,N_15138);
nand U18415 (N_18415,N_17461,N_16607);
or U18416 (N_18416,N_16003,N_16990);
nand U18417 (N_18417,N_15124,N_15706);
and U18418 (N_18418,N_15990,N_15244);
xor U18419 (N_18419,N_16803,N_15768);
nand U18420 (N_18420,N_15888,N_16638);
or U18421 (N_18421,N_15564,N_15028);
and U18422 (N_18422,N_15689,N_15337);
nand U18423 (N_18423,N_17439,N_15728);
nor U18424 (N_18424,N_15260,N_17459);
nand U18425 (N_18425,N_15848,N_15193);
nor U18426 (N_18426,N_16067,N_15872);
and U18427 (N_18427,N_15283,N_17110);
and U18428 (N_18428,N_16813,N_15060);
nand U18429 (N_18429,N_17430,N_16691);
or U18430 (N_18430,N_16194,N_16478);
and U18431 (N_18431,N_16405,N_16260);
nand U18432 (N_18432,N_15940,N_15051);
nand U18433 (N_18433,N_16718,N_15735);
xnor U18434 (N_18434,N_15824,N_15097);
or U18435 (N_18435,N_17480,N_15050);
or U18436 (N_18436,N_15593,N_15618);
or U18437 (N_18437,N_17203,N_15420);
xor U18438 (N_18438,N_16907,N_15215);
and U18439 (N_18439,N_15903,N_15257);
nand U18440 (N_18440,N_16934,N_17494);
or U18441 (N_18441,N_17424,N_17291);
nand U18442 (N_18442,N_16177,N_15771);
nand U18443 (N_18443,N_15576,N_17213);
nor U18444 (N_18444,N_16249,N_16359);
or U18445 (N_18445,N_17190,N_15164);
nor U18446 (N_18446,N_15767,N_15560);
and U18447 (N_18447,N_15248,N_16614);
nand U18448 (N_18448,N_15073,N_16584);
and U18449 (N_18449,N_15630,N_15929);
nand U18450 (N_18450,N_17073,N_17403);
or U18451 (N_18451,N_16101,N_17233);
and U18452 (N_18452,N_17405,N_16089);
nor U18453 (N_18453,N_17415,N_16475);
or U18454 (N_18454,N_16388,N_17181);
nor U18455 (N_18455,N_15015,N_15148);
nand U18456 (N_18456,N_15797,N_15219);
or U18457 (N_18457,N_16533,N_15961);
or U18458 (N_18458,N_17006,N_17400);
or U18459 (N_18459,N_15800,N_16278);
nor U18460 (N_18460,N_17269,N_17416);
nand U18461 (N_18461,N_17322,N_15452);
or U18462 (N_18462,N_16557,N_17162);
nand U18463 (N_18463,N_16397,N_17422);
or U18464 (N_18464,N_16715,N_16034);
nand U18465 (N_18465,N_16180,N_15084);
xnor U18466 (N_18466,N_16328,N_16979);
xor U18467 (N_18467,N_15083,N_15782);
and U18468 (N_18468,N_16225,N_16178);
xnor U18469 (N_18469,N_16641,N_15426);
nand U18470 (N_18470,N_15526,N_17367);
nand U18471 (N_18471,N_16928,N_17486);
nand U18472 (N_18472,N_15299,N_16622);
xnor U18473 (N_18473,N_16393,N_16074);
nand U18474 (N_18474,N_15579,N_16142);
nand U18475 (N_18475,N_17308,N_17017);
nor U18476 (N_18476,N_17158,N_15277);
xnor U18477 (N_18477,N_16794,N_15722);
xnor U18478 (N_18478,N_15294,N_15710);
and U18479 (N_18479,N_16235,N_16104);
nor U18480 (N_18480,N_16256,N_15684);
xnor U18481 (N_18481,N_16206,N_15495);
and U18482 (N_18482,N_16022,N_15289);
or U18483 (N_18483,N_15004,N_15812);
nor U18484 (N_18484,N_16777,N_15339);
nor U18485 (N_18485,N_15682,N_16881);
nand U18486 (N_18486,N_15920,N_16939);
or U18487 (N_18487,N_17123,N_17039);
nor U18488 (N_18488,N_16679,N_16847);
nand U18489 (N_18489,N_15656,N_16043);
nand U18490 (N_18490,N_16605,N_15915);
nor U18491 (N_18491,N_17460,N_15382);
nor U18492 (N_18492,N_16472,N_16402);
xnor U18493 (N_18493,N_16914,N_17345);
nand U18494 (N_18494,N_17016,N_17448);
nand U18495 (N_18495,N_16118,N_17387);
nor U18496 (N_18496,N_16288,N_16306);
xnor U18497 (N_18497,N_17046,N_15571);
nand U18498 (N_18498,N_15811,N_15873);
xor U18499 (N_18499,N_15016,N_15424);
and U18500 (N_18500,N_15281,N_16677);
or U18501 (N_18501,N_15555,N_15465);
nor U18502 (N_18502,N_15494,N_16528);
or U18503 (N_18503,N_15132,N_15398);
xnor U18504 (N_18504,N_15026,N_17318);
nor U18505 (N_18505,N_15934,N_15011);
xor U18506 (N_18506,N_15178,N_15860);
and U18507 (N_18507,N_16726,N_17071);
and U18508 (N_18508,N_15391,N_15108);
and U18509 (N_18509,N_15282,N_16529);
nor U18510 (N_18510,N_15666,N_16880);
nor U18511 (N_18511,N_17260,N_16656);
and U18512 (N_18512,N_17276,N_15320);
and U18513 (N_18513,N_15475,N_15445);
xor U18514 (N_18514,N_16527,N_15450);
nor U18515 (N_18515,N_16162,N_16315);
xnor U18516 (N_18516,N_16324,N_15808);
or U18517 (N_18517,N_16343,N_15214);
nor U18518 (N_18518,N_16437,N_16801);
xnor U18519 (N_18519,N_15274,N_15471);
nand U18520 (N_18520,N_17249,N_16125);
xnor U18521 (N_18521,N_16937,N_17174);
xnor U18522 (N_18522,N_16570,N_16852);
nand U18523 (N_18523,N_15544,N_15879);
xnor U18524 (N_18524,N_15205,N_15548);
nand U18525 (N_18525,N_16563,N_15677);
and U18526 (N_18526,N_17304,N_15474);
xor U18527 (N_18527,N_15729,N_15764);
nand U18528 (N_18528,N_15783,N_17209);
nand U18529 (N_18529,N_16387,N_16329);
nand U18530 (N_18530,N_16196,N_15704);
nor U18531 (N_18531,N_15991,N_17402);
or U18532 (N_18532,N_16091,N_16240);
or U18533 (N_18533,N_17169,N_15263);
and U18534 (N_18534,N_16701,N_16692);
and U18535 (N_18535,N_16381,N_15153);
xor U18536 (N_18536,N_15217,N_15639);
or U18537 (N_18537,N_16215,N_17434);
and U18538 (N_18538,N_15483,N_17441);
nor U18539 (N_18539,N_17009,N_15241);
xor U18540 (N_18540,N_17155,N_15532);
and U18541 (N_18541,N_16674,N_15930);
nand U18542 (N_18542,N_16678,N_16896);
or U18543 (N_18543,N_15740,N_15804);
and U18544 (N_18544,N_17283,N_15035);
nor U18545 (N_18545,N_15893,N_16133);
nor U18546 (N_18546,N_16597,N_15415);
xor U18547 (N_18547,N_15400,N_16157);
and U18548 (N_18548,N_16615,N_15696);
and U18549 (N_18549,N_17251,N_17011);
and U18550 (N_18550,N_17084,N_15587);
or U18551 (N_18551,N_16778,N_15170);
nor U18552 (N_18552,N_15801,N_15057);
and U18553 (N_18553,N_16591,N_15549);
or U18554 (N_18554,N_15678,N_15335);
or U18555 (N_18555,N_16075,N_17149);
or U18556 (N_18556,N_15878,N_15724);
nand U18557 (N_18557,N_15505,N_17317);
and U18558 (N_18558,N_15275,N_17007);
nand U18559 (N_18559,N_16998,N_16334);
or U18560 (N_18560,N_16553,N_15430);
nand U18561 (N_18561,N_16086,N_15600);
or U18562 (N_18562,N_15999,N_17468);
or U18563 (N_18563,N_17202,N_15236);
nor U18564 (N_18564,N_16752,N_16645);
nand U18565 (N_18565,N_17297,N_16120);
or U18566 (N_18566,N_15091,N_17466);
xor U18567 (N_18567,N_15216,N_15351);
or U18568 (N_18568,N_15884,N_15653);
xnor U18569 (N_18569,N_17216,N_17000);
nand U18570 (N_18570,N_17385,N_17003);
and U18571 (N_18571,N_15032,N_15142);
xor U18572 (N_18572,N_15829,N_16468);
xnor U18573 (N_18573,N_16840,N_17312);
and U18574 (N_18574,N_16510,N_16183);
or U18575 (N_18575,N_17022,N_17319);
or U18576 (N_18576,N_16292,N_15226);
xor U18577 (N_18577,N_16893,N_17492);
or U18578 (N_18578,N_16971,N_16543);
xnor U18579 (N_18579,N_17102,N_16056);
nor U18580 (N_18580,N_16026,N_15721);
xor U18581 (N_18581,N_16033,N_15925);
nand U18582 (N_18582,N_17449,N_15904);
nand U18583 (N_18583,N_15090,N_17491);
nand U18584 (N_18584,N_16502,N_16654);
nand U18585 (N_18585,N_17292,N_16725);
nand U18586 (N_18586,N_15998,N_15210);
or U18587 (N_18587,N_16969,N_15841);
xnor U18588 (N_18588,N_16110,N_15838);
xnor U18589 (N_18589,N_16242,N_15602);
xnor U18590 (N_18590,N_16447,N_16738);
xnor U18591 (N_18591,N_16241,N_17362);
and U18592 (N_18592,N_16958,N_16586);
or U18593 (N_18593,N_16733,N_15466);
and U18594 (N_18594,N_15750,N_17389);
xnor U18595 (N_18595,N_16265,N_17214);
or U18596 (N_18596,N_16318,N_16301);
xor U18597 (N_18597,N_15519,N_15197);
or U18598 (N_18598,N_15457,N_15816);
and U18599 (N_18599,N_15643,N_17253);
nand U18600 (N_18600,N_16482,N_16518);
nand U18601 (N_18601,N_16272,N_16819);
xnor U18602 (N_18602,N_16129,N_16271);
and U18603 (N_18603,N_16735,N_16061);
nand U18604 (N_18604,N_15944,N_15027);
xor U18605 (N_18605,N_16984,N_16935);
and U18606 (N_18606,N_15397,N_16837);
nor U18607 (N_18607,N_17230,N_15963);
nor U18608 (N_18608,N_16912,N_17349);
nand U18609 (N_18609,N_17425,N_16779);
nor U18610 (N_18610,N_17187,N_15437);
nand U18611 (N_18611,N_16698,N_16649);
and U18612 (N_18612,N_17267,N_15791);
nor U18613 (N_18613,N_15030,N_15301);
nand U18614 (N_18614,N_16233,N_15267);
and U18615 (N_18615,N_16449,N_15203);
xor U18616 (N_18616,N_16571,N_16150);
nand U18617 (N_18617,N_16337,N_16985);
xor U18618 (N_18618,N_15304,N_15835);
xor U18619 (N_18619,N_17014,N_15125);
xnor U18620 (N_18620,N_16491,N_15478);
nand U18621 (N_18621,N_17333,N_16839);
nand U18622 (N_18622,N_16335,N_15232);
nor U18623 (N_18623,N_16322,N_15291);
xor U18624 (N_18624,N_16578,N_15455);
or U18625 (N_18625,N_16802,N_15053);
nand U18626 (N_18626,N_17436,N_17112);
and U18627 (N_18627,N_17012,N_16336);
or U18628 (N_18628,N_16856,N_16007);
xor U18629 (N_18629,N_17302,N_15362);
and U18630 (N_18630,N_15143,N_15785);
nand U18631 (N_18631,N_15080,N_16275);
nand U18632 (N_18632,N_16556,N_16762);
nand U18633 (N_18633,N_16532,N_15237);
xor U18634 (N_18634,N_16202,N_15960);
or U18635 (N_18635,N_15039,N_15490);
nand U18636 (N_18636,N_16080,N_16987);
nand U18637 (N_18637,N_15163,N_16097);
nor U18638 (N_18638,N_16850,N_16699);
or U18639 (N_18639,N_17122,N_17467);
xor U18640 (N_18640,N_17409,N_15668);
or U18641 (N_18641,N_16167,N_16039);
xor U18642 (N_18642,N_16010,N_15404);
or U18643 (N_18643,N_16350,N_15447);
xnor U18644 (N_18644,N_15104,N_16141);
or U18645 (N_18645,N_15166,N_15042);
and U18646 (N_18646,N_16768,N_16446);
or U18647 (N_18647,N_17179,N_15225);
nor U18648 (N_18648,N_17472,N_17429);
nor U18649 (N_18649,N_17343,N_17286);
xnor U18650 (N_18650,N_16789,N_17258);
nor U18651 (N_18651,N_15180,N_17192);
xnor U18652 (N_18652,N_16707,N_17451);
xnor U18653 (N_18653,N_15309,N_15096);
nor U18654 (N_18654,N_17370,N_16357);
nand U18655 (N_18655,N_15732,N_15966);
nand U18656 (N_18656,N_17093,N_15916);
or U18657 (N_18657,N_17098,N_15211);
or U18658 (N_18658,N_16015,N_15627);
and U18659 (N_18659,N_15697,N_17483);
and U18660 (N_18660,N_17019,N_17246);
nor U18661 (N_18661,N_15606,N_15551);
or U18662 (N_18662,N_17119,N_17132);
nor U18663 (N_18663,N_15308,N_16573);
xnor U18664 (N_18664,N_15861,N_15622);
xnor U18665 (N_18665,N_15262,N_15654);
nor U18666 (N_18666,N_16184,N_17340);
nand U18667 (N_18667,N_15253,N_16885);
and U18668 (N_18668,N_15139,N_16600);
or U18669 (N_18669,N_17368,N_15747);
or U18670 (N_18670,N_17065,N_16426);
xnor U18671 (N_18671,N_16027,N_15793);
or U18672 (N_18672,N_15141,N_16991);
and U18673 (N_18673,N_16351,N_16872);
and U18674 (N_18674,N_16526,N_15270);
xor U18675 (N_18675,N_15601,N_17032);
or U18676 (N_18676,N_16681,N_16355);
and U18677 (N_18677,N_17476,N_15374);
nand U18678 (N_18678,N_15103,N_16626);
xnor U18679 (N_18679,N_17412,N_17484);
nand U18680 (N_18680,N_16264,N_15392);
xnor U18681 (N_18681,N_15338,N_17264);
or U18682 (N_18682,N_16219,N_15017);
and U18683 (N_18683,N_16602,N_17372);
or U18684 (N_18684,N_15803,N_17172);
xnor U18685 (N_18685,N_15161,N_15572);
nor U18686 (N_18686,N_15385,N_15605);
and U18687 (N_18687,N_15790,N_17059);
nor U18688 (N_18688,N_17231,N_17113);
nor U18689 (N_18689,N_17481,N_16146);
nand U18690 (N_18690,N_15293,N_15200);
or U18691 (N_18691,N_16099,N_17471);
xor U18692 (N_18692,N_15209,N_16460);
nor U18693 (N_18693,N_17463,N_17050);
nor U18694 (N_18694,N_17357,N_15616);
nor U18695 (N_18695,N_17454,N_17176);
or U18696 (N_18696,N_16463,N_16500);
or U18697 (N_18697,N_15388,N_16575);
xor U18698 (N_18698,N_15321,N_16688);
xnor U18699 (N_18699,N_16836,N_15151);
xnor U18700 (N_18700,N_15718,N_16466);
or U18701 (N_18701,N_15923,N_17002);
and U18702 (N_18702,N_15222,N_16371);
and U18703 (N_18703,N_17401,N_17023);
xor U18704 (N_18704,N_16434,N_15449);
nand U18705 (N_18705,N_15520,N_15586);
xnor U18706 (N_18706,N_15256,N_16719);
or U18707 (N_18707,N_16484,N_16660);
nand U18708 (N_18708,N_15924,N_16047);
or U18709 (N_18709,N_16507,N_15159);
and U18710 (N_18710,N_16018,N_17263);
nand U18711 (N_18711,N_15479,N_15982);
nand U18712 (N_18712,N_16517,N_17355);
nor U18713 (N_18713,N_16620,N_15871);
or U18714 (N_18714,N_16566,N_16923);
and U18715 (N_18715,N_15369,N_16886);
and U18716 (N_18716,N_17338,N_15854);
or U18717 (N_18717,N_16521,N_15514);
and U18718 (N_18718,N_15626,N_16088);
and U18719 (N_18719,N_16189,N_15085);
nor U18720 (N_18720,N_17178,N_16176);
nor U18721 (N_18721,N_15101,N_15418);
nor U18722 (N_18722,N_16530,N_15789);
xnor U18723 (N_18723,N_16902,N_15774);
and U18724 (N_18724,N_16508,N_16567);
nor U18725 (N_18725,N_16547,N_16561);
or U18726 (N_18726,N_16723,N_17487);
nor U18727 (N_18727,N_16915,N_15806);
nor U18728 (N_18728,N_16279,N_16006);
or U18729 (N_18729,N_15663,N_15660);
or U18730 (N_18730,N_15754,N_15329);
xor U18731 (N_18731,N_15953,N_15062);
nor U18732 (N_18732,N_16103,N_15992);
xnor U18733 (N_18733,N_16989,N_15194);
nand U18734 (N_18734,N_15416,N_15305);
nor U18735 (N_18735,N_15227,N_16744);
xor U18736 (N_18736,N_16084,N_16610);
and U18737 (N_18737,N_17458,N_17083);
nor U18738 (N_18738,N_15157,N_17306);
xor U18739 (N_18739,N_15072,N_16903);
xor U18740 (N_18740,N_17053,N_15120);
nor U18741 (N_18741,N_16617,N_16467);
nand U18742 (N_18742,N_16302,N_15898);
xor U18743 (N_18743,N_15910,N_15866);
nor U18744 (N_18744,N_16430,N_15891);
or U18745 (N_18745,N_15366,N_16763);
nor U18746 (N_18746,N_17189,N_16628);
xor U18747 (N_18747,N_16549,N_15075);
nand U18748 (N_18748,N_15646,N_17236);
nand U18749 (N_18749,N_17077,N_15356);
and U18750 (N_18750,N_15149,N_15740);
and U18751 (N_18751,N_15207,N_15173);
or U18752 (N_18752,N_16071,N_16249);
nor U18753 (N_18753,N_15472,N_16308);
and U18754 (N_18754,N_15633,N_15763);
nor U18755 (N_18755,N_15792,N_15840);
xnor U18756 (N_18756,N_15012,N_16194);
nand U18757 (N_18757,N_15274,N_15452);
nor U18758 (N_18758,N_17082,N_15599);
nor U18759 (N_18759,N_17334,N_17432);
xor U18760 (N_18760,N_17427,N_16121);
nor U18761 (N_18761,N_16243,N_15658);
nand U18762 (N_18762,N_15305,N_15646);
or U18763 (N_18763,N_15748,N_17187);
xor U18764 (N_18764,N_15430,N_17154);
or U18765 (N_18765,N_15563,N_15446);
and U18766 (N_18766,N_15572,N_15895);
nand U18767 (N_18767,N_17088,N_17359);
nor U18768 (N_18768,N_16105,N_17202);
and U18769 (N_18769,N_16428,N_17249);
or U18770 (N_18770,N_17058,N_17072);
nand U18771 (N_18771,N_15382,N_16531);
xnor U18772 (N_18772,N_15287,N_15986);
nor U18773 (N_18773,N_15842,N_16217);
xor U18774 (N_18774,N_15848,N_16021);
and U18775 (N_18775,N_16412,N_17180);
nor U18776 (N_18776,N_16621,N_15673);
or U18777 (N_18777,N_16420,N_17313);
nor U18778 (N_18778,N_16118,N_16272);
or U18779 (N_18779,N_17247,N_17391);
and U18780 (N_18780,N_15265,N_15594);
or U18781 (N_18781,N_16245,N_16722);
xor U18782 (N_18782,N_17474,N_15404);
xor U18783 (N_18783,N_16273,N_15929);
or U18784 (N_18784,N_16961,N_16815);
nor U18785 (N_18785,N_15140,N_15314);
nand U18786 (N_18786,N_16020,N_15936);
or U18787 (N_18787,N_17031,N_16481);
and U18788 (N_18788,N_16163,N_15566);
or U18789 (N_18789,N_17093,N_16041);
and U18790 (N_18790,N_16518,N_17390);
nor U18791 (N_18791,N_15106,N_16088);
xnor U18792 (N_18792,N_16962,N_15693);
nand U18793 (N_18793,N_16401,N_17358);
nor U18794 (N_18794,N_17197,N_16380);
or U18795 (N_18795,N_15193,N_16659);
and U18796 (N_18796,N_15366,N_16568);
nand U18797 (N_18797,N_17384,N_17445);
or U18798 (N_18798,N_15196,N_15342);
nor U18799 (N_18799,N_15819,N_17350);
xnor U18800 (N_18800,N_15348,N_16836);
xnor U18801 (N_18801,N_17150,N_17465);
and U18802 (N_18802,N_17100,N_17431);
nor U18803 (N_18803,N_16848,N_15490);
nand U18804 (N_18804,N_17165,N_16921);
nor U18805 (N_18805,N_15540,N_17261);
or U18806 (N_18806,N_15319,N_17378);
xor U18807 (N_18807,N_15688,N_17454);
xnor U18808 (N_18808,N_16489,N_16230);
xor U18809 (N_18809,N_15284,N_15531);
nor U18810 (N_18810,N_16294,N_16171);
xor U18811 (N_18811,N_15686,N_15464);
nand U18812 (N_18812,N_16945,N_15691);
and U18813 (N_18813,N_15848,N_16838);
nor U18814 (N_18814,N_15134,N_16279);
nand U18815 (N_18815,N_16725,N_16065);
nor U18816 (N_18816,N_17422,N_16159);
nand U18817 (N_18817,N_15953,N_16279);
nand U18818 (N_18818,N_17017,N_15185);
xnor U18819 (N_18819,N_17330,N_16655);
xor U18820 (N_18820,N_16296,N_15027);
and U18821 (N_18821,N_15109,N_17362);
nand U18822 (N_18822,N_16308,N_15855);
and U18823 (N_18823,N_17280,N_15183);
nor U18824 (N_18824,N_17220,N_15720);
nand U18825 (N_18825,N_16037,N_16818);
and U18826 (N_18826,N_15308,N_17032);
and U18827 (N_18827,N_17052,N_15694);
nand U18828 (N_18828,N_16820,N_16858);
or U18829 (N_18829,N_16881,N_16892);
nand U18830 (N_18830,N_16861,N_17098);
xnor U18831 (N_18831,N_15355,N_15769);
xor U18832 (N_18832,N_16597,N_15013);
xor U18833 (N_18833,N_16314,N_17051);
and U18834 (N_18834,N_16585,N_16130);
and U18835 (N_18835,N_15589,N_16508);
xnor U18836 (N_18836,N_15072,N_15019);
and U18837 (N_18837,N_17445,N_15255);
or U18838 (N_18838,N_16646,N_17169);
nor U18839 (N_18839,N_17374,N_17137);
xnor U18840 (N_18840,N_16304,N_17457);
xnor U18841 (N_18841,N_16961,N_16012);
nand U18842 (N_18842,N_16435,N_16481);
nor U18843 (N_18843,N_15254,N_16775);
nand U18844 (N_18844,N_16080,N_16726);
and U18845 (N_18845,N_15703,N_16732);
and U18846 (N_18846,N_15833,N_16676);
nand U18847 (N_18847,N_16352,N_16798);
and U18848 (N_18848,N_15688,N_15067);
xor U18849 (N_18849,N_17206,N_15342);
and U18850 (N_18850,N_17220,N_15477);
xnor U18851 (N_18851,N_15837,N_16538);
or U18852 (N_18852,N_16214,N_16953);
nor U18853 (N_18853,N_16082,N_15094);
nor U18854 (N_18854,N_15330,N_16563);
nor U18855 (N_18855,N_15175,N_16261);
and U18856 (N_18856,N_15972,N_15427);
nand U18857 (N_18857,N_16922,N_15686);
or U18858 (N_18858,N_16270,N_16145);
xor U18859 (N_18859,N_15964,N_16454);
and U18860 (N_18860,N_17417,N_17287);
xor U18861 (N_18861,N_15743,N_15424);
nand U18862 (N_18862,N_15187,N_16296);
and U18863 (N_18863,N_16209,N_15990);
nor U18864 (N_18864,N_16828,N_16763);
nand U18865 (N_18865,N_17194,N_15525);
nand U18866 (N_18866,N_16344,N_15423);
and U18867 (N_18867,N_16165,N_17042);
or U18868 (N_18868,N_15788,N_16718);
xor U18869 (N_18869,N_15607,N_16961);
and U18870 (N_18870,N_17339,N_16183);
nor U18871 (N_18871,N_16568,N_15254);
nand U18872 (N_18872,N_16705,N_15062);
nor U18873 (N_18873,N_15338,N_16647);
or U18874 (N_18874,N_16853,N_16829);
and U18875 (N_18875,N_16579,N_15520);
or U18876 (N_18876,N_16012,N_15664);
nor U18877 (N_18877,N_16925,N_15688);
and U18878 (N_18878,N_16789,N_15774);
xnor U18879 (N_18879,N_15695,N_17457);
or U18880 (N_18880,N_17115,N_17370);
or U18881 (N_18881,N_17487,N_16516);
nand U18882 (N_18882,N_17169,N_15749);
nand U18883 (N_18883,N_17184,N_17417);
and U18884 (N_18884,N_16182,N_16567);
xnor U18885 (N_18885,N_15338,N_15930);
or U18886 (N_18886,N_16834,N_15000);
or U18887 (N_18887,N_17073,N_16320);
nor U18888 (N_18888,N_16118,N_16348);
or U18889 (N_18889,N_16016,N_15888);
xor U18890 (N_18890,N_16889,N_15154);
xnor U18891 (N_18891,N_16597,N_15801);
or U18892 (N_18892,N_16511,N_15909);
or U18893 (N_18893,N_16406,N_17040);
nand U18894 (N_18894,N_15376,N_17207);
and U18895 (N_18895,N_15546,N_15529);
or U18896 (N_18896,N_16594,N_17080);
or U18897 (N_18897,N_17260,N_16239);
nor U18898 (N_18898,N_16879,N_16158);
nor U18899 (N_18899,N_16186,N_16684);
nor U18900 (N_18900,N_17482,N_15530);
or U18901 (N_18901,N_16395,N_16814);
nor U18902 (N_18902,N_17094,N_17252);
nand U18903 (N_18903,N_16533,N_16270);
nand U18904 (N_18904,N_15185,N_16578);
nand U18905 (N_18905,N_16781,N_15764);
or U18906 (N_18906,N_16634,N_16563);
and U18907 (N_18907,N_16124,N_16904);
xnor U18908 (N_18908,N_17231,N_16696);
xor U18909 (N_18909,N_16138,N_16599);
and U18910 (N_18910,N_15074,N_17130);
xnor U18911 (N_18911,N_15536,N_15666);
nand U18912 (N_18912,N_15435,N_15128);
nor U18913 (N_18913,N_15618,N_15460);
nand U18914 (N_18914,N_16290,N_16553);
and U18915 (N_18915,N_17129,N_16152);
xor U18916 (N_18916,N_15871,N_16875);
nand U18917 (N_18917,N_15434,N_16863);
and U18918 (N_18918,N_17160,N_17163);
or U18919 (N_18919,N_15770,N_16992);
nor U18920 (N_18920,N_17356,N_15742);
xor U18921 (N_18921,N_16958,N_15108);
or U18922 (N_18922,N_15826,N_15500);
nand U18923 (N_18923,N_15798,N_15060);
nand U18924 (N_18924,N_16118,N_15282);
and U18925 (N_18925,N_15564,N_15345);
nand U18926 (N_18926,N_16581,N_15482);
or U18927 (N_18927,N_16055,N_15256);
nor U18928 (N_18928,N_17423,N_15816);
nor U18929 (N_18929,N_17277,N_15042);
nand U18930 (N_18930,N_16451,N_15174);
nor U18931 (N_18931,N_16122,N_16506);
nor U18932 (N_18932,N_17175,N_15644);
nand U18933 (N_18933,N_16323,N_15173);
nand U18934 (N_18934,N_16172,N_15459);
nand U18935 (N_18935,N_16244,N_17222);
nand U18936 (N_18936,N_15097,N_17055);
nand U18937 (N_18937,N_15820,N_15007);
or U18938 (N_18938,N_17139,N_16916);
nand U18939 (N_18939,N_15102,N_16576);
xor U18940 (N_18940,N_16594,N_15825);
or U18941 (N_18941,N_15067,N_16372);
and U18942 (N_18942,N_17140,N_17174);
xnor U18943 (N_18943,N_16640,N_16495);
nor U18944 (N_18944,N_16417,N_17170);
xor U18945 (N_18945,N_15614,N_16348);
nand U18946 (N_18946,N_15857,N_16567);
nand U18947 (N_18947,N_16718,N_16761);
or U18948 (N_18948,N_16793,N_17359);
xnor U18949 (N_18949,N_15206,N_17346);
and U18950 (N_18950,N_15556,N_16698);
xor U18951 (N_18951,N_17097,N_15407);
nand U18952 (N_18952,N_15565,N_17182);
and U18953 (N_18953,N_16660,N_16840);
nor U18954 (N_18954,N_15011,N_16826);
nor U18955 (N_18955,N_17234,N_15196);
nor U18956 (N_18956,N_16905,N_15744);
and U18957 (N_18957,N_16965,N_17064);
and U18958 (N_18958,N_15211,N_17371);
or U18959 (N_18959,N_15599,N_15892);
nor U18960 (N_18960,N_16332,N_15374);
and U18961 (N_18961,N_16986,N_16467);
and U18962 (N_18962,N_17478,N_16875);
nor U18963 (N_18963,N_15162,N_17193);
nand U18964 (N_18964,N_15053,N_16118);
or U18965 (N_18965,N_17354,N_15692);
and U18966 (N_18966,N_16200,N_15169);
nor U18967 (N_18967,N_15520,N_15443);
or U18968 (N_18968,N_16026,N_15870);
nand U18969 (N_18969,N_16081,N_15152);
nand U18970 (N_18970,N_16431,N_16261);
and U18971 (N_18971,N_17354,N_15750);
or U18972 (N_18972,N_15496,N_15256);
nor U18973 (N_18973,N_16756,N_16666);
nand U18974 (N_18974,N_15594,N_16591);
or U18975 (N_18975,N_17434,N_15669);
nand U18976 (N_18976,N_17358,N_16779);
xor U18977 (N_18977,N_16608,N_16973);
and U18978 (N_18978,N_15044,N_15622);
xor U18979 (N_18979,N_16893,N_15123);
xor U18980 (N_18980,N_15111,N_16313);
nand U18981 (N_18981,N_15702,N_17002);
nor U18982 (N_18982,N_15234,N_17044);
nor U18983 (N_18983,N_15183,N_15411);
nor U18984 (N_18984,N_16567,N_15026);
xor U18985 (N_18985,N_15946,N_16555);
and U18986 (N_18986,N_17216,N_16425);
or U18987 (N_18987,N_15592,N_16236);
nand U18988 (N_18988,N_15647,N_16903);
nor U18989 (N_18989,N_16828,N_15438);
or U18990 (N_18990,N_16257,N_16997);
xor U18991 (N_18991,N_16173,N_16825);
nor U18992 (N_18992,N_16387,N_15372);
and U18993 (N_18993,N_16540,N_16606);
nor U18994 (N_18994,N_17342,N_16569);
xnor U18995 (N_18995,N_16841,N_17200);
xor U18996 (N_18996,N_15040,N_15498);
nor U18997 (N_18997,N_16885,N_15874);
nand U18998 (N_18998,N_16022,N_15303);
nand U18999 (N_18999,N_15153,N_15911);
xor U19000 (N_19000,N_15388,N_17481);
and U19001 (N_19001,N_15431,N_15772);
nand U19002 (N_19002,N_16070,N_16081);
and U19003 (N_19003,N_17330,N_15349);
and U19004 (N_19004,N_16029,N_17204);
or U19005 (N_19005,N_15107,N_17372);
or U19006 (N_19006,N_15422,N_16980);
or U19007 (N_19007,N_17139,N_16377);
nand U19008 (N_19008,N_16126,N_16756);
xor U19009 (N_19009,N_15996,N_15008);
nand U19010 (N_19010,N_16750,N_15695);
nor U19011 (N_19011,N_15601,N_16466);
nor U19012 (N_19012,N_16268,N_17201);
and U19013 (N_19013,N_16408,N_15320);
nand U19014 (N_19014,N_15246,N_16913);
xor U19015 (N_19015,N_17267,N_15074);
xnor U19016 (N_19016,N_17053,N_16242);
xor U19017 (N_19017,N_16895,N_15602);
and U19018 (N_19018,N_16116,N_17065);
nor U19019 (N_19019,N_16222,N_16469);
or U19020 (N_19020,N_17111,N_16487);
nand U19021 (N_19021,N_17326,N_16542);
or U19022 (N_19022,N_15514,N_16578);
xnor U19023 (N_19023,N_16086,N_16273);
nand U19024 (N_19024,N_16028,N_16186);
xnor U19025 (N_19025,N_15246,N_17130);
nand U19026 (N_19026,N_16535,N_17211);
xnor U19027 (N_19027,N_16643,N_15684);
and U19028 (N_19028,N_17391,N_17300);
nand U19029 (N_19029,N_16202,N_15074);
or U19030 (N_19030,N_17441,N_17241);
nor U19031 (N_19031,N_16231,N_15801);
xnor U19032 (N_19032,N_17193,N_16100);
and U19033 (N_19033,N_15142,N_15507);
and U19034 (N_19034,N_16118,N_16722);
nor U19035 (N_19035,N_17101,N_17134);
xnor U19036 (N_19036,N_16882,N_15819);
nor U19037 (N_19037,N_15750,N_16572);
or U19038 (N_19038,N_15564,N_16704);
nor U19039 (N_19039,N_16005,N_16543);
and U19040 (N_19040,N_16115,N_15715);
nor U19041 (N_19041,N_16205,N_17188);
nand U19042 (N_19042,N_17244,N_16420);
nand U19043 (N_19043,N_17171,N_15826);
nand U19044 (N_19044,N_15868,N_15321);
and U19045 (N_19045,N_17030,N_16198);
xor U19046 (N_19046,N_16236,N_17494);
nand U19047 (N_19047,N_16728,N_15988);
or U19048 (N_19048,N_17477,N_15913);
and U19049 (N_19049,N_15823,N_16542);
or U19050 (N_19050,N_15784,N_17215);
and U19051 (N_19051,N_15434,N_16795);
nand U19052 (N_19052,N_16381,N_16006);
xor U19053 (N_19053,N_15450,N_16328);
xnor U19054 (N_19054,N_16666,N_15783);
or U19055 (N_19055,N_17135,N_17219);
and U19056 (N_19056,N_16772,N_16911);
or U19057 (N_19057,N_15789,N_16041);
or U19058 (N_19058,N_16281,N_16638);
xor U19059 (N_19059,N_15332,N_15778);
nor U19060 (N_19060,N_15083,N_17309);
xor U19061 (N_19061,N_15174,N_15873);
nor U19062 (N_19062,N_15193,N_16595);
and U19063 (N_19063,N_15729,N_15093);
and U19064 (N_19064,N_15115,N_16742);
xnor U19065 (N_19065,N_16853,N_15954);
nand U19066 (N_19066,N_16029,N_17271);
or U19067 (N_19067,N_17242,N_15943);
and U19068 (N_19068,N_16082,N_16200);
nor U19069 (N_19069,N_15862,N_17464);
xor U19070 (N_19070,N_16135,N_15392);
and U19071 (N_19071,N_16090,N_17288);
xor U19072 (N_19072,N_15750,N_17009);
or U19073 (N_19073,N_15874,N_17061);
and U19074 (N_19074,N_17446,N_17036);
or U19075 (N_19075,N_16497,N_15516);
or U19076 (N_19076,N_17011,N_15016);
nor U19077 (N_19077,N_15445,N_17430);
xor U19078 (N_19078,N_15457,N_16749);
and U19079 (N_19079,N_16775,N_15099);
nand U19080 (N_19080,N_15977,N_16100);
and U19081 (N_19081,N_16356,N_16237);
nor U19082 (N_19082,N_15499,N_16751);
nor U19083 (N_19083,N_15339,N_17133);
or U19084 (N_19084,N_17320,N_15810);
nand U19085 (N_19085,N_16190,N_16823);
xor U19086 (N_19086,N_16472,N_17333);
xor U19087 (N_19087,N_17079,N_15956);
nor U19088 (N_19088,N_16525,N_16161);
nand U19089 (N_19089,N_16573,N_16943);
nand U19090 (N_19090,N_15362,N_15454);
nand U19091 (N_19091,N_15099,N_15491);
or U19092 (N_19092,N_15059,N_17316);
or U19093 (N_19093,N_16998,N_15585);
nand U19094 (N_19094,N_15781,N_17042);
nor U19095 (N_19095,N_15720,N_15139);
nor U19096 (N_19096,N_16846,N_15748);
or U19097 (N_19097,N_15340,N_16217);
xnor U19098 (N_19098,N_16696,N_16634);
or U19099 (N_19099,N_16238,N_16557);
or U19100 (N_19100,N_15444,N_15238);
or U19101 (N_19101,N_17497,N_15957);
nor U19102 (N_19102,N_16994,N_17366);
or U19103 (N_19103,N_15852,N_15325);
nor U19104 (N_19104,N_16851,N_15633);
nand U19105 (N_19105,N_17482,N_16292);
xnor U19106 (N_19106,N_15427,N_16507);
and U19107 (N_19107,N_15031,N_17303);
or U19108 (N_19108,N_15715,N_16103);
nor U19109 (N_19109,N_16474,N_17026);
nor U19110 (N_19110,N_15272,N_16837);
nor U19111 (N_19111,N_16312,N_17112);
and U19112 (N_19112,N_15750,N_16652);
nor U19113 (N_19113,N_16816,N_17363);
nand U19114 (N_19114,N_16945,N_15921);
nand U19115 (N_19115,N_16325,N_17094);
nor U19116 (N_19116,N_16670,N_15233);
and U19117 (N_19117,N_15405,N_16477);
nor U19118 (N_19118,N_15253,N_16323);
nor U19119 (N_19119,N_16576,N_16739);
nand U19120 (N_19120,N_16292,N_17075);
or U19121 (N_19121,N_17074,N_16711);
xor U19122 (N_19122,N_15497,N_16680);
xor U19123 (N_19123,N_17081,N_17138);
nand U19124 (N_19124,N_17443,N_15937);
nand U19125 (N_19125,N_16986,N_16834);
and U19126 (N_19126,N_15175,N_16045);
xor U19127 (N_19127,N_15638,N_15924);
or U19128 (N_19128,N_15462,N_16481);
xnor U19129 (N_19129,N_15592,N_15314);
nor U19130 (N_19130,N_16395,N_15060);
nor U19131 (N_19131,N_16367,N_15706);
xor U19132 (N_19132,N_15115,N_16539);
and U19133 (N_19133,N_17443,N_15045);
xor U19134 (N_19134,N_16243,N_16091);
nor U19135 (N_19135,N_15370,N_15158);
xor U19136 (N_19136,N_15260,N_15457);
or U19137 (N_19137,N_15814,N_16711);
nor U19138 (N_19138,N_15524,N_16173);
and U19139 (N_19139,N_17093,N_15980);
and U19140 (N_19140,N_17169,N_17161);
nand U19141 (N_19141,N_17427,N_15078);
and U19142 (N_19142,N_16586,N_15312);
xnor U19143 (N_19143,N_16929,N_15883);
xor U19144 (N_19144,N_15836,N_16553);
xor U19145 (N_19145,N_16607,N_16520);
nand U19146 (N_19146,N_15571,N_15499);
nand U19147 (N_19147,N_16447,N_15728);
xnor U19148 (N_19148,N_15319,N_16042);
and U19149 (N_19149,N_17345,N_16920);
or U19150 (N_19150,N_16876,N_15978);
xnor U19151 (N_19151,N_16606,N_16525);
nand U19152 (N_19152,N_17072,N_15731);
nor U19153 (N_19153,N_16748,N_15143);
and U19154 (N_19154,N_16744,N_15152);
xnor U19155 (N_19155,N_16277,N_16394);
nor U19156 (N_19156,N_15369,N_16417);
or U19157 (N_19157,N_16138,N_15388);
xnor U19158 (N_19158,N_16391,N_16583);
or U19159 (N_19159,N_15687,N_16002);
nand U19160 (N_19160,N_17207,N_16866);
nand U19161 (N_19161,N_16381,N_15068);
and U19162 (N_19162,N_16392,N_16115);
nand U19163 (N_19163,N_15990,N_15707);
and U19164 (N_19164,N_15176,N_16873);
or U19165 (N_19165,N_17101,N_15729);
xor U19166 (N_19166,N_16576,N_16657);
nor U19167 (N_19167,N_16762,N_17152);
or U19168 (N_19168,N_17428,N_16183);
or U19169 (N_19169,N_15761,N_17379);
nor U19170 (N_19170,N_17086,N_15992);
nor U19171 (N_19171,N_15511,N_17347);
nand U19172 (N_19172,N_17353,N_16628);
nand U19173 (N_19173,N_17142,N_16543);
xor U19174 (N_19174,N_17140,N_15065);
and U19175 (N_19175,N_15485,N_15934);
nor U19176 (N_19176,N_15529,N_15878);
nand U19177 (N_19177,N_17148,N_15409);
xor U19178 (N_19178,N_16109,N_16430);
or U19179 (N_19179,N_17270,N_16555);
xor U19180 (N_19180,N_15186,N_16848);
nor U19181 (N_19181,N_17195,N_17312);
nand U19182 (N_19182,N_16616,N_16213);
xor U19183 (N_19183,N_16677,N_17422);
and U19184 (N_19184,N_15521,N_16171);
xnor U19185 (N_19185,N_16762,N_15844);
xor U19186 (N_19186,N_16260,N_16001);
nor U19187 (N_19187,N_15457,N_17157);
xnor U19188 (N_19188,N_15291,N_16247);
or U19189 (N_19189,N_16278,N_17490);
xor U19190 (N_19190,N_15213,N_16016);
and U19191 (N_19191,N_15557,N_16452);
or U19192 (N_19192,N_15710,N_15368);
or U19193 (N_19193,N_16805,N_17263);
or U19194 (N_19194,N_15195,N_15450);
and U19195 (N_19195,N_15167,N_16760);
or U19196 (N_19196,N_15778,N_15167);
and U19197 (N_19197,N_15508,N_16299);
nor U19198 (N_19198,N_15635,N_16568);
nand U19199 (N_19199,N_16948,N_17267);
or U19200 (N_19200,N_16249,N_15995);
xor U19201 (N_19201,N_16679,N_16186);
xor U19202 (N_19202,N_16200,N_15353);
or U19203 (N_19203,N_16633,N_15667);
or U19204 (N_19204,N_15246,N_16329);
xor U19205 (N_19205,N_17333,N_17125);
and U19206 (N_19206,N_15631,N_15885);
or U19207 (N_19207,N_17248,N_17143);
and U19208 (N_19208,N_16989,N_17220);
nor U19209 (N_19209,N_16614,N_15494);
xnor U19210 (N_19210,N_15347,N_15177);
and U19211 (N_19211,N_17266,N_15263);
xor U19212 (N_19212,N_17302,N_17022);
xnor U19213 (N_19213,N_17399,N_15392);
or U19214 (N_19214,N_16455,N_16258);
xnor U19215 (N_19215,N_15019,N_15412);
xnor U19216 (N_19216,N_15465,N_16462);
or U19217 (N_19217,N_17459,N_16529);
or U19218 (N_19218,N_17421,N_15482);
nor U19219 (N_19219,N_15656,N_15519);
nand U19220 (N_19220,N_15820,N_16313);
nand U19221 (N_19221,N_16965,N_16917);
or U19222 (N_19222,N_15119,N_16398);
or U19223 (N_19223,N_15884,N_15384);
nor U19224 (N_19224,N_16485,N_16174);
xor U19225 (N_19225,N_15134,N_15894);
or U19226 (N_19226,N_16882,N_17488);
or U19227 (N_19227,N_16428,N_15414);
nor U19228 (N_19228,N_15026,N_15580);
or U19229 (N_19229,N_17057,N_15120);
or U19230 (N_19230,N_17315,N_15390);
nand U19231 (N_19231,N_16832,N_16127);
or U19232 (N_19232,N_15532,N_17017);
and U19233 (N_19233,N_16060,N_15471);
or U19234 (N_19234,N_15277,N_15456);
xor U19235 (N_19235,N_15211,N_16898);
and U19236 (N_19236,N_15376,N_15703);
xor U19237 (N_19237,N_17279,N_17459);
nand U19238 (N_19238,N_16062,N_15440);
xnor U19239 (N_19239,N_15494,N_16720);
xnor U19240 (N_19240,N_15338,N_16043);
nand U19241 (N_19241,N_15272,N_16232);
and U19242 (N_19242,N_16350,N_17127);
nor U19243 (N_19243,N_16357,N_15851);
or U19244 (N_19244,N_15477,N_15382);
or U19245 (N_19245,N_16001,N_15322);
and U19246 (N_19246,N_16445,N_15808);
nand U19247 (N_19247,N_15937,N_15684);
or U19248 (N_19248,N_16896,N_16907);
or U19249 (N_19249,N_16550,N_16463);
xnor U19250 (N_19250,N_17323,N_16767);
and U19251 (N_19251,N_15409,N_15280);
or U19252 (N_19252,N_17310,N_16837);
and U19253 (N_19253,N_15754,N_17282);
or U19254 (N_19254,N_17033,N_15755);
and U19255 (N_19255,N_16764,N_16941);
xor U19256 (N_19256,N_17436,N_15727);
xnor U19257 (N_19257,N_15905,N_15926);
nor U19258 (N_19258,N_16016,N_15682);
xor U19259 (N_19259,N_15487,N_15765);
xnor U19260 (N_19260,N_15163,N_16486);
and U19261 (N_19261,N_15231,N_17142);
or U19262 (N_19262,N_16240,N_17387);
or U19263 (N_19263,N_17425,N_15375);
and U19264 (N_19264,N_16294,N_15354);
or U19265 (N_19265,N_17382,N_16065);
nand U19266 (N_19266,N_17112,N_15109);
and U19267 (N_19267,N_17085,N_15084);
and U19268 (N_19268,N_15797,N_15687);
nand U19269 (N_19269,N_16501,N_17404);
xnor U19270 (N_19270,N_16418,N_16948);
nor U19271 (N_19271,N_16153,N_17066);
xor U19272 (N_19272,N_15706,N_16768);
xor U19273 (N_19273,N_16749,N_15143);
and U19274 (N_19274,N_16125,N_15947);
nand U19275 (N_19275,N_16270,N_16351);
xnor U19276 (N_19276,N_16970,N_15948);
and U19277 (N_19277,N_17190,N_15050);
or U19278 (N_19278,N_17152,N_15643);
and U19279 (N_19279,N_17090,N_15651);
and U19280 (N_19280,N_15919,N_16540);
nand U19281 (N_19281,N_17321,N_15834);
nand U19282 (N_19282,N_15887,N_15797);
nor U19283 (N_19283,N_16800,N_16879);
xnor U19284 (N_19284,N_15835,N_17129);
nor U19285 (N_19285,N_15236,N_15543);
or U19286 (N_19286,N_15612,N_15532);
xnor U19287 (N_19287,N_17082,N_16773);
xnor U19288 (N_19288,N_15903,N_16769);
nand U19289 (N_19289,N_17032,N_16353);
xnor U19290 (N_19290,N_17370,N_15683);
nand U19291 (N_19291,N_15051,N_15518);
xnor U19292 (N_19292,N_15887,N_17100);
or U19293 (N_19293,N_16567,N_17290);
and U19294 (N_19294,N_15086,N_17058);
or U19295 (N_19295,N_15728,N_15836);
nor U19296 (N_19296,N_15458,N_15200);
or U19297 (N_19297,N_15257,N_15332);
xor U19298 (N_19298,N_16054,N_15296);
nand U19299 (N_19299,N_15923,N_17181);
xnor U19300 (N_19300,N_16513,N_17473);
or U19301 (N_19301,N_16590,N_16240);
xor U19302 (N_19302,N_16253,N_16873);
or U19303 (N_19303,N_16550,N_16242);
or U19304 (N_19304,N_15803,N_17204);
or U19305 (N_19305,N_16721,N_16451);
and U19306 (N_19306,N_15492,N_16501);
nor U19307 (N_19307,N_16192,N_17248);
nand U19308 (N_19308,N_17264,N_16331);
nor U19309 (N_19309,N_17459,N_16646);
xor U19310 (N_19310,N_15888,N_16398);
nand U19311 (N_19311,N_16871,N_16609);
xor U19312 (N_19312,N_15227,N_15598);
nand U19313 (N_19313,N_16009,N_16367);
xor U19314 (N_19314,N_15418,N_17448);
xnor U19315 (N_19315,N_17257,N_15069);
nor U19316 (N_19316,N_16963,N_16835);
xor U19317 (N_19317,N_15428,N_15736);
or U19318 (N_19318,N_16262,N_15734);
or U19319 (N_19319,N_16061,N_17019);
nor U19320 (N_19320,N_16980,N_16429);
xor U19321 (N_19321,N_15160,N_15259);
or U19322 (N_19322,N_17362,N_16903);
and U19323 (N_19323,N_16297,N_15442);
or U19324 (N_19324,N_15642,N_15930);
and U19325 (N_19325,N_15722,N_15870);
xnor U19326 (N_19326,N_15043,N_15168);
or U19327 (N_19327,N_15209,N_15375);
xor U19328 (N_19328,N_16307,N_16722);
and U19329 (N_19329,N_17416,N_15923);
nand U19330 (N_19330,N_16088,N_16241);
nand U19331 (N_19331,N_16617,N_15045);
and U19332 (N_19332,N_15363,N_16406);
xnor U19333 (N_19333,N_17275,N_16742);
and U19334 (N_19334,N_16776,N_16830);
nor U19335 (N_19335,N_16095,N_16212);
and U19336 (N_19336,N_16205,N_17158);
nand U19337 (N_19337,N_16366,N_16670);
xor U19338 (N_19338,N_16209,N_16311);
and U19339 (N_19339,N_15037,N_16969);
nor U19340 (N_19340,N_16650,N_15506);
nand U19341 (N_19341,N_15735,N_16272);
nand U19342 (N_19342,N_16973,N_15144);
nand U19343 (N_19343,N_16348,N_15420);
nand U19344 (N_19344,N_16383,N_16116);
and U19345 (N_19345,N_16065,N_15683);
nand U19346 (N_19346,N_17023,N_16827);
or U19347 (N_19347,N_15304,N_15289);
nand U19348 (N_19348,N_15825,N_15323);
nand U19349 (N_19349,N_17447,N_16000);
nand U19350 (N_19350,N_16700,N_15482);
and U19351 (N_19351,N_16176,N_15961);
and U19352 (N_19352,N_17341,N_16244);
or U19353 (N_19353,N_16596,N_15047);
or U19354 (N_19354,N_15493,N_16988);
and U19355 (N_19355,N_16505,N_16428);
nand U19356 (N_19356,N_16152,N_16275);
xor U19357 (N_19357,N_16301,N_15564);
xor U19358 (N_19358,N_15750,N_17155);
or U19359 (N_19359,N_15407,N_16389);
nor U19360 (N_19360,N_16831,N_15331);
nand U19361 (N_19361,N_15593,N_17364);
nor U19362 (N_19362,N_17202,N_15410);
or U19363 (N_19363,N_16529,N_16269);
and U19364 (N_19364,N_15458,N_16701);
and U19365 (N_19365,N_15802,N_15765);
and U19366 (N_19366,N_16415,N_15631);
xnor U19367 (N_19367,N_17185,N_15008);
nor U19368 (N_19368,N_17211,N_17480);
and U19369 (N_19369,N_15274,N_17043);
xor U19370 (N_19370,N_16695,N_16499);
nor U19371 (N_19371,N_15277,N_17303);
or U19372 (N_19372,N_16402,N_16725);
and U19373 (N_19373,N_15024,N_17272);
xnor U19374 (N_19374,N_17266,N_17412);
nor U19375 (N_19375,N_17316,N_17148);
xor U19376 (N_19376,N_15830,N_15844);
nor U19377 (N_19377,N_16081,N_15420);
and U19378 (N_19378,N_15025,N_15520);
nand U19379 (N_19379,N_17083,N_17274);
and U19380 (N_19380,N_17492,N_17418);
nor U19381 (N_19381,N_15135,N_15573);
xnor U19382 (N_19382,N_15671,N_15079);
xor U19383 (N_19383,N_16014,N_16059);
nor U19384 (N_19384,N_16086,N_15839);
or U19385 (N_19385,N_16187,N_17445);
or U19386 (N_19386,N_16895,N_16183);
nor U19387 (N_19387,N_15904,N_15797);
and U19388 (N_19388,N_15861,N_16043);
xor U19389 (N_19389,N_16947,N_15750);
nor U19390 (N_19390,N_15232,N_15920);
nor U19391 (N_19391,N_15818,N_17036);
nor U19392 (N_19392,N_16855,N_15260);
nand U19393 (N_19393,N_16117,N_17362);
or U19394 (N_19394,N_17250,N_16521);
nand U19395 (N_19395,N_15240,N_15632);
nand U19396 (N_19396,N_17440,N_15532);
or U19397 (N_19397,N_17485,N_16497);
nor U19398 (N_19398,N_15516,N_15694);
or U19399 (N_19399,N_16279,N_17003);
and U19400 (N_19400,N_16062,N_15285);
nand U19401 (N_19401,N_15630,N_15757);
nand U19402 (N_19402,N_16758,N_16477);
nand U19403 (N_19403,N_15071,N_17308);
and U19404 (N_19404,N_15787,N_17205);
xor U19405 (N_19405,N_15885,N_16432);
or U19406 (N_19406,N_15138,N_16922);
nand U19407 (N_19407,N_15296,N_16122);
nor U19408 (N_19408,N_17167,N_16969);
and U19409 (N_19409,N_16321,N_16696);
nor U19410 (N_19410,N_16183,N_15194);
nand U19411 (N_19411,N_15113,N_17096);
nor U19412 (N_19412,N_16314,N_16596);
and U19413 (N_19413,N_16460,N_16477);
xor U19414 (N_19414,N_16307,N_15692);
nor U19415 (N_19415,N_15390,N_15289);
or U19416 (N_19416,N_16165,N_15241);
nor U19417 (N_19417,N_15713,N_15588);
nor U19418 (N_19418,N_15112,N_16430);
and U19419 (N_19419,N_15279,N_15498);
or U19420 (N_19420,N_17206,N_17156);
or U19421 (N_19421,N_15778,N_16575);
nand U19422 (N_19422,N_16882,N_16381);
or U19423 (N_19423,N_17456,N_16408);
and U19424 (N_19424,N_16392,N_16043);
nor U19425 (N_19425,N_15420,N_15644);
and U19426 (N_19426,N_17467,N_16680);
nor U19427 (N_19427,N_15039,N_15550);
or U19428 (N_19428,N_16326,N_16076);
or U19429 (N_19429,N_15323,N_16446);
and U19430 (N_19430,N_17047,N_16398);
and U19431 (N_19431,N_16671,N_16285);
nand U19432 (N_19432,N_17468,N_15109);
or U19433 (N_19433,N_16762,N_15247);
nor U19434 (N_19434,N_15422,N_16246);
and U19435 (N_19435,N_16963,N_16011);
or U19436 (N_19436,N_16069,N_16919);
nand U19437 (N_19437,N_16815,N_16925);
and U19438 (N_19438,N_16616,N_15546);
and U19439 (N_19439,N_15056,N_17358);
xnor U19440 (N_19440,N_15339,N_16729);
nand U19441 (N_19441,N_15657,N_16382);
nor U19442 (N_19442,N_15188,N_16897);
nor U19443 (N_19443,N_17128,N_15591);
or U19444 (N_19444,N_16729,N_15693);
nand U19445 (N_19445,N_15184,N_15244);
and U19446 (N_19446,N_15620,N_15328);
xnor U19447 (N_19447,N_15838,N_16105);
nand U19448 (N_19448,N_15537,N_16229);
nand U19449 (N_19449,N_16234,N_15370);
or U19450 (N_19450,N_15465,N_15699);
xnor U19451 (N_19451,N_16457,N_15631);
and U19452 (N_19452,N_15892,N_15977);
xnor U19453 (N_19453,N_15295,N_16645);
nand U19454 (N_19454,N_15213,N_16518);
or U19455 (N_19455,N_15481,N_17376);
nor U19456 (N_19456,N_16008,N_16559);
nor U19457 (N_19457,N_15999,N_15455);
nor U19458 (N_19458,N_15538,N_15851);
or U19459 (N_19459,N_15402,N_15930);
or U19460 (N_19460,N_15288,N_17044);
and U19461 (N_19461,N_15147,N_16330);
or U19462 (N_19462,N_17116,N_16631);
nor U19463 (N_19463,N_17011,N_16112);
xor U19464 (N_19464,N_15483,N_16658);
or U19465 (N_19465,N_15360,N_16853);
and U19466 (N_19466,N_17216,N_16051);
and U19467 (N_19467,N_15078,N_16165);
nand U19468 (N_19468,N_15843,N_16374);
or U19469 (N_19469,N_15797,N_15161);
nor U19470 (N_19470,N_17318,N_16654);
and U19471 (N_19471,N_17064,N_16202);
nand U19472 (N_19472,N_16192,N_16984);
nor U19473 (N_19473,N_16148,N_16760);
and U19474 (N_19474,N_17257,N_17342);
or U19475 (N_19475,N_16253,N_16368);
and U19476 (N_19476,N_15134,N_15219);
xor U19477 (N_19477,N_15812,N_16932);
xnor U19478 (N_19478,N_16672,N_16960);
and U19479 (N_19479,N_15742,N_16938);
or U19480 (N_19480,N_17264,N_16132);
xor U19481 (N_19481,N_15371,N_15728);
nor U19482 (N_19482,N_15542,N_16879);
nand U19483 (N_19483,N_16888,N_15597);
nor U19484 (N_19484,N_16796,N_15185);
or U19485 (N_19485,N_16735,N_16317);
and U19486 (N_19486,N_15852,N_17022);
nor U19487 (N_19487,N_16877,N_15738);
xor U19488 (N_19488,N_15119,N_16888);
or U19489 (N_19489,N_15801,N_16585);
and U19490 (N_19490,N_16574,N_15926);
and U19491 (N_19491,N_15180,N_17233);
or U19492 (N_19492,N_16132,N_16996);
xor U19493 (N_19493,N_15988,N_16318);
nor U19494 (N_19494,N_16318,N_17101);
xnor U19495 (N_19495,N_16620,N_16931);
nor U19496 (N_19496,N_16713,N_16822);
and U19497 (N_19497,N_16861,N_16839);
xor U19498 (N_19498,N_16813,N_16728);
nand U19499 (N_19499,N_15268,N_16801);
nand U19500 (N_19500,N_15456,N_17205);
nand U19501 (N_19501,N_15843,N_16656);
or U19502 (N_19502,N_16291,N_15893);
nor U19503 (N_19503,N_16380,N_16009);
nand U19504 (N_19504,N_17495,N_17326);
or U19505 (N_19505,N_15743,N_15088);
and U19506 (N_19506,N_16153,N_15031);
nand U19507 (N_19507,N_16298,N_16614);
nor U19508 (N_19508,N_17124,N_16117);
or U19509 (N_19509,N_16487,N_15917);
nand U19510 (N_19510,N_16995,N_16689);
nor U19511 (N_19511,N_16907,N_16302);
xor U19512 (N_19512,N_15120,N_15685);
nor U19513 (N_19513,N_17372,N_16250);
and U19514 (N_19514,N_15978,N_17258);
nand U19515 (N_19515,N_16274,N_16337);
nor U19516 (N_19516,N_17214,N_17139);
and U19517 (N_19517,N_15856,N_16538);
and U19518 (N_19518,N_16112,N_16740);
xor U19519 (N_19519,N_15394,N_15581);
or U19520 (N_19520,N_16063,N_15053);
nand U19521 (N_19521,N_17357,N_17182);
nand U19522 (N_19522,N_15349,N_15645);
or U19523 (N_19523,N_15847,N_17171);
xor U19524 (N_19524,N_16810,N_16207);
or U19525 (N_19525,N_16437,N_16255);
nand U19526 (N_19526,N_15021,N_15236);
nor U19527 (N_19527,N_16774,N_15859);
nor U19528 (N_19528,N_17409,N_16694);
and U19529 (N_19529,N_16724,N_15048);
nor U19530 (N_19530,N_16113,N_16602);
nand U19531 (N_19531,N_16997,N_15593);
and U19532 (N_19532,N_16756,N_17187);
xor U19533 (N_19533,N_15297,N_16491);
nor U19534 (N_19534,N_15390,N_15590);
or U19535 (N_19535,N_16148,N_15887);
or U19536 (N_19536,N_16159,N_16009);
and U19537 (N_19537,N_15563,N_17267);
and U19538 (N_19538,N_15682,N_16449);
and U19539 (N_19539,N_16415,N_16494);
or U19540 (N_19540,N_17130,N_15709);
and U19541 (N_19541,N_16948,N_16979);
and U19542 (N_19542,N_15459,N_16408);
nand U19543 (N_19543,N_17260,N_17433);
and U19544 (N_19544,N_15884,N_17272);
or U19545 (N_19545,N_16307,N_15128);
and U19546 (N_19546,N_16072,N_15884);
nor U19547 (N_19547,N_15572,N_16334);
and U19548 (N_19548,N_16698,N_15939);
and U19549 (N_19549,N_16428,N_16091);
and U19550 (N_19550,N_15842,N_16608);
xnor U19551 (N_19551,N_16096,N_16524);
or U19552 (N_19552,N_17171,N_16116);
and U19553 (N_19553,N_15476,N_17128);
xnor U19554 (N_19554,N_17497,N_16505);
nor U19555 (N_19555,N_15761,N_15782);
nor U19556 (N_19556,N_15686,N_15620);
or U19557 (N_19557,N_15349,N_15490);
and U19558 (N_19558,N_17041,N_16807);
nand U19559 (N_19559,N_17081,N_16880);
and U19560 (N_19560,N_16322,N_16522);
xnor U19561 (N_19561,N_15101,N_15618);
and U19562 (N_19562,N_17258,N_15430);
nor U19563 (N_19563,N_16838,N_16682);
and U19564 (N_19564,N_17112,N_16148);
and U19565 (N_19565,N_15084,N_15159);
xor U19566 (N_19566,N_17000,N_17424);
xnor U19567 (N_19567,N_16095,N_15066);
and U19568 (N_19568,N_16102,N_15782);
and U19569 (N_19569,N_17067,N_16841);
and U19570 (N_19570,N_16273,N_16208);
and U19571 (N_19571,N_16154,N_16638);
nor U19572 (N_19572,N_16799,N_17443);
nor U19573 (N_19573,N_16529,N_16818);
or U19574 (N_19574,N_17455,N_15543);
and U19575 (N_19575,N_16950,N_15676);
nor U19576 (N_19576,N_15958,N_17065);
and U19577 (N_19577,N_15089,N_15574);
nor U19578 (N_19578,N_17366,N_15694);
xnor U19579 (N_19579,N_15661,N_16829);
or U19580 (N_19580,N_15519,N_17198);
nor U19581 (N_19581,N_15001,N_15818);
xor U19582 (N_19582,N_15045,N_15308);
xor U19583 (N_19583,N_16744,N_15757);
xnor U19584 (N_19584,N_15496,N_16451);
nand U19585 (N_19585,N_16472,N_16940);
or U19586 (N_19586,N_16977,N_15273);
nor U19587 (N_19587,N_16647,N_15792);
and U19588 (N_19588,N_15946,N_16579);
or U19589 (N_19589,N_16213,N_15536);
xor U19590 (N_19590,N_15928,N_15536);
nand U19591 (N_19591,N_16918,N_17336);
and U19592 (N_19592,N_15157,N_15769);
nand U19593 (N_19593,N_16389,N_17114);
or U19594 (N_19594,N_15350,N_16958);
xor U19595 (N_19595,N_15392,N_17092);
or U19596 (N_19596,N_16951,N_16047);
or U19597 (N_19597,N_16470,N_17065);
nand U19598 (N_19598,N_17165,N_16183);
nor U19599 (N_19599,N_15111,N_16419);
or U19600 (N_19600,N_15129,N_16106);
nor U19601 (N_19601,N_16239,N_15202);
and U19602 (N_19602,N_16482,N_15029);
and U19603 (N_19603,N_16336,N_16245);
and U19604 (N_19604,N_15553,N_15307);
nor U19605 (N_19605,N_16348,N_16491);
xor U19606 (N_19606,N_16646,N_16872);
nand U19607 (N_19607,N_15257,N_15287);
nor U19608 (N_19608,N_16372,N_17136);
nor U19609 (N_19609,N_16872,N_16891);
xor U19610 (N_19610,N_15557,N_17468);
nand U19611 (N_19611,N_16139,N_16699);
xnor U19612 (N_19612,N_17233,N_17192);
xor U19613 (N_19613,N_16714,N_15880);
nand U19614 (N_19614,N_17105,N_15065);
nand U19615 (N_19615,N_16948,N_15140);
nor U19616 (N_19616,N_15431,N_17415);
and U19617 (N_19617,N_17260,N_16115);
nand U19618 (N_19618,N_15397,N_16128);
and U19619 (N_19619,N_16856,N_16628);
nor U19620 (N_19620,N_15533,N_16025);
xor U19621 (N_19621,N_15307,N_16501);
and U19622 (N_19622,N_16911,N_15976);
nand U19623 (N_19623,N_16122,N_16985);
and U19624 (N_19624,N_15447,N_15648);
or U19625 (N_19625,N_15162,N_15577);
nor U19626 (N_19626,N_15528,N_16334);
xnor U19627 (N_19627,N_15972,N_16810);
nand U19628 (N_19628,N_17097,N_16484);
nor U19629 (N_19629,N_16966,N_16643);
or U19630 (N_19630,N_16652,N_16260);
nor U19631 (N_19631,N_15713,N_16873);
or U19632 (N_19632,N_16608,N_15495);
xor U19633 (N_19633,N_17245,N_16577);
or U19634 (N_19634,N_17323,N_17124);
xnor U19635 (N_19635,N_15076,N_15327);
or U19636 (N_19636,N_15288,N_16419);
xnor U19637 (N_19637,N_17015,N_15364);
nor U19638 (N_19638,N_16108,N_15546);
nand U19639 (N_19639,N_15486,N_17254);
nor U19640 (N_19640,N_15859,N_17378);
nand U19641 (N_19641,N_15267,N_15060);
nand U19642 (N_19642,N_16500,N_15904);
nand U19643 (N_19643,N_15222,N_16028);
nand U19644 (N_19644,N_17352,N_16178);
nor U19645 (N_19645,N_15127,N_17272);
or U19646 (N_19646,N_17239,N_15880);
xor U19647 (N_19647,N_15701,N_16122);
nor U19648 (N_19648,N_16289,N_15079);
or U19649 (N_19649,N_15562,N_16638);
and U19650 (N_19650,N_16181,N_16865);
or U19651 (N_19651,N_17237,N_16507);
nor U19652 (N_19652,N_15622,N_15534);
and U19653 (N_19653,N_16473,N_16759);
and U19654 (N_19654,N_15687,N_16301);
and U19655 (N_19655,N_15854,N_16317);
and U19656 (N_19656,N_16658,N_15679);
nor U19657 (N_19657,N_16664,N_15917);
or U19658 (N_19658,N_15112,N_15383);
xnor U19659 (N_19659,N_16912,N_16977);
nand U19660 (N_19660,N_15598,N_15139);
nand U19661 (N_19661,N_16094,N_17199);
or U19662 (N_19662,N_16513,N_16907);
nand U19663 (N_19663,N_16768,N_15280);
or U19664 (N_19664,N_15521,N_16660);
nor U19665 (N_19665,N_15984,N_15202);
or U19666 (N_19666,N_16848,N_17117);
nand U19667 (N_19667,N_16029,N_16489);
nand U19668 (N_19668,N_15304,N_16470);
and U19669 (N_19669,N_16299,N_15365);
or U19670 (N_19670,N_15109,N_15738);
and U19671 (N_19671,N_16080,N_17179);
and U19672 (N_19672,N_16269,N_15296);
nand U19673 (N_19673,N_15404,N_17106);
or U19674 (N_19674,N_17220,N_15970);
nor U19675 (N_19675,N_15611,N_15311);
xnor U19676 (N_19676,N_16929,N_17226);
or U19677 (N_19677,N_16300,N_16013);
nand U19678 (N_19678,N_15146,N_16152);
nand U19679 (N_19679,N_15232,N_16393);
nand U19680 (N_19680,N_15438,N_15067);
and U19681 (N_19681,N_17199,N_16425);
or U19682 (N_19682,N_15917,N_16173);
and U19683 (N_19683,N_15097,N_16262);
nand U19684 (N_19684,N_15960,N_16510);
nor U19685 (N_19685,N_16601,N_17171);
nor U19686 (N_19686,N_17339,N_16333);
nand U19687 (N_19687,N_16610,N_16047);
and U19688 (N_19688,N_17177,N_16390);
nand U19689 (N_19689,N_16173,N_16366);
or U19690 (N_19690,N_15809,N_16694);
nand U19691 (N_19691,N_16700,N_16582);
xor U19692 (N_19692,N_15454,N_16390);
and U19693 (N_19693,N_16251,N_16539);
or U19694 (N_19694,N_17062,N_16082);
or U19695 (N_19695,N_15901,N_15398);
or U19696 (N_19696,N_15228,N_16338);
and U19697 (N_19697,N_15032,N_15383);
xnor U19698 (N_19698,N_16196,N_15685);
nor U19699 (N_19699,N_16314,N_16544);
or U19700 (N_19700,N_15475,N_16039);
and U19701 (N_19701,N_17180,N_15303);
nand U19702 (N_19702,N_16077,N_15979);
nor U19703 (N_19703,N_15161,N_16500);
or U19704 (N_19704,N_15207,N_16093);
or U19705 (N_19705,N_15920,N_16175);
xnor U19706 (N_19706,N_15375,N_15560);
nand U19707 (N_19707,N_15975,N_17169);
nand U19708 (N_19708,N_15197,N_16883);
xor U19709 (N_19709,N_16330,N_15674);
and U19710 (N_19710,N_15925,N_15061);
and U19711 (N_19711,N_17087,N_16468);
nor U19712 (N_19712,N_15332,N_16048);
nand U19713 (N_19713,N_16504,N_17441);
nand U19714 (N_19714,N_15724,N_15810);
nor U19715 (N_19715,N_15735,N_16754);
xor U19716 (N_19716,N_16643,N_17226);
or U19717 (N_19717,N_16546,N_16768);
or U19718 (N_19718,N_15514,N_16861);
and U19719 (N_19719,N_16363,N_15260);
nor U19720 (N_19720,N_15518,N_17219);
xnor U19721 (N_19721,N_16936,N_15924);
nor U19722 (N_19722,N_15291,N_16740);
and U19723 (N_19723,N_16685,N_16124);
nand U19724 (N_19724,N_16075,N_16707);
and U19725 (N_19725,N_15019,N_15830);
xnor U19726 (N_19726,N_16632,N_15773);
xnor U19727 (N_19727,N_17235,N_15587);
and U19728 (N_19728,N_17053,N_15459);
xnor U19729 (N_19729,N_15804,N_15525);
nand U19730 (N_19730,N_16241,N_17282);
xnor U19731 (N_19731,N_15744,N_15296);
and U19732 (N_19732,N_16347,N_16063);
xnor U19733 (N_19733,N_16561,N_15451);
and U19734 (N_19734,N_17216,N_15736);
or U19735 (N_19735,N_16212,N_15870);
nor U19736 (N_19736,N_15280,N_15746);
nand U19737 (N_19737,N_16017,N_15623);
nand U19738 (N_19738,N_16854,N_15415);
and U19739 (N_19739,N_15517,N_16720);
or U19740 (N_19740,N_17453,N_16374);
or U19741 (N_19741,N_15521,N_17033);
and U19742 (N_19742,N_16418,N_15853);
or U19743 (N_19743,N_16552,N_16600);
xnor U19744 (N_19744,N_17103,N_16461);
and U19745 (N_19745,N_15482,N_15693);
xnor U19746 (N_19746,N_15382,N_16743);
nand U19747 (N_19747,N_16959,N_16444);
nand U19748 (N_19748,N_15327,N_16527);
nand U19749 (N_19749,N_15633,N_16434);
or U19750 (N_19750,N_16602,N_15198);
nor U19751 (N_19751,N_17143,N_15812);
and U19752 (N_19752,N_17194,N_17431);
and U19753 (N_19753,N_15420,N_16186);
and U19754 (N_19754,N_15655,N_16892);
xor U19755 (N_19755,N_15539,N_17423);
xnor U19756 (N_19756,N_15265,N_15537);
xor U19757 (N_19757,N_16601,N_15695);
xnor U19758 (N_19758,N_16456,N_15426);
nand U19759 (N_19759,N_15033,N_16842);
or U19760 (N_19760,N_16553,N_15940);
xor U19761 (N_19761,N_16041,N_16801);
xor U19762 (N_19762,N_16025,N_16373);
nor U19763 (N_19763,N_17271,N_17480);
nor U19764 (N_19764,N_16477,N_17169);
nand U19765 (N_19765,N_15595,N_15082);
nor U19766 (N_19766,N_16936,N_16333);
xnor U19767 (N_19767,N_17125,N_17324);
xnor U19768 (N_19768,N_15422,N_15717);
nor U19769 (N_19769,N_15033,N_16722);
xnor U19770 (N_19770,N_15051,N_17477);
nand U19771 (N_19771,N_15298,N_17008);
xnor U19772 (N_19772,N_16402,N_16199);
xnor U19773 (N_19773,N_16858,N_15874);
nor U19774 (N_19774,N_15798,N_15955);
nand U19775 (N_19775,N_15304,N_17248);
nand U19776 (N_19776,N_17107,N_16025);
and U19777 (N_19777,N_15548,N_15766);
xnor U19778 (N_19778,N_17273,N_15180);
nand U19779 (N_19779,N_17345,N_17170);
xor U19780 (N_19780,N_15067,N_15788);
xnor U19781 (N_19781,N_16743,N_16264);
or U19782 (N_19782,N_15759,N_15236);
nand U19783 (N_19783,N_17438,N_15091);
nand U19784 (N_19784,N_15781,N_15424);
nor U19785 (N_19785,N_16218,N_15920);
nor U19786 (N_19786,N_15364,N_15280);
and U19787 (N_19787,N_15371,N_16380);
xnor U19788 (N_19788,N_15152,N_15034);
xnor U19789 (N_19789,N_15600,N_15787);
nor U19790 (N_19790,N_17093,N_15338);
or U19791 (N_19791,N_15688,N_16115);
nand U19792 (N_19792,N_17212,N_15791);
nand U19793 (N_19793,N_17012,N_16492);
nand U19794 (N_19794,N_15779,N_15692);
nand U19795 (N_19795,N_16211,N_15604);
nand U19796 (N_19796,N_15836,N_15135);
and U19797 (N_19797,N_16039,N_15160);
nand U19798 (N_19798,N_15289,N_15482);
and U19799 (N_19799,N_16917,N_15482);
xor U19800 (N_19800,N_15821,N_15149);
nor U19801 (N_19801,N_17053,N_15411);
or U19802 (N_19802,N_15516,N_16214);
xnor U19803 (N_19803,N_17469,N_15040);
nor U19804 (N_19804,N_16311,N_16166);
nor U19805 (N_19805,N_15198,N_16126);
or U19806 (N_19806,N_16635,N_16868);
nand U19807 (N_19807,N_15918,N_15753);
xor U19808 (N_19808,N_16537,N_17413);
xor U19809 (N_19809,N_16377,N_16020);
nand U19810 (N_19810,N_15685,N_15812);
and U19811 (N_19811,N_15877,N_15739);
and U19812 (N_19812,N_15849,N_15769);
and U19813 (N_19813,N_15356,N_17122);
nand U19814 (N_19814,N_16637,N_15067);
nand U19815 (N_19815,N_16755,N_16688);
nor U19816 (N_19816,N_15063,N_16742);
nor U19817 (N_19817,N_16740,N_15901);
xor U19818 (N_19818,N_16016,N_15152);
xor U19819 (N_19819,N_16085,N_15711);
xor U19820 (N_19820,N_16281,N_15679);
nand U19821 (N_19821,N_15392,N_16462);
nor U19822 (N_19822,N_15423,N_17063);
nand U19823 (N_19823,N_15812,N_16529);
nor U19824 (N_19824,N_16918,N_16151);
xnor U19825 (N_19825,N_16791,N_15844);
nand U19826 (N_19826,N_16108,N_15964);
and U19827 (N_19827,N_16326,N_16915);
and U19828 (N_19828,N_15829,N_16233);
or U19829 (N_19829,N_15548,N_17322);
and U19830 (N_19830,N_17190,N_17204);
nand U19831 (N_19831,N_15721,N_17350);
and U19832 (N_19832,N_15737,N_17199);
xor U19833 (N_19833,N_16497,N_16396);
and U19834 (N_19834,N_16064,N_16326);
nand U19835 (N_19835,N_15580,N_17337);
nor U19836 (N_19836,N_16828,N_15372);
xor U19837 (N_19837,N_17300,N_16657);
xnor U19838 (N_19838,N_15280,N_17042);
and U19839 (N_19839,N_15921,N_16412);
and U19840 (N_19840,N_16491,N_16384);
nor U19841 (N_19841,N_16947,N_15501);
or U19842 (N_19842,N_15088,N_16737);
xor U19843 (N_19843,N_15261,N_15169);
nor U19844 (N_19844,N_16936,N_15173);
xor U19845 (N_19845,N_16502,N_15005);
nor U19846 (N_19846,N_17324,N_16535);
xor U19847 (N_19847,N_17154,N_17321);
xor U19848 (N_19848,N_17288,N_16079);
and U19849 (N_19849,N_16692,N_15233);
or U19850 (N_19850,N_15468,N_17272);
nand U19851 (N_19851,N_17124,N_16189);
nand U19852 (N_19852,N_15000,N_17246);
nor U19853 (N_19853,N_17448,N_15259);
nor U19854 (N_19854,N_16574,N_17498);
and U19855 (N_19855,N_17105,N_17154);
and U19856 (N_19856,N_16512,N_17224);
xnor U19857 (N_19857,N_15904,N_16792);
nand U19858 (N_19858,N_16976,N_16370);
and U19859 (N_19859,N_16123,N_16709);
and U19860 (N_19860,N_15465,N_17149);
xor U19861 (N_19861,N_15565,N_15016);
and U19862 (N_19862,N_17126,N_17165);
nor U19863 (N_19863,N_15891,N_15169);
nand U19864 (N_19864,N_15523,N_17379);
or U19865 (N_19865,N_17384,N_15334);
and U19866 (N_19866,N_15885,N_15913);
and U19867 (N_19867,N_15228,N_17197);
nand U19868 (N_19868,N_15766,N_16061);
nor U19869 (N_19869,N_16246,N_15185);
nand U19870 (N_19870,N_15160,N_16215);
nor U19871 (N_19871,N_17495,N_15377);
or U19872 (N_19872,N_16034,N_15126);
xnor U19873 (N_19873,N_15662,N_15895);
nand U19874 (N_19874,N_15684,N_17013);
nor U19875 (N_19875,N_17166,N_15756);
nand U19876 (N_19876,N_16741,N_15352);
or U19877 (N_19877,N_17352,N_17097);
nand U19878 (N_19878,N_15330,N_15414);
and U19879 (N_19879,N_16975,N_15996);
or U19880 (N_19880,N_15719,N_16332);
nand U19881 (N_19881,N_16633,N_17369);
xnor U19882 (N_19882,N_16484,N_15166);
nor U19883 (N_19883,N_15279,N_15200);
nor U19884 (N_19884,N_16783,N_16032);
nand U19885 (N_19885,N_16255,N_16100);
and U19886 (N_19886,N_16727,N_16434);
xnor U19887 (N_19887,N_16028,N_16639);
nor U19888 (N_19888,N_17497,N_15605);
or U19889 (N_19889,N_15099,N_15942);
nand U19890 (N_19890,N_15878,N_17404);
nor U19891 (N_19891,N_16234,N_15724);
nor U19892 (N_19892,N_16855,N_16430);
xnor U19893 (N_19893,N_17296,N_15377);
nand U19894 (N_19894,N_16315,N_16512);
and U19895 (N_19895,N_16224,N_16863);
xnor U19896 (N_19896,N_16302,N_16630);
or U19897 (N_19897,N_15508,N_15267);
xnor U19898 (N_19898,N_16396,N_17316);
xor U19899 (N_19899,N_16717,N_16007);
and U19900 (N_19900,N_17409,N_15588);
xor U19901 (N_19901,N_15165,N_15458);
nand U19902 (N_19902,N_15618,N_15871);
nand U19903 (N_19903,N_15276,N_16454);
xnor U19904 (N_19904,N_17248,N_16392);
and U19905 (N_19905,N_17383,N_16854);
nand U19906 (N_19906,N_15484,N_16150);
and U19907 (N_19907,N_16354,N_16950);
and U19908 (N_19908,N_16196,N_16498);
and U19909 (N_19909,N_16864,N_15007);
nor U19910 (N_19910,N_17141,N_17018);
xnor U19911 (N_19911,N_17020,N_16025);
and U19912 (N_19912,N_16415,N_16893);
xor U19913 (N_19913,N_16793,N_16962);
nand U19914 (N_19914,N_16071,N_15785);
nor U19915 (N_19915,N_17236,N_17376);
xnor U19916 (N_19916,N_15238,N_17042);
xnor U19917 (N_19917,N_16008,N_16463);
or U19918 (N_19918,N_15596,N_16603);
nor U19919 (N_19919,N_15008,N_15588);
nand U19920 (N_19920,N_16337,N_16517);
and U19921 (N_19921,N_17156,N_15895);
nor U19922 (N_19922,N_15217,N_15942);
nand U19923 (N_19923,N_15299,N_15653);
nor U19924 (N_19924,N_17154,N_16711);
nand U19925 (N_19925,N_16709,N_15587);
xnor U19926 (N_19926,N_15767,N_17289);
or U19927 (N_19927,N_16492,N_17162);
nand U19928 (N_19928,N_16897,N_15463);
nor U19929 (N_19929,N_16787,N_17240);
nand U19930 (N_19930,N_16118,N_16369);
nand U19931 (N_19931,N_16717,N_16536);
nor U19932 (N_19932,N_15881,N_15834);
and U19933 (N_19933,N_15056,N_15592);
nand U19934 (N_19934,N_17343,N_15126);
and U19935 (N_19935,N_17117,N_15231);
or U19936 (N_19936,N_15930,N_15621);
xnor U19937 (N_19937,N_16278,N_16034);
and U19938 (N_19938,N_15812,N_16166);
and U19939 (N_19939,N_17048,N_16644);
nand U19940 (N_19940,N_17222,N_15401);
or U19941 (N_19941,N_16358,N_15382);
xnor U19942 (N_19942,N_17211,N_16181);
and U19943 (N_19943,N_16060,N_15482);
and U19944 (N_19944,N_16559,N_15491);
xnor U19945 (N_19945,N_17380,N_16413);
nand U19946 (N_19946,N_15973,N_16602);
nand U19947 (N_19947,N_16869,N_16419);
nand U19948 (N_19948,N_16760,N_16557);
xnor U19949 (N_19949,N_16681,N_15032);
or U19950 (N_19950,N_16516,N_15963);
and U19951 (N_19951,N_15374,N_15091);
and U19952 (N_19952,N_16626,N_16097);
and U19953 (N_19953,N_17068,N_15183);
and U19954 (N_19954,N_17423,N_16826);
or U19955 (N_19955,N_17397,N_16565);
and U19956 (N_19956,N_16765,N_16377);
nand U19957 (N_19957,N_15307,N_16648);
nor U19958 (N_19958,N_15388,N_17152);
xnor U19959 (N_19959,N_15807,N_17070);
and U19960 (N_19960,N_16530,N_17158);
or U19961 (N_19961,N_16227,N_15752);
nor U19962 (N_19962,N_17107,N_15424);
nor U19963 (N_19963,N_15444,N_15477);
and U19964 (N_19964,N_16563,N_16050);
xnor U19965 (N_19965,N_17387,N_16563);
nand U19966 (N_19966,N_17492,N_15806);
nand U19967 (N_19967,N_15042,N_17113);
nand U19968 (N_19968,N_15162,N_15044);
nand U19969 (N_19969,N_16173,N_16663);
nor U19970 (N_19970,N_16096,N_15878);
nor U19971 (N_19971,N_15732,N_15827);
nand U19972 (N_19972,N_16598,N_16221);
or U19973 (N_19973,N_15695,N_16407);
or U19974 (N_19974,N_16204,N_16431);
xor U19975 (N_19975,N_16397,N_15184);
and U19976 (N_19976,N_16244,N_17039);
nor U19977 (N_19977,N_17131,N_15287);
nand U19978 (N_19978,N_16796,N_17215);
and U19979 (N_19979,N_15664,N_15322);
and U19980 (N_19980,N_15076,N_16461);
or U19981 (N_19981,N_15150,N_16139);
nand U19982 (N_19982,N_16238,N_17314);
nand U19983 (N_19983,N_15760,N_15255);
xor U19984 (N_19984,N_17170,N_16828);
or U19985 (N_19985,N_16367,N_15894);
and U19986 (N_19986,N_15973,N_15217);
nor U19987 (N_19987,N_16228,N_15055);
or U19988 (N_19988,N_15221,N_16529);
and U19989 (N_19989,N_15911,N_16429);
nor U19990 (N_19990,N_15460,N_16529);
and U19991 (N_19991,N_16858,N_16574);
nand U19992 (N_19992,N_16810,N_16598);
nor U19993 (N_19993,N_16579,N_17470);
xor U19994 (N_19994,N_16821,N_15176);
and U19995 (N_19995,N_17371,N_16211);
xnor U19996 (N_19996,N_15187,N_15742);
nor U19997 (N_19997,N_15382,N_16836);
nor U19998 (N_19998,N_16829,N_16306);
and U19999 (N_19999,N_16370,N_17488);
nor U20000 (N_20000,N_19012,N_19103);
nand U20001 (N_20001,N_17856,N_17719);
and U20002 (N_20002,N_19604,N_19701);
nor U20003 (N_20003,N_19951,N_19430);
and U20004 (N_20004,N_18491,N_19128);
nor U20005 (N_20005,N_18978,N_19227);
xor U20006 (N_20006,N_19585,N_19337);
nor U20007 (N_20007,N_18734,N_17620);
nor U20008 (N_20008,N_19613,N_19184);
nor U20009 (N_20009,N_18932,N_19733);
xnor U20010 (N_20010,N_17544,N_18582);
and U20011 (N_20011,N_19414,N_18028);
nand U20012 (N_20012,N_19026,N_18051);
or U20013 (N_20013,N_18435,N_19727);
nor U20014 (N_20014,N_18164,N_18276);
and U20015 (N_20015,N_19299,N_19856);
and U20016 (N_20016,N_19794,N_19191);
nor U20017 (N_20017,N_17823,N_19519);
xnor U20018 (N_20018,N_18090,N_18778);
xor U20019 (N_20019,N_18065,N_18887);
nand U20020 (N_20020,N_19360,N_19922);
nor U20021 (N_20021,N_18635,N_18528);
xor U20022 (N_20022,N_19446,N_18976);
or U20023 (N_20023,N_19106,N_19135);
nor U20024 (N_20024,N_19435,N_19488);
nand U20025 (N_20025,N_19441,N_18686);
or U20026 (N_20026,N_19837,N_18705);
xor U20027 (N_20027,N_18257,N_18063);
nor U20028 (N_20028,N_19901,N_17597);
xnor U20029 (N_20029,N_17560,N_19217);
nand U20030 (N_20030,N_19882,N_19054);
nand U20031 (N_20031,N_19405,N_17899);
or U20032 (N_20032,N_19551,N_17523);
nor U20033 (N_20033,N_18977,N_17845);
nand U20034 (N_20034,N_17642,N_17783);
nand U20035 (N_20035,N_17501,N_18747);
and U20036 (N_20036,N_19208,N_18071);
nand U20037 (N_20037,N_19316,N_18833);
and U20038 (N_20038,N_19445,N_18758);
nand U20039 (N_20039,N_17502,N_19174);
nand U20040 (N_20040,N_19900,N_18264);
xor U20041 (N_20041,N_19529,N_19437);
xnor U20042 (N_20042,N_19828,N_17881);
xor U20043 (N_20043,N_19830,N_19603);
nand U20044 (N_20044,N_18263,N_19630);
xor U20045 (N_20045,N_17584,N_18757);
or U20046 (N_20046,N_18658,N_18406);
xor U20047 (N_20047,N_19472,N_17741);
xor U20048 (N_20048,N_17831,N_17649);
or U20049 (N_20049,N_17759,N_19980);
nand U20050 (N_20050,N_19835,N_18381);
nor U20051 (N_20051,N_18768,N_19561);
xnor U20052 (N_20052,N_19996,N_19530);
and U20053 (N_20053,N_18606,N_17655);
xor U20054 (N_20054,N_18692,N_18238);
or U20055 (N_20055,N_18323,N_17825);
nand U20056 (N_20056,N_18846,N_19760);
nor U20057 (N_20057,N_19100,N_19974);
or U20058 (N_20058,N_19332,N_18086);
or U20059 (N_20059,N_19817,N_19018);
and U20060 (N_20060,N_19237,N_17706);
nand U20061 (N_20061,N_18810,N_17768);
nand U20062 (N_20062,N_19508,N_18564);
nor U20063 (N_20063,N_19489,N_18300);
nand U20064 (N_20064,N_19089,N_18313);
nor U20065 (N_20065,N_19984,N_18001);
xor U20066 (N_20066,N_18923,N_18600);
or U20067 (N_20067,N_17808,N_18183);
nor U20068 (N_20068,N_19321,N_17625);
nor U20069 (N_20069,N_19612,N_19444);
and U20070 (N_20070,N_19627,N_18842);
xor U20071 (N_20071,N_18973,N_18384);
nand U20072 (N_20072,N_19411,N_17563);
nand U20073 (N_20073,N_18645,N_18219);
and U20074 (N_20074,N_19496,N_19595);
nand U20075 (N_20075,N_19077,N_18785);
or U20076 (N_20076,N_18530,N_18291);
or U20077 (N_20077,N_19214,N_18542);
or U20078 (N_20078,N_17636,N_18558);
xor U20079 (N_20079,N_19861,N_18492);
nand U20080 (N_20080,N_17925,N_18649);
and U20081 (N_20081,N_17593,N_19156);
nand U20082 (N_20082,N_19243,N_17959);
xnor U20083 (N_20083,N_19509,N_19206);
or U20084 (N_20084,N_18270,N_19544);
or U20085 (N_20085,N_18037,N_18287);
nor U20086 (N_20086,N_18819,N_18557);
nand U20087 (N_20087,N_17628,N_18460);
nor U20088 (N_20088,N_18925,N_19300);
nor U20089 (N_20089,N_18548,N_17911);
nor U20090 (N_20090,N_17954,N_19200);
or U20091 (N_20091,N_19873,N_19049);
nor U20092 (N_20092,N_18652,N_17772);
nand U20093 (N_20093,N_18822,N_18898);
or U20094 (N_20094,N_19824,N_19578);
nand U20095 (N_20095,N_19201,N_19847);
or U20096 (N_20096,N_19897,N_19236);
nor U20097 (N_20097,N_19678,N_18911);
xnor U20098 (N_20098,N_19165,N_18428);
and U20099 (N_20099,N_17851,N_19306);
or U20100 (N_20100,N_19718,N_19312);
nand U20101 (N_20101,N_17773,N_19550);
xor U20102 (N_20102,N_19254,N_18275);
or U20103 (N_20103,N_17562,N_19584);
or U20104 (N_20104,N_19110,N_17503);
nand U20105 (N_20105,N_19057,N_19129);
or U20106 (N_20106,N_19914,N_19563);
or U20107 (N_20107,N_18870,N_19173);
or U20108 (N_20108,N_19891,N_19916);
and U20109 (N_20109,N_19231,N_17529);
nor U20110 (N_20110,N_18117,N_18500);
nor U20111 (N_20111,N_19015,N_17777);
nand U20112 (N_20112,N_18958,N_19849);
nand U20113 (N_20113,N_18578,N_18707);
nor U20114 (N_20114,N_18472,N_19044);
nand U20115 (N_20115,N_18029,N_18902);
or U20116 (N_20116,N_17952,N_19759);
nor U20117 (N_20117,N_18943,N_18912);
nand U20118 (N_20118,N_17565,N_19566);
and U20119 (N_20119,N_19786,N_19216);
nor U20120 (N_20120,N_19674,N_18620);
xnor U20121 (N_20121,N_19687,N_19671);
or U20122 (N_20122,N_17608,N_18084);
nand U20123 (N_20123,N_18788,N_18163);
xnor U20124 (N_20124,N_17530,N_19634);
xor U20125 (N_20125,N_18807,N_18538);
nor U20126 (N_20126,N_18505,N_18191);
and U20127 (N_20127,N_19399,N_17550);
nor U20128 (N_20128,N_18439,N_19620);
or U20129 (N_20129,N_17985,N_19278);
and U20130 (N_20130,N_19248,N_17590);
and U20131 (N_20131,N_18688,N_17964);
nor U20132 (N_20132,N_18205,N_17585);
nand U20133 (N_20133,N_18698,N_17622);
nand U20134 (N_20134,N_17754,N_19742);
nor U20135 (N_20135,N_18279,N_19662);
and U20136 (N_20136,N_19137,N_17752);
nand U20137 (N_20137,N_19118,N_19475);
nand U20138 (N_20138,N_19862,N_18123);
nor U20139 (N_20139,N_17779,N_19815);
nor U20140 (N_20140,N_19267,N_17519);
and U20141 (N_20141,N_18229,N_18927);
xnor U20142 (N_20142,N_19543,N_17941);
xor U20143 (N_20143,N_17857,N_19463);
or U20144 (N_20144,N_19004,N_17796);
or U20145 (N_20145,N_17760,N_18585);
nor U20146 (N_20146,N_19386,N_19814);
xnor U20147 (N_20147,N_19945,N_19887);
or U20148 (N_20148,N_19999,N_19281);
nand U20149 (N_20149,N_19571,N_17824);
or U20150 (N_20150,N_19518,N_18610);
xor U20151 (N_20151,N_17533,N_19654);
nand U20152 (N_20152,N_19436,N_19601);
or U20153 (N_20153,N_18333,N_18507);
or U20154 (N_20154,N_18162,N_19498);
nand U20155 (N_20155,N_19130,N_18465);
xnor U20156 (N_20156,N_18345,N_19669);
xor U20157 (N_20157,N_19136,N_19064);
nand U20158 (N_20158,N_18572,N_18240);
nor U20159 (N_20159,N_18653,N_18498);
nor U20160 (N_20160,N_18702,N_17929);
xor U20161 (N_20161,N_19774,N_19829);
xnor U20162 (N_20162,N_19164,N_18856);
nand U20163 (N_20163,N_19481,N_19765);
and U20164 (N_20164,N_18827,N_19749);
nor U20165 (N_20165,N_18242,N_18952);
nand U20166 (N_20166,N_19942,N_19473);
xnor U20167 (N_20167,N_18933,N_19694);
or U20168 (N_20168,N_18659,N_17897);
nor U20169 (N_20169,N_17787,N_19908);
nand U20170 (N_20170,N_17835,N_19607);
and U20171 (N_20171,N_19176,N_19697);
nand U20172 (N_20172,N_18105,N_19597);
nand U20173 (N_20173,N_18330,N_18170);
nor U20174 (N_20174,N_19389,N_18249);
and U20175 (N_20175,N_17663,N_18203);
and U20176 (N_20176,N_17898,N_19238);
nor U20177 (N_20177,N_18125,N_17506);
and U20178 (N_20178,N_18178,N_18012);
nor U20179 (N_20179,N_18825,N_18996);
nand U20180 (N_20180,N_17748,N_19875);
nand U20181 (N_20181,N_17589,N_18357);
nor U20182 (N_20182,N_18109,N_18258);
nand U20183 (N_20183,N_19286,N_17886);
nand U20184 (N_20184,N_17617,N_18751);
or U20185 (N_20185,N_17861,N_17974);
and U20186 (N_20186,N_18875,N_17686);
nand U20187 (N_20187,N_19113,N_18244);
or U20188 (N_20188,N_18399,N_18231);
nand U20189 (N_20189,N_19717,N_19123);
and U20190 (N_20190,N_18871,N_19767);
nor U20191 (N_20191,N_19703,N_18780);
nor U20192 (N_20192,N_18383,N_19808);
nand U20193 (N_20193,N_18614,N_17666);
nand U20194 (N_20194,N_17871,N_19677);
xnor U20195 (N_20195,N_17609,N_19894);
or U20196 (N_20196,N_18717,N_18389);
and U20197 (N_20197,N_19284,N_19482);
nand U20198 (N_20198,N_19071,N_19290);
or U20199 (N_20199,N_18536,N_17551);
and U20200 (N_20200,N_17721,N_18963);
xnor U20201 (N_20201,N_19138,N_18391);
or U20202 (N_20202,N_19259,N_19741);
nor U20203 (N_20203,N_18941,N_18022);
nand U20204 (N_20204,N_18294,N_18760);
xnor U20205 (N_20205,N_19329,N_18643);
and U20206 (N_20206,N_18742,N_19981);
xnor U20207 (N_20207,N_18277,N_19081);
nand U20208 (N_20208,N_19361,N_19415);
xor U20209 (N_20209,N_18867,N_19143);
or U20210 (N_20210,N_18803,N_17943);
and U20211 (N_20211,N_18395,N_19338);
nor U20212 (N_20212,N_19960,N_19953);
nor U20213 (N_20213,N_18031,N_18718);
nand U20214 (N_20214,N_19085,N_17801);
nand U20215 (N_20215,N_18451,N_19624);
and U20216 (N_20216,N_19573,N_18550);
xor U20217 (N_20217,N_18302,N_18743);
nand U20218 (N_20218,N_19426,N_19258);
xor U20219 (N_20219,N_19975,N_19119);
nand U20220 (N_20220,N_19852,N_19069);
xnor U20221 (N_20221,N_18618,N_18414);
and U20222 (N_20222,N_17673,N_17643);
and U20223 (N_20223,N_18306,N_18096);
nand U20224 (N_20224,N_17766,N_17958);
nand U20225 (N_20225,N_19826,N_19275);
nand U20226 (N_20226,N_18847,N_18859);
nand U20227 (N_20227,N_18408,N_18225);
or U20228 (N_20228,N_18000,N_17605);
xnor U20229 (N_20229,N_18891,N_19652);
or U20230 (N_20230,N_18570,N_17792);
and U20231 (N_20231,N_17648,N_17917);
nor U20232 (N_20232,N_17924,N_18590);
and U20233 (N_20233,N_17578,N_19531);
xnor U20234 (N_20234,N_19311,N_17664);
nor U20235 (N_20235,N_19401,N_18982);
nor U20236 (N_20236,N_19163,N_17645);
and U20237 (N_20237,N_19402,N_19594);
xnor U20238 (N_20238,N_19189,N_18672);
or U20239 (N_20239,N_18464,N_19387);
xnor U20240 (N_20240,N_18995,N_19950);
nor U20241 (N_20241,N_18915,N_17697);
or U20242 (N_20242,N_18918,N_17668);
xnor U20243 (N_20243,N_19889,N_18056);
and U20244 (N_20244,N_17803,N_18556);
nor U20245 (N_20245,N_19993,N_18657);
and U20246 (N_20246,N_17905,N_18765);
and U20247 (N_20247,N_19913,N_18047);
and U20248 (N_20248,N_18221,N_18754);
or U20249 (N_20249,N_18209,N_18454);
nor U20250 (N_20250,N_18437,N_18166);
nor U20251 (N_20251,N_19038,N_18727);
and U20252 (N_20252,N_18429,N_18104);
or U20253 (N_20253,N_18903,N_19973);
or U20254 (N_20254,N_18905,N_19845);
nand U20255 (N_20255,N_17987,N_19215);
nor U20256 (N_20256,N_19707,N_19159);
and U20257 (N_20257,N_17883,N_19379);
and U20258 (N_20258,N_19340,N_18970);
and U20259 (N_20259,N_19721,N_18188);
nand U20260 (N_20260,N_18795,N_19099);
or U20261 (N_20261,N_18685,N_18741);
nor U20262 (N_20262,N_18971,N_18896);
and U20263 (N_20263,N_19339,N_19046);
nand U20264 (N_20264,N_17726,N_17969);
nor U20265 (N_20265,N_19801,N_19858);
or U20266 (N_20266,N_19907,N_18295);
nand U20267 (N_20267,N_19255,N_19536);
and U20268 (N_20268,N_18985,N_19593);
or U20269 (N_20269,N_18093,N_18928);
or U20270 (N_20270,N_17603,N_18623);
xnor U20271 (N_20271,N_19879,N_18523);
xor U20272 (N_20272,N_19121,N_18664);
and U20273 (N_20273,N_19515,N_17576);
nor U20274 (N_20274,N_19155,N_19377);
nor U20275 (N_20275,N_19423,N_17855);
xor U20276 (N_20276,N_18850,N_19307);
nand U20277 (N_20277,N_19181,N_19649);
nor U20278 (N_20278,N_17976,N_19380);
or U20279 (N_20279,N_18514,N_19425);
xnor U20280 (N_20280,N_19068,N_17681);
or U20281 (N_20281,N_17940,N_19003);
xnor U20282 (N_20282,N_18246,N_18529);
nor U20283 (N_20283,N_19892,N_17999);
nor U20284 (N_20284,N_19149,N_19538);
and U20285 (N_20285,N_19618,N_18050);
xnor U20286 (N_20286,N_19455,N_18425);
nand U20287 (N_20287,N_18866,N_19850);
nand U20288 (N_20288,N_17580,N_18869);
nor U20289 (N_20289,N_18766,N_19079);
xnor U20290 (N_20290,N_19699,N_19520);
and U20291 (N_20291,N_19513,N_19836);
or U20292 (N_20292,N_19154,N_19395);
nor U20293 (N_20293,N_18215,N_18314);
and U20294 (N_20294,N_19785,N_19842);
or U20295 (N_20295,N_19447,N_19418);
and U20296 (N_20296,N_19366,N_17715);
xor U20297 (N_20297,N_19228,N_18272);
xor U20298 (N_20298,N_19764,N_19692);
or U20299 (N_20299,N_19151,N_19608);
nand U20300 (N_20300,N_19368,N_18380);
nand U20301 (N_20301,N_19647,N_17827);
or U20302 (N_20302,N_19196,N_17549);
nor U20303 (N_20303,N_19626,N_18210);
xnor U20304 (N_20304,N_19072,N_18501);
nand U20305 (N_20305,N_17979,N_18651);
nor U20306 (N_20306,N_18052,N_19457);
and U20307 (N_20307,N_19884,N_19588);
nand U20308 (N_20308,N_19964,N_19915);
xnor U20309 (N_20309,N_19272,N_18673);
or U20310 (N_20310,N_19883,N_18180);
nor U20311 (N_20311,N_19190,N_19797);
nand U20312 (N_20312,N_19712,N_17650);
and U20313 (N_20313,N_17699,N_18444);
xnor U20314 (N_20314,N_19170,N_19541);
xor U20315 (N_20315,N_18633,N_18604);
nor U20316 (N_20316,N_19091,N_18083);
nand U20317 (N_20317,N_18650,N_18177);
or U20318 (N_20318,N_18171,N_17908);
xor U20319 (N_20319,N_18924,N_19912);
or U20320 (N_20320,N_18390,N_19393);
nand U20321 (N_20321,N_19433,N_18715);
xor U20322 (N_20322,N_19698,N_19905);
nor U20323 (N_20323,N_17811,N_17832);
nand U20324 (N_20324,N_18248,N_17654);
nand U20325 (N_20325,N_18235,N_17504);
and U20326 (N_20326,N_18640,N_19642);
nor U20327 (N_20327,N_18331,N_18228);
nor U20328 (N_20328,N_18066,N_17505);
xor U20329 (N_20329,N_18288,N_18350);
nor U20330 (N_20330,N_18243,N_19140);
or U20331 (N_20331,N_19331,N_17880);
nor U20332 (N_20332,N_19706,N_18445);
and U20333 (N_20333,N_17938,N_17511);
and U20334 (N_20334,N_18894,N_19070);
nor U20335 (N_20335,N_19367,N_18844);
and U20336 (N_20336,N_17739,N_17631);
xor U20337 (N_20337,N_18520,N_17842);
or U20338 (N_20338,N_19806,N_19737);
nand U20339 (N_20339,N_19511,N_18811);
xnor U20340 (N_20340,N_18290,N_17630);
or U20341 (N_20341,N_17747,N_18931);
or U20342 (N_20342,N_18722,N_18865);
nand U20343 (N_20343,N_17862,N_19666);
and U20344 (N_20344,N_18363,N_18549);
nand U20345 (N_20345,N_19325,N_19169);
and U20346 (N_20346,N_17984,N_17695);
nand U20347 (N_20347,N_19632,N_18048);
nor U20348 (N_20348,N_17942,N_19280);
or U20349 (N_20349,N_18317,N_18626);
nor U20350 (N_20350,N_17579,N_18689);
nand U20351 (N_20351,N_18988,N_19714);
nand U20352 (N_20352,N_19276,N_17877);
and U20353 (N_20353,N_18617,N_19371);
nor U20354 (N_20354,N_19252,N_19709);
and U20355 (N_20355,N_19633,N_18152);
xor U20356 (N_20356,N_17966,N_17844);
xnor U20357 (N_20357,N_19179,N_18085);
or U20358 (N_20358,N_17574,N_19125);
and U20359 (N_20359,N_17646,N_18021);
or U20360 (N_20360,N_18335,N_18944);
xnor U20361 (N_20361,N_18914,N_17607);
or U20362 (N_20362,N_18254,N_18426);
xor U20363 (N_20363,N_19047,N_18592);
and U20364 (N_20364,N_17778,N_18438);
xor U20365 (N_20365,N_17710,N_18655);
nor U20366 (N_20366,N_19150,N_17534);
nand U20367 (N_20367,N_17690,N_18077);
or U20368 (N_20368,N_18237,N_19713);
and U20369 (N_20369,N_18608,N_18304);
or U20370 (N_20370,N_18457,N_19194);
or U20371 (N_20371,N_17556,N_17949);
nand U20372 (N_20372,N_19686,N_19370);
or U20373 (N_20373,N_18448,N_18509);
or U20374 (N_20374,N_19977,N_17800);
and U20375 (N_20375,N_17815,N_19670);
and U20376 (N_20376,N_18661,N_19333);
nor U20377 (N_20377,N_19723,N_18665);
or U20378 (N_20378,N_18624,N_19857);
xor U20379 (N_20379,N_17781,N_19202);
nand U20380 (N_20380,N_19895,N_17889);
and U20381 (N_20381,N_18876,N_18956);
xor U20382 (N_20382,N_18379,N_19045);
xor U20383 (N_20383,N_18946,N_17854);
xnor U20384 (N_20384,N_17716,N_18597);
or U20385 (N_20385,N_19302,N_19198);
and U20386 (N_20386,N_19141,N_18675);
or U20387 (N_20387,N_18119,N_18274);
xor U20388 (N_20388,N_19636,N_19289);
and U20389 (N_20389,N_18490,N_19577);
xnor U20390 (N_20390,N_18127,N_18034);
and U20391 (N_20391,N_18587,N_18216);
nand U20392 (N_20392,N_18857,N_18654);
nor U20393 (N_20393,N_19898,N_18443);
and U20394 (N_20394,N_17890,N_18309);
nand U20395 (N_20395,N_19598,N_17948);
nor U20396 (N_20396,N_19506,N_19590);
nand U20397 (N_20397,N_18816,N_18725);
nand U20398 (N_20398,N_18571,N_18311);
and U20399 (N_20399,N_17931,N_19735);
and U20400 (N_20400,N_17517,N_18573);
xor U20401 (N_20401,N_18212,N_19242);
and U20402 (N_20402,N_17928,N_19930);
and U20403 (N_20403,N_19833,N_19443);
or U20404 (N_20404,N_19043,N_18732);
or U20405 (N_20405,N_18292,N_17914);
or U20406 (N_20406,N_19494,N_18772);
xor U20407 (N_20407,N_19251,N_17986);
xor U20408 (N_20408,N_19462,N_19524);
and U20409 (N_20409,N_18843,N_18328);
and U20410 (N_20410,N_19985,N_18069);
nor U20411 (N_20411,N_19514,N_18415);
nor U20412 (N_20412,N_19988,N_18756);
and U20413 (N_20413,N_18186,N_18382);
and U20414 (N_20414,N_18680,N_17878);
nor U20415 (N_20415,N_17991,N_17515);
nand U20416 (N_20416,N_17713,N_19702);
and U20417 (N_20417,N_18502,N_17573);
nor U20418 (N_20418,N_18830,N_17906);
nand U20419 (N_20419,N_17960,N_17972);
nor U20420 (N_20420,N_18273,N_19568);
nor U20421 (N_20421,N_18853,N_17733);
or U20422 (N_20422,N_18139,N_19344);
and U20423 (N_20423,N_18682,N_18094);
xor U20424 (N_20424,N_19766,N_18194);
xnor U20425 (N_20425,N_19501,N_18775);
nand U20426 (N_20426,N_19024,N_19396);
or U20427 (N_20427,N_17676,N_18628);
and U20428 (N_20428,N_19998,N_19868);
and U20429 (N_20429,N_17892,N_19803);
nor U20430 (N_20430,N_19969,N_18959);
nor U20431 (N_20431,N_18910,N_17936);
and U20432 (N_20432,N_19233,N_19665);
nand U20433 (N_20433,N_19619,N_18364);
or U20434 (N_20434,N_18002,N_19075);
or U20435 (N_20435,N_18873,N_19540);
and U20436 (N_20436,N_18591,N_19458);
or U20437 (N_20437,N_19639,N_17980);
nor U20438 (N_20438,N_19664,N_17723);
nor U20439 (N_20439,N_19213,N_18082);
nor U20440 (N_20440,N_19449,N_19909);
and U20441 (N_20441,N_19693,N_18296);
or U20442 (N_20442,N_18339,N_19673);
or U20443 (N_20443,N_18883,N_18196);
and U20444 (N_20444,N_18906,N_19245);
xor U20445 (N_20445,N_19438,N_19825);
xor U20446 (N_20446,N_18569,N_19681);
nand U20447 (N_20447,N_19592,N_18005);
and U20448 (N_20448,N_18058,N_19287);
nor U20449 (N_20449,N_18080,N_18632);
xnor U20450 (N_20450,N_18115,N_19084);
nand U20451 (N_20451,N_19199,N_18336);
nor U20452 (N_20452,N_18010,N_18638);
xor U20453 (N_20453,N_18267,N_19827);
or U20454 (N_20454,N_17975,N_19050);
and U20455 (N_20455,N_19616,N_18187);
and U20456 (N_20456,N_18957,N_18478);
nand U20457 (N_20457,N_18043,N_19505);
nand U20458 (N_20458,N_19746,N_18147);
nand U20459 (N_20459,N_17750,N_18947);
and U20460 (N_20460,N_19002,N_18458);
and U20461 (N_20461,N_19350,N_19008);
xnor U20462 (N_20462,N_18561,N_19220);
and U20463 (N_20463,N_19708,N_17947);
and U20464 (N_20464,N_17957,N_18851);
and U20465 (N_20465,N_17817,N_18070);
xor U20466 (N_20466,N_18482,N_18326);
and U20467 (N_20467,N_19093,N_18407);
and U20468 (N_20468,N_19203,N_18981);
xnor U20469 (N_20469,N_18631,N_17635);
and U20470 (N_20470,N_19821,N_18806);
and U20471 (N_20471,N_19657,N_18964);
or U20472 (N_20472,N_19142,N_18567);
nor U20473 (N_20473,N_17662,N_17812);
and U20474 (N_20474,N_17627,N_18195);
nand U20475 (N_20475,N_18563,N_19989);
or U20476 (N_20476,N_19439,N_18513);
nor U20477 (N_20477,N_19863,N_19516);
nor U20478 (N_20478,N_18862,N_17882);
and U20479 (N_20479,N_17522,N_18471);
xnor U20480 (N_20480,N_19831,N_19754);
nand U20481 (N_20481,N_18220,N_18987);
nor U20482 (N_20482,N_18308,N_19111);
nand U20483 (N_20483,N_18098,N_19095);
nor U20484 (N_20484,N_19104,N_19192);
nor U20485 (N_20485,N_19838,N_19185);
and U20486 (N_20486,N_19997,N_17967);
nor U20487 (N_20487,N_17731,N_19552);
and U20488 (N_20488,N_17867,N_18159);
nand U20489 (N_20489,N_18485,N_19569);
nor U20490 (N_20490,N_19467,N_19144);
nor U20491 (N_20491,N_19471,N_19661);
or U20492 (N_20492,N_19734,N_18202);
xor U20493 (N_20493,N_18226,N_19929);
xor U20494 (N_20494,N_18551,N_17629);
or U20495 (N_20495,N_18360,N_18936);
nand U20496 (N_20496,N_17582,N_18839);
xor U20497 (N_20497,N_19105,N_18285);
and U20498 (N_20498,N_19625,N_19832);
or U20499 (N_20499,N_18088,N_17895);
or U20500 (N_20500,N_17794,N_18821);
xor U20501 (N_20501,N_18684,N_19166);
nand U20502 (N_20502,N_18033,N_19429);
and U20503 (N_20503,N_19000,N_18253);
or U20504 (N_20504,N_18792,N_19621);
nor U20505 (N_20505,N_19788,N_18813);
and U20506 (N_20506,N_17995,N_17753);
nand U20507 (N_20507,N_19326,N_17771);
nor U20508 (N_20508,N_18484,N_18255);
or U20509 (N_20509,N_17740,N_19921);
nor U20510 (N_20510,N_18452,N_19465);
or U20511 (N_20511,N_18468,N_17685);
or U20512 (N_20512,N_17640,N_18763);
or U20513 (N_20513,N_17775,N_18945);
nor U20514 (N_20514,N_19270,N_19381);
or U20515 (N_20515,N_18543,N_19187);
nand U20516 (N_20516,N_18138,N_19212);
nand U20517 (N_20517,N_18469,N_17722);
nand U20518 (N_20518,N_19959,N_19062);
or U20519 (N_20519,N_19623,N_18241);
or U20520 (N_20520,N_19027,N_19016);
nand U20521 (N_20521,N_17513,N_19517);
and U20522 (N_20522,N_17891,N_18793);
or U20523 (N_20523,N_18738,N_18544);
and U20524 (N_20524,N_17894,N_18211);
nor U20525 (N_20525,N_18128,N_19021);
and U20526 (N_20526,N_18749,N_18899);
nand U20527 (N_20527,N_19851,N_18854);
or U20528 (N_20528,N_18133,N_18895);
and U20529 (N_20529,N_19152,N_18134);
xor U20530 (N_20530,N_19087,N_19637);
or U20531 (N_20531,N_17982,N_18385);
or U20532 (N_20532,N_18179,N_17807);
nor U20533 (N_20533,N_17819,N_19055);
xnor U20534 (N_20534,N_17558,N_19704);
nor U20535 (N_20535,N_18006,N_19605);
or U20536 (N_20536,N_18124,N_19911);
or U20537 (N_20537,N_18790,N_19933);
and U20538 (N_20538,N_18662,N_18184);
or U20539 (N_20539,N_19839,N_18307);
or U20540 (N_20540,N_18344,N_19059);
nor U20541 (N_20541,N_18122,N_18753);
nor U20542 (N_20542,N_18455,N_19936);
nor U20543 (N_20543,N_17683,N_19451);
or U20544 (N_20544,N_18496,N_18983);
nor U20545 (N_20545,N_19770,N_19548);
nand U20546 (N_20546,N_17896,N_19943);
xnor U20547 (N_20547,N_19745,N_19406);
nand U20548 (N_20548,N_18808,N_19534);
nand U20549 (N_20549,N_19172,N_17919);
nor U20550 (N_20550,N_18861,N_19298);
nor U20551 (N_20551,N_18420,N_19101);
xor U20552 (N_20552,N_18731,N_18748);
or U20553 (N_20553,N_19813,N_18713);
xnor U20554 (N_20554,N_17717,N_17728);
and U20555 (N_20555,N_18190,N_18112);
nand U20556 (N_20556,N_18142,N_18319);
nand U20557 (N_20557,N_19133,N_18789);
or U20558 (N_20558,N_19266,N_19995);
nand U20559 (N_20559,N_18055,N_17552);
and U20560 (N_20560,N_19205,N_17566);
xor U20561 (N_20561,N_19188,N_19296);
nand U20562 (N_20562,N_17763,N_19586);
xnor U20563 (N_20563,N_19994,N_18297);
nand U20564 (N_20564,N_17512,N_19247);
and U20565 (N_20565,N_19263,N_19048);
nand U20566 (N_20566,N_19063,N_17828);
nor U20567 (N_20567,N_19822,N_17510);
nand U20568 (N_20568,N_19646,N_17737);
or U20569 (N_20569,N_18735,N_18840);
xnor U20570 (N_20570,N_17840,N_18271);
or U20571 (N_20571,N_18641,N_17672);
nor U20572 (N_20572,N_18260,N_17884);
and U20573 (N_20573,N_18568,N_19320);
nand U20574 (N_20574,N_19503,N_18135);
or U20575 (N_20575,N_19575,N_18516);
or U20576 (N_20576,N_17548,N_17538);
nor U20577 (N_20577,N_19351,N_19274);
xor U20578 (N_20578,N_18595,N_18365);
and U20579 (N_20579,N_19195,N_17614);
nand U20580 (N_20580,N_18036,N_18656);
nand U20581 (N_20581,N_18615,N_19609);
nor U20582 (N_20582,N_18683,N_19342);
or U20583 (N_20583,N_19291,N_17596);
nand U20584 (N_20584,N_18555,N_19581);
and U20585 (N_20585,N_19322,N_18016);
nor U20586 (N_20586,N_18213,N_19510);
nand U20587 (N_20587,N_18522,N_19768);
or U20588 (N_20588,N_18646,N_18064);
and U20589 (N_20589,N_17521,N_19116);
and U20590 (N_20590,N_19223,N_18679);
or U20591 (N_20591,N_17536,N_19240);
and U20592 (N_20592,N_18701,N_18018);
or U20593 (N_20593,N_18798,N_19617);
nor U20594 (N_20594,N_17600,N_19747);
or U20595 (N_20595,N_18990,N_18504);
and U20596 (N_20596,N_17816,N_19523);
nor U20597 (N_20597,N_18318,N_18320);
or U20598 (N_20598,N_18832,N_17705);
or U20599 (N_20599,N_18678,N_17698);
xor U20600 (N_20600,N_17788,N_19304);
xor U20601 (N_20601,N_19971,N_18761);
or U20602 (N_20602,N_18078,N_18913);
or U20603 (N_20603,N_17789,N_18477);
nand U20604 (N_20604,N_18329,N_19628);
nor U20605 (N_20605,N_18369,N_18189);
nand U20606 (N_20606,N_19323,N_18347);
or U20607 (N_20607,N_18723,N_18579);
nor U20608 (N_20608,N_19352,N_18975);
xnor U20609 (N_20609,N_17809,N_18440);
or U20610 (N_20610,N_17592,N_19318);
or U20611 (N_20611,N_19880,N_18517);
and U20612 (N_20612,N_17945,N_17933);
nand U20613 (N_20613,N_19207,N_19744);
nor U20614 (N_20614,N_19309,N_19877);
nand U20615 (N_20615,N_18670,N_19305);
nor U20616 (N_20616,N_19348,N_17746);
nor U20617 (N_20617,N_19067,N_19941);
nand U20618 (N_20618,N_18025,N_18966);
or U20619 (N_20619,N_18771,N_17764);
nor U20620 (N_20620,N_19341,N_19917);
xnor U20621 (N_20621,N_19294,N_18175);
or U20622 (N_20622,N_18208,N_17757);
nor U20623 (N_20623,N_18459,N_18167);
and U20624 (N_20624,N_19522,N_18103);
xnor U20625 (N_20625,N_17677,N_19464);
or U20626 (N_20626,N_19773,N_17688);
xnor U20627 (N_20627,N_18720,N_18030);
nor U20628 (N_20628,N_18824,N_19691);
xnor U20629 (N_20629,N_17915,N_17532);
nor U20630 (N_20630,N_19453,N_18515);
nor U20631 (N_20631,N_18247,N_18054);
nand U20632 (N_20632,N_17708,N_19796);
nand U20633 (N_20633,N_17876,N_19991);
xnor U20634 (N_20634,N_18759,N_19899);
xor U20635 (N_20635,N_18948,N_19182);
or U20636 (N_20636,N_18421,N_17559);
or U20637 (N_20637,N_18584,N_17852);
nor U20638 (N_20638,N_17661,N_19282);
nand U20639 (N_20639,N_17604,N_18126);
nand U20640 (N_20640,N_18447,N_19394);
and U20641 (N_20641,N_18168,N_19421);
nand U20642 (N_20642,N_18422,N_18265);
nand U20643 (N_20643,N_19972,N_18197);
nor U20644 (N_20644,N_17749,N_18545);
or U20645 (N_20645,N_17612,N_17939);
nor U20646 (N_20646,N_18634,N_18233);
nor U20647 (N_20647,N_19818,N_18015);
xor U20648 (N_20648,N_18325,N_19587);
and U20649 (N_20649,N_17946,N_18648);
xor U20650 (N_20650,N_19937,N_19365);
or U20651 (N_20651,N_19400,N_18728);
nand U20652 (N_20652,N_17526,N_18967);
nor U20653 (N_20653,N_19407,N_18750);
nand U20654 (N_20654,N_17514,N_18372);
nand U20655 (N_20655,N_18596,N_17822);
nor U20656 (N_20656,N_18917,N_18493);
and U20657 (N_20657,N_18993,N_17725);
nor U20658 (N_20658,N_18009,N_18565);
nand U20659 (N_20659,N_18629,N_17784);
or U20660 (N_20660,N_18937,N_19007);
xnor U20661 (N_20661,N_19009,N_19096);
nor U20662 (N_20662,N_18547,N_19397);
nor U20663 (N_20663,N_18261,N_19958);
nand U20664 (N_20664,N_17996,N_19583);
and U20665 (N_20665,N_18140,N_17850);
or U20666 (N_20666,N_19986,N_19314);
nand U20667 (N_20667,N_18525,N_19614);
nor U20668 (N_20668,N_17702,N_19582);
xor U20669 (N_20669,N_18462,N_18881);
or U20670 (N_20670,N_19952,N_19022);
nand U20671 (N_20671,N_17599,N_18298);
xnor U20672 (N_20672,N_17618,N_19345);
nand U20673 (N_20673,N_19576,N_19060);
and U20674 (N_20674,N_18836,N_19477);
nand U20675 (N_20675,N_18603,N_19869);
nand U20676 (N_20676,N_19058,N_19798);
nand U20677 (N_20677,N_19147,N_17968);
or U20678 (N_20678,N_19032,N_18695);
and U20679 (N_20679,N_19743,N_19250);
and U20680 (N_20680,N_18907,N_19779);
nand U20681 (N_20681,N_18436,N_19724);
nand U20682 (N_20682,N_19968,N_18432);
xor U20683 (N_20683,N_19820,N_19013);
nand U20684 (N_20684,N_18442,N_17724);
or U20685 (N_20685,N_18062,N_17537);
nand U20686 (N_20686,N_18370,N_19728);
nand U20687 (N_20687,N_19596,N_18540);
nor U20688 (N_20688,N_19073,N_18575);
nand U20689 (N_20689,N_18594,N_19422);
and U20690 (N_20690,N_19074,N_17564);
nand U20691 (N_20691,N_18834,N_18950);
or U20692 (N_20692,N_19492,N_18479);
nand U20693 (N_20693,N_18521,N_17665);
nor U20694 (N_20694,N_19931,N_18972);
or U20695 (N_20695,N_18150,N_19035);
xnor U20696 (N_20696,N_17902,N_19572);
or U20697 (N_20697,N_17774,N_17577);
and U20698 (N_20698,N_19656,N_18463);
nor U20699 (N_20699,N_19992,N_18607);
and U20700 (N_20700,N_18214,N_19967);
nor U20701 (N_20701,N_17810,N_18155);
or U20702 (N_20702,N_19755,N_19385);
nand U20703 (N_20703,N_17507,N_17826);
nand U20704 (N_20704,N_18378,N_19645);
nor U20705 (N_20705,N_18791,N_18256);
nor U20706 (N_20706,N_19934,N_18511);
nor U20707 (N_20707,N_18397,N_18979);
xor U20708 (N_20708,N_17546,N_17813);
and U20709 (N_20709,N_19148,N_19239);
xor U20710 (N_20710,N_19787,N_18398);
nand U20711 (N_20711,N_17953,N_17838);
or U20712 (N_20712,N_19521,N_17595);
nand U20713 (N_20713,N_18800,N_19292);
nand U20714 (N_20714,N_19039,N_17761);
and U20715 (N_20715,N_18546,N_19736);
nor U20716 (N_20716,N_17909,N_17660);
nand U20717 (N_20717,N_19303,N_19098);
xor U20718 (N_20718,N_18935,N_19356);
and U20719 (N_20719,N_19819,N_18131);
xor U20720 (N_20720,N_18158,N_18769);
or U20721 (N_20721,N_18049,N_19011);
xor U20722 (N_20722,N_19651,N_19269);
nand U20723 (N_20723,N_18745,N_19641);
nand U20724 (N_20724,N_19440,N_19667);
or U20725 (N_20725,N_19086,N_18994);
and U20726 (N_20726,N_18157,N_19982);
or U20727 (N_20727,N_19690,N_18897);
nor U20728 (N_20728,N_19854,N_18450);
xor U20729 (N_20729,N_17934,N_17841);
nand U20730 (N_20730,N_19979,N_19805);
or U20731 (N_20731,N_17606,N_18998);
nor U20732 (N_20732,N_18616,N_18690);
or U20733 (N_20733,N_18642,N_19112);
nor U20734 (N_20734,N_18355,N_19398);
or U20735 (N_20735,N_19843,N_17581);
nor U20736 (N_20736,N_17879,N_19493);
or U20737 (N_20737,N_19478,N_18232);
xor U20738 (N_20738,N_17587,N_17821);
nor U20739 (N_20739,N_18020,N_18352);
nor U20740 (N_20740,N_19558,N_19487);
xnor U20741 (N_20741,N_17802,N_18299);
or U20742 (N_20742,N_18884,N_17547);
nor U20743 (N_20743,N_18639,N_19757);
xor U20744 (N_20744,N_19946,N_19748);
nor U20745 (N_20745,N_18153,N_19328);
and U20746 (N_20746,N_18730,N_19781);
nand U20747 (N_20747,N_19042,N_17540);
nand U20748 (N_20748,N_18102,N_17634);
or U20749 (N_20749,N_19512,N_19615);
nand U20750 (N_20750,N_19484,N_18893);
nor U20751 (N_20751,N_17859,N_18411);
nor U20752 (N_20752,N_19716,N_18736);
nand U20753 (N_20753,N_18781,N_19602);
nand U20754 (N_20754,N_18201,N_19193);
xor U20755 (N_20755,N_19685,N_19903);
and U20756 (N_20756,N_19756,N_19944);
xor U20757 (N_20757,N_18663,N_19053);
xnor U20758 (N_20758,N_19893,N_17711);
nor U20759 (N_20759,N_17712,N_18704);
and U20760 (N_20760,N_19006,N_19978);
nor U20761 (N_20761,N_18583,N_17734);
and U20762 (N_20762,N_19987,N_19738);
and U20763 (N_20763,N_19364,N_19555);
nor U20764 (N_20764,N_19384,N_19295);
nor U20765 (N_20765,N_19313,N_18393);
or U20766 (N_20766,N_18154,N_18353);
nand U20767 (N_20767,N_18826,N_18222);
or U20768 (N_20768,N_18236,N_19761);
and U20769 (N_20769,N_17950,N_18405);
and U20770 (N_20770,N_19065,N_18845);
nor U20771 (N_20771,N_17543,N_18986);
nor U20772 (N_20772,N_19410,N_19688);
nor U20773 (N_20773,N_17973,N_18630);
nand U20774 (N_20774,N_19476,N_19454);
and U20775 (N_20775,N_18003,N_17962);
or U20776 (N_20776,N_18637,N_17583);
and U20777 (N_20777,N_19222,N_19769);
nor U20778 (N_20778,N_18506,N_19940);
nand U20779 (N_20779,N_17720,N_19122);
nand U20780 (N_20780,N_17743,N_18099);
nor U20781 (N_20781,N_18074,N_19961);
nand U20782 (N_20782,N_17769,N_18181);
nand U20783 (N_20783,N_19888,N_18042);
or U20784 (N_20784,N_18744,N_18348);
xor U20785 (N_20785,N_18818,N_17798);
nand U20786 (N_20786,N_19056,N_17704);
nand U20787 (N_20787,N_17570,N_18467);
nand U20788 (N_20788,N_18709,N_19485);
and U20789 (N_20789,N_18040,N_19680);
and U20790 (N_20790,N_19256,N_19565);
and U20791 (N_20791,N_18027,N_19431);
nor U20792 (N_20792,N_17539,N_19346);
or U20793 (N_20793,N_19567,N_18860);
nand U20794 (N_20794,N_18706,N_19840);
and U20795 (N_20795,N_19622,N_18719);
xor U20796 (N_20796,N_19177,N_18281);
or U20797 (N_20797,N_19066,N_19127);
and U20798 (N_20798,N_18809,N_19474);
or U20799 (N_20799,N_18729,N_18711);
or U20800 (N_20800,N_17756,N_19158);
nand U20801 (N_20801,N_19167,N_19705);
xor U20802 (N_20802,N_18940,N_19029);
nand U20803 (N_20803,N_19947,N_18494);
xor U20804 (N_20804,N_19369,N_18676);
nor U20805 (N_20805,N_19120,N_17820);
nor U20806 (N_20806,N_18799,N_18340);
nor U20807 (N_20807,N_18560,N_19579);
xnor U20808 (N_20808,N_19762,N_19235);
xor U20809 (N_20809,N_19375,N_18714);
nor U20810 (N_20810,N_19780,N_19183);
or U20811 (N_20811,N_19273,N_18343);
nand U20812 (N_20812,N_18636,N_19948);
nor U20813 (N_20813,N_18045,N_18962);
and U20814 (N_20814,N_19658,N_18474);
xnor U20815 (N_20815,N_18453,N_19799);
nor U20816 (N_20816,N_19663,N_18067);
and U20817 (N_20817,N_18674,N_18968);
nor U20818 (N_20818,N_18481,N_18700);
and U20819 (N_20819,N_17961,N_17870);
xor U20820 (N_20820,N_18703,N_19726);
nor U20821 (N_20821,N_17518,N_17927);
nor U20822 (N_20822,N_19041,N_18855);
nand U20823 (N_20823,N_18668,N_18531);
and U20824 (N_20824,N_18605,N_17567);
or U20825 (N_20825,N_18039,N_18227);
xor U20826 (N_20826,N_18577,N_17872);
and U20827 (N_20827,N_18519,N_18149);
nand U20828 (N_20828,N_17770,N_18007);
nor U20829 (N_20829,N_17707,N_19500);
or U20830 (N_20830,N_19867,N_19938);
and U20831 (N_20831,N_17684,N_18409);
nand U20832 (N_20832,N_18527,N_19023);
nand U20833 (N_20833,N_17951,N_19775);
nand U20834 (N_20834,N_18625,N_18699);
xnor U20835 (N_20835,N_18796,N_17647);
or U20836 (N_20836,N_17696,N_17693);
nor U20837 (N_20837,N_19461,N_17913);
or U20838 (N_20838,N_19391,N_19354);
or U20839 (N_20839,N_17839,N_19126);
and U20840 (N_20840,N_19336,N_18376);
nand U20841 (N_20841,N_18114,N_19146);
xnor U20842 (N_20842,N_17525,N_17633);
xnor U20843 (N_20843,N_17818,N_17616);
xor U20844 (N_20844,N_18388,N_18011);
or U20845 (N_20845,N_18400,N_18057);
and U20846 (N_20846,N_19802,N_17780);
nor U20847 (N_20847,N_18351,N_17853);
nand U20848 (N_20848,N_19355,N_19428);
nor U20849 (N_20849,N_18293,N_18359);
nor U20850 (N_20850,N_18217,N_18441);
nand U20851 (N_20851,N_17626,N_18137);
or U20852 (N_20852,N_19218,N_18278);
xnor U20853 (N_20853,N_19672,N_19812);
and U20854 (N_20854,N_17615,N_18622);
or U20855 (N_20855,N_17926,N_19230);
and U20856 (N_20856,N_18877,N_18268);
nor U20857 (N_20857,N_19253,N_19750);
nand U20858 (N_20858,N_19537,N_19920);
xor U20859 (N_20859,N_17610,N_18053);
xnor U20860 (N_20860,N_18121,N_19139);
or U20861 (N_20861,N_19499,N_19382);
nand U20862 (N_20862,N_19886,N_19450);
nor U20863 (N_20863,N_17793,N_18953);
nand U20864 (N_20864,N_18802,N_18315);
nor U20865 (N_20865,N_19720,N_17997);
nand U20866 (N_20866,N_19752,N_17830);
nand U20867 (N_20867,N_18475,N_18518);
nor U20868 (N_20868,N_18346,N_18386);
xnor U20869 (N_20869,N_18739,N_18532);
or U20870 (N_20870,N_18023,N_17795);
xor U20871 (N_20871,N_18892,N_19528);
nand U20872 (N_20872,N_18044,N_19841);
nand U20873 (N_20873,N_18143,N_17866);
xnor U20874 (N_20874,N_19020,N_17956);
nand U20875 (N_20875,N_18332,N_19301);
nor U20876 (N_20876,N_19679,N_18434);
and U20877 (N_20877,N_17639,N_18136);
and U20878 (N_20878,N_18283,N_18470);
nor U20879 (N_20879,N_17736,N_18185);
nor U20880 (N_20880,N_18666,N_18334);
xor U20881 (N_20881,N_17758,N_18890);
and U20882 (N_20882,N_18794,N_18687);
nand U20883 (N_20883,N_19479,N_19288);
and U20884 (N_20884,N_19676,N_17569);
or U20885 (N_20885,N_19466,N_18286);
xor U20886 (N_20886,N_19751,N_18904);
nand U20887 (N_20887,N_19161,N_18305);
nor U20888 (N_20888,N_18974,N_18537);
or U20889 (N_20889,N_17641,N_19082);
and U20890 (N_20890,N_18373,N_18430);
nand U20891 (N_20891,N_17837,N_18710);
xor U20892 (N_20892,N_18019,N_19556);
or U20893 (N_20893,N_19271,N_18427);
and U20894 (N_20894,N_17955,N_19362);
or U20895 (N_20895,N_18259,N_19507);
or U20896 (N_20896,N_18145,N_19564);
xnor U20897 (N_20897,N_19076,N_19442);
or U20898 (N_20898,N_18361,N_17651);
or U20899 (N_20899,N_19244,N_17680);
and U20900 (N_20900,N_18612,N_17671);
or U20901 (N_20901,N_18838,N_19610);
nor U20902 (N_20902,N_18901,N_19031);
xnor U20903 (N_20903,N_19229,N_19918);
nor U20904 (N_20904,N_19549,N_19866);
and U20905 (N_20905,N_19327,N_19010);
or U20906 (N_20906,N_18419,N_17834);
or U20907 (N_20907,N_19495,N_18316);
xnor U20908 (N_20908,N_19378,N_19317);
and U20909 (N_20909,N_18176,N_19589);
nor U20910 (N_20910,N_18097,N_18234);
nor U20911 (N_20911,N_18106,N_19134);
nor U20912 (N_20912,N_18413,N_17755);
nor U20913 (N_20913,N_19925,N_19878);
nand U20914 (N_20914,N_18726,N_18599);
xor U20915 (N_20915,N_19180,N_19359);
nor U20916 (N_20916,N_19160,N_18541);
nand U20917 (N_20917,N_18250,N_17653);
and U20918 (N_20918,N_17971,N_17682);
nor U20919 (N_20919,N_19533,N_19432);
nand U20920 (N_20920,N_19221,N_17970);
or U20921 (N_20921,N_19783,N_19696);
xnor U20922 (N_20922,N_19335,N_18251);
nor U20923 (N_20923,N_19427,N_19848);
and U20924 (N_20924,N_18872,N_17804);
or U20925 (N_20925,N_18553,N_18466);
xor U20926 (N_20926,N_17691,N_19885);
and U20927 (N_20927,N_18092,N_19776);
xnor U20928 (N_20928,N_19224,N_18303);
nor U20929 (N_20929,N_18169,N_19373);
nand U20930 (N_20930,N_19460,N_19553);
xnor U20931 (N_20931,N_17738,N_19777);
xnor U20932 (N_20932,N_18920,N_19559);
nor U20933 (N_20933,N_18960,N_18691);
or U20934 (N_20934,N_18671,N_19497);
nor U20935 (N_20935,N_18991,N_19131);
nand U20936 (N_20936,N_18014,N_18965);
nand U20937 (N_20937,N_17782,N_19210);
or U20938 (N_20938,N_19241,N_18199);
nand U20939 (N_20939,N_18367,N_17689);
nand U20940 (N_20940,N_17553,N_18076);
xor U20941 (N_20941,N_17885,N_19452);
xor U20942 (N_20942,N_18402,N_19153);
and U20943 (N_20943,N_18598,N_18863);
nand U20944 (N_20944,N_18120,N_18301);
nand U20945 (N_20945,N_17888,N_18589);
and U20946 (N_20946,N_19051,N_19990);
xor U20947 (N_20947,N_19504,N_17916);
and U20948 (N_20948,N_19926,N_19257);
xor U20949 (N_20949,N_19874,N_18489);
and U20950 (N_20950,N_18602,N_19700);
xnor U20951 (N_20951,N_19539,N_18554);
xor U20952 (N_20952,N_18805,N_19906);
nand U20953 (N_20953,N_19502,N_18193);
xnor U20954 (N_20954,N_17718,N_19689);
nor U20955 (N_20955,N_18262,N_19631);
nor U20956 (N_20956,N_19283,N_18919);
and U20957 (N_20957,N_18198,N_17865);
nor U20958 (N_20958,N_19409,N_19860);
nand U20959 (N_20959,N_19034,N_19293);
and U20960 (N_20960,N_18874,N_19546);
xor U20961 (N_20961,N_19711,N_17848);
xor U20962 (N_20962,N_19910,N_18776);
nand U20963 (N_20963,N_18423,N_19730);
xnor U20964 (N_20964,N_17846,N_19890);
nand U20965 (N_20965,N_18697,N_18694);
or U20966 (N_20966,N_19525,N_18204);
or U20967 (N_20967,N_18324,N_19265);
nor U20968 (N_20968,N_18173,N_17944);
or U20969 (N_20969,N_17751,N_18132);
and U20970 (N_20970,N_19434,N_19643);
xor U20971 (N_20971,N_19809,N_19739);
and U20972 (N_20972,N_18404,N_19107);
and U20973 (N_20973,N_17602,N_19080);
or U20974 (N_20974,N_19014,N_18752);
nor U20975 (N_20975,N_19793,N_18041);
nand U20976 (N_20976,N_19480,N_19570);
nor U20977 (N_20977,N_18387,N_17745);
or U20978 (N_20978,N_18113,N_19668);
nor U20979 (N_20979,N_18669,N_18733);
and U20980 (N_20980,N_17799,N_17703);
nand U20981 (N_20981,N_19935,N_18693);
xor U20982 (N_20982,N_18172,N_17591);
and U20983 (N_20983,N_19800,N_18322);
and U20984 (N_20984,N_19408,N_17594);
nand U20985 (N_20985,N_19600,N_19795);
xor U20986 (N_20986,N_17790,N_17847);
nor U20987 (N_20987,N_17692,N_17805);
xor U20988 (N_20988,N_18916,N_19547);
xnor U20989 (N_20989,N_19638,N_18997);
and U20990 (N_20990,N_19315,N_19374);
xor U20991 (N_20991,N_19413,N_19297);
and U20992 (N_20992,N_19881,N_19545);
or U20993 (N_20993,N_18611,N_18269);
nand U20994 (N_20994,N_18245,N_18371);
nand U20995 (N_20995,N_17571,N_18223);
or U20996 (N_20996,N_18508,N_18342);
and U20997 (N_20997,N_17912,N_19823);
or U20998 (N_20998,N_19114,N_18559);
xnor U20999 (N_20999,N_17541,N_18797);
xor U21000 (N_21000,N_17776,N_19807);
and U21001 (N_21001,N_17555,N_18708);
nand U21002 (N_21002,N_18207,N_19955);
xor U21003 (N_21003,N_18284,N_18424);
nand U21004 (N_21004,N_18160,N_18644);
and U21005 (N_21005,N_19772,N_19715);
nand U21006 (N_21006,N_18192,N_18206);
and U21007 (N_21007,N_18581,N_17624);
nor U21008 (N_21008,N_19001,N_19939);
nor U21009 (N_21009,N_18984,N_17762);
nand U21010 (N_21010,N_19949,N_18909);
or U21011 (N_21011,N_17674,N_19640);
nand U21012 (N_21012,N_18456,N_18908);
and U21013 (N_21013,N_19865,N_19319);
and U21014 (N_21014,N_19030,N_19902);
or U21015 (N_21015,N_18182,N_19083);
and U21016 (N_21016,N_19904,N_18885);
and U21017 (N_21017,N_17742,N_17588);
nand U21018 (N_21018,N_19178,N_18483);
and U21019 (N_21019,N_18321,N_18392);
xor U21020 (N_21020,N_17932,N_19846);
or U21021 (N_21021,N_18110,N_17744);
and U21022 (N_21022,N_19330,N_18486);
xor U21023 (N_21023,N_17998,N_17557);
and U21024 (N_21024,N_19763,N_18488);
xnor U21025 (N_21025,N_17520,N_19088);
or U21026 (N_21026,N_18613,N_19963);
and U21027 (N_21027,N_17963,N_19782);
or U21028 (N_21028,N_18151,N_18562);
nand U21029 (N_21029,N_19962,N_18035);
nor U21030 (N_21030,N_19683,N_18804);
nor U21031 (N_21031,N_19976,N_18366);
xnor U21032 (N_21032,N_19532,N_17727);
nand U21033 (N_21033,N_17729,N_18141);
or U21034 (N_21034,N_19470,N_19005);
nand U21035 (N_21035,N_17930,N_19115);
nor U21036 (N_21036,N_18939,N_18889);
xor U21037 (N_21037,N_17575,N_17923);
nor U21038 (N_21038,N_17981,N_17921);
nand U21039 (N_21039,N_19353,N_19791);
xor U21040 (N_21040,N_18480,N_18767);
or U21041 (N_21041,N_17658,N_19542);
nor U21042 (N_21042,N_18148,N_18358);
nor U21043 (N_21043,N_19876,N_19025);
xor U21044 (N_21044,N_17843,N_19486);
xor U21045 (N_21045,N_19376,N_18593);
nor U21046 (N_21046,N_19811,N_19753);
nor U21047 (N_21047,N_18108,N_18374);
xnor U21048 (N_21048,N_17893,N_17922);
nand U21049 (N_21049,N_19562,N_17767);
nand U21050 (N_21050,N_19684,N_18770);
and U21051 (N_21051,N_17637,N_17545);
xor U21052 (N_21052,N_18783,N_19644);
and U21053 (N_21053,N_19804,N_18524);
or U21054 (N_21054,N_18431,N_18779);
nand U21055 (N_21055,N_18534,N_18929);
nor U21056 (N_21056,N_17611,N_17586);
nand U21057 (N_21057,N_18696,N_19040);
xor U21058 (N_21058,N_18858,N_17701);
nor U21059 (N_21059,N_18224,N_18095);
nor U21060 (N_21060,N_17524,N_17977);
or U21061 (N_21061,N_19246,N_18864);
xor U21062 (N_21062,N_19778,N_18886);
nand U21063 (N_21063,N_19279,N_19162);
nor U21064 (N_21064,N_18004,N_18252);
or U21065 (N_21065,N_18510,N_19574);
nand U21066 (N_21066,N_17791,N_19919);
xor U21067 (N_21067,N_18764,N_18837);
and U21068 (N_21068,N_19599,N_19334);
and U21069 (N_21069,N_18026,N_17869);
xor U21070 (N_21070,N_18013,N_17656);
nor U21071 (N_21071,N_19285,N_17935);
nor U21072 (N_21072,N_17900,N_19758);
or U21073 (N_21073,N_18930,N_17887);
xor U21074 (N_21074,N_17572,N_19729);
or U21075 (N_21075,N_19655,N_19731);
xnor U21076 (N_21076,N_19372,N_19052);
and U21077 (N_21077,N_18338,N_19197);
nand U21078 (N_21078,N_19970,N_18310);
nand U21079 (N_21079,N_18814,N_19611);
nand U21080 (N_21080,N_19792,N_17601);
nand U21081 (N_21081,N_19932,N_18512);
xnor U21082 (N_21082,N_18539,N_19580);
or U21083 (N_21083,N_17613,N_19725);
and U21084 (N_21084,N_19965,N_17903);
or U21085 (N_21085,N_18774,N_18829);
xor U21086 (N_21086,N_17873,N_18552);
xnor U21087 (N_21087,N_18200,N_18280);
and U21088 (N_21088,N_19416,N_17918);
and U21089 (N_21089,N_18473,N_17621);
nand U21090 (N_21090,N_19324,N_17993);
nand U21091 (N_21091,N_17675,N_18130);
nand U21092 (N_21092,N_17509,N_19277);
nand U21093 (N_21093,N_17814,N_18446);
xor U21094 (N_21094,N_17659,N_18046);
nor U21095 (N_21095,N_19424,N_18061);
xor U21096 (N_21096,N_19310,N_19308);
and U21097 (N_21097,N_19357,N_18535);
or U21098 (N_21098,N_18681,N_19261);
or U21099 (N_21099,N_19816,N_19388);
and U21100 (N_21100,N_19490,N_19695);
nor U21101 (N_21101,N_18667,N_17864);
and U21102 (N_21102,N_18487,N_19347);
nand U21103 (N_21103,N_18712,N_18503);
and U21104 (N_21104,N_18619,N_19226);
nand U21105 (N_21105,N_17542,N_17508);
nand U21106 (N_21106,N_19448,N_19186);
nor U21107 (N_21107,N_18880,N_18576);
or U21108 (N_21108,N_19483,N_18377);
and U21109 (N_21109,N_18412,N_18716);
and U21110 (N_21110,N_18072,N_18762);
and U21111 (N_21111,N_19468,N_18949);
nand U21112 (N_21112,N_19211,N_19660);
xnor U21113 (N_21113,N_17765,N_18091);
xor U21114 (N_21114,N_18418,N_19092);
nor U21115 (N_21115,N_19682,N_18801);
nand U21116 (N_21116,N_18356,N_19417);
nand U21117 (N_21117,N_19872,N_19102);
or U21118 (N_21118,N_17990,N_19635);
or U21119 (N_21119,N_17806,N_17978);
and U21120 (N_21120,N_18165,N_18938);
and U21121 (N_21121,N_17735,N_17994);
or U21122 (N_21122,N_18942,N_18073);
nor U21123 (N_21123,N_18087,N_17901);
and U21124 (N_21124,N_19535,N_19966);
nand U21125 (N_21125,N_18461,N_18129);
nand U21126 (N_21126,N_19078,N_18934);
xor U21127 (N_21127,N_17785,N_17632);
or U21128 (N_21128,N_19420,N_18526);
nand U21129 (N_21129,N_18312,N_18349);
nand U21130 (N_21130,N_18787,N_18101);
or U21131 (N_21131,N_19629,N_17786);
and U21132 (N_21132,N_19871,N_19648);
nand U21133 (N_21133,N_19896,N_19403);
xor U21134 (N_21134,N_18961,N_19859);
and U21135 (N_21135,N_19526,N_19109);
and U21136 (N_21136,N_18401,N_18156);
nor U21137 (N_21137,N_18969,N_18218);
nor U21138 (N_21138,N_19928,N_19168);
and U21139 (N_21139,N_19554,N_17531);
nor U21140 (N_21140,N_17989,N_18403);
and U21141 (N_21141,N_18823,N_18921);
nor U21142 (N_21142,N_18161,N_19591);
nor U21143 (N_21143,N_18174,N_17652);
xor U21144 (N_21144,N_19094,N_18416);
or U21145 (N_21145,N_18849,N_17694);
nor U21146 (N_21146,N_18079,N_19853);
and U21147 (N_21147,N_18954,N_18586);
and U21148 (N_21148,N_18647,N_17732);
or U21149 (N_21149,N_18396,N_19171);
or U21150 (N_21150,N_17527,N_19358);
or U21151 (N_21151,N_19419,N_17554);
and U21152 (N_21152,N_17561,N_18815);
nand U21153 (N_21153,N_18878,N_18410);
nand U21154 (N_21154,N_18089,N_18341);
xnor U21155 (N_21155,N_18627,N_18282);
or U21156 (N_21156,N_17730,N_18951);
and U21157 (N_21157,N_19234,N_19363);
nor U21158 (N_21158,N_19412,N_19710);
or U21159 (N_21159,N_17874,N_18660);
nor U21160 (N_21160,N_18817,N_19789);
nor U21161 (N_21161,N_18417,N_19036);
xnor U21162 (N_21162,N_18266,N_19719);
or U21163 (N_21163,N_17714,N_19349);
or U21164 (N_21164,N_18038,N_18017);
nand U21165 (N_21165,N_18008,N_18989);
and U21166 (N_21166,N_19784,N_18476);
xnor U21167 (N_21167,N_17992,N_18841);
and U21168 (N_21168,N_19090,N_17904);
or U21169 (N_21169,N_18922,N_18068);
nand U21170 (N_21170,N_19225,N_18992);
nor U21171 (N_21171,N_17623,N_17863);
nor U21172 (N_21172,N_18081,N_19232);
xnor U21173 (N_21173,N_18777,N_18601);
nor U21174 (N_21174,N_17619,N_18327);
or U21175 (N_21175,N_18588,N_18980);
or U21176 (N_21176,N_17670,N_18782);
or U21177 (N_21177,N_18449,N_18580);
and U21178 (N_21178,N_18900,N_19219);
xnor U21179 (N_21179,N_19864,N_18882);
and U21180 (N_21180,N_19249,N_18820);
and U21181 (N_21181,N_18848,N_17598);
and U21182 (N_21182,N_18879,N_18812);
and U21183 (N_21183,N_17983,N_19983);
nor U21184 (N_21184,N_17833,N_19924);
xor U21185 (N_21185,N_18609,N_19844);
and U21186 (N_21186,N_18118,N_18773);
nand U21187 (N_21187,N_18024,N_19037);
nand U21188 (N_21188,N_19456,N_18737);
nor U21189 (N_21189,N_17988,N_17678);
and U21190 (N_21190,N_19209,N_17937);
or U21191 (N_21191,N_17875,N_19033);
or U21192 (N_21192,N_19404,N_19954);
nor U21193 (N_21193,N_17920,N_19957);
and U21194 (N_21194,N_17868,N_19175);
xnor U21195 (N_21195,N_17829,N_19834);
xor U21196 (N_21196,N_19061,N_17528);
or U21197 (N_21197,N_17669,N_17500);
or U21198 (N_21198,N_18566,N_17797);
nor U21199 (N_21199,N_18146,N_19491);
nand U21200 (N_21200,N_18362,N_18394);
xnor U21201 (N_21201,N_17709,N_19870);
nor U21202 (N_21202,N_18999,N_19810);
nor U21203 (N_21203,N_19264,N_18107);
xnor U21204 (N_21204,N_18533,N_19028);
and U21205 (N_21205,N_18740,N_17644);
and U21206 (N_21206,N_18852,N_19268);
or U21207 (N_21207,N_19132,N_19145);
xnor U21208 (N_21208,N_18677,N_18784);
nand U21209 (N_21209,N_18060,N_17638);
xnor U21210 (N_21210,N_17907,N_19469);
xor U21211 (N_21211,N_18574,N_19124);
nand U21212 (N_21212,N_18786,N_19262);
or U21213 (N_21213,N_18835,N_18144);
and U21214 (N_21214,N_17965,N_19560);
xnor U21215 (N_21215,N_18075,N_18621);
and U21216 (N_21216,N_18755,N_19392);
or U21217 (N_21217,N_17667,N_19675);
xor U21218 (N_21218,N_18032,N_19606);
or U21219 (N_21219,N_19157,N_18116);
xnor U21220 (N_21220,N_19557,N_19790);
and U21221 (N_21221,N_18724,N_18495);
xor U21222 (N_21222,N_18499,N_17858);
nand U21223 (N_21223,N_19097,N_19204);
xor U21224 (N_21224,N_19390,N_18721);
nand U21225 (N_21225,N_19527,N_17849);
nand U21226 (N_21226,N_19927,N_18375);
nand U21227 (N_21227,N_19956,N_17568);
nor U21228 (N_21228,N_17516,N_19653);
nand U21229 (N_21229,N_19855,N_18354);
nand U21230 (N_21230,N_18111,N_19343);
or U21231 (N_21231,N_18239,N_19108);
nand U21232 (N_21232,N_19383,N_18828);
nor U21233 (N_21233,N_19017,N_17836);
nand U21234 (N_21234,N_19260,N_17679);
or U21235 (N_21235,N_18230,N_18289);
nor U21236 (N_21236,N_17700,N_17860);
xor U21237 (N_21237,N_18831,N_19771);
and U21238 (N_21238,N_19659,N_19117);
and U21239 (N_21239,N_19740,N_17535);
nor U21240 (N_21240,N_17687,N_19650);
and U21241 (N_21241,N_18497,N_18059);
xor U21242 (N_21242,N_18433,N_18926);
nor U21243 (N_21243,N_17910,N_19923);
nor U21244 (N_21244,N_18337,N_18100);
nor U21245 (N_21245,N_19732,N_18955);
nor U21246 (N_21246,N_18868,N_18746);
nor U21247 (N_21247,N_19722,N_17657);
or U21248 (N_21248,N_19019,N_19459);
xnor U21249 (N_21249,N_18888,N_18368);
nand U21250 (N_21250,N_19236,N_19416);
nor U21251 (N_21251,N_19608,N_18350);
or U21252 (N_21252,N_19439,N_18073);
xnor U21253 (N_21253,N_18308,N_19211);
nor U21254 (N_21254,N_19734,N_19928);
xor U21255 (N_21255,N_19629,N_19476);
nor U21256 (N_21256,N_18013,N_18044);
nand U21257 (N_21257,N_19171,N_18667);
xnor U21258 (N_21258,N_17927,N_18285);
or U21259 (N_21259,N_18866,N_19579);
and U21260 (N_21260,N_18356,N_18235);
nand U21261 (N_21261,N_19649,N_17938);
nor U21262 (N_21262,N_18176,N_19471);
nand U21263 (N_21263,N_19870,N_18728);
nor U21264 (N_21264,N_19418,N_18796);
or U21265 (N_21265,N_19871,N_17852);
nor U21266 (N_21266,N_17634,N_18649);
nand U21267 (N_21267,N_17975,N_19313);
and U21268 (N_21268,N_19518,N_18207);
or U21269 (N_21269,N_17860,N_18959);
or U21270 (N_21270,N_17767,N_18165);
nor U21271 (N_21271,N_18562,N_19418);
nor U21272 (N_21272,N_18022,N_18188);
nor U21273 (N_21273,N_18973,N_19541);
xor U21274 (N_21274,N_19273,N_17951);
or U21275 (N_21275,N_19730,N_17973);
nand U21276 (N_21276,N_18442,N_19488);
and U21277 (N_21277,N_18108,N_18519);
nand U21278 (N_21278,N_18580,N_18722);
xnor U21279 (N_21279,N_17875,N_19722);
xor U21280 (N_21280,N_19447,N_18576);
or U21281 (N_21281,N_19969,N_18693);
nor U21282 (N_21282,N_18229,N_17807);
or U21283 (N_21283,N_17598,N_18421);
xor U21284 (N_21284,N_19815,N_17861);
nor U21285 (N_21285,N_19854,N_19270);
or U21286 (N_21286,N_17777,N_19370);
and U21287 (N_21287,N_19347,N_17657);
nor U21288 (N_21288,N_19239,N_18789);
and U21289 (N_21289,N_19385,N_19864);
xnor U21290 (N_21290,N_17795,N_18531);
nor U21291 (N_21291,N_18931,N_18459);
and U21292 (N_21292,N_19029,N_19419);
xor U21293 (N_21293,N_19297,N_17714);
or U21294 (N_21294,N_19663,N_18133);
nor U21295 (N_21295,N_18809,N_19803);
or U21296 (N_21296,N_17781,N_19325);
or U21297 (N_21297,N_18239,N_18866);
nand U21298 (N_21298,N_18238,N_19022);
xor U21299 (N_21299,N_17906,N_19882);
xnor U21300 (N_21300,N_17934,N_17908);
or U21301 (N_21301,N_19330,N_18788);
and U21302 (N_21302,N_17588,N_17959);
xor U21303 (N_21303,N_18383,N_19802);
nor U21304 (N_21304,N_17978,N_18007);
and U21305 (N_21305,N_17656,N_18118);
or U21306 (N_21306,N_18634,N_19638);
or U21307 (N_21307,N_18274,N_17721);
nand U21308 (N_21308,N_18884,N_18059);
xor U21309 (N_21309,N_18677,N_19632);
and U21310 (N_21310,N_18615,N_19458);
and U21311 (N_21311,N_18068,N_19879);
or U21312 (N_21312,N_18901,N_18154);
nor U21313 (N_21313,N_18862,N_17815);
nor U21314 (N_21314,N_19368,N_18215);
xor U21315 (N_21315,N_19116,N_18567);
or U21316 (N_21316,N_17766,N_19870);
xnor U21317 (N_21317,N_19113,N_19964);
nor U21318 (N_21318,N_19483,N_18252);
nand U21319 (N_21319,N_18535,N_18799);
and U21320 (N_21320,N_19423,N_18682);
and U21321 (N_21321,N_19976,N_17933);
or U21322 (N_21322,N_18590,N_18358);
nand U21323 (N_21323,N_18865,N_19447);
nand U21324 (N_21324,N_19640,N_17731);
and U21325 (N_21325,N_18055,N_18140);
xor U21326 (N_21326,N_18840,N_17655);
xor U21327 (N_21327,N_18302,N_19811);
nand U21328 (N_21328,N_17543,N_19177);
xnor U21329 (N_21329,N_18020,N_18535);
xor U21330 (N_21330,N_18792,N_19166);
and U21331 (N_21331,N_17550,N_19736);
nand U21332 (N_21332,N_17535,N_19664);
or U21333 (N_21333,N_18068,N_18351);
nor U21334 (N_21334,N_17787,N_18519);
or U21335 (N_21335,N_18659,N_18792);
or U21336 (N_21336,N_18576,N_19497);
xnor U21337 (N_21337,N_18972,N_19335);
nand U21338 (N_21338,N_19644,N_18085);
or U21339 (N_21339,N_19573,N_17700);
xnor U21340 (N_21340,N_18323,N_17750);
or U21341 (N_21341,N_18299,N_17934);
and U21342 (N_21342,N_19000,N_19741);
xnor U21343 (N_21343,N_19072,N_19411);
nand U21344 (N_21344,N_18902,N_19852);
nand U21345 (N_21345,N_17500,N_18134);
xnor U21346 (N_21346,N_18020,N_19194);
nor U21347 (N_21347,N_18549,N_19905);
xnor U21348 (N_21348,N_18031,N_19714);
xnor U21349 (N_21349,N_19465,N_18256);
and U21350 (N_21350,N_19648,N_19211);
and U21351 (N_21351,N_19357,N_17952);
nand U21352 (N_21352,N_18005,N_19132);
or U21353 (N_21353,N_19623,N_18673);
xor U21354 (N_21354,N_17775,N_18448);
xor U21355 (N_21355,N_19255,N_17700);
or U21356 (N_21356,N_19518,N_18504);
and U21357 (N_21357,N_18761,N_18590);
nand U21358 (N_21358,N_19846,N_18365);
and U21359 (N_21359,N_18574,N_19025);
and U21360 (N_21360,N_18872,N_19130);
nand U21361 (N_21361,N_18888,N_19524);
xor U21362 (N_21362,N_19376,N_18944);
nor U21363 (N_21363,N_19697,N_18700);
nor U21364 (N_21364,N_19491,N_18074);
or U21365 (N_21365,N_19484,N_18097);
or U21366 (N_21366,N_19670,N_17554);
and U21367 (N_21367,N_19626,N_18851);
nor U21368 (N_21368,N_18196,N_18505);
and U21369 (N_21369,N_19381,N_17573);
nor U21370 (N_21370,N_18831,N_19546);
xnor U21371 (N_21371,N_18903,N_18797);
and U21372 (N_21372,N_18228,N_17548);
nor U21373 (N_21373,N_18936,N_19096);
and U21374 (N_21374,N_18457,N_17900);
or U21375 (N_21375,N_18995,N_18042);
nand U21376 (N_21376,N_18445,N_19073);
xnor U21377 (N_21377,N_19465,N_19968);
and U21378 (N_21378,N_17699,N_19355);
nor U21379 (N_21379,N_17727,N_18248);
or U21380 (N_21380,N_17821,N_18683);
nor U21381 (N_21381,N_17885,N_19585);
xor U21382 (N_21382,N_18857,N_18241);
nor U21383 (N_21383,N_19996,N_18608);
or U21384 (N_21384,N_19646,N_17866);
or U21385 (N_21385,N_19270,N_19992);
or U21386 (N_21386,N_17913,N_19043);
nand U21387 (N_21387,N_19340,N_18244);
nand U21388 (N_21388,N_18822,N_17825);
nor U21389 (N_21389,N_17774,N_18221);
xor U21390 (N_21390,N_17886,N_19819);
xor U21391 (N_21391,N_19267,N_18446);
or U21392 (N_21392,N_19303,N_18618);
nand U21393 (N_21393,N_18105,N_18026);
xor U21394 (N_21394,N_19380,N_17517);
and U21395 (N_21395,N_17726,N_18789);
nor U21396 (N_21396,N_18264,N_19871);
nor U21397 (N_21397,N_18452,N_18252);
nand U21398 (N_21398,N_19170,N_17812);
xor U21399 (N_21399,N_19746,N_19314);
and U21400 (N_21400,N_17568,N_18400);
and U21401 (N_21401,N_19660,N_19461);
nor U21402 (N_21402,N_18046,N_18365);
nor U21403 (N_21403,N_18665,N_17534);
or U21404 (N_21404,N_18599,N_19379);
or U21405 (N_21405,N_18684,N_19539);
nand U21406 (N_21406,N_19437,N_19293);
nor U21407 (N_21407,N_18386,N_18476);
and U21408 (N_21408,N_18533,N_18558);
and U21409 (N_21409,N_17739,N_17982);
and U21410 (N_21410,N_18687,N_17924);
nor U21411 (N_21411,N_18313,N_19442);
xnor U21412 (N_21412,N_19605,N_19064);
xor U21413 (N_21413,N_19719,N_19430);
or U21414 (N_21414,N_18320,N_18956);
or U21415 (N_21415,N_18367,N_18682);
and U21416 (N_21416,N_18197,N_18373);
or U21417 (N_21417,N_19563,N_18980);
nor U21418 (N_21418,N_19630,N_17997);
xnor U21419 (N_21419,N_19302,N_18062);
nor U21420 (N_21420,N_18164,N_19883);
or U21421 (N_21421,N_19840,N_18802);
and U21422 (N_21422,N_18746,N_19933);
nand U21423 (N_21423,N_18226,N_18277);
xnor U21424 (N_21424,N_18103,N_19056);
nand U21425 (N_21425,N_19762,N_18679);
xor U21426 (N_21426,N_17592,N_18370);
xor U21427 (N_21427,N_18385,N_18778);
and U21428 (N_21428,N_19081,N_17615);
nand U21429 (N_21429,N_18656,N_18306);
nand U21430 (N_21430,N_18167,N_18143);
xor U21431 (N_21431,N_18479,N_17964);
xor U21432 (N_21432,N_18736,N_17807);
or U21433 (N_21433,N_19255,N_19272);
nor U21434 (N_21434,N_18997,N_18881);
xnor U21435 (N_21435,N_17580,N_18240);
or U21436 (N_21436,N_18987,N_19763);
xnor U21437 (N_21437,N_18352,N_18076);
nor U21438 (N_21438,N_17737,N_17892);
or U21439 (N_21439,N_18694,N_19545);
nor U21440 (N_21440,N_18561,N_19113);
xnor U21441 (N_21441,N_19812,N_19304);
nand U21442 (N_21442,N_19130,N_19851);
or U21443 (N_21443,N_17682,N_19404);
and U21444 (N_21444,N_19842,N_18197);
xor U21445 (N_21445,N_18883,N_17956);
nor U21446 (N_21446,N_19935,N_19395);
and U21447 (N_21447,N_18397,N_17797);
or U21448 (N_21448,N_19514,N_19717);
xnor U21449 (N_21449,N_17697,N_18121);
or U21450 (N_21450,N_18238,N_19794);
and U21451 (N_21451,N_19469,N_18138);
and U21452 (N_21452,N_17692,N_19750);
and U21453 (N_21453,N_19317,N_18992);
nand U21454 (N_21454,N_18857,N_18503);
or U21455 (N_21455,N_18822,N_17557);
and U21456 (N_21456,N_19539,N_18665);
and U21457 (N_21457,N_18940,N_18935);
nor U21458 (N_21458,N_17626,N_19027);
and U21459 (N_21459,N_19357,N_18432);
xnor U21460 (N_21460,N_18265,N_18685);
nand U21461 (N_21461,N_19825,N_19372);
xor U21462 (N_21462,N_18557,N_18033);
nand U21463 (N_21463,N_18385,N_18254);
nor U21464 (N_21464,N_19506,N_18065);
and U21465 (N_21465,N_19132,N_17506);
or U21466 (N_21466,N_18844,N_18047);
nor U21467 (N_21467,N_19338,N_19880);
nor U21468 (N_21468,N_17850,N_19806);
nor U21469 (N_21469,N_17883,N_17905);
or U21470 (N_21470,N_19553,N_19578);
xnor U21471 (N_21471,N_19869,N_18937);
or U21472 (N_21472,N_17779,N_17504);
or U21473 (N_21473,N_17791,N_19565);
or U21474 (N_21474,N_19495,N_17629);
nand U21475 (N_21475,N_18027,N_19695);
or U21476 (N_21476,N_19434,N_19244);
xnor U21477 (N_21477,N_18828,N_18597);
and U21478 (N_21478,N_17995,N_18173);
xnor U21479 (N_21479,N_18250,N_18100);
xor U21480 (N_21480,N_17971,N_17543);
or U21481 (N_21481,N_18628,N_18445);
or U21482 (N_21482,N_17884,N_18262);
xnor U21483 (N_21483,N_19009,N_19782);
nand U21484 (N_21484,N_19303,N_17578);
nand U21485 (N_21485,N_17939,N_19445);
nor U21486 (N_21486,N_19701,N_18236);
nand U21487 (N_21487,N_19640,N_17708);
xnor U21488 (N_21488,N_19831,N_17587);
and U21489 (N_21489,N_19598,N_19654);
nand U21490 (N_21490,N_18712,N_17509);
nand U21491 (N_21491,N_19566,N_18970);
xor U21492 (N_21492,N_17704,N_17624);
xor U21493 (N_21493,N_19616,N_17723);
nor U21494 (N_21494,N_18405,N_19469);
nand U21495 (N_21495,N_19569,N_19950);
nor U21496 (N_21496,N_19385,N_19338);
or U21497 (N_21497,N_17990,N_18556);
nand U21498 (N_21498,N_19447,N_19547);
nor U21499 (N_21499,N_19565,N_19216);
nor U21500 (N_21500,N_18392,N_17890);
nand U21501 (N_21501,N_17732,N_17884);
and U21502 (N_21502,N_19616,N_18368);
xnor U21503 (N_21503,N_18707,N_17886);
or U21504 (N_21504,N_19530,N_17748);
and U21505 (N_21505,N_18263,N_18145);
nand U21506 (N_21506,N_18984,N_18951);
nand U21507 (N_21507,N_19111,N_19339);
and U21508 (N_21508,N_17784,N_19032);
nor U21509 (N_21509,N_18485,N_18720);
nor U21510 (N_21510,N_17914,N_18514);
nand U21511 (N_21511,N_18853,N_17804);
and U21512 (N_21512,N_19744,N_18465);
nor U21513 (N_21513,N_18564,N_19446);
xnor U21514 (N_21514,N_17776,N_19970);
nor U21515 (N_21515,N_18315,N_19913);
nand U21516 (N_21516,N_18514,N_19954);
or U21517 (N_21517,N_19639,N_18984);
nand U21518 (N_21518,N_19726,N_18502);
xnor U21519 (N_21519,N_17858,N_19121);
xnor U21520 (N_21520,N_19680,N_17642);
or U21521 (N_21521,N_19383,N_19761);
nor U21522 (N_21522,N_19869,N_19729);
nand U21523 (N_21523,N_19717,N_17923);
and U21524 (N_21524,N_19699,N_19222);
nand U21525 (N_21525,N_19257,N_19165);
or U21526 (N_21526,N_18027,N_18595);
or U21527 (N_21527,N_18067,N_19130);
or U21528 (N_21528,N_18429,N_18367);
xnor U21529 (N_21529,N_19331,N_18404);
and U21530 (N_21530,N_19010,N_19506);
or U21531 (N_21531,N_18147,N_18496);
nor U21532 (N_21532,N_19989,N_19401);
xnor U21533 (N_21533,N_19496,N_18973);
or U21534 (N_21534,N_18819,N_18921);
nand U21535 (N_21535,N_18162,N_19724);
nor U21536 (N_21536,N_17508,N_19626);
nand U21537 (N_21537,N_18326,N_19535);
xor U21538 (N_21538,N_19727,N_17727);
xor U21539 (N_21539,N_17696,N_19689);
nor U21540 (N_21540,N_18722,N_19568);
nor U21541 (N_21541,N_18245,N_19137);
xor U21542 (N_21542,N_19472,N_19417);
nand U21543 (N_21543,N_18406,N_19254);
or U21544 (N_21544,N_18836,N_19837);
nor U21545 (N_21545,N_18268,N_17811);
nand U21546 (N_21546,N_17571,N_17621);
nand U21547 (N_21547,N_19316,N_19854);
nor U21548 (N_21548,N_17520,N_19780);
nor U21549 (N_21549,N_19917,N_19589);
or U21550 (N_21550,N_17614,N_19019);
or U21551 (N_21551,N_18327,N_17866);
nor U21552 (N_21552,N_17581,N_18688);
xor U21553 (N_21553,N_19527,N_17955);
nand U21554 (N_21554,N_19747,N_18001);
nor U21555 (N_21555,N_18355,N_17892);
or U21556 (N_21556,N_17589,N_18000);
nand U21557 (N_21557,N_18165,N_19450);
nand U21558 (N_21558,N_19859,N_18461);
and U21559 (N_21559,N_18986,N_18740);
and U21560 (N_21560,N_19600,N_19140);
or U21561 (N_21561,N_18751,N_19688);
or U21562 (N_21562,N_19539,N_19376);
xor U21563 (N_21563,N_18138,N_19951);
xor U21564 (N_21564,N_19204,N_19069);
nand U21565 (N_21565,N_19130,N_19832);
nor U21566 (N_21566,N_18187,N_18142);
nor U21567 (N_21567,N_18303,N_18396);
nor U21568 (N_21568,N_19968,N_19061);
nand U21569 (N_21569,N_19673,N_19731);
and U21570 (N_21570,N_17926,N_19647);
nor U21571 (N_21571,N_18880,N_19602);
nor U21572 (N_21572,N_18404,N_19252);
nand U21573 (N_21573,N_17881,N_17987);
xnor U21574 (N_21574,N_17606,N_17803);
nor U21575 (N_21575,N_17690,N_18440);
xor U21576 (N_21576,N_19627,N_18824);
and U21577 (N_21577,N_17688,N_17746);
and U21578 (N_21578,N_19195,N_18975);
xor U21579 (N_21579,N_18898,N_18472);
xor U21580 (N_21580,N_17821,N_19138);
xnor U21581 (N_21581,N_18975,N_17878);
nor U21582 (N_21582,N_19336,N_18403);
nand U21583 (N_21583,N_19572,N_18872);
xor U21584 (N_21584,N_17576,N_18491);
nor U21585 (N_21585,N_18549,N_19276);
or U21586 (N_21586,N_18279,N_18464);
and U21587 (N_21587,N_18808,N_19382);
nand U21588 (N_21588,N_19336,N_18836);
nand U21589 (N_21589,N_18867,N_17611);
nor U21590 (N_21590,N_19566,N_17953);
nand U21591 (N_21591,N_17720,N_18508);
and U21592 (N_21592,N_18770,N_18418);
nand U21593 (N_21593,N_17634,N_19123);
xnor U21594 (N_21594,N_17708,N_18904);
nand U21595 (N_21595,N_17665,N_17977);
nor U21596 (N_21596,N_19092,N_19753);
nand U21597 (N_21597,N_17929,N_19764);
nor U21598 (N_21598,N_17726,N_18529);
nor U21599 (N_21599,N_18150,N_19912);
or U21600 (N_21600,N_18938,N_17515);
or U21601 (N_21601,N_19705,N_19821);
and U21602 (N_21602,N_19678,N_17604);
xnor U21603 (N_21603,N_17935,N_18939);
nand U21604 (N_21604,N_19830,N_19667);
and U21605 (N_21605,N_18492,N_19726);
or U21606 (N_21606,N_19229,N_19386);
nor U21607 (N_21607,N_18650,N_18212);
xor U21608 (N_21608,N_17506,N_18813);
nand U21609 (N_21609,N_17520,N_19491);
or U21610 (N_21610,N_19775,N_17844);
nor U21611 (N_21611,N_18823,N_19087);
nor U21612 (N_21612,N_19829,N_19101);
and U21613 (N_21613,N_18687,N_18169);
nand U21614 (N_21614,N_17518,N_19728);
nand U21615 (N_21615,N_18922,N_17526);
xnor U21616 (N_21616,N_18115,N_19732);
nand U21617 (N_21617,N_18310,N_18516);
or U21618 (N_21618,N_19868,N_19427);
and U21619 (N_21619,N_17940,N_19123);
nor U21620 (N_21620,N_17752,N_18203);
nand U21621 (N_21621,N_17986,N_18059);
xor U21622 (N_21622,N_18225,N_18577);
nand U21623 (N_21623,N_19664,N_19204);
and U21624 (N_21624,N_19865,N_18800);
and U21625 (N_21625,N_18170,N_18888);
xnor U21626 (N_21626,N_18457,N_18283);
nand U21627 (N_21627,N_18349,N_19234);
and U21628 (N_21628,N_19907,N_19526);
or U21629 (N_21629,N_19141,N_18518);
nor U21630 (N_21630,N_18389,N_18571);
xnor U21631 (N_21631,N_19413,N_17765);
and U21632 (N_21632,N_19005,N_18562);
nand U21633 (N_21633,N_19869,N_18546);
nor U21634 (N_21634,N_19654,N_18742);
or U21635 (N_21635,N_18495,N_19500);
xnor U21636 (N_21636,N_18647,N_17803);
or U21637 (N_21637,N_19701,N_18350);
nand U21638 (N_21638,N_17597,N_18259);
and U21639 (N_21639,N_18429,N_17638);
or U21640 (N_21640,N_18116,N_18597);
or U21641 (N_21641,N_19035,N_18917);
nand U21642 (N_21642,N_19483,N_19066);
or U21643 (N_21643,N_19067,N_18805);
and U21644 (N_21644,N_19480,N_19991);
and U21645 (N_21645,N_19100,N_18390);
or U21646 (N_21646,N_19687,N_17835);
or U21647 (N_21647,N_18279,N_18158);
nand U21648 (N_21648,N_18341,N_19629);
and U21649 (N_21649,N_19588,N_19792);
xor U21650 (N_21650,N_18908,N_18647);
nand U21651 (N_21651,N_19557,N_19301);
nand U21652 (N_21652,N_17828,N_18259);
xnor U21653 (N_21653,N_18450,N_18177);
nand U21654 (N_21654,N_19675,N_19831);
xnor U21655 (N_21655,N_18584,N_17540);
nand U21656 (N_21656,N_17597,N_18962);
nor U21657 (N_21657,N_19289,N_19685);
nor U21658 (N_21658,N_19249,N_19978);
xor U21659 (N_21659,N_18901,N_19711);
xnor U21660 (N_21660,N_18532,N_19927);
nor U21661 (N_21661,N_18156,N_18292);
or U21662 (N_21662,N_18374,N_19087);
nor U21663 (N_21663,N_18676,N_18008);
and U21664 (N_21664,N_18074,N_18408);
nand U21665 (N_21665,N_18481,N_19044);
or U21666 (N_21666,N_17977,N_19901);
nand U21667 (N_21667,N_18533,N_17551);
and U21668 (N_21668,N_19227,N_19509);
nand U21669 (N_21669,N_19874,N_18597);
xnor U21670 (N_21670,N_18616,N_18531);
and U21671 (N_21671,N_19999,N_19403);
nor U21672 (N_21672,N_18758,N_17949);
or U21673 (N_21673,N_17624,N_19220);
nand U21674 (N_21674,N_17963,N_19784);
and U21675 (N_21675,N_17960,N_19611);
nand U21676 (N_21676,N_18727,N_19817);
nand U21677 (N_21677,N_18080,N_18146);
and U21678 (N_21678,N_18455,N_19077);
xor U21679 (N_21679,N_19366,N_19835);
nor U21680 (N_21680,N_18280,N_18051);
nor U21681 (N_21681,N_18486,N_17694);
or U21682 (N_21682,N_19080,N_19749);
and U21683 (N_21683,N_17685,N_17519);
nand U21684 (N_21684,N_17512,N_17904);
and U21685 (N_21685,N_18662,N_17625);
nand U21686 (N_21686,N_19903,N_19999);
nand U21687 (N_21687,N_19191,N_19808);
xnor U21688 (N_21688,N_18249,N_19325);
xor U21689 (N_21689,N_19793,N_17542);
xnor U21690 (N_21690,N_19527,N_18581);
nand U21691 (N_21691,N_18309,N_19332);
xnor U21692 (N_21692,N_18856,N_19917);
xor U21693 (N_21693,N_19581,N_18789);
xnor U21694 (N_21694,N_17701,N_18356);
and U21695 (N_21695,N_18568,N_18497);
xor U21696 (N_21696,N_18485,N_17963);
and U21697 (N_21697,N_18948,N_19948);
or U21698 (N_21698,N_19926,N_19335);
nor U21699 (N_21699,N_18327,N_17572);
and U21700 (N_21700,N_19345,N_18372);
xnor U21701 (N_21701,N_18599,N_18050);
nor U21702 (N_21702,N_19229,N_19721);
nor U21703 (N_21703,N_19056,N_19232);
and U21704 (N_21704,N_19823,N_19588);
nand U21705 (N_21705,N_18653,N_18922);
nor U21706 (N_21706,N_18089,N_19800);
and U21707 (N_21707,N_19980,N_19814);
xor U21708 (N_21708,N_18986,N_18713);
and U21709 (N_21709,N_18457,N_18603);
nor U21710 (N_21710,N_19446,N_18824);
xnor U21711 (N_21711,N_19007,N_18706);
nand U21712 (N_21712,N_18819,N_17891);
and U21713 (N_21713,N_17514,N_18904);
nand U21714 (N_21714,N_17629,N_18139);
nand U21715 (N_21715,N_19355,N_19241);
xnor U21716 (N_21716,N_17777,N_17952);
or U21717 (N_21717,N_17714,N_19647);
and U21718 (N_21718,N_18903,N_18290);
or U21719 (N_21719,N_17729,N_19698);
nor U21720 (N_21720,N_19401,N_18698);
and U21721 (N_21721,N_17899,N_17875);
or U21722 (N_21722,N_18650,N_18202);
and U21723 (N_21723,N_18103,N_19953);
nand U21724 (N_21724,N_19679,N_19348);
nor U21725 (N_21725,N_18511,N_17860);
nand U21726 (N_21726,N_18608,N_17682);
nand U21727 (N_21727,N_19333,N_19447);
nor U21728 (N_21728,N_19375,N_18412);
nand U21729 (N_21729,N_19082,N_18510);
nand U21730 (N_21730,N_17874,N_18610);
nand U21731 (N_21731,N_19904,N_17623);
nand U21732 (N_21732,N_18324,N_18956);
xnor U21733 (N_21733,N_19765,N_19860);
and U21734 (N_21734,N_17994,N_18785);
and U21735 (N_21735,N_19253,N_19181);
nor U21736 (N_21736,N_18275,N_19594);
nand U21737 (N_21737,N_18221,N_18330);
or U21738 (N_21738,N_17981,N_18201);
nand U21739 (N_21739,N_19022,N_18951);
nand U21740 (N_21740,N_18822,N_17975);
or U21741 (N_21741,N_19078,N_19950);
xor U21742 (N_21742,N_18277,N_18654);
xnor U21743 (N_21743,N_18928,N_18161);
xor U21744 (N_21744,N_18826,N_19218);
nand U21745 (N_21745,N_18248,N_18842);
and U21746 (N_21746,N_17918,N_18507);
xnor U21747 (N_21747,N_17787,N_18529);
and U21748 (N_21748,N_19840,N_17770);
xnor U21749 (N_21749,N_19709,N_17859);
xnor U21750 (N_21750,N_18130,N_18816);
nor U21751 (N_21751,N_18901,N_19544);
and U21752 (N_21752,N_18026,N_17781);
nand U21753 (N_21753,N_17850,N_19560);
nor U21754 (N_21754,N_18250,N_18858);
or U21755 (N_21755,N_17988,N_17669);
and U21756 (N_21756,N_19773,N_17614);
or U21757 (N_21757,N_19828,N_19961);
and U21758 (N_21758,N_19537,N_17809);
and U21759 (N_21759,N_18699,N_19380);
or U21760 (N_21760,N_18617,N_17644);
nor U21761 (N_21761,N_19318,N_19616);
nor U21762 (N_21762,N_19772,N_18851);
or U21763 (N_21763,N_18104,N_19220);
and U21764 (N_21764,N_17952,N_19514);
and U21765 (N_21765,N_18155,N_19740);
or U21766 (N_21766,N_18316,N_18682);
nand U21767 (N_21767,N_19747,N_19873);
nor U21768 (N_21768,N_19608,N_17624);
or U21769 (N_21769,N_18169,N_18542);
nand U21770 (N_21770,N_19319,N_19170);
or U21771 (N_21771,N_18887,N_19788);
and U21772 (N_21772,N_18667,N_19854);
and U21773 (N_21773,N_19056,N_17694);
and U21774 (N_21774,N_18156,N_19575);
xor U21775 (N_21775,N_17681,N_17617);
or U21776 (N_21776,N_18932,N_19138);
and U21777 (N_21777,N_18807,N_18567);
nand U21778 (N_21778,N_17695,N_18980);
nand U21779 (N_21779,N_19422,N_19259);
nand U21780 (N_21780,N_18955,N_19204);
nor U21781 (N_21781,N_18346,N_19986);
and U21782 (N_21782,N_18934,N_18875);
and U21783 (N_21783,N_17740,N_19491);
and U21784 (N_21784,N_19152,N_17781);
xor U21785 (N_21785,N_18977,N_19297);
or U21786 (N_21786,N_18872,N_18657);
xor U21787 (N_21787,N_18564,N_18338);
and U21788 (N_21788,N_19365,N_19312);
xnor U21789 (N_21789,N_18467,N_19482);
or U21790 (N_21790,N_19711,N_19870);
or U21791 (N_21791,N_19589,N_17899);
and U21792 (N_21792,N_18346,N_19293);
and U21793 (N_21793,N_18099,N_17831);
xnor U21794 (N_21794,N_19329,N_18542);
or U21795 (N_21795,N_19644,N_18527);
nand U21796 (N_21796,N_17876,N_19267);
xnor U21797 (N_21797,N_19640,N_18500);
nor U21798 (N_21798,N_19927,N_17778);
nor U21799 (N_21799,N_18481,N_17782);
xor U21800 (N_21800,N_19901,N_18590);
or U21801 (N_21801,N_18476,N_19069);
nand U21802 (N_21802,N_17921,N_19427);
xor U21803 (N_21803,N_18782,N_18721);
or U21804 (N_21804,N_18921,N_18111);
nor U21805 (N_21805,N_18770,N_18105);
and U21806 (N_21806,N_18307,N_17795);
or U21807 (N_21807,N_18529,N_19986);
or U21808 (N_21808,N_17781,N_19209);
and U21809 (N_21809,N_17557,N_19392);
nand U21810 (N_21810,N_19522,N_18432);
or U21811 (N_21811,N_19440,N_19066);
xnor U21812 (N_21812,N_19903,N_18569);
and U21813 (N_21813,N_18093,N_18679);
nor U21814 (N_21814,N_18830,N_19313);
nor U21815 (N_21815,N_17584,N_18537);
or U21816 (N_21816,N_19328,N_18843);
nand U21817 (N_21817,N_18420,N_18893);
nor U21818 (N_21818,N_17544,N_19067);
nor U21819 (N_21819,N_19542,N_19970);
and U21820 (N_21820,N_18827,N_17705);
or U21821 (N_21821,N_19563,N_18653);
and U21822 (N_21822,N_17972,N_19071);
nor U21823 (N_21823,N_19591,N_19545);
xor U21824 (N_21824,N_18282,N_18845);
nor U21825 (N_21825,N_18500,N_18057);
and U21826 (N_21826,N_19906,N_19575);
nor U21827 (N_21827,N_18217,N_19490);
and U21828 (N_21828,N_18150,N_18877);
or U21829 (N_21829,N_18084,N_19820);
nand U21830 (N_21830,N_19258,N_18896);
xnor U21831 (N_21831,N_17712,N_17582);
nor U21832 (N_21832,N_17571,N_18441);
xnor U21833 (N_21833,N_17701,N_17940);
and U21834 (N_21834,N_17501,N_18562);
and U21835 (N_21835,N_18792,N_18277);
nor U21836 (N_21836,N_18904,N_19618);
xor U21837 (N_21837,N_18726,N_18191);
xnor U21838 (N_21838,N_18139,N_19671);
and U21839 (N_21839,N_19400,N_19312);
and U21840 (N_21840,N_18796,N_19435);
and U21841 (N_21841,N_19551,N_19384);
nand U21842 (N_21842,N_18928,N_19231);
nor U21843 (N_21843,N_19671,N_18930);
xnor U21844 (N_21844,N_18389,N_18179);
and U21845 (N_21845,N_19560,N_19577);
xor U21846 (N_21846,N_19061,N_19999);
and U21847 (N_21847,N_17647,N_19982);
or U21848 (N_21848,N_18645,N_19537);
and U21849 (N_21849,N_18026,N_18046);
nand U21850 (N_21850,N_19114,N_18014);
xnor U21851 (N_21851,N_17972,N_18854);
nor U21852 (N_21852,N_19182,N_18119);
nor U21853 (N_21853,N_19054,N_18018);
and U21854 (N_21854,N_19481,N_18673);
nor U21855 (N_21855,N_17912,N_17530);
xnor U21856 (N_21856,N_18736,N_17628);
xnor U21857 (N_21857,N_19917,N_17764);
nand U21858 (N_21858,N_19872,N_17934);
and U21859 (N_21859,N_17874,N_18875);
or U21860 (N_21860,N_19614,N_19985);
nand U21861 (N_21861,N_18137,N_17531);
or U21862 (N_21862,N_19041,N_18322);
xor U21863 (N_21863,N_18697,N_19204);
or U21864 (N_21864,N_18988,N_19871);
nor U21865 (N_21865,N_18475,N_17735);
nand U21866 (N_21866,N_18369,N_18361);
nor U21867 (N_21867,N_19581,N_18997);
or U21868 (N_21868,N_19556,N_18195);
xor U21869 (N_21869,N_18483,N_17610);
nor U21870 (N_21870,N_18522,N_19341);
and U21871 (N_21871,N_18473,N_17930);
nand U21872 (N_21872,N_19600,N_19295);
nand U21873 (N_21873,N_19435,N_17511);
nor U21874 (N_21874,N_19905,N_18889);
nand U21875 (N_21875,N_17994,N_17908);
nor U21876 (N_21876,N_19774,N_17777);
or U21877 (N_21877,N_19503,N_19940);
xnor U21878 (N_21878,N_17988,N_19335);
nand U21879 (N_21879,N_18829,N_19145);
nand U21880 (N_21880,N_18356,N_17686);
nor U21881 (N_21881,N_19899,N_17794);
and U21882 (N_21882,N_17628,N_18202);
nor U21883 (N_21883,N_18703,N_19176);
nor U21884 (N_21884,N_18111,N_18827);
nand U21885 (N_21885,N_17726,N_19119);
and U21886 (N_21886,N_18680,N_19629);
and U21887 (N_21887,N_18094,N_19303);
nand U21888 (N_21888,N_19628,N_18258);
or U21889 (N_21889,N_18898,N_17961);
or U21890 (N_21890,N_18443,N_19721);
xor U21891 (N_21891,N_19178,N_17508);
or U21892 (N_21892,N_19196,N_18781);
nand U21893 (N_21893,N_17512,N_19909);
nand U21894 (N_21894,N_17790,N_19854);
and U21895 (N_21895,N_17745,N_18493);
nor U21896 (N_21896,N_18704,N_19086);
and U21897 (N_21897,N_17669,N_19866);
nor U21898 (N_21898,N_18067,N_17667);
or U21899 (N_21899,N_18219,N_19345);
and U21900 (N_21900,N_19716,N_17503);
nand U21901 (N_21901,N_18562,N_17573);
nor U21902 (N_21902,N_18198,N_19205);
xor U21903 (N_21903,N_17560,N_18716);
and U21904 (N_21904,N_19866,N_18839);
nor U21905 (N_21905,N_19566,N_17622);
xnor U21906 (N_21906,N_18751,N_18825);
nand U21907 (N_21907,N_17968,N_19721);
and U21908 (N_21908,N_18821,N_18226);
or U21909 (N_21909,N_19866,N_19570);
xnor U21910 (N_21910,N_18825,N_19970);
or U21911 (N_21911,N_19877,N_18002);
xor U21912 (N_21912,N_18953,N_18275);
nand U21913 (N_21913,N_18731,N_17644);
xnor U21914 (N_21914,N_17945,N_19367);
and U21915 (N_21915,N_17920,N_18815);
xnor U21916 (N_21916,N_18857,N_18332);
xnor U21917 (N_21917,N_19931,N_19291);
nor U21918 (N_21918,N_17787,N_18507);
and U21919 (N_21919,N_19517,N_17664);
or U21920 (N_21920,N_18373,N_18274);
nor U21921 (N_21921,N_19350,N_19536);
nor U21922 (N_21922,N_19266,N_19568);
or U21923 (N_21923,N_19585,N_18086);
or U21924 (N_21924,N_18351,N_19401);
nor U21925 (N_21925,N_18535,N_18873);
nand U21926 (N_21926,N_17898,N_17657);
and U21927 (N_21927,N_18675,N_19803);
nor U21928 (N_21928,N_18347,N_17816);
xor U21929 (N_21929,N_17625,N_19450);
nand U21930 (N_21930,N_17621,N_17572);
nor U21931 (N_21931,N_18025,N_19734);
xor U21932 (N_21932,N_18216,N_18541);
and U21933 (N_21933,N_19460,N_17597);
nand U21934 (N_21934,N_18672,N_18544);
xor U21935 (N_21935,N_19874,N_18990);
or U21936 (N_21936,N_17513,N_19987);
xnor U21937 (N_21937,N_17743,N_17824);
nand U21938 (N_21938,N_19418,N_19962);
nor U21939 (N_21939,N_17508,N_18119);
nand U21940 (N_21940,N_18802,N_18720);
and U21941 (N_21941,N_19306,N_18453);
xnor U21942 (N_21942,N_19337,N_19308);
and U21943 (N_21943,N_18229,N_18403);
nor U21944 (N_21944,N_19997,N_19595);
or U21945 (N_21945,N_19425,N_19054);
or U21946 (N_21946,N_19150,N_17718);
or U21947 (N_21947,N_18638,N_19783);
or U21948 (N_21948,N_18225,N_19622);
or U21949 (N_21949,N_17579,N_19951);
nand U21950 (N_21950,N_19674,N_19619);
nor U21951 (N_21951,N_18439,N_18300);
nand U21952 (N_21952,N_18652,N_19092);
and U21953 (N_21953,N_19397,N_19072);
or U21954 (N_21954,N_17626,N_19287);
xnor U21955 (N_21955,N_17751,N_19123);
or U21956 (N_21956,N_17750,N_18676);
nand U21957 (N_21957,N_19421,N_18695);
and U21958 (N_21958,N_18847,N_19888);
and U21959 (N_21959,N_18146,N_18634);
nand U21960 (N_21960,N_17872,N_18066);
xor U21961 (N_21961,N_17705,N_18416);
xnor U21962 (N_21962,N_18388,N_18091);
nand U21963 (N_21963,N_17707,N_19851);
and U21964 (N_21964,N_17710,N_19072);
and U21965 (N_21965,N_18971,N_18216);
and U21966 (N_21966,N_19823,N_19960);
xnor U21967 (N_21967,N_18624,N_19981);
nand U21968 (N_21968,N_19989,N_18186);
xnor U21969 (N_21969,N_18694,N_18350);
and U21970 (N_21970,N_18386,N_19992);
nor U21971 (N_21971,N_17624,N_18109);
nor U21972 (N_21972,N_19898,N_19058);
or U21973 (N_21973,N_18755,N_18916);
or U21974 (N_21974,N_17811,N_18284);
and U21975 (N_21975,N_18725,N_19817);
nand U21976 (N_21976,N_19064,N_17764);
xnor U21977 (N_21977,N_19406,N_18536);
or U21978 (N_21978,N_17808,N_18857);
and U21979 (N_21979,N_17632,N_19821);
or U21980 (N_21980,N_19368,N_19111);
and U21981 (N_21981,N_18511,N_19143);
and U21982 (N_21982,N_19443,N_17852);
nand U21983 (N_21983,N_18110,N_19103);
xnor U21984 (N_21984,N_17507,N_18275);
or U21985 (N_21985,N_19500,N_17843);
xnor U21986 (N_21986,N_18108,N_17776);
nor U21987 (N_21987,N_17715,N_18050);
nor U21988 (N_21988,N_18231,N_19785);
and U21989 (N_21989,N_18837,N_18482);
and U21990 (N_21990,N_18335,N_19296);
or U21991 (N_21991,N_19440,N_17709);
nand U21992 (N_21992,N_19034,N_19333);
and U21993 (N_21993,N_17741,N_18633);
nor U21994 (N_21994,N_17806,N_18996);
or U21995 (N_21995,N_19109,N_19118);
and U21996 (N_21996,N_19750,N_18555);
nand U21997 (N_21997,N_19008,N_19553);
or U21998 (N_21998,N_17962,N_18063);
and U21999 (N_21999,N_18616,N_19739);
and U22000 (N_22000,N_18425,N_17621);
or U22001 (N_22001,N_17509,N_18709);
nand U22002 (N_22002,N_17888,N_18132);
nand U22003 (N_22003,N_17786,N_18762);
and U22004 (N_22004,N_18467,N_17586);
nor U22005 (N_22005,N_18962,N_18940);
nor U22006 (N_22006,N_18656,N_19465);
or U22007 (N_22007,N_19632,N_19912);
or U22008 (N_22008,N_18263,N_17562);
and U22009 (N_22009,N_17872,N_19125);
nand U22010 (N_22010,N_19991,N_19037);
nand U22011 (N_22011,N_19577,N_18061);
xnor U22012 (N_22012,N_19561,N_18944);
nor U22013 (N_22013,N_17965,N_19939);
xor U22014 (N_22014,N_19239,N_18071);
nor U22015 (N_22015,N_19457,N_18745);
and U22016 (N_22016,N_19054,N_18485);
or U22017 (N_22017,N_18699,N_19370);
nand U22018 (N_22018,N_18589,N_18175);
or U22019 (N_22019,N_18839,N_18332);
xor U22020 (N_22020,N_19697,N_19129);
xnor U22021 (N_22021,N_17673,N_18717);
nand U22022 (N_22022,N_17850,N_17655);
or U22023 (N_22023,N_19635,N_19222);
xnor U22024 (N_22024,N_18221,N_17512);
xor U22025 (N_22025,N_18196,N_17880);
or U22026 (N_22026,N_18102,N_19971);
nand U22027 (N_22027,N_19897,N_18423);
and U22028 (N_22028,N_19191,N_19801);
nand U22029 (N_22029,N_19493,N_18515);
xor U22030 (N_22030,N_18315,N_19836);
nor U22031 (N_22031,N_17770,N_18760);
nand U22032 (N_22032,N_19041,N_19419);
nand U22033 (N_22033,N_18127,N_18907);
nor U22034 (N_22034,N_18858,N_19420);
and U22035 (N_22035,N_17871,N_18017);
nand U22036 (N_22036,N_18772,N_17515);
and U22037 (N_22037,N_19468,N_17939);
nand U22038 (N_22038,N_18444,N_19186);
or U22039 (N_22039,N_17819,N_17834);
or U22040 (N_22040,N_19261,N_18139);
or U22041 (N_22041,N_19470,N_19453);
nor U22042 (N_22042,N_19038,N_19394);
or U22043 (N_22043,N_18987,N_19092);
nor U22044 (N_22044,N_18080,N_18279);
xnor U22045 (N_22045,N_19826,N_19624);
nand U22046 (N_22046,N_18505,N_18983);
nor U22047 (N_22047,N_19844,N_19001);
xor U22048 (N_22048,N_18512,N_19124);
nand U22049 (N_22049,N_19454,N_19450);
or U22050 (N_22050,N_18945,N_19733);
xnor U22051 (N_22051,N_18802,N_18500);
nor U22052 (N_22052,N_19918,N_19984);
nor U22053 (N_22053,N_18901,N_17647);
nand U22054 (N_22054,N_17760,N_17674);
xnor U22055 (N_22055,N_18857,N_18566);
nor U22056 (N_22056,N_18485,N_17730);
or U22057 (N_22057,N_18273,N_18708);
xor U22058 (N_22058,N_18725,N_19545);
and U22059 (N_22059,N_18873,N_18170);
nand U22060 (N_22060,N_17640,N_17747);
nand U22061 (N_22061,N_18653,N_19641);
xnor U22062 (N_22062,N_19912,N_17748);
nor U22063 (N_22063,N_19383,N_19577);
and U22064 (N_22064,N_19152,N_19191);
or U22065 (N_22065,N_19499,N_19405);
nor U22066 (N_22066,N_19357,N_18962);
and U22067 (N_22067,N_17864,N_19151);
or U22068 (N_22068,N_18313,N_19778);
nand U22069 (N_22069,N_18579,N_17547);
xor U22070 (N_22070,N_19333,N_19337);
nand U22071 (N_22071,N_17688,N_18929);
nor U22072 (N_22072,N_18174,N_18054);
or U22073 (N_22073,N_17668,N_17850);
or U22074 (N_22074,N_18828,N_18765);
nand U22075 (N_22075,N_18562,N_17867);
xor U22076 (N_22076,N_18408,N_18815);
and U22077 (N_22077,N_18516,N_18355);
nand U22078 (N_22078,N_18665,N_19876);
and U22079 (N_22079,N_17908,N_19268);
or U22080 (N_22080,N_19538,N_19824);
xor U22081 (N_22081,N_19743,N_19314);
xor U22082 (N_22082,N_19761,N_19360);
xor U22083 (N_22083,N_19883,N_18699);
nor U22084 (N_22084,N_19945,N_17804);
xnor U22085 (N_22085,N_18648,N_18586);
and U22086 (N_22086,N_18503,N_19326);
nand U22087 (N_22087,N_19214,N_18808);
and U22088 (N_22088,N_17602,N_19953);
and U22089 (N_22089,N_19174,N_17558);
nand U22090 (N_22090,N_18643,N_19478);
or U22091 (N_22091,N_18663,N_19790);
and U22092 (N_22092,N_17645,N_19207);
and U22093 (N_22093,N_19597,N_19855);
nor U22094 (N_22094,N_17743,N_19944);
or U22095 (N_22095,N_18715,N_18597);
nand U22096 (N_22096,N_17567,N_18014);
or U22097 (N_22097,N_19239,N_19537);
nand U22098 (N_22098,N_18662,N_19896);
or U22099 (N_22099,N_18385,N_18233);
xor U22100 (N_22100,N_17786,N_19893);
xnor U22101 (N_22101,N_18188,N_17789);
nand U22102 (N_22102,N_19880,N_19849);
nand U22103 (N_22103,N_19392,N_19298);
xnor U22104 (N_22104,N_18401,N_19767);
and U22105 (N_22105,N_18003,N_18405);
xnor U22106 (N_22106,N_19446,N_18907);
and U22107 (N_22107,N_18977,N_18473);
nor U22108 (N_22108,N_17689,N_18987);
xnor U22109 (N_22109,N_19266,N_18547);
nor U22110 (N_22110,N_18263,N_17661);
xnor U22111 (N_22111,N_19890,N_18031);
and U22112 (N_22112,N_18369,N_18455);
nand U22113 (N_22113,N_18452,N_17821);
and U22114 (N_22114,N_18265,N_18722);
xnor U22115 (N_22115,N_18486,N_19919);
xnor U22116 (N_22116,N_17689,N_17838);
nand U22117 (N_22117,N_17895,N_18276);
nor U22118 (N_22118,N_18951,N_19863);
and U22119 (N_22119,N_19067,N_18579);
nand U22120 (N_22120,N_18233,N_18242);
or U22121 (N_22121,N_18236,N_18723);
or U22122 (N_22122,N_19871,N_19219);
or U22123 (N_22123,N_19076,N_18004);
xnor U22124 (N_22124,N_18643,N_19011);
nor U22125 (N_22125,N_18657,N_18433);
nand U22126 (N_22126,N_19049,N_19161);
nor U22127 (N_22127,N_17724,N_19609);
or U22128 (N_22128,N_18542,N_18297);
and U22129 (N_22129,N_18621,N_17942);
and U22130 (N_22130,N_17899,N_19260);
nor U22131 (N_22131,N_19265,N_19874);
nor U22132 (N_22132,N_17699,N_19940);
nand U22133 (N_22133,N_17931,N_17569);
nand U22134 (N_22134,N_19750,N_19058);
xor U22135 (N_22135,N_19954,N_18757);
xor U22136 (N_22136,N_19693,N_19329);
and U22137 (N_22137,N_18560,N_18097);
nor U22138 (N_22138,N_19169,N_18209);
nand U22139 (N_22139,N_19913,N_18110);
or U22140 (N_22140,N_17909,N_18871);
and U22141 (N_22141,N_18505,N_19662);
nand U22142 (N_22142,N_17696,N_17993);
nand U22143 (N_22143,N_17780,N_19863);
nand U22144 (N_22144,N_17916,N_18461);
xor U22145 (N_22145,N_18109,N_18466);
and U22146 (N_22146,N_17774,N_17758);
nand U22147 (N_22147,N_18409,N_18820);
nand U22148 (N_22148,N_19063,N_18056);
nand U22149 (N_22149,N_19897,N_19393);
or U22150 (N_22150,N_19858,N_17809);
xor U22151 (N_22151,N_19244,N_19205);
or U22152 (N_22152,N_19082,N_18909);
xnor U22153 (N_22153,N_19109,N_18898);
nor U22154 (N_22154,N_17516,N_19123);
nor U22155 (N_22155,N_18904,N_18436);
and U22156 (N_22156,N_18599,N_18150);
nand U22157 (N_22157,N_19789,N_18117);
nor U22158 (N_22158,N_19613,N_17718);
and U22159 (N_22159,N_17845,N_18790);
and U22160 (N_22160,N_17560,N_19711);
nor U22161 (N_22161,N_19900,N_18962);
or U22162 (N_22162,N_19797,N_18023);
nor U22163 (N_22163,N_18487,N_19869);
or U22164 (N_22164,N_19046,N_19992);
or U22165 (N_22165,N_18721,N_18986);
nor U22166 (N_22166,N_18133,N_17809);
or U22167 (N_22167,N_18935,N_17862);
xor U22168 (N_22168,N_18851,N_18506);
or U22169 (N_22169,N_17747,N_18626);
nand U22170 (N_22170,N_17850,N_19923);
nor U22171 (N_22171,N_18709,N_17723);
xnor U22172 (N_22172,N_18123,N_17937);
nand U22173 (N_22173,N_19900,N_19095);
and U22174 (N_22174,N_19122,N_18017);
xor U22175 (N_22175,N_19260,N_19419);
nor U22176 (N_22176,N_18201,N_19957);
nand U22177 (N_22177,N_19160,N_19526);
nand U22178 (N_22178,N_17538,N_17749);
xnor U22179 (N_22179,N_19156,N_19252);
xor U22180 (N_22180,N_17936,N_19155);
xor U22181 (N_22181,N_18802,N_18576);
and U22182 (N_22182,N_17505,N_18371);
or U22183 (N_22183,N_18404,N_18012);
nand U22184 (N_22184,N_18329,N_17763);
and U22185 (N_22185,N_19633,N_19374);
nor U22186 (N_22186,N_18872,N_17528);
or U22187 (N_22187,N_19591,N_19018);
nor U22188 (N_22188,N_18294,N_18665);
and U22189 (N_22189,N_18599,N_18960);
nor U22190 (N_22190,N_18373,N_18731);
nand U22191 (N_22191,N_19222,N_19076);
nand U22192 (N_22192,N_18533,N_19678);
nand U22193 (N_22193,N_19807,N_18138);
nor U22194 (N_22194,N_19429,N_18404);
nand U22195 (N_22195,N_17918,N_19734);
or U22196 (N_22196,N_19114,N_18773);
and U22197 (N_22197,N_17874,N_18352);
or U22198 (N_22198,N_18494,N_17994);
and U22199 (N_22199,N_18588,N_19224);
xnor U22200 (N_22200,N_18523,N_19023);
or U22201 (N_22201,N_19135,N_18960);
and U22202 (N_22202,N_17742,N_17558);
xnor U22203 (N_22203,N_18771,N_17802);
nand U22204 (N_22204,N_19578,N_19001);
xnor U22205 (N_22205,N_18748,N_17926);
and U22206 (N_22206,N_18323,N_19479);
and U22207 (N_22207,N_19035,N_17781);
nand U22208 (N_22208,N_18057,N_18326);
nand U22209 (N_22209,N_18782,N_19769);
xor U22210 (N_22210,N_19209,N_19301);
nand U22211 (N_22211,N_19718,N_19509);
nor U22212 (N_22212,N_19857,N_17894);
xnor U22213 (N_22213,N_18215,N_19135);
nor U22214 (N_22214,N_17883,N_19224);
or U22215 (N_22215,N_18165,N_19524);
xor U22216 (N_22216,N_17823,N_18027);
and U22217 (N_22217,N_19946,N_19031);
and U22218 (N_22218,N_17824,N_17623);
or U22219 (N_22219,N_17778,N_19457);
or U22220 (N_22220,N_18537,N_19732);
xor U22221 (N_22221,N_18568,N_19581);
xor U22222 (N_22222,N_19592,N_19658);
nand U22223 (N_22223,N_18903,N_18034);
and U22224 (N_22224,N_17734,N_19199);
nor U22225 (N_22225,N_18755,N_19428);
xor U22226 (N_22226,N_19008,N_17664);
nor U22227 (N_22227,N_17625,N_18369);
xnor U22228 (N_22228,N_19185,N_18688);
nor U22229 (N_22229,N_17791,N_17561);
or U22230 (N_22230,N_19188,N_17746);
or U22231 (N_22231,N_19966,N_18830);
xor U22232 (N_22232,N_19217,N_19129);
or U22233 (N_22233,N_18697,N_19054);
nand U22234 (N_22234,N_18564,N_19993);
and U22235 (N_22235,N_19106,N_18780);
nor U22236 (N_22236,N_19587,N_18071);
nor U22237 (N_22237,N_17893,N_19937);
nand U22238 (N_22238,N_18011,N_19966);
and U22239 (N_22239,N_18447,N_18009);
or U22240 (N_22240,N_17781,N_18993);
and U22241 (N_22241,N_19036,N_19214);
and U22242 (N_22242,N_19628,N_18751);
xnor U22243 (N_22243,N_19780,N_19867);
nor U22244 (N_22244,N_17919,N_19276);
xor U22245 (N_22245,N_19078,N_19867);
and U22246 (N_22246,N_19389,N_19778);
nor U22247 (N_22247,N_18143,N_19936);
and U22248 (N_22248,N_19056,N_19340);
or U22249 (N_22249,N_19828,N_18871);
and U22250 (N_22250,N_19667,N_17578);
nor U22251 (N_22251,N_18932,N_17941);
nor U22252 (N_22252,N_17702,N_19418);
nand U22253 (N_22253,N_17686,N_17795);
nor U22254 (N_22254,N_18858,N_17691);
nor U22255 (N_22255,N_19626,N_18282);
nor U22256 (N_22256,N_18814,N_18310);
or U22257 (N_22257,N_18573,N_18604);
nor U22258 (N_22258,N_18591,N_19649);
nor U22259 (N_22259,N_19953,N_19606);
or U22260 (N_22260,N_18267,N_19265);
nand U22261 (N_22261,N_17973,N_19035);
nand U22262 (N_22262,N_18953,N_18260);
or U22263 (N_22263,N_19460,N_18270);
or U22264 (N_22264,N_18350,N_17876);
nand U22265 (N_22265,N_18956,N_17710);
xnor U22266 (N_22266,N_18549,N_19264);
and U22267 (N_22267,N_18781,N_18168);
nand U22268 (N_22268,N_17504,N_17807);
and U22269 (N_22269,N_19160,N_18986);
and U22270 (N_22270,N_19477,N_19167);
nand U22271 (N_22271,N_18779,N_18414);
nor U22272 (N_22272,N_17890,N_18617);
nor U22273 (N_22273,N_18613,N_19120);
nand U22274 (N_22274,N_18292,N_19632);
or U22275 (N_22275,N_19219,N_17567);
and U22276 (N_22276,N_19996,N_18897);
or U22277 (N_22277,N_19198,N_19860);
or U22278 (N_22278,N_18385,N_19144);
or U22279 (N_22279,N_17526,N_17655);
xnor U22280 (N_22280,N_18233,N_18225);
nand U22281 (N_22281,N_18154,N_18799);
xor U22282 (N_22282,N_19912,N_17660);
or U22283 (N_22283,N_18493,N_19692);
xor U22284 (N_22284,N_17587,N_18198);
nor U22285 (N_22285,N_17790,N_19193);
nand U22286 (N_22286,N_19028,N_19791);
xor U22287 (N_22287,N_19697,N_19206);
or U22288 (N_22288,N_18150,N_19306);
or U22289 (N_22289,N_18970,N_18701);
and U22290 (N_22290,N_19130,N_19653);
and U22291 (N_22291,N_17982,N_18363);
or U22292 (N_22292,N_17691,N_18820);
or U22293 (N_22293,N_18107,N_19779);
or U22294 (N_22294,N_19361,N_18447);
xnor U22295 (N_22295,N_19015,N_18617);
nand U22296 (N_22296,N_19566,N_17611);
and U22297 (N_22297,N_19092,N_18928);
xnor U22298 (N_22298,N_19138,N_17655);
or U22299 (N_22299,N_19601,N_18008);
nand U22300 (N_22300,N_18516,N_18246);
xnor U22301 (N_22301,N_18570,N_18450);
or U22302 (N_22302,N_18976,N_19938);
nand U22303 (N_22303,N_17689,N_19714);
xnor U22304 (N_22304,N_18408,N_18730);
nor U22305 (N_22305,N_18934,N_19055);
and U22306 (N_22306,N_17844,N_18383);
xor U22307 (N_22307,N_17919,N_18021);
nor U22308 (N_22308,N_18350,N_19131);
nand U22309 (N_22309,N_17796,N_18320);
nor U22310 (N_22310,N_19499,N_19297);
and U22311 (N_22311,N_18588,N_17945);
or U22312 (N_22312,N_17797,N_18239);
nor U22313 (N_22313,N_17514,N_18542);
nor U22314 (N_22314,N_19289,N_18439);
nand U22315 (N_22315,N_17752,N_19270);
nor U22316 (N_22316,N_18235,N_18725);
xor U22317 (N_22317,N_19126,N_18110);
xnor U22318 (N_22318,N_18707,N_18119);
and U22319 (N_22319,N_19021,N_18377);
or U22320 (N_22320,N_19297,N_19266);
xnor U22321 (N_22321,N_18143,N_19471);
or U22322 (N_22322,N_19115,N_19876);
and U22323 (N_22323,N_19226,N_18342);
nor U22324 (N_22324,N_18164,N_19103);
nor U22325 (N_22325,N_18385,N_17663);
nand U22326 (N_22326,N_19291,N_18095);
xor U22327 (N_22327,N_18038,N_18308);
and U22328 (N_22328,N_17889,N_18195);
or U22329 (N_22329,N_19875,N_19696);
nor U22330 (N_22330,N_18151,N_18539);
xnor U22331 (N_22331,N_19880,N_18021);
or U22332 (N_22332,N_18494,N_18834);
nand U22333 (N_22333,N_19425,N_18958);
nand U22334 (N_22334,N_18550,N_18134);
nand U22335 (N_22335,N_19453,N_18501);
or U22336 (N_22336,N_18652,N_17623);
and U22337 (N_22337,N_18394,N_19511);
xnor U22338 (N_22338,N_17813,N_18319);
xnor U22339 (N_22339,N_17785,N_18921);
nand U22340 (N_22340,N_19487,N_17647);
nand U22341 (N_22341,N_19626,N_19573);
xor U22342 (N_22342,N_19320,N_18425);
or U22343 (N_22343,N_19768,N_17962);
nor U22344 (N_22344,N_18119,N_19002);
xor U22345 (N_22345,N_19219,N_18993);
nor U22346 (N_22346,N_18590,N_18624);
and U22347 (N_22347,N_19654,N_18194);
xor U22348 (N_22348,N_19858,N_17526);
nand U22349 (N_22349,N_17613,N_19591);
and U22350 (N_22350,N_19815,N_17934);
and U22351 (N_22351,N_19597,N_17988);
nor U22352 (N_22352,N_19491,N_18728);
or U22353 (N_22353,N_17507,N_18610);
nor U22354 (N_22354,N_18606,N_17629);
xor U22355 (N_22355,N_18745,N_17991);
nor U22356 (N_22356,N_19475,N_19708);
or U22357 (N_22357,N_18995,N_18047);
nor U22358 (N_22358,N_19887,N_19334);
or U22359 (N_22359,N_17722,N_19524);
nand U22360 (N_22360,N_17881,N_19347);
nand U22361 (N_22361,N_17658,N_18716);
or U22362 (N_22362,N_18471,N_17954);
nor U22363 (N_22363,N_19682,N_19369);
nor U22364 (N_22364,N_19943,N_17825);
nand U22365 (N_22365,N_18856,N_18346);
nand U22366 (N_22366,N_18854,N_19895);
or U22367 (N_22367,N_19797,N_18397);
nor U22368 (N_22368,N_18627,N_17781);
nor U22369 (N_22369,N_18374,N_19304);
nand U22370 (N_22370,N_19274,N_17887);
nor U22371 (N_22371,N_19158,N_17750);
nor U22372 (N_22372,N_18204,N_17994);
xor U22373 (N_22373,N_19172,N_19113);
or U22374 (N_22374,N_17738,N_17729);
xor U22375 (N_22375,N_18148,N_19893);
nor U22376 (N_22376,N_19352,N_17788);
xnor U22377 (N_22377,N_19454,N_19715);
nor U22378 (N_22378,N_19311,N_19273);
nand U22379 (N_22379,N_17850,N_18584);
and U22380 (N_22380,N_18610,N_18076);
nand U22381 (N_22381,N_18944,N_17897);
nand U22382 (N_22382,N_18378,N_18244);
or U22383 (N_22383,N_19310,N_17649);
and U22384 (N_22384,N_18834,N_17572);
nor U22385 (N_22385,N_17603,N_17946);
or U22386 (N_22386,N_17522,N_19106);
nor U22387 (N_22387,N_17918,N_19695);
and U22388 (N_22388,N_18244,N_19822);
or U22389 (N_22389,N_17602,N_18650);
xor U22390 (N_22390,N_17918,N_17731);
xnor U22391 (N_22391,N_18455,N_17504);
xor U22392 (N_22392,N_19026,N_17561);
nor U22393 (N_22393,N_17867,N_19548);
xor U22394 (N_22394,N_18931,N_18141);
and U22395 (N_22395,N_19613,N_18486);
nand U22396 (N_22396,N_17657,N_17835);
xnor U22397 (N_22397,N_19546,N_17521);
or U22398 (N_22398,N_19729,N_18461);
xor U22399 (N_22399,N_19552,N_18686);
nor U22400 (N_22400,N_19725,N_17572);
xor U22401 (N_22401,N_19442,N_19999);
and U22402 (N_22402,N_18338,N_19743);
xor U22403 (N_22403,N_19708,N_19670);
nand U22404 (N_22404,N_17694,N_17928);
or U22405 (N_22405,N_18104,N_18730);
and U22406 (N_22406,N_17691,N_19946);
nand U22407 (N_22407,N_18997,N_18833);
nand U22408 (N_22408,N_17800,N_18527);
nand U22409 (N_22409,N_18750,N_18820);
nor U22410 (N_22410,N_18275,N_17855);
nand U22411 (N_22411,N_18254,N_19729);
nor U22412 (N_22412,N_19768,N_19160);
xnor U22413 (N_22413,N_19736,N_18531);
and U22414 (N_22414,N_17657,N_17551);
xnor U22415 (N_22415,N_19194,N_18523);
xnor U22416 (N_22416,N_19222,N_18348);
xor U22417 (N_22417,N_17591,N_19491);
and U22418 (N_22418,N_18688,N_19938);
nor U22419 (N_22419,N_18857,N_18236);
and U22420 (N_22420,N_18775,N_19850);
nor U22421 (N_22421,N_18102,N_19206);
and U22422 (N_22422,N_19339,N_18883);
nand U22423 (N_22423,N_18778,N_18473);
or U22424 (N_22424,N_18423,N_19853);
xor U22425 (N_22425,N_19376,N_19601);
nor U22426 (N_22426,N_17725,N_19668);
or U22427 (N_22427,N_17717,N_19107);
or U22428 (N_22428,N_19958,N_17611);
xor U22429 (N_22429,N_18075,N_18484);
and U22430 (N_22430,N_19346,N_19500);
nand U22431 (N_22431,N_19719,N_18367);
and U22432 (N_22432,N_19897,N_18246);
nor U22433 (N_22433,N_18196,N_17771);
and U22434 (N_22434,N_17745,N_19718);
nand U22435 (N_22435,N_17613,N_17768);
nor U22436 (N_22436,N_18006,N_17943);
and U22437 (N_22437,N_17560,N_17741);
nand U22438 (N_22438,N_19939,N_19744);
xor U22439 (N_22439,N_17862,N_18100);
nand U22440 (N_22440,N_19604,N_19617);
nor U22441 (N_22441,N_17560,N_19170);
xnor U22442 (N_22442,N_18437,N_19401);
nor U22443 (N_22443,N_18466,N_18797);
xor U22444 (N_22444,N_17855,N_18196);
xor U22445 (N_22445,N_19869,N_19208);
or U22446 (N_22446,N_19924,N_18599);
nand U22447 (N_22447,N_19322,N_18970);
nand U22448 (N_22448,N_18130,N_19196);
xor U22449 (N_22449,N_17976,N_18394);
nand U22450 (N_22450,N_18560,N_17817);
or U22451 (N_22451,N_17969,N_17636);
and U22452 (N_22452,N_19625,N_18821);
nand U22453 (N_22453,N_19196,N_17777);
nand U22454 (N_22454,N_18694,N_17829);
or U22455 (N_22455,N_19267,N_19792);
nand U22456 (N_22456,N_17871,N_17642);
nand U22457 (N_22457,N_17788,N_19710);
xor U22458 (N_22458,N_19634,N_17558);
and U22459 (N_22459,N_17726,N_18354);
or U22460 (N_22460,N_18008,N_18674);
or U22461 (N_22461,N_17690,N_19727);
and U22462 (N_22462,N_18391,N_19013);
nand U22463 (N_22463,N_17871,N_18883);
nor U22464 (N_22464,N_19160,N_19285);
and U22465 (N_22465,N_18128,N_19041);
nand U22466 (N_22466,N_19743,N_17708);
and U22467 (N_22467,N_19458,N_19026);
or U22468 (N_22468,N_19932,N_18109);
nor U22469 (N_22469,N_18727,N_19927);
nor U22470 (N_22470,N_19365,N_18148);
nand U22471 (N_22471,N_19673,N_19923);
xnor U22472 (N_22472,N_17600,N_19649);
xor U22473 (N_22473,N_19991,N_18285);
and U22474 (N_22474,N_19233,N_17923);
nor U22475 (N_22475,N_19509,N_19189);
and U22476 (N_22476,N_18628,N_18871);
nor U22477 (N_22477,N_18407,N_18641);
nand U22478 (N_22478,N_18306,N_19740);
or U22479 (N_22479,N_19875,N_19631);
nor U22480 (N_22480,N_19107,N_18867);
nor U22481 (N_22481,N_19363,N_19184);
nor U22482 (N_22482,N_17978,N_18449);
nor U22483 (N_22483,N_18945,N_17918);
nor U22484 (N_22484,N_17891,N_18257);
nor U22485 (N_22485,N_19515,N_18990);
and U22486 (N_22486,N_19163,N_18824);
or U22487 (N_22487,N_17531,N_17835);
or U22488 (N_22488,N_18047,N_18370);
xnor U22489 (N_22489,N_19544,N_17666);
nor U22490 (N_22490,N_17693,N_18777);
or U22491 (N_22491,N_19006,N_19145);
nand U22492 (N_22492,N_18048,N_17943);
or U22493 (N_22493,N_19395,N_19716);
and U22494 (N_22494,N_18788,N_18700);
xnor U22495 (N_22495,N_18791,N_18376);
or U22496 (N_22496,N_18541,N_19889);
and U22497 (N_22497,N_18355,N_17802);
nand U22498 (N_22498,N_18867,N_18165);
xnor U22499 (N_22499,N_18638,N_17800);
xor U22500 (N_22500,N_20014,N_22072);
and U22501 (N_22501,N_22489,N_21126);
nand U22502 (N_22502,N_22119,N_20318);
nor U22503 (N_22503,N_21395,N_21927);
nand U22504 (N_22504,N_21243,N_22005);
or U22505 (N_22505,N_20310,N_20814);
or U22506 (N_22506,N_20294,N_20855);
xnor U22507 (N_22507,N_21599,N_21042);
nor U22508 (N_22508,N_20158,N_20772);
and U22509 (N_22509,N_20234,N_22090);
xnor U22510 (N_22510,N_21319,N_20382);
nor U22511 (N_22511,N_21058,N_21655);
xnor U22512 (N_22512,N_20571,N_20677);
nand U22513 (N_22513,N_20725,N_20612);
nand U22514 (N_22514,N_20625,N_21161);
or U22515 (N_22515,N_21962,N_21949);
or U22516 (N_22516,N_20050,N_21290);
and U22517 (N_22517,N_20694,N_20272);
and U22518 (N_22518,N_21553,N_22162);
and U22519 (N_22519,N_20140,N_21940);
nor U22520 (N_22520,N_21190,N_22246);
nor U22521 (N_22521,N_21063,N_20912);
nand U22522 (N_22522,N_20941,N_21637);
xnor U22523 (N_22523,N_20371,N_22327);
or U22524 (N_22524,N_22415,N_20184);
nand U22525 (N_22525,N_21414,N_20920);
or U22526 (N_22526,N_21011,N_21277);
xnor U22527 (N_22527,N_21019,N_20118);
and U22528 (N_22528,N_21153,N_20560);
or U22529 (N_22529,N_20596,N_20918);
nand U22530 (N_22530,N_21304,N_21178);
and U22531 (N_22531,N_20674,N_22031);
xnor U22532 (N_22532,N_22495,N_21846);
nor U22533 (N_22533,N_20385,N_21323);
or U22534 (N_22534,N_20559,N_20619);
nand U22535 (N_22535,N_22432,N_21998);
nand U22536 (N_22536,N_22224,N_20945);
or U22537 (N_22537,N_20651,N_21095);
or U22538 (N_22538,N_21316,N_20105);
or U22539 (N_22539,N_20406,N_21738);
or U22540 (N_22540,N_20628,N_20750);
or U22541 (N_22541,N_22176,N_20740);
nand U22542 (N_22542,N_20066,N_21746);
nand U22543 (N_22543,N_20217,N_22186);
and U22544 (N_22544,N_21369,N_21374);
nand U22545 (N_22545,N_20802,N_20017);
and U22546 (N_22546,N_21474,N_20472);
xnor U22547 (N_22547,N_22120,N_20925);
nor U22548 (N_22548,N_22267,N_20878);
and U22549 (N_22549,N_22397,N_20732);
xor U22550 (N_22550,N_21873,N_21657);
nand U22551 (N_22551,N_20201,N_20028);
or U22552 (N_22552,N_20317,N_21834);
and U22553 (N_22553,N_22488,N_21735);
nand U22554 (N_22554,N_21496,N_21222);
nor U22555 (N_22555,N_20891,N_20273);
or U22556 (N_22556,N_20783,N_22076);
and U22557 (N_22557,N_21983,N_21191);
nand U22558 (N_22558,N_22034,N_22033);
and U22559 (N_22559,N_21170,N_20726);
and U22560 (N_22560,N_20069,N_21164);
xor U22561 (N_22561,N_21779,N_20654);
or U22562 (N_22562,N_20096,N_20136);
or U22563 (N_22563,N_22190,N_20083);
nor U22564 (N_22564,N_21418,N_21267);
xor U22565 (N_22565,N_21969,N_21557);
or U22566 (N_22566,N_21495,N_20377);
xor U22567 (N_22567,N_21090,N_21810);
nor U22568 (N_22568,N_22434,N_22043);
xor U22569 (N_22569,N_20652,N_20845);
xnor U22570 (N_22570,N_22418,N_20718);
or U22571 (N_22571,N_21607,N_22215);
and U22572 (N_22572,N_20686,N_21223);
nor U22573 (N_22573,N_21163,N_20443);
nor U22574 (N_22574,N_22378,N_20530);
nand U22575 (N_22575,N_22467,N_21679);
and U22576 (N_22576,N_20582,N_21526);
and U22577 (N_22577,N_22278,N_21275);
xnor U22578 (N_22578,N_20984,N_21710);
xnor U22579 (N_22579,N_21150,N_22200);
nand U22580 (N_22580,N_21539,N_22030);
xor U22581 (N_22581,N_21087,N_21531);
nand U22582 (N_22582,N_21225,N_22406);
nor U22583 (N_22583,N_21786,N_21322);
and U22584 (N_22584,N_21360,N_21477);
or U22585 (N_22585,N_21855,N_21524);
xnor U22586 (N_22586,N_20216,N_21832);
or U22587 (N_22587,N_21601,N_20424);
or U22588 (N_22588,N_21705,N_22170);
xor U22589 (N_22589,N_22045,N_20521);
nor U22590 (N_22590,N_20550,N_21475);
and U22591 (N_22591,N_20238,N_21022);
xnor U22592 (N_22592,N_20678,N_22414);
or U22593 (N_22593,N_22386,N_20806);
nor U22594 (N_22594,N_21835,N_21159);
nor U22595 (N_22595,N_21118,N_20329);
and U22596 (N_22596,N_22004,N_21939);
xnor U22597 (N_22597,N_21938,N_22317);
xnor U22598 (N_22598,N_21264,N_20270);
xnor U22599 (N_22599,N_20825,N_20497);
and U22600 (N_22600,N_22331,N_20246);
nor U22601 (N_22601,N_20460,N_21140);
or U22602 (N_22602,N_20994,N_21535);
and U22603 (N_22603,N_21291,N_21997);
nor U22604 (N_22604,N_22067,N_21181);
or U22605 (N_22605,N_22302,N_20901);
nand U22606 (N_22606,N_21842,N_21550);
or U22607 (N_22607,N_22460,N_21032);
nor U22608 (N_22608,N_21651,N_21500);
xnor U22609 (N_22609,N_21551,N_20015);
nand U22610 (N_22610,N_21213,N_20191);
and U22611 (N_22611,N_21650,N_22011);
and U22612 (N_22612,N_21902,N_22055);
nor U22613 (N_22613,N_20759,N_21094);
and U22614 (N_22614,N_22124,N_21035);
or U22615 (N_22615,N_22354,N_22191);
or U22616 (N_22616,N_20624,N_22337);
nor U22617 (N_22617,N_20008,N_22214);
nand U22618 (N_22618,N_22376,N_20151);
xnor U22619 (N_22619,N_22227,N_21238);
nand U22620 (N_22620,N_21209,N_21807);
nand U22621 (N_22621,N_22147,N_21904);
xnor U22622 (N_22622,N_21695,N_20417);
and U22623 (N_22623,N_20692,N_20762);
xor U22624 (N_22624,N_22493,N_21003);
xnor U22625 (N_22625,N_22371,N_20477);
and U22626 (N_22626,N_21525,N_20256);
xnor U22627 (N_22627,N_20785,N_20033);
and U22628 (N_22628,N_21463,N_22219);
and U22629 (N_22629,N_21077,N_20658);
nand U22630 (N_22630,N_20663,N_20404);
or U22631 (N_22631,N_20450,N_22187);
or U22632 (N_22632,N_20489,N_20573);
nand U22633 (N_22633,N_20282,N_22143);
and U22634 (N_22634,N_20533,N_21859);
nor U22635 (N_22635,N_20304,N_21093);
and U22636 (N_22636,N_21759,N_20865);
or U22637 (N_22637,N_20353,N_22204);
nand U22638 (N_22638,N_21881,N_20869);
xnor U22639 (N_22639,N_20570,N_20598);
and U22640 (N_22640,N_20222,N_21244);
or U22641 (N_22641,N_22396,N_21700);
or U22642 (N_22642,N_20586,N_21625);
nand U22643 (N_22643,N_21734,N_21990);
nor U22644 (N_22644,N_21335,N_21929);
nand U22645 (N_22645,N_21727,N_20449);
or U22646 (N_22646,N_21624,N_21951);
xnor U22647 (N_22647,N_21593,N_21189);
nand U22648 (N_22648,N_21465,N_21690);
nor U22649 (N_22649,N_21389,N_21719);
or U22650 (N_22650,N_21424,N_21194);
and U22651 (N_22651,N_20671,N_21652);
and U22652 (N_22652,N_21543,N_21200);
xor U22653 (N_22653,N_21613,N_21483);
nor U22654 (N_22654,N_21603,N_21754);
xor U22655 (N_22655,N_21005,N_21208);
and U22656 (N_22656,N_21177,N_21670);
and U22657 (N_22657,N_20911,N_20539);
and U22658 (N_22658,N_20073,N_22341);
nor U22659 (N_22659,N_20463,N_22091);
and U22660 (N_22660,N_22066,N_22348);
nand U22661 (N_22661,N_21425,N_21409);
nand U22662 (N_22662,N_20055,N_20837);
nor U22663 (N_22663,N_22151,N_20087);
nand U22664 (N_22664,N_21351,N_22401);
nand U22665 (N_22665,N_21545,N_21952);
xor U22666 (N_22666,N_21664,N_21080);
nand U22667 (N_22667,N_20668,N_20286);
and U22668 (N_22668,N_20542,N_21503);
nor U22669 (N_22669,N_22457,N_20041);
or U22670 (N_22670,N_20811,N_20940);
or U22671 (N_22671,N_22122,N_20336);
and U22672 (N_22672,N_22047,N_20132);
nor U22673 (N_22673,N_20193,N_22367);
and U22674 (N_22674,N_20187,N_21328);
nor U22675 (N_22675,N_21074,N_20647);
nand U22676 (N_22676,N_20511,N_22350);
or U22677 (N_22677,N_21822,N_20858);
nor U22678 (N_22678,N_21179,N_22330);
nand U22679 (N_22679,N_21675,N_21894);
nand U22680 (N_22680,N_20564,N_21386);
and U22681 (N_22681,N_21686,N_21202);
and U22682 (N_22682,N_21906,N_20829);
nand U22683 (N_22683,N_20293,N_21453);
nor U22684 (N_22684,N_20192,N_20676);
or U22685 (N_22685,N_20793,N_21081);
nand U22686 (N_22686,N_20574,N_21012);
or U22687 (N_22687,N_20791,N_21052);
or U22688 (N_22688,N_20607,N_20048);
and U22689 (N_22689,N_21050,N_20646);
xor U22690 (N_22690,N_20251,N_20895);
nor U22691 (N_22691,N_21507,N_22430);
and U22692 (N_22692,N_20296,N_20749);
nor U22693 (N_22693,N_22058,N_20495);
nand U22694 (N_22694,N_21854,N_22356);
or U22695 (N_22695,N_22440,N_20266);
nand U22696 (N_22696,N_20152,N_20632);
or U22697 (N_22697,N_20233,N_20504);
nor U22698 (N_22698,N_21796,N_20473);
xnor U22699 (N_22699,N_21533,N_22276);
or U22700 (N_22700,N_20758,N_22225);
or U22701 (N_22701,N_20139,N_22394);
xor U22702 (N_22702,N_21556,N_20125);
xnor U22703 (N_22703,N_22455,N_22182);
or U22704 (N_22704,N_21896,N_21368);
nand U22705 (N_22705,N_21914,N_22138);
and U22706 (N_22706,N_22026,N_20703);
nor U22707 (N_22707,N_21692,N_22099);
or U22708 (N_22708,N_20219,N_20985);
or U22709 (N_22709,N_21795,N_20926);
nand U22710 (N_22710,N_21586,N_20892);
or U22711 (N_22711,N_21790,N_22484);
nand U22712 (N_22712,N_21887,N_20403);
xor U22713 (N_22713,N_21907,N_21611);
or U22714 (N_22714,N_21402,N_21614);
or U22715 (N_22715,N_21174,N_22286);
or U22716 (N_22716,N_21433,N_20171);
xnor U22717 (N_22717,N_20428,N_22336);
and U22718 (N_22718,N_21427,N_21132);
nor U22719 (N_22719,N_22156,N_22145);
nor U22720 (N_22720,N_21660,N_20226);
or U22721 (N_22721,N_20198,N_21774);
and U22722 (N_22722,N_20934,N_21214);
nor U22723 (N_22723,N_20381,N_21247);
or U22724 (N_22724,N_20434,N_20374);
or U22725 (N_22725,N_21687,N_21055);
or U22726 (N_22726,N_20595,N_22315);
xnor U22727 (N_22727,N_21278,N_20103);
and U22728 (N_22728,N_21138,N_21918);
or U22729 (N_22729,N_20267,N_22471);
or U22730 (N_22730,N_21871,N_20669);
xor U22731 (N_22731,N_20370,N_20760);
nor U22732 (N_22732,N_20655,N_22256);
nand U22733 (N_22733,N_21644,N_20117);
or U22734 (N_22734,N_21930,N_20405);
xor U22735 (N_22735,N_20590,N_21852);
and U22736 (N_22736,N_20035,N_21813);
xor U22737 (N_22737,N_20834,N_21327);
xor U22738 (N_22738,N_20401,N_22079);
nor U22739 (N_22739,N_20684,N_21956);
or U22740 (N_22740,N_20735,N_22291);
or U22741 (N_22741,N_20730,N_21124);
nand U22742 (N_22742,N_21146,N_22253);
or U22743 (N_22743,N_22318,N_21337);
xor U22744 (N_22744,N_21827,N_20391);
xor U22745 (N_22745,N_20448,N_21714);
nand U22746 (N_22746,N_21765,N_22051);
and U22747 (N_22747,N_22353,N_20765);
or U22748 (N_22748,N_20700,N_20976);
or U22749 (N_22749,N_20998,N_20383);
xnor U22750 (N_22750,N_21302,N_21037);
and U22751 (N_22751,N_21621,N_21410);
nand U22752 (N_22752,N_21885,N_21296);
and U22753 (N_22753,N_21048,N_22183);
and U22754 (N_22754,N_21935,N_21580);
xor U22755 (N_22755,N_21818,N_22194);
and U22756 (N_22756,N_21339,N_22134);
or U22757 (N_22757,N_20387,N_20471);
nand U22758 (N_22758,N_20326,N_22259);
or U22759 (N_22759,N_20906,N_22313);
nor U22760 (N_22760,N_21421,N_20408);
xnor U22761 (N_22761,N_22333,N_21950);
and U22762 (N_22762,N_22114,N_20621);
or U22763 (N_22763,N_22305,N_21242);
and U22764 (N_22764,N_21770,N_20797);
and U22765 (N_22765,N_21515,N_22048);
or U22766 (N_22766,N_21884,N_21145);
nor U22767 (N_22767,N_20633,N_21009);
or U22768 (N_22768,N_21271,N_21555);
or U22769 (N_22769,N_22377,N_21349);
nand U22770 (N_22770,N_22111,N_20341);
nor U22771 (N_22771,N_20250,N_21583);
xor U22772 (N_22772,N_21441,N_20741);
nor U22773 (N_22773,N_22482,N_20629);
and U22774 (N_22774,N_20968,N_20996);
and U22775 (N_22775,N_20464,N_20160);
and U22776 (N_22776,N_21732,N_20138);
and U22777 (N_22777,N_20788,N_20531);
nor U22778 (N_22778,N_20922,N_22464);
nor U22779 (N_22779,N_21036,N_20955);
and U22780 (N_22780,N_20465,N_21733);
and U22781 (N_22781,N_20733,N_20884);
or U22782 (N_22782,N_20290,N_22322);
xnor U22783 (N_22783,N_20334,N_20864);
and U22784 (N_22784,N_20257,N_21762);
and U22785 (N_22785,N_20130,N_20437);
nor U22786 (N_22786,N_20927,N_21348);
nor U22787 (N_22787,N_22074,N_22444);
or U22788 (N_22788,N_20642,N_20862);
or U22789 (N_22789,N_22184,N_20322);
xnor U22790 (N_22790,N_22042,N_20232);
nor U22791 (N_22791,N_21091,N_22496);
and U22792 (N_22792,N_20094,N_21618);
nor U22793 (N_22793,N_20012,N_22448);
xnor U22794 (N_22794,N_20121,N_20062);
nor U22795 (N_22795,N_21253,N_21073);
nand U22796 (N_22796,N_21870,N_20079);
nor U22797 (N_22797,N_20795,N_22177);
nand U22798 (N_22798,N_20074,N_20611);
xnor U22799 (N_22799,N_20425,N_20679);
nor U22800 (N_22800,N_22153,N_22295);
xor U22801 (N_22801,N_20543,N_20185);
nor U22802 (N_22802,N_21212,N_21713);
nand U22803 (N_22803,N_21313,N_21512);
xor U22804 (N_22804,N_20128,N_21847);
nand U22805 (N_22805,N_22468,N_21711);
or U22806 (N_22806,N_21979,N_20992);
or U22807 (N_22807,N_20662,N_20681);
nor U22808 (N_22808,N_22157,N_22059);
nor U22809 (N_22809,N_20291,N_21317);
nor U22810 (N_22810,N_20122,N_20606);
or U22811 (N_22811,N_21173,N_20631);
nand U22812 (N_22812,N_21666,N_21234);
nor U22813 (N_22813,N_21219,N_20091);
or U22814 (N_22814,N_22491,N_22198);
or U22815 (N_22815,N_22346,N_21176);
xnor U22816 (N_22816,N_21298,N_21324);
nor U22817 (N_22817,N_22492,N_21113);
xnor U22818 (N_22818,N_21973,N_20274);
nand U22819 (N_22819,N_20053,N_22379);
and U22820 (N_22820,N_20565,N_20687);
xor U22821 (N_22821,N_20436,N_22311);
nand U22822 (N_22822,N_21261,N_22352);
nor U22823 (N_22823,N_21403,N_22069);
xor U22824 (N_22824,N_22274,N_20980);
and U22825 (N_22825,N_21038,N_22439);
or U22826 (N_22826,N_20106,N_20958);
xor U22827 (N_22827,N_20828,N_21537);
xor U22828 (N_22828,N_22438,N_20853);
or U22829 (N_22829,N_20311,N_21696);
nand U22830 (N_22830,N_21128,N_21588);
or U22831 (N_22831,N_21925,N_20966);
and U22832 (N_22832,N_21008,N_21673);
nand U22833 (N_22833,N_21851,N_22381);
nand U22834 (N_22834,N_20637,N_20279);
and U22835 (N_22835,N_20905,N_20615);
or U22836 (N_22836,N_20908,N_21928);
nand U22837 (N_22837,N_20883,N_21782);
nor U22838 (N_22838,N_20551,N_20609);
xor U22839 (N_22839,N_21344,N_20340);
nand U22840 (N_22840,N_20076,N_21186);
xor U22841 (N_22841,N_21706,N_20235);
nand U22842 (N_22842,N_20721,N_20812);
xnor U22843 (N_22843,N_20876,N_20656);
and U22844 (N_22844,N_20157,N_20777);
and U22845 (N_22845,N_21623,N_20422);
nand U22846 (N_22846,N_20145,N_22310);
xnor U22847 (N_22847,N_22155,N_21819);
xor U22848 (N_22848,N_21800,N_20593);
nand U22849 (N_22849,N_20474,N_21964);
nand U22850 (N_22850,N_21781,N_22044);
or U22851 (N_22851,N_21385,N_20162);
xor U22852 (N_22852,N_21263,N_21991);
nand U22853 (N_22853,N_21722,N_21046);
or U22854 (N_22854,N_21047,N_21338);
or U22855 (N_22855,N_22245,N_20362);
and U22856 (N_22856,N_21815,N_21875);
nor U22857 (N_22857,N_21070,N_21988);
and U22858 (N_22858,N_21099,N_21443);
or U22859 (N_22859,N_20969,N_21667);
nor U22860 (N_22860,N_20835,N_21789);
xor U22861 (N_22861,N_21578,N_21488);
and U22862 (N_22862,N_21629,N_20163);
xor U22863 (N_22863,N_21634,N_20255);
and U22864 (N_22864,N_22027,N_21858);
nor U22865 (N_22865,N_20854,N_22233);
xor U22866 (N_22866,N_20380,N_21872);
nand U22867 (N_22867,N_20115,N_22264);
xor U22868 (N_22868,N_20887,N_21609);
or U22869 (N_22869,N_20525,N_20209);
nand U22870 (N_22870,N_22080,N_20119);
nor U22871 (N_22871,N_21325,N_21104);
or U22872 (N_22872,N_21699,N_21289);
xor U22873 (N_22873,N_20359,N_21996);
xnor U22874 (N_22874,N_22266,N_22387);
and U22875 (N_22875,N_22097,N_21994);
xnor U22876 (N_22876,N_20042,N_20644);
and U22877 (N_22877,N_20603,N_20188);
xor U22878 (N_22878,N_21857,N_20572);
nand U22879 (N_22879,N_22445,N_20397);
xnor U22880 (N_22880,N_21769,N_22092);
nor U22881 (N_22881,N_21083,N_21282);
nand U22882 (N_22882,N_20566,N_21228);
and U22883 (N_22883,N_20554,N_20723);
xnor U22884 (N_22884,N_21948,N_20614);
and U22885 (N_22885,N_20517,N_22240);
and U22886 (N_22886,N_20709,N_21350);
and U22887 (N_22887,N_22073,N_22021);
nor U22888 (N_22888,N_21910,N_20870);
or U22889 (N_22889,N_21198,N_20761);
xnor U22890 (N_22890,N_20826,N_22018);
nor U22891 (N_22891,N_20046,N_21435);
or U22892 (N_22892,N_21879,N_21162);
and U22893 (N_22893,N_20358,N_20180);
nand U22894 (N_22894,N_20207,N_21026);
nor U22895 (N_22895,N_21715,N_21221);
xnor U22896 (N_22896,N_22297,N_20342);
or U22897 (N_22897,N_20886,N_21768);
nor U22898 (N_22898,N_20532,N_21466);
nor U22899 (N_22899,N_22241,N_21799);
or U22900 (N_22900,N_22083,N_20898);
nand U22901 (N_22901,N_20774,N_21509);
and U22902 (N_22902,N_22158,N_21197);
or U22903 (N_22903,N_20931,N_20365);
or U22904 (N_22904,N_20816,N_20492);
xor U22905 (N_22905,N_21482,N_20693);
nand U22906 (N_22906,N_20833,N_21230);
nand U22907 (N_22907,N_21201,N_22193);
and U22908 (N_22908,N_21256,N_20779);
nand U22909 (N_22909,N_21361,N_21334);
and U22910 (N_22910,N_21367,N_22181);
and U22911 (N_22911,N_21971,N_21404);
nand U22912 (N_22912,N_21000,N_22025);
and U22913 (N_22913,N_20084,N_20452);
and U22914 (N_22914,N_20275,N_22425);
nor U22915 (N_22915,N_21522,N_22049);
nand U22916 (N_22916,N_20600,N_20831);
nand U22917 (N_22917,N_21916,N_21773);
and U22918 (N_22918,N_20610,N_22231);
or U22919 (N_22919,N_21249,N_21147);
nand U22920 (N_22920,N_21476,N_21508);
nand U22921 (N_22921,N_20373,N_20879);
nand U22922 (N_22922,N_20454,N_21571);
nor U22923 (N_22923,N_21582,N_20722);
xnor U22924 (N_22924,N_20089,N_20004);
nand U22925 (N_22925,N_21183,N_22068);
or U22926 (N_22926,N_20240,N_20203);
or U22927 (N_22927,N_21137,N_22405);
and U22928 (N_22928,N_22168,N_20839);
or U22929 (N_22929,N_21144,N_21478);
xor U22930 (N_22930,N_20178,N_21382);
or U22931 (N_22931,N_21490,N_21702);
or U22932 (N_22932,N_20634,N_21469);
nor U22933 (N_22933,N_21210,N_22481);
nor U22934 (N_22934,N_21061,N_20769);
nand U22935 (N_22935,N_21772,N_20348);
and U22936 (N_22936,N_20278,N_21442);
or U22937 (N_22937,N_20483,N_21756);
or U22938 (N_22938,N_22016,N_22334);
or U22939 (N_22939,N_20061,N_21266);
and U22940 (N_22940,N_20713,N_22209);
nor U22941 (N_22941,N_21965,N_20248);
or U22942 (N_22942,N_20426,N_22262);
xnor U22943 (N_22943,N_22343,N_21764);
or U22944 (N_22944,N_22273,N_20951);
or U22945 (N_22945,N_22161,N_22062);
xnor U22946 (N_22946,N_22417,N_22179);
and U22947 (N_22947,N_20844,N_21913);
and U22948 (N_22948,N_22232,N_21109);
or U22949 (N_22949,N_20071,N_20848);
and U22950 (N_22950,N_22008,N_21027);
xor U22951 (N_22951,N_20714,N_21241);
nor U22952 (N_22952,N_21518,N_21824);
xnor U22953 (N_22953,N_22281,N_21065);
nor U22954 (N_22954,N_21749,N_22171);
or U22955 (N_22955,N_20349,N_21649);
or U22956 (N_22956,N_22402,N_21584);
nand U22957 (N_22957,N_22071,N_20746);
nand U22958 (N_22958,N_21744,N_20031);
xnor U22959 (N_22959,N_22441,N_20345);
or U22960 (N_22960,N_22100,N_21287);
xnor U22961 (N_22961,N_21236,N_20253);
or U22962 (N_22962,N_20337,N_21028);
nor U22963 (N_22963,N_20081,N_20667);
nor U22964 (N_22964,N_21257,N_20505);
nor U22965 (N_22965,N_21568,N_21577);
xnor U22966 (N_22966,N_20970,N_22329);
and U22967 (N_22967,N_22244,N_21078);
nand U22968 (N_22968,N_20493,N_21320);
nand U22969 (N_22969,N_21787,N_21459);
xnor U22970 (N_22970,N_21076,N_21122);
nand U22971 (N_22971,N_20688,N_21130);
or U22972 (N_22972,N_21057,N_20503);
and U22973 (N_22973,N_21724,N_20418);
nor U22974 (N_22974,N_20939,N_21510);
xor U22975 (N_22975,N_22222,N_20153);
or U22976 (N_22976,N_20455,N_20189);
and U22977 (N_22977,N_20195,N_21610);
and U22978 (N_22978,N_20221,N_21457);
nand U22979 (N_22979,N_20419,N_21152);
and U22980 (N_22980,N_21203,N_20241);
xor U22981 (N_22981,N_20242,N_21079);
nand U22982 (N_22982,N_20894,N_20830);
nor U22983 (N_22983,N_22165,N_20569);
xor U22984 (N_22984,N_21279,N_21922);
nand U22985 (N_22985,N_21691,N_21534);
nand U22986 (N_22986,N_21101,N_21620);
xor U22987 (N_22987,N_22197,N_22096);
xor U22988 (N_22988,N_20528,N_21920);
xor U22989 (N_22989,N_21863,N_21276);
or U22990 (N_22990,N_21541,N_21372);
or U22991 (N_22991,N_21297,N_21010);
xor U22992 (N_22992,N_20330,N_22054);
xor U22993 (N_22993,N_21269,N_21089);
nand U22994 (N_22994,N_21393,N_20040);
nor U22995 (N_22995,N_20617,N_21729);
nand U22996 (N_22996,N_20881,N_22131);
nand U22997 (N_22997,N_21636,N_20952);
or U22998 (N_22998,N_22490,N_21559);
or U22999 (N_22999,N_21294,N_20010);
or U23000 (N_23000,N_21172,N_21292);
or U23001 (N_23001,N_20095,N_20284);
xnor U23002 (N_23002,N_21473,N_21565);
nand U23003 (N_23003,N_21067,N_21844);
and U23004 (N_23004,N_22442,N_21436);
nor U23005 (N_23005,N_21116,N_22082);
nand U23006 (N_23006,N_21516,N_21671);
and U23007 (N_23007,N_22252,N_20431);
or U23008 (N_23008,N_21345,N_20302);
xnor U23009 (N_23009,N_20974,N_22247);
xnor U23010 (N_23010,N_20989,N_21575);
xor U23011 (N_23011,N_21487,N_20410);
nand U23012 (N_23012,N_22413,N_22172);
xnor U23013 (N_23013,N_21086,N_20456);
nor U23014 (N_23014,N_21936,N_20982);
or U23015 (N_23015,N_21750,N_20776);
and U23016 (N_23016,N_20928,N_22189);
or U23017 (N_23017,N_21023,N_21255);
and U23018 (N_23018,N_21984,N_20548);
and U23019 (N_23019,N_22110,N_22087);
xor U23020 (N_23020,N_20491,N_22314);
xnor U23021 (N_23021,N_22038,N_21188);
nor U23022 (N_23022,N_21272,N_21448);
or U23023 (N_23023,N_22095,N_20309);
xor U23024 (N_23024,N_20043,N_21184);
and U23025 (N_23025,N_20680,N_21798);
nand U23026 (N_23026,N_21654,N_20737);
nor U23027 (N_23027,N_21802,N_22388);
and U23028 (N_23028,N_21347,N_22357);
nor U23029 (N_23029,N_21942,N_20796);
xnor U23030 (N_23030,N_20281,N_21663);
xnor U23031 (N_23031,N_20836,N_20352);
nor U23032 (N_23032,N_20011,N_21968);
nand U23033 (N_23033,N_21723,N_21303);
and U23034 (N_23034,N_20446,N_20482);
xor U23035 (N_23035,N_21899,N_21187);
xnor U23036 (N_23036,N_20077,N_21370);
nor U23037 (N_23037,N_20001,N_21995);
nor U23038 (N_23038,N_22001,N_22384);
nor U23039 (N_23039,N_20556,N_21446);
xor U23040 (N_23040,N_21830,N_20781);
xor U23041 (N_23041,N_21103,N_22050);
or U23042 (N_23042,N_21977,N_20792);
nand U23043 (N_23043,N_20239,N_21185);
nor U23044 (N_23044,N_20224,N_20327);
nand U23045 (N_23045,N_21932,N_21604);
and U23046 (N_23046,N_20102,N_20627);
xor U23047 (N_23047,N_20075,N_20972);
or U23048 (N_23048,N_21600,N_20960);
or U23049 (N_23049,N_21293,N_21954);
or U23050 (N_23050,N_20468,N_20488);
xor U23051 (N_23051,N_21105,N_22462);
nor U23052 (N_23052,N_20995,N_22133);
xor U23053 (N_23053,N_22358,N_22238);
nand U23054 (N_23054,N_22185,N_21001);
and U23055 (N_23055,N_21030,N_20440);
xnor U23056 (N_23056,N_21985,N_22152);
xnor U23057 (N_23057,N_20333,N_20480);
nand U23058 (N_23058,N_20752,N_22202);
nor U23059 (N_23059,N_21882,N_20639);
nand U23060 (N_23060,N_21299,N_22323);
and U23061 (N_23061,N_20963,N_20457);
xnor U23062 (N_23062,N_21353,N_22070);
nand U23063 (N_23063,N_20997,N_21332);
nor U23064 (N_23064,N_20120,N_20832);
or U23065 (N_23065,N_21839,N_20840);
nor U23066 (N_23066,N_22173,N_20100);
or U23067 (N_23067,N_22303,N_21044);
nor U23068 (N_23068,N_21814,N_22195);
nor U23069 (N_23069,N_20524,N_21740);
or U23070 (N_23070,N_21725,N_21590);
nand U23071 (N_23071,N_20236,N_21751);
or U23072 (N_23072,N_20872,N_20023);
and U23073 (N_23073,N_21743,N_21574);
nor U23074 (N_23074,N_21888,N_20137);
or U23075 (N_23075,N_22287,N_20947);
or U23076 (N_23076,N_21972,N_21112);
or U23077 (N_23077,N_20786,N_20414);
nor U23078 (N_23078,N_21029,N_21069);
nand U23079 (N_23079,N_20086,N_22399);
or U23080 (N_23080,N_22280,N_20479);
xor U23081 (N_23081,N_21396,N_21383);
xnor U23082 (N_23082,N_20312,N_20805);
nand U23083 (N_23083,N_21923,N_22012);
nand U23084 (N_23084,N_20824,N_22013);
nand U23085 (N_23085,N_20127,N_21376);
and U23086 (N_23086,N_21045,N_22312);
nand U23087 (N_23087,N_21489,N_22324);
nand U23088 (N_23088,N_20375,N_22239);
xor U23089 (N_23089,N_21890,N_20131);
nand U23090 (N_23090,N_22056,N_20973);
nor U23091 (N_23091,N_21521,N_20818);
nor U23092 (N_23092,N_20451,N_21561);
nor U23093 (N_23093,N_22307,N_20344);
or U23094 (N_23094,N_22077,N_21391);
and U23095 (N_23095,N_22359,N_21680);
xnor U23096 (N_23096,N_21398,N_22258);
xnor U23097 (N_23097,N_21919,N_22023);
nor U23098 (N_23098,N_20104,N_21615);
xor U23099 (N_23099,N_20182,N_21633);
nand U23100 (N_23100,N_20357,N_20315);
nor U23101 (N_23101,N_20490,N_22308);
nand U23102 (N_23102,N_20179,N_22089);
nor U23103 (N_23103,N_21547,N_20164);
and U23104 (N_23104,N_22366,N_21326);
xor U23105 (N_23105,N_20838,N_21237);
xnor U23106 (N_23106,N_21021,N_21218);
nor U23107 (N_23107,N_20738,N_20975);
nand U23108 (N_23108,N_21817,N_20500);
and U23109 (N_23109,N_22180,N_21429);
or U23110 (N_23110,N_20961,N_20124);
and U23111 (N_23111,N_20245,N_21755);
and U23112 (N_23112,N_21420,N_20948);
xnor U23113 (N_23113,N_21897,N_21004);
or U23114 (N_23114,N_21133,N_22029);
xnor U23115 (N_23115,N_21564,N_20949);
xnor U23116 (N_23116,N_21801,N_20946);
nand U23117 (N_23117,N_20843,N_21974);
and U23118 (N_23118,N_22426,N_20575);
xnor U23119 (N_23119,N_21273,N_22166);
xor U23120 (N_23120,N_20935,N_21542);
nand U23121 (N_23121,N_22349,N_21462);
xnor U23122 (N_23122,N_20300,N_20763);
or U23123 (N_23123,N_22470,N_21379);
nand U23124 (N_23124,N_21363,N_22345);
or U23125 (N_23125,N_22389,N_21576);
xnor U23126 (N_23126,N_20165,N_21100);
or U23127 (N_23127,N_22205,N_20476);
nor U23128 (N_23128,N_20767,N_20599);
xnor U23129 (N_23129,N_21841,N_21643);
and U23130 (N_23130,N_21136,N_20072);
xnor U23131 (N_23131,N_21157,N_22279);
xor U23132 (N_23132,N_20957,N_22107);
nand U23133 (N_23133,N_20361,N_21794);
xnor U23134 (N_23134,N_20977,N_21158);
nand U23135 (N_23135,N_21454,N_20372);
nand U23136 (N_23136,N_20690,N_20594);
nor U23137 (N_23137,N_21431,N_21926);
xor U23138 (N_23138,N_20399,N_22309);
or U23139 (N_23139,N_20196,N_20716);
xnor U23140 (N_23140,N_21097,N_21437);
or U23141 (N_23141,N_21430,N_21934);
and U23142 (N_23142,N_20335,N_20343);
and U23143 (N_23143,N_22487,N_21560);
xnor U23144 (N_23144,N_21108,N_21662);
and U23145 (N_23145,N_22459,N_21783);
nand U23146 (N_23146,N_22347,N_21054);
and U23147 (N_23147,N_22395,N_20308);
xor U23148 (N_23148,N_20218,N_21869);
nor U23149 (N_23149,N_20850,N_20673);
or U23150 (N_23150,N_21387,N_22424);
xor U23151 (N_23151,N_22458,N_20285);
xnor U23152 (N_23152,N_20698,N_20707);
xnor U23153 (N_23153,N_20323,N_20540);
nand U23154 (N_23154,N_21893,N_22419);
nor U23155 (N_23155,N_22411,N_22255);
or U23156 (N_23156,N_20766,N_21793);
nand U23157 (N_23157,N_21394,N_22431);
and U23158 (N_23158,N_21479,N_22409);
nor U23159 (N_23159,N_20964,N_21707);
nand U23160 (N_23160,N_20620,N_20156);
or U23161 (N_23161,N_20823,N_20394);
nand U23162 (N_23162,N_21321,N_20366);
nand U23163 (N_23163,N_20260,N_21642);
xor U23164 (N_23164,N_20641,N_20186);
nor U23165 (N_23165,N_21778,N_21284);
and U23166 (N_23166,N_22125,N_21880);
nor U23167 (N_23167,N_20301,N_21329);
nor U23168 (N_23168,N_20501,N_21684);
nand U23169 (N_23169,N_21989,N_21286);
or U23170 (N_23170,N_21791,N_20133);
nand U23171 (N_23171,N_21596,N_21821);
or U23172 (N_23172,N_20389,N_21622);
xor U23173 (N_23173,N_20780,N_21017);
and U23174 (N_23174,N_22485,N_20636);
and U23175 (N_23175,N_20400,N_21129);
xor U23176 (N_23176,N_22463,N_20181);
nor U23177 (N_23177,N_20407,N_22020);
or U23178 (N_23178,N_20885,N_21270);
and U23179 (N_23179,N_22098,N_20683);
and U23180 (N_23180,N_21502,N_20332);
and U23181 (N_23181,N_21504,N_21912);
nand U23182 (N_23182,N_21532,N_20204);
xnor U23183 (N_23183,N_21826,N_20507);
nand U23184 (N_23184,N_22223,N_20470);
nor U23185 (N_23185,N_22285,N_20527);
or U23186 (N_23186,N_20847,N_21944);
or U23187 (N_23187,N_20863,N_21788);
nand U23188 (N_23188,N_22294,N_21456);
nand U23189 (N_23189,N_20981,N_20710);
nor U23190 (N_23190,N_21196,N_21468);
or U23191 (N_23191,N_20388,N_22392);
and U23192 (N_23192,N_21068,N_20415);
and U23193 (N_23193,N_22041,N_20168);
and U23194 (N_23194,N_22422,N_22497);
and U23195 (N_23195,N_21889,N_20049);
xnor U23196 (N_23196,N_20328,N_22002);
xnor U23197 (N_23197,N_21876,N_20601);
or U23198 (N_23198,N_20549,N_21232);
and U23199 (N_23199,N_21484,N_20092);
or U23200 (N_23200,N_20080,N_21281);
and U23201 (N_23201,N_21536,N_22052);
nor U23202 (N_23202,N_20613,N_22254);
or U23203 (N_23203,N_21761,N_21064);
or U23204 (N_23204,N_21986,N_20305);
and U23205 (N_23205,N_20956,N_21943);
nor U23206 (N_23206,N_20051,N_20258);
xnor U23207 (N_23207,N_20044,N_20356);
xor U23208 (N_23208,N_20496,N_20696);
or U23209 (N_23209,N_21992,N_21540);
nand U23210 (N_23210,N_22275,N_20129);
xnor U23211 (N_23211,N_21121,N_21428);
or U23212 (N_23212,N_22249,N_22351);
or U23213 (N_23213,N_22250,N_22217);
nor U23214 (N_23214,N_20553,N_21730);
and U23215 (N_23215,N_20744,N_20666);
xnor U23216 (N_23216,N_20154,N_22075);
nand U23217 (N_23217,N_20699,N_21892);
xnor U23218 (N_23218,N_21742,N_20113);
xnor U23219 (N_23219,N_21250,N_21288);
xnor U23220 (N_23220,N_21579,N_21165);
xor U23221 (N_23221,N_21688,N_21224);
and U23222 (N_23222,N_21592,N_21408);
xor U23223 (N_23223,N_21911,N_21594);
and U23224 (N_23224,N_21597,N_20640);
and U23225 (N_23225,N_21259,N_22364);
xnor U23226 (N_23226,N_21280,N_22117);
xnor U23227 (N_23227,N_22160,N_22270);
or U23228 (N_23228,N_21406,N_21235);
nand U23229 (N_23229,N_20914,N_20205);
and U23230 (N_23230,N_20430,N_20800);
xor U23231 (N_23231,N_21848,N_22226);
and U23232 (N_23232,N_21831,N_21685);
xor U23233 (N_23233,N_21767,N_20576);
and U23234 (N_23234,N_22398,N_21432);
xor U23235 (N_23235,N_21451,N_20445);
nor U23236 (N_23236,N_22289,N_22220);
xnor U23237 (N_23237,N_20938,N_20577);
nand U23238 (N_23238,N_20808,N_20754);
and U23239 (N_23239,N_22228,N_20541);
nor U23240 (N_23240,N_20499,N_22235);
and U23241 (N_23241,N_20849,N_22140);
nor U23242 (N_23242,N_21683,N_20421);
xor U23243 (N_23243,N_20494,N_20265);
or U23244 (N_23244,N_22000,N_21548);
and U23245 (N_23245,N_20225,N_20288);
and U23246 (N_23246,N_20261,N_21681);
xor U23247 (N_23247,N_20314,N_21708);
nor U23248 (N_23248,N_22282,N_21737);
nand U23249 (N_23249,N_21970,N_20324);
nor U23250 (N_23250,N_22453,N_21694);
nand U23251 (N_23251,N_22306,N_20243);
nand U23252 (N_23252,N_21135,N_20546);
nor U23253 (N_23253,N_21566,N_20354);
nor U23254 (N_23254,N_21311,N_20280);
xor U23255 (N_23255,N_20584,N_20986);
and U23256 (N_23256,N_21647,N_20579);
xnor U23257 (N_23257,N_21498,N_21677);
xor U23258 (N_23258,N_21307,N_21240);
and U23259 (N_23259,N_22473,N_22298);
nor U23260 (N_23260,N_20999,N_20856);
nor U23261 (N_23261,N_21612,N_20478);
and U23262 (N_23262,N_20773,N_21567);
nor U23263 (N_23263,N_20896,N_21423);
or U23264 (N_23264,N_20561,N_21336);
nand U23265 (N_23265,N_22036,N_22210);
nand U23266 (N_23266,N_20866,N_20875);
and U23267 (N_23267,N_22480,N_21331);
nand U23268 (N_23268,N_21955,N_21908);
nor U23269 (N_23269,N_20237,N_22407);
and U23270 (N_23270,N_20029,N_21066);
xnor U23271 (N_23271,N_20672,N_21780);
and U23272 (N_23272,N_20558,N_20857);
nor U23273 (N_23273,N_20888,N_20439);
xor U23274 (N_23274,N_21314,N_21874);
xor U23275 (N_23275,N_20190,N_21439);
nand U23276 (N_23276,N_20799,N_20817);
xor U23277 (N_23277,N_21602,N_21572);
nor U23278 (N_23278,N_20842,N_20923);
xnor U23279 (N_23279,N_21812,N_20583);
nor U23280 (N_23280,N_20303,N_20522);
or U23281 (N_23281,N_20320,N_22251);
or U23282 (N_23282,N_20529,N_21248);
xor U23283 (N_23283,N_22391,N_20319);
nand U23284 (N_23284,N_22208,N_21709);
or U23285 (N_23285,N_21668,N_21246);
xnor U23286 (N_23286,N_20535,N_20259);
nor U23287 (N_23287,N_21356,N_22115);
nor U23288 (N_23288,N_20339,N_21033);
nand U23289 (N_23289,N_21739,N_22475);
xor U23290 (N_23290,N_21458,N_21501);
or U23291 (N_23291,N_20648,N_21352);
nand U23292 (N_23292,N_20367,N_20623);
xnor U23293 (N_23293,N_21720,N_22212);
or U23294 (N_23294,N_20653,N_20351);
nor U23295 (N_23295,N_20429,N_21569);
xnor U23296 (N_23296,N_21310,N_21513);
and U23297 (N_23297,N_20088,N_22498);
or U23298 (N_23298,N_21511,N_20562);
xnor U23299 (N_23299,N_21626,N_21399);
and U23300 (N_23300,N_21154,N_20299);
nand U23301 (N_23301,N_20009,N_20537);
nor U23302 (N_23302,N_22201,N_21726);
nand U23303 (N_23303,N_20743,N_21400);
and U23304 (N_23304,N_20262,N_20210);
and U23305 (N_23305,N_20295,N_21422);
or U23306 (N_23306,N_21031,N_21562);
xor U23307 (N_23307,N_22009,N_22372);
nor U23308 (N_23308,N_21156,N_21803);
and U23309 (N_23309,N_21886,N_21006);
nor U23310 (N_23310,N_22447,N_20036);
xor U23311 (N_23311,N_21845,N_20591);
or U23312 (N_23312,N_21946,N_21552);
and U23313 (N_23313,N_21371,N_22094);
nand U23314 (N_23314,N_20991,N_20413);
nor U23315 (N_23315,N_20416,N_20790);
nand U23316 (N_23316,N_21239,N_21776);
xor U23317 (N_23317,N_20536,N_21606);
xnor U23318 (N_23318,N_21318,N_22014);
xor U23319 (N_23319,N_20244,N_20719);
xor U23320 (N_23320,N_20432,N_22320);
nor U23321 (N_23321,N_21499,N_22218);
and U23322 (N_23322,N_22236,N_21085);
or U23323 (N_23323,N_20200,N_21254);
xnor U23324 (N_23324,N_21689,N_21811);
or U23325 (N_23325,N_21354,N_21229);
xnor U23326 (N_23326,N_21252,N_20630);
nand U23327 (N_23327,N_22237,N_22335);
xor U23328 (N_23328,N_21849,N_20717);
nor U23329 (N_23329,N_20231,N_21619);
and U23330 (N_23330,N_20567,N_21804);
and U23331 (N_23331,N_21850,N_22380);
xor U23332 (N_23332,N_20682,N_22164);
xnor U23333 (N_23333,N_22476,N_20484);
or U23334 (N_23334,N_21127,N_20930);
xnor U23335 (N_23335,N_21205,N_20212);
xor U23336 (N_23336,N_20987,N_20943);
xnor U23337 (N_23337,N_20228,N_20099);
xnor U23338 (N_23338,N_22242,N_20386);
or U23339 (N_23339,N_22472,N_20045);
or U23340 (N_23340,N_20962,N_20037);
nand U23341 (N_23341,N_20264,N_22088);
nor U23342 (N_23342,N_20027,N_21412);
nor U23343 (N_23343,N_21570,N_22271);
nor U23344 (N_23344,N_21963,N_22410);
nor U23345 (N_23345,N_21530,N_20701);
nor U23346 (N_23346,N_20466,N_20635);
or U23347 (N_23347,N_21365,N_21792);
or U23348 (N_23348,N_20727,N_20252);
nor U23349 (N_23349,N_20002,N_21160);
nand U23350 (N_23350,N_21110,N_22369);
xor U23351 (N_23351,N_21837,N_22149);
nor U23352 (N_23352,N_21960,N_22301);
and U23353 (N_23353,N_22065,N_20271);
xor U23354 (N_23354,N_21877,N_21366);
xor U23355 (N_23355,N_20907,N_21285);
or U23356 (N_23356,N_21283,N_21816);
or U23357 (N_23357,N_20254,N_21505);
or U23358 (N_23358,N_20675,N_22283);
and U23359 (N_23359,N_21672,N_22006);
or U23360 (N_23360,N_20670,N_22450);
xnor U23361 (N_23361,N_20070,N_21357);
and U23362 (N_23362,N_20039,N_20770);
or U23363 (N_23363,N_20846,N_20768);
and U23364 (N_23364,N_20728,N_20979);
nor U23365 (N_23365,N_21766,N_22207);
xnor U23366 (N_23366,N_21415,N_21966);
and U23367 (N_23367,N_20959,N_20032);
nor U23368 (N_23368,N_22456,N_20360);
nor U23369 (N_23369,N_21151,N_20433);
xor U23370 (N_23370,N_21797,N_20060);
xnor U23371 (N_23371,N_20148,N_21538);
or U23372 (N_23372,N_22499,N_22429);
and U23373 (N_23373,N_22408,N_22300);
nand U23374 (N_23374,N_21362,N_22035);
nor U23375 (N_23375,N_22474,N_21823);
xor U23376 (N_23376,N_21616,N_22427);
nand U23377 (N_23377,N_21120,N_21669);
nor U23378 (N_23378,N_20538,N_21405);
and U23379 (N_23379,N_21661,N_21340);
and U23380 (N_23380,N_20392,N_22229);
or U23381 (N_23381,N_21075,N_20487);
nand U23382 (N_23382,N_22040,N_20820);
nand U23383 (N_23383,N_21865,N_20988);
xnor U23384 (N_23384,N_22230,N_21485);
and U23385 (N_23385,N_22269,N_22084);
and U23386 (N_23386,N_21931,N_20110);
xnor U23387 (N_23387,N_22469,N_22154);
nand U23388 (N_23388,N_22248,N_20936);
and U23389 (N_23389,N_20518,N_22316);
xnor U23390 (N_23390,N_22435,N_20398);
and U23391 (N_23391,N_22130,N_20174);
or U23392 (N_23392,N_21728,N_22174);
or U23393 (N_23393,N_20734,N_20297);
xnor U23394 (N_23394,N_22102,N_20890);
and U23395 (N_23395,N_20702,N_21295);
xor U23396 (N_23396,N_22113,N_20057);
and U23397 (N_23397,N_20882,N_22081);
or U23398 (N_23398,N_20161,N_21748);
nor U23399 (N_23399,N_20462,N_21315);
xnor U23400 (N_23400,N_20065,N_22368);
xnor U23401 (N_23401,N_20007,N_21268);
nand U23402 (N_23402,N_21829,N_20321);
nand U23403 (N_23403,N_21450,N_21062);
nor U23404 (N_23404,N_20813,N_20054);
xnor U23405 (N_23405,N_20141,N_22086);
or U23406 (N_23406,N_20919,N_21712);
nand U23407 (N_23407,N_21937,N_20547);
nand U23408 (N_23408,N_20932,N_20396);
nand U23409 (N_23409,N_20112,N_21180);
xnor U23410 (N_23410,N_21546,N_21378);
or U23411 (N_23411,N_21115,N_21967);
nor U23412 (N_23412,N_21840,N_20363);
and U23413 (N_23413,N_22452,N_22175);
xor U23414 (N_23414,N_22403,N_20116);
or U23415 (N_23415,N_21617,N_21895);
and U23416 (N_23416,N_22039,N_20904);
or U23417 (N_23417,N_22137,N_21809);
or U23418 (N_23418,N_21736,N_21072);
nor U23419 (N_23419,N_21155,N_22159);
and U23420 (N_23420,N_20880,N_21388);
nor U23421 (N_23421,N_21581,N_20909);
or U23422 (N_23422,N_20005,N_20801);
or U23423 (N_23423,N_20563,N_21226);
nand U23424 (N_23424,N_20705,N_20755);
nor U23425 (N_23425,N_22465,N_22375);
nor U23426 (N_23426,N_21051,N_20841);
xor U23427 (N_23427,N_21039,N_20971);
and U23428 (N_23428,N_21598,N_20506);
nor U23429 (N_23429,N_22478,N_21013);
nand U23430 (N_23430,N_22135,N_22015);
and U23431 (N_23431,N_21646,N_21549);
nor U23432 (N_23432,N_21757,N_22383);
nand U23433 (N_23433,N_21674,N_21745);
xnor U23434 (N_23434,N_22443,N_22265);
xnor U23435 (N_23435,N_20384,N_21492);
xor U23436 (N_23436,N_20860,N_21697);
xnor U23437 (N_23437,N_20787,N_21864);
nor U23438 (N_23438,N_21589,N_21976);
or U23439 (N_23439,N_21375,N_22385);
nand U23440 (N_23440,N_20019,N_22163);
nand U23441 (N_23441,N_20064,N_20109);
or U23442 (N_23442,N_21341,N_20438);
nor U23443 (N_23443,N_20249,N_22393);
nand U23444 (N_23444,N_21631,N_20822);
nor U23445 (N_23445,N_20798,N_20058);
or U23446 (N_23446,N_20022,N_21878);
or U23447 (N_23447,N_21245,N_21656);
or U23448 (N_23448,N_20871,N_21460);
nor U23449 (N_23449,N_20025,N_20877);
and U23450 (N_23450,N_21472,N_20578);
or U23451 (N_23451,N_20661,N_21843);
xnor U23452 (N_23452,N_21207,N_20933);
and U23453 (N_23453,N_21752,N_21957);
nand U23454 (N_23454,N_21805,N_20706);
nor U23455 (N_23455,N_20444,N_20937);
nor U23456 (N_23456,N_21941,N_20967);
and U23457 (N_23457,N_21407,N_20123);
nor U23458 (N_23458,N_21481,N_22342);
xor U23459 (N_23459,N_20807,N_21640);
or U23460 (N_23460,N_22057,N_20147);
xor U23461 (N_23461,N_20508,N_22109);
and U23462 (N_23462,N_20368,N_20485);
and U23463 (N_23463,N_21193,N_21330);
nor U23464 (N_23464,N_21416,N_20177);
or U23465 (N_23465,N_20819,N_21519);
nor U23466 (N_23466,N_22112,N_20915);
or U23467 (N_23467,N_20000,N_20552);
xor U23468 (N_23468,N_21924,N_21909);
xor U23469 (N_23469,N_20442,N_21227);
xor U23470 (N_23470,N_22483,N_20229);
nor U23471 (N_23471,N_21486,N_20461);
nand U23472 (N_23472,N_22003,N_21082);
nor U23473 (N_23473,N_22325,N_22268);
and U23474 (N_23474,N_20376,N_20622);
or U23475 (N_23475,N_20659,N_20736);
xor U23476 (N_23476,N_21216,N_21953);
and U23477 (N_23477,N_20134,N_20664);
or U23478 (N_23478,N_20910,N_22420);
and U23479 (N_23479,N_21049,N_22451);
nor U23480 (N_23480,N_22211,N_21856);
or U23481 (N_23481,N_20592,N_21753);
or U23482 (N_23482,N_22449,N_21698);
nor U23483 (N_23483,N_22093,N_20953);
nor U23484 (N_23484,N_20516,N_21771);
and U23485 (N_23485,N_21461,N_21471);
nand U23486 (N_23486,N_20412,N_20874);
xnor U23487 (N_23487,N_22365,N_20649);
nor U23488 (N_23488,N_21220,N_22321);
and U23489 (N_23489,N_20954,N_22178);
nor U23490 (N_23490,N_20942,N_21862);
and U23491 (N_23491,N_20745,N_21544);
nor U23492 (N_23492,N_20917,N_20873);
xor U23493 (N_23493,N_21088,N_20287);
nor U23494 (N_23494,N_22339,N_21861);
nor U23495 (N_23495,N_21384,N_21820);
xor U23496 (N_23496,N_20523,N_20742);
nand U23497 (N_23497,N_20739,N_21141);
xnor U23498 (N_23498,N_22400,N_22213);
or U23499 (N_23499,N_20512,N_22446);
xor U23500 (N_23500,N_21860,N_20784);
and U23501 (N_23501,N_21961,N_20338);
nand U23502 (N_23502,N_21381,N_20021);
xnor U23503 (N_23503,N_21444,N_20292);
xor U23504 (N_23504,N_22319,N_20026);
and U23505 (N_23505,N_22326,N_21445);
nand U23506 (N_23506,N_21828,N_20068);
nand U23507 (N_23507,N_22167,N_20211);
nand U23508 (N_23508,N_20213,N_22362);
xor U23509 (N_23509,N_20608,N_20660);
nor U23510 (N_23510,N_20711,N_21265);
nor U23511 (N_23511,N_21262,N_20775);
xnor U23512 (N_23512,N_20097,N_21682);
and U23513 (N_23513,N_20167,N_22132);
or U23514 (N_23514,N_20018,N_21171);
nand U23515 (N_23515,N_22141,N_20889);
or U23516 (N_23516,N_21747,N_22260);
xnor U23517 (N_23517,N_20899,N_21199);
or U23518 (N_23518,N_21233,N_20913);
nor U23519 (N_23519,N_20126,N_22216);
and U23520 (N_23520,N_20650,N_21573);
xor U23521 (N_23521,N_20379,N_21731);
or U23522 (N_23522,N_20289,N_21364);
and U23523 (N_23523,N_21015,N_20897);
and U23524 (N_23524,N_21417,N_22338);
nand U23525 (N_23525,N_22421,N_20588);
or U23526 (N_23526,N_22390,N_21659);
xnor U23527 (N_23527,N_21494,N_21758);
or U23528 (N_23528,N_22373,N_20047);
nand U23529 (N_23529,N_21785,N_20427);
or U23530 (N_23530,N_21464,N_20194);
nand U23531 (N_23531,N_21853,N_20090);
nor U23532 (N_23532,N_21470,N_21016);
nand U23533 (N_23533,N_21591,N_21628);
nor U23534 (N_23534,N_21517,N_22433);
or U23535 (N_23535,N_21959,N_22261);
nand U23536 (N_23536,N_22284,N_21401);
and U23537 (N_23537,N_22061,N_21678);
and U23538 (N_23538,N_22272,N_20006);
and U23539 (N_23539,N_20618,N_21497);
and U23540 (N_23540,N_20307,N_21717);
and U23541 (N_23541,N_22142,N_20067);
xor U23542 (N_23542,N_21305,N_21106);
nor U23543 (N_23543,N_20020,N_22019);
and U23544 (N_23544,N_22328,N_21231);
or U23545 (N_23545,N_22126,N_20544);
nand U23546 (N_23546,N_20306,N_22064);
nand U23547 (N_23547,N_21309,N_21704);
xnor U23548 (N_23548,N_20467,N_21390);
nor U23549 (N_23549,N_21168,N_20355);
nand U23550 (N_23550,N_20809,N_22150);
and U23551 (N_23551,N_21741,N_20861);
nand U23552 (N_23552,N_21413,N_20155);
and U23553 (N_23553,N_20183,N_21467);
nor U23554 (N_23554,N_20206,N_20526);
nor U23555 (N_23555,N_21520,N_21491);
xor U23556 (N_23556,N_21359,N_20520);
and U23557 (N_23557,N_20756,N_21342);
nor U23558 (N_23558,N_20900,N_20030);
nand U23559 (N_23559,N_20346,N_20078);
or U23560 (N_23560,N_21182,N_22374);
or U23561 (N_23561,N_21056,N_22332);
and U23562 (N_23562,N_21251,N_20921);
xnor U23563 (N_23563,N_22108,N_22288);
xor U23564 (N_23564,N_21440,N_22127);
nor U23565 (N_23565,N_20782,N_21040);
nand U23566 (N_23566,N_22296,N_21648);
nor U23567 (N_23567,N_20214,N_20325);
nand U23568 (N_23568,N_20056,N_21148);
and U23569 (N_23569,N_21211,N_21703);
nand U23570 (N_23570,N_21866,N_20657);
nor U23571 (N_23571,N_20197,N_21092);
nand U23572 (N_23572,N_21836,N_21630);
nand U23573 (N_23573,N_21945,N_20230);
nor U23574 (N_23574,N_20420,N_22404);
xnor U23575 (N_23575,N_21166,N_20269);
and U23576 (N_23576,N_22128,N_21018);
nor U23577 (N_23577,N_20983,N_21306);
xor U23578 (N_23578,N_22078,N_20459);
and U23579 (N_23579,N_21868,N_20514);
and U23580 (N_23580,N_20268,N_20150);
and U23581 (N_23581,N_20135,N_22382);
nor U23582 (N_23582,N_22053,N_21891);
nand U23583 (N_23583,N_21114,N_21119);
or U23584 (N_23584,N_20498,N_20585);
xor U23585 (N_23585,N_20587,N_20283);
xor U23586 (N_23586,N_20685,N_20146);
nor U23587 (N_23587,N_22148,N_20616);
nand U23588 (N_23588,N_20085,N_21585);
or U23589 (N_23589,N_20350,N_22169);
and U23590 (N_23590,N_21825,N_21921);
or U23591 (N_23591,N_21901,N_22299);
and U23592 (N_23592,N_20903,N_22277);
and U23593 (N_23593,N_21377,N_21808);
nand U23594 (N_23594,N_21346,N_22104);
or U23595 (N_23595,N_21900,N_20175);
or U23596 (N_23596,N_22139,N_20704);
and U23597 (N_23597,N_21411,N_22370);
nand U23598 (N_23598,N_21447,N_22101);
xnor U23599 (N_23599,N_20502,N_21139);
xor U23600 (N_23600,N_20747,N_20176);
nand U23601 (N_23601,N_21060,N_21716);
or U23602 (N_23602,N_22454,N_21111);
nor U23603 (N_23603,N_21506,N_20108);
or U23604 (N_23604,N_21653,N_21760);
or U23605 (N_23605,N_21333,N_21300);
nor U23606 (N_23606,N_21605,N_20458);
nand U23607 (N_23607,N_21981,N_21380);
nor U23608 (N_23608,N_21024,N_21143);
nand U23609 (N_23609,N_21025,N_21041);
nor U23610 (N_23610,N_20929,N_21434);
xnor U23611 (N_23611,N_22129,N_22243);
or U23612 (N_23612,N_22060,N_21806);
nor U23613 (N_23613,N_21123,N_22416);
and U23614 (N_23614,N_20316,N_20144);
and U23615 (N_23615,N_20810,N_20509);
and U23616 (N_23616,N_20978,N_20893);
nand U23617 (N_23617,N_20568,N_21455);
or U23618 (N_23618,N_21676,N_20107);
xor U23619 (N_23619,N_21206,N_21096);
nor U23620 (N_23620,N_20557,N_20215);
and U23621 (N_23621,N_21632,N_21693);
or U23622 (N_23622,N_21947,N_21514);
and U23623 (N_23623,N_22203,N_22118);
xnor U23624 (N_23624,N_21355,N_21639);
xor U23625 (N_23625,N_22103,N_22479);
xnor U23626 (N_23626,N_22494,N_21059);
or U23627 (N_23627,N_20441,N_20771);
xnor U23628 (N_23628,N_22105,N_20170);
or U23629 (N_23629,N_21493,N_20729);
xor U23630 (N_23630,N_20364,N_21169);
xor U23631 (N_23631,N_21867,N_20277);
nor U23632 (N_23632,N_20757,N_21933);
xor U23633 (N_23633,N_20034,N_20534);
nand U23634 (N_23634,N_20411,N_21833);
or U23635 (N_23635,N_22340,N_20689);
and U23636 (N_23636,N_22257,N_20220);
or U23637 (N_23637,N_20276,N_20944);
nand U23638 (N_23638,N_22437,N_20149);
nand U23639 (N_23639,N_21523,N_20965);
or U23640 (N_23640,N_21665,N_21978);
and U23641 (N_23641,N_21999,N_22123);
nor U23642 (N_23642,N_20227,N_21195);
nand U23643 (N_23643,N_22206,N_22024);
nor U23644 (N_23644,N_20589,N_20202);
nand U23645 (N_23645,N_20638,N_21274);
xor U23646 (N_23646,N_20143,N_20331);
nand U23647 (N_23647,N_22363,N_20378);
or U23648 (N_23648,N_20313,N_20748);
nand U23649 (N_23649,N_20580,N_21204);
nand U23650 (N_23650,N_20597,N_21217);
or U23651 (N_23651,N_20916,N_20298);
and U23652 (N_23652,N_20604,N_22121);
nor U23653 (N_23653,N_20052,N_20665);
nand U23654 (N_23654,N_22263,N_21167);
or U23655 (N_23655,N_22412,N_21915);
nand U23656 (N_23656,N_20447,N_21192);
or U23657 (N_23657,N_22192,N_21883);
or U23658 (N_23658,N_22344,N_20545);
nand U23659 (N_23659,N_20486,N_21134);
xnor U23660 (N_23660,N_20990,N_20789);
xnor U23661 (N_23661,N_20038,N_20867);
nand U23662 (N_23662,N_21343,N_20208);
and U23663 (N_23663,N_20024,N_22304);
nand U23664 (N_23664,N_20645,N_21993);
or U23665 (N_23665,N_20114,N_20347);
nor U23666 (N_23666,N_22221,N_20731);
or U23667 (N_23667,N_20510,N_20063);
or U23668 (N_23668,N_21419,N_20423);
nor U23669 (N_23669,N_20515,N_21125);
and U23670 (N_23670,N_20101,N_22106);
or U23671 (N_23671,N_21131,N_21358);
xor U23672 (N_23672,N_21903,N_20390);
xnor U23673 (N_23673,N_22199,N_21260);
and U23674 (N_23674,N_22144,N_20093);
nor U23675 (N_23675,N_20751,N_21563);
nand U23676 (N_23676,N_22032,N_20082);
or U23677 (N_23677,N_22046,N_22085);
nor U23678 (N_23678,N_21301,N_22196);
nor U23679 (N_23679,N_22028,N_21701);
and U23680 (N_23680,N_20409,N_22477);
and U23681 (N_23681,N_21641,N_20626);
or U23682 (N_23682,N_21635,N_20111);
or U23683 (N_23683,N_21838,N_20602);
nand U23684 (N_23684,N_21438,N_20555);
or U23685 (N_23685,N_21558,N_21071);
nand U23686 (N_23686,N_20435,N_21258);
nand U23687 (N_23687,N_21905,N_22017);
nor U23688 (N_23688,N_21397,N_20402);
or U23689 (N_23689,N_20868,N_20453);
and U23690 (N_23690,N_22355,N_21777);
or U23691 (N_23691,N_21449,N_21308);
xor U23692 (N_23692,N_21718,N_20852);
nand U23693 (N_23693,N_22063,N_20395);
and U23694 (N_23694,N_21142,N_20708);
or U23695 (N_23695,N_21528,N_20778);
and U23696 (N_23696,N_21587,N_20481);
nor U23697 (N_23697,N_21149,N_21102);
or U23698 (N_23698,N_20098,N_22116);
nand U23699 (N_23699,N_21452,N_20016);
or U23700 (N_23700,N_20003,N_22428);
nand U23701 (N_23701,N_21392,N_21898);
xnor U23702 (N_23702,N_21098,N_20513);
nand U23703 (N_23703,N_20142,N_21107);
xnor U23704 (N_23704,N_21982,N_20605);
nand U23705 (N_23705,N_22436,N_22423);
xor U23706 (N_23706,N_20724,N_20753);
nor U23707 (N_23707,N_21721,N_20720);
xor U23708 (N_23708,N_22461,N_20902);
nor U23709 (N_23709,N_21373,N_22136);
and U23710 (N_23710,N_20581,N_20013);
or U23711 (N_23711,N_22010,N_20804);
nand U23712 (N_23712,N_22290,N_20827);
or U23713 (N_23713,N_20173,N_21312);
and U23714 (N_23714,N_21784,N_22466);
nand U23715 (N_23715,N_21034,N_20691);
xnor U23716 (N_23716,N_22146,N_21917);
nor U23717 (N_23717,N_20169,N_20475);
and U23718 (N_23718,N_21987,N_20794);
or U23719 (N_23719,N_21426,N_22037);
xor U23720 (N_23720,N_21638,N_22188);
xor U23721 (N_23721,N_21627,N_22007);
nor U23722 (N_23722,N_20950,N_21554);
nand U23723 (N_23723,N_20369,N_20159);
nand U23724 (N_23724,N_21775,N_21595);
nand U23725 (N_23725,N_22360,N_21975);
and U23726 (N_23726,N_20172,N_21608);
xor U23727 (N_23727,N_21014,N_20643);
or U23728 (N_23728,N_21480,N_22022);
nand U23729 (N_23729,N_22234,N_21117);
and U23730 (N_23730,N_21175,N_20821);
nor U23731 (N_23731,N_22486,N_21053);
nor U23732 (N_23732,N_22361,N_20697);
or U23733 (N_23733,N_20715,N_22292);
nand U23734 (N_23734,N_21763,N_20993);
nor U23735 (N_23735,N_20223,N_21020);
nor U23736 (N_23736,N_20695,N_20469);
or U23737 (N_23737,N_20166,N_20712);
nor U23738 (N_23738,N_21002,N_20059);
nor U23739 (N_23739,N_20247,N_21645);
nand U23740 (N_23740,N_20263,N_20803);
nor U23741 (N_23741,N_21043,N_20924);
and U23742 (N_23742,N_21084,N_20851);
xnor U23743 (N_23743,N_22293,N_20393);
or U23744 (N_23744,N_21980,N_21527);
nand U23745 (N_23745,N_21658,N_21215);
xnor U23746 (N_23746,N_20764,N_20815);
and U23747 (N_23747,N_21958,N_21007);
nor U23748 (N_23748,N_20199,N_20859);
and U23749 (N_23749,N_21529,N_20519);
xnor U23750 (N_23750,N_21534,N_21823);
xnor U23751 (N_23751,N_20342,N_21630);
nor U23752 (N_23752,N_20905,N_21569);
and U23753 (N_23753,N_22111,N_21127);
and U23754 (N_23754,N_20764,N_20362);
or U23755 (N_23755,N_20289,N_20917);
nor U23756 (N_23756,N_22152,N_20946);
and U23757 (N_23757,N_20123,N_20406);
nand U23758 (N_23758,N_20589,N_21910);
nand U23759 (N_23759,N_20281,N_20211);
and U23760 (N_23760,N_21586,N_21678);
nand U23761 (N_23761,N_21261,N_20515);
nand U23762 (N_23762,N_21924,N_22092);
or U23763 (N_23763,N_20321,N_20931);
nand U23764 (N_23764,N_22452,N_22321);
or U23765 (N_23765,N_22200,N_21656);
nand U23766 (N_23766,N_21579,N_20693);
xor U23767 (N_23767,N_21378,N_21266);
xor U23768 (N_23768,N_20155,N_20160);
xnor U23769 (N_23769,N_20109,N_21425);
nor U23770 (N_23770,N_20310,N_20577);
nand U23771 (N_23771,N_21982,N_21186);
or U23772 (N_23772,N_20147,N_20591);
nor U23773 (N_23773,N_22452,N_21430);
nand U23774 (N_23774,N_22397,N_22324);
or U23775 (N_23775,N_20561,N_22342);
or U23776 (N_23776,N_21398,N_21514);
and U23777 (N_23777,N_22040,N_20985);
or U23778 (N_23778,N_20697,N_21352);
nor U23779 (N_23779,N_21995,N_21058);
or U23780 (N_23780,N_20659,N_20903);
and U23781 (N_23781,N_21923,N_20513);
or U23782 (N_23782,N_22489,N_20951);
nand U23783 (N_23783,N_22020,N_20400);
and U23784 (N_23784,N_20586,N_21841);
xnor U23785 (N_23785,N_21153,N_21555);
xnor U23786 (N_23786,N_20406,N_21160);
and U23787 (N_23787,N_20969,N_21065);
nor U23788 (N_23788,N_20514,N_22402);
xor U23789 (N_23789,N_21702,N_22259);
nor U23790 (N_23790,N_20066,N_21175);
and U23791 (N_23791,N_21827,N_21384);
and U23792 (N_23792,N_21956,N_21144);
nor U23793 (N_23793,N_21907,N_22109);
nor U23794 (N_23794,N_21913,N_22146);
xnor U23795 (N_23795,N_22350,N_21381);
xor U23796 (N_23796,N_21571,N_21171);
nand U23797 (N_23797,N_21941,N_21594);
and U23798 (N_23798,N_20823,N_21553);
xnor U23799 (N_23799,N_21165,N_20834);
or U23800 (N_23800,N_21504,N_20766);
or U23801 (N_23801,N_20848,N_21174);
nand U23802 (N_23802,N_20321,N_21217);
xor U23803 (N_23803,N_21362,N_21821);
xnor U23804 (N_23804,N_21850,N_20230);
xnor U23805 (N_23805,N_20438,N_20360);
or U23806 (N_23806,N_20379,N_20695);
or U23807 (N_23807,N_21092,N_21722);
nor U23808 (N_23808,N_21046,N_20571);
nor U23809 (N_23809,N_20291,N_21370);
xor U23810 (N_23810,N_21684,N_20797);
and U23811 (N_23811,N_20111,N_22088);
xor U23812 (N_23812,N_21665,N_21523);
nand U23813 (N_23813,N_22220,N_21162);
nor U23814 (N_23814,N_20475,N_21917);
xnor U23815 (N_23815,N_20623,N_20727);
nor U23816 (N_23816,N_21039,N_22213);
nand U23817 (N_23817,N_21988,N_21974);
or U23818 (N_23818,N_21023,N_21636);
nor U23819 (N_23819,N_20589,N_21234);
or U23820 (N_23820,N_22113,N_21089);
or U23821 (N_23821,N_20377,N_20043);
and U23822 (N_23822,N_21561,N_21191);
nor U23823 (N_23823,N_20856,N_20536);
nor U23824 (N_23824,N_21661,N_21837);
nand U23825 (N_23825,N_20165,N_22364);
nor U23826 (N_23826,N_20865,N_21295);
nor U23827 (N_23827,N_22175,N_21343);
nand U23828 (N_23828,N_20429,N_20292);
and U23829 (N_23829,N_21086,N_20545);
nand U23830 (N_23830,N_20614,N_21578);
xor U23831 (N_23831,N_20980,N_20787);
nor U23832 (N_23832,N_20862,N_20293);
nor U23833 (N_23833,N_20999,N_21589);
and U23834 (N_23834,N_20312,N_20858);
nand U23835 (N_23835,N_21963,N_22281);
and U23836 (N_23836,N_20261,N_22315);
and U23837 (N_23837,N_20961,N_20316);
nor U23838 (N_23838,N_20986,N_21205);
xnor U23839 (N_23839,N_21391,N_22213);
nand U23840 (N_23840,N_20529,N_22427);
xor U23841 (N_23841,N_20612,N_20935);
nor U23842 (N_23842,N_20690,N_20392);
xnor U23843 (N_23843,N_22194,N_20581);
nand U23844 (N_23844,N_21844,N_20346);
xnor U23845 (N_23845,N_21732,N_21123);
and U23846 (N_23846,N_21697,N_20136);
nand U23847 (N_23847,N_22164,N_22223);
xor U23848 (N_23848,N_20198,N_20296);
and U23849 (N_23849,N_21326,N_20764);
and U23850 (N_23850,N_20615,N_21912);
and U23851 (N_23851,N_21255,N_21892);
xor U23852 (N_23852,N_22238,N_20516);
nand U23853 (N_23853,N_20494,N_21366);
or U23854 (N_23854,N_20685,N_21365);
or U23855 (N_23855,N_20430,N_21690);
nor U23856 (N_23856,N_22034,N_21476);
or U23857 (N_23857,N_21358,N_21841);
xnor U23858 (N_23858,N_22255,N_20404);
or U23859 (N_23859,N_21705,N_21710);
or U23860 (N_23860,N_20776,N_20288);
or U23861 (N_23861,N_22424,N_22020);
and U23862 (N_23862,N_20406,N_20978);
and U23863 (N_23863,N_21857,N_22306);
and U23864 (N_23864,N_22046,N_20198);
nor U23865 (N_23865,N_22134,N_20790);
or U23866 (N_23866,N_22062,N_21803);
xor U23867 (N_23867,N_20878,N_22467);
and U23868 (N_23868,N_20139,N_20239);
or U23869 (N_23869,N_20265,N_20204);
xnor U23870 (N_23870,N_21922,N_21663);
nor U23871 (N_23871,N_20091,N_21117);
nand U23872 (N_23872,N_21294,N_20589);
xnor U23873 (N_23873,N_21348,N_22406);
nor U23874 (N_23874,N_21237,N_20653);
and U23875 (N_23875,N_20519,N_22201);
nor U23876 (N_23876,N_20763,N_20983);
xnor U23877 (N_23877,N_22201,N_22198);
and U23878 (N_23878,N_22116,N_21011);
xnor U23879 (N_23879,N_20816,N_21332);
and U23880 (N_23880,N_22235,N_20525);
or U23881 (N_23881,N_21721,N_20893);
nand U23882 (N_23882,N_21329,N_20568);
or U23883 (N_23883,N_20710,N_20971);
xnor U23884 (N_23884,N_20296,N_20450);
or U23885 (N_23885,N_20793,N_20318);
and U23886 (N_23886,N_21474,N_20903);
nand U23887 (N_23887,N_20889,N_20176);
or U23888 (N_23888,N_20842,N_20517);
xor U23889 (N_23889,N_20385,N_21242);
nand U23890 (N_23890,N_21233,N_20993);
nand U23891 (N_23891,N_21885,N_21591);
nand U23892 (N_23892,N_20469,N_22374);
xor U23893 (N_23893,N_21427,N_21595);
or U23894 (N_23894,N_20737,N_20611);
nor U23895 (N_23895,N_22007,N_20414);
and U23896 (N_23896,N_20636,N_20803);
xor U23897 (N_23897,N_20810,N_20859);
and U23898 (N_23898,N_21776,N_21337);
and U23899 (N_23899,N_22026,N_21302);
or U23900 (N_23900,N_21416,N_20318);
and U23901 (N_23901,N_21357,N_21043);
and U23902 (N_23902,N_20098,N_20505);
nand U23903 (N_23903,N_21977,N_20156);
xor U23904 (N_23904,N_22073,N_21220);
nand U23905 (N_23905,N_21384,N_21774);
or U23906 (N_23906,N_22475,N_21507);
and U23907 (N_23907,N_22044,N_21656);
or U23908 (N_23908,N_22059,N_22036);
or U23909 (N_23909,N_21029,N_20646);
or U23910 (N_23910,N_21554,N_20829);
xor U23911 (N_23911,N_21651,N_22338);
or U23912 (N_23912,N_21135,N_21540);
nand U23913 (N_23913,N_21176,N_21676);
or U23914 (N_23914,N_20008,N_20919);
xor U23915 (N_23915,N_20812,N_21452);
and U23916 (N_23916,N_20486,N_22235);
nand U23917 (N_23917,N_22333,N_21607);
xnor U23918 (N_23918,N_21209,N_21805);
nand U23919 (N_23919,N_20473,N_20928);
nand U23920 (N_23920,N_20999,N_20700);
nor U23921 (N_23921,N_20746,N_21606);
nand U23922 (N_23922,N_21943,N_21196);
and U23923 (N_23923,N_22130,N_22499);
nand U23924 (N_23924,N_21494,N_20037);
nand U23925 (N_23925,N_21665,N_21470);
nor U23926 (N_23926,N_20963,N_21044);
xor U23927 (N_23927,N_22258,N_20206);
or U23928 (N_23928,N_21972,N_22461);
or U23929 (N_23929,N_21635,N_20175);
and U23930 (N_23930,N_22252,N_20173);
nand U23931 (N_23931,N_21016,N_21218);
nand U23932 (N_23932,N_20380,N_22336);
nand U23933 (N_23933,N_21918,N_21873);
xor U23934 (N_23934,N_21468,N_20359);
nor U23935 (N_23935,N_21650,N_20794);
or U23936 (N_23936,N_20330,N_21992);
nor U23937 (N_23937,N_22017,N_21080);
and U23938 (N_23938,N_21646,N_21918);
nor U23939 (N_23939,N_21392,N_20053);
nand U23940 (N_23940,N_20921,N_20199);
or U23941 (N_23941,N_21541,N_20002);
and U23942 (N_23942,N_21624,N_21401);
or U23943 (N_23943,N_20010,N_20404);
or U23944 (N_23944,N_22299,N_21592);
nor U23945 (N_23945,N_21538,N_20568);
or U23946 (N_23946,N_20425,N_21286);
or U23947 (N_23947,N_20973,N_20937);
and U23948 (N_23948,N_20019,N_20064);
or U23949 (N_23949,N_21629,N_20246);
and U23950 (N_23950,N_21036,N_20427);
and U23951 (N_23951,N_21091,N_20492);
or U23952 (N_23952,N_21343,N_20603);
and U23953 (N_23953,N_22094,N_21067);
and U23954 (N_23954,N_21591,N_21541);
nor U23955 (N_23955,N_21961,N_21437);
and U23956 (N_23956,N_20507,N_21584);
nand U23957 (N_23957,N_20704,N_22154);
xor U23958 (N_23958,N_21333,N_21004);
nor U23959 (N_23959,N_21785,N_21648);
xnor U23960 (N_23960,N_20723,N_22394);
or U23961 (N_23961,N_20324,N_20716);
and U23962 (N_23962,N_21665,N_20363);
nand U23963 (N_23963,N_20273,N_21896);
and U23964 (N_23964,N_20898,N_20949);
xor U23965 (N_23965,N_20548,N_20845);
xor U23966 (N_23966,N_21108,N_21757);
xor U23967 (N_23967,N_21069,N_20614);
nor U23968 (N_23968,N_21569,N_21062);
nand U23969 (N_23969,N_21341,N_21721);
nor U23970 (N_23970,N_20223,N_22235);
and U23971 (N_23971,N_20372,N_20205);
nand U23972 (N_23972,N_22005,N_20898);
xor U23973 (N_23973,N_21915,N_22211);
xor U23974 (N_23974,N_21537,N_21637);
or U23975 (N_23975,N_21821,N_20306);
nand U23976 (N_23976,N_22428,N_20872);
or U23977 (N_23977,N_20071,N_20751);
nor U23978 (N_23978,N_22224,N_21563);
or U23979 (N_23979,N_21215,N_21969);
and U23980 (N_23980,N_22225,N_21068);
xnor U23981 (N_23981,N_21003,N_21133);
nor U23982 (N_23982,N_20888,N_20854);
nand U23983 (N_23983,N_22063,N_20043);
xnor U23984 (N_23984,N_22305,N_21419);
or U23985 (N_23985,N_22457,N_20595);
nor U23986 (N_23986,N_21296,N_21107);
nand U23987 (N_23987,N_20466,N_21177);
xnor U23988 (N_23988,N_20316,N_22364);
xor U23989 (N_23989,N_20124,N_20265);
or U23990 (N_23990,N_20244,N_22375);
nand U23991 (N_23991,N_20101,N_21967);
nor U23992 (N_23992,N_20639,N_20741);
and U23993 (N_23993,N_20649,N_20783);
nand U23994 (N_23994,N_21108,N_22043);
and U23995 (N_23995,N_20978,N_20065);
and U23996 (N_23996,N_22116,N_22471);
or U23997 (N_23997,N_22303,N_21418);
or U23998 (N_23998,N_20136,N_21872);
nor U23999 (N_23999,N_20449,N_20930);
nor U24000 (N_24000,N_22443,N_20788);
or U24001 (N_24001,N_21635,N_20267);
and U24002 (N_24002,N_21988,N_22044);
nor U24003 (N_24003,N_21406,N_21597);
nand U24004 (N_24004,N_21041,N_20733);
nor U24005 (N_24005,N_20143,N_20404);
or U24006 (N_24006,N_21761,N_22141);
and U24007 (N_24007,N_20647,N_20844);
xnor U24008 (N_24008,N_22267,N_22004);
and U24009 (N_24009,N_21469,N_21823);
or U24010 (N_24010,N_21744,N_21475);
and U24011 (N_24011,N_21615,N_20630);
nand U24012 (N_24012,N_20613,N_20624);
nor U24013 (N_24013,N_20956,N_20346);
xor U24014 (N_24014,N_21823,N_20265);
nor U24015 (N_24015,N_21978,N_22211);
and U24016 (N_24016,N_21430,N_21582);
and U24017 (N_24017,N_21653,N_22222);
xor U24018 (N_24018,N_21347,N_22258);
xor U24019 (N_24019,N_20742,N_22293);
nand U24020 (N_24020,N_20378,N_22269);
xor U24021 (N_24021,N_21505,N_20231);
or U24022 (N_24022,N_21048,N_20831);
nor U24023 (N_24023,N_21507,N_20876);
nand U24024 (N_24024,N_20391,N_21228);
or U24025 (N_24025,N_20410,N_21745);
nand U24026 (N_24026,N_20973,N_21758);
or U24027 (N_24027,N_20421,N_21741);
xor U24028 (N_24028,N_20207,N_21764);
nor U24029 (N_24029,N_21653,N_21898);
nand U24030 (N_24030,N_21519,N_20251);
nor U24031 (N_24031,N_21090,N_20338);
nor U24032 (N_24032,N_20560,N_21787);
or U24033 (N_24033,N_21446,N_20155);
nand U24034 (N_24034,N_20315,N_21641);
xor U24035 (N_24035,N_21244,N_20156);
or U24036 (N_24036,N_21998,N_21814);
nand U24037 (N_24037,N_20876,N_21672);
and U24038 (N_24038,N_20429,N_21262);
nor U24039 (N_24039,N_21942,N_21501);
and U24040 (N_24040,N_21070,N_20940);
nand U24041 (N_24041,N_22329,N_20282);
or U24042 (N_24042,N_20967,N_21600);
nor U24043 (N_24043,N_21400,N_20700);
and U24044 (N_24044,N_20343,N_21670);
nand U24045 (N_24045,N_20643,N_21368);
xnor U24046 (N_24046,N_21672,N_21610);
and U24047 (N_24047,N_21652,N_21538);
and U24048 (N_24048,N_20909,N_20310);
or U24049 (N_24049,N_21066,N_21815);
or U24050 (N_24050,N_22026,N_20178);
nor U24051 (N_24051,N_20110,N_20554);
nand U24052 (N_24052,N_22058,N_21116);
nand U24053 (N_24053,N_22498,N_22380);
and U24054 (N_24054,N_21495,N_20473);
nor U24055 (N_24055,N_20852,N_20638);
or U24056 (N_24056,N_21889,N_20965);
nor U24057 (N_24057,N_21917,N_20841);
or U24058 (N_24058,N_21646,N_22003);
and U24059 (N_24059,N_21233,N_22096);
nor U24060 (N_24060,N_20805,N_22040);
nand U24061 (N_24061,N_21119,N_20328);
and U24062 (N_24062,N_20564,N_21709);
or U24063 (N_24063,N_22183,N_20708);
xnor U24064 (N_24064,N_21946,N_21428);
or U24065 (N_24065,N_21502,N_21494);
nand U24066 (N_24066,N_22056,N_20289);
or U24067 (N_24067,N_22363,N_22184);
or U24068 (N_24068,N_21858,N_21771);
nand U24069 (N_24069,N_21005,N_21171);
and U24070 (N_24070,N_22246,N_20904);
or U24071 (N_24071,N_20329,N_21599);
or U24072 (N_24072,N_20147,N_20176);
or U24073 (N_24073,N_20979,N_21721);
xor U24074 (N_24074,N_20404,N_20265);
nor U24075 (N_24075,N_20325,N_22057);
nand U24076 (N_24076,N_20078,N_22294);
or U24077 (N_24077,N_21098,N_21609);
and U24078 (N_24078,N_21500,N_21301);
xor U24079 (N_24079,N_21006,N_20059);
xnor U24080 (N_24080,N_21348,N_20049);
nor U24081 (N_24081,N_21590,N_20248);
nor U24082 (N_24082,N_20981,N_21070);
xnor U24083 (N_24083,N_21597,N_21672);
and U24084 (N_24084,N_21857,N_21851);
nor U24085 (N_24085,N_21423,N_20174);
or U24086 (N_24086,N_21824,N_20268);
nand U24087 (N_24087,N_21955,N_22456);
nand U24088 (N_24088,N_20031,N_20143);
or U24089 (N_24089,N_20407,N_20760);
nor U24090 (N_24090,N_20240,N_21317);
and U24091 (N_24091,N_21694,N_20668);
or U24092 (N_24092,N_22022,N_20317);
nand U24093 (N_24093,N_20857,N_21246);
and U24094 (N_24094,N_21355,N_22412);
xor U24095 (N_24095,N_22356,N_20150);
xnor U24096 (N_24096,N_20503,N_22306);
or U24097 (N_24097,N_21770,N_20151);
and U24098 (N_24098,N_21327,N_21212);
and U24099 (N_24099,N_21212,N_21665);
xor U24100 (N_24100,N_22397,N_21377);
and U24101 (N_24101,N_20550,N_21031);
nor U24102 (N_24102,N_22379,N_21231);
nand U24103 (N_24103,N_22294,N_21961);
nor U24104 (N_24104,N_20760,N_20791);
and U24105 (N_24105,N_21154,N_21187);
and U24106 (N_24106,N_20714,N_21537);
nor U24107 (N_24107,N_20006,N_21027);
nand U24108 (N_24108,N_20165,N_20960);
nand U24109 (N_24109,N_22262,N_21192);
or U24110 (N_24110,N_20673,N_20032);
and U24111 (N_24111,N_20165,N_20601);
or U24112 (N_24112,N_20022,N_22360);
xnor U24113 (N_24113,N_20061,N_22345);
or U24114 (N_24114,N_21982,N_20294);
and U24115 (N_24115,N_20289,N_20214);
nor U24116 (N_24116,N_20831,N_22314);
nor U24117 (N_24117,N_20717,N_20521);
xor U24118 (N_24118,N_20155,N_20792);
and U24119 (N_24119,N_21628,N_22215);
or U24120 (N_24120,N_21873,N_21686);
xor U24121 (N_24121,N_21373,N_20131);
xnor U24122 (N_24122,N_21593,N_21271);
nor U24123 (N_24123,N_22015,N_20737);
and U24124 (N_24124,N_22271,N_20359);
nor U24125 (N_24125,N_21357,N_22498);
and U24126 (N_24126,N_21471,N_20839);
and U24127 (N_24127,N_20715,N_20482);
and U24128 (N_24128,N_21599,N_20252);
or U24129 (N_24129,N_21110,N_20169);
xnor U24130 (N_24130,N_22345,N_21435);
and U24131 (N_24131,N_21800,N_22130);
or U24132 (N_24132,N_21427,N_22252);
xor U24133 (N_24133,N_21044,N_21112);
nor U24134 (N_24134,N_21546,N_20177);
and U24135 (N_24135,N_20392,N_22120);
and U24136 (N_24136,N_21612,N_22171);
nor U24137 (N_24137,N_20339,N_21743);
and U24138 (N_24138,N_20390,N_20376);
nor U24139 (N_24139,N_22273,N_21609);
and U24140 (N_24140,N_22247,N_21777);
xnor U24141 (N_24141,N_20081,N_21378);
xor U24142 (N_24142,N_22386,N_20217);
and U24143 (N_24143,N_20157,N_22142);
nor U24144 (N_24144,N_21396,N_21891);
xor U24145 (N_24145,N_20582,N_21687);
or U24146 (N_24146,N_21030,N_22298);
nand U24147 (N_24147,N_21650,N_22488);
nand U24148 (N_24148,N_21292,N_21703);
nor U24149 (N_24149,N_21245,N_21779);
and U24150 (N_24150,N_21395,N_20034);
xnor U24151 (N_24151,N_20663,N_20532);
nand U24152 (N_24152,N_21104,N_21008);
nand U24153 (N_24153,N_22176,N_21030);
xnor U24154 (N_24154,N_21142,N_20586);
nand U24155 (N_24155,N_22260,N_20294);
and U24156 (N_24156,N_21289,N_20365);
xor U24157 (N_24157,N_20069,N_21310);
or U24158 (N_24158,N_20681,N_20724);
and U24159 (N_24159,N_21400,N_20462);
and U24160 (N_24160,N_20023,N_20634);
or U24161 (N_24161,N_21129,N_21487);
or U24162 (N_24162,N_20191,N_22358);
xor U24163 (N_24163,N_20413,N_22151);
or U24164 (N_24164,N_20207,N_20527);
and U24165 (N_24165,N_21829,N_21091);
xor U24166 (N_24166,N_22478,N_21044);
xnor U24167 (N_24167,N_20653,N_21385);
xor U24168 (N_24168,N_20275,N_22495);
nand U24169 (N_24169,N_21433,N_21789);
nor U24170 (N_24170,N_21201,N_21175);
nand U24171 (N_24171,N_20189,N_21580);
nand U24172 (N_24172,N_20866,N_20045);
xor U24173 (N_24173,N_21052,N_20847);
and U24174 (N_24174,N_21678,N_20873);
nand U24175 (N_24175,N_22169,N_21065);
nand U24176 (N_24176,N_22073,N_21446);
or U24177 (N_24177,N_21138,N_21804);
and U24178 (N_24178,N_20354,N_21015);
or U24179 (N_24179,N_20003,N_21615);
or U24180 (N_24180,N_22411,N_21831);
or U24181 (N_24181,N_20585,N_21750);
nand U24182 (N_24182,N_21490,N_22017);
nand U24183 (N_24183,N_21485,N_21738);
and U24184 (N_24184,N_20438,N_20938);
xor U24185 (N_24185,N_21365,N_22042);
nand U24186 (N_24186,N_20857,N_21535);
nand U24187 (N_24187,N_20804,N_20432);
nor U24188 (N_24188,N_20968,N_21392);
nor U24189 (N_24189,N_21608,N_21229);
nand U24190 (N_24190,N_20408,N_21759);
or U24191 (N_24191,N_22216,N_20790);
or U24192 (N_24192,N_22210,N_20386);
or U24193 (N_24193,N_20505,N_22232);
or U24194 (N_24194,N_21064,N_20055);
nand U24195 (N_24195,N_21263,N_22243);
nand U24196 (N_24196,N_21983,N_21425);
or U24197 (N_24197,N_21940,N_21117);
or U24198 (N_24198,N_20587,N_21622);
and U24199 (N_24199,N_22030,N_20642);
or U24200 (N_24200,N_20608,N_21048);
and U24201 (N_24201,N_22231,N_22185);
xor U24202 (N_24202,N_20597,N_21864);
and U24203 (N_24203,N_21328,N_21045);
and U24204 (N_24204,N_22216,N_20183);
and U24205 (N_24205,N_21943,N_21675);
nor U24206 (N_24206,N_21592,N_21522);
and U24207 (N_24207,N_21852,N_22240);
or U24208 (N_24208,N_21542,N_21144);
nand U24209 (N_24209,N_22355,N_21679);
nand U24210 (N_24210,N_21464,N_20753);
nand U24211 (N_24211,N_20689,N_20060);
and U24212 (N_24212,N_21802,N_20159);
and U24213 (N_24213,N_22063,N_21623);
xnor U24214 (N_24214,N_21619,N_20925);
nand U24215 (N_24215,N_20658,N_22194);
xnor U24216 (N_24216,N_21766,N_20720);
and U24217 (N_24217,N_21771,N_22458);
nand U24218 (N_24218,N_22460,N_22286);
nand U24219 (N_24219,N_21958,N_21071);
and U24220 (N_24220,N_20284,N_21774);
and U24221 (N_24221,N_21443,N_20723);
and U24222 (N_24222,N_21590,N_21510);
xor U24223 (N_24223,N_21642,N_20745);
xor U24224 (N_24224,N_20025,N_22479);
xnor U24225 (N_24225,N_20381,N_21043);
and U24226 (N_24226,N_22355,N_21774);
or U24227 (N_24227,N_22109,N_20385);
nand U24228 (N_24228,N_20925,N_21978);
nand U24229 (N_24229,N_20368,N_21243);
and U24230 (N_24230,N_21287,N_21677);
or U24231 (N_24231,N_21948,N_22419);
or U24232 (N_24232,N_21426,N_22047);
or U24233 (N_24233,N_21785,N_21546);
xor U24234 (N_24234,N_21434,N_21297);
or U24235 (N_24235,N_20973,N_20684);
or U24236 (N_24236,N_20424,N_20915);
nand U24237 (N_24237,N_22226,N_20564);
nor U24238 (N_24238,N_21549,N_21228);
or U24239 (N_24239,N_20779,N_20115);
or U24240 (N_24240,N_20153,N_20661);
and U24241 (N_24241,N_20172,N_20338);
nand U24242 (N_24242,N_20746,N_21748);
or U24243 (N_24243,N_21844,N_21699);
nor U24244 (N_24244,N_22384,N_21949);
or U24245 (N_24245,N_20475,N_22028);
nand U24246 (N_24246,N_20715,N_20945);
xnor U24247 (N_24247,N_22217,N_21624);
nand U24248 (N_24248,N_20364,N_21674);
or U24249 (N_24249,N_21087,N_21674);
xnor U24250 (N_24250,N_20846,N_22257);
xor U24251 (N_24251,N_21244,N_22004);
and U24252 (N_24252,N_21842,N_21718);
nor U24253 (N_24253,N_21983,N_21729);
or U24254 (N_24254,N_22180,N_21875);
xor U24255 (N_24255,N_21049,N_20578);
xnor U24256 (N_24256,N_20148,N_20102);
xor U24257 (N_24257,N_20558,N_20072);
nand U24258 (N_24258,N_22131,N_20426);
nand U24259 (N_24259,N_22231,N_22339);
xnor U24260 (N_24260,N_21020,N_21082);
or U24261 (N_24261,N_20146,N_21255);
or U24262 (N_24262,N_21484,N_20918);
xnor U24263 (N_24263,N_21400,N_21479);
or U24264 (N_24264,N_20235,N_20660);
xor U24265 (N_24265,N_21770,N_20637);
nor U24266 (N_24266,N_21733,N_22082);
xor U24267 (N_24267,N_20829,N_20404);
xnor U24268 (N_24268,N_21387,N_22137);
and U24269 (N_24269,N_22158,N_20376);
nor U24270 (N_24270,N_21761,N_20281);
xnor U24271 (N_24271,N_22085,N_21357);
and U24272 (N_24272,N_22351,N_21928);
nand U24273 (N_24273,N_22244,N_20342);
xor U24274 (N_24274,N_21512,N_22301);
nor U24275 (N_24275,N_21970,N_22173);
nand U24276 (N_24276,N_21037,N_20272);
and U24277 (N_24277,N_21645,N_20825);
nor U24278 (N_24278,N_21840,N_20955);
or U24279 (N_24279,N_22249,N_22430);
nor U24280 (N_24280,N_20012,N_21374);
or U24281 (N_24281,N_21602,N_21244);
or U24282 (N_24282,N_20398,N_22456);
nand U24283 (N_24283,N_22358,N_20083);
nor U24284 (N_24284,N_21489,N_21854);
and U24285 (N_24285,N_21656,N_20382);
nor U24286 (N_24286,N_20575,N_22355);
and U24287 (N_24287,N_21698,N_20388);
and U24288 (N_24288,N_20008,N_22339);
nor U24289 (N_24289,N_22180,N_21919);
nor U24290 (N_24290,N_21612,N_22156);
and U24291 (N_24291,N_21712,N_20662);
nand U24292 (N_24292,N_21816,N_21895);
nor U24293 (N_24293,N_21513,N_20050);
nor U24294 (N_24294,N_21544,N_22214);
and U24295 (N_24295,N_21504,N_20557);
and U24296 (N_24296,N_20749,N_22192);
or U24297 (N_24297,N_21892,N_20499);
or U24298 (N_24298,N_20944,N_20926);
xnor U24299 (N_24299,N_20377,N_20662);
nand U24300 (N_24300,N_22415,N_20418);
or U24301 (N_24301,N_20313,N_21036);
xnor U24302 (N_24302,N_20069,N_21146);
nor U24303 (N_24303,N_22186,N_21783);
and U24304 (N_24304,N_21055,N_22029);
xnor U24305 (N_24305,N_21070,N_21492);
or U24306 (N_24306,N_21556,N_20051);
xor U24307 (N_24307,N_20423,N_21073);
xnor U24308 (N_24308,N_20631,N_22474);
xor U24309 (N_24309,N_20424,N_20967);
nand U24310 (N_24310,N_20446,N_20424);
nor U24311 (N_24311,N_20003,N_21496);
and U24312 (N_24312,N_20082,N_21746);
nand U24313 (N_24313,N_20894,N_20821);
or U24314 (N_24314,N_20274,N_21156);
nand U24315 (N_24315,N_20850,N_22315);
and U24316 (N_24316,N_20133,N_20646);
nand U24317 (N_24317,N_20287,N_22007);
nor U24318 (N_24318,N_20473,N_21566);
nor U24319 (N_24319,N_20131,N_20755);
or U24320 (N_24320,N_20963,N_21251);
or U24321 (N_24321,N_21507,N_22412);
nor U24322 (N_24322,N_21347,N_21051);
nand U24323 (N_24323,N_21477,N_20311);
xnor U24324 (N_24324,N_21794,N_21429);
or U24325 (N_24325,N_20001,N_20479);
xor U24326 (N_24326,N_21646,N_22009);
nand U24327 (N_24327,N_21171,N_20998);
xnor U24328 (N_24328,N_20118,N_22037);
or U24329 (N_24329,N_20513,N_22347);
nor U24330 (N_24330,N_20166,N_21455);
and U24331 (N_24331,N_20075,N_22272);
or U24332 (N_24332,N_20210,N_21178);
nor U24333 (N_24333,N_20247,N_22117);
or U24334 (N_24334,N_20020,N_20372);
xnor U24335 (N_24335,N_21618,N_21702);
and U24336 (N_24336,N_20866,N_22268);
nor U24337 (N_24337,N_21940,N_20952);
nor U24338 (N_24338,N_20757,N_20511);
nor U24339 (N_24339,N_20217,N_20477);
or U24340 (N_24340,N_21471,N_21466);
xnor U24341 (N_24341,N_21083,N_20754);
or U24342 (N_24342,N_22297,N_22179);
xor U24343 (N_24343,N_20210,N_21389);
or U24344 (N_24344,N_20105,N_21137);
nor U24345 (N_24345,N_21918,N_22117);
or U24346 (N_24346,N_22059,N_20877);
and U24347 (N_24347,N_20427,N_21600);
nand U24348 (N_24348,N_20528,N_20592);
xnor U24349 (N_24349,N_22303,N_21701);
nor U24350 (N_24350,N_20197,N_21095);
nor U24351 (N_24351,N_22296,N_21857);
nand U24352 (N_24352,N_20879,N_21904);
nor U24353 (N_24353,N_21472,N_20334);
nor U24354 (N_24354,N_22390,N_20230);
nand U24355 (N_24355,N_21006,N_20515);
xnor U24356 (N_24356,N_21838,N_20365);
xor U24357 (N_24357,N_20344,N_21856);
nor U24358 (N_24358,N_21365,N_20674);
and U24359 (N_24359,N_21751,N_21049);
and U24360 (N_24360,N_20892,N_20777);
xor U24361 (N_24361,N_21874,N_21451);
nor U24362 (N_24362,N_20048,N_21788);
or U24363 (N_24363,N_21506,N_22389);
and U24364 (N_24364,N_21377,N_20902);
nor U24365 (N_24365,N_20023,N_20031);
nand U24366 (N_24366,N_21731,N_21349);
nor U24367 (N_24367,N_21890,N_22024);
nor U24368 (N_24368,N_22340,N_20164);
or U24369 (N_24369,N_20845,N_22349);
xor U24370 (N_24370,N_22225,N_20994);
and U24371 (N_24371,N_20936,N_21767);
xnor U24372 (N_24372,N_21347,N_21976);
nor U24373 (N_24373,N_22039,N_20770);
xnor U24374 (N_24374,N_21686,N_22125);
and U24375 (N_24375,N_21762,N_20044);
nor U24376 (N_24376,N_21009,N_20596);
nand U24377 (N_24377,N_21351,N_20318);
or U24378 (N_24378,N_22081,N_22097);
xor U24379 (N_24379,N_20095,N_20036);
or U24380 (N_24380,N_20262,N_21829);
xnor U24381 (N_24381,N_21429,N_20568);
xor U24382 (N_24382,N_20713,N_20584);
or U24383 (N_24383,N_20002,N_22341);
and U24384 (N_24384,N_21309,N_20830);
and U24385 (N_24385,N_20468,N_21173);
nand U24386 (N_24386,N_22420,N_20560);
nand U24387 (N_24387,N_20121,N_20976);
nand U24388 (N_24388,N_20072,N_22236);
nor U24389 (N_24389,N_21699,N_21621);
or U24390 (N_24390,N_21010,N_20863);
nor U24391 (N_24391,N_22278,N_22029);
xnor U24392 (N_24392,N_22489,N_20132);
nand U24393 (N_24393,N_22136,N_20148);
nor U24394 (N_24394,N_21840,N_22439);
xnor U24395 (N_24395,N_21101,N_21938);
or U24396 (N_24396,N_20373,N_20474);
nand U24397 (N_24397,N_21286,N_20683);
and U24398 (N_24398,N_21830,N_22225);
nand U24399 (N_24399,N_21283,N_20911);
nand U24400 (N_24400,N_20498,N_20789);
nand U24401 (N_24401,N_21306,N_21529);
nor U24402 (N_24402,N_20230,N_21921);
xor U24403 (N_24403,N_21903,N_22381);
and U24404 (N_24404,N_21529,N_22011);
nand U24405 (N_24405,N_20952,N_22385);
nand U24406 (N_24406,N_21820,N_22347);
or U24407 (N_24407,N_21485,N_20629);
or U24408 (N_24408,N_20510,N_21981);
nand U24409 (N_24409,N_20702,N_20987);
nor U24410 (N_24410,N_20040,N_21846);
or U24411 (N_24411,N_21040,N_21843);
or U24412 (N_24412,N_21595,N_21394);
and U24413 (N_24413,N_20107,N_21923);
or U24414 (N_24414,N_21934,N_21346);
nor U24415 (N_24415,N_22007,N_21843);
or U24416 (N_24416,N_22481,N_21119);
nor U24417 (N_24417,N_21481,N_22158);
and U24418 (N_24418,N_21828,N_20450);
nand U24419 (N_24419,N_21335,N_21265);
nand U24420 (N_24420,N_20136,N_21992);
xnor U24421 (N_24421,N_21518,N_22183);
nand U24422 (N_24422,N_20240,N_20677);
nor U24423 (N_24423,N_21018,N_20623);
nor U24424 (N_24424,N_20405,N_22094);
and U24425 (N_24425,N_21447,N_21792);
or U24426 (N_24426,N_21943,N_21107);
nand U24427 (N_24427,N_20298,N_20956);
and U24428 (N_24428,N_20700,N_20152);
nand U24429 (N_24429,N_20046,N_20555);
nand U24430 (N_24430,N_20197,N_20831);
nand U24431 (N_24431,N_21185,N_20424);
and U24432 (N_24432,N_20235,N_21384);
nor U24433 (N_24433,N_21074,N_21726);
xor U24434 (N_24434,N_21473,N_20361);
nand U24435 (N_24435,N_21579,N_21656);
nor U24436 (N_24436,N_21461,N_20289);
nor U24437 (N_24437,N_21313,N_21746);
nor U24438 (N_24438,N_20400,N_20053);
and U24439 (N_24439,N_21062,N_20283);
nand U24440 (N_24440,N_20471,N_21967);
or U24441 (N_24441,N_22123,N_22167);
nand U24442 (N_24442,N_20824,N_20873);
or U24443 (N_24443,N_21664,N_21377);
nand U24444 (N_24444,N_21254,N_21441);
or U24445 (N_24445,N_20633,N_21747);
nand U24446 (N_24446,N_22107,N_20879);
nand U24447 (N_24447,N_21051,N_21663);
or U24448 (N_24448,N_21274,N_21240);
and U24449 (N_24449,N_21884,N_22012);
nor U24450 (N_24450,N_20762,N_20629);
nor U24451 (N_24451,N_20696,N_20632);
nand U24452 (N_24452,N_21044,N_21088);
or U24453 (N_24453,N_22214,N_22438);
and U24454 (N_24454,N_20613,N_21085);
and U24455 (N_24455,N_20905,N_20274);
xor U24456 (N_24456,N_21491,N_20681);
nor U24457 (N_24457,N_22393,N_20771);
and U24458 (N_24458,N_21151,N_22001);
xnor U24459 (N_24459,N_20482,N_21298);
or U24460 (N_24460,N_20049,N_20819);
and U24461 (N_24461,N_21951,N_21712);
and U24462 (N_24462,N_21675,N_21953);
nand U24463 (N_24463,N_20308,N_20779);
or U24464 (N_24464,N_20856,N_20135);
nor U24465 (N_24465,N_20543,N_20299);
xor U24466 (N_24466,N_21665,N_20566);
nand U24467 (N_24467,N_21008,N_21659);
nand U24468 (N_24468,N_21351,N_20035);
or U24469 (N_24469,N_21559,N_21640);
nand U24470 (N_24470,N_20214,N_21296);
or U24471 (N_24471,N_22071,N_21282);
and U24472 (N_24472,N_20586,N_21928);
nor U24473 (N_24473,N_20376,N_20977);
xor U24474 (N_24474,N_21793,N_22356);
nand U24475 (N_24475,N_21978,N_21358);
nand U24476 (N_24476,N_22432,N_22428);
and U24477 (N_24477,N_22211,N_20250);
nand U24478 (N_24478,N_21631,N_20474);
nand U24479 (N_24479,N_21100,N_20291);
nor U24480 (N_24480,N_21522,N_20709);
xor U24481 (N_24481,N_20318,N_20285);
nor U24482 (N_24482,N_21525,N_22116);
or U24483 (N_24483,N_21861,N_20422);
nand U24484 (N_24484,N_20304,N_20801);
or U24485 (N_24485,N_21448,N_22470);
and U24486 (N_24486,N_22027,N_22078);
and U24487 (N_24487,N_22067,N_22486);
and U24488 (N_24488,N_21228,N_20502);
and U24489 (N_24489,N_22039,N_22370);
nor U24490 (N_24490,N_21990,N_21433);
xor U24491 (N_24491,N_22312,N_20640);
xor U24492 (N_24492,N_20406,N_22301);
and U24493 (N_24493,N_20598,N_21636);
and U24494 (N_24494,N_20760,N_20651);
or U24495 (N_24495,N_22485,N_20443);
nor U24496 (N_24496,N_22171,N_21337);
xnor U24497 (N_24497,N_20493,N_21121);
or U24498 (N_24498,N_22125,N_20593);
nand U24499 (N_24499,N_22340,N_21875);
and U24500 (N_24500,N_20881,N_22077);
nor U24501 (N_24501,N_20391,N_22202);
nor U24502 (N_24502,N_20778,N_20491);
or U24503 (N_24503,N_21458,N_20424);
nand U24504 (N_24504,N_21857,N_20847);
xnor U24505 (N_24505,N_20072,N_20619);
nor U24506 (N_24506,N_20013,N_20850);
nand U24507 (N_24507,N_20435,N_22280);
xor U24508 (N_24508,N_20597,N_22395);
xnor U24509 (N_24509,N_21190,N_21030);
nand U24510 (N_24510,N_21043,N_21544);
nand U24511 (N_24511,N_20406,N_20998);
nand U24512 (N_24512,N_21560,N_20319);
nand U24513 (N_24513,N_21146,N_21086);
or U24514 (N_24514,N_20516,N_20512);
nand U24515 (N_24515,N_21835,N_20672);
xor U24516 (N_24516,N_21633,N_21708);
nor U24517 (N_24517,N_20145,N_22053);
and U24518 (N_24518,N_20684,N_21375);
or U24519 (N_24519,N_20428,N_20062);
xnor U24520 (N_24520,N_22003,N_20573);
xor U24521 (N_24521,N_20241,N_20219);
nor U24522 (N_24522,N_20850,N_21398);
nand U24523 (N_24523,N_20374,N_20688);
or U24524 (N_24524,N_21008,N_21690);
or U24525 (N_24525,N_21772,N_20142);
xor U24526 (N_24526,N_22008,N_20275);
and U24527 (N_24527,N_20105,N_20040);
xnor U24528 (N_24528,N_21998,N_20251);
nand U24529 (N_24529,N_22171,N_21693);
xnor U24530 (N_24530,N_22109,N_20200);
or U24531 (N_24531,N_21031,N_22246);
nand U24532 (N_24532,N_20279,N_22028);
and U24533 (N_24533,N_20221,N_22418);
and U24534 (N_24534,N_20474,N_22151);
nor U24535 (N_24535,N_22157,N_22418);
or U24536 (N_24536,N_20811,N_21854);
xnor U24537 (N_24537,N_21485,N_21559);
nand U24538 (N_24538,N_20658,N_20052);
xnor U24539 (N_24539,N_21546,N_20011);
or U24540 (N_24540,N_20872,N_20540);
nand U24541 (N_24541,N_22480,N_21783);
xor U24542 (N_24542,N_21426,N_22048);
or U24543 (N_24543,N_20716,N_21318);
or U24544 (N_24544,N_20930,N_20765);
nor U24545 (N_24545,N_21868,N_20518);
nor U24546 (N_24546,N_20689,N_20866);
and U24547 (N_24547,N_21037,N_22163);
nor U24548 (N_24548,N_22129,N_21772);
nand U24549 (N_24549,N_21910,N_21387);
xor U24550 (N_24550,N_22457,N_21052);
and U24551 (N_24551,N_20978,N_20966);
or U24552 (N_24552,N_20676,N_20755);
nor U24553 (N_24553,N_20293,N_20549);
nor U24554 (N_24554,N_20919,N_20478);
nand U24555 (N_24555,N_20170,N_21451);
nand U24556 (N_24556,N_20197,N_20040);
nor U24557 (N_24557,N_20707,N_20261);
xor U24558 (N_24558,N_21374,N_20288);
xnor U24559 (N_24559,N_21626,N_21645);
nand U24560 (N_24560,N_21246,N_21143);
or U24561 (N_24561,N_21980,N_20983);
xor U24562 (N_24562,N_21573,N_21132);
nand U24563 (N_24563,N_21717,N_21137);
nor U24564 (N_24564,N_21710,N_22069);
or U24565 (N_24565,N_20476,N_20761);
or U24566 (N_24566,N_21895,N_21162);
xor U24567 (N_24567,N_22389,N_21768);
and U24568 (N_24568,N_20004,N_21051);
and U24569 (N_24569,N_21491,N_20649);
nand U24570 (N_24570,N_20087,N_21305);
xnor U24571 (N_24571,N_21898,N_21091);
or U24572 (N_24572,N_20630,N_21895);
or U24573 (N_24573,N_20068,N_21062);
xnor U24574 (N_24574,N_20092,N_22028);
xnor U24575 (N_24575,N_20526,N_20708);
nand U24576 (N_24576,N_20367,N_21559);
or U24577 (N_24577,N_20192,N_21256);
xor U24578 (N_24578,N_20714,N_21084);
nor U24579 (N_24579,N_22165,N_20496);
nand U24580 (N_24580,N_22295,N_20604);
nand U24581 (N_24581,N_20271,N_21772);
xor U24582 (N_24582,N_20044,N_22285);
xor U24583 (N_24583,N_22072,N_20279);
xnor U24584 (N_24584,N_21133,N_20761);
and U24585 (N_24585,N_20720,N_20267);
or U24586 (N_24586,N_21071,N_21760);
xor U24587 (N_24587,N_21447,N_21049);
nand U24588 (N_24588,N_21316,N_20200);
nand U24589 (N_24589,N_20212,N_20585);
and U24590 (N_24590,N_21391,N_22462);
and U24591 (N_24591,N_21428,N_21463);
or U24592 (N_24592,N_21621,N_20506);
or U24593 (N_24593,N_21413,N_22292);
or U24594 (N_24594,N_20886,N_20157);
nand U24595 (N_24595,N_20487,N_20875);
xnor U24596 (N_24596,N_21501,N_20207);
nand U24597 (N_24597,N_20866,N_20928);
or U24598 (N_24598,N_20573,N_21740);
and U24599 (N_24599,N_22046,N_21070);
and U24600 (N_24600,N_21692,N_21135);
nor U24601 (N_24601,N_22464,N_21146);
nor U24602 (N_24602,N_22034,N_21358);
or U24603 (N_24603,N_21814,N_22468);
nor U24604 (N_24604,N_21589,N_22346);
nand U24605 (N_24605,N_22473,N_22117);
nor U24606 (N_24606,N_20055,N_22007);
nor U24607 (N_24607,N_21130,N_20354);
xor U24608 (N_24608,N_22489,N_21476);
nand U24609 (N_24609,N_21125,N_22373);
nand U24610 (N_24610,N_21651,N_22038);
and U24611 (N_24611,N_20637,N_22319);
nand U24612 (N_24612,N_21962,N_21148);
nand U24613 (N_24613,N_20773,N_21465);
or U24614 (N_24614,N_21227,N_22443);
xor U24615 (N_24615,N_22242,N_20984);
nor U24616 (N_24616,N_20366,N_21349);
xor U24617 (N_24617,N_20662,N_21160);
xnor U24618 (N_24618,N_20872,N_20906);
xnor U24619 (N_24619,N_20834,N_20581);
or U24620 (N_24620,N_22239,N_20347);
nand U24621 (N_24621,N_20550,N_21954);
and U24622 (N_24622,N_20142,N_21032);
or U24623 (N_24623,N_21315,N_22010);
nand U24624 (N_24624,N_20932,N_20558);
nor U24625 (N_24625,N_20091,N_20295);
nand U24626 (N_24626,N_21725,N_20583);
nand U24627 (N_24627,N_21327,N_21357);
or U24628 (N_24628,N_20365,N_21740);
xnor U24629 (N_24629,N_21044,N_21798);
and U24630 (N_24630,N_21071,N_22396);
nor U24631 (N_24631,N_21474,N_21795);
nor U24632 (N_24632,N_21727,N_21161);
or U24633 (N_24633,N_20185,N_20225);
and U24634 (N_24634,N_21622,N_21760);
xnor U24635 (N_24635,N_20175,N_21246);
xor U24636 (N_24636,N_20344,N_21972);
or U24637 (N_24637,N_21019,N_20053);
nand U24638 (N_24638,N_21923,N_21553);
nor U24639 (N_24639,N_21123,N_21144);
nand U24640 (N_24640,N_20167,N_20605);
or U24641 (N_24641,N_22272,N_22385);
and U24642 (N_24642,N_20107,N_21662);
and U24643 (N_24643,N_21544,N_20365);
nor U24644 (N_24644,N_21961,N_20853);
or U24645 (N_24645,N_21759,N_21847);
nor U24646 (N_24646,N_21144,N_22402);
nand U24647 (N_24647,N_22119,N_21774);
and U24648 (N_24648,N_20570,N_21243);
nor U24649 (N_24649,N_20390,N_21008);
nor U24650 (N_24650,N_21356,N_21480);
or U24651 (N_24651,N_22079,N_21538);
and U24652 (N_24652,N_20089,N_20543);
nand U24653 (N_24653,N_20315,N_20431);
and U24654 (N_24654,N_21848,N_22278);
and U24655 (N_24655,N_20379,N_21342);
xnor U24656 (N_24656,N_21653,N_21830);
and U24657 (N_24657,N_22388,N_20416);
and U24658 (N_24658,N_20673,N_21188);
nor U24659 (N_24659,N_22285,N_22189);
nand U24660 (N_24660,N_21486,N_22071);
xnor U24661 (N_24661,N_21715,N_20279);
xor U24662 (N_24662,N_20733,N_21786);
xor U24663 (N_24663,N_21563,N_20166);
and U24664 (N_24664,N_22042,N_21415);
or U24665 (N_24665,N_20807,N_20097);
xor U24666 (N_24666,N_21686,N_21194);
xnor U24667 (N_24667,N_21683,N_20866);
nor U24668 (N_24668,N_20493,N_20861);
and U24669 (N_24669,N_21464,N_21160);
xor U24670 (N_24670,N_20649,N_20374);
nor U24671 (N_24671,N_20311,N_20567);
or U24672 (N_24672,N_21774,N_20451);
or U24673 (N_24673,N_21500,N_20529);
and U24674 (N_24674,N_20728,N_21838);
xnor U24675 (N_24675,N_20395,N_20272);
nor U24676 (N_24676,N_21718,N_20101);
nand U24677 (N_24677,N_20635,N_20895);
xor U24678 (N_24678,N_20836,N_20593);
nor U24679 (N_24679,N_21249,N_21965);
nor U24680 (N_24680,N_22147,N_20336);
nor U24681 (N_24681,N_22261,N_21671);
nor U24682 (N_24682,N_20894,N_21864);
or U24683 (N_24683,N_20730,N_20747);
and U24684 (N_24684,N_22297,N_20789);
xnor U24685 (N_24685,N_20620,N_20780);
or U24686 (N_24686,N_20935,N_20379);
nand U24687 (N_24687,N_21696,N_20662);
nand U24688 (N_24688,N_21291,N_20312);
xor U24689 (N_24689,N_20370,N_20546);
nor U24690 (N_24690,N_20663,N_20619);
and U24691 (N_24691,N_21118,N_21063);
nand U24692 (N_24692,N_20063,N_22490);
or U24693 (N_24693,N_21838,N_20791);
nand U24694 (N_24694,N_21343,N_21339);
xnor U24695 (N_24695,N_21345,N_21203);
nor U24696 (N_24696,N_20700,N_20964);
and U24697 (N_24697,N_22120,N_20143);
nor U24698 (N_24698,N_20067,N_20543);
and U24699 (N_24699,N_20891,N_21407);
or U24700 (N_24700,N_21803,N_20793);
xor U24701 (N_24701,N_20562,N_20226);
nor U24702 (N_24702,N_20361,N_21186);
and U24703 (N_24703,N_20503,N_20903);
nor U24704 (N_24704,N_20859,N_22129);
nand U24705 (N_24705,N_20982,N_20492);
nor U24706 (N_24706,N_20506,N_21507);
nand U24707 (N_24707,N_21540,N_20424);
and U24708 (N_24708,N_22461,N_21704);
or U24709 (N_24709,N_21566,N_20993);
or U24710 (N_24710,N_22346,N_21471);
xnor U24711 (N_24711,N_20708,N_22243);
xnor U24712 (N_24712,N_21133,N_20178);
nor U24713 (N_24713,N_22323,N_22261);
or U24714 (N_24714,N_20684,N_21527);
and U24715 (N_24715,N_21719,N_21528);
and U24716 (N_24716,N_21032,N_22380);
or U24717 (N_24717,N_21792,N_20697);
nor U24718 (N_24718,N_20572,N_22209);
nor U24719 (N_24719,N_21317,N_22201);
xor U24720 (N_24720,N_22001,N_20448);
nor U24721 (N_24721,N_21794,N_21947);
or U24722 (N_24722,N_21955,N_22486);
xnor U24723 (N_24723,N_20170,N_21047);
nor U24724 (N_24724,N_21134,N_21055);
nand U24725 (N_24725,N_20080,N_20361);
nor U24726 (N_24726,N_21840,N_22184);
xnor U24727 (N_24727,N_20081,N_20303);
nand U24728 (N_24728,N_22026,N_22257);
xor U24729 (N_24729,N_20982,N_22146);
and U24730 (N_24730,N_22396,N_20440);
nor U24731 (N_24731,N_22475,N_20423);
or U24732 (N_24732,N_20141,N_22172);
xor U24733 (N_24733,N_22263,N_20110);
nand U24734 (N_24734,N_22307,N_22291);
and U24735 (N_24735,N_20836,N_22110);
or U24736 (N_24736,N_22076,N_22024);
xor U24737 (N_24737,N_20081,N_20654);
nor U24738 (N_24738,N_20383,N_21420);
xnor U24739 (N_24739,N_21251,N_22199);
nor U24740 (N_24740,N_20779,N_20735);
nand U24741 (N_24741,N_20033,N_20797);
xnor U24742 (N_24742,N_20823,N_21473);
nor U24743 (N_24743,N_21850,N_20366);
nor U24744 (N_24744,N_21641,N_22291);
nor U24745 (N_24745,N_22473,N_22415);
xnor U24746 (N_24746,N_20044,N_22107);
or U24747 (N_24747,N_20799,N_20631);
or U24748 (N_24748,N_21654,N_21972);
nand U24749 (N_24749,N_21742,N_22462);
xnor U24750 (N_24750,N_21365,N_21680);
nand U24751 (N_24751,N_22439,N_21787);
and U24752 (N_24752,N_21469,N_21010);
or U24753 (N_24753,N_21613,N_22353);
nand U24754 (N_24754,N_20153,N_20067);
xnor U24755 (N_24755,N_20209,N_21784);
or U24756 (N_24756,N_20916,N_22366);
nor U24757 (N_24757,N_21094,N_20681);
or U24758 (N_24758,N_21192,N_20151);
or U24759 (N_24759,N_22397,N_21091);
xor U24760 (N_24760,N_20970,N_21875);
xor U24761 (N_24761,N_21036,N_22148);
xor U24762 (N_24762,N_20059,N_20734);
xor U24763 (N_24763,N_20965,N_21347);
and U24764 (N_24764,N_20657,N_21632);
and U24765 (N_24765,N_20477,N_21977);
nand U24766 (N_24766,N_20039,N_20622);
xor U24767 (N_24767,N_20995,N_21916);
nand U24768 (N_24768,N_20968,N_22301);
or U24769 (N_24769,N_20728,N_20334);
nand U24770 (N_24770,N_22297,N_22329);
xor U24771 (N_24771,N_20069,N_20484);
and U24772 (N_24772,N_20081,N_22428);
nand U24773 (N_24773,N_20386,N_20004);
and U24774 (N_24774,N_22094,N_20535);
xor U24775 (N_24775,N_20458,N_21889);
nor U24776 (N_24776,N_22410,N_20283);
xor U24777 (N_24777,N_20154,N_21469);
nand U24778 (N_24778,N_20096,N_20230);
and U24779 (N_24779,N_22096,N_21983);
xor U24780 (N_24780,N_22270,N_20534);
or U24781 (N_24781,N_21976,N_21554);
xnor U24782 (N_24782,N_20592,N_21651);
and U24783 (N_24783,N_21974,N_20131);
nand U24784 (N_24784,N_21356,N_20845);
nand U24785 (N_24785,N_21741,N_20192);
xnor U24786 (N_24786,N_20407,N_20657);
or U24787 (N_24787,N_21191,N_20719);
or U24788 (N_24788,N_20232,N_20385);
xnor U24789 (N_24789,N_21808,N_20778);
or U24790 (N_24790,N_20027,N_21074);
xor U24791 (N_24791,N_20485,N_22374);
nor U24792 (N_24792,N_21482,N_20376);
xnor U24793 (N_24793,N_22415,N_21654);
and U24794 (N_24794,N_21961,N_21370);
or U24795 (N_24795,N_22462,N_21368);
nor U24796 (N_24796,N_20284,N_22049);
or U24797 (N_24797,N_20541,N_21488);
nand U24798 (N_24798,N_22345,N_21862);
and U24799 (N_24799,N_21244,N_20627);
and U24800 (N_24800,N_20096,N_21430);
or U24801 (N_24801,N_21411,N_20726);
nand U24802 (N_24802,N_22031,N_20783);
or U24803 (N_24803,N_21322,N_22452);
or U24804 (N_24804,N_20021,N_21015);
nand U24805 (N_24805,N_20526,N_21142);
nor U24806 (N_24806,N_21452,N_20422);
or U24807 (N_24807,N_21631,N_21496);
nand U24808 (N_24808,N_22137,N_21355);
xnor U24809 (N_24809,N_22154,N_20968);
nand U24810 (N_24810,N_20864,N_21794);
xor U24811 (N_24811,N_21038,N_22156);
nand U24812 (N_24812,N_22263,N_20764);
and U24813 (N_24813,N_22137,N_21522);
nand U24814 (N_24814,N_20745,N_20877);
xor U24815 (N_24815,N_21193,N_20788);
nor U24816 (N_24816,N_20519,N_21391);
xnor U24817 (N_24817,N_22129,N_21166);
nand U24818 (N_24818,N_20236,N_20442);
nor U24819 (N_24819,N_21391,N_22482);
and U24820 (N_24820,N_21925,N_20499);
nand U24821 (N_24821,N_21685,N_20259);
nand U24822 (N_24822,N_21932,N_20525);
xnor U24823 (N_24823,N_22414,N_20028);
nand U24824 (N_24824,N_21541,N_20881);
or U24825 (N_24825,N_21618,N_21529);
or U24826 (N_24826,N_21379,N_20379);
xnor U24827 (N_24827,N_20172,N_21424);
or U24828 (N_24828,N_22022,N_21570);
nand U24829 (N_24829,N_22265,N_22340);
and U24830 (N_24830,N_21652,N_21088);
nand U24831 (N_24831,N_21919,N_22067);
xnor U24832 (N_24832,N_21123,N_20878);
nand U24833 (N_24833,N_21129,N_22374);
nor U24834 (N_24834,N_21625,N_20899);
nor U24835 (N_24835,N_22228,N_20988);
xnor U24836 (N_24836,N_20957,N_20385);
nor U24837 (N_24837,N_20668,N_21690);
nand U24838 (N_24838,N_21689,N_21628);
or U24839 (N_24839,N_22248,N_20581);
or U24840 (N_24840,N_20012,N_21603);
and U24841 (N_24841,N_20773,N_21665);
and U24842 (N_24842,N_22398,N_20232);
or U24843 (N_24843,N_20357,N_22350);
and U24844 (N_24844,N_20767,N_21593);
or U24845 (N_24845,N_22233,N_21499);
nor U24846 (N_24846,N_22463,N_21777);
nand U24847 (N_24847,N_21912,N_21330);
nor U24848 (N_24848,N_21127,N_22136);
nor U24849 (N_24849,N_21089,N_22274);
nand U24850 (N_24850,N_22185,N_20192);
and U24851 (N_24851,N_21462,N_21114);
nand U24852 (N_24852,N_21359,N_20042);
nand U24853 (N_24853,N_20144,N_21471);
and U24854 (N_24854,N_20528,N_20998);
nand U24855 (N_24855,N_20830,N_21170);
nor U24856 (N_24856,N_20586,N_21763);
nand U24857 (N_24857,N_21167,N_21537);
nor U24858 (N_24858,N_20939,N_22170);
or U24859 (N_24859,N_20050,N_21108);
xor U24860 (N_24860,N_21261,N_20423);
and U24861 (N_24861,N_20155,N_21631);
and U24862 (N_24862,N_20430,N_21652);
xor U24863 (N_24863,N_21524,N_21027);
nor U24864 (N_24864,N_22309,N_20863);
xnor U24865 (N_24865,N_20337,N_21379);
nand U24866 (N_24866,N_21732,N_20316);
and U24867 (N_24867,N_22055,N_20130);
and U24868 (N_24868,N_21022,N_21906);
nand U24869 (N_24869,N_20456,N_22434);
and U24870 (N_24870,N_21593,N_20683);
nand U24871 (N_24871,N_20133,N_21608);
xnor U24872 (N_24872,N_20074,N_22329);
or U24873 (N_24873,N_21535,N_21868);
nor U24874 (N_24874,N_20842,N_21121);
or U24875 (N_24875,N_22202,N_21626);
xnor U24876 (N_24876,N_20314,N_21743);
nor U24877 (N_24877,N_20958,N_20399);
or U24878 (N_24878,N_21185,N_20313);
and U24879 (N_24879,N_20639,N_20372);
xnor U24880 (N_24880,N_22323,N_22418);
nand U24881 (N_24881,N_20523,N_21859);
nand U24882 (N_24882,N_21336,N_20202);
and U24883 (N_24883,N_22013,N_21368);
xor U24884 (N_24884,N_22232,N_21761);
nand U24885 (N_24885,N_22407,N_22011);
nor U24886 (N_24886,N_20115,N_21484);
xnor U24887 (N_24887,N_21928,N_20365);
xor U24888 (N_24888,N_21974,N_21108);
nand U24889 (N_24889,N_22474,N_21959);
nand U24890 (N_24890,N_21465,N_20210);
and U24891 (N_24891,N_20663,N_20922);
nor U24892 (N_24892,N_20251,N_20603);
nor U24893 (N_24893,N_20900,N_20123);
nor U24894 (N_24894,N_22091,N_20117);
nor U24895 (N_24895,N_22473,N_20193);
xnor U24896 (N_24896,N_22489,N_21815);
or U24897 (N_24897,N_21813,N_20837);
nand U24898 (N_24898,N_22175,N_22404);
xor U24899 (N_24899,N_21942,N_20497);
and U24900 (N_24900,N_20546,N_20143);
or U24901 (N_24901,N_22231,N_21204);
xnor U24902 (N_24902,N_20290,N_20362);
nor U24903 (N_24903,N_21554,N_21741);
or U24904 (N_24904,N_20309,N_20660);
and U24905 (N_24905,N_21812,N_21769);
and U24906 (N_24906,N_21364,N_21785);
nand U24907 (N_24907,N_21198,N_22119);
or U24908 (N_24908,N_20559,N_20569);
or U24909 (N_24909,N_21262,N_22392);
nand U24910 (N_24910,N_20813,N_20750);
nand U24911 (N_24911,N_21674,N_22292);
nand U24912 (N_24912,N_20384,N_20530);
xnor U24913 (N_24913,N_22353,N_22268);
or U24914 (N_24914,N_22168,N_20147);
and U24915 (N_24915,N_21595,N_21268);
and U24916 (N_24916,N_21308,N_21251);
nor U24917 (N_24917,N_21419,N_20334);
nor U24918 (N_24918,N_21594,N_21258);
xnor U24919 (N_24919,N_20411,N_21424);
nand U24920 (N_24920,N_21705,N_22147);
nor U24921 (N_24921,N_21897,N_20798);
nand U24922 (N_24922,N_20891,N_20390);
or U24923 (N_24923,N_20733,N_20454);
xnor U24924 (N_24924,N_21824,N_22310);
xnor U24925 (N_24925,N_20024,N_21842);
xnor U24926 (N_24926,N_20448,N_21049);
nor U24927 (N_24927,N_22072,N_22362);
or U24928 (N_24928,N_21381,N_20214);
nor U24929 (N_24929,N_21768,N_21893);
nand U24930 (N_24930,N_20342,N_21388);
nor U24931 (N_24931,N_20071,N_21402);
nor U24932 (N_24932,N_20422,N_22400);
or U24933 (N_24933,N_20402,N_20841);
nand U24934 (N_24934,N_21834,N_20502);
nor U24935 (N_24935,N_21082,N_22040);
nand U24936 (N_24936,N_22183,N_21292);
or U24937 (N_24937,N_22466,N_20600);
nor U24938 (N_24938,N_22184,N_20575);
xnor U24939 (N_24939,N_21605,N_20721);
or U24940 (N_24940,N_22256,N_20939);
nand U24941 (N_24941,N_21489,N_22343);
xnor U24942 (N_24942,N_21059,N_20388);
nor U24943 (N_24943,N_20851,N_21820);
nor U24944 (N_24944,N_22421,N_22383);
and U24945 (N_24945,N_20865,N_21134);
or U24946 (N_24946,N_20031,N_21999);
nor U24947 (N_24947,N_21320,N_20683);
xnor U24948 (N_24948,N_21790,N_21758);
nand U24949 (N_24949,N_21900,N_22086);
and U24950 (N_24950,N_20667,N_21602);
nor U24951 (N_24951,N_22111,N_22034);
xor U24952 (N_24952,N_21683,N_20752);
or U24953 (N_24953,N_20829,N_20865);
and U24954 (N_24954,N_20429,N_20433);
and U24955 (N_24955,N_20816,N_22310);
or U24956 (N_24956,N_20368,N_22463);
nor U24957 (N_24957,N_21251,N_20329);
or U24958 (N_24958,N_21425,N_20364);
nand U24959 (N_24959,N_22440,N_20192);
and U24960 (N_24960,N_22008,N_21595);
and U24961 (N_24961,N_20512,N_20326);
nor U24962 (N_24962,N_21945,N_20834);
and U24963 (N_24963,N_20458,N_21017);
or U24964 (N_24964,N_21908,N_20664);
nor U24965 (N_24965,N_21755,N_21542);
nand U24966 (N_24966,N_21875,N_21853);
xnor U24967 (N_24967,N_20727,N_21688);
or U24968 (N_24968,N_22451,N_21476);
and U24969 (N_24969,N_21532,N_21039);
and U24970 (N_24970,N_21881,N_21261);
nor U24971 (N_24971,N_21837,N_21628);
xnor U24972 (N_24972,N_21253,N_20668);
and U24973 (N_24973,N_20209,N_20624);
nor U24974 (N_24974,N_20414,N_21911);
or U24975 (N_24975,N_21507,N_22380);
nand U24976 (N_24976,N_22063,N_20767);
or U24977 (N_24977,N_22106,N_21305);
or U24978 (N_24978,N_22171,N_22183);
nor U24979 (N_24979,N_20452,N_20394);
nand U24980 (N_24980,N_21997,N_20408);
xnor U24981 (N_24981,N_21621,N_21107);
or U24982 (N_24982,N_21814,N_21377);
nand U24983 (N_24983,N_21744,N_21756);
nor U24984 (N_24984,N_21607,N_21340);
nand U24985 (N_24985,N_21456,N_20526);
or U24986 (N_24986,N_22293,N_22398);
nor U24987 (N_24987,N_21223,N_21881);
xnor U24988 (N_24988,N_20907,N_20271);
and U24989 (N_24989,N_20928,N_22048);
or U24990 (N_24990,N_20883,N_20642);
and U24991 (N_24991,N_21537,N_21320);
and U24992 (N_24992,N_21955,N_20238);
nor U24993 (N_24993,N_22257,N_22480);
and U24994 (N_24994,N_21682,N_22093);
and U24995 (N_24995,N_21685,N_21376);
nor U24996 (N_24996,N_20809,N_22055);
or U24997 (N_24997,N_20138,N_21100);
or U24998 (N_24998,N_20407,N_21842);
and U24999 (N_24999,N_20247,N_20468);
xnor UO_0 (O_0,N_24080,N_23887);
xnor UO_1 (O_1,N_23133,N_24611);
xor UO_2 (O_2,N_24746,N_23114);
nor UO_3 (O_3,N_22523,N_22678);
or UO_4 (O_4,N_23246,N_24526);
xor UO_5 (O_5,N_24258,N_23762);
nor UO_6 (O_6,N_24351,N_22725);
nor UO_7 (O_7,N_23351,N_24141);
or UO_8 (O_8,N_23200,N_23863);
xnor UO_9 (O_9,N_24082,N_22676);
or UO_10 (O_10,N_23140,N_22784);
or UO_11 (O_11,N_24578,N_22954);
nor UO_12 (O_12,N_23593,N_22842);
xor UO_13 (O_13,N_24135,N_24548);
nor UO_14 (O_14,N_24888,N_22720);
and UO_15 (O_15,N_22824,N_24992);
xnor UO_16 (O_16,N_23992,N_24843);
xnor UO_17 (O_17,N_23331,N_23987);
and UO_18 (O_18,N_24382,N_23010);
or UO_19 (O_19,N_24534,N_23672);
nand UO_20 (O_20,N_23929,N_23945);
and UO_21 (O_21,N_23067,N_23038);
nand UO_22 (O_22,N_24453,N_23658);
xnor UO_23 (O_23,N_22960,N_22828);
nor UO_24 (O_24,N_23991,N_22592);
and UO_25 (O_25,N_22501,N_24057);
or UO_26 (O_26,N_23306,N_23235);
and UO_27 (O_27,N_24220,N_22922);
xnor UO_28 (O_28,N_24076,N_24620);
xor UO_29 (O_29,N_23746,N_23237);
and UO_30 (O_30,N_23125,N_24879);
nor UO_31 (O_31,N_22950,N_22831);
nand UO_32 (O_32,N_24873,N_23288);
or UO_33 (O_33,N_22779,N_24188);
or UO_34 (O_34,N_23685,N_24416);
nand UO_35 (O_35,N_23305,N_23357);
or UO_36 (O_36,N_24550,N_24538);
nor UO_37 (O_37,N_24431,N_24376);
nand UO_38 (O_38,N_22655,N_23382);
or UO_39 (O_39,N_22743,N_24629);
and UO_40 (O_40,N_22808,N_24711);
nor UO_41 (O_41,N_24657,N_24918);
xor UO_42 (O_42,N_24841,N_24844);
nor UO_43 (O_43,N_24830,N_23142);
or UO_44 (O_44,N_23725,N_23183);
xnor UO_45 (O_45,N_23779,N_23997);
or UO_46 (O_46,N_22812,N_24460);
or UO_47 (O_47,N_23944,N_22846);
nand UO_48 (O_48,N_24506,N_24365);
xnor UO_49 (O_49,N_23961,N_23290);
and UO_50 (O_50,N_23111,N_24591);
and UO_51 (O_51,N_23513,N_22834);
or UO_52 (O_52,N_23749,N_23511);
xnor UO_53 (O_53,N_23708,N_24681);
nand UO_54 (O_54,N_22538,N_23325);
or UO_55 (O_55,N_23555,N_22674);
nor UO_56 (O_56,N_24688,N_23259);
or UO_57 (O_57,N_22794,N_24304);
xor UO_58 (O_58,N_24555,N_22845);
xor UO_59 (O_59,N_24853,N_22543);
or UO_60 (O_60,N_23766,N_24372);
xor UO_61 (O_61,N_24925,N_23374);
nand UO_62 (O_62,N_23247,N_24755);
xnor UO_63 (O_63,N_24329,N_24280);
xor UO_64 (O_64,N_22836,N_24838);
nand UO_65 (O_65,N_24274,N_23633);
xor UO_66 (O_66,N_24763,N_24010);
and UO_67 (O_67,N_23359,N_23248);
or UO_68 (O_68,N_23283,N_23786);
and UO_69 (O_69,N_24923,N_24784);
xnor UO_70 (O_70,N_24997,N_23487);
and UO_71 (O_71,N_24565,N_22588);
and UO_72 (O_72,N_23723,N_24848);
or UO_73 (O_73,N_24725,N_22769);
nand UO_74 (O_74,N_24972,N_22558);
or UO_75 (O_75,N_24263,N_24492);
nor UO_76 (O_76,N_22724,N_23229);
xnor UO_77 (O_77,N_23811,N_22587);
nand UO_78 (O_78,N_24355,N_23320);
or UO_79 (O_79,N_24970,N_23644);
xnor UO_80 (O_80,N_23241,N_22885);
nor UO_81 (O_81,N_22669,N_23315);
nor UO_82 (O_82,N_22618,N_22790);
nand UO_83 (O_83,N_22708,N_24302);
and UO_84 (O_84,N_23437,N_24891);
nand UO_85 (O_85,N_23829,N_23905);
xnor UO_86 (O_86,N_24142,N_23254);
or UO_87 (O_87,N_24562,N_24630);
and UO_88 (O_88,N_23302,N_24227);
nor UO_89 (O_89,N_24648,N_22915);
nand UO_90 (O_90,N_23420,N_24640);
or UO_91 (O_91,N_22946,N_23195);
xor UO_92 (O_92,N_24477,N_24757);
and UO_93 (O_93,N_24101,N_23386);
xnor UO_94 (O_94,N_22966,N_24893);
nand UO_95 (O_95,N_24525,N_24706);
and UO_96 (O_96,N_23457,N_23696);
and UO_97 (O_97,N_23396,N_22536);
and UO_98 (O_98,N_24522,N_23709);
nor UO_99 (O_99,N_22600,N_24267);
and UO_100 (O_100,N_22715,N_23294);
nor UO_101 (O_101,N_23274,N_24641);
and UO_102 (O_102,N_23556,N_24729);
nand UO_103 (O_103,N_24649,N_23323);
xnor UO_104 (O_104,N_23951,N_23353);
xor UO_105 (O_105,N_22874,N_24607);
and UO_106 (O_106,N_24081,N_24249);
and UO_107 (O_107,N_23894,N_24405);
xor UO_108 (O_108,N_24493,N_24250);
nand UO_109 (O_109,N_23406,N_24842);
and UO_110 (O_110,N_23291,N_23980);
and UO_111 (O_111,N_24037,N_24660);
and UO_112 (O_112,N_23415,N_22683);
and UO_113 (O_113,N_23505,N_24875);
nand UO_114 (O_114,N_24087,N_23931);
or UO_115 (O_115,N_23131,N_23895);
xnor UO_116 (O_116,N_23872,N_23604);
nand UO_117 (O_117,N_24732,N_23372);
xor UO_118 (O_118,N_23107,N_24261);
xor UO_119 (O_119,N_24294,N_22728);
and UO_120 (O_120,N_23899,N_23726);
and UO_121 (O_121,N_23673,N_22651);
xor UO_122 (O_122,N_23129,N_23074);
nor UO_123 (O_123,N_22653,N_23682);
nor UO_124 (O_124,N_23733,N_22570);
nor UO_125 (O_125,N_23959,N_22817);
xnor UO_126 (O_126,N_23557,N_24907);
and UO_127 (O_127,N_22502,N_23778);
or UO_128 (O_128,N_23099,N_23871);
or UO_129 (O_129,N_23693,N_24298);
xor UO_130 (O_130,N_23185,N_24066);
nand UO_131 (O_131,N_23212,N_23711);
nor UO_132 (O_132,N_23785,N_23460);
nand UO_133 (O_133,N_24687,N_22519);
or UO_134 (O_134,N_23908,N_24736);
nand UO_135 (O_135,N_22910,N_24117);
nand UO_136 (O_136,N_23023,N_23450);
nand UO_137 (O_137,N_24044,N_24070);
or UO_138 (O_138,N_23047,N_24019);
and UO_139 (O_139,N_24683,N_24960);
or UO_140 (O_140,N_23917,N_23520);
nor UO_141 (O_141,N_24651,N_23958);
nand UO_142 (O_142,N_24001,N_22574);
and UO_143 (O_143,N_22507,N_24028);
and UO_144 (O_144,N_22918,N_24198);
xnor UO_145 (O_145,N_24636,N_22912);
or UO_146 (O_146,N_23414,N_24508);
or UO_147 (O_147,N_22805,N_23289);
and UO_148 (O_148,N_24152,N_24184);
nand UO_149 (O_149,N_23580,N_23238);
xor UO_150 (O_150,N_23928,N_23232);
and UO_151 (O_151,N_24637,N_22888);
and UO_152 (O_152,N_23950,N_24828);
xnor UO_153 (O_153,N_24935,N_24946);
and UO_154 (O_154,N_23497,N_23541);
nor UO_155 (O_155,N_23190,N_24476);
nor UO_156 (O_156,N_23239,N_24664);
xnor UO_157 (O_157,N_24475,N_23592);
xor UO_158 (O_158,N_23692,N_23857);
and UO_159 (O_159,N_23105,N_22907);
nand UO_160 (O_160,N_22762,N_22899);
and UO_161 (O_161,N_22613,N_24390);
and UO_162 (O_162,N_23341,N_23228);
or UO_163 (O_163,N_24443,N_23081);
xor UO_164 (O_164,N_23268,N_23122);
nand UO_165 (O_165,N_24452,N_24074);
or UO_166 (O_166,N_22654,N_23085);
nor UO_167 (O_167,N_23255,N_23002);
nor UO_168 (O_168,N_23157,N_23270);
and UO_169 (O_169,N_24916,N_23784);
xor UO_170 (O_170,N_24332,N_23724);
or UO_171 (O_171,N_24932,N_24507);
or UO_172 (O_172,N_22705,N_22857);
xor UO_173 (O_173,N_23399,N_22598);
nand UO_174 (O_174,N_22809,N_22756);
nand UO_175 (O_175,N_24344,N_24943);
nor UO_176 (O_176,N_23418,N_22897);
and UO_177 (O_177,N_22826,N_24265);
or UO_178 (O_178,N_23301,N_24197);
xnor UO_179 (O_179,N_22871,N_23831);
xnor UO_180 (O_180,N_24792,N_24287);
nand UO_181 (O_181,N_22689,N_24697);
and UO_182 (O_182,N_23595,N_24387);
or UO_183 (O_183,N_22554,N_23751);
and UO_184 (O_184,N_24845,N_23060);
or UO_185 (O_185,N_23594,N_23205);
and UO_186 (O_186,N_22994,N_23411);
and UO_187 (O_187,N_22898,N_22657);
nor UO_188 (O_188,N_24223,N_23702);
or UO_189 (O_189,N_22890,N_24446);
and UO_190 (O_190,N_22594,N_22503);
and UO_191 (O_191,N_24791,N_24404);
and UO_192 (O_192,N_23806,N_23888);
nor UO_193 (O_193,N_23988,N_22564);
or UO_194 (O_194,N_24759,N_24361);
and UO_195 (O_195,N_22636,N_24377);
and UO_196 (O_196,N_24635,N_23001);
xnor UO_197 (O_197,N_24088,N_23168);
nor UO_198 (O_198,N_22546,N_23677);
and UO_199 (O_199,N_23510,N_23271);
xor UO_200 (O_200,N_23083,N_23752);
nand UO_201 (O_201,N_24426,N_24084);
nor UO_202 (O_202,N_24487,N_23518);
nand UO_203 (O_203,N_23665,N_23130);
xnor UO_204 (O_204,N_24724,N_22952);
or UO_205 (O_205,N_22962,N_23602);
nor UO_206 (O_206,N_22516,N_23155);
or UO_207 (O_207,N_24608,N_23890);
and UO_208 (O_208,N_24680,N_23451);
nor UO_209 (O_209,N_24979,N_24642);
or UO_210 (O_210,N_24721,N_24085);
nor UO_211 (O_211,N_22611,N_24872);
xor UO_212 (O_212,N_22601,N_24991);
nor UO_213 (O_213,N_23777,N_24574);
nor UO_214 (O_214,N_24345,N_23470);
nor UO_215 (O_215,N_23879,N_23041);
xor UO_216 (O_216,N_23935,N_23421);
xor UO_217 (O_217,N_24439,N_22512);
nor UO_218 (O_218,N_24586,N_23027);
nand UO_219 (O_219,N_23030,N_24465);
nor UO_220 (O_220,N_23833,N_22875);
nor UO_221 (O_221,N_24868,N_22850);
and UO_222 (O_222,N_24260,N_23071);
nor UO_223 (O_223,N_24884,N_24469);
and UO_224 (O_224,N_24285,N_23953);
nor UO_225 (O_225,N_23536,N_22688);
and UO_226 (O_226,N_23496,N_24108);
xnor UO_227 (O_227,N_24617,N_23612);
nand UO_228 (O_228,N_22742,N_24900);
or UO_229 (O_229,N_23109,N_22518);
nand UO_230 (O_230,N_22620,N_23407);
xnor UO_231 (O_231,N_22729,N_22855);
nand UO_232 (O_232,N_22623,N_23793);
nand UO_233 (O_233,N_24708,N_24251);
or UO_234 (O_234,N_24031,N_23461);
nand UO_235 (O_235,N_24598,N_24097);
xor UO_236 (O_236,N_23443,N_24941);
nand UO_237 (O_237,N_23387,N_24005);
nand UO_238 (O_238,N_23919,N_23150);
nand UO_239 (O_239,N_24034,N_22643);
xor UO_240 (O_240,N_22837,N_22926);
and UO_241 (O_241,N_23990,N_23734);
or UO_242 (O_242,N_23982,N_24324);
nor UO_243 (O_243,N_24145,N_22632);
or UO_244 (O_244,N_22860,N_24363);
and UO_245 (O_245,N_23389,N_22813);
or UO_246 (O_246,N_24275,N_24600);
nor UO_247 (O_247,N_23456,N_23492);
nor UO_248 (O_248,N_24038,N_24381);
nand UO_249 (O_249,N_24413,N_22977);
xnor UO_250 (O_250,N_24758,N_22872);
or UO_251 (O_251,N_23732,N_23203);
xor UO_252 (O_252,N_24242,N_23827);
nand UO_253 (O_253,N_24071,N_24004);
nand UO_254 (O_254,N_24549,N_24911);
nor UO_255 (O_255,N_22789,N_23020);
nand UO_256 (O_256,N_24110,N_22883);
or UO_257 (O_257,N_23966,N_24012);
and UO_258 (O_258,N_22747,N_24962);
nand UO_259 (O_259,N_22895,N_24560);
nor UO_260 (O_260,N_23812,N_23661);
xor UO_261 (O_261,N_23787,N_23075);
xor UO_262 (O_262,N_24462,N_23159);
or UO_263 (O_263,N_22555,N_24839);
xnor UO_264 (O_264,N_22917,N_24384);
and UO_265 (O_265,N_23652,N_22886);
or UO_266 (O_266,N_22989,N_22755);
and UO_267 (O_267,N_23930,N_24217);
xnor UO_268 (O_268,N_24064,N_22644);
nor UO_269 (O_269,N_24334,N_24221);
nor UO_270 (O_270,N_24222,N_23098);
or UO_271 (O_271,N_22510,N_23610);
or UO_272 (O_272,N_23675,N_22741);
and UO_273 (O_273,N_24335,N_24995);
nand UO_274 (O_274,N_23574,N_24908);
nor UO_275 (O_275,N_24890,N_24238);
or UO_276 (O_276,N_24824,N_24113);
nor UO_277 (O_277,N_23586,N_24816);
nor UO_278 (O_278,N_24394,N_24429);
xnor UO_279 (O_279,N_24726,N_24621);
nor UO_280 (O_280,N_24581,N_24051);
and UO_281 (O_281,N_23120,N_24350);
nand UO_282 (O_282,N_24160,N_23668);
xnor UO_283 (O_283,N_23713,N_22616);
and UO_284 (O_284,N_22707,N_24914);
or UO_285 (O_285,N_22983,N_24825);
nand UO_286 (O_286,N_24318,N_22569);
xor UO_287 (O_287,N_23838,N_22854);
nand UO_288 (O_288,N_23840,N_24449);
and UO_289 (O_289,N_23458,N_24107);
or UO_290 (O_290,N_24819,N_23576);
xor UO_291 (O_291,N_24322,N_24194);
and UO_292 (O_292,N_24667,N_23646);
or UO_293 (O_293,N_23442,N_24437);
nand UO_294 (O_294,N_22691,N_23172);
nand UO_295 (O_295,N_24389,N_24986);
nand UO_296 (O_296,N_24418,N_24849);
nor UO_297 (O_297,N_24073,N_22740);
nand UO_298 (O_298,N_22722,N_24112);
nor UO_299 (O_299,N_23334,N_22582);
xnor UO_300 (O_300,N_23759,N_22819);
or UO_301 (O_301,N_24360,N_23329);
nor UO_302 (O_302,N_24055,N_23921);
or UO_303 (O_303,N_24472,N_24403);
nor UO_304 (O_304,N_23662,N_23321);
xnor UO_305 (O_305,N_23391,N_23710);
nand UO_306 (O_306,N_22648,N_24720);
nand UO_307 (O_307,N_24915,N_22619);
nand UO_308 (O_308,N_24132,N_23589);
nor UO_309 (O_309,N_23358,N_22816);
or UO_310 (O_310,N_24502,N_24357);
or UO_311 (O_311,N_24447,N_22701);
nor UO_312 (O_312,N_23554,N_24366);
xor UO_313 (O_313,N_24775,N_24597);
nor UO_314 (O_314,N_24924,N_22635);
or UO_315 (O_315,N_23512,N_22697);
or UO_316 (O_316,N_23490,N_24823);
xnor UO_317 (O_317,N_23163,N_23119);
xor UO_318 (O_318,N_24628,N_24847);
nand UO_319 (O_319,N_23666,N_22630);
or UO_320 (O_320,N_24341,N_24414);
nor UO_321 (O_321,N_24471,N_22903);
nor UO_322 (O_322,N_22757,N_22979);
nand UO_323 (O_323,N_24499,N_22980);
and UO_324 (O_324,N_23342,N_24273);
and UO_325 (O_325,N_22971,N_23210);
xnor UO_326 (O_326,N_23714,N_23836);
nand UO_327 (O_327,N_24068,N_24699);
xnor UO_328 (O_328,N_23043,N_24910);
xor UO_329 (O_329,N_22963,N_24143);
nand UO_330 (O_330,N_23994,N_23715);
xnor UO_331 (O_331,N_24990,N_24735);
nor UO_332 (O_332,N_23346,N_22578);
nand UO_333 (O_333,N_24902,N_24419);
nor UO_334 (O_334,N_23606,N_24407);
or UO_335 (O_335,N_24870,N_23343);
and UO_336 (O_336,N_23467,N_22718);
nor UO_337 (O_337,N_24129,N_24252);
or UO_338 (O_338,N_24086,N_24121);
and UO_339 (O_339,N_22672,N_24645);
or UO_340 (O_340,N_24587,N_23699);
or UO_341 (O_341,N_24148,N_23036);
xnor UO_342 (O_342,N_23138,N_23340);
nand UO_343 (O_343,N_24147,N_24204);
xnor UO_344 (O_344,N_24459,N_23862);
or UO_345 (O_345,N_22716,N_22851);
xnor UO_346 (O_346,N_23565,N_24457);
or UO_347 (O_347,N_22702,N_24386);
and UO_348 (O_348,N_22914,N_22560);
and UO_349 (O_349,N_23638,N_24619);
nand UO_350 (O_350,N_23167,N_23585);
nor UO_351 (O_351,N_22739,N_24211);
nand UO_352 (O_352,N_22717,N_22624);
and UO_353 (O_353,N_23146,N_22690);
xor UO_354 (O_354,N_22995,N_23514);
nor UO_355 (O_355,N_24006,N_22902);
xor UO_356 (O_356,N_23169,N_24500);
nor UO_357 (O_357,N_24430,N_22556);
nor UO_358 (O_358,N_22833,N_24190);
or UO_359 (O_359,N_24488,N_23540);
nor UO_360 (O_360,N_24782,N_23643);
xnor UO_361 (O_361,N_23976,N_23227);
nand UO_362 (O_362,N_24936,N_23128);
or UO_363 (O_363,N_23025,N_24832);
and UO_364 (O_364,N_22736,N_23756);
or UO_365 (O_365,N_23446,N_23145);
nor UO_366 (O_366,N_24676,N_23181);
nor UO_367 (O_367,N_22709,N_22732);
or UO_368 (O_368,N_24594,N_24359);
nand UO_369 (O_369,N_22645,N_24323);
or UO_370 (O_370,N_23940,N_23705);
nand UO_371 (O_371,N_23021,N_22887);
or UO_372 (O_372,N_23077,N_22964);
nor UO_373 (O_373,N_23768,N_23299);
nand UO_374 (O_374,N_24123,N_22581);
or UO_375 (O_375,N_23597,N_23729);
or UO_376 (O_376,N_24177,N_23369);
and UO_377 (O_377,N_23121,N_24903);
and UO_378 (O_378,N_22713,N_22767);
and UO_379 (O_379,N_24632,N_24002);
xnor UO_380 (O_380,N_22792,N_22988);
nand UO_381 (O_381,N_24813,N_23975);
nor UO_382 (O_382,N_24993,N_22776);
xnor UO_383 (O_383,N_24539,N_22770);
or UO_384 (O_384,N_24196,N_24761);
nand UO_385 (O_385,N_23886,N_23765);
nand UO_386 (O_386,N_24138,N_24542);
or UO_387 (O_387,N_23066,N_23250);
xor UO_388 (O_388,N_24569,N_22606);
or UO_389 (O_389,N_24672,N_23230);
xnor UO_390 (O_390,N_23013,N_24599);
xnor UO_391 (O_391,N_23877,N_23376);
and UO_392 (O_392,N_24185,N_24186);
nand UO_393 (O_393,N_24246,N_24650);
and UO_394 (O_394,N_23671,N_23095);
xor UO_395 (O_395,N_23883,N_23267);
and UO_396 (O_396,N_22921,N_22913);
nand UO_397 (O_397,N_22923,N_22684);
xnor UO_398 (O_398,N_24834,N_24480);
or UO_399 (O_399,N_23617,N_24880);
nand UO_400 (O_400,N_22559,N_24279);
nand UO_401 (O_401,N_23932,N_23544);
or UO_402 (O_402,N_23984,N_23681);
nand UO_403 (O_403,N_22524,N_22765);
xor UO_404 (O_404,N_24036,N_23149);
nand UO_405 (O_405,N_24253,N_23689);
nand UO_406 (O_406,N_23654,N_23647);
xnor UO_407 (O_407,N_23375,N_22877);
and UO_408 (O_408,N_23100,N_24510);
and UO_409 (O_409,N_23007,N_23616);
and UO_410 (O_410,N_24235,N_23328);
or UO_411 (O_411,N_23403,N_24815);
and UO_412 (O_412,N_23116,N_24056);
nor UO_413 (O_413,N_23924,N_23719);
nand UO_414 (O_414,N_22766,N_24370);
nand UO_415 (O_415,N_23416,N_24625);
and UO_416 (O_416,N_23814,N_23324);
or UO_417 (O_417,N_24929,N_23542);
or UO_418 (O_418,N_22513,N_22692);
nand UO_419 (O_419,N_24367,N_23327);
nand UO_420 (O_420,N_24913,N_24385);
nand UO_421 (O_421,N_23903,N_24638);
or UO_422 (O_422,N_22928,N_24321);
nor UO_423 (O_423,N_23981,N_23304);
xnor UO_424 (O_424,N_23087,N_22754);
xnor UO_425 (O_425,N_23998,N_24181);
xnor UO_426 (O_426,N_24931,N_22773);
xor UO_427 (O_427,N_23018,N_23096);
nor UO_428 (O_428,N_23308,N_22640);
nor UO_429 (O_429,N_24543,N_23855);
and UO_430 (O_430,N_23154,N_24206);
nand UO_431 (O_431,N_22704,N_23307);
or UO_432 (O_432,N_24652,N_24114);
or UO_433 (O_433,N_22638,N_24199);
nand UO_434 (O_434,N_24067,N_24616);
and UO_435 (O_435,N_22804,N_24976);
or UO_436 (O_436,N_23180,N_23084);
and UO_437 (O_437,N_24778,N_24982);
and UO_438 (O_438,N_23669,N_23426);
nor UO_439 (O_439,N_24703,N_24781);
or UO_440 (O_440,N_23664,N_22542);
or UO_441 (O_441,N_22956,N_24213);
or UO_442 (O_442,N_22589,N_24799);
or UO_443 (O_443,N_23608,N_22951);
xnor UO_444 (O_444,N_23963,N_23293);
nor UO_445 (O_445,N_23667,N_23567);
nand UO_446 (O_446,N_24662,N_22968);
xnor UO_447 (O_447,N_23048,N_23964);
and UO_448 (O_448,N_24723,N_24175);
and UO_449 (O_449,N_22807,N_24750);
nor UO_450 (O_450,N_22565,N_23427);
nand UO_451 (O_451,N_22737,N_22942);
nand UO_452 (O_452,N_23206,N_24079);
nand UO_453 (O_453,N_24698,N_23280);
and UO_454 (O_454,N_23763,N_23712);
xnor UO_455 (O_455,N_23424,N_24944);
xnor UO_456 (O_456,N_23438,N_23506);
or UO_457 (O_457,N_23285,N_24679);
nor UO_458 (O_458,N_22806,N_23436);
and UO_459 (O_459,N_23819,N_24187);
xor UO_460 (O_460,N_24859,N_24558);
xnor UO_461 (O_461,N_23475,N_24647);
xnor UO_462 (O_462,N_22858,N_22802);
nor UO_463 (O_463,N_22869,N_22832);
and UO_464 (O_464,N_22567,N_23423);
nor UO_465 (O_465,N_22778,N_24707);
nand UO_466 (O_466,N_22529,N_24283);
nor UO_467 (O_467,N_24214,N_22525);
or UO_468 (O_468,N_24963,N_23772);
nand UO_469 (O_469,N_23607,N_23639);
or UO_470 (O_470,N_24496,N_24580);
nand UO_471 (O_471,N_23123,N_23508);
and UO_472 (O_472,N_22835,N_23912);
or UO_473 (O_473,N_24754,N_22626);
or UO_474 (O_474,N_22585,N_23253);
xor UO_475 (O_475,N_24505,N_23575);
and UO_476 (O_476,N_22793,N_23502);
nor UO_477 (O_477,N_23286,N_23611);
nor UO_478 (O_478,N_23810,N_23471);
xor UO_479 (O_479,N_23545,N_22852);
and UO_480 (O_480,N_23388,N_24803);
and UO_481 (O_481,N_22763,N_24852);
and UO_482 (O_482,N_24300,N_24326);
nor UO_483 (O_483,N_24953,N_23564);
nor UO_484 (O_484,N_23058,N_23535);
or UO_485 (O_485,N_23648,N_24874);
or UO_486 (O_486,N_24244,N_24980);
nand UO_487 (O_487,N_23298,N_24861);
and UO_488 (O_488,N_22612,N_24677);
xor UO_489 (O_489,N_22970,N_23697);
or UO_490 (O_490,N_24061,N_23045);
xnor UO_491 (O_491,N_22520,N_23993);
nor UO_492 (O_492,N_22659,N_24833);
nor UO_493 (O_493,N_23017,N_22514);
nor UO_494 (O_494,N_24882,N_23031);
and UO_495 (O_495,N_22810,N_22974);
or UO_496 (O_496,N_23977,N_24276);
xor UO_497 (O_497,N_23880,N_24975);
xnor UO_498 (O_498,N_23052,N_24395);
xnor UO_499 (O_499,N_23151,N_24776);
nor UO_500 (O_500,N_23559,N_24523);
and UO_501 (O_501,N_24928,N_23823);
or UO_502 (O_502,N_24466,N_24172);
nand UO_503 (O_503,N_24127,N_22840);
nand UO_504 (O_504,N_22999,N_24965);
nand UO_505 (O_505,N_23706,N_22505);
nor UO_506 (O_506,N_24643,N_22986);
xnor UO_507 (O_507,N_23718,N_23640);
xnor UO_508 (O_508,N_24314,N_22786);
or UO_509 (O_509,N_22976,N_24337);
nor UO_510 (O_510,N_24765,N_24865);
nand UO_511 (O_511,N_24728,N_23645);
and UO_512 (O_512,N_23971,N_23596);
or UO_513 (O_513,N_22865,N_24846);
xnor UO_514 (O_514,N_23852,N_22909);
or UO_515 (O_515,N_24013,N_24827);
xor UO_516 (O_516,N_23318,N_23598);
xnor UO_517 (O_517,N_23878,N_23362);
and UO_518 (O_518,N_24531,N_23166);
nor UO_519 (O_519,N_23209,N_24571);
nand UO_520 (O_520,N_22590,N_23737);
nand UO_521 (O_521,N_24553,N_22694);
xor UO_522 (O_522,N_24053,N_23798);
xor UO_523 (O_523,N_22880,N_23563);
or UO_524 (O_524,N_24896,N_24602);
nor UO_525 (O_525,N_24517,N_23419);
and UO_526 (O_526,N_23408,N_23780);
or UO_527 (O_527,N_23428,N_23741);
xnor UO_528 (O_528,N_23224,N_23000);
nand UO_529 (O_529,N_23859,N_23922);
or UO_530 (O_530,N_24388,N_23281);
and UO_531 (O_531,N_24489,N_22751);
or UO_532 (O_532,N_24857,N_24358);
and UO_533 (O_533,N_22661,N_23478);
nor UO_534 (O_534,N_24561,N_22904);
nand UO_535 (O_535,N_23258,N_24049);
nand UO_536 (O_536,N_24340,N_24375);
nand UO_537 (O_537,N_23019,N_24131);
nand UO_538 (O_538,N_24105,N_24753);
nand UO_539 (O_539,N_23882,N_24041);
xor UO_540 (O_540,N_23952,N_23549);
xor UO_541 (O_541,N_24441,N_22531);
nor UO_542 (O_542,N_24983,N_23521);
xor UO_543 (O_543,N_22973,N_24878);
and UO_544 (O_544,N_24644,N_22749);
xnor UO_545 (O_545,N_22634,N_24521);
nand UO_546 (O_546,N_24551,N_23498);
or UO_547 (O_547,N_23338,N_23135);
and UO_548 (O_548,N_23995,N_24867);
nor UO_549 (O_549,N_24093,N_23333);
nand UO_550 (O_550,N_22595,N_24590);
nand UO_551 (O_551,N_22723,N_23215);
nand UO_552 (O_552,N_23941,N_22815);
nor UO_553 (O_553,N_23584,N_24584);
or UO_554 (O_554,N_24719,N_24552);
and UO_555 (O_555,N_24008,N_23493);
and UO_556 (O_556,N_24556,N_22878);
or UO_557 (O_557,N_23960,N_24045);
or UO_558 (O_558,N_24501,N_23875);
nand UO_559 (O_559,N_22545,N_23350);
xnor UO_560 (O_560,N_24593,N_24670);
or UO_561 (O_561,N_24768,N_24544);
nor UO_562 (O_562,N_24150,N_23158);
or UO_563 (O_563,N_24748,N_22782);
or UO_564 (O_564,N_24665,N_23925);
xnor UO_565 (O_565,N_24762,N_23311);
nand UO_566 (O_566,N_23870,N_24727);
or UO_567 (O_567,N_23447,N_22937);
nand UO_568 (O_568,N_23721,N_24490);
and UO_569 (O_569,N_23820,N_24092);
or UO_570 (O_570,N_24116,N_22673);
nor UO_571 (O_571,N_23068,N_23193);
nand UO_572 (O_572,N_23704,N_23226);
xor UO_573 (O_573,N_23817,N_24954);
nor UO_574 (O_574,N_24656,N_23275);
nor UO_575 (O_575,N_23885,N_22719);
xor UO_576 (O_576,N_23853,N_23495);
nor UO_577 (O_577,N_23192,N_23024);
and UO_578 (O_578,N_24790,N_23401);
nand UO_579 (O_579,N_24731,N_23690);
and UO_580 (O_580,N_22726,N_22629);
and UO_581 (O_581,N_22953,N_22760);
and UO_582 (O_582,N_24678,N_24812);
or UO_583 (O_583,N_23244,N_23171);
xor UO_584 (O_584,N_23679,N_23745);
or UO_585 (O_585,N_23700,N_24378);
and UO_586 (O_586,N_22730,N_23546);
xor UO_587 (O_587,N_22597,N_22712);
and UO_588 (O_588,N_24785,N_23916);
or UO_589 (O_589,N_23989,N_23261);
or UO_590 (O_590,N_24658,N_23796);
and UO_591 (O_591,N_24682,N_22665);
xor UO_592 (O_592,N_23578,N_24423);
xor UO_593 (O_593,N_24428,N_23747);
or UO_594 (O_594,N_23986,N_22500);
and UO_595 (O_595,N_24673,N_22553);
and UO_596 (O_596,N_24512,N_23587);
nor UO_597 (O_597,N_22870,N_22745);
and UO_598 (O_598,N_24926,N_24173);
nand UO_599 (O_599,N_24100,N_23523);
and UO_600 (O_600,N_23866,N_22511);
xor UO_601 (O_601,N_24346,N_23663);
and UO_602 (O_602,N_23174,N_24933);
xnor UO_603 (O_603,N_23804,N_24444);
xor UO_604 (O_604,N_24745,N_22647);
and UO_605 (O_605,N_22948,N_24596);
or UO_606 (O_606,N_24686,N_24922);
and UO_607 (O_607,N_24165,N_22670);
or UO_608 (O_608,N_24938,N_23251);
and UO_609 (O_609,N_24897,N_22509);
nand UO_610 (O_610,N_24033,N_24069);
xnor UO_611 (O_611,N_24210,N_24851);
xor UO_612 (O_612,N_23864,N_24802);
xnor UO_613 (O_613,N_23090,N_24987);
xnor UO_614 (O_614,N_24722,N_23326);
xnor UO_615 (O_615,N_23094,N_23354);
nand UO_616 (O_616,N_22664,N_23985);
xnor UO_617 (O_617,N_24610,N_23202);
nor UO_618 (O_618,N_24171,N_23278);
or UO_619 (O_619,N_23876,N_24529);
or UO_620 (O_620,N_22591,N_23425);
xor UO_621 (O_621,N_23322,N_24343);
nor UO_622 (O_622,N_22607,N_24497);
nand UO_623 (O_623,N_24764,N_24089);
and UO_624 (O_624,N_23256,N_22978);
nor UO_625 (O_625,N_23364,N_23955);
and UO_626 (O_626,N_24011,N_24520);
nor UO_627 (O_627,N_24484,N_23972);
nand UO_628 (O_628,N_24296,N_23453);
xor UO_629 (O_629,N_23701,N_23035);
xnor UO_630 (O_630,N_22539,N_23051);
and UO_631 (O_631,N_23509,N_23064);
and UO_632 (O_632,N_24541,N_23454);
nand UO_633 (O_633,N_23141,N_24509);
nor UO_634 (O_634,N_23431,N_24060);
xor UO_635 (O_635,N_22799,N_24866);
nand UO_636 (O_636,N_24479,N_24478);
nand UO_637 (O_637,N_23355,N_22981);
or UO_638 (O_638,N_22625,N_23393);
xnor UO_639 (O_639,N_23761,N_23091);
nor UO_640 (O_640,N_23479,N_23092);
nand UO_641 (O_641,N_23108,N_23469);
and UO_642 (O_642,N_24483,N_22521);
and UO_643 (O_643,N_24532,N_24193);
or UO_644 (O_644,N_23055,N_23757);
nor UO_645 (O_645,N_24917,N_23057);
and UO_646 (O_646,N_24320,N_22571);
and UO_647 (O_647,N_24313,N_22530);
xnor UO_648 (O_648,N_24383,N_22610);
nand UO_649 (O_649,N_22527,N_24436);
xnor UO_650 (O_650,N_22771,N_23016);
nand UO_651 (O_651,N_24927,N_24730);
nor UO_652 (O_652,N_24025,N_22733);
nand UO_653 (O_653,N_24099,N_24291);
nand UO_654 (O_654,N_23760,N_23348);
nand UO_655 (O_655,N_24236,N_23053);
nor UO_656 (O_656,N_24024,N_23869);
nor UO_657 (O_657,N_24125,N_22955);
and UO_658 (O_658,N_23636,N_23184);
nor UO_659 (O_659,N_24806,N_24277);
and UO_660 (O_660,N_23194,N_22541);
and UO_661 (O_661,N_22896,N_23452);
and UO_662 (O_662,N_22892,N_24248);
or UO_663 (O_663,N_24327,N_22924);
and UO_664 (O_664,N_23562,N_24380);
nand UO_665 (O_665,N_24424,N_22533);
nand UO_666 (O_666,N_24690,N_23371);
or UO_667 (O_667,N_24072,N_24631);
nor UO_668 (O_668,N_23139,N_24115);
and UO_669 (O_669,N_22881,N_22882);
and UO_670 (O_670,N_24091,N_23818);
nor UO_671 (O_671,N_24039,N_23605);
or UO_672 (O_672,N_24118,N_23848);
nand UO_673 (O_673,N_23620,N_23983);
nand UO_674 (O_674,N_23136,N_22628);
xnor UO_675 (O_675,N_23211,N_23264);
or UO_676 (O_676,N_24981,N_22814);
nand UO_677 (O_677,N_23776,N_22894);
and UO_678 (O_678,N_24968,N_23439);
nor UO_679 (O_679,N_24281,N_24786);
xnor UO_680 (O_680,N_23629,N_23260);
nand UO_681 (O_681,N_22534,N_22752);
nor UO_682 (O_682,N_22528,N_24822);
and UO_683 (O_683,N_24042,N_24240);
nand UO_684 (O_684,N_23365,N_23548);
nand UO_685 (O_685,N_23079,N_24189);
and UO_686 (O_686,N_24779,N_24615);
and UO_687 (O_687,N_22957,N_24601);
and UO_688 (O_688,N_23552,N_24693);
xnor UO_689 (O_689,N_22841,N_22698);
nor UO_690 (O_690,N_22679,N_24464);
nor UO_691 (O_691,N_24482,N_23480);
xor UO_692 (O_692,N_24062,N_24144);
nor UO_693 (O_693,N_22938,N_24714);
nand UO_694 (O_694,N_24009,N_24440);
nor UO_695 (O_695,N_23117,N_23967);
nor UO_696 (O_696,N_24554,N_24826);
xnor UO_697 (O_697,N_23191,N_23494);
or UO_698 (O_698,N_23243,N_24589);
and UO_699 (O_699,N_23588,N_23352);
nand UO_700 (O_700,N_23435,N_23394);
or UO_701 (O_701,N_23946,N_23901);
and UO_702 (O_702,N_23771,N_23694);
xor UO_703 (O_703,N_23754,N_23769);
nand UO_704 (O_704,N_22532,N_24048);
xor UO_705 (O_705,N_23530,N_24756);
xor UO_706 (O_706,N_24234,N_22800);
and UO_707 (O_707,N_23735,N_23473);
xor UO_708 (O_708,N_24015,N_22579);
nand UO_709 (O_709,N_22932,N_23707);
and UO_710 (O_710,N_24485,N_22738);
xnor UO_711 (O_711,N_24338,N_24226);
or UO_712 (O_712,N_24237,N_22656);
nand UO_713 (O_713,N_24032,N_24162);
nand UO_714 (O_714,N_24623,N_24612);
nand UO_715 (O_715,N_24075,N_23947);
xor UO_716 (O_716,N_24887,N_24043);
or UO_717 (O_717,N_24518,N_24958);
nor UO_718 (O_718,N_24964,N_22642);
and UO_719 (O_719,N_23579,N_23954);
and UO_720 (O_720,N_23160,N_24153);
nand UO_721 (O_721,N_23379,N_24869);
nand UO_722 (O_722,N_23164,N_24513);
or UO_723 (O_723,N_24978,N_22547);
xnor UO_724 (O_724,N_23196,N_22744);
xor UO_725 (O_725,N_23844,N_22504);
xor UO_726 (O_726,N_24977,N_23628);
and UO_727 (O_727,N_24284,N_23279);
xor UO_728 (O_728,N_23551,N_23273);
nand UO_729 (O_729,N_23516,N_23086);
or UO_730 (O_730,N_24537,N_24353);
nor UO_731 (O_731,N_22868,N_23942);
or UO_732 (O_732,N_23050,N_23911);
and UO_733 (O_733,N_23126,N_23147);
xnor UO_734 (O_734,N_24701,N_24230);
and UO_735 (O_735,N_24576,N_24831);
nor UO_736 (O_736,N_23843,N_22873);
xor UO_737 (O_737,N_24241,N_24572);
or UO_738 (O_738,N_23717,N_23858);
nand UO_739 (O_739,N_22580,N_22818);
xor UO_740 (O_740,N_23065,N_23649);
and UO_741 (O_741,N_24691,N_24894);
or UO_742 (O_742,N_23432,N_24176);
nand UO_743 (O_743,N_24268,N_23356);
or UO_744 (O_744,N_24342,N_23269);
xor UO_745 (O_745,N_23618,N_23910);
or UO_746 (O_746,N_24417,N_23061);
nor UO_747 (O_747,N_22844,N_22699);
and UO_748 (O_748,N_24798,N_23913);
nand UO_749 (O_749,N_22711,N_22522);
nand UO_750 (O_750,N_24829,N_24788);
nor UO_751 (O_751,N_22615,N_24881);
xor UO_752 (O_752,N_24411,N_23825);
nor UO_753 (O_753,N_22939,N_24741);
xor UO_754 (O_754,N_22596,N_23527);
or UO_755 (O_755,N_23214,N_24811);
and UO_756 (O_756,N_23655,N_23909);
nand UO_757 (O_757,N_23774,N_23014);
nor UO_758 (O_758,N_24864,N_24710);
nor UO_759 (O_759,N_23319,N_23344);
and UO_760 (O_760,N_24225,N_23501);
nand UO_761 (O_761,N_24445,N_22961);
nand UO_762 (O_762,N_22710,N_22929);
and UO_763 (O_763,N_24454,N_23590);
nor UO_764 (O_764,N_24668,N_24696);
xor UO_765 (O_765,N_24063,N_24255);
nor UO_766 (O_766,N_24371,N_23801);
nand UO_767 (O_767,N_24809,N_23115);
and UO_768 (O_768,N_24016,N_24409);
nor UO_769 (O_769,N_24583,N_24540);
xor UO_770 (O_770,N_24524,N_24709);
or UO_771 (O_771,N_24959,N_23688);
nand UO_772 (O_772,N_22803,N_24399);
and UO_773 (O_773,N_24704,N_23404);
nand UO_774 (O_774,N_23300,N_24026);
or UO_775 (O_775,N_22652,N_24018);
xor UO_776 (O_776,N_24862,N_23037);
and UO_777 (O_777,N_24369,N_22925);
and UO_778 (O_778,N_23626,N_24559);
nor UO_779 (O_779,N_23902,N_22838);
or UO_780 (O_780,N_23623,N_23380);
or UO_781 (O_781,N_24546,N_24807);
nor UO_782 (O_782,N_24336,N_23634);
xnor UO_783 (O_783,N_24134,N_24022);
or UO_784 (O_784,N_23137,N_24767);
nor UO_785 (O_785,N_23245,N_24795);
nor UO_786 (O_786,N_23005,N_23660);
or UO_787 (O_787,N_24017,N_23296);
nor UO_788 (O_788,N_23063,N_22992);
or UO_789 (O_789,N_23515,N_23609);
nand UO_790 (O_790,N_23148,N_23472);
nor UO_791 (O_791,N_23402,N_24218);
or UO_792 (O_792,N_23571,N_24675);
nor UO_793 (O_793,N_23740,N_24934);
or UO_794 (O_794,N_23089,N_22603);
nor UO_795 (O_795,N_24940,N_24801);
nor UO_796 (O_796,N_24514,N_22550);
or UO_797 (O_797,N_24047,N_24468);
xor UO_798 (O_798,N_24128,N_24169);
nand UO_799 (O_799,N_23973,N_23968);
nor UO_800 (O_800,N_23923,N_24023);
nand UO_801 (O_801,N_24438,N_24442);
nor UO_802 (O_802,N_24259,N_24219);
nand UO_803 (O_803,N_24603,N_22668);
xnor UO_804 (O_804,N_22920,N_24156);
nand UO_805 (O_805,N_24974,N_24805);
nand UO_806 (O_806,N_22900,N_23132);
and UO_807 (O_807,N_23178,N_23462);
or UO_808 (O_808,N_23182,N_23782);
xnor UO_809 (O_809,N_22775,N_24751);
or UO_810 (O_810,N_23455,N_24328);
and UO_811 (O_811,N_24159,N_24948);
xor UO_812 (O_812,N_24789,N_24769);
and UO_813 (O_813,N_24120,N_23770);
xor UO_814 (O_814,N_24059,N_23078);
nand UO_815 (O_815,N_23813,N_23390);
or UO_816 (O_816,N_24733,N_24921);
nand UO_817 (O_817,N_23507,N_24820);
nor UO_818 (O_818,N_22682,N_23698);
and UO_819 (O_819,N_24461,N_23006);
and UO_820 (O_820,N_24573,N_23788);
nor UO_821 (O_821,N_22506,N_24567);
xor UO_822 (O_822,N_23828,N_23750);
nor UO_823 (O_823,N_23034,N_23599);
xor UO_824 (O_824,N_23113,N_24515);
nand UO_825 (O_825,N_23847,N_23920);
nand UO_826 (O_826,N_23824,N_23854);
and UO_827 (O_827,N_24393,N_23272);
and UO_828 (O_828,N_23795,N_24473);
or UO_829 (O_829,N_23312,N_24796);
or UO_830 (O_830,N_24654,N_24027);
and UO_831 (O_831,N_23349,N_22859);
nor UO_832 (O_832,N_23309,N_23284);
nor UO_833 (O_833,N_23332,N_24570);
nor UO_834 (O_834,N_22662,N_22646);
nand UO_835 (O_835,N_23466,N_24973);
and UO_836 (O_836,N_23482,N_23361);
and UO_837 (O_837,N_24030,N_22930);
or UO_838 (O_838,N_23397,N_23943);
or UO_839 (O_839,N_22864,N_22982);
and UO_840 (O_840,N_24392,N_24191);
and UO_841 (O_841,N_23722,N_24209);
nand UO_842 (O_842,N_23070,N_22622);
and UO_843 (O_843,N_23794,N_24528);
or UO_844 (O_844,N_23363,N_23225);
nand UO_845 (O_845,N_24999,N_22633);
nand UO_846 (O_846,N_22990,N_23124);
nand UO_847 (O_847,N_23860,N_24899);
or UO_848 (O_848,N_23028,N_24800);
or UO_849 (O_849,N_23687,N_24702);
nand UO_850 (O_850,N_24663,N_24895);
nor UO_851 (O_851,N_22843,N_24817);
nor UO_852 (O_852,N_22785,N_23489);
nor UO_853 (O_853,N_22801,N_24694);
nand UO_854 (O_854,N_23742,N_23103);
nand UO_855 (O_855,N_22696,N_24939);
or UO_856 (O_856,N_24634,N_22876);
nor UO_857 (O_857,N_24742,N_24050);
and UO_858 (O_858,N_23676,N_23400);
xor UO_859 (O_859,N_24232,N_24474);
and UO_860 (O_860,N_22787,N_22575);
and UO_861 (O_861,N_23881,N_23674);
or UO_862 (O_862,N_22641,N_24000);
nand UO_863 (O_863,N_23345,N_22965);
nand UO_864 (O_864,N_23499,N_23127);
xor UO_865 (O_865,N_22758,N_24096);
or UO_866 (O_866,N_23651,N_23101);
nor UO_867 (O_867,N_22853,N_24787);
xor UO_868 (O_868,N_24130,N_24195);
or UO_869 (O_869,N_23800,N_24950);
nor UO_870 (O_870,N_23834,N_24614);
or UO_871 (O_871,N_23900,N_23969);
and UO_872 (O_872,N_23835,N_23204);
and UO_873 (O_873,N_24622,N_24470);
and UO_874 (O_874,N_24289,N_23276);
and UO_875 (O_875,N_22602,N_24364);
nor UO_876 (O_876,N_24919,N_22526);
or UO_877 (O_877,N_24046,N_22830);
or UO_878 (O_878,N_23753,N_24835);
nor UO_879 (O_879,N_24349,N_22572);
and UO_880 (O_880,N_23622,N_22649);
nand UO_881 (O_881,N_24655,N_24170);
or UO_882 (O_882,N_24307,N_23965);
and UO_883 (O_883,N_23790,N_23560);
or UO_884 (O_884,N_24208,N_23653);
nand UO_885 (O_885,N_23347,N_24886);
nand UO_886 (O_886,N_23039,N_23242);
and UO_887 (O_887,N_22829,N_23748);
nor UO_888 (O_888,N_23731,N_24224);
or UO_889 (O_889,N_23736,N_24303);
nor UO_890 (O_890,N_24618,N_23684);
or UO_891 (O_891,N_24078,N_24739);
xor UO_892 (O_892,N_23444,N_23962);
and UO_893 (O_893,N_23069,N_23410);
xor UO_894 (O_894,N_24952,N_24095);
nand UO_895 (O_895,N_23615,N_23029);
nand UO_896 (O_896,N_22753,N_23933);
or UO_897 (O_897,N_24401,N_24330);
and UO_898 (O_898,N_23889,N_23577);
or UO_899 (O_899,N_22573,N_23082);
xnor UO_900 (O_900,N_24955,N_23767);
or UO_901 (O_901,N_24398,N_22919);
nor UO_902 (O_902,N_23948,N_23336);
nand UO_903 (O_903,N_24231,N_24685);
nor UO_904 (O_904,N_23789,N_24889);
or UO_905 (O_905,N_22568,N_24278);
nand UO_906 (O_906,N_23485,N_23764);
and UO_907 (O_907,N_23805,N_24333);
nor UO_908 (O_908,N_24290,N_23059);
or UO_909 (O_909,N_23867,N_24971);
and UO_910 (O_910,N_24860,N_24040);
nor UO_911 (O_911,N_23445,N_24606);
nand UO_912 (O_912,N_24373,N_23476);
nand UO_913 (O_913,N_23891,N_23650);
and UO_914 (O_914,N_24348,N_23199);
and UO_915 (O_915,N_23367,N_24661);
and UO_916 (O_916,N_22552,N_24391);
nand UO_917 (O_917,N_23996,N_24967);
and UO_918 (O_918,N_23691,N_24451);
nand UO_919 (O_919,N_24310,N_24669);
or UO_920 (O_920,N_22943,N_23213);
and UO_921 (O_921,N_24498,N_24689);
or UO_922 (O_922,N_24090,N_23188);
xnor UO_923 (O_923,N_24122,N_23528);
and UO_924 (O_924,N_22944,N_24773);
and UO_925 (O_925,N_24136,N_24293);
nor UO_926 (O_926,N_23143,N_23792);
nand UO_927 (O_927,N_23175,N_22996);
xnor UO_928 (O_928,N_24212,N_23392);
nor UO_929 (O_929,N_22780,N_22515);
nand UO_930 (O_930,N_23517,N_22931);
xor UO_931 (O_931,N_23441,N_23197);
xnor UO_932 (O_932,N_23381,N_24821);
xor UO_933 (O_933,N_24065,N_23670);
nand UO_934 (O_934,N_24312,N_23832);
xor UO_935 (O_935,N_24306,N_24579);
or UO_936 (O_936,N_24738,N_23850);
nor UO_937 (O_937,N_24988,N_24557);
nor UO_938 (O_938,N_24705,N_23093);
or UO_939 (O_939,N_23583,N_24536);
and UO_940 (O_940,N_23187,N_24305);
and UO_941 (O_941,N_22687,N_23856);
or UO_942 (O_942,N_22820,N_22945);
xor UO_943 (O_943,N_23526,N_24292);
or UO_944 (O_944,N_24163,N_22791);
nand UO_945 (O_945,N_24533,N_24605);
nand UO_946 (O_946,N_24052,N_24966);
nand UO_947 (O_947,N_24157,N_24077);
nand UO_948 (O_948,N_24947,N_24158);
and UO_949 (O_949,N_22593,N_24969);
and UO_950 (O_950,N_23775,N_24174);
or UO_951 (O_951,N_23815,N_24511);
xor UO_952 (O_952,N_24309,N_24203);
nand UO_953 (O_953,N_23465,N_24771);
or UO_954 (O_954,N_23474,N_23641);
or UO_955 (O_955,N_23657,N_23896);
nor UO_956 (O_956,N_22959,N_23816);
nand UO_957 (O_957,N_22693,N_24951);
or UO_958 (O_958,N_23463,N_23808);
xnor UO_959 (O_959,N_22985,N_23366);
nor UO_960 (O_960,N_24945,N_23046);
and UO_961 (O_961,N_24229,N_23054);
xor UO_962 (O_962,N_23384,N_22935);
or UO_963 (O_963,N_23591,N_23282);
or UO_964 (O_964,N_23898,N_24202);
nand UO_965 (O_965,N_22663,N_22721);
and UO_966 (O_966,N_24684,N_23893);
nand UO_967 (O_967,N_22774,N_23222);
and UO_968 (O_968,N_24491,N_22731);
nor UO_969 (O_969,N_24585,N_24317);
and UO_970 (O_970,N_23603,N_23619);
xnor UO_971 (O_971,N_22540,N_24717);
and UO_972 (O_972,N_24102,N_22891);
and UO_973 (O_973,N_24566,N_22759);
and UO_974 (O_974,N_24626,N_23543);
nor UO_975 (O_975,N_23488,N_24998);
xor UO_976 (O_976,N_23004,N_23956);
and UO_977 (O_977,N_24653,N_24760);
and UO_978 (O_978,N_24633,N_24106);
and UO_979 (O_979,N_24288,N_23637);
and UO_980 (O_980,N_22734,N_23566);
and UO_981 (O_981,N_24301,N_24737);
xnor UO_982 (O_982,N_24140,N_23849);
nand UO_983 (O_983,N_24957,N_23601);
or UO_984 (O_984,N_23938,N_24588);
or UO_985 (O_985,N_23572,N_24021);
xnor UO_986 (O_986,N_23803,N_22821);
nor UO_987 (O_987,N_24577,N_23678);
or UO_988 (O_988,N_23022,N_24167);
nor UO_989 (O_989,N_23330,N_23026);
or UO_990 (O_990,N_23865,N_23218);
nand UO_991 (O_991,N_23360,N_24695);
or UO_992 (O_992,N_23846,N_24269);
or UO_993 (O_993,N_23207,N_24858);
or UO_994 (O_994,N_23758,N_23303);
nor UO_995 (O_995,N_24777,N_24119);
nand UO_996 (O_996,N_23799,N_24744);
or UO_997 (O_997,N_24793,N_23680);
nor UO_998 (O_998,N_23049,N_24718);
or UO_999 (O_999,N_24639,N_23252);
nor UO_1000 (O_1000,N_24901,N_24161);
nand UO_1001 (O_1001,N_24883,N_24271);
nand UO_1002 (O_1002,N_22576,N_24396);
or UO_1003 (O_1003,N_23072,N_24712);
or UO_1004 (O_1004,N_22941,N_24243);
nor UO_1005 (O_1005,N_24448,N_24347);
and UO_1006 (O_1006,N_23170,N_24455);
or UO_1007 (O_1007,N_24168,N_22609);
nand UO_1008 (O_1008,N_23491,N_24856);
nor UO_1009 (O_1009,N_24503,N_23378);
nand UO_1010 (O_1010,N_23531,N_24354);
and UO_1011 (O_1011,N_23173,N_24311);
xnor UO_1012 (O_1012,N_23683,N_23897);
nor UO_1013 (O_1013,N_24692,N_24700);
nor UO_1014 (O_1014,N_23582,N_23189);
or UO_1015 (O_1015,N_24247,N_24646);
xor UO_1016 (O_1016,N_24837,N_23477);
and UO_1017 (O_1017,N_24613,N_23003);
and UO_1018 (O_1018,N_23630,N_22772);
and UO_1019 (O_1019,N_24984,N_22566);
nor UO_1020 (O_1020,N_24434,N_22686);
xnor UO_1021 (O_1021,N_22768,N_23553);
nand UO_1022 (O_1022,N_23568,N_23503);
nand UO_1023 (O_1023,N_24504,N_24519);
and UO_1024 (O_1024,N_22916,N_24808);
and UO_1025 (O_1025,N_24794,N_22798);
nor UO_1026 (O_1026,N_22879,N_24149);
xnor UO_1027 (O_1027,N_24495,N_23464);
and UO_1028 (O_1028,N_22748,N_23161);
xnor UO_1029 (O_1029,N_24420,N_24920);
and UO_1030 (O_1030,N_24905,N_23177);
or UO_1031 (O_1031,N_24003,N_23573);
or UO_1032 (O_1032,N_24804,N_24904);
nor UO_1033 (O_1033,N_24797,N_23624);
or UO_1034 (O_1034,N_24547,N_23009);
xnor UO_1035 (O_1035,N_24433,N_24286);
or UO_1036 (O_1036,N_23257,N_22796);
xnor UO_1037 (O_1037,N_23915,N_23297);
nand UO_1038 (O_1038,N_23631,N_24535);
or UO_1039 (O_1039,N_24985,N_24406);
or UO_1040 (O_1040,N_22940,N_23632);
and UO_1041 (O_1041,N_24956,N_22781);
xnor UO_1042 (O_1042,N_22908,N_23686);
nor UO_1043 (O_1043,N_23373,N_23625);
or UO_1044 (O_1044,N_22906,N_22614);
nor UO_1045 (O_1045,N_23538,N_23263);
or UO_1046 (O_1046,N_23449,N_23313);
xnor UO_1047 (O_1047,N_22667,N_24989);
or UO_1048 (O_1048,N_24766,N_23539);
nand UO_1049 (O_1049,N_24545,N_24245);
nor UO_1050 (O_1050,N_24425,N_24871);
nor UO_1051 (O_1051,N_23153,N_24400);
nor UO_1052 (O_1052,N_24850,N_23483);
nor UO_1053 (O_1053,N_23314,N_24270);
and UO_1054 (O_1054,N_24299,N_22727);
or UO_1055 (O_1055,N_23957,N_22867);
and UO_1056 (O_1056,N_23395,N_22637);
xor UO_1057 (O_1057,N_23335,N_22998);
xor UO_1058 (O_1058,N_23459,N_23012);
or UO_1059 (O_1059,N_23934,N_24568);
xor UO_1060 (O_1060,N_24752,N_23234);
nand UO_1061 (O_1061,N_23486,N_24020);
or UO_1062 (O_1062,N_23216,N_24109);
or UO_1063 (O_1063,N_24035,N_23413);
or UO_1064 (O_1064,N_23703,N_24319);
xor UO_1065 (O_1065,N_24256,N_23755);
and UO_1066 (O_1066,N_22551,N_22947);
and UO_1067 (O_1067,N_22761,N_22561);
nor UO_1068 (O_1068,N_22671,N_23500);
or UO_1069 (O_1069,N_23999,N_24216);
and UO_1070 (O_1070,N_24402,N_23845);
xnor UO_1071 (O_1071,N_22695,N_22889);
nor UO_1072 (O_1072,N_22535,N_23600);
nand UO_1073 (O_1073,N_22627,N_24494);
nor UO_1074 (O_1074,N_23532,N_24743);
or UO_1075 (O_1075,N_22958,N_24937);
or UO_1076 (O_1076,N_23504,N_23110);
or UO_1077 (O_1077,N_24239,N_24104);
nor UO_1078 (O_1078,N_22849,N_23695);
nand UO_1079 (O_1079,N_22984,N_23581);
nor UO_1080 (O_1080,N_24582,N_22822);
nor UO_1081 (O_1081,N_23522,N_23156);
nand UO_1082 (O_1082,N_24467,N_23716);
nor UO_1083 (O_1083,N_23240,N_22675);
or UO_1084 (O_1084,N_24994,N_24854);
and UO_1085 (O_1085,N_23979,N_23176);
nand UO_1086 (O_1086,N_24659,N_23550);
or UO_1087 (O_1087,N_23783,N_24368);
nor UO_1088 (O_1088,N_24961,N_24379);
and UO_1089 (O_1089,N_24527,N_24421);
or UO_1090 (O_1090,N_23949,N_22936);
or UO_1091 (O_1091,N_24146,N_24339);
nor UO_1092 (O_1092,N_23970,N_23430);
or UO_1093 (O_1093,N_24233,N_22839);
or UO_1094 (O_1094,N_23738,N_24316);
and UO_1095 (O_1095,N_23015,N_24262);
and UO_1096 (O_1096,N_23370,N_24098);
or UO_1097 (O_1097,N_22783,N_23433);
or UO_1098 (O_1098,N_22660,N_24716);
and UO_1099 (O_1099,N_23939,N_23524);
nor UO_1100 (O_1100,N_23118,N_23621);
xor UO_1101 (O_1101,N_23076,N_24412);
xor UO_1102 (O_1102,N_22658,N_23851);
nand UO_1103 (O_1103,N_22544,N_23165);
or UO_1104 (O_1104,N_22584,N_23097);
xnor UO_1105 (O_1105,N_24435,N_23295);
xnor UO_1106 (O_1106,N_23233,N_24410);
and UO_1107 (O_1107,N_24192,N_22617);
nand UO_1108 (O_1108,N_23830,N_24295);
nor UO_1109 (O_1109,N_24054,N_24151);
nor UO_1110 (O_1110,N_24182,N_24254);
and UO_1111 (O_1111,N_24840,N_22893);
nand UO_1112 (O_1112,N_23635,N_24810);
and UO_1113 (O_1113,N_24331,N_22677);
nand UO_1114 (O_1114,N_24575,N_22680);
nor UO_1115 (O_1115,N_22746,N_22927);
xnor UO_1116 (O_1116,N_24266,N_23219);
or UO_1117 (O_1117,N_24126,N_23266);
xor UO_1118 (O_1118,N_22975,N_22666);
xnor UO_1119 (O_1119,N_24178,N_24137);
and UO_1120 (O_1120,N_23892,N_23429);
xnor UO_1121 (O_1121,N_24362,N_24747);
or UO_1122 (O_1122,N_23292,N_24892);
nand UO_1123 (O_1123,N_22764,N_23008);
nor UO_1124 (O_1124,N_22997,N_23907);
xor UO_1125 (O_1125,N_23088,N_24516);
nor UO_1126 (O_1126,N_24674,N_23104);
xor UO_1127 (O_1127,N_23797,N_22884);
or UO_1128 (O_1128,N_22825,N_23821);
nor UO_1129 (O_1129,N_23422,N_23112);
nand UO_1130 (O_1130,N_22993,N_22905);
and UO_1131 (O_1131,N_22706,N_23398);
or UO_1132 (O_1132,N_24297,N_22700);
nand UO_1133 (O_1133,N_24201,N_22861);
nor UO_1134 (O_1134,N_22967,N_23033);
xnor UO_1135 (O_1135,N_23405,N_23073);
and UO_1136 (O_1136,N_22987,N_22972);
xnor UO_1137 (O_1137,N_23412,N_22608);
xor UO_1138 (O_1138,N_24909,N_23223);
and UO_1139 (O_1139,N_23316,N_24671);
and UO_1140 (O_1140,N_23656,N_23873);
xnor UO_1141 (O_1141,N_24713,N_22586);
xnor UO_1142 (O_1142,N_24408,N_24780);
and UO_1143 (O_1143,N_23781,N_22827);
and UO_1144 (O_1144,N_22969,N_24124);
nor UO_1145 (O_1145,N_24783,N_24094);
xnor UO_1146 (O_1146,N_23642,N_24356);
nand UO_1147 (O_1147,N_23744,N_23385);
xnor UO_1148 (O_1148,N_23525,N_24666);
nor UO_1149 (O_1149,N_23809,N_23773);
nor UO_1150 (O_1150,N_23974,N_23720);
nand UO_1151 (O_1151,N_22848,N_24592);
or UO_1152 (O_1152,N_23383,N_24007);
xnor UO_1153 (O_1153,N_23440,N_23377);
or UO_1154 (O_1154,N_24397,N_24530);
or UO_1155 (O_1155,N_22949,N_23743);
nand UO_1156 (O_1156,N_24029,N_24083);
nand UO_1157 (O_1157,N_24264,N_22811);
nand UO_1158 (O_1158,N_23468,N_24930);
or UO_1159 (O_1159,N_23561,N_24257);
nor UO_1160 (O_1160,N_23417,N_22562);
and UO_1161 (O_1161,N_22599,N_23011);
nor UO_1162 (O_1162,N_22862,N_24563);
xnor UO_1163 (O_1163,N_22991,N_24432);
and UO_1164 (O_1164,N_22735,N_24749);
xor UO_1165 (O_1165,N_23040,N_23842);
or UO_1166 (O_1166,N_24609,N_23042);
nor UO_1167 (O_1167,N_24207,N_22650);
or UO_1168 (O_1168,N_23547,N_24180);
nand UO_1169 (O_1169,N_24876,N_24228);
xnor UO_1170 (O_1170,N_23221,N_24058);
or UO_1171 (O_1171,N_23839,N_22537);
and UO_1172 (O_1172,N_24770,N_22563);
and UO_1173 (O_1173,N_23533,N_24179);
nor UO_1174 (O_1174,N_22856,N_23802);
xnor UO_1175 (O_1175,N_23481,N_23236);
and UO_1176 (O_1176,N_24604,N_24427);
and UO_1177 (O_1177,N_22797,N_24155);
nand UO_1178 (O_1178,N_24624,N_23868);
xor UO_1179 (O_1179,N_23727,N_23265);
nor UO_1180 (O_1180,N_23927,N_23277);
or UO_1181 (O_1181,N_24374,N_22714);
nor UO_1182 (O_1182,N_23837,N_24166);
nor UO_1183 (O_1183,N_23434,N_23529);
nand UO_1184 (O_1184,N_23884,N_23080);
nor UO_1185 (O_1185,N_23841,N_24164);
nand UO_1186 (O_1186,N_24836,N_23102);
and UO_1187 (O_1187,N_24282,N_23409);
nand UO_1188 (O_1188,N_22788,N_24308);
and UO_1189 (O_1189,N_24450,N_24885);
nand UO_1190 (O_1190,N_24942,N_23730);
nand UO_1191 (O_1191,N_23904,N_23739);
xor UO_1192 (O_1192,N_24863,N_24111);
or UO_1193 (O_1193,N_24595,N_24463);
nand UO_1194 (O_1194,N_22631,N_23337);
or UO_1195 (O_1195,N_23978,N_22703);
or UO_1196 (O_1196,N_24315,N_23368);
nor UO_1197 (O_1197,N_24139,N_24855);
and UO_1198 (O_1198,N_23310,N_24996);
or UO_1199 (O_1199,N_22863,N_23822);
and UO_1200 (O_1200,N_23448,N_22605);
nand UO_1201 (O_1201,N_24486,N_24564);
and UO_1202 (O_1202,N_24272,N_22777);
or UO_1203 (O_1203,N_23807,N_23570);
nor UO_1204 (O_1204,N_23220,N_23791);
and UO_1205 (O_1205,N_22750,N_23728);
and UO_1206 (O_1206,N_23186,N_22681);
xnor UO_1207 (O_1207,N_24325,N_24906);
and UO_1208 (O_1208,N_23926,N_24481);
nor UO_1209 (O_1209,N_23936,N_24456);
xnor UO_1210 (O_1210,N_24352,N_24154);
xnor UO_1211 (O_1211,N_24422,N_24458);
and UO_1212 (O_1212,N_23874,N_22549);
or UO_1213 (O_1213,N_23262,N_23659);
xnor UO_1214 (O_1214,N_22933,N_23144);
nand UO_1215 (O_1215,N_22621,N_23106);
xnor UO_1216 (O_1216,N_23558,N_24740);
xor UO_1217 (O_1217,N_22823,N_24774);
nor UO_1218 (O_1218,N_23918,N_22934);
and UO_1219 (O_1219,N_22577,N_23198);
and UO_1220 (O_1220,N_22795,N_24205);
nand UO_1221 (O_1221,N_22583,N_24877);
nand UO_1222 (O_1222,N_24818,N_24215);
nand UO_1223 (O_1223,N_24014,N_24133);
and UO_1224 (O_1224,N_24103,N_23614);
nor UO_1225 (O_1225,N_24772,N_23231);
and UO_1226 (O_1226,N_22548,N_23152);
or UO_1227 (O_1227,N_23519,N_23937);
or UO_1228 (O_1228,N_23569,N_23056);
and UO_1229 (O_1229,N_23317,N_24415);
and UO_1230 (O_1230,N_24814,N_24200);
or UO_1231 (O_1231,N_24627,N_22866);
nor UO_1232 (O_1232,N_24898,N_24949);
nor UO_1233 (O_1233,N_23032,N_22685);
or UO_1234 (O_1234,N_23906,N_22639);
or UO_1235 (O_1235,N_22557,N_23179);
and UO_1236 (O_1236,N_24715,N_23861);
or UO_1237 (O_1237,N_23914,N_22901);
or UO_1238 (O_1238,N_24912,N_22517);
nand UO_1239 (O_1239,N_23339,N_23044);
and UO_1240 (O_1240,N_23217,N_23162);
nand UO_1241 (O_1241,N_23287,N_23627);
xor UO_1242 (O_1242,N_23134,N_22911);
xor UO_1243 (O_1243,N_23062,N_23826);
nand UO_1244 (O_1244,N_24183,N_23613);
or UO_1245 (O_1245,N_23537,N_23201);
nand UO_1246 (O_1246,N_23534,N_22604);
and UO_1247 (O_1247,N_22847,N_23208);
or UO_1248 (O_1248,N_22508,N_23484);
or UO_1249 (O_1249,N_23249,N_24734);
or UO_1250 (O_1250,N_23496,N_24730);
nor UO_1251 (O_1251,N_24203,N_23400);
nor UO_1252 (O_1252,N_22941,N_23950);
xnor UO_1253 (O_1253,N_24759,N_23113);
xor UO_1254 (O_1254,N_24645,N_23011);
xor UO_1255 (O_1255,N_23259,N_23305);
and UO_1256 (O_1256,N_24986,N_24823);
or UO_1257 (O_1257,N_24661,N_22640);
and UO_1258 (O_1258,N_23397,N_24970);
nor UO_1259 (O_1259,N_24855,N_23999);
nor UO_1260 (O_1260,N_23761,N_24268);
nand UO_1261 (O_1261,N_23923,N_23916);
nand UO_1262 (O_1262,N_24427,N_24554);
nor UO_1263 (O_1263,N_24550,N_23050);
nand UO_1264 (O_1264,N_23081,N_23880);
xor UO_1265 (O_1265,N_24445,N_23843);
or UO_1266 (O_1266,N_24902,N_24797);
or UO_1267 (O_1267,N_23018,N_23505);
nand UO_1268 (O_1268,N_22862,N_24605);
xnor UO_1269 (O_1269,N_24636,N_23952);
or UO_1270 (O_1270,N_22738,N_24262);
nand UO_1271 (O_1271,N_24559,N_24011);
nor UO_1272 (O_1272,N_23199,N_23432);
xor UO_1273 (O_1273,N_24182,N_23522);
xor UO_1274 (O_1274,N_24820,N_22519);
nand UO_1275 (O_1275,N_23928,N_24416);
and UO_1276 (O_1276,N_23776,N_23393);
xor UO_1277 (O_1277,N_23057,N_24964);
xor UO_1278 (O_1278,N_24074,N_22939);
xor UO_1279 (O_1279,N_23602,N_23680);
and UO_1280 (O_1280,N_24179,N_22622);
or UO_1281 (O_1281,N_24272,N_23523);
xnor UO_1282 (O_1282,N_22982,N_24612);
nor UO_1283 (O_1283,N_22585,N_24149);
xnor UO_1284 (O_1284,N_24854,N_22732);
and UO_1285 (O_1285,N_23883,N_24030);
nor UO_1286 (O_1286,N_23642,N_23305);
and UO_1287 (O_1287,N_24937,N_24556);
nand UO_1288 (O_1288,N_23687,N_24535);
or UO_1289 (O_1289,N_24915,N_23996);
nor UO_1290 (O_1290,N_24609,N_24241);
xnor UO_1291 (O_1291,N_23615,N_22585);
nand UO_1292 (O_1292,N_24142,N_23850);
nor UO_1293 (O_1293,N_24545,N_24704);
nor UO_1294 (O_1294,N_22710,N_24905);
and UO_1295 (O_1295,N_23835,N_24732);
nor UO_1296 (O_1296,N_23316,N_22509);
and UO_1297 (O_1297,N_22908,N_24047);
and UO_1298 (O_1298,N_24738,N_22513);
nand UO_1299 (O_1299,N_23985,N_24531);
nand UO_1300 (O_1300,N_22762,N_22673);
or UO_1301 (O_1301,N_23006,N_23266);
and UO_1302 (O_1302,N_23495,N_24022);
xor UO_1303 (O_1303,N_22763,N_23284);
nand UO_1304 (O_1304,N_22856,N_24849);
and UO_1305 (O_1305,N_22582,N_23218);
nor UO_1306 (O_1306,N_24709,N_24855);
or UO_1307 (O_1307,N_22632,N_23837);
xor UO_1308 (O_1308,N_23371,N_24010);
nand UO_1309 (O_1309,N_23081,N_24210);
nand UO_1310 (O_1310,N_24119,N_24307);
nor UO_1311 (O_1311,N_23412,N_22527);
nor UO_1312 (O_1312,N_23438,N_23779);
xnor UO_1313 (O_1313,N_23428,N_23005);
nor UO_1314 (O_1314,N_22759,N_23642);
nand UO_1315 (O_1315,N_23091,N_23961);
or UO_1316 (O_1316,N_24894,N_23157);
nand UO_1317 (O_1317,N_23449,N_24078);
nand UO_1318 (O_1318,N_24121,N_22649);
nor UO_1319 (O_1319,N_24120,N_23227);
and UO_1320 (O_1320,N_22608,N_24573);
and UO_1321 (O_1321,N_23578,N_24021);
or UO_1322 (O_1322,N_24410,N_22820);
nor UO_1323 (O_1323,N_22685,N_22872);
xnor UO_1324 (O_1324,N_23216,N_23562);
nand UO_1325 (O_1325,N_22525,N_24164);
nor UO_1326 (O_1326,N_23489,N_23050);
xor UO_1327 (O_1327,N_22721,N_23885);
nand UO_1328 (O_1328,N_23313,N_24758);
nor UO_1329 (O_1329,N_23290,N_22760);
nand UO_1330 (O_1330,N_24776,N_24456);
nor UO_1331 (O_1331,N_23918,N_23561);
or UO_1332 (O_1332,N_23505,N_23756);
nor UO_1333 (O_1333,N_23350,N_23337);
nor UO_1334 (O_1334,N_23647,N_23122);
xor UO_1335 (O_1335,N_22745,N_23815);
xnor UO_1336 (O_1336,N_22573,N_23792);
nor UO_1337 (O_1337,N_23439,N_22725);
and UO_1338 (O_1338,N_24769,N_24518);
nor UO_1339 (O_1339,N_22824,N_24666);
and UO_1340 (O_1340,N_23693,N_23285);
nand UO_1341 (O_1341,N_24320,N_24731);
xnor UO_1342 (O_1342,N_24565,N_24981);
and UO_1343 (O_1343,N_23055,N_24133);
xnor UO_1344 (O_1344,N_23624,N_23982);
nand UO_1345 (O_1345,N_23592,N_22763);
and UO_1346 (O_1346,N_24826,N_24702);
nand UO_1347 (O_1347,N_23711,N_22716);
and UO_1348 (O_1348,N_23812,N_23836);
xnor UO_1349 (O_1349,N_24046,N_24470);
nor UO_1350 (O_1350,N_23962,N_24953);
nor UO_1351 (O_1351,N_22590,N_24164);
or UO_1352 (O_1352,N_23214,N_23439);
nor UO_1353 (O_1353,N_23652,N_23371);
and UO_1354 (O_1354,N_24548,N_23401);
or UO_1355 (O_1355,N_23529,N_22857);
xor UO_1356 (O_1356,N_23334,N_23660);
and UO_1357 (O_1357,N_24686,N_24986);
nand UO_1358 (O_1358,N_23802,N_24022);
nand UO_1359 (O_1359,N_24112,N_22685);
nor UO_1360 (O_1360,N_22793,N_23826);
xor UO_1361 (O_1361,N_22969,N_24201);
or UO_1362 (O_1362,N_24095,N_22863);
nand UO_1363 (O_1363,N_24000,N_23081);
or UO_1364 (O_1364,N_22810,N_24259);
and UO_1365 (O_1365,N_23182,N_23125);
or UO_1366 (O_1366,N_23676,N_23795);
nand UO_1367 (O_1367,N_24393,N_24182);
nor UO_1368 (O_1368,N_24553,N_23144);
and UO_1369 (O_1369,N_24780,N_22971);
xor UO_1370 (O_1370,N_23602,N_24004);
and UO_1371 (O_1371,N_23663,N_23234);
or UO_1372 (O_1372,N_22761,N_23166);
and UO_1373 (O_1373,N_23196,N_24300);
or UO_1374 (O_1374,N_22936,N_22878);
and UO_1375 (O_1375,N_23532,N_24103);
or UO_1376 (O_1376,N_22725,N_22546);
nor UO_1377 (O_1377,N_24241,N_23992);
and UO_1378 (O_1378,N_24855,N_22870);
nand UO_1379 (O_1379,N_23159,N_23217);
nor UO_1380 (O_1380,N_22861,N_22965);
or UO_1381 (O_1381,N_22551,N_23219);
xor UO_1382 (O_1382,N_23032,N_23817);
xor UO_1383 (O_1383,N_23431,N_24316);
xnor UO_1384 (O_1384,N_23906,N_22941);
nor UO_1385 (O_1385,N_23179,N_23107);
nor UO_1386 (O_1386,N_23285,N_23964);
nand UO_1387 (O_1387,N_24993,N_22617);
xor UO_1388 (O_1388,N_22638,N_24615);
and UO_1389 (O_1389,N_22717,N_23400);
and UO_1390 (O_1390,N_24696,N_23851);
or UO_1391 (O_1391,N_24665,N_24182);
and UO_1392 (O_1392,N_23924,N_22571);
nor UO_1393 (O_1393,N_24447,N_24263);
xor UO_1394 (O_1394,N_22509,N_24454);
and UO_1395 (O_1395,N_23765,N_22807);
nor UO_1396 (O_1396,N_24686,N_23459);
xor UO_1397 (O_1397,N_23642,N_23294);
nor UO_1398 (O_1398,N_24968,N_23673);
and UO_1399 (O_1399,N_23789,N_24933);
xnor UO_1400 (O_1400,N_24842,N_24767);
or UO_1401 (O_1401,N_23522,N_22695);
nand UO_1402 (O_1402,N_24607,N_22533);
or UO_1403 (O_1403,N_22531,N_23055);
nand UO_1404 (O_1404,N_24791,N_23849);
nand UO_1405 (O_1405,N_24702,N_23488);
nand UO_1406 (O_1406,N_24881,N_22585);
nor UO_1407 (O_1407,N_23627,N_24436);
nor UO_1408 (O_1408,N_24986,N_24815);
nor UO_1409 (O_1409,N_24424,N_24707);
nor UO_1410 (O_1410,N_24186,N_22768);
or UO_1411 (O_1411,N_23737,N_22969);
xor UO_1412 (O_1412,N_24537,N_22742);
xor UO_1413 (O_1413,N_23495,N_23267);
or UO_1414 (O_1414,N_23040,N_22869);
nand UO_1415 (O_1415,N_23366,N_23809);
xnor UO_1416 (O_1416,N_24845,N_22757);
nor UO_1417 (O_1417,N_23732,N_23696);
nor UO_1418 (O_1418,N_24171,N_23005);
nor UO_1419 (O_1419,N_23050,N_24267);
nor UO_1420 (O_1420,N_23541,N_22894);
or UO_1421 (O_1421,N_24128,N_24804);
nor UO_1422 (O_1422,N_23095,N_22877);
nor UO_1423 (O_1423,N_23499,N_22789);
nand UO_1424 (O_1424,N_23417,N_23054);
and UO_1425 (O_1425,N_23503,N_23268);
and UO_1426 (O_1426,N_24414,N_22771);
xor UO_1427 (O_1427,N_23211,N_24428);
or UO_1428 (O_1428,N_23902,N_23247);
and UO_1429 (O_1429,N_22970,N_23400);
nand UO_1430 (O_1430,N_24907,N_23592);
and UO_1431 (O_1431,N_23029,N_22588);
xnor UO_1432 (O_1432,N_23926,N_22740);
and UO_1433 (O_1433,N_23090,N_24496);
and UO_1434 (O_1434,N_23145,N_23631);
nand UO_1435 (O_1435,N_24573,N_23226);
nor UO_1436 (O_1436,N_24621,N_23234);
nor UO_1437 (O_1437,N_24497,N_22855);
or UO_1438 (O_1438,N_24652,N_24130);
nor UO_1439 (O_1439,N_23771,N_23263);
nand UO_1440 (O_1440,N_23580,N_22628);
nand UO_1441 (O_1441,N_23906,N_24395);
nand UO_1442 (O_1442,N_22762,N_23874);
and UO_1443 (O_1443,N_24858,N_24447);
nor UO_1444 (O_1444,N_24710,N_23625);
nand UO_1445 (O_1445,N_24822,N_24255);
or UO_1446 (O_1446,N_24139,N_23371);
nor UO_1447 (O_1447,N_24849,N_24909);
or UO_1448 (O_1448,N_24496,N_23777);
nand UO_1449 (O_1449,N_24048,N_23812);
xor UO_1450 (O_1450,N_23534,N_24848);
nand UO_1451 (O_1451,N_24658,N_24099);
xor UO_1452 (O_1452,N_23386,N_22763);
nor UO_1453 (O_1453,N_23431,N_24988);
xnor UO_1454 (O_1454,N_23584,N_22658);
or UO_1455 (O_1455,N_23926,N_22867);
and UO_1456 (O_1456,N_24871,N_24560);
nor UO_1457 (O_1457,N_23896,N_24781);
nand UO_1458 (O_1458,N_24841,N_22644);
nand UO_1459 (O_1459,N_24175,N_23174);
and UO_1460 (O_1460,N_23630,N_24030);
or UO_1461 (O_1461,N_23654,N_24371);
nand UO_1462 (O_1462,N_22784,N_23534);
or UO_1463 (O_1463,N_22523,N_23897);
or UO_1464 (O_1464,N_23352,N_24855);
or UO_1465 (O_1465,N_24368,N_23922);
and UO_1466 (O_1466,N_22733,N_23003);
or UO_1467 (O_1467,N_24823,N_24449);
and UO_1468 (O_1468,N_23000,N_22530);
and UO_1469 (O_1469,N_24931,N_22869);
or UO_1470 (O_1470,N_23994,N_22885);
nor UO_1471 (O_1471,N_24662,N_22987);
and UO_1472 (O_1472,N_24020,N_24379);
or UO_1473 (O_1473,N_23761,N_23217);
nand UO_1474 (O_1474,N_24766,N_24893);
nor UO_1475 (O_1475,N_23609,N_22730);
xor UO_1476 (O_1476,N_23439,N_24370);
or UO_1477 (O_1477,N_23091,N_22830);
nand UO_1478 (O_1478,N_22946,N_24435);
xnor UO_1479 (O_1479,N_24893,N_23654);
and UO_1480 (O_1480,N_23275,N_24207);
nand UO_1481 (O_1481,N_24966,N_24513);
or UO_1482 (O_1482,N_24861,N_23326);
nor UO_1483 (O_1483,N_24979,N_22666);
or UO_1484 (O_1484,N_24998,N_22821);
and UO_1485 (O_1485,N_22743,N_24329);
or UO_1486 (O_1486,N_23610,N_23786);
nor UO_1487 (O_1487,N_24457,N_23505);
nand UO_1488 (O_1488,N_23025,N_24212);
xor UO_1489 (O_1489,N_24861,N_23660);
nand UO_1490 (O_1490,N_23540,N_24779);
nand UO_1491 (O_1491,N_23619,N_24381);
nand UO_1492 (O_1492,N_24919,N_22772);
and UO_1493 (O_1493,N_22628,N_23084);
nor UO_1494 (O_1494,N_24257,N_23983);
and UO_1495 (O_1495,N_24208,N_23503);
or UO_1496 (O_1496,N_23059,N_22594);
and UO_1497 (O_1497,N_23399,N_23957);
nand UO_1498 (O_1498,N_23744,N_22628);
xnor UO_1499 (O_1499,N_23348,N_24554);
xor UO_1500 (O_1500,N_22952,N_24373);
xor UO_1501 (O_1501,N_22841,N_24108);
nand UO_1502 (O_1502,N_22534,N_24848);
nor UO_1503 (O_1503,N_22507,N_22644);
nand UO_1504 (O_1504,N_24463,N_23583);
nand UO_1505 (O_1505,N_23213,N_23959);
nor UO_1506 (O_1506,N_23081,N_24561);
xnor UO_1507 (O_1507,N_23959,N_24653);
nand UO_1508 (O_1508,N_23217,N_24641);
nor UO_1509 (O_1509,N_24628,N_23573);
xor UO_1510 (O_1510,N_24743,N_24523);
nor UO_1511 (O_1511,N_24888,N_23069);
or UO_1512 (O_1512,N_22876,N_24905);
nor UO_1513 (O_1513,N_23973,N_22542);
and UO_1514 (O_1514,N_23355,N_23170);
or UO_1515 (O_1515,N_24205,N_23693);
or UO_1516 (O_1516,N_23708,N_23736);
nand UO_1517 (O_1517,N_23456,N_23719);
and UO_1518 (O_1518,N_24615,N_23708);
xnor UO_1519 (O_1519,N_24805,N_23065);
and UO_1520 (O_1520,N_23806,N_22526);
and UO_1521 (O_1521,N_24080,N_23525);
nor UO_1522 (O_1522,N_22917,N_24225);
or UO_1523 (O_1523,N_23196,N_23314);
nor UO_1524 (O_1524,N_24641,N_24596);
nand UO_1525 (O_1525,N_24708,N_22661);
xor UO_1526 (O_1526,N_23634,N_22576);
nand UO_1527 (O_1527,N_24556,N_23305);
and UO_1528 (O_1528,N_24665,N_24957);
or UO_1529 (O_1529,N_23128,N_24627);
and UO_1530 (O_1530,N_23012,N_23424);
nand UO_1531 (O_1531,N_22799,N_22512);
and UO_1532 (O_1532,N_23696,N_23594);
nor UO_1533 (O_1533,N_23265,N_24210);
nand UO_1534 (O_1534,N_24111,N_23412);
and UO_1535 (O_1535,N_23124,N_24863);
or UO_1536 (O_1536,N_24112,N_24732);
xnor UO_1537 (O_1537,N_24186,N_23294);
and UO_1538 (O_1538,N_23002,N_22740);
nand UO_1539 (O_1539,N_24819,N_24048);
nand UO_1540 (O_1540,N_22696,N_24519);
nand UO_1541 (O_1541,N_22825,N_24478);
xor UO_1542 (O_1542,N_23505,N_23582);
xor UO_1543 (O_1543,N_23146,N_22779);
and UO_1544 (O_1544,N_22559,N_22827);
xnor UO_1545 (O_1545,N_23520,N_22830);
and UO_1546 (O_1546,N_24705,N_24664);
nand UO_1547 (O_1547,N_24215,N_23153);
and UO_1548 (O_1548,N_23036,N_24665);
nor UO_1549 (O_1549,N_24418,N_24599);
and UO_1550 (O_1550,N_24215,N_24649);
nand UO_1551 (O_1551,N_24162,N_23390);
and UO_1552 (O_1552,N_24277,N_23203);
nor UO_1553 (O_1553,N_23599,N_22538);
and UO_1554 (O_1554,N_24383,N_23112);
nand UO_1555 (O_1555,N_24428,N_24321);
xnor UO_1556 (O_1556,N_24021,N_22821);
nand UO_1557 (O_1557,N_22677,N_23572);
nand UO_1558 (O_1558,N_24748,N_23507);
xnor UO_1559 (O_1559,N_23339,N_24279);
nand UO_1560 (O_1560,N_23492,N_23865);
or UO_1561 (O_1561,N_23632,N_23136);
xor UO_1562 (O_1562,N_22943,N_24898);
nand UO_1563 (O_1563,N_23361,N_22601);
nor UO_1564 (O_1564,N_22641,N_24544);
nand UO_1565 (O_1565,N_23090,N_24199);
nand UO_1566 (O_1566,N_23577,N_23972);
and UO_1567 (O_1567,N_22952,N_23572);
and UO_1568 (O_1568,N_22700,N_23829);
nand UO_1569 (O_1569,N_24194,N_24016);
nor UO_1570 (O_1570,N_22710,N_22515);
or UO_1571 (O_1571,N_24719,N_22689);
xor UO_1572 (O_1572,N_23178,N_23625);
xor UO_1573 (O_1573,N_23850,N_23044);
nand UO_1574 (O_1574,N_23308,N_24361);
nand UO_1575 (O_1575,N_23922,N_22576);
and UO_1576 (O_1576,N_24751,N_23623);
nor UO_1577 (O_1577,N_24930,N_24066);
nor UO_1578 (O_1578,N_22687,N_23236);
nand UO_1579 (O_1579,N_24158,N_23641);
and UO_1580 (O_1580,N_22576,N_23824);
and UO_1581 (O_1581,N_24319,N_23221);
nand UO_1582 (O_1582,N_23190,N_24496);
and UO_1583 (O_1583,N_23634,N_24689);
or UO_1584 (O_1584,N_23069,N_24012);
nor UO_1585 (O_1585,N_24939,N_24452);
or UO_1586 (O_1586,N_24708,N_22589);
and UO_1587 (O_1587,N_23367,N_24875);
and UO_1588 (O_1588,N_23087,N_23172);
nor UO_1589 (O_1589,N_23371,N_23869);
nor UO_1590 (O_1590,N_22832,N_24316);
nand UO_1591 (O_1591,N_23207,N_23486);
nand UO_1592 (O_1592,N_24428,N_24170);
xnor UO_1593 (O_1593,N_23781,N_23626);
nor UO_1594 (O_1594,N_23438,N_22674);
nand UO_1595 (O_1595,N_23676,N_22510);
and UO_1596 (O_1596,N_24181,N_24095);
or UO_1597 (O_1597,N_23258,N_23651);
and UO_1598 (O_1598,N_24018,N_24924);
xor UO_1599 (O_1599,N_24931,N_24348);
xor UO_1600 (O_1600,N_23721,N_23927);
xor UO_1601 (O_1601,N_23248,N_22676);
nor UO_1602 (O_1602,N_23804,N_23155);
and UO_1603 (O_1603,N_24030,N_24161);
or UO_1604 (O_1604,N_23980,N_22824);
nand UO_1605 (O_1605,N_23661,N_24839);
xor UO_1606 (O_1606,N_24242,N_24000);
nand UO_1607 (O_1607,N_22805,N_23922);
or UO_1608 (O_1608,N_23191,N_22794);
xnor UO_1609 (O_1609,N_22690,N_24615);
or UO_1610 (O_1610,N_23692,N_23843);
xnor UO_1611 (O_1611,N_23394,N_23997);
or UO_1612 (O_1612,N_23668,N_24599);
xnor UO_1613 (O_1613,N_22807,N_22775);
nand UO_1614 (O_1614,N_23108,N_22973);
nand UO_1615 (O_1615,N_23224,N_22559);
nor UO_1616 (O_1616,N_22931,N_24055);
or UO_1617 (O_1617,N_24489,N_24235);
nand UO_1618 (O_1618,N_24437,N_23087);
nand UO_1619 (O_1619,N_23116,N_23056);
nor UO_1620 (O_1620,N_24019,N_24857);
nand UO_1621 (O_1621,N_22730,N_24051);
and UO_1622 (O_1622,N_24287,N_23329);
nand UO_1623 (O_1623,N_22653,N_24247);
or UO_1624 (O_1624,N_23482,N_22734);
xor UO_1625 (O_1625,N_22835,N_23773);
or UO_1626 (O_1626,N_24775,N_23569);
xnor UO_1627 (O_1627,N_23265,N_24557);
or UO_1628 (O_1628,N_24457,N_23099);
xnor UO_1629 (O_1629,N_23947,N_24729);
and UO_1630 (O_1630,N_22807,N_23507);
or UO_1631 (O_1631,N_23967,N_23897);
xnor UO_1632 (O_1632,N_24894,N_24159);
and UO_1633 (O_1633,N_22964,N_23662);
nor UO_1634 (O_1634,N_22990,N_24857);
nand UO_1635 (O_1635,N_23703,N_24018);
or UO_1636 (O_1636,N_22693,N_22865);
xnor UO_1637 (O_1637,N_24038,N_23096);
xnor UO_1638 (O_1638,N_23150,N_24210);
nand UO_1639 (O_1639,N_22852,N_23634);
or UO_1640 (O_1640,N_24848,N_23737);
and UO_1641 (O_1641,N_24458,N_24454);
nand UO_1642 (O_1642,N_22589,N_23039);
nor UO_1643 (O_1643,N_24605,N_23623);
xor UO_1644 (O_1644,N_23539,N_24588);
nor UO_1645 (O_1645,N_23422,N_22723);
and UO_1646 (O_1646,N_24736,N_23134);
or UO_1647 (O_1647,N_24591,N_24842);
and UO_1648 (O_1648,N_22925,N_23944);
nand UO_1649 (O_1649,N_23643,N_24036);
nand UO_1650 (O_1650,N_24935,N_23424);
nand UO_1651 (O_1651,N_23881,N_22517);
and UO_1652 (O_1652,N_24683,N_24797);
xor UO_1653 (O_1653,N_23767,N_24039);
or UO_1654 (O_1654,N_23161,N_24335);
nor UO_1655 (O_1655,N_22615,N_24865);
nor UO_1656 (O_1656,N_24702,N_22804);
xnor UO_1657 (O_1657,N_23267,N_22809);
and UO_1658 (O_1658,N_23141,N_22751);
xor UO_1659 (O_1659,N_23353,N_22766);
nor UO_1660 (O_1660,N_23838,N_23355);
xnor UO_1661 (O_1661,N_23918,N_23706);
and UO_1662 (O_1662,N_23805,N_24256);
xnor UO_1663 (O_1663,N_22968,N_22771);
nor UO_1664 (O_1664,N_24975,N_22799);
and UO_1665 (O_1665,N_23206,N_23230);
or UO_1666 (O_1666,N_24718,N_23920);
nand UO_1667 (O_1667,N_23949,N_22594);
and UO_1668 (O_1668,N_24583,N_24832);
xor UO_1669 (O_1669,N_22723,N_24409);
xnor UO_1670 (O_1670,N_24619,N_24598);
xnor UO_1671 (O_1671,N_24602,N_24070);
nor UO_1672 (O_1672,N_22965,N_23019);
and UO_1673 (O_1673,N_22619,N_24635);
nand UO_1674 (O_1674,N_23042,N_24201);
nor UO_1675 (O_1675,N_22713,N_23321);
nor UO_1676 (O_1676,N_23649,N_24582);
nand UO_1677 (O_1677,N_23270,N_24903);
or UO_1678 (O_1678,N_24699,N_23921);
or UO_1679 (O_1679,N_23128,N_24398);
xnor UO_1680 (O_1680,N_23623,N_24416);
or UO_1681 (O_1681,N_23032,N_24164);
and UO_1682 (O_1682,N_23154,N_23443);
or UO_1683 (O_1683,N_24654,N_23709);
nor UO_1684 (O_1684,N_23079,N_23645);
xor UO_1685 (O_1685,N_24431,N_22871);
nor UO_1686 (O_1686,N_24867,N_24289);
or UO_1687 (O_1687,N_23890,N_24618);
xnor UO_1688 (O_1688,N_23975,N_23120);
and UO_1689 (O_1689,N_22895,N_22726);
xnor UO_1690 (O_1690,N_23853,N_24016);
nor UO_1691 (O_1691,N_22916,N_24565);
nand UO_1692 (O_1692,N_24067,N_23380);
nand UO_1693 (O_1693,N_23488,N_22803);
xor UO_1694 (O_1694,N_24096,N_22575);
or UO_1695 (O_1695,N_23131,N_23330);
xor UO_1696 (O_1696,N_22998,N_24439);
or UO_1697 (O_1697,N_23947,N_22990);
xor UO_1698 (O_1698,N_24860,N_23308);
or UO_1699 (O_1699,N_22862,N_23791);
xnor UO_1700 (O_1700,N_23426,N_23133);
nor UO_1701 (O_1701,N_24937,N_23887);
nor UO_1702 (O_1702,N_24149,N_22855);
or UO_1703 (O_1703,N_24223,N_24190);
xnor UO_1704 (O_1704,N_23217,N_22815);
and UO_1705 (O_1705,N_24431,N_24586);
nand UO_1706 (O_1706,N_24917,N_24924);
xnor UO_1707 (O_1707,N_24959,N_23802);
xor UO_1708 (O_1708,N_23052,N_22846);
nand UO_1709 (O_1709,N_24298,N_22769);
xor UO_1710 (O_1710,N_23091,N_22930);
nor UO_1711 (O_1711,N_24607,N_23281);
nand UO_1712 (O_1712,N_22569,N_23746);
xor UO_1713 (O_1713,N_24514,N_24528);
nor UO_1714 (O_1714,N_24980,N_24398);
xor UO_1715 (O_1715,N_24366,N_23733);
nor UO_1716 (O_1716,N_23787,N_22836);
xor UO_1717 (O_1717,N_23602,N_23941);
nand UO_1718 (O_1718,N_23063,N_22813);
nor UO_1719 (O_1719,N_23323,N_24199);
nand UO_1720 (O_1720,N_24767,N_24419);
xor UO_1721 (O_1721,N_22935,N_24042);
or UO_1722 (O_1722,N_23002,N_23631);
xor UO_1723 (O_1723,N_23682,N_23202);
or UO_1724 (O_1724,N_22808,N_24518);
or UO_1725 (O_1725,N_24008,N_24660);
nor UO_1726 (O_1726,N_23247,N_24664);
xor UO_1727 (O_1727,N_24155,N_23877);
xnor UO_1728 (O_1728,N_22877,N_23401);
nand UO_1729 (O_1729,N_24403,N_24715);
and UO_1730 (O_1730,N_24781,N_22688);
nor UO_1731 (O_1731,N_23933,N_22804);
xnor UO_1732 (O_1732,N_23425,N_24177);
nand UO_1733 (O_1733,N_23362,N_22654);
nor UO_1734 (O_1734,N_24933,N_23657);
and UO_1735 (O_1735,N_24806,N_23492);
and UO_1736 (O_1736,N_24060,N_24057);
xor UO_1737 (O_1737,N_23321,N_23919);
nand UO_1738 (O_1738,N_23852,N_23892);
nand UO_1739 (O_1739,N_24956,N_24182);
and UO_1740 (O_1740,N_22649,N_24323);
nor UO_1741 (O_1741,N_23096,N_22594);
or UO_1742 (O_1742,N_24439,N_23534);
or UO_1743 (O_1743,N_22516,N_24651);
nor UO_1744 (O_1744,N_23167,N_22574);
nor UO_1745 (O_1745,N_24143,N_24996);
and UO_1746 (O_1746,N_23524,N_24108);
and UO_1747 (O_1747,N_23422,N_24613);
or UO_1748 (O_1748,N_23510,N_22505);
xor UO_1749 (O_1749,N_22693,N_24820);
and UO_1750 (O_1750,N_24462,N_23584);
xnor UO_1751 (O_1751,N_24291,N_24218);
or UO_1752 (O_1752,N_24081,N_24573);
nand UO_1753 (O_1753,N_23315,N_23219);
nor UO_1754 (O_1754,N_22973,N_23064);
xnor UO_1755 (O_1755,N_24284,N_23923);
and UO_1756 (O_1756,N_24933,N_24165);
nor UO_1757 (O_1757,N_24451,N_24577);
and UO_1758 (O_1758,N_23427,N_23167);
nand UO_1759 (O_1759,N_22814,N_24036);
and UO_1760 (O_1760,N_23374,N_22743);
xor UO_1761 (O_1761,N_24972,N_23015);
or UO_1762 (O_1762,N_24907,N_24787);
xor UO_1763 (O_1763,N_23188,N_23767);
and UO_1764 (O_1764,N_22839,N_23753);
xor UO_1765 (O_1765,N_23454,N_23398);
and UO_1766 (O_1766,N_22573,N_23248);
or UO_1767 (O_1767,N_24518,N_24111);
or UO_1768 (O_1768,N_24505,N_23215);
xnor UO_1769 (O_1769,N_23642,N_23549);
and UO_1770 (O_1770,N_23942,N_22607);
or UO_1771 (O_1771,N_23027,N_22563);
nor UO_1772 (O_1772,N_22967,N_23576);
nand UO_1773 (O_1773,N_24395,N_22694);
xnor UO_1774 (O_1774,N_23519,N_23581);
and UO_1775 (O_1775,N_23048,N_24349);
xor UO_1776 (O_1776,N_24773,N_23599);
xor UO_1777 (O_1777,N_23719,N_24496);
nand UO_1778 (O_1778,N_22877,N_22655);
nor UO_1779 (O_1779,N_22521,N_24912);
and UO_1780 (O_1780,N_23559,N_23759);
nand UO_1781 (O_1781,N_23590,N_24924);
xnor UO_1782 (O_1782,N_22866,N_23667);
nor UO_1783 (O_1783,N_23010,N_24365);
nor UO_1784 (O_1784,N_23451,N_24343);
nand UO_1785 (O_1785,N_22729,N_22647);
nand UO_1786 (O_1786,N_23079,N_24835);
xnor UO_1787 (O_1787,N_23124,N_23004);
nor UO_1788 (O_1788,N_23447,N_23079);
nor UO_1789 (O_1789,N_23581,N_22757);
and UO_1790 (O_1790,N_24651,N_23929);
or UO_1791 (O_1791,N_23368,N_23053);
nor UO_1792 (O_1792,N_23923,N_22874);
nor UO_1793 (O_1793,N_24286,N_22934);
and UO_1794 (O_1794,N_23793,N_22516);
xnor UO_1795 (O_1795,N_23886,N_23467);
or UO_1796 (O_1796,N_22790,N_23983);
nor UO_1797 (O_1797,N_22604,N_23592);
and UO_1798 (O_1798,N_24973,N_24368);
nand UO_1799 (O_1799,N_24785,N_23070);
or UO_1800 (O_1800,N_22761,N_22851);
nand UO_1801 (O_1801,N_23195,N_24599);
xor UO_1802 (O_1802,N_22946,N_23819);
xnor UO_1803 (O_1803,N_23800,N_24461);
nand UO_1804 (O_1804,N_23909,N_24324);
or UO_1805 (O_1805,N_22958,N_23565);
nor UO_1806 (O_1806,N_24429,N_23582);
and UO_1807 (O_1807,N_24979,N_23646);
xnor UO_1808 (O_1808,N_23509,N_24186);
xor UO_1809 (O_1809,N_23813,N_22620);
and UO_1810 (O_1810,N_23305,N_23718);
nor UO_1811 (O_1811,N_22654,N_23443);
nand UO_1812 (O_1812,N_23788,N_22707);
or UO_1813 (O_1813,N_23206,N_22505);
and UO_1814 (O_1814,N_23331,N_23279);
xor UO_1815 (O_1815,N_23307,N_24426);
nand UO_1816 (O_1816,N_22887,N_22539);
nor UO_1817 (O_1817,N_22687,N_22583);
nand UO_1818 (O_1818,N_23817,N_23549);
nor UO_1819 (O_1819,N_22506,N_23576);
xor UO_1820 (O_1820,N_23454,N_24096);
or UO_1821 (O_1821,N_23061,N_22567);
nor UO_1822 (O_1822,N_22500,N_24759);
nand UO_1823 (O_1823,N_23223,N_23312);
xnor UO_1824 (O_1824,N_23077,N_22716);
nor UO_1825 (O_1825,N_23158,N_23679);
xor UO_1826 (O_1826,N_23446,N_24251);
or UO_1827 (O_1827,N_24941,N_24240);
nand UO_1828 (O_1828,N_24045,N_23496);
xnor UO_1829 (O_1829,N_23718,N_23410);
nor UO_1830 (O_1830,N_22534,N_24418);
nor UO_1831 (O_1831,N_24701,N_23511);
nor UO_1832 (O_1832,N_24785,N_24045);
and UO_1833 (O_1833,N_24127,N_24457);
nor UO_1834 (O_1834,N_24857,N_24348);
or UO_1835 (O_1835,N_23733,N_22838);
and UO_1836 (O_1836,N_23084,N_24173);
xnor UO_1837 (O_1837,N_22754,N_22582);
and UO_1838 (O_1838,N_23179,N_22877);
xnor UO_1839 (O_1839,N_23297,N_23838);
xnor UO_1840 (O_1840,N_24670,N_24511);
or UO_1841 (O_1841,N_24506,N_23466);
and UO_1842 (O_1842,N_24886,N_22862);
and UO_1843 (O_1843,N_24991,N_23944);
nand UO_1844 (O_1844,N_24438,N_24607);
or UO_1845 (O_1845,N_24156,N_23321);
nand UO_1846 (O_1846,N_23622,N_24322);
and UO_1847 (O_1847,N_24040,N_24873);
and UO_1848 (O_1848,N_23930,N_23636);
and UO_1849 (O_1849,N_23783,N_23280);
and UO_1850 (O_1850,N_24124,N_23355);
nor UO_1851 (O_1851,N_23318,N_22682);
nor UO_1852 (O_1852,N_24724,N_24556);
and UO_1853 (O_1853,N_23753,N_24085);
and UO_1854 (O_1854,N_23969,N_24293);
nand UO_1855 (O_1855,N_23060,N_24237);
xor UO_1856 (O_1856,N_23363,N_23240);
and UO_1857 (O_1857,N_23430,N_22951);
nand UO_1858 (O_1858,N_23450,N_23134);
nor UO_1859 (O_1859,N_22589,N_24525);
xor UO_1860 (O_1860,N_23009,N_22886);
nand UO_1861 (O_1861,N_22514,N_23703);
nor UO_1862 (O_1862,N_23034,N_23024);
or UO_1863 (O_1863,N_24068,N_24234);
or UO_1864 (O_1864,N_24792,N_22552);
xnor UO_1865 (O_1865,N_24666,N_23904);
nand UO_1866 (O_1866,N_23282,N_24993);
or UO_1867 (O_1867,N_24773,N_22886);
nand UO_1868 (O_1868,N_24028,N_23487);
and UO_1869 (O_1869,N_24931,N_24014);
nor UO_1870 (O_1870,N_23222,N_23879);
or UO_1871 (O_1871,N_23350,N_24947);
nor UO_1872 (O_1872,N_23847,N_24997);
and UO_1873 (O_1873,N_23423,N_23016);
and UO_1874 (O_1874,N_22860,N_22767);
or UO_1875 (O_1875,N_23771,N_23613);
nor UO_1876 (O_1876,N_24881,N_24783);
and UO_1877 (O_1877,N_24926,N_24710);
and UO_1878 (O_1878,N_24676,N_24208);
nand UO_1879 (O_1879,N_23090,N_23207);
nand UO_1880 (O_1880,N_23622,N_23867);
nor UO_1881 (O_1881,N_22651,N_23927);
nand UO_1882 (O_1882,N_23183,N_24453);
or UO_1883 (O_1883,N_24059,N_23158);
nor UO_1884 (O_1884,N_23434,N_24842);
xor UO_1885 (O_1885,N_24925,N_24850);
nand UO_1886 (O_1886,N_22586,N_22608);
nor UO_1887 (O_1887,N_23446,N_22572);
xnor UO_1888 (O_1888,N_24701,N_24060);
or UO_1889 (O_1889,N_22592,N_23069);
nor UO_1890 (O_1890,N_24392,N_22686);
nor UO_1891 (O_1891,N_23404,N_22525);
xor UO_1892 (O_1892,N_24080,N_23035);
nand UO_1893 (O_1893,N_24404,N_24582);
and UO_1894 (O_1894,N_24356,N_22549);
and UO_1895 (O_1895,N_24294,N_24689);
and UO_1896 (O_1896,N_24066,N_23748);
nor UO_1897 (O_1897,N_24327,N_24622);
or UO_1898 (O_1898,N_23631,N_22537);
nor UO_1899 (O_1899,N_23952,N_24373);
xnor UO_1900 (O_1900,N_22632,N_23870);
nor UO_1901 (O_1901,N_24272,N_23415);
nor UO_1902 (O_1902,N_24996,N_24110);
and UO_1903 (O_1903,N_23624,N_23652);
nand UO_1904 (O_1904,N_23980,N_23784);
and UO_1905 (O_1905,N_22789,N_24272);
nand UO_1906 (O_1906,N_24134,N_24030);
nor UO_1907 (O_1907,N_24610,N_24318);
and UO_1908 (O_1908,N_24053,N_23626);
or UO_1909 (O_1909,N_24140,N_24422);
nand UO_1910 (O_1910,N_24385,N_22898);
nand UO_1911 (O_1911,N_24688,N_24905);
nand UO_1912 (O_1912,N_23591,N_23519);
and UO_1913 (O_1913,N_22572,N_22687);
and UO_1914 (O_1914,N_24779,N_23890);
xor UO_1915 (O_1915,N_24506,N_23919);
nor UO_1916 (O_1916,N_24873,N_24846);
nor UO_1917 (O_1917,N_23748,N_22729);
and UO_1918 (O_1918,N_23902,N_23506);
xnor UO_1919 (O_1919,N_23291,N_23915);
or UO_1920 (O_1920,N_24835,N_23872);
xor UO_1921 (O_1921,N_22823,N_24445);
and UO_1922 (O_1922,N_23110,N_24460);
or UO_1923 (O_1923,N_22839,N_22937);
or UO_1924 (O_1924,N_23333,N_24161);
or UO_1925 (O_1925,N_24458,N_24660);
or UO_1926 (O_1926,N_23050,N_24119);
xnor UO_1927 (O_1927,N_24252,N_24249);
nand UO_1928 (O_1928,N_23708,N_24296);
and UO_1929 (O_1929,N_24199,N_24496);
nand UO_1930 (O_1930,N_23301,N_23916);
xor UO_1931 (O_1931,N_22920,N_24148);
nor UO_1932 (O_1932,N_23516,N_23328);
and UO_1933 (O_1933,N_23132,N_24747);
xnor UO_1934 (O_1934,N_22810,N_24433);
or UO_1935 (O_1935,N_23891,N_24593);
or UO_1936 (O_1936,N_24862,N_23985);
or UO_1937 (O_1937,N_24498,N_23991);
xor UO_1938 (O_1938,N_24025,N_23360);
and UO_1939 (O_1939,N_22936,N_23852);
or UO_1940 (O_1940,N_24098,N_23746);
xnor UO_1941 (O_1941,N_22591,N_22827);
xnor UO_1942 (O_1942,N_22551,N_24246);
and UO_1943 (O_1943,N_24738,N_23473);
and UO_1944 (O_1944,N_24911,N_24245);
xnor UO_1945 (O_1945,N_23796,N_23974);
nand UO_1946 (O_1946,N_23086,N_23854);
nand UO_1947 (O_1947,N_22627,N_24285);
xor UO_1948 (O_1948,N_24298,N_23532);
nand UO_1949 (O_1949,N_24973,N_24114);
or UO_1950 (O_1950,N_23512,N_22624);
or UO_1951 (O_1951,N_24210,N_24077);
and UO_1952 (O_1952,N_23919,N_22954);
nor UO_1953 (O_1953,N_22941,N_24674);
or UO_1954 (O_1954,N_23937,N_23998);
nand UO_1955 (O_1955,N_23362,N_24640);
or UO_1956 (O_1956,N_23615,N_24113);
nand UO_1957 (O_1957,N_22925,N_22557);
or UO_1958 (O_1958,N_23505,N_23451);
or UO_1959 (O_1959,N_24554,N_22847);
and UO_1960 (O_1960,N_23484,N_24309);
nand UO_1961 (O_1961,N_24437,N_22536);
and UO_1962 (O_1962,N_24683,N_23014);
and UO_1963 (O_1963,N_24692,N_23397);
or UO_1964 (O_1964,N_23470,N_22992);
or UO_1965 (O_1965,N_22962,N_24036);
nand UO_1966 (O_1966,N_24166,N_22582);
and UO_1967 (O_1967,N_22550,N_23606);
nand UO_1968 (O_1968,N_23802,N_22677);
and UO_1969 (O_1969,N_23294,N_24646);
xor UO_1970 (O_1970,N_22760,N_24750);
nand UO_1971 (O_1971,N_24976,N_23208);
nor UO_1972 (O_1972,N_22579,N_23537);
nor UO_1973 (O_1973,N_22803,N_22597);
nor UO_1974 (O_1974,N_24378,N_23271);
and UO_1975 (O_1975,N_23030,N_23648);
xnor UO_1976 (O_1976,N_24987,N_24454);
xor UO_1977 (O_1977,N_24577,N_24020);
and UO_1978 (O_1978,N_24320,N_23031);
and UO_1979 (O_1979,N_23797,N_23833);
and UO_1980 (O_1980,N_22602,N_23830);
and UO_1981 (O_1981,N_24775,N_23660);
nor UO_1982 (O_1982,N_23333,N_23321);
xor UO_1983 (O_1983,N_24116,N_24545);
xor UO_1984 (O_1984,N_24966,N_24185);
or UO_1985 (O_1985,N_24211,N_23147);
nand UO_1986 (O_1986,N_22862,N_24241);
or UO_1987 (O_1987,N_22604,N_23374);
nand UO_1988 (O_1988,N_23152,N_23680);
nor UO_1989 (O_1989,N_22711,N_23386);
or UO_1990 (O_1990,N_22993,N_22661);
and UO_1991 (O_1991,N_23229,N_23826);
or UO_1992 (O_1992,N_24787,N_23214);
xnor UO_1993 (O_1993,N_23324,N_23273);
xor UO_1994 (O_1994,N_24916,N_22904);
xor UO_1995 (O_1995,N_23155,N_23680);
or UO_1996 (O_1996,N_24409,N_24434);
nand UO_1997 (O_1997,N_23940,N_23175);
or UO_1998 (O_1998,N_23166,N_23845);
or UO_1999 (O_1999,N_24303,N_22645);
and UO_2000 (O_2000,N_24841,N_24419);
and UO_2001 (O_2001,N_23350,N_22938);
nand UO_2002 (O_2002,N_24853,N_22751);
or UO_2003 (O_2003,N_24064,N_22521);
or UO_2004 (O_2004,N_23034,N_23604);
xnor UO_2005 (O_2005,N_23116,N_23512);
and UO_2006 (O_2006,N_24435,N_23474);
or UO_2007 (O_2007,N_24043,N_24415);
nand UO_2008 (O_2008,N_23341,N_22951);
nand UO_2009 (O_2009,N_23422,N_24286);
nor UO_2010 (O_2010,N_24838,N_23363);
and UO_2011 (O_2011,N_23496,N_23153);
and UO_2012 (O_2012,N_24041,N_23622);
or UO_2013 (O_2013,N_23590,N_24310);
nand UO_2014 (O_2014,N_24154,N_23608);
nand UO_2015 (O_2015,N_24491,N_24649);
and UO_2016 (O_2016,N_23891,N_24592);
and UO_2017 (O_2017,N_23534,N_22513);
nand UO_2018 (O_2018,N_23199,N_22820);
nand UO_2019 (O_2019,N_23360,N_24088);
nand UO_2020 (O_2020,N_24852,N_22713);
nand UO_2021 (O_2021,N_23705,N_24802);
xnor UO_2022 (O_2022,N_22745,N_23771);
and UO_2023 (O_2023,N_23138,N_24030);
or UO_2024 (O_2024,N_22526,N_23603);
nor UO_2025 (O_2025,N_23652,N_23559);
nand UO_2026 (O_2026,N_23138,N_23551);
and UO_2027 (O_2027,N_24660,N_23901);
nor UO_2028 (O_2028,N_24388,N_23962);
nor UO_2029 (O_2029,N_23188,N_22785);
xnor UO_2030 (O_2030,N_23584,N_24848);
xor UO_2031 (O_2031,N_23479,N_24649);
nor UO_2032 (O_2032,N_23974,N_24759);
nor UO_2033 (O_2033,N_24337,N_23408);
nor UO_2034 (O_2034,N_24306,N_24940);
xnor UO_2035 (O_2035,N_22816,N_23290);
nor UO_2036 (O_2036,N_24638,N_23591);
or UO_2037 (O_2037,N_22842,N_23372);
nor UO_2038 (O_2038,N_23114,N_24066);
and UO_2039 (O_2039,N_23119,N_24801);
xor UO_2040 (O_2040,N_23793,N_24941);
nand UO_2041 (O_2041,N_22982,N_22949);
nor UO_2042 (O_2042,N_22903,N_24088);
or UO_2043 (O_2043,N_24904,N_23499);
xnor UO_2044 (O_2044,N_24006,N_23044);
or UO_2045 (O_2045,N_23028,N_24244);
xnor UO_2046 (O_2046,N_24410,N_23012);
nor UO_2047 (O_2047,N_23894,N_24441);
or UO_2048 (O_2048,N_24019,N_23860);
xor UO_2049 (O_2049,N_22780,N_23068);
nor UO_2050 (O_2050,N_23766,N_24211);
and UO_2051 (O_2051,N_24486,N_23498);
nand UO_2052 (O_2052,N_23749,N_22624);
and UO_2053 (O_2053,N_24496,N_23352);
or UO_2054 (O_2054,N_23209,N_22656);
nor UO_2055 (O_2055,N_24811,N_24021);
and UO_2056 (O_2056,N_23841,N_22741);
and UO_2057 (O_2057,N_22514,N_23964);
or UO_2058 (O_2058,N_24034,N_23275);
and UO_2059 (O_2059,N_22551,N_24160);
and UO_2060 (O_2060,N_23668,N_23164);
xor UO_2061 (O_2061,N_23745,N_23868);
nor UO_2062 (O_2062,N_23570,N_23785);
xor UO_2063 (O_2063,N_22871,N_24242);
xnor UO_2064 (O_2064,N_23598,N_24548);
nand UO_2065 (O_2065,N_24871,N_22696);
nand UO_2066 (O_2066,N_22598,N_23781);
and UO_2067 (O_2067,N_23882,N_23873);
and UO_2068 (O_2068,N_24087,N_24729);
and UO_2069 (O_2069,N_24477,N_22614);
nor UO_2070 (O_2070,N_24188,N_23299);
and UO_2071 (O_2071,N_22757,N_23784);
nor UO_2072 (O_2072,N_23799,N_23240);
and UO_2073 (O_2073,N_23921,N_22510);
nand UO_2074 (O_2074,N_23130,N_24242);
and UO_2075 (O_2075,N_23027,N_23263);
or UO_2076 (O_2076,N_23264,N_22691);
and UO_2077 (O_2077,N_23196,N_23829);
xor UO_2078 (O_2078,N_24657,N_23402);
or UO_2079 (O_2079,N_22743,N_22970);
and UO_2080 (O_2080,N_24672,N_23864);
nor UO_2081 (O_2081,N_23867,N_24635);
and UO_2082 (O_2082,N_22770,N_24969);
nand UO_2083 (O_2083,N_24758,N_24984);
nand UO_2084 (O_2084,N_24719,N_24603);
or UO_2085 (O_2085,N_24467,N_24293);
nand UO_2086 (O_2086,N_22548,N_24197);
and UO_2087 (O_2087,N_24921,N_24306);
and UO_2088 (O_2088,N_23814,N_22518);
and UO_2089 (O_2089,N_24142,N_24975);
xnor UO_2090 (O_2090,N_24669,N_24677);
nand UO_2091 (O_2091,N_24403,N_23245);
or UO_2092 (O_2092,N_23313,N_24822);
or UO_2093 (O_2093,N_23642,N_24749);
nor UO_2094 (O_2094,N_22661,N_23633);
xor UO_2095 (O_2095,N_23328,N_23582);
and UO_2096 (O_2096,N_22561,N_23430);
or UO_2097 (O_2097,N_22862,N_22707);
or UO_2098 (O_2098,N_24546,N_23478);
xor UO_2099 (O_2099,N_23935,N_23719);
and UO_2100 (O_2100,N_23287,N_23199);
or UO_2101 (O_2101,N_23873,N_24282);
xor UO_2102 (O_2102,N_24145,N_24199);
nand UO_2103 (O_2103,N_22610,N_22581);
xnor UO_2104 (O_2104,N_23405,N_22569);
xnor UO_2105 (O_2105,N_22564,N_24874);
or UO_2106 (O_2106,N_23930,N_24901);
and UO_2107 (O_2107,N_22873,N_23850);
nor UO_2108 (O_2108,N_24028,N_23092);
nor UO_2109 (O_2109,N_24626,N_24353);
nand UO_2110 (O_2110,N_22980,N_23784);
nand UO_2111 (O_2111,N_23262,N_22539);
xor UO_2112 (O_2112,N_24753,N_23524);
and UO_2113 (O_2113,N_23673,N_23893);
nor UO_2114 (O_2114,N_23449,N_23173);
or UO_2115 (O_2115,N_24301,N_24455);
or UO_2116 (O_2116,N_23279,N_24583);
nor UO_2117 (O_2117,N_23347,N_22804);
or UO_2118 (O_2118,N_23443,N_24059);
nor UO_2119 (O_2119,N_23891,N_23246);
xnor UO_2120 (O_2120,N_23644,N_24549);
nand UO_2121 (O_2121,N_23757,N_22798);
nor UO_2122 (O_2122,N_22808,N_23955);
nand UO_2123 (O_2123,N_24649,N_24285);
nand UO_2124 (O_2124,N_23356,N_22907);
nand UO_2125 (O_2125,N_24251,N_23691);
xnor UO_2126 (O_2126,N_22537,N_24431);
xor UO_2127 (O_2127,N_24147,N_24011);
or UO_2128 (O_2128,N_23237,N_22733);
xnor UO_2129 (O_2129,N_22712,N_22777);
nand UO_2130 (O_2130,N_23943,N_24856);
nand UO_2131 (O_2131,N_23823,N_23877);
xnor UO_2132 (O_2132,N_24813,N_24958);
xnor UO_2133 (O_2133,N_22684,N_22898);
and UO_2134 (O_2134,N_23337,N_22826);
nand UO_2135 (O_2135,N_22822,N_24204);
nand UO_2136 (O_2136,N_24585,N_24218);
and UO_2137 (O_2137,N_24676,N_24617);
xnor UO_2138 (O_2138,N_24906,N_22549);
nand UO_2139 (O_2139,N_24392,N_23266);
xor UO_2140 (O_2140,N_23410,N_23118);
and UO_2141 (O_2141,N_23112,N_22884);
and UO_2142 (O_2142,N_24990,N_23057);
nand UO_2143 (O_2143,N_24340,N_22619);
xnor UO_2144 (O_2144,N_23210,N_24144);
xor UO_2145 (O_2145,N_24453,N_23225);
nand UO_2146 (O_2146,N_23931,N_24059);
and UO_2147 (O_2147,N_23358,N_23367);
or UO_2148 (O_2148,N_24839,N_24859);
nor UO_2149 (O_2149,N_23882,N_24062);
and UO_2150 (O_2150,N_24398,N_23808);
nor UO_2151 (O_2151,N_23435,N_24755);
or UO_2152 (O_2152,N_24013,N_24922);
nand UO_2153 (O_2153,N_23601,N_23416);
and UO_2154 (O_2154,N_22501,N_24058);
or UO_2155 (O_2155,N_24678,N_22941);
or UO_2156 (O_2156,N_23122,N_24894);
or UO_2157 (O_2157,N_23299,N_24971);
nor UO_2158 (O_2158,N_23334,N_23800);
or UO_2159 (O_2159,N_22883,N_24693);
nand UO_2160 (O_2160,N_24720,N_23762);
or UO_2161 (O_2161,N_24673,N_24863);
nand UO_2162 (O_2162,N_23987,N_23072);
xor UO_2163 (O_2163,N_24531,N_23670);
xor UO_2164 (O_2164,N_24087,N_24795);
nand UO_2165 (O_2165,N_24985,N_24669);
nor UO_2166 (O_2166,N_24945,N_22735);
or UO_2167 (O_2167,N_22993,N_23562);
and UO_2168 (O_2168,N_23855,N_22540);
and UO_2169 (O_2169,N_23035,N_23603);
xor UO_2170 (O_2170,N_22573,N_23898);
nor UO_2171 (O_2171,N_23765,N_23284);
nand UO_2172 (O_2172,N_23435,N_24465);
nand UO_2173 (O_2173,N_24816,N_24123);
and UO_2174 (O_2174,N_22667,N_23650);
nor UO_2175 (O_2175,N_23690,N_24377);
and UO_2176 (O_2176,N_24363,N_24359);
nand UO_2177 (O_2177,N_24907,N_24103);
and UO_2178 (O_2178,N_23769,N_24239);
or UO_2179 (O_2179,N_23452,N_23415);
nand UO_2180 (O_2180,N_24200,N_24071);
nand UO_2181 (O_2181,N_24600,N_22786);
and UO_2182 (O_2182,N_23191,N_23767);
xor UO_2183 (O_2183,N_22794,N_22929);
xnor UO_2184 (O_2184,N_23936,N_23479);
and UO_2185 (O_2185,N_24577,N_22827);
nand UO_2186 (O_2186,N_23130,N_23437);
nor UO_2187 (O_2187,N_23100,N_23875);
xor UO_2188 (O_2188,N_23290,N_24857);
nor UO_2189 (O_2189,N_24804,N_24223);
nor UO_2190 (O_2190,N_23413,N_22604);
and UO_2191 (O_2191,N_23959,N_24811);
nor UO_2192 (O_2192,N_24411,N_24794);
xor UO_2193 (O_2193,N_23283,N_24787);
xor UO_2194 (O_2194,N_24710,N_23978);
xnor UO_2195 (O_2195,N_24808,N_23730);
or UO_2196 (O_2196,N_24317,N_24931);
and UO_2197 (O_2197,N_22673,N_23141);
nor UO_2198 (O_2198,N_24145,N_24429);
and UO_2199 (O_2199,N_23748,N_22627);
or UO_2200 (O_2200,N_24915,N_24576);
xor UO_2201 (O_2201,N_24306,N_24769);
nor UO_2202 (O_2202,N_24746,N_24154);
nand UO_2203 (O_2203,N_22832,N_24378);
nand UO_2204 (O_2204,N_22678,N_24853);
or UO_2205 (O_2205,N_23587,N_24027);
nor UO_2206 (O_2206,N_23163,N_22787);
xor UO_2207 (O_2207,N_24767,N_22571);
xnor UO_2208 (O_2208,N_23818,N_24128);
nor UO_2209 (O_2209,N_23528,N_23702);
xnor UO_2210 (O_2210,N_24210,N_23176);
and UO_2211 (O_2211,N_23762,N_24001);
xor UO_2212 (O_2212,N_24387,N_23587);
and UO_2213 (O_2213,N_24297,N_23120);
nand UO_2214 (O_2214,N_22522,N_23656);
and UO_2215 (O_2215,N_24945,N_23405);
xnor UO_2216 (O_2216,N_24505,N_22576);
and UO_2217 (O_2217,N_24249,N_24012);
nand UO_2218 (O_2218,N_23019,N_23414);
or UO_2219 (O_2219,N_24852,N_22647);
nand UO_2220 (O_2220,N_22774,N_23610);
xor UO_2221 (O_2221,N_23199,N_24449);
or UO_2222 (O_2222,N_22832,N_24071);
nand UO_2223 (O_2223,N_24521,N_23514);
nor UO_2224 (O_2224,N_24020,N_23424);
or UO_2225 (O_2225,N_24033,N_23353);
nand UO_2226 (O_2226,N_24221,N_22751);
and UO_2227 (O_2227,N_23041,N_24299);
nand UO_2228 (O_2228,N_23492,N_23042);
xor UO_2229 (O_2229,N_23221,N_23826);
xnor UO_2230 (O_2230,N_23294,N_24304);
xor UO_2231 (O_2231,N_23038,N_24170);
or UO_2232 (O_2232,N_24884,N_23239);
xor UO_2233 (O_2233,N_24652,N_23993);
or UO_2234 (O_2234,N_24531,N_24212);
nand UO_2235 (O_2235,N_24299,N_23120);
and UO_2236 (O_2236,N_23655,N_23363);
and UO_2237 (O_2237,N_23326,N_23816);
and UO_2238 (O_2238,N_23289,N_22904);
and UO_2239 (O_2239,N_24654,N_24952);
nor UO_2240 (O_2240,N_23794,N_24725);
or UO_2241 (O_2241,N_23816,N_23561);
or UO_2242 (O_2242,N_23249,N_23408);
or UO_2243 (O_2243,N_22783,N_23451);
xnor UO_2244 (O_2244,N_24872,N_23694);
nor UO_2245 (O_2245,N_23834,N_23287);
nand UO_2246 (O_2246,N_22671,N_24006);
nor UO_2247 (O_2247,N_23534,N_23367);
and UO_2248 (O_2248,N_23974,N_23086);
nor UO_2249 (O_2249,N_24085,N_23712);
nor UO_2250 (O_2250,N_23113,N_24443);
or UO_2251 (O_2251,N_22765,N_24460);
nand UO_2252 (O_2252,N_24023,N_22814);
or UO_2253 (O_2253,N_23138,N_24901);
or UO_2254 (O_2254,N_24818,N_23568);
nor UO_2255 (O_2255,N_23181,N_22566);
xor UO_2256 (O_2256,N_23559,N_24268);
and UO_2257 (O_2257,N_23000,N_22571);
nor UO_2258 (O_2258,N_23345,N_24621);
or UO_2259 (O_2259,N_23508,N_23461);
nand UO_2260 (O_2260,N_22994,N_23543);
nor UO_2261 (O_2261,N_24142,N_23445);
nor UO_2262 (O_2262,N_24677,N_23157);
nand UO_2263 (O_2263,N_23449,N_24739);
xor UO_2264 (O_2264,N_22516,N_23375);
nand UO_2265 (O_2265,N_24313,N_23090);
or UO_2266 (O_2266,N_23943,N_24357);
nand UO_2267 (O_2267,N_24614,N_23063);
or UO_2268 (O_2268,N_23114,N_24203);
nor UO_2269 (O_2269,N_23754,N_24220);
nand UO_2270 (O_2270,N_23082,N_24159);
nor UO_2271 (O_2271,N_23961,N_23951);
xnor UO_2272 (O_2272,N_23550,N_22697);
nand UO_2273 (O_2273,N_24812,N_23180);
nand UO_2274 (O_2274,N_24172,N_23465);
or UO_2275 (O_2275,N_23446,N_24105);
xnor UO_2276 (O_2276,N_24344,N_24710);
xor UO_2277 (O_2277,N_24702,N_24756);
xnor UO_2278 (O_2278,N_23480,N_24115);
xor UO_2279 (O_2279,N_24731,N_22565);
nor UO_2280 (O_2280,N_24833,N_23227);
and UO_2281 (O_2281,N_23959,N_23065);
and UO_2282 (O_2282,N_23881,N_22833);
xor UO_2283 (O_2283,N_22965,N_23011);
nor UO_2284 (O_2284,N_23451,N_22594);
nor UO_2285 (O_2285,N_23352,N_22837);
or UO_2286 (O_2286,N_24687,N_22682);
or UO_2287 (O_2287,N_24339,N_23296);
nor UO_2288 (O_2288,N_24537,N_23457);
or UO_2289 (O_2289,N_22638,N_22650);
and UO_2290 (O_2290,N_23361,N_23363);
and UO_2291 (O_2291,N_23269,N_23664);
xor UO_2292 (O_2292,N_24686,N_22870);
nor UO_2293 (O_2293,N_23392,N_24744);
nor UO_2294 (O_2294,N_22781,N_24532);
xnor UO_2295 (O_2295,N_24506,N_24494);
and UO_2296 (O_2296,N_22558,N_23285);
nand UO_2297 (O_2297,N_23809,N_24138);
xor UO_2298 (O_2298,N_24650,N_24953);
or UO_2299 (O_2299,N_24705,N_24499);
nand UO_2300 (O_2300,N_24302,N_23954);
nand UO_2301 (O_2301,N_24403,N_24836);
nor UO_2302 (O_2302,N_23059,N_24799);
xor UO_2303 (O_2303,N_24817,N_24579);
nor UO_2304 (O_2304,N_24787,N_23871);
xor UO_2305 (O_2305,N_23733,N_23317);
xor UO_2306 (O_2306,N_23174,N_23635);
and UO_2307 (O_2307,N_24384,N_23689);
xnor UO_2308 (O_2308,N_24295,N_24468);
and UO_2309 (O_2309,N_24619,N_23045);
and UO_2310 (O_2310,N_23978,N_24087);
or UO_2311 (O_2311,N_22905,N_24129);
and UO_2312 (O_2312,N_24480,N_24243);
or UO_2313 (O_2313,N_24960,N_23106);
and UO_2314 (O_2314,N_23486,N_22883);
and UO_2315 (O_2315,N_23510,N_24657);
xor UO_2316 (O_2316,N_24313,N_23641);
or UO_2317 (O_2317,N_23136,N_22700);
or UO_2318 (O_2318,N_23991,N_22600);
nand UO_2319 (O_2319,N_24773,N_24262);
xnor UO_2320 (O_2320,N_23042,N_24834);
nor UO_2321 (O_2321,N_24007,N_23515);
xnor UO_2322 (O_2322,N_24601,N_23676);
nand UO_2323 (O_2323,N_23075,N_23518);
nand UO_2324 (O_2324,N_23174,N_23097);
or UO_2325 (O_2325,N_24007,N_23812);
and UO_2326 (O_2326,N_24976,N_24999);
xnor UO_2327 (O_2327,N_23761,N_24656);
or UO_2328 (O_2328,N_24022,N_24907);
nand UO_2329 (O_2329,N_24534,N_23061);
or UO_2330 (O_2330,N_24059,N_24693);
nor UO_2331 (O_2331,N_23250,N_23587);
or UO_2332 (O_2332,N_24057,N_23378);
xor UO_2333 (O_2333,N_22699,N_22859);
nor UO_2334 (O_2334,N_23516,N_24810);
nand UO_2335 (O_2335,N_24481,N_23192);
nand UO_2336 (O_2336,N_22987,N_23710);
and UO_2337 (O_2337,N_23363,N_24332);
nand UO_2338 (O_2338,N_24523,N_23676);
nor UO_2339 (O_2339,N_22584,N_24051);
nor UO_2340 (O_2340,N_24884,N_23832);
and UO_2341 (O_2341,N_22506,N_24729);
nand UO_2342 (O_2342,N_23371,N_24119);
nor UO_2343 (O_2343,N_24454,N_23839);
nand UO_2344 (O_2344,N_23906,N_22677);
or UO_2345 (O_2345,N_23061,N_23898);
and UO_2346 (O_2346,N_22887,N_22582);
and UO_2347 (O_2347,N_22659,N_24648);
xor UO_2348 (O_2348,N_23339,N_24608);
and UO_2349 (O_2349,N_24106,N_24220);
xnor UO_2350 (O_2350,N_23485,N_23404);
nand UO_2351 (O_2351,N_23127,N_24611);
nor UO_2352 (O_2352,N_22752,N_24509);
and UO_2353 (O_2353,N_23403,N_23784);
xnor UO_2354 (O_2354,N_22519,N_24168);
xnor UO_2355 (O_2355,N_24055,N_24750);
nand UO_2356 (O_2356,N_23273,N_23416);
xnor UO_2357 (O_2357,N_22912,N_24996);
nor UO_2358 (O_2358,N_24584,N_24718);
xnor UO_2359 (O_2359,N_24900,N_22635);
nand UO_2360 (O_2360,N_24295,N_23903);
or UO_2361 (O_2361,N_23008,N_23033);
nor UO_2362 (O_2362,N_23737,N_23496);
xor UO_2363 (O_2363,N_22729,N_24681);
or UO_2364 (O_2364,N_24541,N_24172);
nand UO_2365 (O_2365,N_24308,N_22985);
xor UO_2366 (O_2366,N_22800,N_24406);
nand UO_2367 (O_2367,N_24865,N_23856);
or UO_2368 (O_2368,N_24528,N_24238);
xnor UO_2369 (O_2369,N_24056,N_24847);
or UO_2370 (O_2370,N_24872,N_24556);
or UO_2371 (O_2371,N_23652,N_24523);
nand UO_2372 (O_2372,N_23074,N_23168);
nor UO_2373 (O_2373,N_22915,N_23181);
xnor UO_2374 (O_2374,N_24692,N_24323);
nor UO_2375 (O_2375,N_23572,N_22566);
xnor UO_2376 (O_2376,N_23146,N_23409);
xor UO_2377 (O_2377,N_22833,N_22821);
xnor UO_2378 (O_2378,N_23249,N_24217);
nor UO_2379 (O_2379,N_24647,N_24277);
nand UO_2380 (O_2380,N_23533,N_24949);
xor UO_2381 (O_2381,N_24533,N_24146);
and UO_2382 (O_2382,N_23010,N_23185);
nor UO_2383 (O_2383,N_23755,N_23482);
xor UO_2384 (O_2384,N_24967,N_23212);
nand UO_2385 (O_2385,N_24193,N_23813);
or UO_2386 (O_2386,N_23364,N_24124);
xor UO_2387 (O_2387,N_22508,N_22959);
nor UO_2388 (O_2388,N_23612,N_22839);
xor UO_2389 (O_2389,N_23203,N_22914);
and UO_2390 (O_2390,N_24376,N_24226);
nor UO_2391 (O_2391,N_24939,N_24670);
and UO_2392 (O_2392,N_23471,N_23062);
xor UO_2393 (O_2393,N_24887,N_23542);
and UO_2394 (O_2394,N_22637,N_24704);
nand UO_2395 (O_2395,N_24126,N_23132);
and UO_2396 (O_2396,N_24327,N_23380);
nor UO_2397 (O_2397,N_23548,N_22692);
xor UO_2398 (O_2398,N_24919,N_24124);
xnor UO_2399 (O_2399,N_24508,N_23714);
nand UO_2400 (O_2400,N_23619,N_24003);
nand UO_2401 (O_2401,N_24460,N_23823);
nand UO_2402 (O_2402,N_23613,N_22929);
nor UO_2403 (O_2403,N_23248,N_22977);
and UO_2404 (O_2404,N_23260,N_23382);
xnor UO_2405 (O_2405,N_23333,N_22951);
and UO_2406 (O_2406,N_23568,N_23971);
xor UO_2407 (O_2407,N_22820,N_24093);
xnor UO_2408 (O_2408,N_24935,N_23434);
and UO_2409 (O_2409,N_23691,N_23484);
nor UO_2410 (O_2410,N_24177,N_22795);
nor UO_2411 (O_2411,N_23330,N_24396);
nand UO_2412 (O_2412,N_24675,N_24238);
and UO_2413 (O_2413,N_23221,N_23116);
nand UO_2414 (O_2414,N_24896,N_22835);
or UO_2415 (O_2415,N_24196,N_22586);
and UO_2416 (O_2416,N_22686,N_23953);
nor UO_2417 (O_2417,N_24003,N_23277);
and UO_2418 (O_2418,N_23821,N_23420);
xnor UO_2419 (O_2419,N_23021,N_24700);
nand UO_2420 (O_2420,N_23843,N_23874);
xor UO_2421 (O_2421,N_23207,N_22544);
and UO_2422 (O_2422,N_22612,N_22650);
or UO_2423 (O_2423,N_24671,N_23219);
nand UO_2424 (O_2424,N_23644,N_23756);
nor UO_2425 (O_2425,N_23426,N_23788);
and UO_2426 (O_2426,N_23591,N_23088);
and UO_2427 (O_2427,N_22781,N_22630);
or UO_2428 (O_2428,N_24861,N_23092);
xor UO_2429 (O_2429,N_24754,N_23088);
nor UO_2430 (O_2430,N_24017,N_24584);
or UO_2431 (O_2431,N_24110,N_22980);
or UO_2432 (O_2432,N_22821,N_22575);
nor UO_2433 (O_2433,N_24492,N_24696);
xor UO_2434 (O_2434,N_24501,N_24276);
nand UO_2435 (O_2435,N_24176,N_22964);
nand UO_2436 (O_2436,N_24549,N_24551);
or UO_2437 (O_2437,N_22573,N_24541);
and UO_2438 (O_2438,N_24473,N_22917);
nor UO_2439 (O_2439,N_24733,N_24768);
or UO_2440 (O_2440,N_22637,N_23725);
and UO_2441 (O_2441,N_23504,N_23738);
and UO_2442 (O_2442,N_23770,N_23191);
nor UO_2443 (O_2443,N_24069,N_22745);
and UO_2444 (O_2444,N_22944,N_23191);
and UO_2445 (O_2445,N_22841,N_23326);
or UO_2446 (O_2446,N_22549,N_23801);
xnor UO_2447 (O_2447,N_23497,N_23706);
nor UO_2448 (O_2448,N_23518,N_24430);
or UO_2449 (O_2449,N_24681,N_23918);
and UO_2450 (O_2450,N_24731,N_24423);
xnor UO_2451 (O_2451,N_22734,N_23724);
or UO_2452 (O_2452,N_23028,N_23090);
nand UO_2453 (O_2453,N_23083,N_24870);
nand UO_2454 (O_2454,N_24648,N_22684);
and UO_2455 (O_2455,N_23103,N_23746);
nand UO_2456 (O_2456,N_23098,N_24508);
xnor UO_2457 (O_2457,N_23525,N_23945);
nand UO_2458 (O_2458,N_22786,N_24883);
and UO_2459 (O_2459,N_23406,N_22936);
and UO_2460 (O_2460,N_22811,N_23844);
nand UO_2461 (O_2461,N_23694,N_24543);
xnor UO_2462 (O_2462,N_24116,N_24791);
xnor UO_2463 (O_2463,N_23509,N_24945);
xor UO_2464 (O_2464,N_24311,N_24479);
nand UO_2465 (O_2465,N_22975,N_22899);
xnor UO_2466 (O_2466,N_23887,N_24436);
nand UO_2467 (O_2467,N_22529,N_23232);
xnor UO_2468 (O_2468,N_24005,N_22707);
nor UO_2469 (O_2469,N_22946,N_24288);
nor UO_2470 (O_2470,N_23114,N_24874);
and UO_2471 (O_2471,N_24297,N_22858);
nor UO_2472 (O_2472,N_22542,N_22545);
or UO_2473 (O_2473,N_24465,N_23031);
and UO_2474 (O_2474,N_24115,N_23980);
and UO_2475 (O_2475,N_24423,N_24403);
and UO_2476 (O_2476,N_23740,N_23885);
xor UO_2477 (O_2477,N_23849,N_23431);
nand UO_2478 (O_2478,N_24786,N_24619);
or UO_2479 (O_2479,N_22990,N_24046);
nand UO_2480 (O_2480,N_24755,N_22507);
xnor UO_2481 (O_2481,N_22757,N_24417);
and UO_2482 (O_2482,N_24317,N_22554);
and UO_2483 (O_2483,N_22815,N_23507);
nor UO_2484 (O_2484,N_22952,N_23548);
and UO_2485 (O_2485,N_23477,N_24023);
xor UO_2486 (O_2486,N_22777,N_24842);
and UO_2487 (O_2487,N_23592,N_24073);
or UO_2488 (O_2488,N_23852,N_23119);
nor UO_2489 (O_2489,N_24867,N_23895);
or UO_2490 (O_2490,N_23071,N_23035);
xor UO_2491 (O_2491,N_23515,N_23896);
nor UO_2492 (O_2492,N_24163,N_23115);
xnor UO_2493 (O_2493,N_23473,N_22579);
nand UO_2494 (O_2494,N_23781,N_22953);
xor UO_2495 (O_2495,N_23011,N_24275);
xor UO_2496 (O_2496,N_23711,N_24220);
nand UO_2497 (O_2497,N_24693,N_22568);
xor UO_2498 (O_2498,N_23464,N_24651);
and UO_2499 (O_2499,N_24068,N_23455);
nand UO_2500 (O_2500,N_22982,N_23238);
and UO_2501 (O_2501,N_24885,N_22884);
and UO_2502 (O_2502,N_23934,N_23220);
nand UO_2503 (O_2503,N_22712,N_23175);
or UO_2504 (O_2504,N_24158,N_24470);
or UO_2505 (O_2505,N_24037,N_24166);
nor UO_2506 (O_2506,N_23880,N_24522);
nor UO_2507 (O_2507,N_23071,N_22831);
xor UO_2508 (O_2508,N_24086,N_22932);
or UO_2509 (O_2509,N_22571,N_23814);
nand UO_2510 (O_2510,N_23410,N_23377);
and UO_2511 (O_2511,N_22541,N_23261);
and UO_2512 (O_2512,N_23262,N_23566);
xnor UO_2513 (O_2513,N_24914,N_22531);
nand UO_2514 (O_2514,N_22616,N_24800);
xnor UO_2515 (O_2515,N_23767,N_23979);
nor UO_2516 (O_2516,N_24655,N_24432);
nor UO_2517 (O_2517,N_23844,N_24233);
nand UO_2518 (O_2518,N_23095,N_23841);
and UO_2519 (O_2519,N_24267,N_24505);
xnor UO_2520 (O_2520,N_24862,N_24757);
nand UO_2521 (O_2521,N_24081,N_23935);
xnor UO_2522 (O_2522,N_22712,N_23752);
xor UO_2523 (O_2523,N_22825,N_22777);
xor UO_2524 (O_2524,N_24875,N_22833);
and UO_2525 (O_2525,N_23761,N_22702);
or UO_2526 (O_2526,N_22629,N_22840);
nand UO_2527 (O_2527,N_24681,N_24113);
and UO_2528 (O_2528,N_22904,N_23063);
nor UO_2529 (O_2529,N_24697,N_23659);
or UO_2530 (O_2530,N_24086,N_24362);
xnor UO_2531 (O_2531,N_23853,N_23485);
or UO_2532 (O_2532,N_24104,N_24653);
nor UO_2533 (O_2533,N_22689,N_24017);
and UO_2534 (O_2534,N_23392,N_24622);
and UO_2535 (O_2535,N_23399,N_24030);
and UO_2536 (O_2536,N_22826,N_24643);
and UO_2537 (O_2537,N_22654,N_24986);
nand UO_2538 (O_2538,N_22821,N_22945);
xor UO_2539 (O_2539,N_24633,N_24273);
or UO_2540 (O_2540,N_22833,N_24622);
or UO_2541 (O_2541,N_22755,N_23091);
nand UO_2542 (O_2542,N_23184,N_23264);
or UO_2543 (O_2543,N_22564,N_24946);
nand UO_2544 (O_2544,N_23751,N_23673);
or UO_2545 (O_2545,N_24439,N_24098);
xnor UO_2546 (O_2546,N_23473,N_23993);
nor UO_2547 (O_2547,N_24059,N_23715);
nor UO_2548 (O_2548,N_22916,N_23799);
nor UO_2549 (O_2549,N_23144,N_24552);
nand UO_2550 (O_2550,N_22938,N_22807);
or UO_2551 (O_2551,N_24334,N_24061);
xor UO_2552 (O_2552,N_24788,N_23373);
nor UO_2553 (O_2553,N_23704,N_24925);
or UO_2554 (O_2554,N_24364,N_24958);
xnor UO_2555 (O_2555,N_23720,N_24449);
nor UO_2556 (O_2556,N_24453,N_24112);
or UO_2557 (O_2557,N_24686,N_24642);
nand UO_2558 (O_2558,N_24459,N_24345);
nor UO_2559 (O_2559,N_23912,N_23828);
or UO_2560 (O_2560,N_23039,N_24441);
nor UO_2561 (O_2561,N_23418,N_22631);
or UO_2562 (O_2562,N_23263,N_23366);
xnor UO_2563 (O_2563,N_23774,N_22585);
xor UO_2564 (O_2564,N_24583,N_24071);
nor UO_2565 (O_2565,N_22920,N_22590);
or UO_2566 (O_2566,N_24041,N_24249);
and UO_2567 (O_2567,N_24692,N_24420);
nand UO_2568 (O_2568,N_24320,N_23342);
nor UO_2569 (O_2569,N_23232,N_22598);
and UO_2570 (O_2570,N_24009,N_24073);
nand UO_2571 (O_2571,N_24192,N_24510);
and UO_2572 (O_2572,N_22569,N_22961);
nor UO_2573 (O_2573,N_23156,N_22618);
nor UO_2574 (O_2574,N_23864,N_23961);
nor UO_2575 (O_2575,N_23880,N_23558);
nor UO_2576 (O_2576,N_22953,N_23227);
nand UO_2577 (O_2577,N_23129,N_24861);
and UO_2578 (O_2578,N_23849,N_22895);
or UO_2579 (O_2579,N_22833,N_23659);
and UO_2580 (O_2580,N_23172,N_23474);
or UO_2581 (O_2581,N_23499,N_23524);
and UO_2582 (O_2582,N_24902,N_24222);
nor UO_2583 (O_2583,N_23351,N_22546);
and UO_2584 (O_2584,N_23164,N_23947);
xor UO_2585 (O_2585,N_23085,N_22971);
and UO_2586 (O_2586,N_22893,N_24030);
and UO_2587 (O_2587,N_22752,N_24620);
or UO_2588 (O_2588,N_24133,N_24141);
and UO_2589 (O_2589,N_23009,N_22801);
and UO_2590 (O_2590,N_22638,N_24318);
and UO_2591 (O_2591,N_23449,N_23730);
or UO_2592 (O_2592,N_24393,N_24932);
nor UO_2593 (O_2593,N_24362,N_24336);
nor UO_2594 (O_2594,N_23975,N_22546);
nand UO_2595 (O_2595,N_23971,N_23174);
and UO_2596 (O_2596,N_23916,N_24675);
nor UO_2597 (O_2597,N_23731,N_24279);
nand UO_2598 (O_2598,N_23777,N_24705);
nand UO_2599 (O_2599,N_24582,N_24959);
xnor UO_2600 (O_2600,N_23073,N_23254);
nand UO_2601 (O_2601,N_23923,N_24838);
and UO_2602 (O_2602,N_24184,N_22909);
nor UO_2603 (O_2603,N_23919,N_23114);
xnor UO_2604 (O_2604,N_22876,N_24716);
nand UO_2605 (O_2605,N_23344,N_22610);
or UO_2606 (O_2606,N_22667,N_23943);
xor UO_2607 (O_2607,N_23989,N_23005);
nand UO_2608 (O_2608,N_23803,N_24221);
nor UO_2609 (O_2609,N_22857,N_23180);
or UO_2610 (O_2610,N_24275,N_24627);
or UO_2611 (O_2611,N_24321,N_23674);
nor UO_2612 (O_2612,N_24100,N_23955);
or UO_2613 (O_2613,N_24886,N_24528);
and UO_2614 (O_2614,N_24802,N_24480);
xnor UO_2615 (O_2615,N_24423,N_24723);
xor UO_2616 (O_2616,N_23499,N_22935);
or UO_2617 (O_2617,N_22731,N_23344);
nor UO_2618 (O_2618,N_24397,N_22910);
or UO_2619 (O_2619,N_24654,N_24915);
nand UO_2620 (O_2620,N_23809,N_24598);
nor UO_2621 (O_2621,N_23662,N_22671);
nand UO_2622 (O_2622,N_23785,N_24927);
nand UO_2623 (O_2623,N_24150,N_23813);
nand UO_2624 (O_2624,N_23571,N_24909);
xor UO_2625 (O_2625,N_22751,N_23258);
xor UO_2626 (O_2626,N_24970,N_23934);
and UO_2627 (O_2627,N_24981,N_24808);
nor UO_2628 (O_2628,N_22774,N_24578);
nand UO_2629 (O_2629,N_23736,N_24220);
nor UO_2630 (O_2630,N_23135,N_23920);
or UO_2631 (O_2631,N_24544,N_23200);
nor UO_2632 (O_2632,N_23723,N_24227);
nand UO_2633 (O_2633,N_24663,N_24373);
nor UO_2634 (O_2634,N_22501,N_24122);
nor UO_2635 (O_2635,N_22501,N_24526);
nor UO_2636 (O_2636,N_24443,N_24257);
xnor UO_2637 (O_2637,N_24192,N_24314);
xor UO_2638 (O_2638,N_24643,N_24031);
and UO_2639 (O_2639,N_23688,N_23193);
and UO_2640 (O_2640,N_23613,N_23671);
nand UO_2641 (O_2641,N_23619,N_22975);
or UO_2642 (O_2642,N_24146,N_24032);
and UO_2643 (O_2643,N_23790,N_24061);
or UO_2644 (O_2644,N_23179,N_22649);
nor UO_2645 (O_2645,N_23180,N_23598);
or UO_2646 (O_2646,N_23918,N_24444);
xnor UO_2647 (O_2647,N_22579,N_24806);
and UO_2648 (O_2648,N_23703,N_24061);
and UO_2649 (O_2649,N_23121,N_22891);
and UO_2650 (O_2650,N_24222,N_22888);
or UO_2651 (O_2651,N_23982,N_23820);
or UO_2652 (O_2652,N_23326,N_23917);
nor UO_2653 (O_2653,N_23366,N_22647);
and UO_2654 (O_2654,N_23080,N_24953);
or UO_2655 (O_2655,N_22659,N_22736);
or UO_2656 (O_2656,N_23400,N_24991);
and UO_2657 (O_2657,N_22576,N_23730);
or UO_2658 (O_2658,N_23499,N_22787);
nand UO_2659 (O_2659,N_24704,N_24629);
xor UO_2660 (O_2660,N_23991,N_24632);
nor UO_2661 (O_2661,N_23848,N_23611);
and UO_2662 (O_2662,N_24426,N_23644);
xor UO_2663 (O_2663,N_24555,N_23215);
xnor UO_2664 (O_2664,N_23933,N_22915);
xnor UO_2665 (O_2665,N_22535,N_24948);
xnor UO_2666 (O_2666,N_23385,N_22970);
or UO_2667 (O_2667,N_24786,N_22837);
xor UO_2668 (O_2668,N_24814,N_23380);
xnor UO_2669 (O_2669,N_24164,N_23328);
or UO_2670 (O_2670,N_23378,N_24653);
and UO_2671 (O_2671,N_24176,N_24940);
nor UO_2672 (O_2672,N_23698,N_22622);
nor UO_2673 (O_2673,N_22613,N_24713);
or UO_2674 (O_2674,N_24544,N_23183);
nand UO_2675 (O_2675,N_24941,N_24610);
nor UO_2676 (O_2676,N_24373,N_23149);
or UO_2677 (O_2677,N_23620,N_23059);
xnor UO_2678 (O_2678,N_24813,N_23961);
or UO_2679 (O_2679,N_23041,N_22548);
xnor UO_2680 (O_2680,N_23726,N_23763);
xnor UO_2681 (O_2681,N_23899,N_24735);
nor UO_2682 (O_2682,N_24259,N_22964);
nor UO_2683 (O_2683,N_24052,N_24556);
xor UO_2684 (O_2684,N_22964,N_23589);
nand UO_2685 (O_2685,N_24090,N_24172);
nor UO_2686 (O_2686,N_24672,N_22724);
nand UO_2687 (O_2687,N_23888,N_24254);
and UO_2688 (O_2688,N_23934,N_23963);
nand UO_2689 (O_2689,N_23042,N_23570);
xor UO_2690 (O_2690,N_24349,N_23471);
nor UO_2691 (O_2691,N_23174,N_24800);
xnor UO_2692 (O_2692,N_24195,N_22951);
or UO_2693 (O_2693,N_24156,N_24349);
nand UO_2694 (O_2694,N_22532,N_23479);
nor UO_2695 (O_2695,N_22785,N_24681);
nand UO_2696 (O_2696,N_22957,N_24652);
nand UO_2697 (O_2697,N_24860,N_22725);
nor UO_2698 (O_2698,N_24059,N_23151);
xor UO_2699 (O_2699,N_23375,N_24139);
or UO_2700 (O_2700,N_24524,N_24810);
and UO_2701 (O_2701,N_24503,N_23036);
or UO_2702 (O_2702,N_23890,N_23174);
nor UO_2703 (O_2703,N_24883,N_23510);
or UO_2704 (O_2704,N_23825,N_24842);
nor UO_2705 (O_2705,N_24823,N_23555);
nand UO_2706 (O_2706,N_23812,N_24877);
and UO_2707 (O_2707,N_23397,N_23522);
nor UO_2708 (O_2708,N_23010,N_24287);
or UO_2709 (O_2709,N_23558,N_24261);
xnor UO_2710 (O_2710,N_24487,N_23814);
nor UO_2711 (O_2711,N_24238,N_24174);
nor UO_2712 (O_2712,N_24384,N_24135);
nor UO_2713 (O_2713,N_24352,N_24372);
xnor UO_2714 (O_2714,N_22684,N_24167);
nand UO_2715 (O_2715,N_22534,N_23191);
xor UO_2716 (O_2716,N_24832,N_24167);
and UO_2717 (O_2717,N_23605,N_22833);
and UO_2718 (O_2718,N_22982,N_23800);
xor UO_2719 (O_2719,N_24007,N_22798);
nand UO_2720 (O_2720,N_23111,N_22730);
or UO_2721 (O_2721,N_22637,N_23196);
and UO_2722 (O_2722,N_24646,N_24558);
xor UO_2723 (O_2723,N_23907,N_24422);
and UO_2724 (O_2724,N_24401,N_23149);
and UO_2725 (O_2725,N_24493,N_24439);
and UO_2726 (O_2726,N_23276,N_24133);
nor UO_2727 (O_2727,N_23368,N_23856);
xor UO_2728 (O_2728,N_24554,N_23488);
and UO_2729 (O_2729,N_22970,N_22880);
nand UO_2730 (O_2730,N_23675,N_24410);
or UO_2731 (O_2731,N_23389,N_23833);
nor UO_2732 (O_2732,N_24072,N_24380);
and UO_2733 (O_2733,N_24296,N_23876);
or UO_2734 (O_2734,N_23700,N_22922);
and UO_2735 (O_2735,N_24866,N_23070);
nor UO_2736 (O_2736,N_23854,N_23294);
nand UO_2737 (O_2737,N_23781,N_22514);
xnor UO_2738 (O_2738,N_22677,N_23115);
xnor UO_2739 (O_2739,N_24007,N_24421);
nand UO_2740 (O_2740,N_22738,N_23894);
xnor UO_2741 (O_2741,N_22952,N_24264);
nand UO_2742 (O_2742,N_23458,N_23598);
and UO_2743 (O_2743,N_22813,N_22843);
or UO_2744 (O_2744,N_24878,N_23176);
xnor UO_2745 (O_2745,N_24237,N_23977);
or UO_2746 (O_2746,N_23451,N_22821);
nor UO_2747 (O_2747,N_24712,N_24264);
nand UO_2748 (O_2748,N_23978,N_23030);
nor UO_2749 (O_2749,N_24417,N_24232);
xor UO_2750 (O_2750,N_24377,N_23393);
xor UO_2751 (O_2751,N_23106,N_22513);
and UO_2752 (O_2752,N_24689,N_22558);
or UO_2753 (O_2753,N_23858,N_24267);
or UO_2754 (O_2754,N_23707,N_22649);
nand UO_2755 (O_2755,N_24397,N_23744);
xor UO_2756 (O_2756,N_22949,N_24021);
and UO_2757 (O_2757,N_24482,N_23813);
or UO_2758 (O_2758,N_24781,N_24945);
nor UO_2759 (O_2759,N_24260,N_24188);
or UO_2760 (O_2760,N_23050,N_23340);
nor UO_2761 (O_2761,N_23811,N_23893);
nor UO_2762 (O_2762,N_22810,N_23607);
and UO_2763 (O_2763,N_24377,N_22788);
or UO_2764 (O_2764,N_24938,N_23273);
nor UO_2765 (O_2765,N_24231,N_23960);
nand UO_2766 (O_2766,N_24828,N_24850);
nand UO_2767 (O_2767,N_23871,N_24404);
or UO_2768 (O_2768,N_24645,N_24463);
or UO_2769 (O_2769,N_23696,N_23260);
or UO_2770 (O_2770,N_24843,N_24126);
xnor UO_2771 (O_2771,N_24815,N_23713);
nand UO_2772 (O_2772,N_23042,N_23875);
nand UO_2773 (O_2773,N_23503,N_22670);
xor UO_2774 (O_2774,N_24085,N_24089);
xor UO_2775 (O_2775,N_23373,N_23159);
nor UO_2776 (O_2776,N_23133,N_24133);
nor UO_2777 (O_2777,N_23185,N_23731);
and UO_2778 (O_2778,N_23374,N_23263);
xor UO_2779 (O_2779,N_22647,N_23517);
nor UO_2780 (O_2780,N_24834,N_23632);
and UO_2781 (O_2781,N_24319,N_24839);
xnor UO_2782 (O_2782,N_23839,N_24210);
nor UO_2783 (O_2783,N_22753,N_24188);
nor UO_2784 (O_2784,N_24707,N_24862);
and UO_2785 (O_2785,N_22662,N_22990);
or UO_2786 (O_2786,N_22790,N_23053);
nand UO_2787 (O_2787,N_23033,N_22777);
or UO_2788 (O_2788,N_22527,N_23446);
nand UO_2789 (O_2789,N_23368,N_24445);
xor UO_2790 (O_2790,N_24999,N_23944);
nand UO_2791 (O_2791,N_24328,N_22524);
xor UO_2792 (O_2792,N_23729,N_23860);
or UO_2793 (O_2793,N_24564,N_24587);
or UO_2794 (O_2794,N_23789,N_23359);
nand UO_2795 (O_2795,N_23128,N_23675);
and UO_2796 (O_2796,N_23816,N_23864);
or UO_2797 (O_2797,N_22807,N_22708);
nor UO_2798 (O_2798,N_22836,N_24637);
nor UO_2799 (O_2799,N_24974,N_23335);
xor UO_2800 (O_2800,N_23380,N_24653);
xor UO_2801 (O_2801,N_23451,N_23904);
nor UO_2802 (O_2802,N_23674,N_24583);
or UO_2803 (O_2803,N_23899,N_24169);
or UO_2804 (O_2804,N_24085,N_24926);
nor UO_2805 (O_2805,N_22567,N_24233);
or UO_2806 (O_2806,N_24802,N_24442);
nand UO_2807 (O_2807,N_23346,N_22711);
nand UO_2808 (O_2808,N_22863,N_23459);
and UO_2809 (O_2809,N_24976,N_24598);
xor UO_2810 (O_2810,N_22965,N_24541);
xnor UO_2811 (O_2811,N_23762,N_24113);
or UO_2812 (O_2812,N_23089,N_24540);
nor UO_2813 (O_2813,N_22770,N_24543);
nor UO_2814 (O_2814,N_23430,N_22719);
or UO_2815 (O_2815,N_24162,N_23383);
and UO_2816 (O_2816,N_22632,N_23710);
nand UO_2817 (O_2817,N_24168,N_24354);
nor UO_2818 (O_2818,N_24630,N_23111);
xor UO_2819 (O_2819,N_22569,N_23273);
nand UO_2820 (O_2820,N_23377,N_24669);
nor UO_2821 (O_2821,N_24521,N_23064);
or UO_2822 (O_2822,N_22759,N_24955);
nor UO_2823 (O_2823,N_24014,N_22681);
and UO_2824 (O_2824,N_24594,N_24791);
or UO_2825 (O_2825,N_22984,N_24058);
nor UO_2826 (O_2826,N_24670,N_23798);
xnor UO_2827 (O_2827,N_24847,N_23619);
nor UO_2828 (O_2828,N_24211,N_22876);
or UO_2829 (O_2829,N_23918,N_22918);
nand UO_2830 (O_2830,N_23501,N_24454);
nor UO_2831 (O_2831,N_24113,N_23321);
nor UO_2832 (O_2832,N_24915,N_24587);
or UO_2833 (O_2833,N_24102,N_22588);
nor UO_2834 (O_2834,N_24377,N_24893);
or UO_2835 (O_2835,N_24365,N_24279);
nor UO_2836 (O_2836,N_23621,N_24796);
nand UO_2837 (O_2837,N_24361,N_24572);
nand UO_2838 (O_2838,N_23732,N_24579);
or UO_2839 (O_2839,N_23789,N_23045);
nand UO_2840 (O_2840,N_23463,N_24065);
nor UO_2841 (O_2841,N_24384,N_23238);
or UO_2842 (O_2842,N_24308,N_22827);
and UO_2843 (O_2843,N_22582,N_23752);
and UO_2844 (O_2844,N_24349,N_24813);
xnor UO_2845 (O_2845,N_23787,N_23163);
xor UO_2846 (O_2846,N_23756,N_23381);
nand UO_2847 (O_2847,N_24909,N_24968);
xor UO_2848 (O_2848,N_22880,N_24209);
xnor UO_2849 (O_2849,N_24287,N_22838);
nand UO_2850 (O_2850,N_23608,N_23813);
nand UO_2851 (O_2851,N_22874,N_23774);
or UO_2852 (O_2852,N_23823,N_23232);
xnor UO_2853 (O_2853,N_24153,N_24325);
and UO_2854 (O_2854,N_24635,N_22627);
or UO_2855 (O_2855,N_22651,N_24778);
xnor UO_2856 (O_2856,N_23100,N_23337);
and UO_2857 (O_2857,N_23827,N_23915);
and UO_2858 (O_2858,N_24833,N_23507);
nor UO_2859 (O_2859,N_24239,N_23930);
nor UO_2860 (O_2860,N_22862,N_23892);
nor UO_2861 (O_2861,N_24153,N_23620);
and UO_2862 (O_2862,N_24344,N_24768);
nand UO_2863 (O_2863,N_24474,N_24480);
or UO_2864 (O_2864,N_22696,N_24445);
nor UO_2865 (O_2865,N_23070,N_23572);
and UO_2866 (O_2866,N_22605,N_23032);
xnor UO_2867 (O_2867,N_24934,N_23545);
and UO_2868 (O_2868,N_24693,N_22760);
xor UO_2869 (O_2869,N_24648,N_22629);
nor UO_2870 (O_2870,N_24736,N_24767);
nor UO_2871 (O_2871,N_22557,N_22526);
nor UO_2872 (O_2872,N_24929,N_22784);
nand UO_2873 (O_2873,N_24952,N_23108);
xnor UO_2874 (O_2874,N_24042,N_24387);
nor UO_2875 (O_2875,N_24963,N_24232);
xnor UO_2876 (O_2876,N_24645,N_23203);
nor UO_2877 (O_2877,N_24111,N_22673);
nor UO_2878 (O_2878,N_22890,N_23545);
nand UO_2879 (O_2879,N_23419,N_23504);
xor UO_2880 (O_2880,N_24280,N_23120);
or UO_2881 (O_2881,N_23783,N_23790);
nand UO_2882 (O_2882,N_23001,N_23650);
and UO_2883 (O_2883,N_22575,N_22762);
nand UO_2884 (O_2884,N_24089,N_22759);
xnor UO_2885 (O_2885,N_24832,N_22954);
nand UO_2886 (O_2886,N_24424,N_22692);
or UO_2887 (O_2887,N_22522,N_23807);
nor UO_2888 (O_2888,N_24962,N_22930);
and UO_2889 (O_2889,N_24875,N_23755);
nor UO_2890 (O_2890,N_24307,N_23946);
nand UO_2891 (O_2891,N_24215,N_24861);
xor UO_2892 (O_2892,N_23508,N_24744);
xnor UO_2893 (O_2893,N_22840,N_24138);
or UO_2894 (O_2894,N_22878,N_24342);
nand UO_2895 (O_2895,N_24922,N_23464);
xnor UO_2896 (O_2896,N_24571,N_22695);
and UO_2897 (O_2897,N_23815,N_24166);
or UO_2898 (O_2898,N_24787,N_23540);
and UO_2899 (O_2899,N_23714,N_23541);
xor UO_2900 (O_2900,N_23539,N_23552);
xor UO_2901 (O_2901,N_24358,N_24106);
and UO_2902 (O_2902,N_24573,N_24365);
xor UO_2903 (O_2903,N_22776,N_23412);
nand UO_2904 (O_2904,N_22730,N_23061);
nand UO_2905 (O_2905,N_24675,N_23324);
and UO_2906 (O_2906,N_22734,N_23650);
nor UO_2907 (O_2907,N_22594,N_24938);
and UO_2908 (O_2908,N_24792,N_22897);
or UO_2909 (O_2909,N_23861,N_24893);
and UO_2910 (O_2910,N_24674,N_23575);
xor UO_2911 (O_2911,N_23111,N_22773);
and UO_2912 (O_2912,N_24558,N_24200);
nor UO_2913 (O_2913,N_23397,N_24185);
and UO_2914 (O_2914,N_23069,N_22544);
and UO_2915 (O_2915,N_24400,N_22710);
nand UO_2916 (O_2916,N_24442,N_24940);
nand UO_2917 (O_2917,N_23960,N_23182);
or UO_2918 (O_2918,N_24883,N_23164);
and UO_2919 (O_2919,N_24028,N_23281);
nand UO_2920 (O_2920,N_22916,N_22923);
nand UO_2921 (O_2921,N_24172,N_23850);
nand UO_2922 (O_2922,N_23087,N_24425);
nor UO_2923 (O_2923,N_22614,N_24053);
or UO_2924 (O_2924,N_24855,N_23665);
and UO_2925 (O_2925,N_23161,N_24659);
and UO_2926 (O_2926,N_22567,N_24745);
or UO_2927 (O_2927,N_23988,N_24502);
or UO_2928 (O_2928,N_24064,N_22732);
nand UO_2929 (O_2929,N_24465,N_23428);
nor UO_2930 (O_2930,N_23287,N_23812);
nand UO_2931 (O_2931,N_23676,N_23078);
xnor UO_2932 (O_2932,N_24790,N_24448);
nor UO_2933 (O_2933,N_23945,N_22544);
nor UO_2934 (O_2934,N_24179,N_23382);
xnor UO_2935 (O_2935,N_24292,N_23973);
nor UO_2936 (O_2936,N_24794,N_23311);
nand UO_2937 (O_2937,N_24965,N_24202);
or UO_2938 (O_2938,N_24480,N_22554);
or UO_2939 (O_2939,N_24025,N_23812);
nand UO_2940 (O_2940,N_24744,N_22795);
nor UO_2941 (O_2941,N_22752,N_22524);
or UO_2942 (O_2942,N_22945,N_24968);
xor UO_2943 (O_2943,N_23131,N_24360);
xor UO_2944 (O_2944,N_22597,N_23800);
or UO_2945 (O_2945,N_23867,N_24870);
or UO_2946 (O_2946,N_23947,N_22676);
and UO_2947 (O_2947,N_23443,N_23285);
xor UO_2948 (O_2948,N_24531,N_23818);
xnor UO_2949 (O_2949,N_23079,N_22714);
and UO_2950 (O_2950,N_23756,N_23895);
nor UO_2951 (O_2951,N_23884,N_23831);
or UO_2952 (O_2952,N_23289,N_23161);
nor UO_2953 (O_2953,N_24194,N_23021);
or UO_2954 (O_2954,N_24054,N_23350);
nor UO_2955 (O_2955,N_23889,N_23217);
or UO_2956 (O_2956,N_23389,N_23295);
or UO_2957 (O_2957,N_24446,N_24652);
or UO_2958 (O_2958,N_23728,N_24756);
nand UO_2959 (O_2959,N_23945,N_24876);
or UO_2960 (O_2960,N_24056,N_23578);
xnor UO_2961 (O_2961,N_24471,N_24762);
or UO_2962 (O_2962,N_23061,N_22942);
or UO_2963 (O_2963,N_23987,N_22527);
xor UO_2964 (O_2964,N_23306,N_23737);
or UO_2965 (O_2965,N_24522,N_23570);
nor UO_2966 (O_2966,N_24140,N_24822);
and UO_2967 (O_2967,N_22571,N_24526);
xnor UO_2968 (O_2968,N_24928,N_23251);
nand UO_2969 (O_2969,N_22906,N_24729);
nand UO_2970 (O_2970,N_24600,N_23011);
nand UO_2971 (O_2971,N_24402,N_23400);
or UO_2972 (O_2972,N_24919,N_24307);
xor UO_2973 (O_2973,N_23215,N_23852);
nand UO_2974 (O_2974,N_22695,N_23065);
xnor UO_2975 (O_2975,N_24195,N_22501);
or UO_2976 (O_2976,N_23826,N_24127);
nand UO_2977 (O_2977,N_23982,N_22642);
or UO_2978 (O_2978,N_23111,N_24938);
xor UO_2979 (O_2979,N_23770,N_23606);
xnor UO_2980 (O_2980,N_22934,N_23706);
and UO_2981 (O_2981,N_23865,N_24230);
and UO_2982 (O_2982,N_23911,N_23727);
nand UO_2983 (O_2983,N_22945,N_23211);
and UO_2984 (O_2984,N_23356,N_24445);
or UO_2985 (O_2985,N_24136,N_23160);
xor UO_2986 (O_2986,N_23522,N_24548);
nor UO_2987 (O_2987,N_24684,N_22930);
or UO_2988 (O_2988,N_22598,N_22964);
and UO_2989 (O_2989,N_24725,N_23544);
nor UO_2990 (O_2990,N_22648,N_24588);
or UO_2991 (O_2991,N_22872,N_24467);
nand UO_2992 (O_2992,N_23327,N_23840);
and UO_2993 (O_2993,N_22997,N_24127);
nor UO_2994 (O_2994,N_22856,N_22652);
xnor UO_2995 (O_2995,N_23773,N_23245);
or UO_2996 (O_2996,N_24521,N_24725);
or UO_2997 (O_2997,N_23283,N_23043);
xor UO_2998 (O_2998,N_24417,N_24659);
and UO_2999 (O_2999,N_24122,N_23514);
endmodule