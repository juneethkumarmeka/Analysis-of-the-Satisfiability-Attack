module basic_500_3000_500_50_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_37,In_34);
xnor U1 (N_1,In_156,In_47);
nand U2 (N_2,In_381,In_5);
or U3 (N_3,In_451,In_84);
nand U4 (N_4,In_103,In_295);
nand U5 (N_5,In_127,In_106);
or U6 (N_6,In_361,In_355);
and U7 (N_7,In_120,In_462);
and U8 (N_8,In_291,In_278);
nor U9 (N_9,In_341,In_323);
and U10 (N_10,In_174,In_369);
or U11 (N_11,In_318,In_82);
nand U12 (N_12,In_245,In_170);
and U13 (N_13,In_426,In_439);
nand U14 (N_14,In_296,In_350);
and U15 (N_15,In_403,In_93);
or U16 (N_16,In_219,In_16);
nand U17 (N_17,In_372,In_370);
or U18 (N_18,In_179,In_115);
or U19 (N_19,In_181,In_480);
or U20 (N_20,In_160,In_412);
nand U21 (N_21,In_385,In_119);
xnor U22 (N_22,In_141,In_499);
xor U23 (N_23,In_293,In_66);
or U24 (N_24,In_283,In_70);
nand U25 (N_25,In_69,In_325);
and U26 (N_26,In_228,In_198);
and U27 (N_27,In_236,In_270);
nand U28 (N_28,In_314,In_105);
and U29 (N_29,In_63,In_159);
nand U30 (N_30,In_108,In_216);
and U31 (N_31,In_229,In_334);
nand U32 (N_32,In_64,In_377);
nor U33 (N_33,In_389,In_254);
or U34 (N_34,In_413,In_49);
nand U35 (N_35,In_336,In_60);
or U36 (N_36,In_475,In_476);
nand U37 (N_37,In_315,In_365);
and U38 (N_38,In_279,In_102);
and U39 (N_39,In_186,In_77);
nor U40 (N_40,In_444,In_155);
or U41 (N_41,In_477,In_55);
nand U42 (N_42,In_438,In_153);
and U43 (N_43,In_187,In_422);
and U44 (N_44,In_252,In_137);
and U45 (N_45,In_484,In_392);
or U46 (N_46,In_332,In_429);
nor U47 (N_47,In_235,In_146);
xnor U48 (N_48,In_259,In_405);
nor U49 (N_49,In_195,In_399);
and U50 (N_50,In_7,In_428);
nor U51 (N_51,In_147,In_297);
nor U52 (N_52,In_249,In_189);
xnor U53 (N_53,In_437,In_328);
or U54 (N_54,In_423,In_363);
or U55 (N_55,In_209,In_414);
nand U56 (N_56,In_359,In_465);
or U57 (N_57,In_131,In_220);
or U58 (N_58,In_455,In_497);
xor U59 (N_59,In_339,In_237);
and U60 (N_60,In_255,In_322);
nor U61 (N_61,In_133,In_308);
and U62 (N_62,N_29,In_261);
nor U63 (N_63,In_83,In_408);
and U64 (N_64,In_330,In_267);
or U65 (N_65,In_163,In_118);
nor U66 (N_66,In_194,In_280);
or U67 (N_67,N_9,In_299);
or U68 (N_68,In_498,In_86);
or U69 (N_69,In_394,In_492);
nor U70 (N_70,In_320,In_74);
nor U71 (N_71,N_23,In_391);
nand U72 (N_72,In_446,N_57);
and U73 (N_73,N_1,In_301);
or U74 (N_74,In_264,In_321);
nand U75 (N_75,In_42,In_393);
and U76 (N_76,In_288,In_116);
and U77 (N_77,In_20,In_104);
or U78 (N_78,In_324,In_57);
and U79 (N_79,In_402,In_436);
or U80 (N_80,In_39,In_284);
and U81 (N_81,In_352,In_166);
xor U82 (N_82,In_326,In_274);
nor U83 (N_83,In_425,In_199);
nand U84 (N_84,N_41,In_26);
nor U85 (N_85,In_192,In_300);
and U86 (N_86,N_20,In_313);
or U87 (N_87,In_109,In_117);
or U88 (N_88,In_305,In_184);
nand U89 (N_89,In_79,In_362);
nand U90 (N_90,In_67,In_27);
nor U91 (N_91,N_42,In_483);
or U92 (N_92,In_342,N_8);
or U93 (N_93,In_125,In_65);
or U94 (N_94,N_43,In_230);
or U95 (N_95,In_256,In_58);
and U96 (N_96,In_126,In_317);
nand U97 (N_97,In_474,In_11);
nand U98 (N_98,In_286,In_347);
and U99 (N_99,In_172,In_193);
or U100 (N_100,In_205,In_15);
or U101 (N_101,In_445,In_260);
nor U102 (N_102,In_238,N_18);
nor U103 (N_103,In_373,In_382);
nand U104 (N_104,In_24,In_22);
nor U105 (N_105,In_62,In_466);
nor U106 (N_106,In_387,In_407);
or U107 (N_107,In_6,N_2);
nand U108 (N_108,N_35,In_210);
or U109 (N_109,In_234,N_28);
nand U110 (N_110,In_152,In_178);
nand U111 (N_111,In_99,In_461);
and U112 (N_112,In_398,N_54);
nor U113 (N_113,In_72,In_8);
nand U114 (N_114,In_277,In_247);
nor U115 (N_115,In_447,In_306);
and U116 (N_116,In_167,In_138);
or U117 (N_117,N_26,In_1);
nand U118 (N_118,In_467,In_182);
or U119 (N_119,In_73,In_243);
or U120 (N_120,N_72,In_489);
nand U121 (N_121,In_139,N_84);
nor U122 (N_122,In_95,N_14);
nor U123 (N_123,N_64,In_463);
nand U124 (N_124,N_3,In_143);
nand U125 (N_125,In_397,In_395);
xor U126 (N_126,In_50,In_433);
xnor U127 (N_127,In_4,N_113);
nand U128 (N_128,In_383,In_107);
nor U129 (N_129,In_435,In_168);
nor U130 (N_130,In_345,In_241);
or U131 (N_131,In_418,In_51);
nor U132 (N_132,In_150,In_17);
nor U133 (N_133,N_77,N_118);
or U134 (N_134,In_122,N_37);
or U135 (N_135,In_452,In_424);
nand U136 (N_136,N_101,In_38);
and U137 (N_137,In_176,In_98);
nor U138 (N_138,In_233,In_364);
nor U139 (N_139,N_40,In_43);
and U140 (N_140,In_61,In_396);
nand U141 (N_141,In_188,N_94);
nor U142 (N_142,In_303,N_117);
nand U143 (N_143,In_53,In_269);
nand U144 (N_144,In_248,In_459);
and U145 (N_145,N_33,In_89);
or U146 (N_146,N_51,N_83);
nand U147 (N_147,In_449,In_207);
nand U148 (N_148,In_204,In_427);
nor U149 (N_149,In_78,N_0);
nand U150 (N_150,In_458,In_289);
and U151 (N_151,In_130,In_56);
or U152 (N_152,In_290,N_114);
or U153 (N_153,N_32,In_390);
nand U154 (N_154,In_154,N_89);
xnor U155 (N_155,In_164,In_457);
xor U156 (N_156,N_66,In_46);
or U157 (N_157,N_47,In_97);
and U158 (N_158,In_257,In_36);
or U159 (N_159,In_453,In_351);
and U160 (N_160,In_185,In_276);
or U161 (N_161,In_23,In_374);
nor U162 (N_162,In_333,In_419);
nor U163 (N_163,N_88,In_35);
and U164 (N_164,N_19,In_470);
and U165 (N_165,In_379,In_145);
nor U166 (N_166,In_92,In_353);
nor U167 (N_167,N_24,In_222);
nor U168 (N_168,In_41,In_443);
xor U169 (N_169,In_211,In_460);
nand U170 (N_170,N_25,In_287);
or U171 (N_171,In_409,In_171);
or U172 (N_172,N_50,In_31);
or U173 (N_173,In_265,N_109);
and U174 (N_174,In_226,In_494);
nand U175 (N_175,In_430,In_368);
nand U176 (N_176,In_486,In_48);
or U177 (N_177,In_404,In_273);
nand U178 (N_178,In_215,N_102);
nor U179 (N_179,In_416,In_124);
nor U180 (N_180,In_183,In_140);
xor U181 (N_181,N_160,In_158);
nand U182 (N_182,N_121,N_36);
and U183 (N_183,In_144,N_81);
xor U184 (N_184,N_149,In_358);
xnor U185 (N_185,In_488,In_191);
nor U186 (N_186,In_448,In_263);
and U187 (N_187,N_168,In_173);
nor U188 (N_188,In_169,In_162);
xor U189 (N_189,In_196,In_380);
xor U190 (N_190,N_150,N_38);
and U191 (N_191,N_79,N_126);
or U192 (N_192,N_96,N_98);
and U193 (N_193,In_44,In_68);
xnor U194 (N_194,In_478,N_46);
and U195 (N_195,N_52,N_136);
nor U196 (N_196,In_110,N_110);
or U197 (N_197,N_174,In_2);
nand U198 (N_198,In_479,N_59);
and U199 (N_199,In_354,In_214);
or U200 (N_200,N_45,In_468);
and U201 (N_201,In_440,In_357);
xnor U202 (N_202,In_410,N_49);
or U203 (N_203,N_135,N_91);
nand U204 (N_204,In_203,N_104);
xor U205 (N_205,N_95,N_159);
nor U206 (N_206,N_179,N_156);
or U207 (N_207,In_400,In_90);
and U208 (N_208,N_73,In_9);
nor U209 (N_209,In_100,N_80);
and U210 (N_210,In_246,In_327);
and U211 (N_211,In_456,In_85);
xnor U212 (N_212,In_177,N_106);
and U213 (N_213,In_388,N_157);
and U214 (N_214,In_464,In_384);
nor U215 (N_215,N_134,N_78);
xor U216 (N_216,N_56,N_172);
nand U217 (N_217,In_376,In_201);
or U218 (N_218,N_177,In_135);
and U219 (N_219,In_471,In_490);
and U220 (N_220,N_162,In_329);
and U221 (N_221,In_231,In_253);
and U222 (N_222,N_127,N_10);
nor U223 (N_223,In_111,In_268);
or U224 (N_224,In_485,N_139);
and U225 (N_225,In_493,In_221);
or U226 (N_226,In_190,In_224);
or U227 (N_227,In_496,In_149);
or U228 (N_228,N_155,In_420);
nor U229 (N_229,In_469,In_240);
and U230 (N_230,In_96,In_275);
xor U231 (N_231,N_154,N_152);
nor U232 (N_232,In_87,N_116);
nand U233 (N_233,N_16,N_99);
xor U234 (N_234,In_33,In_218);
and U235 (N_235,N_68,In_3);
and U236 (N_236,N_74,N_145);
nor U237 (N_237,In_442,N_87);
and U238 (N_238,N_133,In_223);
and U239 (N_239,In_319,N_69);
and U240 (N_240,In_32,N_176);
nor U241 (N_241,N_232,N_186);
and U242 (N_242,In_344,N_187);
nor U243 (N_243,In_200,In_304);
and U244 (N_244,In_371,In_285);
nor U245 (N_245,In_40,In_348);
and U246 (N_246,In_421,N_142);
nor U247 (N_247,In_121,N_191);
and U248 (N_248,In_312,In_213);
nand U249 (N_249,N_207,In_142);
or U250 (N_250,N_239,N_163);
nor U251 (N_251,N_131,N_164);
xnor U252 (N_252,In_113,In_175);
or U253 (N_253,N_151,N_211);
or U254 (N_254,N_67,In_29);
or U255 (N_255,N_63,N_61);
or U256 (N_256,In_52,N_30);
nand U257 (N_257,In_91,N_230);
nand U258 (N_258,N_200,In_415);
nor U259 (N_259,In_294,N_238);
nor U260 (N_260,N_148,In_81);
nor U261 (N_261,In_316,N_205);
nor U262 (N_262,N_22,N_4);
and U263 (N_263,N_225,In_482);
nand U264 (N_264,In_206,N_137);
or U265 (N_265,N_11,N_192);
nor U266 (N_266,In_165,N_100);
nand U267 (N_267,N_215,In_310);
or U268 (N_268,In_262,N_34);
xor U269 (N_269,N_115,In_432);
nor U270 (N_270,N_171,In_161);
nor U271 (N_271,In_335,N_138);
nand U272 (N_272,In_45,In_12);
nand U273 (N_273,N_107,N_44);
or U274 (N_274,In_0,N_108);
nand U275 (N_275,In_298,N_226);
nand U276 (N_276,In_212,In_281);
and U277 (N_277,In_367,In_309);
and U278 (N_278,N_233,In_202);
and U279 (N_279,N_132,N_6);
nand U280 (N_280,N_75,In_18);
xnor U281 (N_281,In_378,In_80);
nor U282 (N_282,N_125,In_282);
nand U283 (N_283,In_244,In_251);
or U284 (N_284,In_360,N_224);
and U285 (N_285,N_173,In_30);
nand U286 (N_286,In_134,N_48);
nor U287 (N_287,In_366,N_122);
nand U288 (N_288,In_208,N_93);
xor U289 (N_289,N_141,N_90);
and U290 (N_290,N_198,In_239);
nand U291 (N_291,In_250,N_76);
nor U292 (N_292,N_92,N_216);
xnor U293 (N_293,In_129,N_70);
or U294 (N_294,N_235,N_204);
nand U295 (N_295,N_237,In_10);
nor U296 (N_296,N_55,In_472);
and U297 (N_297,N_129,In_331);
or U298 (N_298,N_123,In_225);
nor U299 (N_299,N_85,N_195);
or U300 (N_300,N_297,In_21);
or U301 (N_301,N_274,N_276);
nand U302 (N_302,N_62,N_58);
or U303 (N_303,In_311,In_157);
or U304 (N_304,N_53,In_13);
or U305 (N_305,N_182,N_120);
nand U306 (N_306,N_294,In_25);
or U307 (N_307,N_252,N_245);
nand U308 (N_308,N_140,N_248);
nor U309 (N_309,N_288,In_495);
nor U310 (N_310,N_254,N_279);
xor U311 (N_311,In_346,N_124);
or U312 (N_312,In_75,In_232);
nor U313 (N_313,N_287,N_203);
or U314 (N_314,N_282,N_263);
or U315 (N_315,N_277,In_28);
nand U316 (N_316,N_169,N_208);
nand U317 (N_317,N_227,N_146);
nand U318 (N_318,In_271,N_218);
nor U319 (N_319,N_247,N_119);
nand U320 (N_320,N_167,In_411);
and U321 (N_321,N_210,N_231);
and U322 (N_322,N_265,N_97);
and U323 (N_323,N_253,N_130);
nand U324 (N_324,N_286,N_242);
or U325 (N_325,N_241,N_273);
or U326 (N_326,N_13,In_128);
and U327 (N_327,N_111,N_293);
nor U328 (N_328,In_54,N_65);
and U329 (N_329,In_227,N_166);
nand U330 (N_330,In_302,N_181);
nand U331 (N_331,N_275,N_266);
nor U332 (N_332,In_123,In_59);
nand U333 (N_333,N_188,N_103);
or U334 (N_334,N_213,In_197);
and U335 (N_335,N_17,N_234);
or U336 (N_336,N_240,N_229);
nand U337 (N_337,In_76,N_5);
nor U338 (N_338,In_258,In_266);
or U339 (N_339,N_283,In_343);
and U340 (N_340,N_249,N_189);
nand U341 (N_341,In_375,N_269);
or U342 (N_342,In_340,N_60);
nor U343 (N_343,N_153,N_219);
xor U344 (N_344,N_259,N_271);
nor U345 (N_345,N_144,N_217);
xor U346 (N_346,N_158,In_386);
and U347 (N_347,N_222,N_184);
and U348 (N_348,In_338,In_491);
nand U349 (N_349,In_148,N_228);
nand U350 (N_350,N_251,N_261);
nor U351 (N_351,In_151,N_243);
and U352 (N_352,N_272,N_175);
or U353 (N_353,N_199,In_180);
xnor U354 (N_354,N_15,N_183);
nand U355 (N_355,N_202,N_255);
or U356 (N_356,N_82,N_270);
nor U357 (N_357,N_201,N_281);
and U358 (N_358,N_291,In_356);
nor U359 (N_359,N_299,N_267);
nand U360 (N_360,N_333,N_170);
xnor U361 (N_361,N_193,N_310);
nand U362 (N_362,N_196,N_359);
nand U363 (N_363,N_334,N_236);
and U364 (N_364,N_340,N_326);
and U365 (N_365,N_312,N_343);
nor U366 (N_366,N_295,N_39);
or U367 (N_367,N_190,In_217);
or U368 (N_368,N_206,In_94);
nand U369 (N_369,N_358,N_320);
nand U370 (N_370,N_319,N_317);
nor U371 (N_371,In_88,In_112);
nand U372 (N_372,N_314,N_313);
or U373 (N_373,In_242,N_262);
and U374 (N_374,N_278,N_285);
nand U375 (N_375,N_244,N_197);
or U376 (N_376,N_307,N_349);
or U377 (N_377,N_344,N_338);
xor U378 (N_378,N_346,N_328);
xor U379 (N_379,N_322,N_357);
and U380 (N_380,In_307,N_143);
xor U381 (N_381,N_327,N_308);
nor U382 (N_382,In_450,In_454);
nor U383 (N_383,N_323,N_180);
or U384 (N_384,N_325,N_348);
nor U385 (N_385,In_19,N_315);
or U386 (N_386,N_27,N_128);
nand U387 (N_387,In_434,N_305);
or U388 (N_388,N_220,N_264);
and U389 (N_389,In_349,N_7);
xnor U390 (N_390,N_178,In_401);
nor U391 (N_391,N_280,N_311);
nand U392 (N_392,N_258,N_329);
nor U393 (N_393,N_223,N_31);
nor U394 (N_394,N_147,In_132);
or U395 (N_395,N_301,N_221);
nor U396 (N_396,N_289,N_292);
and U397 (N_397,N_268,N_246);
nor U398 (N_398,N_318,N_290);
or U399 (N_399,In_431,N_284);
and U400 (N_400,N_336,N_298);
xor U401 (N_401,In_481,N_324);
nand U402 (N_402,N_250,In_417);
and U403 (N_403,In_292,N_304);
nand U404 (N_404,In_487,In_71);
nand U405 (N_405,N_356,N_337);
and U406 (N_406,In_272,N_332);
xnor U407 (N_407,N_354,N_302);
or U408 (N_408,N_214,N_256);
and U409 (N_409,N_321,N_257);
nand U410 (N_410,N_71,N_353);
nor U411 (N_411,In_473,In_441);
nor U412 (N_412,N_347,N_185);
nor U413 (N_413,In_337,N_165);
or U414 (N_414,N_350,N_86);
xor U415 (N_415,N_352,N_209);
nand U416 (N_416,N_355,In_14);
or U417 (N_417,In_101,N_112);
and U418 (N_418,N_303,N_260);
nand U419 (N_419,N_309,In_406);
and U420 (N_420,N_384,N_366);
nand U421 (N_421,N_370,N_374);
or U422 (N_422,N_411,N_389);
nand U423 (N_423,N_403,N_367);
and U424 (N_424,N_372,N_405);
and U425 (N_425,N_415,N_105);
xnor U426 (N_426,N_391,N_386);
or U427 (N_427,N_161,N_381);
xor U428 (N_428,N_373,N_365);
nand U429 (N_429,N_300,N_385);
or U430 (N_430,N_360,N_375);
or U431 (N_431,N_408,N_419);
and U432 (N_432,N_306,N_418);
or U433 (N_433,N_414,N_12);
nand U434 (N_434,N_393,N_296);
or U435 (N_435,N_400,N_368);
nand U436 (N_436,N_341,N_390);
and U437 (N_437,N_392,N_377);
and U438 (N_438,N_404,In_114);
nor U439 (N_439,N_395,N_331);
or U440 (N_440,N_409,N_397);
and U441 (N_441,N_398,N_378);
nand U442 (N_442,N_330,N_212);
nor U443 (N_443,N_406,N_396);
nor U444 (N_444,N_399,N_361);
and U445 (N_445,N_339,N_412);
nor U446 (N_446,N_21,N_388);
or U447 (N_447,N_410,N_364);
nor U448 (N_448,In_136,N_383);
nor U449 (N_449,N_369,N_194);
or U450 (N_450,N_335,N_379);
and U451 (N_451,N_362,N_345);
nor U452 (N_452,N_382,N_376);
nor U453 (N_453,N_351,N_387);
xnor U454 (N_454,N_371,N_394);
nand U455 (N_455,N_416,N_402);
and U456 (N_456,N_316,N_407);
nand U457 (N_457,N_342,N_363);
nor U458 (N_458,N_417,N_413);
and U459 (N_459,N_380,N_401);
nor U460 (N_460,N_367,N_388);
and U461 (N_461,N_405,N_365);
xnor U462 (N_462,N_366,N_416);
xnor U463 (N_463,N_360,N_331);
xnor U464 (N_464,N_398,N_408);
xor U465 (N_465,N_300,N_383);
and U466 (N_466,N_306,N_402);
nand U467 (N_467,N_351,N_212);
nor U468 (N_468,N_416,N_414);
xor U469 (N_469,N_415,N_416);
nand U470 (N_470,N_351,N_371);
nand U471 (N_471,N_373,N_296);
or U472 (N_472,N_418,N_410);
and U473 (N_473,N_413,N_387);
nor U474 (N_474,N_381,N_405);
and U475 (N_475,N_335,N_380);
and U476 (N_476,N_408,N_105);
and U477 (N_477,N_330,N_402);
nor U478 (N_478,N_410,N_380);
or U479 (N_479,N_406,N_415);
and U480 (N_480,N_437,N_467);
nand U481 (N_481,N_453,N_474);
and U482 (N_482,N_423,N_478);
and U483 (N_483,N_473,N_421);
nand U484 (N_484,N_428,N_440);
or U485 (N_485,N_472,N_462);
nor U486 (N_486,N_438,N_426);
and U487 (N_487,N_422,N_420);
xnor U488 (N_488,N_441,N_458);
nor U489 (N_489,N_452,N_446);
nand U490 (N_490,N_457,N_470);
nor U491 (N_491,N_448,N_460);
nor U492 (N_492,N_475,N_479);
or U493 (N_493,N_471,N_434);
or U494 (N_494,N_469,N_459);
or U495 (N_495,N_477,N_465);
and U496 (N_496,N_464,N_439);
nor U497 (N_497,N_425,N_443);
nor U498 (N_498,N_430,N_432);
and U499 (N_499,N_435,N_447);
nor U500 (N_500,N_445,N_424);
nor U501 (N_501,N_455,N_444);
nand U502 (N_502,N_429,N_427);
and U503 (N_503,N_450,N_468);
or U504 (N_504,N_431,N_451);
nor U505 (N_505,N_466,N_442);
and U506 (N_506,N_454,N_461);
or U507 (N_507,N_433,N_476);
and U508 (N_508,N_456,N_436);
nor U509 (N_509,N_449,N_463);
and U510 (N_510,N_453,N_458);
or U511 (N_511,N_424,N_421);
and U512 (N_512,N_429,N_467);
or U513 (N_513,N_461,N_473);
xnor U514 (N_514,N_432,N_457);
nand U515 (N_515,N_455,N_445);
xnor U516 (N_516,N_420,N_478);
and U517 (N_517,N_434,N_456);
xnor U518 (N_518,N_452,N_450);
xor U519 (N_519,N_440,N_438);
nand U520 (N_520,N_423,N_458);
nand U521 (N_521,N_448,N_450);
nand U522 (N_522,N_447,N_448);
and U523 (N_523,N_438,N_429);
and U524 (N_524,N_461,N_443);
nand U525 (N_525,N_476,N_423);
nand U526 (N_526,N_460,N_437);
nand U527 (N_527,N_421,N_431);
or U528 (N_528,N_446,N_434);
nand U529 (N_529,N_461,N_463);
xnor U530 (N_530,N_420,N_432);
nor U531 (N_531,N_479,N_457);
and U532 (N_532,N_467,N_470);
and U533 (N_533,N_453,N_447);
xnor U534 (N_534,N_454,N_426);
or U535 (N_535,N_450,N_435);
or U536 (N_536,N_463,N_471);
nor U537 (N_537,N_477,N_430);
or U538 (N_538,N_437,N_431);
nand U539 (N_539,N_436,N_437);
nand U540 (N_540,N_533,N_488);
nor U541 (N_541,N_539,N_534);
or U542 (N_542,N_528,N_486);
and U543 (N_543,N_491,N_493);
xnor U544 (N_544,N_482,N_518);
nand U545 (N_545,N_496,N_520);
or U546 (N_546,N_489,N_490);
nand U547 (N_547,N_527,N_532);
nor U548 (N_548,N_500,N_494);
nand U549 (N_549,N_513,N_509);
or U550 (N_550,N_526,N_525);
xor U551 (N_551,N_516,N_481);
or U552 (N_552,N_511,N_524);
or U553 (N_553,N_523,N_514);
nor U554 (N_554,N_530,N_510);
and U555 (N_555,N_503,N_495);
nand U556 (N_556,N_507,N_499);
and U557 (N_557,N_504,N_531);
nand U558 (N_558,N_498,N_484);
or U559 (N_559,N_505,N_502);
and U560 (N_560,N_537,N_515);
and U561 (N_561,N_480,N_519);
nor U562 (N_562,N_521,N_538);
nand U563 (N_563,N_487,N_517);
and U564 (N_564,N_483,N_522);
and U565 (N_565,N_536,N_529);
and U566 (N_566,N_512,N_492);
and U567 (N_567,N_506,N_501);
nor U568 (N_568,N_535,N_508);
and U569 (N_569,N_497,N_485);
nor U570 (N_570,N_490,N_491);
and U571 (N_571,N_480,N_522);
xnor U572 (N_572,N_512,N_516);
nand U573 (N_573,N_517,N_482);
nand U574 (N_574,N_494,N_486);
or U575 (N_575,N_506,N_512);
nor U576 (N_576,N_535,N_525);
nor U577 (N_577,N_520,N_488);
nor U578 (N_578,N_532,N_530);
or U579 (N_579,N_493,N_507);
nor U580 (N_580,N_513,N_537);
xnor U581 (N_581,N_496,N_495);
xor U582 (N_582,N_528,N_512);
nor U583 (N_583,N_513,N_504);
or U584 (N_584,N_511,N_537);
and U585 (N_585,N_522,N_516);
nor U586 (N_586,N_517,N_488);
nand U587 (N_587,N_523,N_486);
or U588 (N_588,N_513,N_486);
or U589 (N_589,N_485,N_520);
and U590 (N_590,N_500,N_504);
and U591 (N_591,N_526,N_517);
and U592 (N_592,N_522,N_536);
and U593 (N_593,N_484,N_480);
and U594 (N_594,N_507,N_500);
nor U595 (N_595,N_495,N_506);
nor U596 (N_596,N_538,N_515);
and U597 (N_597,N_504,N_499);
nand U598 (N_598,N_505,N_531);
nand U599 (N_599,N_494,N_523);
or U600 (N_600,N_599,N_575);
nand U601 (N_601,N_572,N_557);
nand U602 (N_602,N_590,N_567);
and U603 (N_603,N_554,N_593);
or U604 (N_604,N_584,N_585);
or U605 (N_605,N_596,N_562);
nand U606 (N_606,N_589,N_551);
nor U607 (N_607,N_566,N_595);
nor U608 (N_608,N_540,N_597);
and U609 (N_609,N_573,N_578);
nor U610 (N_610,N_548,N_582);
nand U611 (N_611,N_580,N_586);
xor U612 (N_612,N_542,N_569);
and U613 (N_613,N_552,N_547);
xor U614 (N_614,N_574,N_594);
nor U615 (N_615,N_565,N_559);
and U616 (N_616,N_579,N_563);
and U617 (N_617,N_550,N_545);
or U618 (N_618,N_553,N_549);
nand U619 (N_619,N_598,N_546);
nor U620 (N_620,N_564,N_576);
nand U621 (N_621,N_568,N_581);
and U622 (N_622,N_587,N_561);
or U623 (N_623,N_591,N_583);
or U624 (N_624,N_555,N_588);
nand U625 (N_625,N_558,N_543);
and U626 (N_626,N_577,N_544);
nand U627 (N_627,N_560,N_592);
or U628 (N_628,N_556,N_571);
xor U629 (N_629,N_541,N_570);
nor U630 (N_630,N_554,N_561);
or U631 (N_631,N_573,N_544);
nor U632 (N_632,N_549,N_588);
and U633 (N_633,N_547,N_595);
nor U634 (N_634,N_582,N_578);
xnor U635 (N_635,N_599,N_582);
and U636 (N_636,N_544,N_587);
nand U637 (N_637,N_547,N_566);
nor U638 (N_638,N_576,N_570);
nor U639 (N_639,N_594,N_543);
nand U640 (N_640,N_554,N_548);
nor U641 (N_641,N_592,N_549);
xor U642 (N_642,N_584,N_595);
nor U643 (N_643,N_577,N_584);
or U644 (N_644,N_543,N_592);
and U645 (N_645,N_552,N_566);
or U646 (N_646,N_546,N_553);
or U647 (N_647,N_564,N_563);
and U648 (N_648,N_562,N_560);
and U649 (N_649,N_551,N_556);
xnor U650 (N_650,N_595,N_545);
or U651 (N_651,N_574,N_558);
xnor U652 (N_652,N_568,N_589);
and U653 (N_653,N_545,N_541);
or U654 (N_654,N_575,N_542);
or U655 (N_655,N_554,N_575);
xnor U656 (N_656,N_591,N_577);
or U657 (N_657,N_558,N_577);
xor U658 (N_658,N_564,N_588);
or U659 (N_659,N_596,N_569);
nor U660 (N_660,N_604,N_633);
and U661 (N_661,N_641,N_610);
nand U662 (N_662,N_608,N_656);
nand U663 (N_663,N_649,N_647);
or U664 (N_664,N_631,N_646);
nor U665 (N_665,N_648,N_636);
nand U666 (N_666,N_637,N_654);
nand U667 (N_667,N_635,N_639);
or U668 (N_668,N_629,N_616);
and U669 (N_669,N_634,N_612);
or U670 (N_670,N_628,N_644);
and U671 (N_671,N_622,N_624);
or U672 (N_672,N_602,N_645);
and U673 (N_673,N_605,N_643);
and U674 (N_674,N_611,N_625);
nor U675 (N_675,N_609,N_627);
or U676 (N_676,N_642,N_603);
xor U677 (N_677,N_621,N_600);
and U678 (N_678,N_601,N_653);
or U679 (N_679,N_626,N_623);
or U680 (N_680,N_659,N_607);
nor U681 (N_681,N_658,N_620);
nor U682 (N_682,N_651,N_650);
nor U683 (N_683,N_655,N_606);
nor U684 (N_684,N_630,N_618);
or U685 (N_685,N_615,N_640);
and U686 (N_686,N_617,N_613);
and U687 (N_687,N_614,N_638);
or U688 (N_688,N_632,N_652);
nor U689 (N_689,N_657,N_619);
nor U690 (N_690,N_649,N_637);
nor U691 (N_691,N_651,N_632);
or U692 (N_692,N_629,N_622);
or U693 (N_693,N_618,N_645);
nor U694 (N_694,N_644,N_631);
nor U695 (N_695,N_645,N_658);
xor U696 (N_696,N_658,N_657);
nand U697 (N_697,N_601,N_628);
nor U698 (N_698,N_604,N_647);
xor U699 (N_699,N_625,N_658);
or U700 (N_700,N_616,N_649);
and U701 (N_701,N_616,N_608);
and U702 (N_702,N_623,N_641);
nor U703 (N_703,N_642,N_637);
nor U704 (N_704,N_605,N_644);
nor U705 (N_705,N_636,N_600);
nand U706 (N_706,N_631,N_649);
and U707 (N_707,N_602,N_654);
xnor U708 (N_708,N_619,N_642);
xnor U709 (N_709,N_641,N_603);
nand U710 (N_710,N_647,N_642);
and U711 (N_711,N_654,N_615);
nor U712 (N_712,N_658,N_632);
or U713 (N_713,N_624,N_628);
or U714 (N_714,N_640,N_603);
nor U715 (N_715,N_613,N_622);
nor U716 (N_716,N_614,N_605);
or U717 (N_717,N_626,N_633);
and U718 (N_718,N_624,N_640);
nand U719 (N_719,N_648,N_605);
nor U720 (N_720,N_682,N_688);
or U721 (N_721,N_697,N_674);
and U722 (N_722,N_708,N_687);
and U723 (N_723,N_678,N_706);
and U724 (N_724,N_713,N_675);
nand U725 (N_725,N_719,N_690);
or U726 (N_726,N_665,N_661);
or U727 (N_727,N_693,N_673);
nor U728 (N_728,N_696,N_676);
or U729 (N_729,N_703,N_662);
and U730 (N_730,N_684,N_667);
or U731 (N_731,N_704,N_709);
nor U732 (N_732,N_717,N_712);
nand U733 (N_733,N_669,N_660);
nand U734 (N_734,N_670,N_715);
xor U735 (N_735,N_701,N_683);
or U736 (N_736,N_689,N_695);
and U737 (N_737,N_710,N_699);
or U738 (N_738,N_714,N_711);
or U739 (N_739,N_705,N_691);
nor U740 (N_740,N_707,N_698);
nand U741 (N_741,N_685,N_718);
nor U742 (N_742,N_671,N_679);
nand U743 (N_743,N_672,N_686);
and U744 (N_744,N_681,N_664);
xnor U745 (N_745,N_680,N_666);
and U746 (N_746,N_716,N_692);
xnor U747 (N_747,N_663,N_702);
xnor U748 (N_748,N_700,N_694);
xor U749 (N_749,N_677,N_668);
nand U750 (N_750,N_688,N_703);
and U751 (N_751,N_662,N_675);
and U752 (N_752,N_717,N_660);
nand U753 (N_753,N_688,N_690);
nand U754 (N_754,N_671,N_660);
nor U755 (N_755,N_694,N_697);
nand U756 (N_756,N_714,N_685);
nand U757 (N_757,N_681,N_695);
and U758 (N_758,N_680,N_676);
nand U759 (N_759,N_716,N_678);
xor U760 (N_760,N_701,N_689);
or U761 (N_761,N_666,N_710);
and U762 (N_762,N_690,N_697);
and U763 (N_763,N_703,N_692);
nand U764 (N_764,N_717,N_680);
xor U765 (N_765,N_702,N_686);
or U766 (N_766,N_695,N_705);
xor U767 (N_767,N_717,N_693);
or U768 (N_768,N_684,N_680);
and U769 (N_769,N_689,N_704);
nand U770 (N_770,N_684,N_677);
or U771 (N_771,N_705,N_699);
xnor U772 (N_772,N_704,N_672);
nor U773 (N_773,N_718,N_686);
and U774 (N_774,N_709,N_671);
or U775 (N_775,N_674,N_662);
and U776 (N_776,N_708,N_710);
xor U777 (N_777,N_674,N_666);
nand U778 (N_778,N_682,N_678);
or U779 (N_779,N_675,N_708);
and U780 (N_780,N_751,N_726);
nor U781 (N_781,N_743,N_760);
or U782 (N_782,N_754,N_775);
nor U783 (N_783,N_729,N_733);
nor U784 (N_784,N_742,N_770);
xor U785 (N_785,N_759,N_769);
and U786 (N_786,N_747,N_721);
nor U787 (N_787,N_737,N_736);
and U788 (N_788,N_725,N_741);
nor U789 (N_789,N_730,N_756);
nand U790 (N_790,N_757,N_763);
nor U791 (N_791,N_746,N_723);
or U792 (N_792,N_749,N_744);
and U793 (N_793,N_777,N_758);
xor U794 (N_794,N_728,N_735);
or U795 (N_795,N_774,N_779);
or U796 (N_796,N_731,N_764);
and U797 (N_797,N_734,N_761);
nor U798 (N_798,N_732,N_762);
or U799 (N_799,N_740,N_776);
and U800 (N_800,N_724,N_753);
nand U801 (N_801,N_778,N_727);
nand U802 (N_802,N_767,N_752);
nor U803 (N_803,N_738,N_722);
nand U804 (N_804,N_750,N_773);
xnor U805 (N_805,N_765,N_748);
and U806 (N_806,N_768,N_771);
or U807 (N_807,N_755,N_766);
and U808 (N_808,N_772,N_739);
nand U809 (N_809,N_720,N_745);
nand U810 (N_810,N_779,N_776);
or U811 (N_811,N_777,N_739);
nor U812 (N_812,N_757,N_727);
nor U813 (N_813,N_752,N_736);
nor U814 (N_814,N_752,N_762);
and U815 (N_815,N_762,N_730);
and U816 (N_816,N_733,N_766);
or U817 (N_817,N_752,N_741);
nand U818 (N_818,N_730,N_736);
nand U819 (N_819,N_753,N_754);
nand U820 (N_820,N_743,N_758);
or U821 (N_821,N_739,N_778);
nand U822 (N_822,N_778,N_746);
nor U823 (N_823,N_748,N_755);
and U824 (N_824,N_747,N_745);
or U825 (N_825,N_777,N_752);
xor U826 (N_826,N_775,N_728);
nor U827 (N_827,N_728,N_737);
nand U828 (N_828,N_769,N_729);
xor U829 (N_829,N_771,N_731);
xor U830 (N_830,N_777,N_723);
nor U831 (N_831,N_723,N_737);
and U832 (N_832,N_738,N_746);
or U833 (N_833,N_768,N_725);
and U834 (N_834,N_731,N_772);
or U835 (N_835,N_741,N_765);
or U836 (N_836,N_730,N_733);
or U837 (N_837,N_721,N_775);
nand U838 (N_838,N_733,N_748);
nand U839 (N_839,N_756,N_754);
nand U840 (N_840,N_784,N_794);
nand U841 (N_841,N_780,N_837);
and U842 (N_842,N_803,N_809);
or U843 (N_843,N_834,N_789);
nor U844 (N_844,N_827,N_822);
nand U845 (N_845,N_835,N_796);
nor U846 (N_846,N_788,N_820);
nor U847 (N_847,N_811,N_808);
nor U848 (N_848,N_830,N_813);
nand U849 (N_849,N_795,N_814);
xnor U850 (N_850,N_812,N_816);
and U851 (N_851,N_823,N_838);
nor U852 (N_852,N_785,N_802);
nor U853 (N_853,N_836,N_782);
or U854 (N_854,N_829,N_832);
and U855 (N_855,N_828,N_824);
and U856 (N_856,N_818,N_791);
nor U857 (N_857,N_801,N_787);
nand U858 (N_858,N_825,N_790);
xnor U859 (N_859,N_839,N_819);
nor U860 (N_860,N_833,N_781);
or U861 (N_861,N_817,N_815);
nand U862 (N_862,N_786,N_826);
and U863 (N_863,N_797,N_783);
nor U864 (N_864,N_807,N_798);
and U865 (N_865,N_799,N_805);
or U866 (N_866,N_810,N_821);
nand U867 (N_867,N_831,N_792);
nand U868 (N_868,N_806,N_804);
and U869 (N_869,N_793,N_800);
or U870 (N_870,N_791,N_836);
nor U871 (N_871,N_801,N_826);
xor U872 (N_872,N_814,N_790);
or U873 (N_873,N_806,N_794);
or U874 (N_874,N_824,N_825);
xnor U875 (N_875,N_816,N_800);
nand U876 (N_876,N_801,N_790);
and U877 (N_877,N_808,N_827);
or U878 (N_878,N_781,N_782);
or U879 (N_879,N_828,N_819);
or U880 (N_880,N_782,N_797);
nand U881 (N_881,N_816,N_785);
or U882 (N_882,N_802,N_822);
or U883 (N_883,N_826,N_781);
nand U884 (N_884,N_790,N_836);
nand U885 (N_885,N_793,N_839);
xor U886 (N_886,N_785,N_810);
or U887 (N_887,N_815,N_792);
xnor U888 (N_888,N_828,N_836);
and U889 (N_889,N_796,N_783);
or U890 (N_890,N_780,N_812);
nand U891 (N_891,N_832,N_795);
or U892 (N_892,N_784,N_789);
nor U893 (N_893,N_788,N_826);
or U894 (N_894,N_806,N_800);
and U895 (N_895,N_792,N_803);
nor U896 (N_896,N_804,N_834);
nand U897 (N_897,N_823,N_812);
and U898 (N_898,N_832,N_830);
xor U899 (N_899,N_789,N_781);
and U900 (N_900,N_887,N_853);
and U901 (N_901,N_865,N_891);
xor U902 (N_902,N_890,N_877);
and U903 (N_903,N_870,N_846);
or U904 (N_904,N_880,N_854);
and U905 (N_905,N_845,N_871);
nand U906 (N_906,N_861,N_883);
or U907 (N_907,N_878,N_898);
and U908 (N_908,N_889,N_888);
nand U909 (N_909,N_858,N_884);
or U910 (N_910,N_862,N_899);
xor U911 (N_911,N_850,N_859);
nor U912 (N_912,N_840,N_841);
xor U913 (N_913,N_860,N_874);
or U914 (N_914,N_842,N_897);
or U915 (N_915,N_896,N_864);
and U916 (N_916,N_856,N_867);
and U917 (N_917,N_847,N_882);
nor U918 (N_918,N_895,N_872);
and U919 (N_919,N_892,N_885);
and U920 (N_920,N_881,N_886);
nor U921 (N_921,N_876,N_868);
and U922 (N_922,N_852,N_855);
nand U923 (N_923,N_851,N_844);
and U924 (N_924,N_875,N_848);
nor U925 (N_925,N_873,N_849);
nand U926 (N_926,N_857,N_843);
or U927 (N_927,N_863,N_879);
nand U928 (N_928,N_893,N_866);
nand U929 (N_929,N_894,N_869);
and U930 (N_930,N_894,N_863);
nor U931 (N_931,N_859,N_876);
and U932 (N_932,N_897,N_890);
and U933 (N_933,N_862,N_871);
nor U934 (N_934,N_848,N_896);
nand U935 (N_935,N_854,N_886);
nand U936 (N_936,N_898,N_861);
and U937 (N_937,N_888,N_898);
or U938 (N_938,N_860,N_898);
nor U939 (N_939,N_885,N_875);
nor U940 (N_940,N_888,N_845);
and U941 (N_941,N_888,N_893);
nand U942 (N_942,N_896,N_884);
and U943 (N_943,N_864,N_880);
nor U944 (N_944,N_857,N_883);
nor U945 (N_945,N_862,N_892);
nand U946 (N_946,N_872,N_870);
nand U947 (N_947,N_879,N_872);
nor U948 (N_948,N_889,N_856);
or U949 (N_949,N_892,N_858);
nand U950 (N_950,N_862,N_870);
nor U951 (N_951,N_897,N_872);
nand U952 (N_952,N_843,N_849);
and U953 (N_953,N_894,N_866);
nor U954 (N_954,N_886,N_899);
nand U955 (N_955,N_881,N_879);
nor U956 (N_956,N_878,N_895);
or U957 (N_957,N_861,N_855);
nand U958 (N_958,N_893,N_865);
and U959 (N_959,N_846,N_871);
or U960 (N_960,N_945,N_957);
nand U961 (N_961,N_906,N_912);
nand U962 (N_962,N_910,N_950);
nand U963 (N_963,N_915,N_952);
and U964 (N_964,N_949,N_937);
nor U965 (N_965,N_956,N_935);
xnor U966 (N_966,N_908,N_904);
or U967 (N_967,N_930,N_932);
nand U968 (N_968,N_921,N_928);
and U969 (N_969,N_925,N_936);
nor U970 (N_970,N_942,N_914);
and U971 (N_971,N_903,N_923);
xnor U972 (N_972,N_948,N_920);
nor U973 (N_973,N_905,N_927);
nor U974 (N_974,N_944,N_900);
and U975 (N_975,N_924,N_913);
nand U976 (N_976,N_901,N_933);
or U977 (N_977,N_931,N_958);
or U978 (N_978,N_929,N_919);
and U979 (N_979,N_947,N_941);
xnor U980 (N_980,N_917,N_938);
nand U981 (N_981,N_922,N_954);
or U982 (N_982,N_959,N_951);
xnor U983 (N_983,N_946,N_909);
and U984 (N_984,N_907,N_934);
and U985 (N_985,N_911,N_918);
nand U986 (N_986,N_939,N_902);
and U987 (N_987,N_943,N_916);
nor U988 (N_988,N_953,N_940);
or U989 (N_989,N_926,N_955);
nor U990 (N_990,N_918,N_931);
nor U991 (N_991,N_924,N_933);
nor U992 (N_992,N_939,N_948);
and U993 (N_993,N_908,N_939);
or U994 (N_994,N_902,N_920);
or U995 (N_995,N_910,N_941);
nor U996 (N_996,N_924,N_912);
or U997 (N_997,N_958,N_929);
and U998 (N_998,N_952,N_941);
nor U999 (N_999,N_937,N_952);
nand U1000 (N_1000,N_947,N_913);
nor U1001 (N_1001,N_904,N_958);
and U1002 (N_1002,N_944,N_921);
or U1003 (N_1003,N_922,N_924);
xnor U1004 (N_1004,N_956,N_947);
xor U1005 (N_1005,N_926,N_911);
nor U1006 (N_1006,N_949,N_938);
or U1007 (N_1007,N_942,N_911);
or U1008 (N_1008,N_925,N_902);
nor U1009 (N_1009,N_904,N_921);
and U1010 (N_1010,N_947,N_911);
or U1011 (N_1011,N_954,N_911);
nand U1012 (N_1012,N_915,N_902);
xnor U1013 (N_1013,N_915,N_935);
nand U1014 (N_1014,N_931,N_950);
xnor U1015 (N_1015,N_932,N_917);
or U1016 (N_1016,N_958,N_909);
nor U1017 (N_1017,N_906,N_910);
xnor U1018 (N_1018,N_908,N_900);
and U1019 (N_1019,N_950,N_955);
nor U1020 (N_1020,N_987,N_993);
or U1021 (N_1021,N_1004,N_998);
xor U1022 (N_1022,N_986,N_1003);
nand U1023 (N_1023,N_964,N_1013);
nand U1024 (N_1024,N_960,N_965);
and U1025 (N_1025,N_999,N_994);
and U1026 (N_1026,N_989,N_979);
nor U1027 (N_1027,N_981,N_1016);
nand U1028 (N_1028,N_996,N_1010);
and U1029 (N_1029,N_1018,N_1019);
nor U1030 (N_1030,N_1001,N_1011);
nor U1031 (N_1031,N_980,N_966);
nand U1032 (N_1032,N_971,N_969);
nor U1033 (N_1033,N_1017,N_972);
nor U1034 (N_1034,N_975,N_1005);
xor U1035 (N_1035,N_1008,N_1012);
nand U1036 (N_1036,N_973,N_992);
and U1037 (N_1037,N_961,N_1002);
nand U1038 (N_1038,N_1000,N_982);
or U1039 (N_1039,N_963,N_1009);
xnor U1040 (N_1040,N_976,N_967);
and U1041 (N_1041,N_995,N_1007);
nor U1042 (N_1042,N_978,N_1015);
and U1043 (N_1043,N_977,N_997);
nor U1044 (N_1044,N_962,N_990);
nand U1045 (N_1045,N_974,N_970);
nor U1046 (N_1046,N_984,N_1006);
nor U1047 (N_1047,N_968,N_983);
and U1048 (N_1048,N_991,N_1014);
nand U1049 (N_1049,N_988,N_985);
or U1050 (N_1050,N_1009,N_969);
or U1051 (N_1051,N_985,N_1006);
and U1052 (N_1052,N_965,N_1004);
nor U1053 (N_1053,N_995,N_963);
nand U1054 (N_1054,N_978,N_961);
or U1055 (N_1055,N_1015,N_1012);
nand U1056 (N_1056,N_986,N_988);
and U1057 (N_1057,N_979,N_1015);
or U1058 (N_1058,N_977,N_981);
and U1059 (N_1059,N_982,N_969);
xor U1060 (N_1060,N_963,N_970);
nand U1061 (N_1061,N_1003,N_990);
xor U1062 (N_1062,N_962,N_993);
nand U1063 (N_1063,N_985,N_1014);
or U1064 (N_1064,N_1005,N_992);
or U1065 (N_1065,N_970,N_1003);
or U1066 (N_1066,N_964,N_962);
nand U1067 (N_1067,N_1019,N_1013);
xnor U1068 (N_1068,N_970,N_969);
or U1069 (N_1069,N_982,N_981);
nand U1070 (N_1070,N_987,N_1008);
nor U1071 (N_1071,N_983,N_990);
and U1072 (N_1072,N_962,N_1008);
nor U1073 (N_1073,N_981,N_1017);
nor U1074 (N_1074,N_974,N_971);
or U1075 (N_1075,N_1014,N_986);
nor U1076 (N_1076,N_975,N_987);
nor U1077 (N_1077,N_1006,N_994);
and U1078 (N_1078,N_1018,N_963);
nor U1079 (N_1079,N_960,N_984);
nand U1080 (N_1080,N_1020,N_1046);
xnor U1081 (N_1081,N_1049,N_1061);
nand U1082 (N_1082,N_1034,N_1031);
and U1083 (N_1083,N_1036,N_1079);
and U1084 (N_1084,N_1040,N_1070);
nand U1085 (N_1085,N_1072,N_1066);
nor U1086 (N_1086,N_1022,N_1058);
and U1087 (N_1087,N_1052,N_1065);
and U1088 (N_1088,N_1045,N_1041);
nand U1089 (N_1089,N_1051,N_1078);
nor U1090 (N_1090,N_1067,N_1060);
and U1091 (N_1091,N_1024,N_1033);
or U1092 (N_1092,N_1025,N_1038);
xnor U1093 (N_1093,N_1043,N_1048);
xor U1094 (N_1094,N_1063,N_1068);
nor U1095 (N_1095,N_1028,N_1064);
or U1096 (N_1096,N_1057,N_1059);
and U1097 (N_1097,N_1056,N_1074);
and U1098 (N_1098,N_1071,N_1021);
and U1099 (N_1099,N_1029,N_1054);
and U1100 (N_1100,N_1023,N_1073);
nand U1101 (N_1101,N_1047,N_1039);
and U1102 (N_1102,N_1050,N_1076);
nand U1103 (N_1103,N_1055,N_1075);
or U1104 (N_1104,N_1032,N_1069);
nand U1105 (N_1105,N_1044,N_1030);
and U1106 (N_1106,N_1027,N_1077);
nand U1107 (N_1107,N_1026,N_1037);
and U1108 (N_1108,N_1062,N_1035);
or U1109 (N_1109,N_1053,N_1042);
nand U1110 (N_1110,N_1025,N_1047);
nand U1111 (N_1111,N_1061,N_1043);
and U1112 (N_1112,N_1052,N_1044);
nand U1113 (N_1113,N_1078,N_1076);
or U1114 (N_1114,N_1041,N_1068);
or U1115 (N_1115,N_1046,N_1028);
and U1116 (N_1116,N_1073,N_1051);
and U1117 (N_1117,N_1072,N_1073);
nor U1118 (N_1118,N_1055,N_1058);
or U1119 (N_1119,N_1053,N_1071);
or U1120 (N_1120,N_1067,N_1057);
and U1121 (N_1121,N_1032,N_1024);
or U1122 (N_1122,N_1029,N_1033);
xor U1123 (N_1123,N_1025,N_1064);
and U1124 (N_1124,N_1029,N_1028);
or U1125 (N_1125,N_1048,N_1036);
nor U1126 (N_1126,N_1063,N_1034);
nand U1127 (N_1127,N_1058,N_1064);
xor U1128 (N_1128,N_1054,N_1026);
nand U1129 (N_1129,N_1065,N_1022);
nor U1130 (N_1130,N_1020,N_1054);
nand U1131 (N_1131,N_1022,N_1050);
nor U1132 (N_1132,N_1057,N_1032);
or U1133 (N_1133,N_1047,N_1030);
or U1134 (N_1134,N_1038,N_1057);
nor U1135 (N_1135,N_1035,N_1032);
xor U1136 (N_1136,N_1061,N_1034);
and U1137 (N_1137,N_1029,N_1062);
nand U1138 (N_1138,N_1076,N_1028);
nand U1139 (N_1139,N_1079,N_1033);
nor U1140 (N_1140,N_1090,N_1111);
and U1141 (N_1141,N_1134,N_1130);
or U1142 (N_1142,N_1119,N_1112);
nand U1143 (N_1143,N_1120,N_1089);
or U1144 (N_1144,N_1087,N_1081);
nor U1145 (N_1145,N_1093,N_1095);
nand U1146 (N_1146,N_1138,N_1137);
nand U1147 (N_1147,N_1126,N_1125);
or U1148 (N_1148,N_1092,N_1105);
or U1149 (N_1149,N_1101,N_1085);
nand U1150 (N_1150,N_1104,N_1121);
nor U1151 (N_1151,N_1096,N_1098);
xnor U1152 (N_1152,N_1100,N_1127);
and U1153 (N_1153,N_1102,N_1103);
xnor U1154 (N_1154,N_1132,N_1131);
or U1155 (N_1155,N_1128,N_1109);
nor U1156 (N_1156,N_1115,N_1116);
nand U1157 (N_1157,N_1082,N_1124);
and U1158 (N_1158,N_1135,N_1091);
nand U1159 (N_1159,N_1080,N_1108);
and U1160 (N_1160,N_1099,N_1133);
nor U1161 (N_1161,N_1123,N_1113);
nor U1162 (N_1162,N_1118,N_1114);
xnor U1163 (N_1163,N_1094,N_1110);
xor U1164 (N_1164,N_1122,N_1107);
nand U1165 (N_1165,N_1088,N_1097);
and U1166 (N_1166,N_1129,N_1106);
or U1167 (N_1167,N_1136,N_1086);
nor U1168 (N_1168,N_1083,N_1139);
or U1169 (N_1169,N_1117,N_1084);
nand U1170 (N_1170,N_1096,N_1106);
nand U1171 (N_1171,N_1115,N_1127);
nand U1172 (N_1172,N_1081,N_1096);
xor U1173 (N_1173,N_1121,N_1081);
nand U1174 (N_1174,N_1093,N_1092);
xnor U1175 (N_1175,N_1114,N_1082);
or U1176 (N_1176,N_1101,N_1096);
and U1177 (N_1177,N_1131,N_1089);
nor U1178 (N_1178,N_1124,N_1101);
or U1179 (N_1179,N_1100,N_1133);
nand U1180 (N_1180,N_1128,N_1134);
nand U1181 (N_1181,N_1126,N_1113);
and U1182 (N_1182,N_1128,N_1102);
nor U1183 (N_1183,N_1116,N_1124);
xor U1184 (N_1184,N_1138,N_1107);
or U1185 (N_1185,N_1114,N_1119);
nor U1186 (N_1186,N_1128,N_1081);
nand U1187 (N_1187,N_1120,N_1100);
nor U1188 (N_1188,N_1130,N_1125);
nand U1189 (N_1189,N_1087,N_1100);
nor U1190 (N_1190,N_1122,N_1098);
nand U1191 (N_1191,N_1111,N_1138);
nor U1192 (N_1192,N_1098,N_1131);
nor U1193 (N_1193,N_1081,N_1089);
and U1194 (N_1194,N_1113,N_1081);
or U1195 (N_1195,N_1124,N_1100);
nand U1196 (N_1196,N_1127,N_1087);
nor U1197 (N_1197,N_1088,N_1132);
and U1198 (N_1198,N_1109,N_1132);
xnor U1199 (N_1199,N_1092,N_1085);
or U1200 (N_1200,N_1143,N_1170);
nand U1201 (N_1201,N_1171,N_1175);
or U1202 (N_1202,N_1162,N_1147);
and U1203 (N_1203,N_1144,N_1195);
nor U1204 (N_1204,N_1156,N_1165);
or U1205 (N_1205,N_1148,N_1153);
or U1206 (N_1206,N_1187,N_1159);
xor U1207 (N_1207,N_1197,N_1188);
nor U1208 (N_1208,N_1146,N_1178);
xor U1209 (N_1209,N_1177,N_1141);
and U1210 (N_1210,N_1183,N_1179);
and U1211 (N_1211,N_1164,N_1180);
or U1212 (N_1212,N_1182,N_1189);
or U1213 (N_1213,N_1199,N_1152);
nand U1214 (N_1214,N_1168,N_1184);
or U1215 (N_1215,N_1169,N_1145);
xnor U1216 (N_1216,N_1173,N_1190);
xnor U1217 (N_1217,N_1174,N_1185);
nand U1218 (N_1218,N_1196,N_1176);
and U1219 (N_1219,N_1154,N_1150);
nand U1220 (N_1220,N_1140,N_1157);
nor U1221 (N_1221,N_1161,N_1163);
xnor U1222 (N_1222,N_1186,N_1191);
and U1223 (N_1223,N_1160,N_1193);
and U1224 (N_1224,N_1149,N_1194);
and U1225 (N_1225,N_1192,N_1158);
xnor U1226 (N_1226,N_1155,N_1181);
and U1227 (N_1227,N_1172,N_1151);
and U1228 (N_1228,N_1167,N_1198);
nand U1229 (N_1229,N_1142,N_1166);
or U1230 (N_1230,N_1190,N_1144);
or U1231 (N_1231,N_1198,N_1194);
and U1232 (N_1232,N_1184,N_1182);
and U1233 (N_1233,N_1140,N_1176);
nor U1234 (N_1234,N_1153,N_1164);
and U1235 (N_1235,N_1182,N_1166);
or U1236 (N_1236,N_1146,N_1151);
or U1237 (N_1237,N_1183,N_1176);
or U1238 (N_1238,N_1165,N_1146);
and U1239 (N_1239,N_1183,N_1190);
nand U1240 (N_1240,N_1194,N_1190);
or U1241 (N_1241,N_1145,N_1151);
nand U1242 (N_1242,N_1198,N_1147);
nor U1243 (N_1243,N_1174,N_1150);
nand U1244 (N_1244,N_1163,N_1185);
and U1245 (N_1245,N_1190,N_1174);
and U1246 (N_1246,N_1188,N_1198);
or U1247 (N_1247,N_1192,N_1145);
nand U1248 (N_1248,N_1145,N_1155);
nand U1249 (N_1249,N_1145,N_1189);
and U1250 (N_1250,N_1194,N_1172);
or U1251 (N_1251,N_1150,N_1189);
nor U1252 (N_1252,N_1155,N_1189);
or U1253 (N_1253,N_1184,N_1193);
nand U1254 (N_1254,N_1177,N_1167);
nor U1255 (N_1255,N_1199,N_1196);
nand U1256 (N_1256,N_1161,N_1177);
and U1257 (N_1257,N_1183,N_1164);
or U1258 (N_1258,N_1145,N_1171);
nor U1259 (N_1259,N_1141,N_1196);
and U1260 (N_1260,N_1219,N_1202);
or U1261 (N_1261,N_1213,N_1224);
xor U1262 (N_1262,N_1238,N_1248);
or U1263 (N_1263,N_1220,N_1246);
nand U1264 (N_1264,N_1235,N_1229);
nand U1265 (N_1265,N_1234,N_1232);
nand U1266 (N_1266,N_1247,N_1209);
nor U1267 (N_1267,N_1255,N_1256);
and U1268 (N_1268,N_1259,N_1236);
or U1269 (N_1269,N_1222,N_1200);
nor U1270 (N_1270,N_1205,N_1206);
or U1271 (N_1271,N_1204,N_1228);
nor U1272 (N_1272,N_1225,N_1245);
and U1273 (N_1273,N_1242,N_1218);
or U1274 (N_1274,N_1231,N_1207);
nor U1275 (N_1275,N_1244,N_1210);
and U1276 (N_1276,N_1211,N_1214);
and U1277 (N_1277,N_1215,N_1203);
nor U1278 (N_1278,N_1254,N_1257);
xor U1279 (N_1279,N_1226,N_1233);
nor U1280 (N_1280,N_1221,N_1237);
or U1281 (N_1281,N_1253,N_1208);
nand U1282 (N_1282,N_1212,N_1239);
nand U1283 (N_1283,N_1230,N_1227);
or U1284 (N_1284,N_1249,N_1241);
nor U1285 (N_1285,N_1223,N_1201);
nor U1286 (N_1286,N_1250,N_1258);
and U1287 (N_1287,N_1217,N_1216);
nand U1288 (N_1288,N_1240,N_1251);
or U1289 (N_1289,N_1243,N_1252);
nor U1290 (N_1290,N_1219,N_1207);
nand U1291 (N_1291,N_1217,N_1245);
nor U1292 (N_1292,N_1211,N_1241);
or U1293 (N_1293,N_1251,N_1234);
nor U1294 (N_1294,N_1233,N_1200);
nand U1295 (N_1295,N_1243,N_1240);
and U1296 (N_1296,N_1226,N_1236);
nand U1297 (N_1297,N_1236,N_1258);
and U1298 (N_1298,N_1205,N_1251);
nor U1299 (N_1299,N_1216,N_1238);
or U1300 (N_1300,N_1235,N_1243);
nor U1301 (N_1301,N_1216,N_1245);
xor U1302 (N_1302,N_1231,N_1214);
nand U1303 (N_1303,N_1253,N_1243);
and U1304 (N_1304,N_1251,N_1256);
and U1305 (N_1305,N_1244,N_1248);
or U1306 (N_1306,N_1228,N_1211);
or U1307 (N_1307,N_1254,N_1219);
and U1308 (N_1308,N_1250,N_1216);
nor U1309 (N_1309,N_1227,N_1249);
nand U1310 (N_1310,N_1208,N_1218);
nand U1311 (N_1311,N_1209,N_1213);
nand U1312 (N_1312,N_1214,N_1222);
nand U1313 (N_1313,N_1240,N_1208);
or U1314 (N_1314,N_1252,N_1222);
or U1315 (N_1315,N_1258,N_1226);
xnor U1316 (N_1316,N_1252,N_1202);
xor U1317 (N_1317,N_1258,N_1208);
and U1318 (N_1318,N_1206,N_1220);
or U1319 (N_1319,N_1250,N_1224);
or U1320 (N_1320,N_1301,N_1313);
or U1321 (N_1321,N_1261,N_1291);
or U1322 (N_1322,N_1309,N_1275);
and U1323 (N_1323,N_1318,N_1312);
xnor U1324 (N_1324,N_1289,N_1311);
nand U1325 (N_1325,N_1284,N_1267);
nor U1326 (N_1326,N_1294,N_1281);
or U1327 (N_1327,N_1306,N_1317);
nor U1328 (N_1328,N_1272,N_1273);
nand U1329 (N_1329,N_1279,N_1304);
nor U1330 (N_1330,N_1305,N_1292);
and U1331 (N_1331,N_1303,N_1315);
and U1332 (N_1332,N_1287,N_1307);
nor U1333 (N_1333,N_1276,N_1268);
xor U1334 (N_1334,N_1269,N_1296);
nor U1335 (N_1335,N_1299,N_1263);
nand U1336 (N_1336,N_1286,N_1297);
xnor U1337 (N_1337,N_1295,N_1271);
or U1338 (N_1338,N_1280,N_1302);
nand U1339 (N_1339,N_1282,N_1319);
or U1340 (N_1340,N_1277,N_1274);
and U1341 (N_1341,N_1310,N_1308);
and U1342 (N_1342,N_1300,N_1265);
nand U1343 (N_1343,N_1262,N_1293);
or U1344 (N_1344,N_1283,N_1266);
nor U1345 (N_1345,N_1314,N_1298);
nand U1346 (N_1346,N_1290,N_1260);
nor U1347 (N_1347,N_1270,N_1264);
xnor U1348 (N_1348,N_1316,N_1285);
nand U1349 (N_1349,N_1278,N_1288);
and U1350 (N_1350,N_1290,N_1275);
or U1351 (N_1351,N_1311,N_1300);
or U1352 (N_1352,N_1292,N_1293);
and U1353 (N_1353,N_1261,N_1273);
or U1354 (N_1354,N_1267,N_1318);
nand U1355 (N_1355,N_1313,N_1305);
and U1356 (N_1356,N_1294,N_1296);
or U1357 (N_1357,N_1291,N_1290);
and U1358 (N_1358,N_1291,N_1287);
nand U1359 (N_1359,N_1266,N_1291);
nand U1360 (N_1360,N_1316,N_1301);
nor U1361 (N_1361,N_1284,N_1270);
or U1362 (N_1362,N_1314,N_1286);
nand U1363 (N_1363,N_1283,N_1280);
and U1364 (N_1364,N_1262,N_1299);
nor U1365 (N_1365,N_1276,N_1311);
nor U1366 (N_1366,N_1282,N_1301);
and U1367 (N_1367,N_1283,N_1303);
and U1368 (N_1368,N_1287,N_1313);
nand U1369 (N_1369,N_1300,N_1318);
and U1370 (N_1370,N_1275,N_1266);
nand U1371 (N_1371,N_1297,N_1318);
xnor U1372 (N_1372,N_1283,N_1285);
nand U1373 (N_1373,N_1314,N_1266);
nand U1374 (N_1374,N_1298,N_1302);
nand U1375 (N_1375,N_1260,N_1301);
and U1376 (N_1376,N_1316,N_1286);
nand U1377 (N_1377,N_1287,N_1282);
or U1378 (N_1378,N_1299,N_1300);
nor U1379 (N_1379,N_1298,N_1285);
nand U1380 (N_1380,N_1343,N_1328);
xor U1381 (N_1381,N_1353,N_1349);
and U1382 (N_1382,N_1355,N_1368);
and U1383 (N_1383,N_1320,N_1377);
nor U1384 (N_1384,N_1366,N_1350);
and U1385 (N_1385,N_1346,N_1324);
or U1386 (N_1386,N_1344,N_1326);
or U1387 (N_1387,N_1338,N_1364);
nor U1388 (N_1388,N_1376,N_1374);
or U1389 (N_1389,N_1321,N_1331);
nor U1390 (N_1390,N_1340,N_1323);
and U1391 (N_1391,N_1357,N_1359);
or U1392 (N_1392,N_1362,N_1334);
and U1393 (N_1393,N_1337,N_1332);
or U1394 (N_1394,N_1341,N_1371);
nor U1395 (N_1395,N_1360,N_1379);
or U1396 (N_1396,N_1347,N_1369);
nand U1397 (N_1397,N_1342,N_1330);
or U1398 (N_1398,N_1329,N_1322);
and U1399 (N_1399,N_1339,N_1367);
nand U1400 (N_1400,N_1361,N_1335);
or U1401 (N_1401,N_1354,N_1351);
or U1402 (N_1402,N_1363,N_1345);
nand U1403 (N_1403,N_1378,N_1348);
and U1404 (N_1404,N_1336,N_1365);
or U1405 (N_1405,N_1373,N_1370);
and U1406 (N_1406,N_1358,N_1333);
and U1407 (N_1407,N_1375,N_1372);
and U1408 (N_1408,N_1325,N_1352);
and U1409 (N_1409,N_1327,N_1356);
nand U1410 (N_1410,N_1339,N_1359);
nor U1411 (N_1411,N_1338,N_1355);
and U1412 (N_1412,N_1370,N_1375);
nand U1413 (N_1413,N_1351,N_1357);
nand U1414 (N_1414,N_1334,N_1340);
and U1415 (N_1415,N_1363,N_1352);
or U1416 (N_1416,N_1350,N_1353);
or U1417 (N_1417,N_1324,N_1378);
or U1418 (N_1418,N_1320,N_1328);
or U1419 (N_1419,N_1358,N_1327);
nor U1420 (N_1420,N_1341,N_1340);
nor U1421 (N_1421,N_1324,N_1367);
or U1422 (N_1422,N_1326,N_1334);
nand U1423 (N_1423,N_1350,N_1364);
and U1424 (N_1424,N_1360,N_1370);
or U1425 (N_1425,N_1343,N_1322);
nand U1426 (N_1426,N_1364,N_1348);
nor U1427 (N_1427,N_1334,N_1342);
nor U1428 (N_1428,N_1329,N_1331);
nand U1429 (N_1429,N_1355,N_1323);
or U1430 (N_1430,N_1368,N_1341);
or U1431 (N_1431,N_1349,N_1345);
and U1432 (N_1432,N_1324,N_1377);
or U1433 (N_1433,N_1344,N_1346);
nand U1434 (N_1434,N_1362,N_1344);
or U1435 (N_1435,N_1347,N_1322);
nor U1436 (N_1436,N_1368,N_1379);
nor U1437 (N_1437,N_1330,N_1359);
nand U1438 (N_1438,N_1336,N_1333);
nand U1439 (N_1439,N_1321,N_1341);
and U1440 (N_1440,N_1399,N_1393);
or U1441 (N_1441,N_1405,N_1434);
and U1442 (N_1442,N_1420,N_1414);
nor U1443 (N_1443,N_1408,N_1438);
nand U1444 (N_1444,N_1400,N_1384);
and U1445 (N_1445,N_1429,N_1423);
xnor U1446 (N_1446,N_1430,N_1404);
and U1447 (N_1447,N_1412,N_1424);
and U1448 (N_1448,N_1388,N_1390);
or U1449 (N_1449,N_1397,N_1401);
nand U1450 (N_1450,N_1421,N_1407);
xor U1451 (N_1451,N_1411,N_1383);
nand U1452 (N_1452,N_1416,N_1437);
and U1453 (N_1453,N_1406,N_1431);
nor U1454 (N_1454,N_1381,N_1417);
or U1455 (N_1455,N_1385,N_1433);
or U1456 (N_1456,N_1382,N_1392);
nor U1457 (N_1457,N_1428,N_1427);
and U1458 (N_1458,N_1389,N_1387);
nand U1459 (N_1459,N_1413,N_1439);
or U1460 (N_1460,N_1432,N_1419);
or U1461 (N_1461,N_1422,N_1394);
or U1462 (N_1462,N_1409,N_1386);
nor U1463 (N_1463,N_1396,N_1395);
or U1464 (N_1464,N_1398,N_1426);
and U1465 (N_1465,N_1435,N_1436);
nand U1466 (N_1466,N_1425,N_1415);
nor U1467 (N_1467,N_1402,N_1418);
and U1468 (N_1468,N_1391,N_1410);
or U1469 (N_1469,N_1403,N_1380);
xnor U1470 (N_1470,N_1423,N_1417);
and U1471 (N_1471,N_1433,N_1401);
or U1472 (N_1472,N_1407,N_1399);
and U1473 (N_1473,N_1412,N_1405);
xnor U1474 (N_1474,N_1383,N_1418);
and U1475 (N_1475,N_1418,N_1412);
nor U1476 (N_1476,N_1382,N_1426);
nor U1477 (N_1477,N_1397,N_1425);
or U1478 (N_1478,N_1393,N_1381);
nor U1479 (N_1479,N_1396,N_1438);
or U1480 (N_1480,N_1435,N_1391);
xor U1481 (N_1481,N_1409,N_1408);
and U1482 (N_1482,N_1387,N_1423);
or U1483 (N_1483,N_1425,N_1406);
nor U1484 (N_1484,N_1403,N_1438);
nand U1485 (N_1485,N_1392,N_1410);
xor U1486 (N_1486,N_1397,N_1423);
xnor U1487 (N_1487,N_1381,N_1426);
nand U1488 (N_1488,N_1433,N_1398);
or U1489 (N_1489,N_1426,N_1387);
and U1490 (N_1490,N_1420,N_1403);
nand U1491 (N_1491,N_1439,N_1389);
xnor U1492 (N_1492,N_1383,N_1386);
nor U1493 (N_1493,N_1428,N_1435);
nor U1494 (N_1494,N_1434,N_1435);
nand U1495 (N_1495,N_1383,N_1391);
and U1496 (N_1496,N_1389,N_1436);
and U1497 (N_1497,N_1432,N_1421);
or U1498 (N_1498,N_1434,N_1404);
nor U1499 (N_1499,N_1427,N_1406);
nor U1500 (N_1500,N_1479,N_1488);
nand U1501 (N_1501,N_1451,N_1462);
or U1502 (N_1502,N_1470,N_1481);
and U1503 (N_1503,N_1473,N_1440);
or U1504 (N_1504,N_1497,N_1461);
and U1505 (N_1505,N_1472,N_1452);
or U1506 (N_1506,N_1478,N_1475);
nor U1507 (N_1507,N_1468,N_1476);
or U1508 (N_1508,N_1477,N_1493);
and U1509 (N_1509,N_1482,N_1474);
and U1510 (N_1510,N_1471,N_1459);
and U1511 (N_1511,N_1490,N_1489);
nor U1512 (N_1512,N_1458,N_1443);
nand U1513 (N_1513,N_1456,N_1445);
and U1514 (N_1514,N_1447,N_1449);
nand U1515 (N_1515,N_1495,N_1467);
or U1516 (N_1516,N_1480,N_1499);
and U1517 (N_1517,N_1454,N_1448);
nand U1518 (N_1518,N_1444,N_1453);
nand U1519 (N_1519,N_1487,N_1483);
and U1520 (N_1520,N_1486,N_1441);
nand U1521 (N_1521,N_1496,N_1469);
or U1522 (N_1522,N_1463,N_1484);
nand U1523 (N_1523,N_1498,N_1464);
nor U1524 (N_1524,N_1465,N_1455);
xor U1525 (N_1525,N_1442,N_1491);
or U1526 (N_1526,N_1457,N_1460);
xor U1527 (N_1527,N_1450,N_1485);
or U1528 (N_1528,N_1492,N_1466);
or U1529 (N_1529,N_1446,N_1494);
nand U1530 (N_1530,N_1489,N_1470);
or U1531 (N_1531,N_1481,N_1477);
nor U1532 (N_1532,N_1478,N_1464);
xor U1533 (N_1533,N_1496,N_1476);
nand U1534 (N_1534,N_1456,N_1459);
or U1535 (N_1535,N_1455,N_1497);
nand U1536 (N_1536,N_1486,N_1488);
xnor U1537 (N_1537,N_1448,N_1474);
nand U1538 (N_1538,N_1451,N_1469);
or U1539 (N_1539,N_1443,N_1483);
or U1540 (N_1540,N_1460,N_1491);
or U1541 (N_1541,N_1452,N_1454);
nand U1542 (N_1542,N_1465,N_1488);
nand U1543 (N_1543,N_1482,N_1484);
nand U1544 (N_1544,N_1486,N_1461);
nand U1545 (N_1545,N_1477,N_1497);
xnor U1546 (N_1546,N_1491,N_1472);
nor U1547 (N_1547,N_1465,N_1444);
nand U1548 (N_1548,N_1478,N_1498);
xnor U1549 (N_1549,N_1473,N_1444);
nand U1550 (N_1550,N_1446,N_1490);
nand U1551 (N_1551,N_1451,N_1496);
nand U1552 (N_1552,N_1471,N_1492);
and U1553 (N_1553,N_1495,N_1487);
and U1554 (N_1554,N_1454,N_1476);
or U1555 (N_1555,N_1466,N_1495);
nor U1556 (N_1556,N_1495,N_1455);
and U1557 (N_1557,N_1449,N_1463);
or U1558 (N_1558,N_1494,N_1484);
nand U1559 (N_1559,N_1498,N_1451);
nor U1560 (N_1560,N_1541,N_1514);
or U1561 (N_1561,N_1557,N_1554);
and U1562 (N_1562,N_1518,N_1517);
xnor U1563 (N_1563,N_1524,N_1539);
nand U1564 (N_1564,N_1513,N_1538);
and U1565 (N_1565,N_1553,N_1529);
or U1566 (N_1566,N_1502,N_1525);
xor U1567 (N_1567,N_1545,N_1531);
nand U1568 (N_1568,N_1543,N_1505);
and U1569 (N_1569,N_1516,N_1537);
and U1570 (N_1570,N_1506,N_1512);
or U1571 (N_1571,N_1503,N_1547);
nor U1572 (N_1572,N_1523,N_1558);
and U1573 (N_1573,N_1542,N_1546);
xor U1574 (N_1574,N_1520,N_1500);
or U1575 (N_1575,N_1530,N_1509);
nor U1576 (N_1576,N_1522,N_1501);
or U1577 (N_1577,N_1526,N_1552);
and U1578 (N_1578,N_1511,N_1544);
or U1579 (N_1579,N_1527,N_1549);
nor U1580 (N_1580,N_1507,N_1533);
and U1581 (N_1581,N_1540,N_1556);
or U1582 (N_1582,N_1534,N_1528);
or U1583 (N_1583,N_1521,N_1510);
and U1584 (N_1584,N_1551,N_1555);
nand U1585 (N_1585,N_1508,N_1504);
nor U1586 (N_1586,N_1519,N_1559);
or U1587 (N_1587,N_1548,N_1535);
or U1588 (N_1588,N_1550,N_1532);
nor U1589 (N_1589,N_1536,N_1515);
xor U1590 (N_1590,N_1521,N_1534);
xnor U1591 (N_1591,N_1524,N_1523);
or U1592 (N_1592,N_1527,N_1515);
or U1593 (N_1593,N_1530,N_1548);
nor U1594 (N_1594,N_1538,N_1539);
nor U1595 (N_1595,N_1508,N_1530);
nand U1596 (N_1596,N_1512,N_1539);
nor U1597 (N_1597,N_1514,N_1516);
or U1598 (N_1598,N_1526,N_1517);
nand U1599 (N_1599,N_1519,N_1546);
or U1600 (N_1600,N_1533,N_1536);
nand U1601 (N_1601,N_1537,N_1548);
and U1602 (N_1602,N_1500,N_1518);
nor U1603 (N_1603,N_1501,N_1500);
or U1604 (N_1604,N_1503,N_1525);
nor U1605 (N_1605,N_1531,N_1505);
nor U1606 (N_1606,N_1517,N_1532);
or U1607 (N_1607,N_1530,N_1500);
or U1608 (N_1608,N_1503,N_1528);
or U1609 (N_1609,N_1505,N_1507);
nand U1610 (N_1610,N_1530,N_1543);
or U1611 (N_1611,N_1536,N_1519);
and U1612 (N_1612,N_1540,N_1535);
or U1613 (N_1613,N_1538,N_1541);
and U1614 (N_1614,N_1500,N_1529);
and U1615 (N_1615,N_1541,N_1554);
nand U1616 (N_1616,N_1525,N_1517);
nor U1617 (N_1617,N_1553,N_1503);
xor U1618 (N_1618,N_1542,N_1524);
nand U1619 (N_1619,N_1505,N_1541);
or U1620 (N_1620,N_1566,N_1585);
nor U1621 (N_1621,N_1613,N_1596);
nor U1622 (N_1622,N_1610,N_1607);
or U1623 (N_1623,N_1570,N_1562);
or U1624 (N_1624,N_1594,N_1615);
or U1625 (N_1625,N_1567,N_1586);
nor U1626 (N_1626,N_1589,N_1600);
nand U1627 (N_1627,N_1606,N_1608);
xnor U1628 (N_1628,N_1599,N_1584);
nand U1629 (N_1629,N_1602,N_1565);
nand U1630 (N_1630,N_1619,N_1590);
or U1631 (N_1631,N_1616,N_1568);
or U1632 (N_1632,N_1593,N_1579);
and U1633 (N_1633,N_1595,N_1601);
nand U1634 (N_1634,N_1614,N_1577);
or U1635 (N_1635,N_1560,N_1603);
or U1636 (N_1636,N_1578,N_1580);
nand U1637 (N_1637,N_1612,N_1597);
nor U1638 (N_1638,N_1588,N_1582);
and U1639 (N_1639,N_1605,N_1575);
and U1640 (N_1640,N_1576,N_1592);
nand U1641 (N_1641,N_1598,N_1587);
nand U1642 (N_1642,N_1573,N_1617);
or U1643 (N_1643,N_1563,N_1583);
or U1644 (N_1644,N_1571,N_1581);
nor U1645 (N_1645,N_1564,N_1561);
xor U1646 (N_1646,N_1604,N_1574);
or U1647 (N_1647,N_1611,N_1609);
nor U1648 (N_1648,N_1618,N_1572);
and U1649 (N_1649,N_1569,N_1591);
and U1650 (N_1650,N_1563,N_1593);
and U1651 (N_1651,N_1609,N_1615);
xnor U1652 (N_1652,N_1586,N_1615);
nand U1653 (N_1653,N_1577,N_1584);
or U1654 (N_1654,N_1563,N_1596);
and U1655 (N_1655,N_1580,N_1592);
or U1656 (N_1656,N_1613,N_1589);
nand U1657 (N_1657,N_1590,N_1609);
nor U1658 (N_1658,N_1615,N_1601);
nor U1659 (N_1659,N_1611,N_1596);
and U1660 (N_1660,N_1568,N_1607);
nand U1661 (N_1661,N_1603,N_1596);
and U1662 (N_1662,N_1612,N_1602);
and U1663 (N_1663,N_1601,N_1596);
nor U1664 (N_1664,N_1567,N_1592);
nand U1665 (N_1665,N_1594,N_1563);
or U1666 (N_1666,N_1617,N_1613);
nand U1667 (N_1667,N_1582,N_1586);
nand U1668 (N_1668,N_1569,N_1618);
nor U1669 (N_1669,N_1613,N_1563);
nand U1670 (N_1670,N_1598,N_1596);
nor U1671 (N_1671,N_1566,N_1571);
nand U1672 (N_1672,N_1591,N_1619);
nand U1673 (N_1673,N_1564,N_1588);
nor U1674 (N_1674,N_1598,N_1562);
xnor U1675 (N_1675,N_1599,N_1560);
nor U1676 (N_1676,N_1570,N_1601);
nor U1677 (N_1677,N_1595,N_1586);
nand U1678 (N_1678,N_1608,N_1586);
nand U1679 (N_1679,N_1596,N_1560);
nand U1680 (N_1680,N_1635,N_1665);
or U1681 (N_1681,N_1669,N_1621);
nand U1682 (N_1682,N_1642,N_1626);
or U1683 (N_1683,N_1667,N_1623);
nand U1684 (N_1684,N_1662,N_1622);
or U1685 (N_1685,N_1633,N_1632);
nor U1686 (N_1686,N_1671,N_1655);
nor U1687 (N_1687,N_1663,N_1627);
or U1688 (N_1688,N_1654,N_1630);
and U1689 (N_1689,N_1638,N_1677);
or U1690 (N_1690,N_1624,N_1674);
and U1691 (N_1691,N_1636,N_1668);
or U1692 (N_1692,N_1678,N_1652);
and U1693 (N_1693,N_1666,N_1649);
and U1694 (N_1694,N_1679,N_1670);
nor U1695 (N_1695,N_1659,N_1631);
nor U1696 (N_1696,N_1629,N_1672);
nand U1697 (N_1697,N_1643,N_1675);
or U1698 (N_1698,N_1637,N_1641);
xor U1699 (N_1699,N_1628,N_1676);
nand U1700 (N_1700,N_1650,N_1647);
nand U1701 (N_1701,N_1661,N_1664);
and U1702 (N_1702,N_1658,N_1625);
and U1703 (N_1703,N_1640,N_1644);
and U1704 (N_1704,N_1645,N_1653);
nand U1705 (N_1705,N_1639,N_1656);
or U1706 (N_1706,N_1634,N_1646);
or U1707 (N_1707,N_1657,N_1651);
or U1708 (N_1708,N_1673,N_1648);
or U1709 (N_1709,N_1620,N_1660);
or U1710 (N_1710,N_1642,N_1676);
and U1711 (N_1711,N_1631,N_1669);
nor U1712 (N_1712,N_1654,N_1621);
and U1713 (N_1713,N_1669,N_1666);
or U1714 (N_1714,N_1643,N_1634);
xnor U1715 (N_1715,N_1633,N_1625);
nor U1716 (N_1716,N_1667,N_1672);
and U1717 (N_1717,N_1669,N_1655);
xor U1718 (N_1718,N_1649,N_1626);
nor U1719 (N_1719,N_1669,N_1667);
and U1720 (N_1720,N_1639,N_1669);
and U1721 (N_1721,N_1628,N_1663);
nand U1722 (N_1722,N_1659,N_1676);
or U1723 (N_1723,N_1636,N_1679);
or U1724 (N_1724,N_1666,N_1641);
nor U1725 (N_1725,N_1635,N_1637);
xnor U1726 (N_1726,N_1653,N_1643);
nand U1727 (N_1727,N_1641,N_1631);
nor U1728 (N_1728,N_1633,N_1638);
nor U1729 (N_1729,N_1634,N_1666);
nand U1730 (N_1730,N_1640,N_1658);
or U1731 (N_1731,N_1622,N_1658);
nor U1732 (N_1732,N_1625,N_1661);
nand U1733 (N_1733,N_1673,N_1663);
nor U1734 (N_1734,N_1628,N_1647);
nand U1735 (N_1735,N_1621,N_1675);
nor U1736 (N_1736,N_1653,N_1623);
nand U1737 (N_1737,N_1655,N_1639);
or U1738 (N_1738,N_1669,N_1664);
or U1739 (N_1739,N_1656,N_1661);
nand U1740 (N_1740,N_1736,N_1708);
nor U1741 (N_1741,N_1689,N_1701);
and U1742 (N_1742,N_1706,N_1735);
or U1743 (N_1743,N_1711,N_1719);
xnor U1744 (N_1744,N_1690,N_1728);
xnor U1745 (N_1745,N_1731,N_1727);
nor U1746 (N_1746,N_1681,N_1702);
and U1747 (N_1747,N_1691,N_1723);
nor U1748 (N_1748,N_1682,N_1713);
nor U1749 (N_1749,N_1704,N_1739);
or U1750 (N_1750,N_1700,N_1717);
nand U1751 (N_1751,N_1707,N_1714);
or U1752 (N_1752,N_1715,N_1693);
nor U1753 (N_1753,N_1709,N_1725);
or U1754 (N_1754,N_1697,N_1685);
nor U1755 (N_1755,N_1712,N_1734);
and U1756 (N_1756,N_1686,N_1683);
nor U1757 (N_1757,N_1732,N_1698);
nand U1758 (N_1758,N_1733,N_1696);
nor U1759 (N_1759,N_1692,N_1699);
xor U1760 (N_1760,N_1738,N_1694);
or U1761 (N_1761,N_1687,N_1724);
nand U1762 (N_1762,N_1710,N_1737);
nor U1763 (N_1763,N_1729,N_1703);
and U1764 (N_1764,N_1695,N_1730);
nand U1765 (N_1765,N_1720,N_1721);
or U1766 (N_1766,N_1705,N_1680);
or U1767 (N_1767,N_1718,N_1684);
xor U1768 (N_1768,N_1688,N_1726);
or U1769 (N_1769,N_1716,N_1722);
xnor U1770 (N_1770,N_1707,N_1694);
xnor U1771 (N_1771,N_1730,N_1737);
nand U1772 (N_1772,N_1732,N_1688);
or U1773 (N_1773,N_1728,N_1704);
or U1774 (N_1774,N_1724,N_1705);
or U1775 (N_1775,N_1726,N_1703);
and U1776 (N_1776,N_1687,N_1736);
nor U1777 (N_1777,N_1709,N_1739);
nand U1778 (N_1778,N_1687,N_1716);
and U1779 (N_1779,N_1726,N_1713);
nand U1780 (N_1780,N_1701,N_1727);
nor U1781 (N_1781,N_1686,N_1701);
or U1782 (N_1782,N_1691,N_1701);
and U1783 (N_1783,N_1733,N_1724);
or U1784 (N_1784,N_1689,N_1700);
and U1785 (N_1785,N_1717,N_1720);
or U1786 (N_1786,N_1721,N_1723);
or U1787 (N_1787,N_1696,N_1686);
or U1788 (N_1788,N_1684,N_1699);
xnor U1789 (N_1789,N_1706,N_1716);
and U1790 (N_1790,N_1694,N_1693);
xnor U1791 (N_1791,N_1737,N_1683);
nor U1792 (N_1792,N_1691,N_1728);
and U1793 (N_1793,N_1724,N_1693);
and U1794 (N_1794,N_1738,N_1722);
nand U1795 (N_1795,N_1726,N_1699);
nand U1796 (N_1796,N_1730,N_1704);
xor U1797 (N_1797,N_1724,N_1696);
and U1798 (N_1798,N_1687,N_1696);
or U1799 (N_1799,N_1682,N_1699);
nand U1800 (N_1800,N_1786,N_1765);
and U1801 (N_1801,N_1789,N_1796);
and U1802 (N_1802,N_1793,N_1764);
or U1803 (N_1803,N_1769,N_1760);
or U1804 (N_1804,N_1773,N_1788);
nand U1805 (N_1805,N_1744,N_1777);
or U1806 (N_1806,N_1785,N_1790);
or U1807 (N_1807,N_1740,N_1795);
or U1808 (N_1808,N_1761,N_1745);
or U1809 (N_1809,N_1757,N_1741);
nor U1810 (N_1810,N_1780,N_1783);
or U1811 (N_1811,N_1799,N_1784);
nand U1812 (N_1812,N_1742,N_1797);
and U1813 (N_1813,N_1794,N_1748);
nor U1814 (N_1814,N_1782,N_1791);
nor U1815 (N_1815,N_1749,N_1752);
nand U1816 (N_1816,N_1746,N_1798);
nand U1817 (N_1817,N_1792,N_1754);
and U1818 (N_1818,N_1778,N_1768);
or U1819 (N_1819,N_1787,N_1771);
and U1820 (N_1820,N_1772,N_1751);
nor U1821 (N_1821,N_1743,N_1762);
nand U1822 (N_1822,N_1759,N_1781);
nor U1823 (N_1823,N_1779,N_1753);
or U1824 (N_1824,N_1776,N_1766);
nand U1825 (N_1825,N_1774,N_1758);
or U1826 (N_1826,N_1770,N_1763);
or U1827 (N_1827,N_1750,N_1767);
xor U1828 (N_1828,N_1747,N_1756);
nor U1829 (N_1829,N_1775,N_1755);
nor U1830 (N_1830,N_1741,N_1774);
or U1831 (N_1831,N_1778,N_1743);
xor U1832 (N_1832,N_1779,N_1747);
nand U1833 (N_1833,N_1775,N_1786);
nand U1834 (N_1834,N_1782,N_1794);
and U1835 (N_1835,N_1788,N_1759);
or U1836 (N_1836,N_1751,N_1759);
nand U1837 (N_1837,N_1772,N_1767);
and U1838 (N_1838,N_1778,N_1755);
nor U1839 (N_1839,N_1747,N_1745);
nor U1840 (N_1840,N_1759,N_1778);
and U1841 (N_1841,N_1790,N_1757);
nand U1842 (N_1842,N_1748,N_1777);
and U1843 (N_1843,N_1780,N_1755);
xnor U1844 (N_1844,N_1762,N_1748);
nand U1845 (N_1845,N_1746,N_1754);
xnor U1846 (N_1846,N_1770,N_1782);
and U1847 (N_1847,N_1777,N_1761);
and U1848 (N_1848,N_1782,N_1758);
nand U1849 (N_1849,N_1783,N_1778);
nor U1850 (N_1850,N_1782,N_1774);
or U1851 (N_1851,N_1760,N_1768);
nand U1852 (N_1852,N_1744,N_1749);
nand U1853 (N_1853,N_1786,N_1742);
and U1854 (N_1854,N_1741,N_1784);
or U1855 (N_1855,N_1746,N_1797);
nand U1856 (N_1856,N_1786,N_1790);
nand U1857 (N_1857,N_1783,N_1758);
or U1858 (N_1858,N_1793,N_1780);
or U1859 (N_1859,N_1790,N_1750);
and U1860 (N_1860,N_1842,N_1850);
and U1861 (N_1861,N_1811,N_1809);
and U1862 (N_1862,N_1859,N_1816);
or U1863 (N_1863,N_1819,N_1808);
nand U1864 (N_1864,N_1838,N_1835);
nor U1865 (N_1865,N_1840,N_1857);
nand U1866 (N_1866,N_1800,N_1803);
or U1867 (N_1867,N_1831,N_1805);
nor U1868 (N_1868,N_1820,N_1814);
or U1869 (N_1869,N_1802,N_1834);
nand U1870 (N_1870,N_1823,N_1806);
or U1871 (N_1871,N_1858,N_1810);
nand U1872 (N_1872,N_1801,N_1822);
or U1873 (N_1873,N_1833,N_1836);
nand U1874 (N_1874,N_1827,N_1813);
nand U1875 (N_1875,N_1841,N_1825);
and U1876 (N_1876,N_1812,N_1843);
nor U1877 (N_1877,N_1837,N_1826);
and U1878 (N_1878,N_1845,N_1815);
and U1879 (N_1879,N_1848,N_1804);
or U1880 (N_1880,N_1854,N_1824);
or U1881 (N_1881,N_1847,N_1853);
xnor U1882 (N_1882,N_1829,N_1828);
or U1883 (N_1883,N_1852,N_1849);
and U1884 (N_1884,N_1846,N_1856);
nand U1885 (N_1885,N_1818,N_1832);
or U1886 (N_1886,N_1807,N_1817);
xor U1887 (N_1887,N_1855,N_1821);
and U1888 (N_1888,N_1844,N_1839);
nand U1889 (N_1889,N_1851,N_1830);
or U1890 (N_1890,N_1837,N_1839);
or U1891 (N_1891,N_1807,N_1832);
and U1892 (N_1892,N_1827,N_1844);
or U1893 (N_1893,N_1826,N_1810);
and U1894 (N_1894,N_1804,N_1845);
and U1895 (N_1895,N_1845,N_1856);
xnor U1896 (N_1896,N_1859,N_1801);
xnor U1897 (N_1897,N_1844,N_1830);
nand U1898 (N_1898,N_1818,N_1847);
and U1899 (N_1899,N_1807,N_1843);
nand U1900 (N_1900,N_1802,N_1822);
nor U1901 (N_1901,N_1827,N_1859);
or U1902 (N_1902,N_1854,N_1843);
or U1903 (N_1903,N_1808,N_1811);
nor U1904 (N_1904,N_1857,N_1825);
nand U1905 (N_1905,N_1850,N_1851);
or U1906 (N_1906,N_1805,N_1832);
xor U1907 (N_1907,N_1832,N_1809);
and U1908 (N_1908,N_1859,N_1831);
xnor U1909 (N_1909,N_1820,N_1852);
and U1910 (N_1910,N_1823,N_1815);
and U1911 (N_1911,N_1835,N_1827);
nor U1912 (N_1912,N_1835,N_1829);
nand U1913 (N_1913,N_1812,N_1831);
and U1914 (N_1914,N_1840,N_1805);
nand U1915 (N_1915,N_1804,N_1813);
and U1916 (N_1916,N_1821,N_1842);
nor U1917 (N_1917,N_1840,N_1842);
nor U1918 (N_1918,N_1802,N_1841);
nand U1919 (N_1919,N_1856,N_1811);
nor U1920 (N_1920,N_1895,N_1907);
xor U1921 (N_1921,N_1918,N_1901);
nor U1922 (N_1922,N_1881,N_1899);
nor U1923 (N_1923,N_1887,N_1904);
xnor U1924 (N_1924,N_1884,N_1885);
xor U1925 (N_1925,N_1894,N_1900);
nor U1926 (N_1926,N_1903,N_1908);
nand U1927 (N_1927,N_1898,N_1917);
nand U1928 (N_1928,N_1875,N_1911);
xnor U1929 (N_1929,N_1862,N_1876);
nor U1930 (N_1930,N_1906,N_1902);
or U1931 (N_1931,N_1860,N_1912);
nor U1932 (N_1932,N_1874,N_1892);
nand U1933 (N_1933,N_1913,N_1896);
and U1934 (N_1934,N_1905,N_1890);
or U1935 (N_1935,N_1868,N_1877);
nand U1936 (N_1936,N_1871,N_1897);
nor U1937 (N_1937,N_1916,N_1909);
nand U1938 (N_1938,N_1865,N_1915);
and U1939 (N_1939,N_1866,N_1910);
and U1940 (N_1940,N_1864,N_1861);
and U1941 (N_1941,N_1872,N_1888);
nor U1942 (N_1942,N_1919,N_1878);
or U1943 (N_1943,N_1867,N_1883);
nand U1944 (N_1944,N_1880,N_1886);
and U1945 (N_1945,N_1889,N_1891);
nand U1946 (N_1946,N_1879,N_1914);
xor U1947 (N_1947,N_1869,N_1863);
and U1948 (N_1948,N_1873,N_1882);
nor U1949 (N_1949,N_1893,N_1870);
and U1950 (N_1950,N_1898,N_1868);
nand U1951 (N_1951,N_1871,N_1876);
or U1952 (N_1952,N_1885,N_1901);
nor U1953 (N_1953,N_1893,N_1860);
and U1954 (N_1954,N_1917,N_1905);
nor U1955 (N_1955,N_1875,N_1862);
nor U1956 (N_1956,N_1885,N_1866);
nand U1957 (N_1957,N_1883,N_1900);
nand U1958 (N_1958,N_1868,N_1863);
and U1959 (N_1959,N_1893,N_1866);
nor U1960 (N_1960,N_1890,N_1910);
and U1961 (N_1961,N_1915,N_1902);
nand U1962 (N_1962,N_1903,N_1875);
and U1963 (N_1963,N_1867,N_1861);
nor U1964 (N_1964,N_1881,N_1904);
and U1965 (N_1965,N_1884,N_1892);
or U1966 (N_1966,N_1909,N_1886);
nand U1967 (N_1967,N_1881,N_1860);
nand U1968 (N_1968,N_1904,N_1878);
and U1969 (N_1969,N_1901,N_1861);
and U1970 (N_1970,N_1888,N_1870);
nor U1971 (N_1971,N_1874,N_1904);
or U1972 (N_1972,N_1871,N_1904);
nand U1973 (N_1973,N_1868,N_1919);
nor U1974 (N_1974,N_1907,N_1863);
nor U1975 (N_1975,N_1901,N_1868);
nor U1976 (N_1976,N_1899,N_1885);
or U1977 (N_1977,N_1915,N_1877);
nand U1978 (N_1978,N_1892,N_1865);
nor U1979 (N_1979,N_1875,N_1868);
nor U1980 (N_1980,N_1960,N_1970);
nor U1981 (N_1981,N_1924,N_1928);
and U1982 (N_1982,N_1929,N_1933);
xor U1983 (N_1983,N_1979,N_1978);
and U1984 (N_1984,N_1935,N_1938);
or U1985 (N_1985,N_1921,N_1959);
or U1986 (N_1986,N_1947,N_1977);
or U1987 (N_1987,N_1930,N_1942);
nor U1988 (N_1988,N_1951,N_1932);
or U1989 (N_1989,N_1952,N_1941);
and U1990 (N_1990,N_1965,N_1948);
or U1991 (N_1991,N_1926,N_1920);
nor U1992 (N_1992,N_1969,N_1976);
nand U1993 (N_1993,N_1923,N_1967);
or U1994 (N_1994,N_1949,N_1937);
or U1995 (N_1995,N_1973,N_1954);
and U1996 (N_1996,N_1944,N_1931);
or U1997 (N_1997,N_1946,N_1972);
nand U1998 (N_1998,N_1975,N_1971);
or U1999 (N_1999,N_1925,N_1974);
and U2000 (N_2000,N_1950,N_1961);
and U2001 (N_2001,N_1955,N_1958);
nand U2002 (N_2002,N_1963,N_1964);
nand U2003 (N_2003,N_1957,N_1953);
nand U2004 (N_2004,N_1968,N_1936);
and U2005 (N_2005,N_1945,N_1943);
and U2006 (N_2006,N_1927,N_1962);
xor U2007 (N_2007,N_1934,N_1966);
or U2008 (N_2008,N_1939,N_1940);
nor U2009 (N_2009,N_1922,N_1956);
nor U2010 (N_2010,N_1946,N_1957);
nor U2011 (N_2011,N_1957,N_1958);
and U2012 (N_2012,N_1968,N_1949);
and U2013 (N_2013,N_1924,N_1937);
xor U2014 (N_2014,N_1968,N_1961);
and U2015 (N_2015,N_1943,N_1964);
nand U2016 (N_2016,N_1966,N_1974);
or U2017 (N_2017,N_1965,N_1971);
and U2018 (N_2018,N_1979,N_1941);
or U2019 (N_2019,N_1939,N_1936);
nor U2020 (N_2020,N_1926,N_1923);
nor U2021 (N_2021,N_1976,N_1947);
or U2022 (N_2022,N_1928,N_1925);
nor U2023 (N_2023,N_1958,N_1975);
nor U2024 (N_2024,N_1953,N_1947);
xnor U2025 (N_2025,N_1932,N_1933);
or U2026 (N_2026,N_1927,N_1977);
xor U2027 (N_2027,N_1946,N_1945);
or U2028 (N_2028,N_1928,N_1945);
or U2029 (N_2029,N_1956,N_1972);
xnor U2030 (N_2030,N_1972,N_1978);
nor U2031 (N_2031,N_1920,N_1942);
and U2032 (N_2032,N_1922,N_1946);
nand U2033 (N_2033,N_1935,N_1947);
and U2034 (N_2034,N_1963,N_1957);
nor U2035 (N_2035,N_1940,N_1942);
nor U2036 (N_2036,N_1948,N_1951);
nor U2037 (N_2037,N_1947,N_1923);
and U2038 (N_2038,N_1968,N_1931);
nand U2039 (N_2039,N_1951,N_1961);
or U2040 (N_2040,N_1995,N_2026);
or U2041 (N_2041,N_2024,N_2004);
and U2042 (N_2042,N_2007,N_2034);
nor U2043 (N_2043,N_2028,N_2008);
and U2044 (N_2044,N_2033,N_2022);
and U2045 (N_2045,N_1986,N_2019);
nor U2046 (N_2046,N_2037,N_1992);
nor U2047 (N_2047,N_1989,N_1998);
nand U2048 (N_2048,N_1982,N_2021);
xnor U2049 (N_2049,N_2039,N_1983);
or U2050 (N_2050,N_2035,N_2002);
or U2051 (N_2051,N_2016,N_1985);
and U2052 (N_2052,N_1996,N_2000);
nor U2053 (N_2053,N_1988,N_1997);
nand U2054 (N_2054,N_1990,N_1981);
nand U2055 (N_2055,N_2015,N_2009);
or U2056 (N_2056,N_2018,N_2010);
nand U2057 (N_2057,N_2013,N_1980);
nand U2058 (N_2058,N_2029,N_2027);
or U2059 (N_2059,N_2017,N_2038);
nor U2060 (N_2060,N_1987,N_1984);
nand U2061 (N_2061,N_2005,N_2030);
nand U2062 (N_2062,N_1993,N_1991);
nand U2063 (N_2063,N_2032,N_1999);
or U2064 (N_2064,N_2001,N_2011);
xnor U2065 (N_2065,N_2025,N_2006);
nand U2066 (N_2066,N_2003,N_2014);
or U2067 (N_2067,N_2036,N_2020);
nor U2068 (N_2068,N_2023,N_1994);
xor U2069 (N_2069,N_2031,N_2012);
nor U2070 (N_2070,N_2020,N_1998);
or U2071 (N_2071,N_2034,N_1987);
nand U2072 (N_2072,N_2004,N_2009);
nor U2073 (N_2073,N_2007,N_1982);
and U2074 (N_2074,N_1987,N_2023);
or U2075 (N_2075,N_1988,N_1999);
nor U2076 (N_2076,N_2016,N_1991);
or U2077 (N_2077,N_2001,N_1986);
nor U2078 (N_2078,N_2011,N_2006);
or U2079 (N_2079,N_2001,N_2036);
nand U2080 (N_2080,N_2029,N_1988);
and U2081 (N_2081,N_1993,N_2033);
nand U2082 (N_2082,N_1997,N_1986);
or U2083 (N_2083,N_2028,N_2006);
nand U2084 (N_2084,N_2038,N_1999);
nor U2085 (N_2085,N_2008,N_2004);
and U2086 (N_2086,N_2021,N_2023);
or U2087 (N_2087,N_2038,N_1983);
or U2088 (N_2088,N_1991,N_2004);
nor U2089 (N_2089,N_1999,N_2028);
nor U2090 (N_2090,N_1988,N_2034);
and U2091 (N_2091,N_2000,N_1997);
or U2092 (N_2092,N_1989,N_1993);
xnor U2093 (N_2093,N_2023,N_2001);
nor U2094 (N_2094,N_2036,N_1989);
nand U2095 (N_2095,N_1984,N_2016);
and U2096 (N_2096,N_1988,N_2006);
and U2097 (N_2097,N_2029,N_1997);
nor U2098 (N_2098,N_2002,N_2030);
and U2099 (N_2099,N_2038,N_2005);
or U2100 (N_2100,N_2092,N_2064);
nand U2101 (N_2101,N_2068,N_2043);
xnor U2102 (N_2102,N_2047,N_2074);
nor U2103 (N_2103,N_2040,N_2069);
xnor U2104 (N_2104,N_2071,N_2086);
xor U2105 (N_2105,N_2063,N_2093);
and U2106 (N_2106,N_2081,N_2080);
or U2107 (N_2107,N_2089,N_2061);
nor U2108 (N_2108,N_2050,N_2075);
nor U2109 (N_2109,N_2044,N_2060);
nand U2110 (N_2110,N_2049,N_2076);
and U2111 (N_2111,N_2082,N_2085);
xnor U2112 (N_2112,N_2087,N_2098);
nand U2113 (N_2113,N_2051,N_2042);
nand U2114 (N_2114,N_2097,N_2083);
xnor U2115 (N_2115,N_2079,N_2090);
or U2116 (N_2116,N_2091,N_2055);
nor U2117 (N_2117,N_2062,N_2067);
or U2118 (N_2118,N_2095,N_2084);
nand U2119 (N_2119,N_2046,N_2059);
xnor U2120 (N_2120,N_2057,N_2072);
nand U2121 (N_2121,N_2078,N_2099);
nand U2122 (N_2122,N_2053,N_2070);
xor U2123 (N_2123,N_2065,N_2094);
and U2124 (N_2124,N_2052,N_2096);
or U2125 (N_2125,N_2048,N_2041);
nor U2126 (N_2126,N_2077,N_2088);
or U2127 (N_2127,N_2045,N_2073);
and U2128 (N_2128,N_2058,N_2066);
and U2129 (N_2129,N_2054,N_2056);
nor U2130 (N_2130,N_2091,N_2079);
nor U2131 (N_2131,N_2042,N_2071);
nand U2132 (N_2132,N_2049,N_2046);
or U2133 (N_2133,N_2041,N_2051);
and U2134 (N_2134,N_2095,N_2044);
and U2135 (N_2135,N_2092,N_2085);
xnor U2136 (N_2136,N_2049,N_2091);
nand U2137 (N_2137,N_2054,N_2092);
nor U2138 (N_2138,N_2070,N_2093);
xnor U2139 (N_2139,N_2074,N_2084);
and U2140 (N_2140,N_2059,N_2068);
nor U2141 (N_2141,N_2090,N_2064);
nor U2142 (N_2142,N_2098,N_2044);
xor U2143 (N_2143,N_2053,N_2084);
and U2144 (N_2144,N_2096,N_2058);
or U2145 (N_2145,N_2040,N_2073);
nand U2146 (N_2146,N_2050,N_2044);
or U2147 (N_2147,N_2054,N_2072);
nand U2148 (N_2148,N_2091,N_2083);
nand U2149 (N_2149,N_2093,N_2040);
nor U2150 (N_2150,N_2061,N_2080);
or U2151 (N_2151,N_2083,N_2045);
nand U2152 (N_2152,N_2042,N_2062);
and U2153 (N_2153,N_2049,N_2096);
xor U2154 (N_2154,N_2064,N_2097);
or U2155 (N_2155,N_2077,N_2090);
nand U2156 (N_2156,N_2095,N_2074);
nand U2157 (N_2157,N_2059,N_2047);
nand U2158 (N_2158,N_2060,N_2065);
nor U2159 (N_2159,N_2055,N_2044);
or U2160 (N_2160,N_2114,N_2147);
nand U2161 (N_2161,N_2153,N_2151);
or U2162 (N_2162,N_2133,N_2122);
nor U2163 (N_2163,N_2116,N_2132);
nor U2164 (N_2164,N_2112,N_2141);
and U2165 (N_2165,N_2146,N_2138);
nor U2166 (N_2166,N_2125,N_2148);
nor U2167 (N_2167,N_2140,N_2123);
nand U2168 (N_2168,N_2113,N_2120);
nand U2169 (N_2169,N_2152,N_2142);
or U2170 (N_2170,N_2104,N_2156);
nand U2171 (N_2171,N_2118,N_2105);
nor U2172 (N_2172,N_2106,N_2108);
nor U2173 (N_2173,N_2115,N_2145);
or U2174 (N_2174,N_2111,N_2149);
or U2175 (N_2175,N_2102,N_2124);
nor U2176 (N_2176,N_2103,N_2150);
nand U2177 (N_2177,N_2127,N_2135);
or U2178 (N_2178,N_2109,N_2130);
xnor U2179 (N_2179,N_2134,N_2159);
xor U2180 (N_2180,N_2137,N_2157);
and U2181 (N_2181,N_2128,N_2129);
and U2182 (N_2182,N_2119,N_2101);
nand U2183 (N_2183,N_2155,N_2107);
nand U2184 (N_2184,N_2144,N_2143);
nor U2185 (N_2185,N_2136,N_2117);
nor U2186 (N_2186,N_2110,N_2139);
nand U2187 (N_2187,N_2158,N_2126);
or U2188 (N_2188,N_2131,N_2154);
nand U2189 (N_2189,N_2121,N_2100);
nand U2190 (N_2190,N_2110,N_2117);
or U2191 (N_2191,N_2118,N_2115);
or U2192 (N_2192,N_2124,N_2127);
xnor U2193 (N_2193,N_2117,N_2113);
nand U2194 (N_2194,N_2145,N_2141);
nor U2195 (N_2195,N_2137,N_2142);
or U2196 (N_2196,N_2132,N_2123);
nand U2197 (N_2197,N_2110,N_2121);
or U2198 (N_2198,N_2155,N_2137);
or U2199 (N_2199,N_2150,N_2108);
or U2200 (N_2200,N_2120,N_2153);
nand U2201 (N_2201,N_2154,N_2143);
and U2202 (N_2202,N_2100,N_2150);
or U2203 (N_2203,N_2146,N_2149);
or U2204 (N_2204,N_2144,N_2158);
or U2205 (N_2205,N_2143,N_2111);
or U2206 (N_2206,N_2147,N_2149);
and U2207 (N_2207,N_2104,N_2136);
nand U2208 (N_2208,N_2119,N_2122);
nor U2209 (N_2209,N_2143,N_2150);
nor U2210 (N_2210,N_2115,N_2135);
and U2211 (N_2211,N_2116,N_2130);
or U2212 (N_2212,N_2131,N_2130);
nand U2213 (N_2213,N_2159,N_2121);
nor U2214 (N_2214,N_2117,N_2143);
or U2215 (N_2215,N_2116,N_2127);
or U2216 (N_2216,N_2156,N_2152);
nand U2217 (N_2217,N_2144,N_2112);
xnor U2218 (N_2218,N_2101,N_2111);
xnor U2219 (N_2219,N_2135,N_2154);
nand U2220 (N_2220,N_2218,N_2211);
xnor U2221 (N_2221,N_2215,N_2202);
and U2222 (N_2222,N_2216,N_2205);
xnor U2223 (N_2223,N_2190,N_2168);
xor U2224 (N_2224,N_2192,N_2176);
xor U2225 (N_2225,N_2167,N_2173);
and U2226 (N_2226,N_2193,N_2179);
or U2227 (N_2227,N_2214,N_2178);
nor U2228 (N_2228,N_2180,N_2194);
and U2229 (N_2229,N_2203,N_2208);
or U2230 (N_2230,N_2166,N_2172);
or U2231 (N_2231,N_2206,N_2177);
xnor U2232 (N_2232,N_2183,N_2219);
nor U2233 (N_2233,N_2164,N_2201);
and U2234 (N_2234,N_2161,N_2182);
nand U2235 (N_2235,N_2162,N_2213);
or U2236 (N_2236,N_2160,N_2191);
xor U2237 (N_2237,N_2204,N_2163);
nand U2238 (N_2238,N_2196,N_2210);
or U2239 (N_2239,N_2212,N_2199);
and U2240 (N_2240,N_2198,N_2197);
and U2241 (N_2241,N_2207,N_2174);
and U2242 (N_2242,N_2186,N_2217);
nand U2243 (N_2243,N_2170,N_2209);
and U2244 (N_2244,N_2200,N_2169);
nor U2245 (N_2245,N_2189,N_2188);
nor U2246 (N_2246,N_2165,N_2187);
nor U2247 (N_2247,N_2171,N_2181);
and U2248 (N_2248,N_2184,N_2195);
or U2249 (N_2249,N_2185,N_2175);
or U2250 (N_2250,N_2201,N_2197);
or U2251 (N_2251,N_2172,N_2162);
nor U2252 (N_2252,N_2219,N_2184);
nor U2253 (N_2253,N_2210,N_2164);
nor U2254 (N_2254,N_2160,N_2216);
nor U2255 (N_2255,N_2199,N_2174);
or U2256 (N_2256,N_2171,N_2173);
nor U2257 (N_2257,N_2174,N_2196);
xnor U2258 (N_2258,N_2209,N_2178);
nand U2259 (N_2259,N_2165,N_2176);
and U2260 (N_2260,N_2169,N_2207);
nor U2261 (N_2261,N_2170,N_2196);
xnor U2262 (N_2262,N_2206,N_2178);
nor U2263 (N_2263,N_2201,N_2204);
nor U2264 (N_2264,N_2162,N_2217);
nor U2265 (N_2265,N_2199,N_2185);
or U2266 (N_2266,N_2169,N_2185);
or U2267 (N_2267,N_2172,N_2180);
or U2268 (N_2268,N_2200,N_2192);
nand U2269 (N_2269,N_2193,N_2189);
xnor U2270 (N_2270,N_2198,N_2190);
nor U2271 (N_2271,N_2199,N_2215);
nand U2272 (N_2272,N_2216,N_2218);
or U2273 (N_2273,N_2201,N_2196);
nand U2274 (N_2274,N_2191,N_2161);
or U2275 (N_2275,N_2203,N_2175);
xnor U2276 (N_2276,N_2174,N_2163);
nand U2277 (N_2277,N_2189,N_2218);
nor U2278 (N_2278,N_2202,N_2191);
nor U2279 (N_2279,N_2166,N_2192);
nor U2280 (N_2280,N_2260,N_2236);
nor U2281 (N_2281,N_2254,N_2239);
nand U2282 (N_2282,N_2259,N_2258);
xnor U2283 (N_2283,N_2263,N_2242);
and U2284 (N_2284,N_2272,N_2257);
nor U2285 (N_2285,N_2221,N_2223);
nand U2286 (N_2286,N_2253,N_2249);
and U2287 (N_2287,N_2277,N_2237);
and U2288 (N_2288,N_2243,N_2271);
nand U2289 (N_2289,N_2251,N_2265);
nand U2290 (N_2290,N_2222,N_2276);
nand U2291 (N_2291,N_2256,N_2246);
and U2292 (N_2292,N_2240,N_2264);
nand U2293 (N_2293,N_2269,N_2231);
nand U2294 (N_2294,N_2274,N_2227);
nor U2295 (N_2295,N_2268,N_2229);
xor U2296 (N_2296,N_2279,N_2241);
nand U2297 (N_2297,N_2225,N_2270);
nand U2298 (N_2298,N_2248,N_2233);
or U2299 (N_2299,N_2275,N_2234);
and U2300 (N_2300,N_2266,N_2228);
nand U2301 (N_2301,N_2226,N_2220);
and U2302 (N_2302,N_2244,N_2273);
nor U2303 (N_2303,N_2252,N_2238);
and U2304 (N_2304,N_2261,N_2235);
or U2305 (N_2305,N_2262,N_2245);
and U2306 (N_2306,N_2255,N_2224);
xor U2307 (N_2307,N_2230,N_2247);
nand U2308 (N_2308,N_2267,N_2278);
nand U2309 (N_2309,N_2250,N_2232);
xor U2310 (N_2310,N_2231,N_2229);
or U2311 (N_2311,N_2226,N_2256);
and U2312 (N_2312,N_2274,N_2263);
xor U2313 (N_2313,N_2265,N_2241);
or U2314 (N_2314,N_2244,N_2260);
or U2315 (N_2315,N_2258,N_2276);
or U2316 (N_2316,N_2245,N_2225);
and U2317 (N_2317,N_2268,N_2252);
and U2318 (N_2318,N_2265,N_2267);
or U2319 (N_2319,N_2262,N_2223);
nor U2320 (N_2320,N_2249,N_2251);
and U2321 (N_2321,N_2225,N_2230);
and U2322 (N_2322,N_2233,N_2235);
or U2323 (N_2323,N_2272,N_2236);
nor U2324 (N_2324,N_2237,N_2230);
nand U2325 (N_2325,N_2238,N_2273);
and U2326 (N_2326,N_2235,N_2240);
nand U2327 (N_2327,N_2242,N_2239);
nand U2328 (N_2328,N_2251,N_2238);
xor U2329 (N_2329,N_2276,N_2271);
nor U2330 (N_2330,N_2262,N_2229);
xor U2331 (N_2331,N_2265,N_2270);
nand U2332 (N_2332,N_2257,N_2271);
and U2333 (N_2333,N_2270,N_2236);
nand U2334 (N_2334,N_2273,N_2225);
xor U2335 (N_2335,N_2261,N_2225);
nand U2336 (N_2336,N_2274,N_2257);
nand U2337 (N_2337,N_2275,N_2251);
and U2338 (N_2338,N_2258,N_2254);
and U2339 (N_2339,N_2277,N_2255);
and U2340 (N_2340,N_2336,N_2294);
nor U2341 (N_2341,N_2327,N_2318);
nor U2342 (N_2342,N_2320,N_2301);
nor U2343 (N_2343,N_2281,N_2300);
and U2344 (N_2344,N_2311,N_2332);
or U2345 (N_2345,N_2289,N_2334);
nand U2346 (N_2346,N_2291,N_2326);
nand U2347 (N_2347,N_2338,N_2297);
or U2348 (N_2348,N_2284,N_2295);
nor U2349 (N_2349,N_2305,N_2337);
nand U2350 (N_2350,N_2283,N_2298);
or U2351 (N_2351,N_2331,N_2299);
nand U2352 (N_2352,N_2319,N_2287);
nand U2353 (N_2353,N_2292,N_2315);
nand U2354 (N_2354,N_2290,N_2302);
and U2355 (N_2355,N_2280,N_2286);
and U2356 (N_2356,N_2328,N_2304);
and U2357 (N_2357,N_2309,N_2325);
or U2358 (N_2358,N_2312,N_2333);
or U2359 (N_2359,N_2310,N_2322);
nand U2360 (N_2360,N_2321,N_2316);
and U2361 (N_2361,N_2324,N_2314);
and U2362 (N_2362,N_2288,N_2282);
nand U2363 (N_2363,N_2323,N_2303);
and U2364 (N_2364,N_2313,N_2307);
nand U2365 (N_2365,N_2339,N_2308);
nand U2366 (N_2366,N_2285,N_2329);
nand U2367 (N_2367,N_2296,N_2317);
nor U2368 (N_2368,N_2306,N_2330);
and U2369 (N_2369,N_2293,N_2335);
nand U2370 (N_2370,N_2288,N_2317);
or U2371 (N_2371,N_2304,N_2280);
nand U2372 (N_2372,N_2339,N_2306);
or U2373 (N_2373,N_2318,N_2316);
or U2374 (N_2374,N_2316,N_2308);
xnor U2375 (N_2375,N_2321,N_2322);
nor U2376 (N_2376,N_2284,N_2325);
xnor U2377 (N_2377,N_2285,N_2287);
nand U2378 (N_2378,N_2296,N_2325);
and U2379 (N_2379,N_2288,N_2319);
nor U2380 (N_2380,N_2319,N_2308);
nor U2381 (N_2381,N_2287,N_2283);
xor U2382 (N_2382,N_2283,N_2324);
or U2383 (N_2383,N_2324,N_2281);
or U2384 (N_2384,N_2291,N_2332);
or U2385 (N_2385,N_2329,N_2284);
and U2386 (N_2386,N_2316,N_2311);
and U2387 (N_2387,N_2301,N_2283);
and U2388 (N_2388,N_2334,N_2286);
or U2389 (N_2389,N_2334,N_2325);
nand U2390 (N_2390,N_2287,N_2335);
or U2391 (N_2391,N_2333,N_2318);
or U2392 (N_2392,N_2294,N_2281);
nand U2393 (N_2393,N_2325,N_2324);
or U2394 (N_2394,N_2304,N_2310);
or U2395 (N_2395,N_2322,N_2298);
xnor U2396 (N_2396,N_2319,N_2332);
and U2397 (N_2397,N_2337,N_2311);
or U2398 (N_2398,N_2295,N_2310);
or U2399 (N_2399,N_2323,N_2316);
nor U2400 (N_2400,N_2385,N_2361);
nand U2401 (N_2401,N_2348,N_2381);
or U2402 (N_2402,N_2367,N_2376);
and U2403 (N_2403,N_2371,N_2347);
and U2404 (N_2404,N_2383,N_2360);
or U2405 (N_2405,N_2344,N_2364);
nor U2406 (N_2406,N_2378,N_2345);
or U2407 (N_2407,N_2370,N_2373);
or U2408 (N_2408,N_2392,N_2353);
and U2409 (N_2409,N_2390,N_2349);
nand U2410 (N_2410,N_2379,N_2350);
or U2411 (N_2411,N_2375,N_2386);
and U2412 (N_2412,N_2363,N_2391);
nand U2413 (N_2413,N_2359,N_2399);
or U2414 (N_2414,N_2374,N_2398);
and U2415 (N_2415,N_2397,N_2356);
nand U2416 (N_2416,N_2382,N_2369);
nor U2417 (N_2417,N_2387,N_2358);
or U2418 (N_2418,N_2341,N_2396);
nor U2419 (N_2419,N_2389,N_2377);
or U2420 (N_2420,N_2380,N_2340);
and U2421 (N_2421,N_2372,N_2354);
nand U2422 (N_2422,N_2394,N_2395);
nor U2423 (N_2423,N_2346,N_2365);
nand U2424 (N_2424,N_2357,N_2368);
or U2425 (N_2425,N_2393,N_2366);
and U2426 (N_2426,N_2355,N_2384);
or U2427 (N_2427,N_2343,N_2342);
xor U2428 (N_2428,N_2388,N_2362);
or U2429 (N_2429,N_2352,N_2351);
or U2430 (N_2430,N_2357,N_2353);
nand U2431 (N_2431,N_2375,N_2353);
and U2432 (N_2432,N_2379,N_2343);
and U2433 (N_2433,N_2380,N_2371);
or U2434 (N_2434,N_2366,N_2355);
or U2435 (N_2435,N_2386,N_2361);
nand U2436 (N_2436,N_2395,N_2379);
or U2437 (N_2437,N_2393,N_2387);
and U2438 (N_2438,N_2353,N_2388);
and U2439 (N_2439,N_2356,N_2350);
nor U2440 (N_2440,N_2378,N_2394);
nand U2441 (N_2441,N_2398,N_2343);
and U2442 (N_2442,N_2371,N_2352);
and U2443 (N_2443,N_2341,N_2386);
or U2444 (N_2444,N_2348,N_2393);
xnor U2445 (N_2445,N_2393,N_2364);
or U2446 (N_2446,N_2361,N_2378);
or U2447 (N_2447,N_2373,N_2354);
and U2448 (N_2448,N_2372,N_2363);
nand U2449 (N_2449,N_2388,N_2378);
nand U2450 (N_2450,N_2353,N_2346);
or U2451 (N_2451,N_2348,N_2355);
nor U2452 (N_2452,N_2382,N_2396);
nand U2453 (N_2453,N_2356,N_2346);
nand U2454 (N_2454,N_2363,N_2366);
or U2455 (N_2455,N_2385,N_2377);
nand U2456 (N_2456,N_2342,N_2371);
nand U2457 (N_2457,N_2378,N_2353);
or U2458 (N_2458,N_2373,N_2383);
or U2459 (N_2459,N_2394,N_2348);
and U2460 (N_2460,N_2445,N_2416);
nor U2461 (N_2461,N_2429,N_2418);
nand U2462 (N_2462,N_2417,N_2442);
or U2463 (N_2463,N_2421,N_2403);
or U2464 (N_2464,N_2407,N_2449);
or U2465 (N_2465,N_2404,N_2406);
or U2466 (N_2466,N_2453,N_2440);
and U2467 (N_2467,N_2424,N_2435);
and U2468 (N_2468,N_2451,N_2413);
nor U2469 (N_2469,N_2428,N_2427);
xnor U2470 (N_2470,N_2405,N_2452);
nor U2471 (N_2471,N_2438,N_2409);
or U2472 (N_2472,N_2426,N_2447);
xnor U2473 (N_2473,N_2411,N_2400);
and U2474 (N_2474,N_2410,N_2457);
xnor U2475 (N_2475,N_2408,N_2455);
or U2476 (N_2476,N_2419,N_2439);
and U2477 (N_2477,N_2437,N_2448);
or U2478 (N_2478,N_2450,N_2459);
nor U2479 (N_2479,N_2454,N_2431);
or U2480 (N_2480,N_2422,N_2441);
or U2481 (N_2481,N_2444,N_2432);
nor U2482 (N_2482,N_2430,N_2420);
nand U2483 (N_2483,N_2434,N_2414);
and U2484 (N_2484,N_2436,N_2433);
nand U2485 (N_2485,N_2412,N_2458);
and U2486 (N_2486,N_2415,N_2456);
nand U2487 (N_2487,N_2402,N_2446);
and U2488 (N_2488,N_2401,N_2423);
and U2489 (N_2489,N_2425,N_2443);
or U2490 (N_2490,N_2425,N_2451);
and U2491 (N_2491,N_2414,N_2403);
nor U2492 (N_2492,N_2424,N_2402);
and U2493 (N_2493,N_2417,N_2441);
and U2494 (N_2494,N_2412,N_2408);
nor U2495 (N_2495,N_2403,N_2426);
nand U2496 (N_2496,N_2449,N_2401);
nand U2497 (N_2497,N_2401,N_2443);
or U2498 (N_2498,N_2419,N_2441);
and U2499 (N_2499,N_2455,N_2404);
nor U2500 (N_2500,N_2437,N_2435);
and U2501 (N_2501,N_2429,N_2415);
nor U2502 (N_2502,N_2402,N_2407);
or U2503 (N_2503,N_2413,N_2414);
xor U2504 (N_2504,N_2411,N_2440);
or U2505 (N_2505,N_2435,N_2436);
and U2506 (N_2506,N_2457,N_2436);
nor U2507 (N_2507,N_2422,N_2431);
nand U2508 (N_2508,N_2402,N_2458);
or U2509 (N_2509,N_2405,N_2449);
nor U2510 (N_2510,N_2452,N_2441);
or U2511 (N_2511,N_2431,N_2450);
nor U2512 (N_2512,N_2420,N_2438);
xnor U2513 (N_2513,N_2427,N_2447);
nor U2514 (N_2514,N_2432,N_2429);
or U2515 (N_2515,N_2415,N_2451);
nand U2516 (N_2516,N_2412,N_2413);
or U2517 (N_2517,N_2442,N_2455);
or U2518 (N_2518,N_2400,N_2427);
xor U2519 (N_2519,N_2459,N_2457);
or U2520 (N_2520,N_2515,N_2505);
or U2521 (N_2521,N_2483,N_2461);
and U2522 (N_2522,N_2482,N_2484);
nand U2523 (N_2523,N_2480,N_2472);
nand U2524 (N_2524,N_2493,N_2491);
xnor U2525 (N_2525,N_2466,N_2502);
or U2526 (N_2526,N_2467,N_2516);
nor U2527 (N_2527,N_2485,N_2500);
xor U2528 (N_2528,N_2497,N_2481);
nand U2529 (N_2529,N_2465,N_2492);
or U2530 (N_2530,N_2518,N_2486);
or U2531 (N_2531,N_2499,N_2508);
nand U2532 (N_2532,N_2474,N_2471);
nor U2533 (N_2533,N_2510,N_2460);
nand U2534 (N_2534,N_2479,N_2477);
nor U2535 (N_2535,N_2490,N_2495);
nand U2536 (N_2536,N_2487,N_2462);
nor U2537 (N_2537,N_2517,N_2498);
nor U2538 (N_2538,N_2506,N_2470);
nor U2539 (N_2539,N_2501,N_2489);
and U2540 (N_2540,N_2504,N_2478);
nand U2541 (N_2541,N_2473,N_2503);
and U2542 (N_2542,N_2494,N_2464);
nor U2543 (N_2543,N_2514,N_2469);
and U2544 (N_2544,N_2511,N_2468);
and U2545 (N_2545,N_2488,N_2519);
or U2546 (N_2546,N_2463,N_2496);
or U2547 (N_2547,N_2507,N_2513);
nor U2548 (N_2548,N_2509,N_2512);
nor U2549 (N_2549,N_2475,N_2476);
nand U2550 (N_2550,N_2494,N_2506);
nor U2551 (N_2551,N_2487,N_2502);
and U2552 (N_2552,N_2500,N_2466);
and U2553 (N_2553,N_2508,N_2504);
and U2554 (N_2554,N_2500,N_2510);
or U2555 (N_2555,N_2487,N_2500);
nor U2556 (N_2556,N_2474,N_2505);
and U2557 (N_2557,N_2465,N_2477);
and U2558 (N_2558,N_2497,N_2507);
nand U2559 (N_2559,N_2495,N_2472);
xor U2560 (N_2560,N_2482,N_2469);
nand U2561 (N_2561,N_2464,N_2470);
nand U2562 (N_2562,N_2480,N_2492);
nor U2563 (N_2563,N_2508,N_2503);
nor U2564 (N_2564,N_2489,N_2490);
or U2565 (N_2565,N_2497,N_2487);
and U2566 (N_2566,N_2478,N_2515);
nor U2567 (N_2567,N_2469,N_2499);
xnor U2568 (N_2568,N_2460,N_2466);
xnor U2569 (N_2569,N_2488,N_2473);
and U2570 (N_2570,N_2494,N_2498);
nand U2571 (N_2571,N_2467,N_2469);
nand U2572 (N_2572,N_2474,N_2508);
nor U2573 (N_2573,N_2488,N_2470);
nor U2574 (N_2574,N_2517,N_2510);
or U2575 (N_2575,N_2474,N_2469);
and U2576 (N_2576,N_2484,N_2469);
or U2577 (N_2577,N_2490,N_2463);
nor U2578 (N_2578,N_2499,N_2470);
and U2579 (N_2579,N_2481,N_2515);
xnor U2580 (N_2580,N_2546,N_2554);
or U2581 (N_2581,N_2532,N_2550);
or U2582 (N_2582,N_2574,N_2570);
xor U2583 (N_2583,N_2568,N_2544);
nand U2584 (N_2584,N_2522,N_2576);
xor U2585 (N_2585,N_2547,N_2565);
nor U2586 (N_2586,N_2560,N_2564);
nand U2587 (N_2587,N_2555,N_2538);
or U2588 (N_2588,N_2575,N_2531);
or U2589 (N_2589,N_2523,N_2571);
nand U2590 (N_2590,N_2542,N_2557);
xor U2591 (N_2591,N_2573,N_2559);
and U2592 (N_2592,N_2553,N_2579);
or U2593 (N_2593,N_2543,N_2540);
or U2594 (N_2594,N_2562,N_2537);
nand U2595 (N_2595,N_2525,N_2561);
or U2596 (N_2596,N_2527,N_2526);
nor U2597 (N_2597,N_2548,N_2578);
nor U2598 (N_2598,N_2566,N_2539);
and U2599 (N_2599,N_2558,N_2545);
nand U2600 (N_2600,N_2563,N_2572);
nor U2601 (N_2601,N_2524,N_2521);
nand U2602 (N_2602,N_2528,N_2533);
and U2603 (N_2603,N_2569,N_2552);
xor U2604 (N_2604,N_2551,N_2535);
nand U2605 (N_2605,N_2577,N_2549);
nand U2606 (N_2606,N_2530,N_2529);
or U2607 (N_2607,N_2534,N_2536);
nor U2608 (N_2608,N_2520,N_2556);
nor U2609 (N_2609,N_2541,N_2567);
or U2610 (N_2610,N_2548,N_2557);
or U2611 (N_2611,N_2559,N_2535);
nor U2612 (N_2612,N_2530,N_2574);
nand U2613 (N_2613,N_2562,N_2577);
nor U2614 (N_2614,N_2540,N_2571);
xnor U2615 (N_2615,N_2546,N_2526);
or U2616 (N_2616,N_2525,N_2575);
and U2617 (N_2617,N_2529,N_2534);
and U2618 (N_2618,N_2569,N_2572);
nand U2619 (N_2619,N_2567,N_2526);
and U2620 (N_2620,N_2575,N_2564);
nand U2621 (N_2621,N_2536,N_2533);
or U2622 (N_2622,N_2566,N_2530);
xor U2623 (N_2623,N_2562,N_2559);
or U2624 (N_2624,N_2565,N_2527);
and U2625 (N_2625,N_2521,N_2573);
nand U2626 (N_2626,N_2538,N_2545);
nor U2627 (N_2627,N_2575,N_2540);
nand U2628 (N_2628,N_2558,N_2548);
nand U2629 (N_2629,N_2544,N_2520);
nand U2630 (N_2630,N_2572,N_2559);
nand U2631 (N_2631,N_2529,N_2541);
and U2632 (N_2632,N_2526,N_2539);
and U2633 (N_2633,N_2558,N_2524);
and U2634 (N_2634,N_2554,N_2533);
nand U2635 (N_2635,N_2539,N_2538);
or U2636 (N_2636,N_2549,N_2536);
or U2637 (N_2637,N_2555,N_2567);
xor U2638 (N_2638,N_2553,N_2535);
nand U2639 (N_2639,N_2536,N_2578);
nand U2640 (N_2640,N_2596,N_2623);
or U2641 (N_2641,N_2601,N_2627);
nand U2642 (N_2642,N_2597,N_2604);
xnor U2643 (N_2643,N_2606,N_2588);
xor U2644 (N_2644,N_2624,N_2595);
nor U2645 (N_2645,N_2584,N_2639);
and U2646 (N_2646,N_2635,N_2593);
and U2647 (N_2647,N_2581,N_2629);
nand U2648 (N_2648,N_2617,N_2599);
and U2649 (N_2649,N_2620,N_2614);
or U2650 (N_2650,N_2636,N_2628);
or U2651 (N_2651,N_2602,N_2630);
or U2652 (N_2652,N_2592,N_2598);
nand U2653 (N_2653,N_2587,N_2608);
nor U2654 (N_2654,N_2582,N_2600);
nand U2655 (N_2655,N_2619,N_2633);
or U2656 (N_2656,N_2638,N_2591);
or U2657 (N_2657,N_2621,N_2610);
and U2658 (N_2658,N_2605,N_2594);
nor U2659 (N_2659,N_2616,N_2607);
or U2660 (N_2660,N_2613,N_2589);
nand U2661 (N_2661,N_2632,N_2631);
xnor U2662 (N_2662,N_2625,N_2612);
nand U2663 (N_2663,N_2590,N_2615);
and U2664 (N_2664,N_2626,N_2583);
nor U2665 (N_2665,N_2634,N_2611);
and U2666 (N_2666,N_2603,N_2637);
and U2667 (N_2667,N_2618,N_2609);
nand U2668 (N_2668,N_2622,N_2586);
nand U2669 (N_2669,N_2580,N_2585);
or U2670 (N_2670,N_2592,N_2614);
nor U2671 (N_2671,N_2619,N_2626);
xor U2672 (N_2672,N_2585,N_2603);
and U2673 (N_2673,N_2619,N_2582);
nor U2674 (N_2674,N_2608,N_2595);
or U2675 (N_2675,N_2622,N_2636);
and U2676 (N_2676,N_2585,N_2632);
nand U2677 (N_2677,N_2591,N_2623);
or U2678 (N_2678,N_2634,N_2594);
and U2679 (N_2679,N_2617,N_2612);
or U2680 (N_2680,N_2594,N_2593);
and U2681 (N_2681,N_2629,N_2613);
or U2682 (N_2682,N_2602,N_2597);
nand U2683 (N_2683,N_2607,N_2608);
or U2684 (N_2684,N_2625,N_2604);
or U2685 (N_2685,N_2621,N_2598);
and U2686 (N_2686,N_2623,N_2585);
xor U2687 (N_2687,N_2638,N_2583);
or U2688 (N_2688,N_2636,N_2614);
nand U2689 (N_2689,N_2584,N_2617);
or U2690 (N_2690,N_2619,N_2597);
nand U2691 (N_2691,N_2639,N_2598);
or U2692 (N_2692,N_2633,N_2626);
and U2693 (N_2693,N_2611,N_2614);
or U2694 (N_2694,N_2608,N_2582);
and U2695 (N_2695,N_2605,N_2634);
nor U2696 (N_2696,N_2626,N_2599);
or U2697 (N_2697,N_2608,N_2614);
nand U2698 (N_2698,N_2620,N_2582);
nand U2699 (N_2699,N_2584,N_2583);
xnor U2700 (N_2700,N_2662,N_2642);
and U2701 (N_2701,N_2690,N_2671);
or U2702 (N_2702,N_2664,N_2655);
or U2703 (N_2703,N_2675,N_2692);
nand U2704 (N_2704,N_2647,N_2640);
or U2705 (N_2705,N_2666,N_2698);
nor U2706 (N_2706,N_2650,N_2689);
or U2707 (N_2707,N_2663,N_2697);
nand U2708 (N_2708,N_2676,N_2688);
nor U2709 (N_2709,N_2659,N_2699);
and U2710 (N_2710,N_2667,N_2649);
nor U2711 (N_2711,N_2686,N_2678);
or U2712 (N_2712,N_2682,N_2661);
nand U2713 (N_2713,N_2693,N_2696);
or U2714 (N_2714,N_2652,N_2643);
and U2715 (N_2715,N_2669,N_2660);
nand U2716 (N_2716,N_2694,N_2644);
xnor U2717 (N_2717,N_2673,N_2654);
nor U2718 (N_2718,N_2681,N_2668);
nand U2719 (N_2719,N_2685,N_2653);
nor U2720 (N_2720,N_2657,N_2677);
and U2721 (N_2721,N_2674,N_2645);
or U2722 (N_2722,N_2641,N_2687);
nand U2723 (N_2723,N_2651,N_2646);
or U2724 (N_2724,N_2680,N_2683);
and U2725 (N_2725,N_2658,N_2679);
xor U2726 (N_2726,N_2648,N_2684);
or U2727 (N_2727,N_2665,N_2695);
or U2728 (N_2728,N_2691,N_2656);
nand U2729 (N_2729,N_2670,N_2672);
nand U2730 (N_2730,N_2672,N_2690);
nand U2731 (N_2731,N_2658,N_2650);
and U2732 (N_2732,N_2690,N_2691);
nor U2733 (N_2733,N_2648,N_2669);
nor U2734 (N_2734,N_2673,N_2640);
xnor U2735 (N_2735,N_2690,N_2681);
and U2736 (N_2736,N_2694,N_2670);
and U2737 (N_2737,N_2696,N_2664);
and U2738 (N_2738,N_2654,N_2686);
or U2739 (N_2739,N_2678,N_2657);
or U2740 (N_2740,N_2682,N_2683);
and U2741 (N_2741,N_2680,N_2652);
nand U2742 (N_2742,N_2640,N_2664);
nor U2743 (N_2743,N_2668,N_2655);
nor U2744 (N_2744,N_2657,N_2644);
and U2745 (N_2745,N_2662,N_2684);
nor U2746 (N_2746,N_2669,N_2646);
or U2747 (N_2747,N_2642,N_2644);
and U2748 (N_2748,N_2654,N_2650);
and U2749 (N_2749,N_2696,N_2683);
and U2750 (N_2750,N_2679,N_2642);
nor U2751 (N_2751,N_2645,N_2655);
and U2752 (N_2752,N_2675,N_2662);
or U2753 (N_2753,N_2671,N_2675);
and U2754 (N_2754,N_2656,N_2672);
nand U2755 (N_2755,N_2654,N_2670);
and U2756 (N_2756,N_2661,N_2695);
nor U2757 (N_2757,N_2694,N_2663);
nor U2758 (N_2758,N_2692,N_2684);
nand U2759 (N_2759,N_2653,N_2661);
nor U2760 (N_2760,N_2747,N_2725);
nor U2761 (N_2761,N_2742,N_2739);
or U2762 (N_2762,N_2741,N_2757);
nand U2763 (N_2763,N_2714,N_2728);
nor U2764 (N_2764,N_2745,N_2730);
or U2765 (N_2765,N_2749,N_2746);
nand U2766 (N_2766,N_2709,N_2744);
xnor U2767 (N_2767,N_2707,N_2721);
nand U2768 (N_2768,N_2731,N_2723);
xnor U2769 (N_2769,N_2722,N_2758);
nor U2770 (N_2770,N_2753,N_2755);
or U2771 (N_2771,N_2743,N_2759);
or U2772 (N_2772,N_2754,N_2718);
nand U2773 (N_2773,N_2748,N_2735);
nor U2774 (N_2774,N_2720,N_2713);
and U2775 (N_2775,N_2703,N_2705);
nand U2776 (N_2776,N_2719,N_2700);
or U2777 (N_2777,N_2717,N_2716);
or U2778 (N_2778,N_2701,N_2710);
or U2779 (N_2779,N_2724,N_2750);
and U2780 (N_2780,N_2738,N_2751);
nor U2781 (N_2781,N_2740,N_2736);
and U2782 (N_2782,N_2715,N_2756);
nor U2783 (N_2783,N_2704,N_2711);
and U2784 (N_2784,N_2702,N_2737);
xnor U2785 (N_2785,N_2752,N_2734);
or U2786 (N_2786,N_2732,N_2712);
nand U2787 (N_2787,N_2727,N_2729);
and U2788 (N_2788,N_2726,N_2733);
nor U2789 (N_2789,N_2706,N_2708);
and U2790 (N_2790,N_2726,N_2743);
nor U2791 (N_2791,N_2709,N_2749);
or U2792 (N_2792,N_2718,N_2729);
or U2793 (N_2793,N_2750,N_2759);
xnor U2794 (N_2794,N_2744,N_2719);
and U2795 (N_2795,N_2716,N_2711);
nand U2796 (N_2796,N_2749,N_2719);
nand U2797 (N_2797,N_2704,N_2751);
nor U2798 (N_2798,N_2722,N_2753);
or U2799 (N_2799,N_2742,N_2710);
and U2800 (N_2800,N_2701,N_2739);
or U2801 (N_2801,N_2717,N_2730);
nand U2802 (N_2802,N_2732,N_2730);
and U2803 (N_2803,N_2721,N_2704);
nor U2804 (N_2804,N_2759,N_2721);
and U2805 (N_2805,N_2743,N_2735);
and U2806 (N_2806,N_2746,N_2717);
or U2807 (N_2807,N_2741,N_2712);
nand U2808 (N_2808,N_2722,N_2703);
xnor U2809 (N_2809,N_2705,N_2711);
or U2810 (N_2810,N_2726,N_2725);
nand U2811 (N_2811,N_2706,N_2755);
and U2812 (N_2812,N_2718,N_2714);
nor U2813 (N_2813,N_2709,N_2726);
nor U2814 (N_2814,N_2714,N_2724);
or U2815 (N_2815,N_2737,N_2713);
xor U2816 (N_2816,N_2730,N_2751);
and U2817 (N_2817,N_2739,N_2738);
nor U2818 (N_2818,N_2746,N_2745);
nand U2819 (N_2819,N_2700,N_2741);
and U2820 (N_2820,N_2772,N_2787);
nand U2821 (N_2821,N_2763,N_2802);
and U2822 (N_2822,N_2771,N_2762);
xor U2823 (N_2823,N_2806,N_2798);
nor U2824 (N_2824,N_2816,N_2810);
nand U2825 (N_2825,N_2797,N_2818);
or U2826 (N_2826,N_2807,N_2800);
and U2827 (N_2827,N_2788,N_2775);
or U2828 (N_2828,N_2781,N_2811);
nand U2829 (N_2829,N_2777,N_2779);
or U2830 (N_2830,N_2782,N_2805);
or U2831 (N_2831,N_2813,N_2814);
nor U2832 (N_2832,N_2794,N_2792);
xor U2833 (N_2833,N_2761,N_2796);
xor U2834 (N_2834,N_2767,N_2790);
xnor U2835 (N_2835,N_2785,N_2799);
nand U2836 (N_2836,N_2786,N_2773);
or U2837 (N_2837,N_2768,N_2801);
or U2838 (N_2838,N_2795,N_2760);
and U2839 (N_2839,N_2809,N_2778);
and U2840 (N_2840,N_2770,N_2812);
nor U2841 (N_2841,N_2803,N_2783);
nand U2842 (N_2842,N_2776,N_2793);
nor U2843 (N_2843,N_2791,N_2780);
nand U2844 (N_2844,N_2804,N_2764);
nor U2845 (N_2845,N_2817,N_2815);
nor U2846 (N_2846,N_2789,N_2766);
xnor U2847 (N_2847,N_2808,N_2765);
nor U2848 (N_2848,N_2819,N_2774);
or U2849 (N_2849,N_2784,N_2769);
nand U2850 (N_2850,N_2774,N_2797);
xnor U2851 (N_2851,N_2799,N_2818);
or U2852 (N_2852,N_2811,N_2800);
nand U2853 (N_2853,N_2789,N_2774);
and U2854 (N_2854,N_2797,N_2781);
nand U2855 (N_2855,N_2787,N_2793);
or U2856 (N_2856,N_2763,N_2773);
or U2857 (N_2857,N_2789,N_2777);
and U2858 (N_2858,N_2807,N_2784);
or U2859 (N_2859,N_2768,N_2811);
or U2860 (N_2860,N_2769,N_2814);
or U2861 (N_2861,N_2763,N_2769);
and U2862 (N_2862,N_2764,N_2779);
xor U2863 (N_2863,N_2763,N_2783);
xor U2864 (N_2864,N_2763,N_2813);
xnor U2865 (N_2865,N_2812,N_2817);
nand U2866 (N_2866,N_2783,N_2817);
or U2867 (N_2867,N_2797,N_2785);
or U2868 (N_2868,N_2812,N_2763);
nand U2869 (N_2869,N_2778,N_2818);
nor U2870 (N_2870,N_2815,N_2770);
or U2871 (N_2871,N_2812,N_2811);
nor U2872 (N_2872,N_2793,N_2765);
xor U2873 (N_2873,N_2803,N_2800);
nand U2874 (N_2874,N_2819,N_2814);
or U2875 (N_2875,N_2783,N_2760);
nand U2876 (N_2876,N_2814,N_2776);
nand U2877 (N_2877,N_2779,N_2762);
or U2878 (N_2878,N_2815,N_2786);
or U2879 (N_2879,N_2760,N_2794);
nand U2880 (N_2880,N_2854,N_2828);
or U2881 (N_2881,N_2852,N_2853);
and U2882 (N_2882,N_2842,N_2872);
nor U2883 (N_2883,N_2825,N_2820);
or U2884 (N_2884,N_2839,N_2836);
nand U2885 (N_2885,N_2849,N_2840);
xor U2886 (N_2886,N_2847,N_2869);
nor U2887 (N_2887,N_2866,N_2870);
nor U2888 (N_2888,N_2832,N_2843);
xnor U2889 (N_2889,N_2837,N_2827);
nand U2890 (N_2890,N_2857,N_2833);
nor U2891 (N_2891,N_2848,N_2878);
or U2892 (N_2892,N_2861,N_2865);
nor U2893 (N_2893,N_2879,N_2844);
or U2894 (N_2894,N_2846,N_2834);
nand U2895 (N_2895,N_2821,N_2874);
or U2896 (N_2896,N_2835,N_2875);
and U2897 (N_2897,N_2855,N_2860);
nor U2898 (N_2898,N_2851,N_2877);
nor U2899 (N_2899,N_2867,N_2826);
nor U2900 (N_2900,N_2822,N_2859);
nand U2901 (N_2901,N_2830,N_2858);
and U2902 (N_2902,N_2841,N_2823);
nand U2903 (N_2903,N_2876,N_2862);
or U2904 (N_2904,N_2873,N_2838);
nor U2905 (N_2905,N_2824,N_2863);
or U2906 (N_2906,N_2864,N_2829);
and U2907 (N_2907,N_2845,N_2831);
nor U2908 (N_2908,N_2856,N_2850);
or U2909 (N_2909,N_2868,N_2871);
or U2910 (N_2910,N_2837,N_2845);
and U2911 (N_2911,N_2844,N_2851);
and U2912 (N_2912,N_2850,N_2863);
nor U2913 (N_2913,N_2820,N_2869);
and U2914 (N_2914,N_2841,N_2826);
and U2915 (N_2915,N_2839,N_2847);
and U2916 (N_2916,N_2843,N_2836);
nand U2917 (N_2917,N_2852,N_2854);
and U2918 (N_2918,N_2820,N_2839);
nor U2919 (N_2919,N_2872,N_2855);
and U2920 (N_2920,N_2866,N_2869);
nand U2921 (N_2921,N_2873,N_2829);
or U2922 (N_2922,N_2830,N_2851);
nor U2923 (N_2923,N_2821,N_2860);
nor U2924 (N_2924,N_2872,N_2852);
or U2925 (N_2925,N_2869,N_2834);
nand U2926 (N_2926,N_2878,N_2857);
nor U2927 (N_2927,N_2836,N_2859);
and U2928 (N_2928,N_2850,N_2878);
and U2929 (N_2929,N_2838,N_2876);
or U2930 (N_2930,N_2867,N_2870);
nor U2931 (N_2931,N_2865,N_2845);
or U2932 (N_2932,N_2840,N_2834);
or U2933 (N_2933,N_2858,N_2869);
and U2934 (N_2934,N_2860,N_2856);
nand U2935 (N_2935,N_2878,N_2869);
nor U2936 (N_2936,N_2863,N_2879);
and U2937 (N_2937,N_2858,N_2852);
nand U2938 (N_2938,N_2855,N_2865);
nand U2939 (N_2939,N_2821,N_2854);
and U2940 (N_2940,N_2912,N_2934);
and U2941 (N_2941,N_2906,N_2932);
nand U2942 (N_2942,N_2889,N_2938);
and U2943 (N_2943,N_2930,N_2902);
xor U2944 (N_2944,N_2898,N_2933);
or U2945 (N_2945,N_2928,N_2909);
nand U2946 (N_2946,N_2913,N_2935);
or U2947 (N_2947,N_2910,N_2900);
nand U2948 (N_2948,N_2911,N_2881);
nor U2949 (N_2949,N_2919,N_2890);
and U2950 (N_2950,N_2884,N_2915);
nand U2951 (N_2951,N_2926,N_2887);
or U2952 (N_2952,N_2882,N_2922);
or U2953 (N_2953,N_2885,N_2916);
xnor U2954 (N_2954,N_2892,N_2937);
nand U2955 (N_2955,N_2891,N_2929);
nand U2956 (N_2956,N_2917,N_2936);
nand U2957 (N_2957,N_2907,N_2895);
xor U2958 (N_2958,N_2893,N_2880);
or U2959 (N_2959,N_2899,N_2894);
or U2960 (N_2960,N_2931,N_2883);
nand U2961 (N_2961,N_2923,N_2914);
xnor U2962 (N_2962,N_2918,N_2927);
nand U2963 (N_2963,N_2896,N_2924);
or U2964 (N_2964,N_2888,N_2908);
or U2965 (N_2965,N_2886,N_2901);
or U2966 (N_2966,N_2925,N_2905);
nor U2967 (N_2967,N_2897,N_2920);
and U2968 (N_2968,N_2921,N_2903);
nor U2969 (N_2969,N_2904,N_2939);
nor U2970 (N_2970,N_2916,N_2938);
and U2971 (N_2971,N_2935,N_2922);
and U2972 (N_2972,N_2921,N_2882);
nor U2973 (N_2973,N_2934,N_2905);
nand U2974 (N_2974,N_2921,N_2918);
and U2975 (N_2975,N_2918,N_2889);
nor U2976 (N_2976,N_2899,N_2927);
nor U2977 (N_2977,N_2911,N_2934);
or U2978 (N_2978,N_2890,N_2917);
and U2979 (N_2979,N_2926,N_2934);
nand U2980 (N_2980,N_2925,N_2921);
or U2981 (N_2981,N_2923,N_2907);
or U2982 (N_2982,N_2913,N_2892);
nand U2983 (N_2983,N_2910,N_2887);
nand U2984 (N_2984,N_2892,N_2901);
and U2985 (N_2985,N_2916,N_2939);
and U2986 (N_2986,N_2922,N_2894);
or U2987 (N_2987,N_2902,N_2882);
and U2988 (N_2988,N_2913,N_2923);
or U2989 (N_2989,N_2915,N_2924);
and U2990 (N_2990,N_2922,N_2905);
or U2991 (N_2991,N_2937,N_2926);
nand U2992 (N_2992,N_2912,N_2899);
xnor U2993 (N_2993,N_2921,N_2915);
and U2994 (N_2994,N_2906,N_2918);
nand U2995 (N_2995,N_2937,N_2882);
and U2996 (N_2996,N_2919,N_2889);
or U2997 (N_2997,N_2891,N_2934);
nor U2998 (N_2998,N_2891,N_2928);
nor U2999 (N_2999,N_2924,N_2936);
nor UO_0 (O_0,N_2971,N_2960);
nand UO_1 (O_1,N_2955,N_2943);
nand UO_2 (O_2,N_2964,N_2980);
xor UO_3 (O_3,N_2976,N_2963);
and UO_4 (O_4,N_2958,N_2979);
nand UO_5 (O_5,N_2949,N_2941);
and UO_6 (O_6,N_2967,N_2981);
or UO_7 (O_7,N_2997,N_2988);
or UO_8 (O_8,N_2942,N_2951);
nand UO_9 (O_9,N_2985,N_2998);
nand UO_10 (O_10,N_2962,N_2992);
and UO_11 (O_11,N_2982,N_2950);
nand UO_12 (O_12,N_2970,N_2975);
nor UO_13 (O_13,N_2953,N_2991);
nor UO_14 (O_14,N_2968,N_2996);
and UO_15 (O_15,N_2974,N_2977);
or UO_16 (O_16,N_2994,N_2947);
nand UO_17 (O_17,N_2965,N_2940);
and UO_18 (O_18,N_2952,N_2948);
nand UO_19 (O_19,N_2978,N_2954);
xnor UO_20 (O_20,N_2986,N_2959);
or UO_21 (O_21,N_2944,N_2972);
or UO_22 (O_22,N_2993,N_2946);
or UO_23 (O_23,N_2956,N_2945);
nor UO_24 (O_24,N_2966,N_2973);
nor UO_25 (O_25,N_2999,N_2957);
and UO_26 (O_26,N_2989,N_2969);
nand UO_27 (O_27,N_2987,N_2983);
nand UO_28 (O_28,N_2961,N_2984);
or UO_29 (O_29,N_2990,N_2995);
nand UO_30 (O_30,N_2941,N_2969);
or UO_31 (O_31,N_2969,N_2988);
or UO_32 (O_32,N_2972,N_2966);
nor UO_33 (O_33,N_2988,N_2951);
nand UO_34 (O_34,N_2978,N_2948);
xnor UO_35 (O_35,N_2971,N_2964);
xnor UO_36 (O_36,N_2959,N_2960);
and UO_37 (O_37,N_2983,N_2974);
nand UO_38 (O_38,N_2970,N_2951);
xor UO_39 (O_39,N_2943,N_2997);
nand UO_40 (O_40,N_2996,N_2971);
or UO_41 (O_41,N_2960,N_2991);
or UO_42 (O_42,N_2964,N_2990);
or UO_43 (O_43,N_2954,N_2977);
or UO_44 (O_44,N_2943,N_2948);
and UO_45 (O_45,N_2967,N_2996);
or UO_46 (O_46,N_2984,N_2957);
xnor UO_47 (O_47,N_2992,N_2979);
nor UO_48 (O_48,N_2949,N_2979);
or UO_49 (O_49,N_2947,N_2948);
nor UO_50 (O_50,N_2986,N_2984);
xnor UO_51 (O_51,N_2979,N_2944);
nand UO_52 (O_52,N_2979,N_2980);
or UO_53 (O_53,N_2988,N_2986);
nand UO_54 (O_54,N_2974,N_2997);
nand UO_55 (O_55,N_2950,N_2989);
and UO_56 (O_56,N_2991,N_2961);
and UO_57 (O_57,N_2981,N_2959);
xor UO_58 (O_58,N_2963,N_2949);
nor UO_59 (O_59,N_2954,N_2942);
xor UO_60 (O_60,N_2964,N_2983);
or UO_61 (O_61,N_2961,N_2952);
nor UO_62 (O_62,N_2997,N_2945);
and UO_63 (O_63,N_2968,N_2962);
nand UO_64 (O_64,N_2968,N_2951);
and UO_65 (O_65,N_2961,N_2965);
nor UO_66 (O_66,N_2953,N_2965);
xnor UO_67 (O_67,N_2986,N_2997);
nand UO_68 (O_68,N_2962,N_2957);
xor UO_69 (O_69,N_2952,N_2943);
nand UO_70 (O_70,N_2955,N_2944);
nor UO_71 (O_71,N_2967,N_2977);
nor UO_72 (O_72,N_2986,N_2953);
and UO_73 (O_73,N_2946,N_2991);
nand UO_74 (O_74,N_2946,N_2974);
nand UO_75 (O_75,N_2961,N_2954);
and UO_76 (O_76,N_2973,N_2971);
nor UO_77 (O_77,N_2979,N_2960);
nor UO_78 (O_78,N_2959,N_2994);
and UO_79 (O_79,N_2980,N_2950);
or UO_80 (O_80,N_2978,N_2989);
nor UO_81 (O_81,N_2970,N_2971);
nand UO_82 (O_82,N_2978,N_2961);
or UO_83 (O_83,N_2965,N_2956);
nor UO_84 (O_84,N_2998,N_2980);
nand UO_85 (O_85,N_2967,N_2961);
nand UO_86 (O_86,N_2990,N_2957);
nand UO_87 (O_87,N_2956,N_2976);
nor UO_88 (O_88,N_2957,N_2996);
or UO_89 (O_89,N_2999,N_2948);
nand UO_90 (O_90,N_2948,N_2997);
or UO_91 (O_91,N_2992,N_2943);
and UO_92 (O_92,N_2979,N_2948);
or UO_93 (O_93,N_2942,N_2953);
and UO_94 (O_94,N_2943,N_2961);
nand UO_95 (O_95,N_2956,N_2980);
and UO_96 (O_96,N_2972,N_2949);
nand UO_97 (O_97,N_2981,N_2969);
or UO_98 (O_98,N_2981,N_2979);
xor UO_99 (O_99,N_2954,N_2988);
and UO_100 (O_100,N_2962,N_2963);
nor UO_101 (O_101,N_2965,N_2946);
or UO_102 (O_102,N_2963,N_2985);
nand UO_103 (O_103,N_2989,N_2963);
nor UO_104 (O_104,N_2986,N_2949);
nand UO_105 (O_105,N_2998,N_2953);
and UO_106 (O_106,N_2957,N_2989);
or UO_107 (O_107,N_2944,N_2986);
and UO_108 (O_108,N_2984,N_2944);
xnor UO_109 (O_109,N_2949,N_2946);
or UO_110 (O_110,N_2995,N_2948);
xor UO_111 (O_111,N_2965,N_2973);
nor UO_112 (O_112,N_2950,N_2966);
or UO_113 (O_113,N_2953,N_2944);
nand UO_114 (O_114,N_2997,N_2959);
nor UO_115 (O_115,N_2974,N_2944);
or UO_116 (O_116,N_2955,N_2946);
nand UO_117 (O_117,N_2959,N_2940);
nor UO_118 (O_118,N_2992,N_2977);
and UO_119 (O_119,N_2992,N_2983);
nor UO_120 (O_120,N_2951,N_2999);
nand UO_121 (O_121,N_2982,N_2983);
xnor UO_122 (O_122,N_2962,N_2949);
and UO_123 (O_123,N_2960,N_2993);
and UO_124 (O_124,N_2961,N_2997);
or UO_125 (O_125,N_2966,N_2984);
and UO_126 (O_126,N_2968,N_2960);
or UO_127 (O_127,N_2999,N_2986);
or UO_128 (O_128,N_2995,N_2989);
nor UO_129 (O_129,N_2943,N_2945);
or UO_130 (O_130,N_2989,N_2961);
nand UO_131 (O_131,N_2973,N_2978);
nor UO_132 (O_132,N_2985,N_2946);
xnor UO_133 (O_133,N_2947,N_2988);
nand UO_134 (O_134,N_2993,N_2940);
nand UO_135 (O_135,N_2986,N_2964);
and UO_136 (O_136,N_2969,N_2986);
nand UO_137 (O_137,N_2944,N_2999);
xnor UO_138 (O_138,N_2960,N_2998);
or UO_139 (O_139,N_2991,N_2947);
or UO_140 (O_140,N_2959,N_2943);
nor UO_141 (O_141,N_2950,N_2994);
nand UO_142 (O_142,N_2989,N_2955);
xnor UO_143 (O_143,N_2986,N_2985);
or UO_144 (O_144,N_2956,N_2949);
nor UO_145 (O_145,N_2990,N_2987);
or UO_146 (O_146,N_2980,N_2997);
nor UO_147 (O_147,N_2987,N_2962);
nor UO_148 (O_148,N_2947,N_2995);
or UO_149 (O_149,N_2984,N_2992);
or UO_150 (O_150,N_2982,N_2973);
nor UO_151 (O_151,N_2985,N_2995);
or UO_152 (O_152,N_2965,N_2993);
nor UO_153 (O_153,N_2947,N_2980);
and UO_154 (O_154,N_2944,N_2943);
nand UO_155 (O_155,N_2970,N_2985);
and UO_156 (O_156,N_2980,N_2977);
or UO_157 (O_157,N_2946,N_2976);
or UO_158 (O_158,N_2968,N_2946);
or UO_159 (O_159,N_2964,N_2957);
nand UO_160 (O_160,N_2958,N_2984);
and UO_161 (O_161,N_2942,N_2940);
nor UO_162 (O_162,N_2996,N_2990);
and UO_163 (O_163,N_2988,N_2983);
and UO_164 (O_164,N_2979,N_2974);
nand UO_165 (O_165,N_2941,N_2971);
nor UO_166 (O_166,N_2998,N_2959);
or UO_167 (O_167,N_2957,N_2949);
nor UO_168 (O_168,N_2971,N_2944);
and UO_169 (O_169,N_2966,N_2987);
nor UO_170 (O_170,N_2960,N_2942);
xnor UO_171 (O_171,N_2976,N_2978);
nand UO_172 (O_172,N_2990,N_2954);
or UO_173 (O_173,N_2966,N_2953);
or UO_174 (O_174,N_2964,N_2972);
and UO_175 (O_175,N_2972,N_2991);
nor UO_176 (O_176,N_2951,N_2987);
or UO_177 (O_177,N_2980,N_2986);
nand UO_178 (O_178,N_2945,N_2990);
or UO_179 (O_179,N_2970,N_2997);
nand UO_180 (O_180,N_2995,N_2960);
or UO_181 (O_181,N_2968,N_2987);
and UO_182 (O_182,N_2956,N_2994);
or UO_183 (O_183,N_2950,N_2965);
nor UO_184 (O_184,N_2994,N_2967);
nand UO_185 (O_185,N_2962,N_2976);
xnor UO_186 (O_186,N_2944,N_2992);
and UO_187 (O_187,N_2961,N_2983);
or UO_188 (O_188,N_2984,N_2991);
nand UO_189 (O_189,N_2950,N_2959);
nand UO_190 (O_190,N_2948,N_2967);
and UO_191 (O_191,N_2976,N_2964);
nor UO_192 (O_192,N_2965,N_2988);
nor UO_193 (O_193,N_2943,N_2976);
nor UO_194 (O_194,N_2974,N_2953);
or UO_195 (O_195,N_2982,N_2999);
or UO_196 (O_196,N_2969,N_2974);
nor UO_197 (O_197,N_2980,N_2983);
nand UO_198 (O_198,N_2959,N_2964);
nor UO_199 (O_199,N_2994,N_2943);
and UO_200 (O_200,N_2964,N_2989);
and UO_201 (O_201,N_2973,N_2987);
or UO_202 (O_202,N_2966,N_2977);
nand UO_203 (O_203,N_2962,N_2990);
nand UO_204 (O_204,N_2976,N_2970);
nand UO_205 (O_205,N_2949,N_2966);
nor UO_206 (O_206,N_2974,N_2998);
nor UO_207 (O_207,N_2985,N_2960);
nand UO_208 (O_208,N_2983,N_2944);
nor UO_209 (O_209,N_2991,N_2963);
or UO_210 (O_210,N_2952,N_2941);
nand UO_211 (O_211,N_2998,N_2996);
nand UO_212 (O_212,N_2998,N_2990);
xor UO_213 (O_213,N_2984,N_2977);
or UO_214 (O_214,N_2959,N_2949);
nor UO_215 (O_215,N_2986,N_2974);
nand UO_216 (O_216,N_2947,N_2981);
and UO_217 (O_217,N_2963,N_2946);
nor UO_218 (O_218,N_2976,N_2945);
nor UO_219 (O_219,N_2989,N_2985);
xnor UO_220 (O_220,N_2977,N_2970);
or UO_221 (O_221,N_2963,N_2966);
and UO_222 (O_222,N_2994,N_2940);
or UO_223 (O_223,N_2987,N_2960);
or UO_224 (O_224,N_2941,N_2984);
nor UO_225 (O_225,N_2953,N_2941);
xor UO_226 (O_226,N_2964,N_2988);
or UO_227 (O_227,N_2985,N_2953);
or UO_228 (O_228,N_2977,N_2945);
or UO_229 (O_229,N_2991,N_2977);
xor UO_230 (O_230,N_2976,N_2991);
or UO_231 (O_231,N_2963,N_2960);
nor UO_232 (O_232,N_2972,N_2973);
and UO_233 (O_233,N_2993,N_2964);
or UO_234 (O_234,N_2991,N_2945);
and UO_235 (O_235,N_2942,N_2994);
nor UO_236 (O_236,N_2966,N_2976);
nor UO_237 (O_237,N_2960,N_2951);
nor UO_238 (O_238,N_2955,N_2997);
nor UO_239 (O_239,N_2975,N_2986);
xor UO_240 (O_240,N_2986,N_2990);
nand UO_241 (O_241,N_2958,N_2970);
or UO_242 (O_242,N_2952,N_2993);
nor UO_243 (O_243,N_2946,N_2961);
or UO_244 (O_244,N_2964,N_2966);
and UO_245 (O_245,N_2943,N_2999);
or UO_246 (O_246,N_2983,N_2995);
nor UO_247 (O_247,N_2947,N_2970);
and UO_248 (O_248,N_2952,N_2963);
nand UO_249 (O_249,N_2995,N_2941);
or UO_250 (O_250,N_2948,N_2986);
or UO_251 (O_251,N_2989,N_2981);
and UO_252 (O_252,N_2964,N_2940);
nor UO_253 (O_253,N_2971,N_2993);
nor UO_254 (O_254,N_2954,N_2951);
and UO_255 (O_255,N_2963,N_2958);
nor UO_256 (O_256,N_2970,N_2949);
nand UO_257 (O_257,N_2968,N_2980);
or UO_258 (O_258,N_2966,N_2999);
nor UO_259 (O_259,N_2991,N_2940);
nand UO_260 (O_260,N_2952,N_2951);
nand UO_261 (O_261,N_2991,N_2982);
nor UO_262 (O_262,N_2947,N_2945);
nor UO_263 (O_263,N_2975,N_2945);
and UO_264 (O_264,N_2980,N_2990);
and UO_265 (O_265,N_2956,N_2989);
nor UO_266 (O_266,N_2956,N_2955);
xnor UO_267 (O_267,N_2979,N_2984);
xor UO_268 (O_268,N_2987,N_2993);
nand UO_269 (O_269,N_2998,N_2986);
nor UO_270 (O_270,N_2984,N_2983);
or UO_271 (O_271,N_2980,N_2943);
or UO_272 (O_272,N_2974,N_2957);
xnor UO_273 (O_273,N_2974,N_2990);
nor UO_274 (O_274,N_2977,N_2986);
nor UO_275 (O_275,N_2953,N_2999);
xnor UO_276 (O_276,N_2952,N_2982);
or UO_277 (O_277,N_2958,N_2995);
nand UO_278 (O_278,N_2965,N_2989);
or UO_279 (O_279,N_2960,N_2940);
and UO_280 (O_280,N_2963,N_2971);
and UO_281 (O_281,N_2973,N_2949);
or UO_282 (O_282,N_2960,N_2982);
nand UO_283 (O_283,N_2987,N_2996);
or UO_284 (O_284,N_2961,N_2942);
and UO_285 (O_285,N_2976,N_2947);
xnor UO_286 (O_286,N_2967,N_2986);
nor UO_287 (O_287,N_2955,N_2999);
and UO_288 (O_288,N_2982,N_2951);
nand UO_289 (O_289,N_2986,N_2972);
nor UO_290 (O_290,N_2948,N_2973);
or UO_291 (O_291,N_2969,N_2992);
nand UO_292 (O_292,N_2991,N_2957);
or UO_293 (O_293,N_2948,N_2990);
nand UO_294 (O_294,N_2968,N_2993);
and UO_295 (O_295,N_2992,N_2989);
or UO_296 (O_296,N_2990,N_2976);
and UO_297 (O_297,N_2971,N_2942);
nor UO_298 (O_298,N_2943,N_2987);
and UO_299 (O_299,N_2997,N_2995);
and UO_300 (O_300,N_2966,N_2982);
and UO_301 (O_301,N_2996,N_2980);
and UO_302 (O_302,N_2980,N_2940);
or UO_303 (O_303,N_2953,N_2960);
nand UO_304 (O_304,N_2954,N_2996);
or UO_305 (O_305,N_2979,N_2988);
nor UO_306 (O_306,N_2999,N_2992);
or UO_307 (O_307,N_2985,N_2959);
nor UO_308 (O_308,N_2994,N_2963);
or UO_309 (O_309,N_2994,N_2970);
and UO_310 (O_310,N_2999,N_2960);
and UO_311 (O_311,N_2983,N_2972);
xnor UO_312 (O_312,N_2970,N_2989);
xnor UO_313 (O_313,N_2992,N_2947);
or UO_314 (O_314,N_2958,N_2975);
or UO_315 (O_315,N_2965,N_2972);
nor UO_316 (O_316,N_2971,N_2980);
xnor UO_317 (O_317,N_2960,N_2977);
nor UO_318 (O_318,N_2972,N_2957);
or UO_319 (O_319,N_2940,N_2968);
and UO_320 (O_320,N_2989,N_2986);
xnor UO_321 (O_321,N_2971,N_2991);
or UO_322 (O_322,N_2986,N_2946);
nand UO_323 (O_323,N_2967,N_2987);
nor UO_324 (O_324,N_2964,N_2960);
nand UO_325 (O_325,N_2979,N_2950);
nor UO_326 (O_326,N_2984,N_2990);
nor UO_327 (O_327,N_2963,N_2981);
and UO_328 (O_328,N_2972,N_2940);
xnor UO_329 (O_329,N_2998,N_2976);
nor UO_330 (O_330,N_2948,N_2991);
nor UO_331 (O_331,N_2959,N_2973);
or UO_332 (O_332,N_2983,N_2949);
nor UO_333 (O_333,N_2980,N_2954);
and UO_334 (O_334,N_2955,N_2994);
or UO_335 (O_335,N_2941,N_2956);
and UO_336 (O_336,N_2967,N_2958);
and UO_337 (O_337,N_2974,N_2964);
xor UO_338 (O_338,N_2966,N_2969);
or UO_339 (O_339,N_2966,N_2956);
and UO_340 (O_340,N_2989,N_2974);
nand UO_341 (O_341,N_2963,N_2995);
or UO_342 (O_342,N_2999,N_2991);
or UO_343 (O_343,N_2998,N_2971);
and UO_344 (O_344,N_2974,N_2966);
nor UO_345 (O_345,N_2975,N_2980);
or UO_346 (O_346,N_2963,N_2992);
xor UO_347 (O_347,N_2967,N_2954);
or UO_348 (O_348,N_2955,N_2979);
xnor UO_349 (O_349,N_2955,N_2992);
and UO_350 (O_350,N_2952,N_2966);
nor UO_351 (O_351,N_2950,N_2991);
or UO_352 (O_352,N_2985,N_2966);
or UO_353 (O_353,N_2945,N_2948);
nor UO_354 (O_354,N_2985,N_2981);
xor UO_355 (O_355,N_2966,N_2958);
or UO_356 (O_356,N_2999,N_2965);
or UO_357 (O_357,N_2953,N_2980);
and UO_358 (O_358,N_2992,N_2991);
nor UO_359 (O_359,N_2944,N_2962);
or UO_360 (O_360,N_2946,N_2948);
or UO_361 (O_361,N_2955,N_2988);
and UO_362 (O_362,N_2950,N_2967);
or UO_363 (O_363,N_2997,N_2977);
nor UO_364 (O_364,N_2993,N_2984);
xor UO_365 (O_365,N_2964,N_2953);
nor UO_366 (O_366,N_2991,N_2969);
xnor UO_367 (O_367,N_2963,N_2998);
nand UO_368 (O_368,N_2958,N_2949);
nor UO_369 (O_369,N_2994,N_2945);
nor UO_370 (O_370,N_2995,N_2980);
xnor UO_371 (O_371,N_2978,N_2977);
or UO_372 (O_372,N_2958,N_2945);
xor UO_373 (O_373,N_2980,N_2957);
and UO_374 (O_374,N_2975,N_2952);
nor UO_375 (O_375,N_2996,N_2977);
nand UO_376 (O_376,N_2948,N_2959);
or UO_377 (O_377,N_2948,N_2987);
and UO_378 (O_378,N_2983,N_2969);
nor UO_379 (O_379,N_2991,N_2965);
and UO_380 (O_380,N_2951,N_2959);
nor UO_381 (O_381,N_2947,N_2985);
xor UO_382 (O_382,N_2986,N_2968);
and UO_383 (O_383,N_2947,N_2987);
nor UO_384 (O_384,N_2972,N_2993);
nor UO_385 (O_385,N_2988,N_2982);
and UO_386 (O_386,N_2993,N_2990);
nand UO_387 (O_387,N_2941,N_2977);
xnor UO_388 (O_388,N_2986,N_2940);
and UO_389 (O_389,N_2971,N_2974);
and UO_390 (O_390,N_2967,N_2944);
nand UO_391 (O_391,N_2951,N_2955);
nand UO_392 (O_392,N_2967,N_2965);
and UO_393 (O_393,N_2979,N_2943);
or UO_394 (O_394,N_2968,N_2947);
and UO_395 (O_395,N_2995,N_2965);
and UO_396 (O_396,N_2987,N_2988);
or UO_397 (O_397,N_2997,N_2990);
nand UO_398 (O_398,N_2942,N_2987);
or UO_399 (O_399,N_2946,N_2975);
or UO_400 (O_400,N_2958,N_2973);
nor UO_401 (O_401,N_2943,N_2953);
or UO_402 (O_402,N_2984,N_2942);
nor UO_403 (O_403,N_2972,N_2967);
and UO_404 (O_404,N_2984,N_2989);
nor UO_405 (O_405,N_2961,N_2998);
nor UO_406 (O_406,N_2975,N_2953);
nand UO_407 (O_407,N_2950,N_2997);
xnor UO_408 (O_408,N_2944,N_2946);
nor UO_409 (O_409,N_2976,N_2982);
xor UO_410 (O_410,N_2960,N_2970);
nor UO_411 (O_411,N_2989,N_2971);
nor UO_412 (O_412,N_2962,N_2966);
nor UO_413 (O_413,N_2985,N_2988);
or UO_414 (O_414,N_2967,N_2942);
nor UO_415 (O_415,N_2994,N_2981);
nor UO_416 (O_416,N_2996,N_2991);
nand UO_417 (O_417,N_2977,N_2946);
and UO_418 (O_418,N_2970,N_2982);
nor UO_419 (O_419,N_2966,N_2980);
and UO_420 (O_420,N_2951,N_2965);
or UO_421 (O_421,N_2995,N_2981);
or UO_422 (O_422,N_2982,N_2971);
nor UO_423 (O_423,N_2966,N_2965);
nor UO_424 (O_424,N_2973,N_2984);
or UO_425 (O_425,N_2954,N_2976);
and UO_426 (O_426,N_2987,N_2961);
nand UO_427 (O_427,N_2967,N_2953);
xor UO_428 (O_428,N_2962,N_2965);
nor UO_429 (O_429,N_2992,N_2941);
or UO_430 (O_430,N_2970,N_2984);
nand UO_431 (O_431,N_2983,N_2989);
nand UO_432 (O_432,N_2986,N_2943);
or UO_433 (O_433,N_2977,N_2955);
and UO_434 (O_434,N_2985,N_2980);
and UO_435 (O_435,N_2983,N_2953);
xnor UO_436 (O_436,N_2945,N_2967);
or UO_437 (O_437,N_2962,N_2950);
nand UO_438 (O_438,N_2948,N_2975);
and UO_439 (O_439,N_2942,N_2970);
or UO_440 (O_440,N_2993,N_2951);
or UO_441 (O_441,N_2994,N_2948);
nor UO_442 (O_442,N_2952,N_2991);
nor UO_443 (O_443,N_2991,N_2942);
nor UO_444 (O_444,N_2962,N_2951);
and UO_445 (O_445,N_2963,N_2975);
and UO_446 (O_446,N_2963,N_2977);
nand UO_447 (O_447,N_2954,N_2960);
and UO_448 (O_448,N_2941,N_2973);
and UO_449 (O_449,N_2972,N_2984);
xnor UO_450 (O_450,N_2960,N_2958);
nand UO_451 (O_451,N_2970,N_2963);
or UO_452 (O_452,N_2971,N_2984);
nand UO_453 (O_453,N_2982,N_2953);
xnor UO_454 (O_454,N_2976,N_2948);
or UO_455 (O_455,N_2943,N_2941);
nor UO_456 (O_456,N_2984,N_2988);
nor UO_457 (O_457,N_2956,N_2969);
or UO_458 (O_458,N_2952,N_2978);
or UO_459 (O_459,N_2992,N_2951);
or UO_460 (O_460,N_2967,N_2946);
and UO_461 (O_461,N_2998,N_2966);
xor UO_462 (O_462,N_2983,N_2940);
or UO_463 (O_463,N_2997,N_2953);
or UO_464 (O_464,N_2971,N_2968);
or UO_465 (O_465,N_2974,N_2958);
nor UO_466 (O_466,N_2993,N_2961);
nor UO_467 (O_467,N_2977,N_2942);
and UO_468 (O_468,N_2944,N_2993);
nand UO_469 (O_469,N_2957,N_2943);
or UO_470 (O_470,N_2981,N_2987);
nand UO_471 (O_471,N_2984,N_2997);
and UO_472 (O_472,N_2977,N_2993);
xor UO_473 (O_473,N_2984,N_2964);
or UO_474 (O_474,N_2993,N_2942);
nor UO_475 (O_475,N_2997,N_2976);
xor UO_476 (O_476,N_2940,N_2956);
nand UO_477 (O_477,N_2943,N_2960);
nand UO_478 (O_478,N_2958,N_2996);
nor UO_479 (O_479,N_2985,N_2955);
nand UO_480 (O_480,N_2979,N_2987);
nand UO_481 (O_481,N_2963,N_2957);
nand UO_482 (O_482,N_2987,N_2944);
nor UO_483 (O_483,N_2989,N_2948);
nor UO_484 (O_484,N_2960,N_2950);
nand UO_485 (O_485,N_2950,N_2940);
and UO_486 (O_486,N_2973,N_2961);
nand UO_487 (O_487,N_2979,N_2972);
nor UO_488 (O_488,N_2988,N_2975);
nand UO_489 (O_489,N_2999,N_2952);
and UO_490 (O_490,N_2980,N_2961);
xor UO_491 (O_491,N_2952,N_2955);
nand UO_492 (O_492,N_2967,N_2998);
and UO_493 (O_493,N_2942,N_2955);
nor UO_494 (O_494,N_2958,N_2989);
nor UO_495 (O_495,N_2961,N_2974);
or UO_496 (O_496,N_2967,N_2941);
nand UO_497 (O_497,N_2952,N_2960);
nand UO_498 (O_498,N_2988,N_2999);
and UO_499 (O_499,N_2953,N_2973);
endmodule