module basic_500_3000_500_3_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_473,In_471);
nor U1 (N_1,In_303,In_2);
and U2 (N_2,In_40,In_42);
nand U3 (N_3,In_219,In_35);
nor U4 (N_4,In_314,In_279);
and U5 (N_5,In_237,In_425);
or U6 (N_6,In_407,In_454);
and U7 (N_7,In_347,In_68);
nor U8 (N_8,In_201,In_298);
and U9 (N_9,In_101,In_385);
nor U10 (N_10,In_334,In_146);
nand U11 (N_11,In_175,In_327);
nor U12 (N_12,In_23,In_284);
or U13 (N_13,In_224,In_433);
or U14 (N_14,In_449,In_56);
or U15 (N_15,In_197,In_411);
or U16 (N_16,In_335,In_300);
or U17 (N_17,In_363,In_481);
and U18 (N_18,In_478,In_104);
nor U19 (N_19,In_404,In_384);
nor U20 (N_20,In_212,In_36);
nand U21 (N_21,In_301,In_368);
nor U22 (N_22,In_450,In_244);
nor U23 (N_23,In_488,In_432);
nand U24 (N_24,In_89,In_390);
and U25 (N_25,In_49,In_359);
and U26 (N_26,In_463,In_345);
xnor U27 (N_27,In_263,In_389);
or U28 (N_28,In_154,In_66);
nor U29 (N_29,In_108,In_491);
nand U30 (N_30,In_34,In_323);
and U31 (N_31,In_32,In_168);
or U32 (N_32,In_325,In_487);
and U33 (N_33,In_235,In_147);
nand U34 (N_34,In_475,In_393);
and U35 (N_35,In_412,In_353);
nor U36 (N_36,In_78,In_214);
nand U37 (N_37,In_349,In_132);
or U38 (N_38,In_13,In_99);
nor U39 (N_39,In_11,In_125);
and U40 (N_40,In_302,In_403);
nor U41 (N_41,In_4,In_150);
or U42 (N_42,In_496,In_14);
nor U43 (N_43,In_110,In_285);
nor U44 (N_44,In_243,In_127);
or U45 (N_45,In_230,In_497);
nor U46 (N_46,In_341,In_374);
and U47 (N_47,In_377,In_228);
or U48 (N_48,In_337,In_129);
nor U49 (N_49,In_207,In_469);
or U50 (N_50,In_198,In_88);
and U51 (N_51,In_131,In_161);
nor U52 (N_52,In_258,In_107);
and U53 (N_53,In_157,In_382);
nor U54 (N_54,In_241,In_142);
and U55 (N_55,In_330,In_152);
nor U56 (N_56,In_85,In_116);
or U57 (N_57,In_402,In_405);
or U58 (N_58,In_238,In_466);
nor U59 (N_59,In_242,In_313);
nor U60 (N_60,In_398,In_455);
nor U61 (N_61,In_416,In_312);
and U62 (N_62,In_311,In_262);
nor U63 (N_63,In_134,In_184);
or U64 (N_64,In_26,In_435);
and U65 (N_65,In_418,In_80);
nor U66 (N_66,In_48,In_268);
and U67 (N_67,In_117,In_60);
and U68 (N_68,In_441,In_401);
or U69 (N_69,In_287,In_145);
nand U70 (N_70,In_222,In_342);
nand U71 (N_71,In_5,In_319);
nand U72 (N_72,In_409,In_159);
nand U73 (N_73,In_153,In_223);
nand U74 (N_74,In_477,In_351);
nor U75 (N_75,In_289,In_255);
or U76 (N_76,In_354,In_379);
and U77 (N_77,In_74,In_278);
or U78 (N_78,In_167,In_249);
nor U79 (N_79,In_442,In_294);
nand U80 (N_80,In_120,In_430);
and U81 (N_81,In_59,In_218);
nand U82 (N_82,In_483,In_364);
or U83 (N_83,In_121,In_71);
nand U84 (N_84,In_163,In_93);
or U85 (N_85,In_63,In_286);
and U86 (N_86,In_424,In_106);
nor U87 (N_87,In_370,In_37);
nand U88 (N_88,In_231,In_20);
or U89 (N_89,In_306,In_188);
and U90 (N_90,In_461,In_98);
or U91 (N_91,In_415,In_148);
nand U92 (N_92,In_67,In_328);
or U93 (N_93,In_87,In_413);
nand U94 (N_94,In_465,In_169);
and U95 (N_95,In_427,In_358);
or U96 (N_96,In_191,In_86);
and U97 (N_97,In_397,In_355);
or U98 (N_98,In_375,In_299);
nor U99 (N_99,In_82,In_220);
nand U100 (N_100,In_408,In_336);
and U101 (N_101,In_250,In_315);
nand U102 (N_102,In_421,In_76);
nand U103 (N_103,In_190,In_348);
and U104 (N_104,In_261,In_304);
or U105 (N_105,In_96,In_25);
or U106 (N_106,In_309,In_266);
or U107 (N_107,In_138,In_317);
nand U108 (N_108,In_44,In_339);
nand U109 (N_109,In_170,In_196);
or U110 (N_110,In_29,In_73);
nor U111 (N_111,In_199,In_492);
or U112 (N_112,In_171,In_137);
nor U113 (N_113,In_77,In_293);
or U114 (N_114,In_136,In_467);
or U115 (N_115,In_6,In_39);
nand U116 (N_116,In_177,In_254);
nand U117 (N_117,In_16,In_352);
or U118 (N_118,In_178,In_124);
or U119 (N_119,In_9,In_431);
and U120 (N_120,In_444,In_360);
nor U121 (N_121,In_308,In_216);
or U122 (N_122,In_46,In_480);
nand U123 (N_123,In_162,In_396);
or U124 (N_124,In_380,In_252);
nand U125 (N_125,In_172,In_484);
and U126 (N_126,In_7,In_156);
and U127 (N_127,In_62,In_0);
and U128 (N_128,In_105,In_346);
and U129 (N_129,In_64,In_19);
nand U130 (N_130,In_386,In_305);
nor U131 (N_131,In_493,In_392);
or U132 (N_132,In_422,In_256);
and U133 (N_133,In_118,In_232);
nand U134 (N_134,In_123,In_217);
nand U135 (N_135,In_61,In_320);
or U136 (N_136,In_221,In_264);
nor U137 (N_137,In_280,In_208);
nor U138 (N_138,In_17,In_155);
or U139 (N_139,In_419,In_183);
nor U140 (N_140,In_369,In_271);
nand U141 (N_141,In_443,In_58);
nand U142 (N_142,In_50,In_179);
and U143 (N_143,In_111,In_437);
and U144 (N_144,In_195,In_367);
nor U145 (N_145,In_438,In_236);
nand U146 (N_146,In_47,In_429);
nor U147 (N_147,In_149,In_55);
nor U148 (N_148,In_53,In_296);
nand U149 (N_149,In_457,In_251);
or U150 (N_150,In_324,In_79);
nor U151 (N_151,In_468,In_187);
nand U152 (N_152,In_69,In_176);
nand U153 (N_153,In_371,In_316);
nand U154 (N_154,In_290,In_119);
nor U155 (N_155,In_267,In_388);
or U156 (N_156,In_229,In_453);
nand U157 (N_157,In_90,In_248);
or U158 (N_158,In_322,In_45);
nor U159 (N_159,In_310,In_372);
nand U160 (N_160,In_344,In_321);
nor U161 (N_161,In_357,In_10);
nor U162 (N_162,In_391,In_452);
nand U163 (N_163,In_213,In_464);
nand U164 (N_164,In_318,In_297);
nor U165 (N_165,In_31,In_54);
nand U166 (N_166,In_362,In_406);
nor U167 (N_167,In_28,In_192);
and U168 (N_168,In_22,In_140);
and U169 (N_169,In_126,In_265);
and U170 (N_170,In_122,In_494);
nand U171 (N_171,In_376,In_259);
or U172 (N_172,In_440,In_102);
and U173 (N_173,In_21,In_165);
nand U174 (N_174,In_194,In_135);
or U175 (N_175,In_30,In_141);
or U176 (N_176,In_246,In_225);
nand U177 (N_177,In_373,In_12);
and U178 (N_178,In_272,In_114);
and U179 (N_179,In_459,In_41);
and U180 (N_180,In_182,In_283);
or U181 (N_181,In_112,In_288);
or U182 (N_182,In_479,In_482);
nand U183 (N_183,In_72,In_245);
nor U184 (N_184,In_203,In_428);
nand U185 (N_185,In_383,In_128);
nor U186 (N_186,In_83,In_498);
or U187 (N_187,In_340,In_326);
or U188 (N_188,In_333,In_151);
nor U189 (N_189,In_164,In_239);
nand U190 (N_190,In_173,In_426);
nand U191 (N_191,In_395,In_206);
and U192 (N_192,In_439,In_174);
and U193 (N_193,In_185,In_276);
nand U194 (N_194,In_269,In_260);
xor U195 (N_195,In_24,In_92);
and U196 (N_196,In_447,In_356);
nor U197 (N_197,In_247,In_281);
and U198 (N_198,In_234,In_350);
nor U199 (N_199,In_144,In_448);
or U200 (N_200,In_489,In_1);
or U201 (N_201,In_109,In_462);
or U202 (N_202,In_410,In_193);
nor U203 (N_203,In_130,In_329);
or U204 (N_204,In_227,In_139);
and U205 (N_205,In_270,In_75);
nor U206 (N_206,In_18,In_15);
nor U207 (N_207,In_434,In_474);
nand U208 (N_208,In_277,In_446);
nor U209 (N_209,In_97,In_233);
and U210 (N_210,In_189,In_52);
nor U211 (N_211,In_70,In_209);
and U212 (N_212,In_282,In_200);
nor U213 (N_213,In_486,In_115);
nor U214 (N_214,In_81,In_181);
or U215 (N_215,In_100,In_8);
or U216 (N_216,In_343,In_51);
or U217 (N_217,In_257,In_458);
or U218 (N_218,In_33,In_275);
and U219 (N_219,In_436,In_166);
and U220 (N_220,In_400,In_451);
and U221 (N_221,In_215,In_361);
or U222 (N_222,In_476,In_253);
and U223 (N_223,In_113,In_186);
xor U224 (N_224,In_160,In_95);
nor U225 (N_225,In_381,In_399);
nor U226 (N_226,In_204,In_133);
nand U227 (N_227,In_211,In_240);
and U228 (N_228,In_91,In_94);
and U229 (N_229,In_423,In_158);
or U230 (N_230,In_365,In_226);
nor U231 (N_231,In_274,In_273);
and U232 (N_232,In_103,In_43);
or U233 (N_233,In_3,In_338);
nand U234 (N_234,In_27,In_490);
or U235 (N_235,In_65,In_84);
nor U236 (N_236,In_472,In_460);
nor U237 (N_237,In_366,In_456);
nand U238 (N_238,In_57,In_485);
nand U239 (N_239,In_394,In_202);
nor U240 (N_240,In_205,In_307);
nor U241 (N_241,In_378,In_414);
nor U242 (N_242,In_499,In_332);
nand U243 (N_243,In_417,In_180);
and U244 (N_244,In_387,In_420);
nand U245 (N_245,In_445,In_291);
nand U246 (N_246,In_38,In_295);
nand U247 (N_247,In_143,In_210);
nand U248 (N_248,In_292,In_331);
nand U249 (N_249,In_470,In_495);
or U250 (N_250,In_284,In_374);
nand U251 (N_251,In_207,In_263);
and U252 (N_252,In_57,In_385);
and U253 (N_253,In_362,In_142);
or U254 (N_254,In_423,In_214);
nand U255 (N_255,In_457,In_376);
nand U256 (N_256,In_403,In_333);
nor U257 (N_257,In_480,In_158);
nand U258 (N_258,In_124,In_148);
or U259 (N_259,In_142,In_147);
nor U260 (N_260,In_448,In_289);
and U261 (N_261,In_450,In_146);
or U262 (N_262,In_320,In_393);
and U263 (N_263,In_421,In_185);
or U264 (N_264,In_274,In_213);
or U265 (N_265,In_214,In_174);
and U266 (N_266,In_64,In_50);
nand U267 (N_267,In_45,In_445);
nand U268 (N_268,In_6,In_43);
and U269 (N_269,In_260,In_476);
nand U270 (N_270,In_240,In_365);
nor U271 (N_271,In_398,In_396);
or U272 (N_272,In_140,In_14);
nand U273 (N_273,In_240,In_434);
and U274 (N_274,In_135,In_410);
nand U275 (N_275,In_38,In_106);
or U276 (N_276,In_56,In_71);
and U277 (N_277,In_32,In_396);
and U278 (N_278,In_132,In_434);
nand U279 (N_279,In_426,In_102);
nand U280 (N_280,In_155,In_470);
nor U281 (N_281,In_302,In_12);
nor U282 (N_282,In_305,In_381);
nand U283 (N_283,In_164,In_63);
nand U284 (N_284,In_368,In_214);
and U285 (N_285,In_118,In_120);
and U286 (N_286,In_189,In_18);
nor U287 (N_287,In_247,In_106);
nand U288 (N_288,In_383,In_356);
nor U289 (N_289,In_45,In_468);
nand U290 (N_290,In_255,In_435);
nand U291 (N_291,In_258,In_105);
or U292 (N_292,In_185,In_44);
and U293 (N_293,In_327,In_99);
and U294 (N_294,In_213,In_226);
nand U295 (N_295,In_241,In_80);
nor U296 (N_296,In_76,In_225);
nor U297 (N_297,In_439,In_180);
nand U298 (N_298,In_385,In_19);
nand U299 (N_299,In_125,In_489);
nand U300 (N_300,In_380,In_243);
or U301 (N_301,In_249,In_282);
xnor U302 (N_302,In_460,In_320);
nor U303 (N_303,In_300,In_228);
nor U304 (N_304,In_72,In_366);
nor U305 (N_305,In_190,In_285);
and U306 (N_306,In_154,In_266);
or U307 (N_307,In_141,In_182);
nor U308 (N_308,In_62,In_80);
and U309 (N_309,In_398,In_118);
nand U310 (N_310,In_164,In_14);
nand U311 (N_311,In_275,In_72);
and U312 (N_312,In_203,In_269);
and U313 (N_313,In_234,In_225);
and U314 (N_314,In_80,In_29);
or U315 (N_315,In_305,In_495);
xnor U316 (N_316,In_46,In_356);
xnor U317 (N_317,In_134,In_395);
and U318 (N_318,In_454,In_54);
nand U319 (N_319,In_189,In_455);
nand U320 (N_320,In_480,In_447);
nor U321 (N_321,In_103,In_466);
and U322 (N_322,In_64,In_122);
and U323 (N_323,In_411,In_17);
or U324 (N_324,In_353,In_63);
or U325 (N_325,In_486,In_7);
nand U326 (N_326,In_88,In_286);
and U327 (N_327,In_227,In_20);
nand U328 (N_328,In_389,In_274);
or U329 (N_329,In_351,In_393);
nor U330 (N_330,In_437,In_399);
or U331 (N_331,In_300,In_80);
or U332 (N_332,In_289,In_433);
nor U333 (N_333,In_391,In_386);
or U334 (N_334,In_277,In_413);
nand U335 (N_335,In_461,In_385);
nor U336 (N_336,In_166,In_373);
nor U337 (N_337,In_380,In_283);
or U338 (N_338,In_352,In_421);
or U339 (N_339,In_164,In_256);
or U340 (N_340,In_57,In_190);
or U341 (N_341,In_112,In_292);
or U342 (N_342,In_244,In_173);
nor U343 (N_343,In_319,In_470);
nand U344 (N_344,In_182,In_204);
nor U345 (N_345,In_333,In_224);
nor U346 (N_346,In_158,In_128);
or U347 (N_347,In_372,In_253);
or U348 (N_348,In_306,In_36);
nor U349 (N_349,In_33,In_142);
or U350 (N_350,In_371,In_320);
and U351 (N_351,In_236,In_279);
and U352 (N_352,In_333,In_42);
nor U353 (N_353,In_157,In_71);
nor U354 (N_354,In_66,In_1);
and U355 (N_355,In_190,In_410);
or U356 (N_356,In_259,In_203);
and U357 (N_357,In_301,In_341);
and U358 (N_358,In_307,In_380);
nand U359 (N_359,In_176,In_82);
or U360 (N_360,In_135,In_29);
or U361 (N_361,In_188,In_284);
xor U362 (N_362,In_299,In_209);
nand U363 (N_363,In_488,In_149);
or U364 (N_364,In_290,In_21);
and U365 (N_365,In_318,In_236);
nand U366 (N_366,In_18,In_242);
nand U367 (N_367,In_238,In_60);
and U368 (N_368,In_471,In_331);
and U369 (N_369,In_287,In_275);
and U370 (N_370,In_105,In_455);
nor U371 (N_371,In_433,In_371);
nand U372 (N_372,In_276,In_445);
or U373 (N_373,In_477,In_92);
nand U374 (N_374,In_476,In_394);
or U375 (N_375,In_53,In_80);
or U376 (N_376,In_257,In_214);
and U377 (N_377,In_162,In_433);
nor U378 (N_378,In_23,In_188);
nor U379 (N_379,In_352,In_97);
or U380 (N_380,In_401,In_74);
or U381 (N_381,In_234,In_424);
nor U382 (N_382,In_195,In_442);
and U383 (N_383,In_237,In_17);
nand U384 (N_384,In_74,In_334);
and U385 (N_385,In_451,In_167);
and U386 (N_386,In_175,In_29);
and U387 (N_387,In_15,In_68);
and U388 (N_388,In_318,In_326);
xnor U389 (N_389,In_55,In_82);
nor U390 (N_390,In_129,In_214);
nor U391 (N_391,In_260,In_238);
nand U392 (N_392,In_339,In_497);
nand U393 (N_393,In_490,In_126);
nor U394 (N_394,In_284,In_269);
or U395 (N_395,In_200,In_147);
nor U396 (N_396,In_407,In_352);
nand U397 (N_397,In_284,In_43);
or U398 (N_398,In_134,In_283);
and U399 (N_399,In_201,In_351);
nor U400 (N_400,In_435,In_278);
or U401 (N_401,In_479,In_8);
or U402 (N_402,In_228,In_134);
nor U403 (N_403,In_216,In_424);
xnor U404 (N_404,In_355,In_475);
or U405 (N_405,In_447,In_335);
nor U406 (N_406,In_122,In_202);
and U407 (N_407,In_259,In_188);
nand U408 (N_408,In_243,In_419);
and U409 (N_409,In_396,In_124);
and U410 (N_410,In_445,In_80);
nand U411 (N_411,In_1,In_392);
or U412 (N_412,In_332,In_329);
nand U413 (N_413,In_386,In_35);
and U414 (N_414,In_364,In_448);
and U415 (N_415,In_339,In_486);
nor U416 (N_416,In_37,In_248);
nand U417 (N_417,In_42,In_344);
nand U418 (N_418,In_480,In_216);
or U419 (N_419,In_128,In_272);
or U420 (N_420,In_201,In_93);
nand U421 (N_421,In_475,In_395);
or U422 (N_422,In_386,In_38);
nor U423 (N_423,In_496,In_6);
and U424 (N_424,In_234,In_412);
nand U425 (N_425,In_483,In_361);
and U426 (N_426,In_400,In_100);
nor U427 (N_427,In_425,In_323);
nor U428 (N_428,In_130,In_231);
nor U429 (N_429,In_40,In_189);
nand U430 (N_430,In_301,In_26);
nor U431 (N_431,In_75,In_493);
nor U432 (N_432,In_176,In_38);
or U433 (N_433,In_497,In_291);
nand U434 (N_434,In_443,In_13);
or U435 (N_435,In_315,In_35);
nor U436 (N_436,In_209,In_49);
nor U437 (N_437,In_240,In_356);
nor U438 (N_438,In_165,In_48);
nand U439 (N_439,In_366,In_77);
nand U440 (N_440,In_319,In_488);
nor U441 (N_441,In_237,In_150);
nor U442 (N_442,In_253,In_347);
or U443 (N_443,In_421,In_439);
nand U444 (N_444,In_257,In_452);
nand U445 (N_445,In_78,In_25);
or U446 (N_446,In_265,In_208);
nand U447 (N_447,In_23,In_262);
nor U448 (N_448,In_261,In_449);
nand U449 (N_449,In_273,In_101);
and U450 (N_450,In_75,In_107);
and U451 (N_451,In_390,In_307);
or U452 (N_452,In_337,In_79);
and U453 (N_453,In_297,In_437);
or U454 (N_454,In_248,In_186);
nand U455 (N_455,In_364,In_41);
nor U456 (N_456,In_332,In_463);
nand U457 (N_457,In_471,In_364);
or U458 (N_458,In_289,In_377);
nand U459 (N_459,In_3,In_229);
nor U460 (N_460,In_128,In_16);
nor U461 (N_461,In_82,In_269);
and U462 (N_462,In_490,In_269);
or U463 (N_463,In_137,In_42);
nand U464 (N_464,In_440,In_33);
nand U465 (N_465,In_196,In_129);
or U466 (N_466,In_117,In_140);
or U467 (N_467,In_14,In_439);
nand U468 (N_468,In_138,In_486);
and U469 (N_469,In_484,In_73);
and U470 (N_470,In_54,In_44);
and U471 (N_471,In_168,In_209);
and U472 (N_472,In_454,In_366);
and U473 (N_473,In_326,In_180);
and U474 (N_474,In_295,In_388);
nor U475 (N_475,In_402,In_353);
or U476 (N_476,In_401,In_247);
and U477 (N_477,In_336,In_199);
nor U478 (N_478,In_457,In_48);
or U479 (N_479,In_406,In_379);
nor U480 (N_480,In_100,In_15);
nor U481 (N_481,In_17,In_454);
nor U482 (N_482,In_72,In_452);
nand U483 (N_483,In_57,In_4);
nor U484 (N_484,In_430,In_241);
and U485 (N_485,In_492,In_410);
nand U486 (N_486,In_31,In_495);
nand U487 (N_487,In_343,In_5);
and U488 (N_488,In_287,In_172);
and U489 (N_489,In_175,In_376);
or U490 (N_490,In_488,In_341);
nor U491 (N_491,In_52,In_214);
nor U492 (N_492,In_335,In_150);
nand U493 (N_493,In_353,In_401);
nand U494 (N_494,In_174,In_36);
or U495 (N_495,In_399,In_319);
nand U496 (N_496,In_303,In_480);
or U497 (N_497,In_104,In_462);
and U498 (N_498,In_479,In_497);
nor U499 (N_499,In_304,In_13);
and U500 (N_500,In_233,In_486);
and U501 (N_501,In_381,In_466);
and U502 (N_502,In_207,In_280);
or U503 (N_503,In_241,In_411);
nor U504 (N_504,In_317,In_483);
or U505 (N_505,In_383,In_150);
nor U506 (N_506,In_413,In_279);
nor U507 (N_507,In_405,In_320);
nor U508 (N_508,In_213,In_279);
or U509 (N_509,In_176,In_374);
nor U510 (N_510,In_113,In_291);
or U511 (N_511,In_169,In_253);
nor U512 (N_512,In_386,In_72);
nor U513 (N_513,In_442,In_74);
nor U514 (N_514,In_7,In_424);
nand U515 (N_515,In_376,In_497);
and U516 (N_516,In_63,In_212);
nand U517 (N_517,In_385,In_288);
nand U518 (N_518,In_372,In_184);
or U519 (N_519,In_211,In_58);
and U520 (N_520,In_57,In_172);
or U521 (N_521,In_487,In_476);
nor U522 (N_522,In_161,In_368);
nand U523 (N_523,In_415,In_122);
nand U524 (N_524,In_59,In_326);
or U525 (N_525,In_81,In_251);
nor U526 (N_526,In_203,In_73);
or U527 (N_527,In_129,In_96);
and U528 (N_528,In_24,In_262);
nor U529 (N_529,In_118,In_449);
nor U530 (N_530,In_102,In_260);
and U531 (N_531,In_291,In_309);
nand U532 (N_532,In_239,In_181);
and U533 (N_533,In_338,In_71);
or U534 (N_534,In_290,In_53);
nor U535 (N_535,In_191,In_471);
or U536 (N_536,In_125,In_19);
nand U537 (N_537,In_170,In_241);
nand U538 (N_538,In_225,In_466);
nand U539 (N_539,In_404,In_306);
nor U540 (N_540,In_350,In_111);
and U541 (N_541,In_474,In_283);
and U542 (N_542,In_158,In_408);
or U543 (N_543,In_264,In_124);
nor U544 (N_544,In_423,In_61);
or U545 (N_545,In_394,In_378);
nand U546 (N_546,In_471,In_301);
or U547 (N_547,In_104,In_223);
and U548 (N_548,In_52,In_347);
nand U549 (N_549,In_438,In_344);
and U550 (N_550,In_178,In_126);
and U551 (N_551,In_84,In_354);
nor U552 (N_552,In_264,In_447);
nand U553 (N_553,In_339,In_58);
or U554 (N_554,In_177,In_89);
nor U555 (N_555,In_440,In_274);
nand U556 (N_556,In_74,In_165);
nor U557 (N_557,In_181,In_246);
nor U558 (N_558,In_213,In_458);
nand U559 (N_559,In_287,In_9);
nand U560 (N_560,In_272,In_256);
nand U561 (N_561,In_120,In_296);
and U562 (N_562,In_469,In_43);
nor U563 (N_563,In_31,In_418);
nor U564 (N_564,In_409,In_94);
nand U565 (N_565,In_66,In_169);
or U566 (N_566,In_398,In_429);
and U567 (N_567,In_248,In_377);
nor U568 (N_568,In_160,In_117);
xor U569 (N_569,In_271,In_496);
nand U570 (N_570,In_159,In_227);
or U571 (N_571,In_416,In_48);
and U572 (N_572,In_109,In_181);
or U573 (N_573,In_177,In_480);
and U574 (N_574,In_325,In_411);
nor U575 (N_575,In_487,In_78);
nand U576 (N_576,In_133,In_360);
xor U577 (N_577,In_422,In_346);
or U578 (N_578,In_413,In_429);
and U579 (N_579,In_490,In_357);
or U580 (N_580,In_485,In_297);
nand U581 (N_581,In_419,In_433);
and U582 (N_582,In_259,In_462);
nor U583 (N_583,In_211,In_193);
nand U584 (N_584,In_176,In_306);
and U585 (N_585,In_251,In_267);
and U586 (N_586,In_7,In_102);
and U587 (N_587,In_334,In_440);
nor U588 (N_588,In_5,In_99);
and U589 (N_589,In_209,In_244);
and U590 (N_590,In_155,In_13);
nor U591 (N_591,In_16,In_332);
and U592 (N_592,In_70,In_81);
nand U593 (N_593,In_223,In_73);
or U594 (N_594,In_446,In_47);
or U595 (N_595,In_165,In_188);
nor U596 (N_596,In_416,In_479);
nand U597 (N_597,In_307,In_376);
nand U598 (N_598,In_385,In_124);
and U599 (N_599,In_200,In_254);
or U600 (N_600,In_44,In_267);
and U601 (N_601,In_464,In_38);
and U602 (N_602,In_259,In_495);
nor U603 (N_603,In_395,In_423);
and U604 (N_604,In_437,In_85);
or U605 (N_605,In_250,In_479);
and U606 (N_606,In_83,In_456);
or U607 (N_607,In_237,In_46);
nor U608 (N_608,In_105,In_112);
nand U609 (N_609,In_111,In_295);
and U610 (N_610,In_202,In_161);
nand U611 (N_611,In_278,In_274);
or U612 (N_612,In_326,In_153);
or U613 (N_613,In_24,In_13);
or U614 (N_614,In_402,In_460);
nand U615 (N_615,In_459,In_342);
or U616 (N_616,In_375,In_124);
or U617 (N_617,In_12,In_37);
nand U618 (N_618,In_327,In_118);
or U619 (N_619,In_59,In_179);
and U620 (N_620,In_402,In_355);
nor U621 (N_621,In_187,In_193);
or U622 (N_622,In_232,In_274);
nand U623 (N_623,In_359,In_110);
and U624 (N_624,In_442,In_467);
and U625 (N_625,In_30,In_441);
nand U626 (N_626,In_157,In_283);
or U627 (N_627,In_114,In_494);
and U628 (N_628,In_269,In_224);
and U629 (N_629,In_254,In_371);
nand U630 (N_630,In_33,In_171);
nor U631 (N_631,In_9,In_17);
nor U632 (N_632,In_135,In_318);
nor U633 (N_633,In_316,In_411);
and U634 (N_634,In_26,In_449);
and U635 (N_635,In_7,In_44);
and U636 (N_636,In_337,In_36);
and U637 (N_637,In_335,In_18);
nand U638 (N_638,In_236,In_129);
nand U639 (N_639,In_50,In_174);
and U640 (N_640,In_265,In_46);
and U641 (N_641,In_0,In_492);
nor U642 (N_642,In_165,In_88);
and U643 (N_643,In_160,In_30);
nor U644 (N_644,In_391,In_484);
nor U645 (N_645,In_108,In_412);
nor U646 (N_646,In_183,In_29);
or U647 (N_647,In_464,In_113);
nand U648 (N_648,In_467,In_343);
nor U649 (N_649,In_140,In_159);
nor U650 (N_650,In_418,In_316);
or U651 (N_651,In_210,In_403);
nor U652 (N_652,In_333,In_186);
nand U653 (N_653,In_56,In_108);
nor U654 (N_654,In_339,In_77);
or U655 (N_655,In_117,In_422);
and U656 (N_656,In_334,In_26);
nor U657 (N_657,In_369,In_140);
nand U658 (N_658,In_360,In_404);
and U659 (N_659,In_457,In_353);
or U660 (N_660,In_289,In_458);
or U661 (N_661,In_414,In_274);
nor U662 (N_662,In_373,In_63);
nand U663 (N_663,In_113,In_326);
nor U664 (N_664,In_51,In_148);
and U665 (N_665,In_259,In_13);
or U666 (N_666,In_158,In_228);
nand U667 (N_667,In_407,In_370);
nand U668 (N_668,In_69,In_114);
or U669 (N_669,In_114,In_453);
nor U670 (N_670,In_163,In_206);
nand U671 (N_671,In_384,In_444);
and U672 (N_672,In_428,In_300);
nor U673 (N_673,In_7,In_455);
nand U674 (N_674,In_349,In_406);
xor U675 (N_675,In_221,In_285);
or U676 (N_676,In_358,In_284);
and U677 (N_677,In_446,In_455);
nor U678 (N_678,In_494,In_242);
nor U679 (N_679,In_19,In_215);
and U680 (N_680,In_346,In_3);
or U681 (N_681,In_196,In_315);
and U682 (N_682,In_351,In_341);
nand U683 (N_683,In_91,In_2);
and U684 (N_684,In_89,In_103);
and U685 (N_685,In_364,In_240);
nor U686 (N_686,In_88,In_25);
nor U687 (N_687,In_221,In_375);
nor U688 (N_688,In_388,In_140);
or U689 (N_689,In_100,In_30);
or U690 (N_690,In_328,In_47);
nand U691 (N_691,In_94,In_432);
nand U692 (N_692,In_60,In_143);
and U693 (N_693,In_8,In_6);
nor U694 (N_694,In_105,In_445);
and U695 (N_695,In_94,In_256);
and U696 (N_696,In_157,In_38);
or U697 (N_697,In_427,In_417);
or U698 (N_698,In_322,In_437);
nor U699 (N_699,In_76,In_244);
nor U700 (N_700,In_164,In_17);
or U701 (N_701,In_455,In_279);
or U702 (N_702,In_240,In_251);
nand U703 (N_703,In_451,In_296);
nor U704 (N_704,In_358,In_48);
or U705 (N_705,In_463,In_25);
nand U706 (N_706,In_145,In_133);
nand U707 (N_707,In_267,In_372);
nor U708 (N_708,In_43,In_106);
and U709 (N_709,In_318,In_206);
or U710 (N_710,In_275,In_180);
nor U711 (N_711,In_385,In_223);
nand U712 (N_712,In_145,In_257);
nand U713 (N_713,In_445,In_328);
nand U714 (N_714,In_454,In_493);
nand U715 (N_715,In_454,In_162);
or U716 (N_716,In_345,In_236);
or U717 (N_717,In_280,In_261);
or U718 (N_718,In_345,In_377);
nand U719 (N_719,In_426,In_441);
nand U720 (N_720,In_132,In_172);
nand U721 (N_721,In_222,In_233);
or U722 (N_722,In_215,In_434);
or U723 (N_723,In_312,In_109);
nand U724 (N_724,In_498,In_265);
nor U725 (N_725,In_117,In_330);
nand U726 (N_726,In_382,In_427);
or U727 (N_727,In_381,In_258);
and U728 (N_728,In_221,In_22);
or U729 (N_729,In_432,In_435);
and U730 (N_730,In_249,In_148);
or U731 (N_731,In_296,In_141);
and U732 (N_732,In_420,In_57);
or U733 (N_733,In_348,In_399);
nor U734 (N_734,In_253,In_243);
or U735 (N_735,In_436,In_25);
nand U736 (N_736,In_156,In_22);
nand U737 (N_737,In_117,In_119);
nand U738 (N_738,In_19,In_487);
or U739 (N_739,In_395,In_192);
or U740 (N_740,In_417,In_7);
nand U741 (N_741,In_233,In_129);
or U742 (N_742,In_427,In_144);
nand U743 (N_743,In_442,In_214);
nor U744 (N_744,In_80,In_338);
nor U745 (N_745,In_157,In_467);
nand U746 (N_746,In_106,In_26);
nor U747 (N_747,In_374,In_433);
nor U748 (N_748,In_316,In_429);
or U749 (N_749,In_127,In_241);
nand U750 (N_750,In_396,In_294);
nor U751 (N_751,In_236,In_84);
nand U752 (N_752,In_7,In_182);
nor U753 (N_753,In_491,In_140);
and U754 (N_754,In_451,In_469);
and U755 (N_755,In_410,In_248);
and U756 (N_756,In_325,In_163);
nor U757 (N_757,In_265,In_206);
and U758 (N_758,In_222,In_412);
nand U759 (N_759,In_482,In_10);
and U760 (N_760,In_15,In_202);
and U761 (N_761,In_70,In_212);
or U762 (N_762,In_136,In_407);
and U763 (N_763,In_253,In_71);
and U764 (N_764,In_299,In_325);
nand U765 (N_765,In_66,In_460);
nor U766 (N_766,In_389,In_479);
or U767 (N_767,In_356,In_178);
and U768 (N_768,In_315,In_39);
and U769 (N_769,In_119,In_24);
and U770 (N_770,In_126,In_14);
or U771 (N_771,In_325,In_9);
nand U772 (N_772,In_52,In_367);
and U773 (N_773,In_337,In_174);
nor U774 (N_774,In_234,In_456);
nor U775 (N_775,In_52,In_421);
nor U776 (N_776,In_297,In_219);
nand U777 (N_777,In_175,In_416);
nor U778 (N_778,In_494,In_444);
and U779 (N_779,In_458,In_47);
or U780 (N_780,In_131,In_28);
and U781 (N_781,In_457,In_151);
or U782 (N_782,In_80,In_323);
nor U783 (N_783,In_394,In_159);
and U784 (N_784,In_337,In_144);
nand U785 (N_785,In_480,In_6);
or U786 (N_786,In_208,In_142);
and U787 (N_787,In_306,In_148);
and U788 (N_788,In_296,In_83);
and U789 (N_789,In_423,In_118);
and U790 (N_790,In_151,In_442);
nor U791 (N_791,In_136,In_372);
or U792 (N_792,In_88,In_299);
nor U793 (N_793,In_320,In_103);
nor U794 (N_794,In_42,In_205);
nand U795 (N_795,In_293,In_393);
nand U796 (N_796,In_18,In_454);
nand U797 (N_797,In_32,In_114);
and U798 (N_798,In_13,In_273);
or U799 (N_799,In_347,In_298);
nor U800 (N_800,In_113,In_232);
or U801 (N_801,In_117,In_350);
and U802 (N_802,In_469,In_186);
and U803 (N_803,In_10,In_236);
nor U804 (N_804,In_320,In_438);
nor U805 (N_805,In_150,In_409);
nand U806 (N_806,In_392,In_342);
nand U807 (N_807,In_359,In_262);
and U808 (N_808,In_404,In_34);
and U809 (N_809,In_44,In_315);
nand U810 (N_810,In_202,In_403);
or U811 (N_811,In_201,In_367);
and U812 (N_812,In_69,In_490);
nand U813 (N_813,In_48,In_447);
nand U814 (N_814,In_299,In_55);
or U815 (N_815,In_22,In_147);
nor U816 (N_816,In_279,In_59);
nor U817 (N_817,In_359,In_395);
nor U818 (N_818,In_453,In_224);
or U819 (N_819,In_102,In_2);
nand U820 (N_820,In_49,In_341);
or U821 (N_821,In_43,In_373);
or U822 (N_822,In_350,In_159);
and U823 (N_823,In_237,In_348);
and U824 (N_824,In_304,In_271);
nor U825 (N_825,In_338,In_6);
nor U826 (N_826,In_251,In_283);
nor U827 (N_827,In_8,In_81);
nand U828 (N_828,In_352,In_254);
or U829 (N_829,In_22,In_430);
nand U830 (N_830,In_340,In_45);
and U831 (N_831,In_161,In_171);
or U832 (N_832,In_384,In_104);
and U833 (N_833,In_468,In_58);
nor U834 (N_834,In_169,In_452);
nand U835 (N_835,In_390,In_23);
nor U836 (N_836,In_124,In_327);
and U837 (N_837,In_488,In_381);
or U838 (N_838,In_350,In_232);
nand U839 (N_839,In_51,In_95);
or U840 (N_840,In_342,In_245);
nor U841 (N_841,In_134,In_470);
nand U842 (N_842,In_10,In_90);
or U843 (N_843,In_454,In_147);
and U844 (N_844,In_209,In_46);
nor U845 (N_845,In_220,In_118);
or U846 (N_846,In_239,In_393);
or U847 (N_847,In_253,In_226);
and U848 (N_848,In_226,In_138);
and U849 (N_849,In_258,In_8);
nor U850 (N_850,In_278,In_75);
nand U851 (N_851,In_236,In_348);
or U852 (N_852,In_217,In_485);
or U853 (N_853,In_275,In_463);
nand U854 (N_854,In_111,In_380);
nor U855 (N_855,In_137,In_282);
and U856 (N_856,In_33,In_332);
nor U857 (N_857,In_299,In_410);
nand U858 (N_858,In_143,In_408);
and U859 (N_859,In_399,In_280);
nor U860 (N_860,In_401,In_264);
and U861 (N_861,In_367,In_236);
nand U862 (N_862,In_396,In_235);
nand U863 (N_863,In_475,In_389);
or U864 (N_864,In_462,In_233);
and U865 (N_865,In_424,In_41);
nand U866 (N_866,In_145,In_321);
nor U867 (N_867,In_271,In_297);
nand U868 (N_868,In_415,In_353);
nor U869 (N_869,In_6,In_273);
nand U870 (N_870,In_410,In_357);
nand U871 (N_871,In_245,In_307);
nand U872 (N_872,In_76,In_445);
or U873 (N_873,In_183,In_145);
nand U874 (N_874,In_399,In_182);
nor U875 (N_875,In_217,In_9);
and U876 (N_876,In_339,In_283);
nand U877 (N_877,In_338,In_53);
nand U878 (N_878,In_304,In_308);
and U879 (N_879,In_14,In_364);
nor U880 (N_880,In_107,In_307);
nand U881 (N_881,In_236,In_444);
nor U882 (N_882,In_134,In_349);
nand U883 (N_883,In_220,In_384);
nor U884 (N_884,In_126,In_284);
and U885 (N_885,In_49,In_298);
or U886 (N_886,In_409,In_99);
nand U887 (N_887,In_100,In_353);
and U888 (N_888,In_286,In_271);
nand U889 (N_889,In_312,In_62);
nor U890 (N_890,In_111,In_145);
or U891 (N_891,In_60,In_257);
or U892 (N_892,In_88,In_18);
and U893 (N_893,In_477,In_9);
and U894 (N_894,In_201,In_231);
nor U895 (N_895,In_242,In_324);
and U896 (N_896,In_201,In_65);
nor U897 (N_897,In_103,In_73);
or U898 (N_898,In_18,In_223);
nand U899 (N_899,In_497,In_88);
nand U900 (N_900,In_202,In_402);
or U901 (N_901,In_297,In_214);
nand U902 (N_902,In_123,In_205);
nor U903 (N_903,In_289,In_94);
and U904 (N_904,In_328,In_285);
nor U905 (N_905,In_497,In_420);
nor U906 (N_906,In_425,In_466);
nor U907 (N_907,In_193,In_297);
nand U908 (N_908,In_6,In_475);
nand U909 (N_909,In_123,In_53);
or U910 (N_910,In_150,In_431);
or U911 (N_911,In_242,In_386);
nand U912 (N_912,In_457,In_64);
or U913 (N_913,In_47,In_18);
nand U914 (N_914,In_340,In_123);
nand U915 (N_915,In_149,In_163);
nand U916 (N_916,In_448,In_145);
and U917 (N_917,In_320,In_65);
nor U918 (N_918,In_309,In_1);
or U919 (N_919,In_401,In_307);
nor U920 (N_920,In_439,In_72);
and U921 (N_921,In_272,In_241);
nand U922 (N_922,In_292,In_105);
nor U923 (N_923,In_410,In_216);
and U924 (N_924,In_285,In_89);
and U925 (N_925,In_159,In_248);
nor U926 (N_926,In_375,In_270);
nand U927 (N_927,In_426,In_394);
nor U928 (N_928,In_429,In_206);
or U929 (N_929,In_86,In_31);
nor U930 (N_930,In_493,In_167);
or U931 (N_931,In_141,In_144);
nor U932 (N_932,In_311,In_190);
nor U933 (N_933,In_472,In_496);
nand U934 (N_934,In_422,In_95);
and U935 (N_935,In_243,In_464);
and U936 (N_936,In_25,In_48);
nand U937 (N_937,In_388,In_216);
nor U938 (N_938,In_449,In_204);
or U939 (N_939,In_478,In_332);
and U940 (N_940,In_40,In_482);
or U941 (N_941,In_127,In_282);
nand U942 (N_942,In_283,In_369);
or U943 (N_943,In_286,In_14);
and U944 (N_944,In_54,In_152);
and U945 (N_945,In_392,In_175);
nor U946 (N_946,In_109,In_152);
and U947 (N_947,In_271,In_456);
nand U948 (N_948,In_298,In_109);
and U949 (N_949,In_324,In_246);
or U950 (N_950,In_149,In_409);
and U951 (N_951,In_131,In_220);
nand U952 (N_952,In_68,In_452);
nand U953 (N_953,In_488,In_277);
or U954 (N_954,In_383,In_487);
and U955 (N_955,In_19,In_222);
and U956 (N_956,In_48,In_173);
nor U957 (N_957,In_354,In_342);
nand U958 (N_958,In_406,In_132);
xor U959 (N_959,In_125,In_287);
nor U960 (N_960,In_253,In_402);
and U961 (N_961,In_24,In_65);
or U962 (N_962,In_495,In_29);
or U963 (N_963,In_8,In_76);
and U964 (N_964,In_331,In_146);
nor U965 (N_965,In_266,In_323);
nand U966 (N_966,In_206,In_60);
and U967 (N_967,In_440,In_482);
or U968 (N_968,In_109,In_17);
or U969 (N_969,In_328,In_460);
nor U970 (N_970,In_434,In_56);
nor U971 (N_971,In_143,In_336);
and U972 (N_972,In_283,In_305);
or U973 (N_973,In_440,In_436);
nand U974 (N_974,In_336,In_264);
nand U975 (N_975,In_269,In_434);
nand U976 (N_976,In_10,In_301);
xor U977 (N_977,In_439,In_11);
or U978 (N_978,In_444,In_289);
and U979 (N_979,In_390,In_70);
nand U980 (N_980,In_12,In_122);
and U981 (N_981,In_197,In_277);
nor U982 (N_982,In_100,In_187);
or U983 (N_983,In_160,In_155);
or U984 (N_984,In_51,In_402);
or U985 (N_985,In_328,In_38);
and U986 (N_986,In_117,In_464);
nor U987 (N_987,In_119,In_183);
or U988 (N_988,In_433,In_96);
nor U989 (N_989,In_324,In_70);
xnor U990 (N_990,In_283,In_396);
or U991 (N_991,In_296,In_455);
nor U992 (N_992,In_274,In_70);
nor U993 (N_993,In_220,In_433);
and U994 (N_994,In_365,In_319);
nand U995 (N_995,In_293,In_64);
and U996 (N_996,In_371,In_70);
or U997 (N_997,In_476,In_63);
nor U998 (N_998,In_240,In_214);
and U999 (N_999,In_10,In_499);
nand U1000 (N_1000,N_5,N_312);
and U1001 (N_1001,N_494,N_245);
nor U1002 (N_1002,N_602,N_256);
nor U1003 (N_1003,N_615,N_448);
nor U1004 (N_1004,N_824,N_529);
or U1005 (N_1005,N_466,N_973);
or U1006 (N_1006,N_74,N_3);
or U1007 (N_1007,N_863,N_777);
or U1008 (N_1008,N_40,N_76);
or U1009 (N_1009,N_928,N_195);
nor U1010 (N_1010,N_301,N_349);
nand U1011 (N_1011,N_225,N_89);
and U1012 (N_1012,N_410,N_649);
nand U1013 (N_1013,N_443,N_482);
nor U1014 (N_1014,N_185,N_730);
nand U1015 (N_1015,N_621,N_158);
and U1016 (N_1016,N_627,N_542);
nor U1017 (N_1017,N_70,N_668);
and U1018 (N_1018,N_951,N_731);
or U1019 (N_1019,N_17,N_960);
nand U1020 (N_1020,N_884,N_120);
nor U1021 (N_1021,N_170,N_947);
or U1022 (N_1022,N_227,N_721);
nand U1023 (N_1023,N_313,N_452);
nand U1024 (N_1024,N_555,N_681);
nand U1025 (N_1025,N_561,N_893);
or U1026 (N_1026,N_530,N_861);
nand U1027 (N_1027,N_444,N_829);
nand U1028 (N_1028,N_100,N_849);
nor U1029 (N_1029,N_573,N_397);
nand U1030 (N_1030,N_98,N_140);
and U1031 (N_1031,N_696,N_125);
and U1032 (N_1032,N_648,N_867);
or U1033 (N_1033,N_713,N_577);
nor U1034 (N_1034,N_953,N_516);
or U1035 (N_1035,N_669,N_702);
and U1036 (N_1036,N_910,N_159);
and U1037 (N_1037,N_266,N_20);
nor U1038 (N_1038,N_436,N_331);
nor U1039 (N_1039,N_923,N_728);
and U1040 (N_1040,N_572,N_263);
nor U1041 (N_1041,N_678,N_854);
nor U1042 (N_1042,N_528,N_205);
and U1043 (N_1043,N_955,N_38);
and U1044 (N_1044,N_833,N_500);
and U1045 (N_1045,N_352,N_241);
and U1046 (N_1046,N_611,N_31);
or U1047 (N_1047,N_33,N_701);
or U1048 (N_1048,N_585,N_134);
xnor U1049 (N_1049,N_468,N_640);
nor U1050 (N_1050,N_624,N_243);
and U1051 (N_1051,N_168,N_109);
or U1052 (N_1052,N_543,N_575);
or U1053 (N_1053,N_985,N_920);
or U1054 (N_1054,N_49,N_71);
nor U1055 (N_1055,N_550,N_831);
or U1056 (N_1056,N_42,N_914);
nand U1057 (N_1057,N_576,N_972);
nor U1058 (N_1058,N_952,N_275);
nor U1059 (N_1059,N_683,N_509);
or U1060 (N_1060,N_641,N_59);
xor U1061 (N_1061,N_864,N_817);
nor U1062 (N_1062,N_161,N_870);
nand U1063 (N_1063,N_82,N_979);
and U1064 (N_1064,N_823,N_63);
and U1065 (N_1065,N_271,N_780);
and U1066 (N_1066,N_167,N_41);
and U1067 (N_1067,N_188,N_877);
and U1068 (N_1068,N_246,N_201);
and U1069 (N_1069,N_866,N_274);
nand U1070 (N_1070,N_321,N_44);
or U1071 (N_1071,N_768,N_304);
and U1072 (N_1072,N_704,N_138);
and U1073 (N_1073,N_881,N_811);
nand U1074 (N_1074,N_694,N_539);
nor U1075 (N_1075,N_19,N_191);
and U1076 (N_1076,N_607,N_414);
nor U1077 (N_1077,N_944,N_897);
and U1078 (N_1078,N_869,N_265);
nand U1079 (N_1079,N_693,N_463);
or U1080 (N_1080,N_868,N_395);
or U1081 (N_1081,N_359,N_236);
nor U1082 (N_1082,N_96,N_630);
nand U1083 (N_1083,N_318,N_93);
or U1084 (N_1084,N_909,N_233);
or U1085 (N_1085,N_420,N_422);
nor U1086 (N_1086,N_320,N_229);
and U1087 (N_1087,N_839,N_633);
or U1088 (N_1088,N_250,N_417);
nor U1089 (N_1089,N_548,N_628);
xnor U1090 (N_1090,N_386,N_964);
and U1091 (N_1091,N_806,N_652);
nand U1092 (N_1092,N_837,N_901);
xor U1093 (N_1093,N_355,N_257);
and U1094 (N_1094,N_921,N_828);
nand U1095 (N_1095,N_128,N_671);
or U1096 (N_1096,N_560,N_9);
nand U1097 (N_1097,N_559,N_978);
and U1098 (N_1098,N_112,N_378);
and U1099 (N_1099,N_315,N_270);
nand U1100 (N_1100,N_778,N_504);
nor U1101 (N_1101,N_200,N_916);
nand U1102 (N_1102,N_165,N_335);
nand U1103 (N_1103,N_298,N_157);
nor U1104 (N_1104,N_812,N_943);
nor U1105 (N_1105,N_458,N_799);
nor U1106 (N_1106,N_949,N_406);
or U1107 (N_1107,N_794,N_892);
nor U1108 (N_1108,N_84,N_154);
and U1109 (N_1109,N_58,N_450);
nand U1110 (N_1110,N_720,N_345);
and U1111 (N_1111,N_249,N_454);
nand U1112 (N_1112,N_589,N_83);
nand U1113 (N_1113,N_166,N_133);
nand U1114 (N_1114,N_363,N_691);
nand U1115 (N_1115,N_647,N_366);
nand U1116 (N_1116,N_551,N_805);
nor U1117 (N_1117,N_541,N_24);
or U1118 (N_1118,N_18,N_10);
nand U1119 (N_1119,N_217,N_762);
and U1120 (N_1120,N_342,N_663);
nand U1121 (N_1121,N_656,N_862);
nor U1122 (N_1122,N_264,N_710);
nand U1123 (N_1123,N_673,N_919);
or U1124 (N_1124,N_618,N_441);
or U1125 (N_1125,N_409,N_16);
or U1126 (N_1126,N_116,N_996);
or U1127 (N_1127,N_278,N_343);
nand U1128 (N_1128,N_876,N_171);
nor U1129 (N_1129,N_251,N_8);
nor U1130 (N_1130,N_103,N_723);
nand U1131 (N_1131,N_4,N_430);
nand U1132 (N_1132,N_418,N_334);
and U1133 (N_1133,N_603,N_660);
or U1134 (N_1134,N_685,N_958);
nor U1135 (N_1135,N_566,N_636);
or U1136 (N_1136,N_771,N_276);
nor U1137 (N_1137,N_362,N_204);
nor U1138 (N_1138,N_612,N_28);
or U1139 (N_1139,N_235,N_724);
nor U1140 (N_1140,N_507,N_287);
or U1141 (N_1141,N_369,N_294);
or U1142 (N_1142,N_101,N_259);
or U1143 (N_1143,N_609,N_725);
and U1144 (N_1144,N_825,N_476);
nand U1145 (N_1145,N_291,N_520);
xor U1146 (N_1146,N_495,N_485);
or U1147 (N_1147,N_986,N_108);
nand U1148 (N_1148,N_904,N_330);
or U1149 (N_1149,N_826,N_769);
or U1150 (N_1150,N_426,N_290);
or U1151 (N_1151,N_999,N_173);
nor U1152 (N_1152,N_481,N_186);
and U1153 (N_1153,N_906,N_992);
nand U1154 (N_1154,N_211,N_984);
nor U1155 (N_1155,N_965,N_682);
and U1156 (N_1156,N_997,N_709);
or U1157 (N_1157,N_122,N_809);
or U1158 (N_1158,N_324,N_908);
or U1159 (N_1159,N_638,N_107);
and U1160 (N_1160,N_853,N_323);
nand U1161 (N_1161,N_85,N_580);
nand U1162 (N_1162,N_765,N_586);
or U1163 (N_1163,N_364,N_929);
nand U1164 (N_1164,N_486,N_6);
nor U1165 (N_1165,N_948,N_78);
nand U1166 (N_1166,N_968,N_461);
and U1167 (N_1167,N_339,N_438);
nor U1168 (N_1168,N_353,N_68);
xnor U1169 (N_1169,N_501,N_48);
nand U1170 (N_1170,N_792,N_55);
and U1171 (N_1171,N_488,N_238);
or U1172 (N_1172,N_213,N_959);
nor U1173 (N_1173,N_686,N_514);
nor U1174 (N_1174,N_147,N_333);
and U1175 (N_1175,N_326,N_130);
nor U1176 (N_1176,N_309,N_797);
nor U1177 (N_1177,N_865,N_976);
nand U1178 (N_1178,N_900,N_684);
or U1179 (N_1179,N_385,N_961);
nor U1180 (N_1180,N_87,N_741);
nor U1181 (N_1181,N_889,N_727);
nand U1182 (N_1182,N_64,N_69);
or U1183 (N_1183,N_111,N_646);
and U1184 (N_1184,N_924,N_830);
or U1185 (N_1185,N_467,N_729);
nand U1186 (N_1186,N_350,N_408);
nor U1187 (N_1187,N_303,N_990);
or U1188 (N_1188,N_505,N_743);
nor U1189 (N_1189,N_759,N_433);
and U1190 (N_1190,N_88,N_493);
or U1191 (N_1191,N_616,N_478);
and U1192 (N_1192,N_12,N_153);
and U1193 (N_1193,N_600,N_155);
nor U1194 (N_1194,N_665,N_124);
and U1195 (N_1195,N_664,N_360);
or U1196 (N_1196,N_706,N_590);
or U1197 (N_1197,N_358,N_295);
nor U1198 (N_1198,N_524,N_570);
or U1199 (N_1199,N_22,N_855);
nand U1200 (N_1200,N_337,N_655);
or U1201 (N_1201,N_736,N_399);
and U1202 (N_1202,N_988,N_14);
and U1203 (N_1203,N_699,N_401);
nand U1204 (N_1204,N_405,N_617);
nand U1205 (N_1205,N_427,N_783);
nor U1206 (N_1206,N_581,N_781);
and U1207 (N_1207,N_610,N_564);
or U1208 (N_1208,N_196,N_286);
nor U1209 (N_1209,N_926,N_383);
or U1210 (N_1210,N_605,N_393);
or U1211 (N_1211,N_712,N_974);
nand U1212 (N_1212,N_941,N_898);
nor U1213 (N_1213,N_372,N_565);
nor U1214 (N_1214,N_894,N_136);
nor U1215 (N_1215,N_65,N_925);
nand U1216 (N_1216,N_273,N_808);
nand U1217 (N_1217,N_875,N_105);
or U1218 (N_1218,N_172,N_832);
nor U1219 (N_1219,N_651,N_54);
and U1220 (N_1220,N_689,N_472);
nand U1221 (N_1221,N_492,N_86);
nor U1222 (N_1222,N_767,N_29);
and U1223 (N_1223,N_761,N_643);
nor U1224 (N_1224,N_141,N_625);
and U1225 (N_1225,N_356,N_338);
or U1226 (N_1226,N_25,N_460);
or U1227 (N_1227,N_178,N_989);
xor U1228 (N_1228,N_253,N_766);
or U1229 (N_1229,N_873,N_796);
or U1230 (N_1230,N_2,N_774);
nand U1231 (N_1231,N_626,N_842);
or U1232 (N_1232,N_786,N_740);
xnor U1233 (N_1233,N_822,N_240);
nor U1234 (N_1234,N_179,N_584);
and U1235 (N_1235,N_465,N_770);
nand U1236 (N_1236,N_162,N_735);
or U1237 (N_1237,N_991,N_659);
nand U1238 (N_1238,N_148,N_527);
or U1239 (N_1239,N_834,N_593);
nor U1240 (N_1240,N_549,N_432);
nor U1241 (N_1241,N_289,N_695);
nor U1242 (N_1242,N_578,N_174);
or U1243 (N_1243,N_252,N_690);
nor U1244 (N_1244,N_187,N_517);
and U1245 (N_1245,N_887,N_428);
nand U1246 (N_1246,N_208,N_747);
and U1247 (N_1247,N_567,N_885);
nand U1248 (N_1248,N_558,N_341);
nor U1249 (N_1249,N_732,N_160);
nor U1250 (N_1250,N_840,N_32);
nor U1251 (N_1251,N_202,N_579);
nand U1252 (N_1252,N_674,N_95);
nor U1253 (N_1253,N_305,N_742);
and U1254 (N_1254,N_218,N_242);
or U1255 (N_1255,N_221,N_431);
and U1256 (N_1256,N_917,N_970);
nand U1257 (N_1257,N_11,N_282);
or U1258 (N_1258,N_679,N_471);
nor U1259 (N_1259,N_637,N_224);
and U1260 (N_1260,N_222,N_220);
and U1261 (N_1261,N_554,N_176);
or U1262 (N_1262,N_268,N_94);
and U1263 (N_1263,N_526,N_599);
and U1264 (N_1264,N_571,N_39);
and U1265 (N_1265,N_857,N_272);
and U1266 (N_1266,N_677,N_503);
and U1267 (N_1267,N_934,N_977);
and U1268 (N_1268,N_895,N_368);
or U1269 (N_1269,N_911,N_110);
nor U1270 (N_1270,N_882,N_963);
nand U1271 (N_1271,N_307,N_464);
or U1272 (N_1272,N_546,N_814);
or U1273 (N_1273,N_27,N_905);
and U1274 (N_1274,N_123,N_328);
or U1275 (N_1275,N_446,N_316);
and U1276 (N_1276,N_143,N_206);
nand U1277 (N_1277,N_102,N_403);
nand U1278 (N_1278,N_210,N_36);
nor U1279 (N_1279,N_545,N_818);
nor U1280 (N_1280,N_827,N_595);
nand U1281 (N_1281,N_254,N_614);
xnor U1282 (N_1282,N_511,N_491);
and U1283 (N_1283,N_670,N_180);
nand U1284 (N_1284,N_795,N_456);
and U1285 (N_1285,N_714,N_707);
and U1286 (N_1286,N_697,N_469);
nor U1287 (N_1287,N_874,N_300);
nand U1288 (N_1288,N_594,N_810);
and U1289 (N_1289,N_962,N_447);
nand U1290 (N_1290,N_751,N_623);
nand U1291 (N_1291,N_361,N_214);
nand U1292 (N_1292,N_135,N_622);
nor U1293 (N_1293,N_223,N_975);
nor U1294 (N_1294,N_878,N_513);
and U1295 (N_1295,N_568,N_376);
nor U1296 (N_1296,N_888,N_329);
nand U1297 (N_1297,N_645,N_932);
and U1298 (N_1298,N_680,N_987);
nor U1299 (N_1299,N_308,N_692);
or U1300 (N_1300,N_336,N_969);
nand U1301 (N_1301,N_983,N_480);
nand U1302 (N_1302,N_498,N_203);
or U1303 (N_1303,N_804,N_382);
nand U1304 (N_1304,N_424,N_700);
or U1305 (N_1305,N_152,N_748);
or U1306 (N_1306,N_502,N_587);
nor U1307 (N_1307,N_15,N_247);
or U1308 (N_1308,N_119,N_474);
nor U1309 (N_1309,N_193,N_995);
xor U1310 (N_1310,N_930,N_705);
nor U1311 (N_1311,N_175,N_421);
nor U1312 (N_1312,N_606,N_752);
nand U1313 (N_1313,N_299,N_588);
nand U1314 (N_1314,N_980,N_145);
nand U1315 (N_1315,N_62,N_556);
and U1316 (N_1316,N_733,N_262);
or U1317 (N_1317,N_91,N_197);
nor U1318 (N_1318,N_288,N_856);
and U1319 (N_1319,N_104,N_234);
nor U1320 (N_1320,N_788,N_327);
nor U1321 (N_1321,N_499,N_845);
nand U1322 (N_1322,N_35,N_45);
nor U1323 (N_1323,N_230,N_667);
and U1324 (N_1324,N_370,N_902);
nand U1325 (N_1325,N_1,N_387);
xnor U1326 (N_1326,N_785,N_97);
and U1327 (N_1327,N_411,N_150);
nand U1328 (N_1328,N_657,N_412);
xor U1329 (N_1329,N_228,N_820);
and U1330 (N_1330,N_532,N_891);
nor U1331 (N_1331,N_843,N_199);
nor U1332 (N_1332,N_484,N_592);
and U1333 (N_1333,N_755,N_760);
nor U1334 (N_1334,N_381,N_90);
or U1335 (N_1335,N_544,N_192);
or U1336 (N_1336,N_407,N_244);
or U1337 (N_1337,N_672,N_413);
nand U1338 (N_1338,N_872,N_716);
or U1339 (N_1339,N_813,N_791);
or U1340 (N_1340,N_838,N_151);
or U1341 (N_1341,N_675,N_890);
nand U1342 (N_1342,N_763,N_896);
nand U1343 (N_1343,N_92,N_114);
nor U1344 (N_1344,N_574,N_429);
or U1345 (N_1345,N_131,N_455);
nand U1346 (N_1346,N_956,N_753);
nand U1347 (N_1347,N_757,N_922);
and U1348 (N_1348,N_604,N_237);
nand U1349 (N_1349,N_666,N_142);
nand U1350 (N_1350,N_519,N_189);
nor U1351 (N_1351,N_547,N_722);
nor U1352 (N_1352,N_277,N_184);
nor U1353 (N_1353,N_129,N_787);
or U1354 (N_1354,N_53,N_982);
nand U1355 (N_1355,N_190,N_37);
nand U1356 (N_1356,N_435,N_164);
nand U1357 (N_1357,N_879,N_538);
and U1358 (N_1358,N_521,N_779);
or U1359 (N_1359,N_357,N_81);
nand U1360 (N_1360,N_703,N_931);
and U1361 (N_1361,N_942,N_23);
nor U1362 (N_1362,N_297,N_182);
and U1363 (N_1363,N_782,N_310);
and U1364 (N_1364,N_351,N_60);
or U1365 (N_1365,N_613,N_676);
or U1366 (N_1366,N_967,N_739);
nor U1367 (N_1367,N_7,N_13);
and U1368 (N_1368,N_216,N_749);
or U1369 (N_1369,N_231,N_354);
or U1370 (N_1370,N_852,N_30);
nand U1371 (N_1371,N_149,N_496);
nand U1372 (N_1372,N_591,N_394);
or U1373 (N_1373,N_423,N_416);
nor U1374 (N_1374,N_841,N_440);
and U1375 (N_1375,N_525,N_425);
and U1376 (N_1376,N_402,N_391);
nand U1377 (N_1377,N_293,N_198);
or U1378 (N_1378,N_708,N_118);
nor U1379 (N_1379,N_283,N_404);
nor U1380 (N_1380,N_859,N_515);
and U1381 (N_1381,N_181,N_661);
or U1382 (N_1382,N_207,N_169);
nand U1383 (N_1383,N_523,N_746);
and U1384 (N_1384,N_209,N_798);
nand U1385 (N_1385,N_819,N_937);
nand U1386 (N_1386,N_535,N_292);
xor U1387 (N_1387,N_415,N_620);
and U1388 (N_1388,N_775,N_284);
or U1389 (N_1389,N_377,N_583);
nand U1390 (N_1390,N_536,N_99);
and U1391 (N_1391,N_936,N_445);
and U1392 (N_1392,N_380,N_314);
nand U1393 (N_1393,N_629,N_886);
and U1394 (N_1394,N_106,N_601);
nand U1395 (N_1395,N_457,N_899);
or U1396 (N_1396,N_177,N_57);
nand U1397 (N_1397,N_927,N_533);
nor U1398 (N_1398,N_772,N_137);
or U1399 (N_1399,N_113,N_258);
nand U1400 (N_1400,N_490,N_758);
or U1401 (N_1401,N_800,N_437);
and U1402 (N_1402,N_510,N_390);
or U1403 (N_1403,N_47,N_255);
nor U1404 (N_1404,N_994,N_365);
and U1405 (N_1405,N_43,N_654);
nor U1406 (N_1406,N_537,N_719);
nor U1407 (N_1407,N_711,N_726);
and U1408 (N_1408,N_462,N_50);
or U1409 (N_1409,N_642,N_619);
nor U1410 (N_1410,N_913,N_608);
nand U1411 (N_1411,N_698,N_453);
or U1412 (N_1412,N_156,N_325);
nor U1413 (N_1413,N_497,N_21);
and U1414 (N_1414,N_398,N_860);
nand U1415 (N_1415,N_718,N_67);
and U1416 (N_1416,N_261,N_632);
and U1417 (N_1417,N_522,N_346);
or U1418 (N_1418,N_658,N_569);
and U1419 (N_1419,N_553,N_734);
or U1420 (N_1420,N_596,N_80);
nand U1421 (N_1421,N_844,N_552);
nand U1422 (N_1422,N_46,N_597);
nor U1423 (N_1423,N_449,N_793);
or U1424 (N_1424,N_846,N_851);
nand U1425 (N_1425,N_939,N_194);
nor U1426 (N_1426,N_993,N_880);
or U1427 (N_1427,N_801,N_802);
nor U1428 (N_1428,N_248,N_562);
and U1429 (N_1429,N_379,N_850);
nor U1430 (N_1430,N_506,N_650);
nor U1431 (N_1431,N_836,N_915);
nor U1432 (N_1432,N_764,N_56);
and U1433 (N_1433,N_470,N_434);
nor U1434 (N_1434,N_479,N_477);
and U1435 (N_1435,N_61,N_0);
nand U1436 (N_1436,N_938,N_717);
and U1437 (N_1437,N_688,N_871);
nand U1438 (N_1438,N_912,N_302);
or U1439 (N_1439,N_419,N_508);
nand U1440 (N_1440,N_212,N_392);
nor U1441 (N_1441,N_907,N_738);
or U1442 (N_1442,N_639,N_998);
or U1443 (N_1443,N_489,N_306);
nand U1444 (N_1444,N_807,N_634);
nand U1445 (N_1445,N_971,N_945);
and U1446 (N_1446,N_183,N_531);
nor U1447 (N_1447,N_750,N_340);
nor U1448 (N_1448,N_582,N_375);
nor U1449 (N_1449,N_483,N_512);
and U1450 (N_1450,N_127,N_439);
nand U1451 (N_1451,N_957,N_773);
and U1452 (N_1452,N_144,N_784);
and U1453 (N_1453,N_239,N_459);
nor U1454 (N_1454,N_662,N_146);
and U1455 (N_1455,N_267,N_117);
nand U1456 (N_1456,N_946,N_598);
nor U1457 (N_1457,N_487,N_821);
or U1458 (N_1458,N_317,N_26);
nand U1459 (N_1459,N_348,N_715);
and U1460 (N_1460,N_557,N_66);
or U1461 (N_1461,N_371,N_121);
and U1462 (N_1462,N_373,N_776);
nor U1463 (N_1463,N_396,N_954);
or U1464 (N_1464,N_280,N_139);
nand U1465 (N_1465,N_835,N_744);
nor U1466 (N_1466,N_226,N_789);
and U1467 (N_1467,N_347,N_933);
and U1468 (N_1468,N_966,N_790);
and U1469 (N_1469,N_756,N_737);
or U1470 (N_1470,N_848,N_260);
nor U1471 (N_1471,N_374,N_126);
or U1472 (N_1472,N_311,N_803);
and U1473 (N_1473,N_815,N_389);
xnor U1474 (N_1474,N_883,N_34);
and U1475 (N_1475,N_644,N_232);
nand U1476 (N_1476,N_319,N_442);
and U1477 (N_1477,N_279,N_132);
xor U1478 (N_1478,N_754,N_653);
or U1479 (N_1479,N_475,N_847);
or U1480 (N_1480,N_816,N_631);
and U1481 (N_1481,N_858,N_79);
nor U1482 (N_1482,N_281,N_563);
nand U1483 (N_1483,N_51,N_115);
nor U1484 (N_1484,N_296,N_73);
nand U1485 (N_1485,N_451,N_473);
and U1486 (N_1486,N_540,N_332);
nand U1487 (N_1487,N_285,N_269);
nor U1488 (N_1488,N_950,N_687);
nand U1489 (N_1489,N_745,N_77);
or U1490 (N_1490,N_344,N_981);
nor U1491 (N_1491,N_534,N_903);
or U1492 (N_1492,N_384,N_72);
nand U1493 (N_1493,N_219,N_388);
or U1494 (N_1494,N_75,N_367);
and U1495 (N_1495,N_322,N_400);
nand U1496 (N_1496,N_635,N_52);
and U1497 (N_1497,N_163,N_935);
nand U1498 (N_1498,N_940,N_918);
nand U1499 (N_1499,N_215,N_518);
nor U1500 (N_1500,N_844,N_349);
nor U1501 (N_1501,N_213,N_319);
nand U1502 (N_1502,N_243,N_61);
nor U1503 (N_1503,N_251,N_203);
nor U1504 (N_1504,N_339,N_887);
or U1505 (N_1505,N_500,N_62);
and U1506 (N_1506,N_810,N_310);
nor U1507 (N_1507,N_592,N_483);
and U1508 (N_1508,N_455,N_433);
and U1509 (N_1509,N_321,N_634);
nand U1510 (N_1510,N_292,N_174);
nor U1511 (N_1511,N_767,N_349);
nor U1512 (N_1512,N_113,N_348);
or U1513 (N_1513,N_362,N_956);
and U1514 (N_1514,N_161,N_828);
or U1515 (N_1515,N_75,N_162);
nor U1516 (N_1516,N_394,N_578);
or U1517 (N_1517,N_916,N_341);
or U1518 (N_1518,N_447,N_275);
or U1519 (N_1519,N_947,N_640);
nor U1520 (N_1520,N_185,N_800);
or U1521 (N_1521,N_12,N_464);
and U1522 (N_1522,N_15,N_663);
nand U1523 (N_1523,N_91,N_241);
nor U1524 (N_1524,N_160,N_673);
nor U1525 (N_1525,N_766,N_42);
and U1526 (N_1526,N_954,N_477);
and U1527 (N_1527,N_257,N_926);
and U1528 (N_1528,N_523,N_255);
or U1529 (N_1529,N_248,N_92);
nand U1530 (N_1530,N_487,N_534);
and U1531 (N_1531,N_354,N_194);
and U1532 (N_1532,N_888,N_151);
and U1533 (N_1533,N_340,N_681);
and U1534 (N_1534,N_614,N_692);
nand U1535 (N_1535,N_670,N_799);
and U1536 (N_1536,N_222,N_368);
nor U1537 (N_1537,N_105,N_734);
and U1538 (N_1538,N_403,N_21);
nor U1539 (N_1539,N_254,N_495);
nor U1540 (N_1540,N_50,N_289);
and U1541 (N_1541,N_105,N_316);
nor U1542 (N_1542,N_837,N_435);
or U1543 (N_1543,N_835,N_858);
nand U1544 (N_1544,N_255,N_315);
nor U1545 (N_1545,N_334,N_683);
nor U1546 (N_1546,N_274,N_409);
or U1547 (N_1547,N_892,N_292);
or U1548 (N_1548,N_829,N_463);
nor U1549 (N_1549,N_538,N_99);
nand U1550 (N_1550,N_593,N_439);
or U1551 (N_1551,N_264,N_98);
and U1552 (N_1552,N_533,N_257);
nand U1553 (N_1553,N_295,N_190);
or U1554 (N_1554,N_833,N_521);
nor U1555 (N_1555,N_200,N_756);
or U1556 (N_1556,N_950,N_612);
and U1557 (N_1557,N_453,N_325);
nand U1558 (N_1558,N_828,N_922);
or U1559 (N_1559,N_421,N_235);
nand U1560 (N_1560,N_971,N_788);
nor U1561 (N_1561,N_539,N_806);
and U1562 (N_1562,N_700,N_259);
nand U1563 (N_1563,N_714,N_551);
nor U1564 (N_1564,N_123,N_526);
nand U1565 (N_1565,N_815,N_45);
or U1566 (N_1566,N_805,N_250);
or U1567 (N_1567,N_332,N_311);
nand U1568 (N_1568,N_339,N_42);
nand U1569 (N_1569,N_840,N_662);
nor U1570 (N_1570,N_627,N_183);
xor U1571 (N_1571,N_648,N_298);
nand U1572 (N_1572,N_426,N_297);
or U1573 (N_1573,N_823,N_894);
or U1574 (N_1574,N_157,N_486);
or U1575 (N_1575,N_870,N_104);
and U1576 (N_1576,N_555,N_219);
and U1577 (N_1577,N_565,N_177);
and U1578 (N_1578,N_172,N_147);
or U1579 (N_1579,N_299,N_40);
and U1580 (N_1580,N_674,N_337);
and U1581 (N_1581,N_189,N_987);
nor U1582 (N_1582,N_689,N_756);
nor U1583 (N_1583,N_598,N_427);
nand U1584 (N_1584,N_288,N_940);
nor U1585 (N_1585,N_739,N_906);
or U1586 (N_1586,N_64,N_824);
nand U1587 (N_1587,N_239,N_736);
or U1588 (N_1588,N_295,N_210);
and U1589 (N_1589,N_621,N_453);
nand U1590 (N_1590,N_170,N_422);
or U1591 (N_1591,N_163,N_589);
or U1592 (N_1592,N_295,N_6);
nor U1593 (N_1593,N_622,N_901);
nor U1594 (N_1594,N_262,N_922);
nand U1595 (N_1595,N_529,N_142);
and U1596 (N_1596,N_793,N_392);
and U1597 (N_1597,N_314,N_940);
nand U1598 (N_1598,N_585,N_235);
nand U1599 (N_1599,N_941,N_915);
or U1600 (N_1600,N_63,N_976);
nand U1601 (N_1601,N_337,N_414);
or U1602 (N_1602,N_589,N_230);
nand U1603 (N_1603,N_691,N_789);
and U1604 (N_1604,N_553,N_210);
nand U1605 (N_1605,N_714,N_112);
nor U1606 (N_1606,N_397,N_923);
nand U1607 (N_1607,N_533,N_250);
and U1608 (N_1608,N_592,N_354);
or U1609 (N_1609,N_164,N_898);
xnor U1610 (N_1610,N_897,N_838);
nor U1611 (N_1611,N_754,N_636);
and U1612 (N_1612,N_106,N_241);
nand U1613 (N_1613,N_794,N_66);
and U1614 (N_1614,N_541,N_744);
nand U1615 (N_1615,N_665,N_223);
and U1616 (N_1616,N_274,N_537);
and U1617 (N_1617,N_343,N_826);
and U1618 (N_1618,N_913,N_689);
and U1619 (N_1619,N_540,N_834);
and U1620 (N_1620,N_327,N_663);
nand U1621 (N_1621,N_873,N_465);
and U1622 (N_1622,N_387,N_834);
nand U1623 (N_1623,N_605,N_178);
or U1624 (N_1624,N_432,N_981);
and U1625 (N_1625,N_307,N_850);
and U1626 (N_1626,N_876,N_222);
nor U1627 (N_1627,N_270,N_99);
and U1628 (N_1628,N_621,N_620);
or U1629 (N_1629,N_341,N_452);
or U1630 (N_1630,N_356,N_336);
xor U1631 (N_1631,N_273,N_435);
nand U1632 (N_1632,N_965,N_707);
nor U1633 (N_1633,N_306,N_303);
nor U1634 (N_1634,N_564,N_322);
or U1635 (N_1635,N_298,N_159);
or U1636 (N_1636,N_858,N_472);
nand U1637 (N_1637,N_654,N_268);
nand U1638 (N_1638,N_415,N_482);
or U1639 (N_1639,N_935,N_787);
nor U1640 (N_1640,N_836,N_228);
nor U1641 (N_1641,N_566,N_830);
nor U1642 (N_1642,N_886,N_193);
and U1643 (N_1643,N_391,N_772);
or U1644 (N_1644,N_538,N_275);
nor U1645 (N_1645,N_257,N_563);
nand U1646 (N_1646,N_765,N_766);
nor U1647 (N_1647,N_385,N_943);
nor U1648 (N_1648,N_6,N_56);
or U1649 (N_1649,N_3,N_246);
nor U1650 (N_1650,N_613,N_152);
nor U1651 (N_1651,N_865,N_831);
nor U1652 (N_1652,N_152,N_883);
or U1653 (N_1653,N_736,N_692);
nor U1654 (N_1654,N_571,N_204);
or U1655 (N_1655,N_407,N_804);
and U1656 (N_1656,N_66,N_648);
nor U1657 (N_1657,N_826,N_254);
and U1658 (N_1658,N_714,N_151);
or U1659 (N_1659,N_749,N_561);
nand U1660 (N_1660,N_350,N_0);
nand U1661 (N_1661,N_139,N_71);
nand U1662 (N_1662,N_650,N_275);
or U1663 (N_1663,N_215,N_113);
nand U1664 (N_1664,N_443,N_992);
and U1665 (N_1665,N_535,N_506);
or U1666 (N_1666,N_179,N_127);
nand U1667 (N_1667,N_353,N_713);
nor U1668 (N_1668,N_535,N_510);
nand U1669 (N_1669,N_723,N_399);
and U1670 (N_1670,N_501,N_356);
and U1671 (N_1671,N_388,N_393);
or U1672 (N_1672,N_943,N_62);
and U1673 (N_1673,N_685,N_768);
nor U1674 (N_1674,N_789,N_545);
or U1675 (N_1675,N_258,N_333);
nand U1676 (N_1676,N_346,N_915);
or U1677 (N_1677,N_989,N_472);
xor U1678 (N_1678,N_420,N_595);
or U1679 (N_1679,N_729,N_682);
or U1680 (N_1680,N_834,N_648);
nand U1681 (N_1681,N_753,N_919);
or U1682 (N_1682,N_471,N_374);
or U1683 (N_1683,N_806,N_59);
or U1684 (N_1684,N_454,N_990);
and U1685 (N_1685,N_153,N_143);
nor U1686 (N_1686,N_606,N_549);
or U1687 (N_1687,N_74,N_411);
and U1688 (N_1688,N_360,N_834);
nand U1689 (N_1689,N_342,N_337);
or U1690 (N_1690,N_223,N_400);
and U1691 (N_1691,N_186,N_697);
and U1692 (N_1692,N_595,N_219);
nor U1693 (N_1693,N_842,N_404);
or U1694 (N_1694,N_368,N_269);
nand U1695 (N_1695,N_361,N_882);
or U1696 (N_1696,N_915,N_991);
and U1697 (N_1697,N_837,N_360);
and U1698 (N_1698,N_298,N_190);
nor U1699 (N_1699,N_714,N_457);
and U1700 (N_1700,N_753,N_982);
nand U1701 (N_1701,N_293,N_626);
and U1702 (N_1702,N_814,N_517);
nand U1703 (N_1703,N_957,N_852);
nand U1704 (N_1704,N_518,N_637);
nor U1705 (N_1705,N_638,N_464);
nand U1706 (N_1706,N_680,N_121);
nand U1707 (N_1707,N_338,N_962);
and U1708 (N_1708,N_645,N_934);
and U1709 (N_1709,N_127,N_119);
or U1710 (N_1710,N_755,N_753);
nand U1711 (N_1711,N_14,N_123);
or U1712 (N_1712,N_47,N_894);
nor U1713 (N_1713,N_196,N_103);
and U1714 (N_1714,N_86,N_930);
nor U1715 (N_1715,N_291,N_789);
and U1716 (N_1716,N_164,N_716);
nand U1717 (N_1717,N_734,N_402);
nand U1718 (N_1718,N_274,N_374);
or U1719 (N_1719,N_697,N_654);
nand U1720 (N_1720,N_63,N_489);
and U1721 (N_1721,N_746,N_618);
nor U1722 (N_1722,N_656,N_727);
nand U1723 (N_1723,N_478,N_27);
nor U1724 (N_1724,N_413,N_603);
nand U1725 (N_1725,N_694,N_818);
nor U1726 (N_1726,N_351,N_781);
and U1727 (N_1727,N_480,N_912);
or U1728 (N_1728,N_957,N_355);
nand U1729 (N_1729,N_558,N_565);
and U1730 (N_1730,N_524,N_748);
nor U1731 (N_1731,N_559,N_222);
nand U1732 (N_1732,N_311,N_282);
or U1733 (N_1733,N_250,N_772);
xnor U1734 (N_1734,N_851,N_941);
nor U1735 (N_1735,N_230,N_96);
or U1736 (N_1736,N_970,N_101);
nand U1737 (N_1737,N_437,N_871);
nand U1738 (N_1738,N_617,N_756);
nand U1739 (N_1739,N_125,N_737);
or U1740 (N_1740,N_392,N_625);
nand U1741 (N_1741,N_303,N_740);
nor U1742 (N_1742,N_433,N_336);
and U1743 (N_1743,N_30,N_281);
and U1744 (N_1744,N_876,N_595);
nor U1745 (N_1745,N_456,N_835);
nand U1746 (N_1746,N_321,N_707);
nor U1747 (N_1747,N_401,N_285);
nand U1748 (N_1748,N_965,N_869);
nand U1749 (N_1749,N_618,N_279);
nor U1750 (N_1750,N_326,N_676);
nand U1751 (N_1751,N_971,N_531);
and U1752 (N_1752,N_423,N_151);
and U1753 (N_1753,N_596,N_213);
and U1754 (N_1754,N_973,N_446);
and U1755 (N_1755,N_198,N_500);
and U1756 (N_1756,N_648,N_790);
or U1757 (N_1757,N_901,N_227);
and U1758 (N_1758,N_282,N_731);
nor U1759 (N_1759,N_236,N_750);
and U1760 (N_1760,N_94,N_656);
nor U1761 (N_1761,N_403,N_841);
nor U1762 (N_1762,N_31,N_949);
and U1763 (N_1763,N_763,N_231);
and U1764 (N_1764,N_780,N_947);
and U1765 (N_1765,N_123,N_989);
nor U1766 (N_1766,N_748,N_199);
nor U1767 (N_1767,N_742,N_435);
nand U1768 (N_1768,N_310,N_342);
or U1769 (N_1769,N_115,N_612);
and U1770 (N_1770,N_735,N_189);
nand U1771 (N_1771,N_633,N_445);
or U1772 (N_1772,N_694,N_504);
and U1773 (N_1773,N_279,N_931);
nor U1774 (N_1774,N_255,N_835);
nor U1775 (N_1775,N_199,N_859);
nor U1776 (N_1776,N_425,N_782);
or U1777 (N_1777,N_225,N_539);
nor U1778 (N_1778,N_980,N_237);
and U1779 (N_1779,N_145,N_408);
and U1780 (N_1780,N_109,N_575);
nor U1781 (N_1781,N_764,N_29);
or U1782 (N_1782,N_263,N_235);
nor U1783 (N_1783,N_27,N_399);
and U1784 (N_1784,N_825,N_865);
nor U1785 (N_1785,N_213,N_548);
or U1786 (N_1786,N_202,N_496);
nor U1787 (N_1787,N_66,N_979);
nor U1788 (N_1788,N_365,N_765);
and U1789 (N_1789,N_732,N_33);
or U1790 (N_1790,N_733,N_989);
nand U1791 (N_1791,N_819,N_812);
nand U1792 (N_1792,N_321,N_48);
or U1793 (N_1793,N_84,N_709);
nand U1794 (N_1794,N_428,N_596);
or U1795 (N_1795,N_755,N_283);
or U1796 (N_1796,N_469,N_998);
nor U1797 (N_1797,N_249,N_371);
and U1798 (N_1798,N_374,N_418);
and U1799 (N_1799,N_628,N_343);
or U1800 (N_1800,N_116,N_487);
nor U1801 (N_1801,N_780,N_299);
and U1802 (N_1802,N_978,N_683);
or U1803 (N_1803,N_76,N_824);
or U1804 (N_1804,N_640,N_649);
and U1805 (N_1805,N_146,N_633);
or U1806 (N_1806,N_147,N_897);
nand U1807 (N_1807,N_191,N_792);
nand U1808 (N_1808,N_565,N_133);
and U1809 (N_1809,N_713,N_674);
and U1810 (N_1810,N_453,N_953);
nand U1811 (N_1811,N_43,N_572);
and U1812 (N_1812,N_304,N_87);
and U1813 (N_1813,N_954,N_296);
or U1814 (N_1814,N_105,N_483);
and U1815 (N_1815,N_793,N_893);
or U1816 (N_1816,N_146,N_239);
nand U1817 (N_1817,N_151,N_63);
or U1818 (N_1818,N_802,N_302);
nand U1819 (N_1819,N_654,N_954);
and U1820 (N_1820,N_706,N_540);
nor U1821 (N_1821,N_723,N_919);
nand U1822 (N_1822,N_318,N_888);
and U1823 (N_1823,N_9,N_586);
nor U1824 (N_1824,N_375,N_105);
nand U1825 (N_1825,N_940,N_623);
or U1826 (N_1826,N_702,N_47);
nor U1827 (N_1827,N_308,N_141);
or U1828 (N_1828,N_298,N_690);
and U1829 (N_1829,N_617,N_312);
and U1830 (N_1830,N_341,N_866);
nor U1831 (N_1831,N_617,N_930);
nor U1832 (N_1832,N_559,N_593);
and U1833 (N_1833,N_321,N_859);
or U1834 (N_1834,N_263,N_421);
or U1835 (N_1835,N_430,N_469);
or U1836 (N_1836,N_831,N_583);
nand U1837 (N_1837,N_564,N_445);
nor U1838 (N_1838,N_928,N_336);
and U1839 (N_1839,N_175,N_92);
nor U1840 (N_1840,N_809,N_801);
nor U1841 (N_1841,N_280,N_463);
nand U1842 (N_1842,N_833,N_990);
or U1843 (N_1843,N_694,N_321);
or U1844 (N_1844,N_608,N_227);
or U1845 (N_1845,N_385,N_364);
and U1846 (N_1846,N_217,N_613);
nor U1847 (N_1847,N_31,N_206);
and U1848 (N_1848,N_777,N_990);
nand U1849 (N_1849,N_764,N_397);
and U1850 (N_1850,N_218,N_441);
and U1851 (N_1851,N_404,N_611);
nor U1852 (N_1852,N_371,N_542);
and U1853 (N_1853,N_296,N_866);
and U1854 (N_1854,N_909,N_852);
nand U1855 (N_1855,N_892,N_248);
nor U1856 (N_1856,N_771,N_420);
or U1857 (N_1857,N_666,N_672);
or U1858 (N_1858,N_504,N_254);
nand U1859 (N_1859,N_187,N_379);
nor U1860 (N_1860,N_948,N_828);
nand U1861 (N_1861,N_659,N_547);
and U1862 (N_1862,N_382,N_583);
nor U1863 (N_1863,N_194,N_836);
nor U1864 (N_1864,N_466,N_344);
nand U1865 (N_1865,N_705,N_351);
or U1866 (N_1866,N_350,N_670);
and U1867 (N_1867,N_544,N_178);
or U1868 (N_1868,N_319,N_638);
or U1869 (N_1869,N_15,N_455);
nand U1870 (N_1870,N_732,N_555);
nor U1871 (N_1871,N_332,N_776);
and U1872 (N_1872,N_800,N_883);
nand U1873 (N_1873,N_25,N_154);
or U1874 (N_1874,N_856,N_619);
or U1875 (N_1875,N_397,N_497);
and U1876 (N_1876,N_81,N_871);
or U1877 (N_1877,N_917,N_526);
and U1878 (N_1878,N_395,N_128);
nor U1879 (N_1879,N_892,N_271);
and U1880 (N_1880,N_479,N_605);
or U1881 (N_1881,N_848,N_275);
nor U1882 (N_1882,N_251,N_545);
nor U1883 (N_1883,N_190,N_121);
nand U1884 (N_1884,N_700,N_627);
or U1885 (N_1885,N_297,N_296);
xor U1886 (N_1886,N_677,N_371);
and U1887 (N_1887,N_679,N_952);
or U1888 (N_1888,N_777,N_928);
nor U1889 (N_1889,N_929,N_998);
and U1890 (N_1890,N_19,N_566);
nor U1891 (N_1891,N_672,N_91);
nand U1892 (N_1892,N_412,N_430);
nand U1893 (N_1893,N_643,N_321);
nor U1894 (N_1894,N_586,N_12);
or U1895 (N_1895,N_781,N_404);
and U1896 (N_1896,N_49,N_422);
or U1897 (N_1897,N_909,N_360);
nor U1898 (N_1898,N_860,N_902);
or U1899 (N_1899,N_551,N_381);
and U1900 (N_1900,N_45,N_984);
nor U1901 (N_1901,N_9,N_378);
and U1902 (N_1902,N_111,N_28);
and U1903 (N_1903,N_456,N_450);
and U1904 (N_1904,N_258,N_316);
or U1905 (N_1905,N_132,N_830);
nor U1906 (N_1906,N_990,N_398);
and U1907 (N_1907,N_200,N_227);
nand U1908 (N_1908,N_178,N_598);
nor U1909 (N_1909,N_150,N_519);
nor U1910 (N_1910,N_828,N_265);
nor U1911 (N_1911,N_955,N_771);
nor U1912 (N_1912,N_488,N_359);
nor U1913 (N_1913,N_994,N_448);
nor U1914 (N_1914,N_573,N_946);
and U1915 (N_1915,N_319,N_470);
nand U1916 (N_1916,N_813,N_79);
nand U1917 (N_1917,N_919,N_475);
nor U1918 (N_1918,N_793,N_989);
or U1919 (N_1919,N_416,N_188);
or U1920 (N_1920,N_849,N_585);
and U1921 (N_1921,N_421,N_462);
and U1922 (N_1922,N_77,N_923);
nand U1923 (N_1923,N_846,N_8);
nor U1924 (N_1924,N_151,N_72);
nand U1925 (N_1925,N_89,N_557);
nor U1926 (N_1926,N_418,N_468);
nand U1927 (N_1927,N_559,N_983);
and U1928 (N_1928,N_946,N_955);
nor U1929 (N_1929,N_669,N_825);
nand U1930 (N_1930,N_896,N_534);
or U1931 (N_1931,N_423,N_604);
nor U1932 (N_1932,N_319,N_238);
or U1933 (N_1933,N_476,N_33);
and U1934 (N_1934,N_893,N_16);
nor U1935 (N_1935,N_63,N_569);
and U1936 (N_1936,N_72,N_785);
nor U1937 (N_1937,N_713,N_400);
or U1938 (N_1938,N_138,N_912);
and U1939 (N_1939,N_696,N_208);
or U1940 (N_1940,N_945,N_70);
and U1941 (N_1941,N_819,N_649);
and U1942 (N_1942,N_205,N_179);
nor U1943 (N_1943,N_324,N_731);
nor U1944 (N_1944,N_612,N_224);
nor U1945 (N_1945,N_439,N_693);
nand U1946 (N_1946,N_91,N_85);
and U1947 (N_1947,N_899,N_224);
nor U1948 (N_1948,N_272,N_540);
nand U1949 (N_1949,N_4,N_330);
and U1950 (N_1950,N_347,N_81);
and U1951 (N_1951,N_545,N_982);
nand U1952 (N_1952,N_558,N_958);
and U1953 (N_1953,N_671,N_963);
nand U1954 (N_1954,N_758,N_829);
or U1955 (N_1955,N_252,N_315);
nor U1956 (N_1956,N_542,N_560);
or U1957 (N_1957,N_577,N_674);
nand U1958 (N_1958,N_949,N_864);
nand U1959 (N_1959,N_268,N_104);
or U1960 (N_1960,N_897,N_829);
nand U1961 (N_1961,N_518,N_403);
nand U1962 (N_1962,N_787,N_972);
and U1963 (N_1963,N_958,N_330);
or U1964 (N_1964,N_508,N_915);
or U1965 (N_1965,N_339,N_575);
or U1966 (N_1966,N_222,N_599);
nand U1967 (N_1967,N_863,N_792);
and U1968 (N_1968,N_744,N_80);
nor U1969 (N_1969,N_133,N_210);
or U1970 (N_1970,N_827,N_230);
nor U1971 (N_1971,N_113,N_464);
nor U1972 (N_1972,N_375,N_177);
or U1973 (N_1973,N_781,N_215);
nand U1974 (N_1974,N_158,N_591);
and U1975 (N_1975,N_815,N_255);
nand U1976 (N_1976,N_756,N_614);
nor U1977 (N_1977,N_248,N_733);
nand U1978 (N_1978,N_383,N_155);
or U1979 (N_1979,N_874,N_551);
nor U1980 (N_1980,N_27,N_407);
and U1981 (N_1981,N_994,N_695);
nor U1982 (N_1982,N_601,N_869);
nor U1983 (N_1983,N_557,N_46);
nor U1984 (N_1984,N_298,N_376);
or U1985 (N_1985,N_425,N_656);
nand U1986 (N_1986,N_691,N_788);
nor U1987 (N_1987,N_233,N_53);
nor U1988 (N_1988,N_685,N_707);
or U1989 (N_1989,N_172,N_540);
and U1990 (N_1990,N_463,N_993);
nand U1991 (N_1991,N_239,N_312);
and U1992 (N_1992,N_157,N_687);
nand U1993 (N_1993,N_287,N_86);
nand U1994 (N_1994,N_876,N_461);
nand U1995 (N_1995,N_591,N_780);
nor U1996 (N_1996,N_664,N_246);
and U1997 (N_1997,N_739,N_659);
or U1998 (N_1998,N_599,N_345);
nand U1999 (N_1999,N_219,N_136);
nor U2000 (N_2000,N_1423,N_1352);
and U2001 (N_2001,N_1492,N_1845);
nor U2002 (N_2002,N_1049,N_1351);
nor U2003 (N_2003,N_1642,N_1228);
nor U2004 (N_2004,N_1505,N_1982);
nor U2005 (N_2005,N_1878,N_1294);
or U2006 (N_2006,N_1712,N_1614);
or U2007 (N_2007,N_1452,N_1446);
nand U2008 (N_2008,N_1732,N_1208);
and U2009 (N_2009,N_1564,N_1115);
or U2010 (N_2010,N_1218,N_1034);
nor U2011 (N_2011,N_1976,N_1170);
or U2012 (N_2012,N_1815,N_1634);
or U2013 (N_2013,N_1187,N_1731);
nor U2014 (N_2014,N_1859,N_1223);
nand U2015 (N_2015,N_1710,N_1511);
or U2016 (N_2016,N_1690,N_1318);
or U2017 (N_2017,N_1464,N_1136);
nand U2018 (N_2018,N_1965,N_1415);
or U2019 (N_2019,N_1281,N_1526);
nor U2020 (N_2020,N_1935,N_1172);
nand U2021 (N_2021,N_1593,N_1366);
nand U2022 (N_2022,N_1933,N_1521);
nand U2023 (N_2023,N_1917,N_1998);
nor U2024 (N_2024,N_1900,N_1451);
nor U2025 (N_2025,N_1814,N_1461);
and U2026 (N_2026,N_1134,N_1552);
and U2027 (N_2027,N_1072,N_1879);
or U2028 (N_2028,N_1680,N_1264);
nand U2029 (N_2029,N_1481,N_1353);
xor U2030 (N_2030,N_1655,N_1055);
nor U2031 (N_2031,N_1988,N_1392);
nand U2032 (N_2032,N_1382,N_1079);
or U2033 (N_2033,N_1818,N_1581);
or U2034 (N_2034,N_1930,N_1458);
nand U2035 (N_2035,N_1506,N_1188);
or U2036 (N_2036,N_1243,N_1307);
and U2037 (N_2037,N_1373,N_1338);
or U2038 (N_2038,N_1271,N_1117);
nand U2039 (N_2039,N_1705,N_1219);
nor U2040 (N_2040,N_1555,N_1590);
nand U2041 (N_2041,N_1334,N_1694);
nand U2042 (N_2042,N_1844,N_1400);
or U2043 (N_2043,N_1911,N_1221);
nor U2044 (N_2044,N_1798,N_1015);
nor U2045 (N_2045,N_1517,N_1257);
or U2046 (N_2046,N_1148,N_1058);
or U2047 (N_2047,N_1527,N_1867);
or U2048 (N_2048,N_1514,N_1191);
nor U2049 (N_2049,N_1490,N_1019);
and U2050 (N_2050,N_1629,N_1355);
nand U2051 (N_2051,N_1702,N_1887);
nand U2052 (N_2052,N_1226,N_1184);
and U2053 (N_2053,N_1291,N_1484);
nor U2054 (N_2054,N_1945,N_1475);
nand U2055 (N_2055,N_1596,N_1606);
nor U2056 (N_2056,N_1745,N_1245);
nand U2057 (N_2057,N_1923,N_1643);
or U2058 (N_2058,N_1996,N_1320);
and U2059 (N_2059,N_1649,N_1599);
and U2060 (N_2060,N_1685,N_1774);
and U2061 (N_2061,N_1362,N_1340);
and U2062 (N_2062,N_1277,N_1151);
and U2063 (N_2063,N_1078,N_1118);
nor U2064 (N_2064,N_1420,N_1825);
nor U2065 (N_2065,N_1431,N_1207);
nor U2066 (N_2066,N_1014,N_1623);
and U2067 (N_2067,N_1794,N_1173);
nor U2068 (N_2068,N_1106,N_1582);
nand U2069 (N_2069,N_1341,N_1906);
and U2070 (N_2070,N_1254,N_1872);
nand U2071 (N_2071,N_1986,N_1220);
nand U2072 (N_2072,N_1765,N_1388);
or U2073 (N_2073,N_1246,N_1928);
nand U2074 (N_2074,N_1678,N_1699);
or U2075 (N_2075,N_1529,N_1293);
and U2076 (N_2076,N_1166,N_1357);
nor U2077 (N_2077,N_1298,N_1323);
nor U2078 (N_2078,N_1720,N_1455);
nor U2079 (N_2079,N_1259,N_1378);
and U2080 (N_2080,N_1403,N_1483);
or U2081 (N_2081,N_1442,N_1723);
or U2082 (N_2082,N_1761,N_1627);
nand U2083 (N_2083,N_1874,N_1537);
nand U2084 (N_2084,N_1750,N_1894);
or U2085 (N_2085,N_1279,N_1572);
nand U2086 (N_2086,N_1578,N_1372);
or U2087 (N_2087,N_1622,N_1729);
or U2088 (N_2088,N_1896,N_1863);
nand U2089 (N_2089,N_1496,N_1493);
or U2090 (N_2090,N_1085,N_1179);
or U2091 (N_2091,N_1213,N_1076);
and U2092 (N_2092,N_1544,N_1441);
or U2093 (N_2093,N_1823,N_1494);
or U2094 (N_2094,N_1401,N_1788);
and U2095 (N_2095,N_1342,N_1531);
nand U2096 (N_2096,N_1503,N_1875);
and U2097 (N_2097,N_1947,N_1060);
or U2098 (N_2098,N_1802,N_1239);
or U2099 (N_2099,N_1405,N_1737);
or U2100 (N_2100,N_1783,N_1399);
or U2101 (N_2101,N_1045,N_1994);
nand U2102 (N_2102,N_1495,N_1656);
nor U2103 (N_2103,N_1465,N_1944);
or U2104 (N_2104,N_1385,N_1093);
nand U2105 (N_2105,N_1889,N_1381);
and U2106 (N_2106,N_1953,N_1591);
nor U2107 (N_2107,N_1430,N_1197);
or U2108 (N_2108,N_1968,N_1449);
nor U2109 (N_2109,N_1849,N_1282);
and U2110 (N_2110,N_1133,N_1891);
and U2111 (N_2111,N_1065,N_1039);
nor U2112 (N_2112,N_1903,N_1651);
and U2113 (N_2113,N_1384,N_1285);
nand U2114 (N_2114,N_1883,N_1274);
or U2115 (N_2115,N_1630,N_1209);
nand U2116 (N_2116,N_1343,N_1296);
nand U2117 (N_2117,N_1297,N_1668);
or U2118 (N_2118,N_1733,N_1325);
nand U2119 (N_2119,N_1198,N_1672);
or U2120 (N_2120,N_1673,N_1006);
nand U2121 (N_2121,N_1562,N_1989);
or U2122 (N_2122,N_1217,N_1892);
or U2123 (N_2123,N_1743,N_1364);
or U2124 (N_2124,N_1909,N_1127);
or U2125 (N_2125,N_1719,N_1434);
and U2126 (N_2126,N_1509,N_1326);
or U2127 (N_2127,N_1156,N_1069);
or U2128 (N_2128,N_1225,N_1063);
nand U2129 (N_2129,N_1235,N_1158);
nor U2130 (N_2130,N_1612,N_1222);
nor U2131 (N_2131,N_1440,N_1489);
nor U2132 (N_2132,N_1135,N_1196);
nor U2133 (N_2133,N_1589,N_1155);
nand U2134 (N_2134,N_1677,N_1515);
nor U2135 (N_2135,N_1328,N_1402);
nand U2136 (N_2136,N_1113,N_1467);
and U2137 (N_2137,N_1309,N_1661);
and U2138 (N_2138,N_1676,N_1966);
and U2139 (N_2139,N_1682,N_1550);
nor U2140 (N_2140,N_1561,N_1653);
or U2141 (N_2141,N_1703,N_1919);
nor U2142 (N_2142,N_1044,N_1299);
and U2143 (N_2143,N_1398,N_1011);
nand U2144 (N_2144,N_1168,N_1358);
xnor U2145 (N_2145,N_1062,N_1631);
nand U2146 (N_2146,N_1791,N_1250);
nand U2147 (N_2147,N_1252,N_1664);
or U2148 (N_2148,N_1871,N_1958);
nor U2149 (N_2149,N_1500,N_1478);
or U2150 (N_2150,N_1329,N_1738);
or U2151 (N_2151,N_1551,N_1626);
nand U2152 (N_2152,N_1967,N_1726);
or U2153 (N_2153,N_1161,N_1230);
or U2154 (N_2154,N_1588,N_1302);
nor U2155 (N_2155,N_1052,N_1033);
nor U2156 (N_2156,N_1510,N_1881);
and U2157 (N_2157,N_1706,N_1920);
and U2158 (N_2158,N_1885,N_1337);
xor U2159 (N_2159,N_1598,N_1051);
nor U2160 (N_2160,N_1059,N_1010);
nand U2161 (N_2161,N_1283,N_1284);
and U2162 (N_2162,N_1713,N_1053);
nand U2163 (N_2163,N_1573,N_1162);
nand U2164 (N_2164,N_1330,N_1110);
and U2165 (N_2165,N_1108,N_1335);
nand U2166 (N_2166,N_1043,N_1803);
nor U2167 (N_2167,N_1576,N_1542);
or U2168 (N_2168,N_1129,N_1025);
or U2169 (N_2169,N_1018,N_1957);
nand U2170 (N_2170,N_1321,N_1541);
nand U2171 (N_2171,N_1955,N_1021);
nand U2172 (N_2172,N_1865,N_1377);
or U2173 (N_2173,N_1313,N_1905);
or U2174 (N_2174,N_1799,N_1102);
nor U2175 (N_2175,N_1404,N_1003);
and U2176 (N_2176,N_1806,N_1406);
nor U2177 (N_2177,N_1012,N_1114);
nor U2178 (N_2178,N_1205,N_1308);
or U2179 (N_2179,N_1587,N_1212);
and U2180 (N_2180,N_1575,N_1766);
and U2181 (N_2181,N_1997,N_1004);
or U2182 (N_2182,N_1075,N_1331);
nor U2183 (N_2183,N_1781,N_1122);
nor U2184 (N_2184,N_1787,N_1499);
and U2185 (N_2185,N_1615,N_1862);
or U2186 (N_2186,N_1776,N_1696);
and U2187 (N_2187,N_1816,N_1670);
or U2188 (N_2188,N_1763,N_1348);
or U2189 (N_2189,N_1407,N_1746);
and U2190 (N_2190,N_1050,N_1350);
or U2191 (N_2191,N_1248,N_1183);
and U2192 (N_2192,N_1240,N_1416);
xor U2193 (N_2193,N_1425,N_1104);
nand U2194 (N_2194,N_1779,N_1876);
nand U2195 (N_2195,N_1586,N_1831);
nand U2196 (N_2196,N_1539,N_1751);
nand U2197 (N_2197,N_1534,N_1370);
nor U2198 (N_2198,N_1826,N_1999);
or U2199 (N_2199,N_1453,N_1669);
nand U2200 (N_2200,N_1456,N_1922);
nor U2201 (N_2201,N_1202,N_1638);
and U2202 (N_2202,N_1064,N_1304);
nor U2203 (N_2203,N_1652,N_1741);
nor U2204 (N_2204,N_1601,N_1460);
or U2205 (N_2205,N_1141,N_1128);
and U2206 (N_2206,N_1360,N_1717);
nand U2207 (N_2207,N_1164,N_1486);
nor U2208 (N_2208,N_1972,N_1345);
or U2209 (N_2209,N_1707,N_1436);
and U2210 (N_2210,N_1178,N_1035);
nand U2211 (N_2211,N_1667,N_1868);
nor U2212 (N_2212,N_1870,N_1090);
nand U2213 (N_2213,N_1447,N_1557);
nor U2214 (N_2214,N_1523,N_1952);
nor U2215 (N_2215,N_1548,N_1083);
nand U2216 (N_2216,N_1175,N_1288);
or U2217 (N_2217,N_1476,N_1227);
or U2218 (N_2218,N_1782,N_1140);
nand U2219 (N_2219,N_1146,N_1639);
nor U2220 (N_2220,N_1971,N_1290);
nor U2221 (N_2221,N_1547,N_1024);
or U2222 (N_2222,N_1468,N_1154);
and U2223 (N_2223,N_1211,N_1962);
and U2224 (N_2224,N_1784,N_1603);
or U2225 (N_2225,N_1995,N_1632);
nand U2226 (N_2226,N_1808,N_1621);
nor U2227 (N_2227,N_1472,N_1890);
nor U2228 (N_2228,N_1897,N_1993);
or U2229 (N_2229,N_1171,N_1267);
nand U2230 (N_2230,N_1736,N_1800);
nand U2231 (N_2231,N_1327,N_1303);
or U2232 (N_2232,N_1098,N_1913);
or U2233 (N_2233,N_1809,N_1269);
or U2234 (N_2234,N_1822,N_1032);
nor U2235 (N_2235,N_1904,N_1444);
nor U2236 (N_2236,N_1827,N_1138);
nor U2237 (N_2237,N_1375,N_1580);
nor U2238 (N_2238,N_1394,N_1908);
and U2239 (N_2239,N_1801,N_1924);
nor U2240 (N_2240,N_1324,N_1253);
or U2241 (N_2241,N_1540,N_1347);
nor U2242 (N_2242,N_1981,N_1443);
or U2243 (N_2243,N_1695,N_1236);
and U2244 (N_2244,N_1866,N_1426);
and U2245 (N_2245,N_1585,N_1925);
nor U2246 (N_2246,N_1459,N_1419);
xnor U2247 (N_2247,N_1869,N_1648);
nand U2248 (N_2248,N_1145,N_1688);
nand U2249 (N_2249,N_1915,N_1657);
nor U2250 (N_2250,N_1747,N_1956);
nor U2251 (N_2251,N_1853,N_1807);
and U2252 (N_2252,N_1939,N_1543);
nand U2253 (N_2253,N_1824,N_1268);
or U2254 (N_2254,N_1675,N_1697);
and U2255 (N_2255,N_1311,N_1275);
nor U2256 (N_2256,N_1821,N_1099);
and U2257 (N_2257,N_1262,N_1984);
nor U2258 (N_2258,N_1777,N_1389);
and U2259 (N_2259,N_1721,N_1316);
nand U2260 (N_2260,N_1463,N_1975);
and U2261 (N_2261,N_1433,N_1435);
or U2262 (N_2262,N_1497,N_1742);
or U2263 (N_2263,N_1735,N_1068);
nor U2264 (N_2264,N_1684,N_1711);
nor U2265 (N_2265,N_1759,N_1837);
nor U2266 (N_2266,N_1216,N_1709);
nor U2267 (N_2267,N_1658,N_1387);
or U2268 (N_2268,N_1546,N_1429);
or U2269 (N_2269,N_1566,N_1718);
nand U2270 (N_2270,N_1786,N_1414);
and U2271 (N_2271,N_1959,N_1026);
and U2272 (N_2272,N_1992,N_1165);
or U2273 (N_2273,N_1292,N_1031);
nand U2274 (N_2274,N_1336,N_1948);
or U2275 (N_2275,N_1409,N_1553);
and U2276 (N_2276,N_1116,N_1570);
nand U2277 (N_2277,N_1176,N_1983);
and U2278 (N_2278,N_1934,N_1773);
or U2279 (N_2279,N_1858,N_1056);
nand U2280 (N_2280,N_1462,N_1757);
nor U2281 (N_2281,N_1636,N_1625);
nor U2282 (N_2282,N_1095,N_1884);
nor U2283 (N_2283,N_1941,N_1528);
or U2284 (N_2284,N_1261,N_1258);
nand U2285 (N_2285,N_1428,N_1371);
nor U2286 (N_2286,N_1954,N_1314);
nor U2287 (N_2287,N_1635,N_1910);
and U2288 (N_2288,N_1856,N_1009);
or U2289 (N_2289,N_1556,N_1042);
or U2290 (N_2290,N_1150,N_1772);
nor U2291 (N_2291,N_1716,N_1109);
or U2292 (N_2292,N_1610,N_1927);
or U2293 (N_2293,N_1628,N_1980);
or U2294 (N_2294,N_1071,N_1130);
or U2295 (N_2295,N_1232,N_1233);
nand U2296 (N_2296,N_1571,N_1811);
or U2297 (N_2297,N_1424,N_1907);
nand U2298 (N_2298,N_1081,N_1990);
and U2299 (N_2299,N_1931,N_1882);
nor U2300 (N_2300,N_1349,N_1144);
or U2301 (N_2301,N_1077,N_1964);
nor U2302 (N_2302,N_1942,N_1091);
nor U2303 (N_2303,N_1790,N_1020);
or U2304 (N_2304,N_1912,N_1665);
or U2305 (N_2305,N_1023,N_1951);
nor U2306 (N_2306,N_1758,N_1181);
nand U2307 (N_2307,N_1082,N_1466);
xor U2308 (N_2308,N_1088,N_1549);
nand U2309 (N_2309,N_1270,N_1877);
or U2310 (N_2310,N_1074,N_1700);
and U2311 (N_2311,N_1383,N_1969);
nand U2312 (N_2312,N_1192,N_1200);
nand U2313 (N_2313,N_1898,N_1963);
nor U2314 (N_2314,N_1251,N_1847);
nor U2315 (N_2315,N_1393,N_1609);
nor U2316 (N_2316,N_1038,N_1391);
nor U2317 (N_2317,N_1397,N_1177);
and U2318 (N_2318,N_1748,N_1839);
nor U2319 (N_2319,N_1123,N_1624);
nand U2320 (N_2320,N_1125,N_1620);
or U2321 (N_2321,N_1785,N_1448);
nand U2322 (N_2322,N_1535,N_1344);
and U2323 (N_2323,N_1554,N_1132);
and U2324 (N_2324,N_1728,N_1600);
and U2325 (N_2325,N_1810,N_1278);
nand U2326 (N_2326,N_1408,N_1244);
or U2327 (N_2327,N_1829,N_1061);
or U2328 (N_2328,N_1880,N_1473);
and U2329 (N_2329,N_1067,N_1092);
and U2330 (N_2330,N_1438,N_1206);
nor U2331 (N_2331,N_1577,N_1796);
and U2332 (N_2332,N_1027,N_1792);
and U2333 (N_2333,N_1595,N_1902);
nand U2334 (N_2334,N_1835,N_1159);
and U2335 (N_2335,N_1522,N_1979);
and U2336 (N_2336,N_1938,N_1396);
nand U2337 (N_2337,N_1502,N_1525);
nand U2338 (N_2338,N_1961,N_1780);
nand U2339 (N_2339,N_1985,N_1753);
nand U2340 (N_2340,N_1359,N_1273);
nor U2341 (N_2341,N_1618,N_1469);
xor U2342 (N_2342,N_1769,N_1182);
and U2343 (N_2343,N_1255,N_1491);
nor U2344 (N_2344,N_1819,N_1932);
and U2345 (N_2345,N_1617,N_1597);
and U2346 (N_2346,N_1756,N_1704);
and U2347 (N_2347,N_1893,N_1265);
and U2348 (N_2348,N_1001,N_1513);
or U2349 (N_2349,N_1137,N_1368);
or U2350 (N_2350,N_1855,N_1616);
or U2351 (N_2351,N_1080,N_1730);
nor U2352 (N_2352,N_1305,N_1760);
nor U2353 (N_2353,N_1508,N_1000);
nor U2354 (N_2354,N_1701,N_1121);
or U2355 (N_2355,N_1861,N_1752);
or U2356 (N_2356,N_1005,N_1584);
nand U2357 (N_2357,N_1937,N_1689);
nand U2358 (N_2358,N_1926,N_1633);
nand U2359 (N_2359,N_1978,N_1229);
nand U2360 (N_2360,N_1480,N_1663);
and U2361 (N_2361,N_1613,N_1147);
nor U2362 (N_2362,N_1852,N_1410);
and U2363 (N_2363,N_1660,N_1214);
nor U2364 (N_2364,N_1411,N_1256);
and U2365 (N_2365,N_1770,N_1160);
nand U2366 (N_2366,N_1247,N_1828);
and U2367 (N_2367,N_1851,N_1841);
or U2368 (N_2368,N_1797,N_1046);
and U2369 (N_2369,N_1659,N_1193);
nor U2370 (N_2370,N_1640,N_1974);
or U2371 (N_2371,N_1120,N_1153);
nand U2372 (N_2372,N_1725,N_1242);
or U2373 (N_2373,N_1771,N_1683);
or U2374 (N_2374,N_1671,N_1300);
nor U2375 (N_2375,N_1666,N_1376);
nor U2376 (N_2376,N_1107,N_1180);
and U2377 (N_2377,N_1873,N_1813);
nor U2378 (N_2378,N_1524,N_1094);
and U2379 (N_2379,N_1795,N_1749);
nand U2380 (N_2380,N_1286,N_1740);
nor U2381 (N_2381,N_1681,N_1111);
nor U2382 (N_2382,N_1174,N_1762);
and U2383 (N_2383,N_1504,N_1210);
and U2384 (N_2384,N_1946,N_1445);
nor U2385 (N_2385,N_1754,N_1778);
nor U2386 (N_2386,N_1189,N_1950);
nand U2387 (N_2387,N_1361,N_1390);
and U2388 (N_2388,N_1276,N_1037);
and U2389 (N_2389,N_1437,N_1804);
and U2390 (N_2390,N_1013,N_1418);
nor U2391 (N_2391,N_1412,N_1022);
and U2392 (N_2392,N_1838,N_1686);
and U2393 (N_2393,N_1558,N_1310);
nor U2394 (N_2394,N_1190,N_1119);
nand U2395 (N_2395,N_1611,N_1936);
and U2396 (N_2396,N_1734,N_1346);
or U2397 (N_2397,N_1674,N_1516);
nand U2398 (N_2398,N_1637,N_1973);
and U2399 (N_2399,N_1567,N_1650);
nor U2400 (N_2400,N_1482,N_1940);
or U2401 (N_2401,N_1843,N_1693);
nor U2402 (N_2402,N_1101,N_1201);
nor U2403 (N_2403,N_1301,N_1096);
or U2404 (N_2404,N_1708,N_1899);
nand U2405 (N_2405,N_1100,N_1722);
nor U2406 (N_2406,N_1916,N_1149);
nor U2407 (N_2407,N_1619,N_1574);
or U2408 (N_2408,N_1047,N_1157);
nor U2409 (N_2409,N_1563,N_1427);
and U2410 (N_2410,N_1084,N_1518);
or U2411 (N_2411,N_1854,N_1817);
nand U2412 (N_2412,N_1860,N_1319);
and U2413 (N_2413,N_1687,N_1016);
nand U2414 (N_2414,N_1260,N_1501);
nand U2415 (N_2415,N_1048,N_1454);
nor U2416 (N_2416,N_1332,N_1089);
and U2417 (N_2417,N_1289,N_1395);
nand U2418 (N_2418,N_1842,N_1103);
or U2419 (N_2419,N_1367,N_1131);
or U2420 (N_2420,N_1186,N_1943);
nor U2421 (N_2421,N_1356,N_1322);
nor U2422 (N_2422,N_1568,N_1602);
or U2423 (N_2423,N_1379,N_1002);
and U2424 (N_2424,N_1266,N_1241);
nand U2425 (N_2425,N_1036,N_1538);
or U2426 (N_2426,N_1365,N_1203);
and U2427 (N_2427,N_1112,N_1775);
xnor U2428 (N_2428,N_1487,N_1057);
and U2429 (N_2429,N_1886,N_1474);
nor U2430 (N_2430,N_1662,N_1724);
or U2431 (N_2431,N_1848,N_1479);
or U2432 (N_2432,N_1317,N_1374);
nand U2433 (N_2433,N_1421,N_1224);
nor U2434 (N_2434,N_1812,N_1040);
nand U2435 (N_2435,N_1169,N_1691);
or U2436 (N_2436,N_1498,N_1805);
nand U2437 (N_2437,N_1139,N_1583);
nor U2438 (N_2438,N_1914,N_1744);
nor U2439 (N_2439,N_1987,N_1512);
nand U2440 (N_2440,N_1354,N_1369);
or U2441 (N_2441,N_1579,N_1030);
nor U2442 (N_2442,N_1830,N_1439);
nor U2443 (N_2443,N_1097,N_1569);
and U2444 (N_2444,N_1087,N_1692);
nor U2445 (N_2445,N_1789,N_1413);
nand U2446 (N_2446,N_1470,N_1295);
nand U2447 (N_2447,N_1231,N_1864);
or U2448 (N_2448,N_1450,N_1565);
and U2449 (N_2449,N_1644,N_1991);
nand U2450 (N_2450,N_1432,N_1477);
and U2451 (N_2451,N_1646,N_1608);
or U2452 (N_2452,N_1507,N_1530);
nand U2453 (N_2453,N_1124,N_1888);
or U2454 (N_2454,N_1857,N_1280);
and U2455 (N_2455,N_1086,N_1380);
nand U2456 (N_2456,N_1533,N_1306);
nor U2457 (N_2457,N_1645,N_1457);
nor U2458 (N_2458,N_1679,N_1417);
or U2459 (N_2459,N_1312,N_1287);
or U2460 (N_2460,N_1833,N_1272);
or U2461 (N_2461,N_1194,N_1921);
nor U2462 (N_2462,N_1768,N_1007);
or U2463 (N_2463,N_1070,N_1850);
or U2464 (N_2464,N_1654,N_1234);
or U2465 (N_2465,N_1846,N_1840);
or U2466 (N_2466,N_1167,N_1755);
or U2467 (N_2467,N_1594,N_1315);
or U2468 (N_2468,N_1714,N_1066);
nor U2469 (N_2469,N_1532,N_1471);
nand U2470 (N_2470,N_1363,N_1054);
nor U2471 (N_2471,N_1767,N_1105);
or U2472 (N_2472,N_1545,N_1901);
nand U2473 (N_2473,N_1764,N_1185);
nor U2474 (N_2474,N_1918,N_1249);
nand U2475 (N_2475,N_1126,N_1488);
nor U2476 (N_2476,N_1029,N_1715);
and U2477 (N_2477,N_1820,N_1143);
and U2478 (N_2478,N_1836,N_1238);
or U2479 (N_2479,N_1028,N_1607);
and U2480 (N_2480,N_1073,N_1339);
xnor U2481 (N_2481,N_1386,N_1017);
or U2482 (N_2482,N_1152,N_1199);
nand U2483 (N_2483,N_1605,N_1041);
nand U2484 (N_2484,N_1739,N_1204);
and U2485 (N_2485,N_1519,N_1536);
nand U2486 (N_2486,N_1727,N_1834);
nor U2487 (N_2487,N_1520,N_1237);
or U2488 (N_2488,N_1422,N_1604);
or U2489 (N_2489,N_1215,N_1832);
or U2490 (N_2490,N_1698,N_1970);
and U2491 (N_2491,N_1163,N_1641);
nor U2492 (N_2492,N_1977,N_1949);
and U2493 (N_2493,N_1142,N_1195);
nor U2494 (N_2494,N_1960,N_1929);
nor U2495 (N_2495,N_1647,N_1793);
nand U2496 (N_2496,N_1333,N_1559);
nand U2497 (N_2497,N_1263,N_1895);
nand U2498 (N_2498,N_1485,N_1008);
and U2499 (N_2499,N_1560,N_1592);
nand U2500 (N_2500,N_1022,N_1839);
or U2501 (N_2501,N_1050,N_1345);
nor U2502 (N_2502,N_1597,N_1192);
and U2503 (N_2503,N_1862,N_1562);
nor U2504 (N_2504,N_1406,N_1923);
or U2505 (N_2505,N_1776,N_1346);
or U2506 (N_2506,N_1288,N_1164);
nor U2507 (N_2507,N_1330,N_1744);
and U2508 (N_2508,N_1803,N_1162);
nor U2509 (N_2509,N_1876,N_1753);
nand U2510 (N_2510,N_1568,N_1064);
and U2511 (N_2511,N_1452,N_1162);
and U2512 (N_2512,N_1112,N_1083);
or U2513 (N_2513,N_1567,N_1485);
nand U2514 (N_2514,N_1786,N_1640);
nand U2515 (N_2515,N_1497,N_1892);
and U2516 (N_2516,N_1681,N_1083);
nor U2517 (N_2517,N_1357,N_1333);
nand U2518 (N_2518,N_1783,N_1106);
and U2519 (N_2519,N_1376,N_1067);
nand U2520 (N_2520,N_1435,N_1401);
and U2521 (N_2521,N_1129,N_1450);
nor U2522 (N_2522,N_1301,N_1571);
nor U2523 (N_2523,N_1956,N_1323);
nand U2524 (N_2524,N_1757,N_1071);
and U2525 (N_2525,N_1525,N_1506);
nand U2526 (N_2526,N_1397,N_1562);
and U2527 (N_2527,N_1763,N_1946);
and U2528 (N_2528,N_1707,N_1358);
nand U2529 (N_2529,N_1863,N_1043);
or U2530 (N_2530,N_1684,N_1465);
nor U2531 (N_2531,N_1269,N_1368);
nand U2532 (N_2532,N_1794,N_1955);
nand U2533 (N_2533,N_1813,N_1277);
nor U2534 (N_2534,N_1107,N_1578);
nor U2535 (N_2535,N_1469,N_1911);
nor U2536 (N_2536,N_1342,N_1929);
or U2537 (N_2537,N_1280,N_1340);
and U2538 (N_2538,N_1083,N_1317);
nor U2539 (N_2539,N_1725,N_1148);
nor U2540 (N_2540,N_1142,N_1408);
nand U2541 (N_2541,N_1996,N_1939);
or U2542 (N_2542,N_1855,N_1040);
and U2543 (N_2543,N_1145,N_1491);
nand U2544 (N_2544,N_1127,N_1545);
nand U2545 (N_2545,N_1126,N_1400);
nand U2546 (N_2546,N_1086,N_1991);
or U2547 (N_2547,N_1617,N_1871);
and U2548 (N_2548,N_1758,N_1926);
and U2549 (N_2549,N_1300,N_1919);
or U2550 (N_2550,N_1398,N_1512);
nand U2551 (N_2551,N_1401,N_1345);
and U2552 (N_2552,N_1661,N_1486);
nand U2553 (N_2553,N_1236,N_1462);
and U2554 (N_2554,N_1687,N_1142);
nor U2555 (N_2555,N_1015,N_1559);
and U2556 (N_2556,N_1918,N_1819);
or U2557 (N_2557,N_1505,N_1417);
nand U2558 (N_2558,N_1505,N_1211);
nand U2559 (N_2559,N_1924,N_1542);
nand U2560 (N_2560,N_1754,N_1528);
or U2561 (N_2561,N_1112,N_1093);
and U2562 (N_2562,N_1648,N_1285);
or U2563 (N_2563,N_1409,N_1449);
and U2564 (N_2564,N_1967,N_1143);
and U2565 (N_2565,N_1235,N_1377);
or U2566 (N_2566,N_1692,N_1241);
nor U2567 (N_2567,N_1445,N_1484);
and U2568 (N_2568,N_1856,N_1425);
nor U2569 (N_2569,N_1252,N_1256);
and U2570 (N_2570,N_1728,N_1070);
nand U2571 (N_2571,N_1262,N_1554);
and U2572 (N_2572,N_1306,N_1375);
nor U2573 (N_2573,N_1350,N_1850);
or U2574 (N_2574,N_1999,N_1940);
or U2575 (N_2575,N_1979,N_1832);
nand U2576 (N_2576,N_1298,N_1493);
nor U2577 (N_2577,N_1660,N_1542);
nand U2578 (N_2578,N_1924,N_1793);
or U2579 (N_2579,N_1505,N_1142);
nand U2580 (N_2580,N_1836,N_1698);
and U2581 (N_2581,N_1256,N_1317);
or U2582 (N_2582,N_1941,N_1532);
and U2583 (N_2583,N_1994,N_1093);
nand U2584 (N_2584,N_1276,N_1027);
nand U2585 (N_2585,N_1403,N_1040);
nand U2586 (N_2586,N_1665,N_1269);
nor U2587 (N_2587,N_1246,N_1520);
and U2588 (N_2588,N_1204,N_1374);
nor U2589 (N_2589,N_1664,N_1130);
nand U2590 (N_2590,N_1914,N_1971);
nor U2591 (N_2591,N_1151,N_1453);
nor U2592 (N_2592,N_1520,N_1275);
nor U2593 (N_2593,N_1851,N_1296);
nand U2594 (N_2594,N_1189,N_1088);
and U2595 (N_2595,N_1213,N_1440);
nand U2596 (N_2596,N_1902,N_1185);
or U2597 (N_2597,N_1208,N_1914);
and U2598 (N_2598,N_1527,N_1183);
or U2599 (N_2599,N_1718,N_1280);
and U2600 (N_2600,N_1069,N_1608);
nor U2601 (N_2601,N_1386,N_1081);
nand U2602 (N_2602,N_1721,N_1717);
nand U2603 (N_2603,N_1533,N_1443);
nor U2604 (N_2604,N_1091,N_1633);
and U2605 (N_2605,N_1468,N_1220);
nand U2606 (N_2606,N_1510,N_1067);
or U2607 (N_2607,N_1112,N_1222);
and U2608 (N_2608,N_1773,N_1351);
nor U2609 (N_2609,N_1701,N_1838);
nand U2610 (N_2610,N_1864,N_1844);
nand U2611 (N_2611,N_1686,N_1533);
and U2612 (N_2612,N_1352,N_1549);
and U2613 (N_2613,N_1716,N_1709);
nand U2614 (N_2614,N_1522,N_1711);
nand U2615 (N_2615,N_1101,N_1010);
or U2616 (N_2616,N_1863,N_1409);
or U2617 (N_2617,N_1928,N_1373);
nor U2618 (N_2618,N_1680,N_1580);
and U2619 (N_2619,N_1385,N_1118);
and U2620 (N_2620,N_1112,N_1396);
or U2621 (N_2621,N_1901,N_1772);
or U2622 (N_2622,N_1340,N_1847);
or U2623 (N_2623,N_1892,N_1524);
nor U2624 (N_2624,N_1485,N_1021);
nand U2625 (N_2625,N_1694,N_1113);
and U2626 (N_2626,N_1347,N_1131);
xor U2627 (N_2627,N_1739,N_1887);
nor U2628 (N_2628,N_1278,N_1913);
or U2629 (N_2629,N_1062,N_1562);
or U2630 (N_2630,N_1382,N_1790);
nand U2631 (N_2631,N_1949,N_1556);
or U2632 (N_2632,N_1735,N_1521);
nor U2633 (N_2633,N_1652,N_1103);
or U2634 (N_2634,N_1357,N_1779);
nand U2635 (N_2635,N_1674,N_1938);
and U2636 (N_2636,N_1529,N_1458);
or U2637 (N_2637,N_1698,N_1159);
nor U2638 (N_2638,N_1072,N_1748);
and U2639 (N_2639,N_1537,N_1660);
and U2640 (N_2640,N_1092,N_1725);
and U2641 (N_2641,N_1789,N_1866);
nor U2642 (N_2642,N_1794,N_1704);
nand U2643 (N_2643,N_1657,N_1397);
xnor U2644 (N_2644,N_1830,N_1468);
nor U2645 (N_2645,N_1814,N_1846);
nor U2646 (N_2646,N_1969,N_1879);
nand U2647 (N_2647,N_1555,N_1750);
or U2648 (N_2648,N_1423,N_1482);
nand U2649 (N_2649,N_1518,N_1531);
nand U2650 (N_2650,N_1915,N_1447);
nor U2651 (N_2651,N_1551,N_1855);
and U2652 (N_2652,N_1981,N_1404);
nor U2653 (N_2653,N_1432,N_1879);
nand U2654 (N_2654,N_1259,N_1208);
nor U2655 (N_2655,N_1999,N_1781);
nor U2656 (N_2656,N_1376,N_1740);
nor U2657 (N_2657,N_1581,N_1844);
and U2658 (N_2658,N_1213,N_1650);
nor U2659 (N_2659,N_1485,N_1701);
and U2660 (N_2660,N_1692,N_1473);
nand U2661 (N_2661,N_1633,N_1884);
nor U2662 (N_2662,N_1623,N_1757);
or U2663 (N_2663,N_1992,N_1186);
and U2664 (N_2664,N_1065,N_1868);
and U2665 (N_2665,N_1366,N_1904);
or U2666 (N_2666,N_1165,N_1473);
or U2667 (N_2667,N_1590,N_1988);
and U2668 (N_2668,N_1489,N_1799);
and U2669 (N_2669,N_1123,N_1856);
nor U2670 (N_2670,N_1346,N_1798);
nand U2671 (N_2671,N_1147,N_1447);
nor U2672 (N_2672,N_1393,N_1051);
nand U2673 (N_2673,N_1101,N_1912);
or U2674 (N_2674,N_1510,N_1352);
or U2675 (N_2675,N_1461,N_1279);
or U2676 (N_2676,N_1508,N_1798);
nand U2677 (N_2677,N_1237,N_1191);
or U2678 (N_2678,N_1837,N_1473);
nor U2679 (N_2679,N_1270,N_1554);
nand U2680 (N_2680,N_1349,N_1661);
and U2681 (N_2681,N_1519,N_1465);
nand U2682 (N_2682,N_1704,N_1397);
xnor U2683 (N_2683,N_1838,N_1019);
nor U2684 (N_2684,N_1596,N_1578);
nor U2685 (N_2685,N_1937,N_1432);
nand U2686 (N_2686,N_1881,N_1614);
nand U2687 (N_2687,N_1223,N_1812);
and U2688 (N_2688,N_1520,N_1736);
nand U2689 (N_2689,N_1259,N_1083);
nor U2690 (N_2690,N_1327,N_1204);
nor U2691 (N_2691,N_1183,N_1976);
nor U2692 (N_2692,N_1617,N_1527);
nor U2693 (N_2693,N_1012,N_1924);
nand U2694 (N_2694,N_1994,N_1429);
nand U2695 (N_2695,N_1601,N_1335);
nor U2696 (N_2696,N_1928,N_1285);
nor U2697 (N_2697,N_1710,N_1276);
nand U2698 (N_2698,N_1860,N_1664);
or U2699 (N_2699,N_1977,N_1015);
and U2700 (N_2700,N_1102,N_1873);
nand U2701 (N_2701,N_1744,N_1794);
and U2702 (N_2702,N_1561,N_1526);
or U2703 (N_2703,N_1474,N_1173);
and U2704 (N_2704,N_1570,N_1131);
nor U2705 (N_2705,N_1769,N_1174);
or U2706 (N_2706,N_1520,N_1352);
nor U2707 (N_2707,N_1602,N_1671);
and U2708 (N_2708,N_1966,N_1036);
or U2709 (N_2709,N_1488,N_1197);
and U2710 (N_2710,N_1393,N_1139);
nand U2711 (N_2711,N_1978,N_1311);
xnor U2712 (N_2712,N_1903,N_1565);
or U2713 (N_2713,N_1408,N_1612);
nor U2714 (N_2714,N_1299,N_1250);
nand U2715 (N_2715,N_1126,N_1523);
and U2716 (N_2716,N_1163,N_1546);
and U2717 (N_2717,N_1865,N_1512);
nor U2718 (N_2718,N_1697,N_1696);
or U2719 (N_2719,N_1931,N_1623);
nor U2720 (N_2720,N_1917,N_1744);
nor U2721 (N_2721,N_1842,N_1649);
nand U2722 (N_2722,N_1799,N_1344);
nor U2723 (N_2723,N_1918,N_1824);
nand U2724 (N_2724,N_1239,N_1220);
nor U2725 (N_2725,N_1301,N_1575);
nor U2726 (N_2726,N_1348,N_1791);
nor U2727 (N_2727,N_1367,N_1243);
nand U2728 (N_2728,N_1530,N_1551);
and U2729 (N_2729,N_1143,N_1132);
or U2730 (N_2730,N_1257,N_1991);
nand U2731 (N_2731,N_1788,N_1074);
or U2732 (N_2732,N_1386,N_1334);
or U2733 (N_2733,N_1494,N_1236);
or U2734 (N_2734,N_1507,N_1451);
nor U2735 (N_2735,N_1812,N_1620);
nand U2736 (N_2736,N_1916,N_1077);
or U2737 (N_2737,N_1291,N_1855);
or U2738 (N_2738,N_1503,N_1022);
nor U2739 (N_2739,N_1006,N_1437);
nand U2740 (N_2740,N_1771,N_1794);
or U2741 (N_2741,N_1754,N_1453);
nor U2742 (N_2742,N_1014,N_1337);
and U2743 (N_2743,N_1597,N_1705);
or U2744 (N_2744,N_1667,N_1914);
nor U2745 (N_2745,N_1357,N_1729);
or U2746 (N_2746,N_1461,N_1354);
or U2747 (N_2747,N_1694,N_1124);
nand U2748 (N_2748,N_1783,N_1057);
nand U2749 (N_2749,N_1848,N_1602);
nor U2750 (N_2750,N_1627,N_1378);
or U2751 (N_2751,N_1824,N_1804);
nand U2752 (N_2752,N_1464,N_1585);
or U2753 (N_2753,N_1104,N_1035);
nand U2754 (N_2754,N_1198,N_1618);
nor U2755 (N_2755,N_1802,N_1417);
nand U2756 (N_2756,N_1366,N_1604);
or U2757 (N_2757,N_1556,N_1517);
nor U2758 (N_2758,N_1849,N_1090);
or U2759 (N_2759,N_1816,N_1548);
nand U2760 (N_2760,N_1693,N_1642);
and U2761 (N_2761,N_1666,N_1916);
nor U2762 (N_2762,N_1492,N_1797);
or U2763 (N_2763,N_1336,N_1080);
or U2764 (N_2764,N_1194,N_1097);
or U2765 (N_2765,N_1075,N_1185);
nand U2766 (N_2766,N_1339,N_1950);
nand U2767 (N_2767,N_1893,N_1326);
nand U2768 (N_2768,N_1165,N_1505);
or U2769 (N_2769,N_1382,N_1750);
and U2770 (N_2770,N_1261,N_1028);
and U2771 (N_2771,N_1456,N_1144);
or U2772 (N_2772,N_1579,N_1524);
and U2773 (N_2773,N_1972,N_1512);
nor U2774 (N_2774,N_1478,N_1687);
nor U2775 (N_2775,N_1276,N_1589);
nor U2776 (N_2776,N_1009,N_1094);
and U2777 (N_2777,N_1967,N_1266);
and U2778 (N_2778,N_1702,N_1655);
xnor U2779 (N_2779,N_1358,N_1766);
nor U2780 (N_2780,N_1546,N_1663);
nand U2781 (N_2781,N_1001,N_1090);
nor U2782 (N_2782,N_1397,N_1822);
or U2783 (N_2783,N_1138,N_1483);
nand U2784 (N_2784,N_1972,N_1416);
and U2785 (N_2785,N_1786,N_1829);
or U2786 (N_2786,N_1446,N_1192);
nor U2787 (N_2787,N_1292,N_1016);
or U2788 (N_2788,N_1701,N_1718);
xnor U2789 (N_2789,N_1140,N_1199);
or U2790 (N_2790,N_1924,N_1435);
nand U2791 (N_2791,N_1031,N_1267);
or U2792 (N_2792,N_1336,N_1160);
nor U2793 (N_2793,N_1711,N_1311);
or U2794 (N_2794,N_1386,N_1453);
nor U2795 (N_2795,N_1070,N_1101);
or U2796 (N_2796,N_1825,N_1697);
nand U2797 (N_2797,N_1890,N_1384);
and U2798 (N_2798,N_1307,N_1213);
or U2799 (N_2799,N_1176,N_1079);
nand U2800 (N_2800,N_1667,N_1948);
nand U2801 (N_2801,N_1674,N_1646);
or U2802 (N_2802,N_1104,N_1389);
nor U2803 (N_2803,N_1332,N_1095);
and U2804 (N_2804,N_1883,N_1536);
nand U2805 (N_2805,N_1819,N_1688);
and U2806 (N_2806,N_1574,N_1448);
or U2807 (N_2807,N_1257,N_1030);
nor U2808 (N_2808,N_1725,N_1274);
nor U2809 (N_2809,N_1053,N_1033);
or U2810 (N_2810,N_1619,N_1851);
nor U2811 (N_2811,N_1000,N_1340);
and U2812 (N_2812,N_1416,N_1180);
or U2813 (N_2813,N_1826,N_1371);
nand U2814 (N_2814,N_1359,N_1768);
nand U2815 (N_2815,N_1313,N_1785);
xnor U2816 (N_2816,N_1264,N_1785);
and U2817 (N_2817,N_1487,N_1370);
and U2818 (N_2818,N_1782,N_1578);
nor U2819 (N_2819,N_1057,N_1551);
or U2820 (N_2820,N_1109,N_1959);
nand U2821 (N_2821,N_1500,N_1562);
or U2822 (N_2822,N_1673,N_1257);
nand U2823 (N_2823,N_1984,N_1571);
or U2824 (N_2824,N_1314,N_1948);
and U2825 (N_2825,N_1036,N_1756);
nand U2826 (N_2826,N_1806,N_1681);
nand U2827 (N_2827,N_1827,N_1193);
nand U2828 (N_2828,N_1474,N_1083);
or U2829 (N_2829,N_1855,N_1809);
nor U2830 (N_2830,N_1677,N_1348);
nor U2831 (N_2831,N_1259,N_1196);
or U2832 (N_2832,N_1318,N_1662);
or U2833 (N_2833,N_1839,N_1169);
nand U2834 (N_2834,N_1296,N_1853);
or U2835 (N_2835,N_1425,N_1044);
and U2836 (N_2836,N_1032,N_1721);
and U2837 (N_2837,N_1474,N_1839);
nand U2838 (N_2838,N_1029,N_1221);
and U2839 (N_2839,N_1258,N_1454);
and U2840 (N_2840,N_1562,N_1502);
nand U2841 (N_2841,N_1850,N_1290);
or U2842 (N_2842,N_1580,N_1007);
nor U2843 (N_2843,N_1996,N_1591);
or U2844 (N_2844,N_1962,N_1733);
nor U2845 (N_2845,N_1646,N_1861);
and U2846 (N_2846,N_1655,N_1923);
nor U2847 (N_2847,N_1643,N_1488);
nor U2848 (N_2848,N_1706,N_1803);
or U2849 (N_2849,N_1429,N_1455);
nor U2850 (N_2850,N_1699,N_1231);
or U2851 (N_2851,N_1545,N_1646);
and U2852 (N_2852,N_1160,N_1066);
nor U2853 (N_2853,N_1380,N_1958);
or U2854 (N_2854,N_1309,N_1405);
nand U2855 (N_2855,N_1132,N_1967);
or U2856 (N_2856,N_1989,N_1736);
and U2857 (N_2857,N_1468,N_1224);
nor U2858 (N_2858,N_1962,N_1664);
nor U2859 (N_2859,N_1764,N_1441);
nor U2860 (N_2860,N_1735,N_1963);
or U2861 (N_2861,N_1591,N_1659);
or U2862 (N_2862,N_1235,N_1248);
nor U2863 (N_2863,N_1529,N_1250);
nor U2864 (N_2864,N_1448,N_1294);
and U2865 (N_2865,N_1653,N_1613);
or U2866 (N_2866,N_1534,N_1884);
nand U2867 (N_2867,N_1015,N_1589);
nor U2868 (N_2868,N_1715,N_1406);
nand U2869 (N_2869,N_1779,N_1984);
and U2870 (N_2870,N_1391,N_1049);
and U2871 (N_2871,N_1690,N_1459);
nor U2872 (N_2872,N_1941,N_1188);
and U2873 (N_2873,N_1943,N_1231);
nor U2874 (N_2874,N_1410,N_1245);
and U2875 (N_2875,N_1138,N_1587);
nand U2876 (N_2876,N_1532,N_1889);
nand U2877 (N_2877,N_1150,N_1928);
nand U2878 (N_2878,N_1551,N_1093);
and U2879 (N_2879,N_1044,N_1469);
nand U2880 (N_2880,N_1953,N_1595);
nand U2881 (N_2881,N_1272,N_1484);
nand U2882 (N_2882,N_1635,N_1658);
nor U2883 (N_2883,N_1658,N_1875);
nand U2884 (N_2884,N_1670,N_1168);
or U2885 (N_2885,N_1048,N_1728);
nor U2886 (N_2886,N_1269,N_1301);
or U2887 (N_2887,N_1101,N_1877);
nor U2888 (N_2888,N_1389,N_1854);
nand U2889 (N_2889,N_1378,N_1974);
and U2890 (N_2890,N_1695,N_1830);
or U2891 (N_2891,N_1869,N_1504);
nor U2892 (N_2892,N_1341,N_1137);
nand U2893 (N_2893,N_1239,N_1275);
and U2894 (N_2894,N_1962,N_1436);
and U2895 (N_2895,N_1241,N_1606);
nor U2896 (N_2896,N_1241,N_1059);
nand U2897 (N_2897,N_1305,N_1518);
nor U2898 (N_2898,N_1759,N_1086);
or U2899 (N_2899,N_1589,N_1673);
and U2900 (N_2900,N_1882,N_1117);
or U2901 (N_2901,N_1439,N_1772);
and U2902 (N_2902,N_1465,N_1296);
and U2903 (N_2903,N_1200,N_1111);
nor U2904 (N_2904,N_1314,N_1928);
or U2905 (N_2905,N_1138,N_1791);
and U2906 (N_2906,N_1624,N_1956);
or U2907 (N_2907,N_1919,N_1489);
and U2908 (N_2908,N_1238,N_1582);
and U2909 (N_2909,N_1033,N_1073);
nor U2910 (N_2910,N_1860,N_1326);
and U2911 (N_2911,N_1109,N_1487);
and U2912 (N_2912,N_1603,N_1417);
nand U2913 (N_2913,N_1559,N_1997);
nand U2914 (N_2914,N_1866,N_1980);
nor U2915 (N_2915,N_1685,N_1854);
nor U2916 (N_2916,N_1391,N_1576);
nor U2917 (N_2917,N_1487,N_1298);
or U2918 (N_2918,N_1324,N_1790);
nor U2919 (N_2919,N_1299,N_1125);
and U2920 (N_2920,N_1883,N_1050);
nand U2921 (N_2921,N_1817,N_1408);
nor U2922 (N_2922,N_1031,N_1627);
nand U2923 (N_2923,N_1964,N_1628);
nor U2924 (N_2924,N_1936,N_1149);
or U2925 (N_2925,N_1233,N_1825);
and U2926 (N_2926,N_1686,N_1163);
and U2927 (N_2927,N_1848,N_1018);
and U2928 (N_2928,N_1446,N_1683);
nor U2929 (N_2929,N_1390,N_1978);
nand U2930 (N_2930,N_1466,N_1597);
and U2931 (N_2931,N_1399,N_1627);
nand U2932 (N_2932,N_1186,N_1422);
and U2933 (N_2933,N_1226,N_1803);
nand U2934 (N_2934,N_1831,N_1920);
nand U2935 (N_2935,N_1612,N_1197);
or U2936 (N_2936,N_1843,N_1951);
nor U2937 (N_2937,N_1561,N_1578);
and U2938 (N_2938,N_1016,N_1559);
nand U2939 (N_2939,N_1365,N_1731);
nand U2940 (N_2940,N_1721,N_1532);
nand U2941 (N_2941,N_1393,N_1983);
and U2942 (N_2942,N_1600,N_1026);
nor U2943 (N_2943,N_1542,N_1930);
nand U2944 (N_2944,N_1953,N_1320);
or U2945 (N_2945,N_1079,N_1925);
or U2946 (N_2946,N_1031,N_1207);
xnor U2947 (N_2947,N_1779,N_1995);
and U2948 (N_2948,N_1841,N_1269);
nand U2949 (N_2949,N_1993,N_1739);
nand U2950 (N_2950,N_1501,N_1644);
nand U2951 (N_2951,N_1713,N_1195);
and U2952 (N_2952,N_1971,N_1664);
and U2953 (N_2953,N_1792,N_1746);
nor U2954 (N_2954,N_1027,N_1459);
and U2955 (N_2955,N_1944,N_1222);
or U2956 (N_2956,N_1468,N_1299);
nor U2957 (N_2957,N_1504,N_1222);
or U2958 (N_2958,N_1455,N_1270);
nor U2959 (N_2959,N_1617,N_1296);
xor U2960 (N_2960,N_1815,N_1319);
or U2961 (N_2961,N_1697,N_1054);
or U2962 (N_2962,N_1158,N_1816);
nand U2963 (N_2963,N_1323,N_1207);
nor U2964 (N_2964,N_1842,N_1014);
or U2965 (N_2965,N_1532,N_1896);
nor U2966 (N_2966,N_1800,N_1599);
nor U2967 (N_2967,N_1015,N_1419);
or U2968 (N_2968,N_1788,N_1147);
or U2969 (N_2969,N_1854,N_1544);
nor U2970 (N_2970,N_1567,N_1837);
nor U2971 (N_2971,N_1377,N_1312);
nand U2972 (N_2972,N_1122,N_1254);
nor U2973 (N_2973,N_1780,N_1986);
or U2974 (N_2974,N_1631,N_1567);
nor U2975 (N_2975,N_1871,N_1264);
or U2976 (N_2976,N_1517,N_1330);
or U2977 (N_2977,N_1561,N_1060);
nand U2978 (N_2978,N_1273,N_1662);
nor U2979 (N_2979,N_1625,N_1620);
nor U2980 (N_2980,N_1892,N_1586);
nor U2981 (N_2981,N_1813,N_1332);
nand U2982 (N_2982,N_1616,N_1275);
nand U2983 (N_2983,N_1978,N_1994);
nor U2984 (N_2984,N_1322,N_1534);
nand U2985 (N_2985,N_1864,N_1621);
and U2986 (N_2986,N_1023,N_1113);
and U2987 (N_2987,N_1208,N_1085);
or U2988 (N_2988,N_1631,N_1655);
nor U2989 (N_2989,N_1481,N_1327);
nor U2990 (N_2990,N_1106,N_1733);
xnor U2991 (N_2991,N_1995,N_1754);
nor U2992 (N_2992,N_1902,N_1050);
and U2993 (N_2993,N_1035,N_1352);
nand U2994 (N_2994,N_1805,N_1317);
and U2995 (N_2995,N_1734,N_1076);
nand U2996 (N_2996,N_1707,N_1869);
nor U2997 (N_2997,N_1116,N_1309);
nor U2998 (N_2998,N_1810,N_1410);
and U2999 (N_2999,N_1236,N_1332);
or UO_0 (O_0,N_2973,N_2551);
nor UO_1 (O_1,N_2979,N_2055);
or UO_2 (O_2,N_2186,N_2522);
nor UO_3 (O_3,N_2119,N_2337);
nor UO_4 (O_4,N_2845,N_2559);
and UO_5 (O_5,N_2224,N_2994);
nand UO_6 (O_6,N_2884,N_2724);
or UO_7 (O_7,N_2447,N_2129);
and UO_8 (O_8,N_2537,N_2817);
and UO_9 (O_9,N_2378,N_2099);
or UO_10 (O_10,N_2439,N_2614);
and UO_11 (O_11,N_2036,N_2197);
or UO_12 (O_12,N_2980,N_2310);
nor UO_13 (O_13,N_2628,N_2667);
and UO_14 (O_14,N_2966,N_2627);
nand UO_15 (O_15,N_2750,N_2606);
nor UO_16 (O_16,N_2235,N_2113);
nor UO_17 (O_17,N_2526,N_2839);
nand UO_18 (O_18,N_2192,N_2883);
nand UO_19 (O_19,N_2577,N_2516);
and UO_20 (O_20,N_2803,N_2266);
and UO_21 (O_21,N_2459,N_2728);
or UO_22 (O_22,N_2366,N_2858);
nor UO_23 (O_23,N_2581,N_2991);
nor UO_24 (O_24,N_2521,N_2073);
or UO_25 (O_25,N_2900,N_2430);
or UO_26 (O_26,N_2511,N_2069);
nand UO_27 (O_27,N_2390,N_2513);
or UO_28 (O_28,N_2475,N_2125);
and UO_29 (O_29,N_2638,N_2322);
and UO_30 (O_30,N_2666,N_2919);
and UO_31 (O_31,N_2643,N_2820);
and UO_32 (O_32,N_2250,N_2589);
xor UO_33 (O_33,N_2792,N_2246);
and UO_34 (O_34,N_2663,N_2751);
and UO_35 (O_35,N_2063,N_2877);
nand UO_36 (O_36,N_2384,N_2339);
nor UO_37 (O_37,N_2917,N_2335);
nor UO_38 (O_38,N_2651,N_2889);
nor UO_39 (O_39,N_2995,N_2670);
and UO_40 (O_40,N_2906,N_2925);
or UO_41 (O_41,N_2901,N_2733);
nand UO_42 (O_42,N_2449,N_2386);
nand UO_43 (O_43,N_2992,N_2054);
and UO_44 (O_44,N_2957,N_2920);
nor UO_45 (O_45,N_2227,N_2950);
nand UO_46 (O_46,N_2615,N_2454);
nor UO_47 (O_47,N_2444,N_2634);
xor UO_48 (O_48,N_2196,N_2239);
or UO_49 (O_49,N_2737,N_2682);
nand UO_50 (O_50,N_2230,N_2466);
or UO_51 (O_51,N_2500,N_2278);
or UO_52 (O_52,N_2044,N_2598);
or UO_53 (O_53,N_2825,N_2968);
and UO_54 (O_54,N_2094,N_2494);
xnor UO_55 (O_55,N_2816,N_2982);
nand UO_56 (O_56,N_2493,N_2954);
and UO_57 (O_57,N_2188,N_2398);
or UO_58 (O_58,N_2918,N_2945);
nor UO_59 (O_59,N_2048,N_2546);
nor UO_60 (O_60,N_2659,N_2706);
and UO_61 (O_61,N_2154,N_2913);
nand UO_62 (O_62,N_2496,N_2397);
or UO_63 (O_63,N_2604,N_2958);
and UO_64 (O_64,N_2132,N_2762);
nor UO_65 (O_65,N_2348,N_2178);
and UO_66 (O_66,N_2201,N_2100);
or UO_67 (O_67,N_2428,N_2865);
nand UO_68 (O_68,N_2130,N_2867);
nand UO_69 (O_69,N_2051,N_2785);
nand UO_70 (O_70,N_2976,N_2861);
or UO_71 (O_71,N_2350,N_2507);
nand UO_72 (O_72,N_2886,N_2258);
xnor UO_73 (O_73,N_2139,N_2106);
nand UO_74 (O_74,N_2838,N_2163);
or UO_75 (O_75,N_2830,N_2394);
or UO_76 (O_76,N_2609,N_2962);
nand UO_77 (O_77,N_2249,N_2332);
nand UO_78 (O_78,N_2757,N_2294);
nand UO_79 (O_79,N_2039,N_2133);
nor UO_80 (O_80,N_2399,N_2436);
or UO_81 (O_81,N_2840,N_2243);
and UO_82 (O_82,N_2946,N_2902);
nor UO_83 (O_83,N_2434,N_2960);
or UO_84 (O_84,N_2531,N_2121);
nor UO_85 (O_85,N_2833,N_2812);
nor UO_86 (O_86,N_2343,N_2126);
and UO_87 (O_87,N_2928,N_2159);
and UO_88 (O_88,N_2116,N_2584);
nand UO_89 (O_89,N_2257,N_2261);
nand UO_90 (O_90,N_2695,N_2574);
or UO_91 (O_91,N_2168,N_2406);
nand UO_92 (O_92,N_2232,N_2713);
nand UO_93 (O_93,N_2468,N_2026);
nor UO_94 (O_94,N_2557,N_2289);
or UO_95 (O_95,N_2520,N_2563);
nand UO_96 (O_96,N_2686,N_2034);
nand UO_97 (O_97,N_2956,N_2318);
or UO_98 (O_98,N_2678,N_2264);
nand UO_99 (O_99,N_2208,N_2417);
or UO_100 (O_100,N_2970,N_2023);
or UO_101 (O_101,N_2710,N_2352);
and UO_102 (O_102,N_2986,N_2095);
nor UO_103 (O_103,N_2087,N_2143);
nand UO_104 (O_104,N_2267,N_2396);
nand UO_105 (O_105,N_2233,N_2420);
nor UO_106 (O_106,N_2619,N_2376);
or UO_107 (O_107,N_2975,N_2618);
nand UO_108 (O_108,N_2527,N_2329);
and UO_109 (O_109,N_2714,N_2076);
or UO_110 (O_110,N_2977,N_2429);
and UO_111 (O_111,N_2798,N_2541);
nand UO_112 (O_112,N_2056,N_2736);
or UO_113 (O_113,N_2117,N_2198);
or UO_114 (O_114,N_2422,N_2897);
nor UO_115 (O_115,N_2864,N_2084);
and UO_116 (O_116,N_2298,N_2972);
and UO_117 (O_117,N_2274,N_2821);
nor UO_118 (O_118,N_2644,N_2810);
nand UO_119 (O_119,N_2277,N_2756);
nand UO_120 (O_120,N_2579,N_2814);
nand UO_121 (O_121,N_2423,N_2880);
and UO_122 (O_122,N_2346,N_2759);
or UO_123 (O_123,N_2115,N_2665);
nand UO_124 (O_124,N_2215,N_2342);
or UO_125 (O_125,N_2488,N_2053);
or UO_126 (O_126,N_2770,N_2797);
nor UO_127 (O_127,N_2984,N_2829);
and UO_128 (O_128,N_2760,N_2842);
nand UO_129 (O_129,N_2734,N_2544);
nor UO_130 (O_130,N_2316,N_2543);
or UO_131 (O_131,N_2911,N_2029);
xnor UO_132 (O_132,N_2899,N_2908);
and UO_133 (O_133,N_2382,N_2501);
nand UO_134 (O_134,N_2974,N_2664);
or UO_135 (O_135,N_2158,N_2641);
nand UO_136 (O_136,N_2532,N_2947);
nor UO_137 (O_137,N_2085,N_2014);
nor UO_138 (O_138,N_2887,N_2823);
or UO_139 (O_139,N_2360,N_2138);
or UO_140 (O_140,N_2012,N_2195);
or UO_141 (O_141,N_2929,N_2391);
or UO_142 (O_142,N_2308,N_2187);
nor UO_143 (O_143,N_2744,N_2875);
xor UO_144 (O_144,N_2131,N_2747);
or UO_145 (O_145,N_2145,N_2834);
or UO_146 (O_146,N_2401,N_2687);
and UO_147 (O_147,N_2170,N_2061);
and UO_148 (O_148,N_2652,N_2755);
nor UO_149 (O_149,N_2912,N_2472);
nor UO_150 (O_150,N_2617,N_2538);
or UO_151 (O_151,N_2699,N_2548);
nand UO_152 (O_152,N_2907,N_2469);
or UO_153 (O_153,N_2487,N_2066);
and UO_154 (O_154,N_2683,N_2005);
nand UO_155 (O_155,N_2328,N_2895);
and UO_156 (O_156,N_2281,N_2037);
or UO_157 (O_157,N_2242,N_2400);
or UO_158 (O_158,N_2273,N_2748);
and UO_159 (O_159,N_2176,N_2743);
nor UO_160 (O_160,N_2746,N_2182);
and UO_161 (O_161,N_2591,N_2971);
and UO_162 (O_162,N_2903,N_2432);
nor UO_163 (O_163,N_2062,N_2509);
or UO_164 (O_164,N_2698,N_2771);
and UO_165 (O_165,N_2361,N_2740);
or UO_166 (O_166,N_2510,N_2435);
or UO_167 (O_167,N_2585,N_2828);
nor UO_168 (O_168,N_2824,N_2616);
and UO_169 (O_169,N_2523,N_2795);
and UO_170 (O_170,N_2373,N_2418);
nor UO_171 (O_171,N_2455,N_2768);
nor UO_172 (O_172,N_2127,N_2403);
or UO_173 (O_173,N_2047,N_2380);
nand UO_174 (O_174,N_2200,N_2720);
or UO_175 (O_175,N_2210,N_2011);
nand UO_176 (O_176,N_2742,N_2203);
nand UO_177 (O_177,N_2671,N_2764);
nor UO_178 (O_178,N_2093,N_2700);
or UO_179 (O_179,N_2878,N_2265);
or UO_180 (O_180,N_2137,N_2850);
or UO_181 (O_181,N_2778,N_2632);
nor UO_182 (O_182,N_2111,N_2114);
and UO_183 (O_183,N_2443,N_2058);
or UO_184 (O_184,N_2575,N_2655);
nor UO_185 (O_185,N_2333,N_2477);
nor UO_186 (O_186,N_2004,N_2456);
and UO_187 (O_187,N_2486,N_2936);
and UO_188 (O_188,N_2882,N_2802);
and UO_189 (O_189,N_2885,N_2402);
or UO_190 (O_190,N_2164,N_2871);
nand UO_191 (O_191,N_2212,N_2582);
xnor UO_192 (O_192,N_2059,N_2288);
nor UO_193 (O_193,N_2465,N_2952);
and UO_194 (O_194,N_2891,N_2324);
and UO_195 (O_195,N_2354,N_2515);
nand UO_196 (O_196,N_2108,N_2939);
or UO_197 (O_197,N_2202,N_2847);
and UO_198 (O_198,N_2152,N_2731);
nor UO_199 (O_199,N_2379,N_2518);
nor UO_200 (O_200,N_2677,N_2122);
or UO_201 (O_201,N_2271,N_2790);
or UO_202 (O_202,N_2782,N_2573);
and UO_203 (O_203,N_2506,N_2171);
nand UO_204 (O_204,N_2844,N_2621);
nor UO_205 (O_205,N_2799,N_2259);
nor UO_206 (O_206,N_2754,N_2718);
or UO_207 (O_207,N_2978,N_2341);
or UO_208 (O_208,N_2779,N_2240);
nand UO_209 (O_209,N_2625,N_2161);
and UO_210 (O_210,N_2852,N_2786);
nand UO_211 (O_211,N_2863,N_2870);
and UO_212 (O_212,N_2179,N_2567);
xnor UO_213 (O_213,N_2022,N_2213);
and UO_214 (O_214,N_2359,N_2112);
nand UO_215 (O_215,N_2514,N_2089);
or UO_216 (O_216,N_2784,N_2098);
nor UO_217 (O_217,N_2789,N_2002);
nand UO_218 (O_218,N_2639,N_2835);
nand UO_219 (O_219,N_2237,N_2461);
or UO_220 (O_220,N_2565,N_2040);
or UO_221 (O_221,N_2254,N_2626);
and UO_222 (O_222,N_2385,N_2943);
or UO_223 (O_223,N_2030,N_2388);
and UO_224 (O_224,N_2876,N_2533);
and UO_225 (O_225,N_2613,N_2938);
nand UO_226 (O_226,N_2220,N_2990);
and UO_227 (O_227,N_2438,N_2482);
nor UO_228 (O_228,N_2872,N_2955);
or UO_229 (O_229,N_2107,N_2204);
and UO_230 (O_230,N_2392,N_2846);
nor UO_231 (O_231,N_2566,N_2175);
or UO_232 (O_232,N_2932,N_2856);
nor UO_233 (O_233,N_2433,N_2826);
xnor UO_234 (O_234,N_2118,N_2097);
nand UO_235 (O_235,N_2753,N_2162);
nand UO_236 (O_236,N_2253,N_2424);
or UO_237 (O_237,N_2989,N_2451);
or UO_238 (O_238,N_2590,N_2964);
or UO_239 (O_239,N_2719,N_2092);
nor UO_240 (O_240,N_2935,N_2916);
or UO_241 (O_241,N_2603,N_2177);
or UO_242 (O_242,N_2416,N_2642);
nand UO_243 (O_243,N_2849,N_2827);
nand UO_244 (O_244,N_2745,N_2715);
and UO_245 (O_245,N_2185,N_2763);
nand UO_246 (O_246,N_2739,N_2460);
nor UO_247 (O_247,N_2286,N_2374);
nand UO_248 (O_248,N_2421,N_2167);
nor UO_249 (O_249,N_2293,N_2951);
or UO_250 (O_250,N_2325,N_2000);
and UO_251 (O_251,N_2189,N_2819);
nand UO_252 (O_252,N_2934,N_2007);
nor UO_253 (O_253,N_2726,N_2776);
and UO_254 (O_254,N_2909,N_2791);
or UO_255 (O_255,N_2080,N_2668);
nand UO_256 (O_256,N_2704,N_2631);
nand UO_257 (O_257,N_2165,N_2749);
or UO_258 (O_258,N_2353,N_2788);
or UO_259 (O_259,N_2305,N_2869);
and UO_260 (O_260,N_2067,N_2234);
nand UO_261 (O_261,N_2411,N_2492);
or UO_262 (O_262,N_2141,N_2291);
and UO_263 (O_263,N_2866,N_2637);
nor UO_264 (O_264,N_2490,N_2610);
nor UO_265 (O_265,N_2387,N_2268);
and UO_266 (O_266,N_2410,N_2180);
or UO_267 (O_267,N_2772,N_2405);
nand UO_268 (O_268,N_2236,N_2136);
or UO_269 (O_269,N_2327,N_2769);
nor UO_270 (O_270,N_2307,N_2295);
nor UO_271 (O_271,N_2629,N_2049);
nor UO_272 (O_272,N_2462,N_2660);
or UO_273 (O_273,N_2851,N_2725);
and UO_274 (O_274,N_2806,N_2583);
nor UO_275 (O_275,N_2857,N_2142);
or UO_276 (O_276,N_2910,N_2680);
or UO_277 (O_277,N_2483,N_2512);
or UO_278 (O_278,N_2471,N_2245);
and UO_279 (O_279,N_2272,N_2045);
and UO_280 (O_280,N_2033,N_2183);
and UO_281 (O_281,N_2599,N_2151);
and UO_282 (O_282,N_2091,N_2244);
nand UO_283 (O_283,N_2003,N_2813);
nand UO_284 (O_284,N_2874,N_2442);
nand UO_285 (O_285,N_2231,N_2156);
or UO_286 (O_286,N_2255,N_2775);
xor UO_287 (O_287,N_2709,N_2931);
nor UO_288 (O_288,N_2256,N_2993);
or UO_289 (O_289,N_2344,N_2160);
nand UO_290 (O_290,N_2306,N_2446);
nor UO_291 (O_291,N_2440,N_2146);
or UO_292 (O_292,N_2153,N_2555);
nor UO_293 (O_293,N_2437,N_2169);
nor UO_294 (O_294,N_2032,N_2331);
or UO_295 (O_295,N_2988,N_2648);
or UO_296 (O_296,N_2653,N_2959);
or UO_297 (O_297,N_2941,N_2340);
nand UO_298 (O_298,N_2630,N_2702);
or UO_299 (O_299,N_2102,N_2600);
or UO_300 (O_300,N_2363,N_2654);
and UO_301 (O_301,N_2081,N_2601);
and UO_302 (O_302,N_2924,N_2470);
nor UO_303 (O_303,N_2135,N_2985);
and UO_304 (O_304,N_2998,N_2279);
nor UO_305 (O_305,N_2028,N_2191);
or UO_306 (O_306,N_2206,N_2334);
nor UO_307 (O_307,N_2948,N_2283);
nand UO_308 (O_308,N_2473,N_2074);
or UO_309 (O_309,N_2721,N_2926);
nand UO_310 (O_310,N_2060,N_2967);
or UO_311 (O_311,N_2696,N_2338);
nand UO_312 (O_312,N_2793,N_2349);
or UO_313 (O_313,N_2898,N_2690);
nor UO_314 (O_314,N_2831,N_2491);
nor UO_315 (O_315,N_2550,N_2767);
or UO_316 (O_316,N_2860,N_2414);
and UO_317 (O_317,N_2190,N_2035);
and UO_318 (O_318,N_2569,N_2319);
nor UO_319 (O_319,N_2174,N_2467);
nand UO_320 (O_320,N_2647,N_2508);
nor UO_321 (O_321,N_2381,N_2303);
and UO_322 (O_322,N_2815,N_2019);
or UO_323 (O_323,N_2669,N_2010);
nand UO_324 (O_324,N_2194,N_2299);
nand UO_325 (O_325,N_2395,N_2357);
nand UO_326 (O_326,N_2578,N_2369);
and UO_327 (O_327,N_2148,N_2561);
and UO_328 (O_328,N_2787,N_2326);
and UO_329 (O_329,N_2684,N_2571);
nor UO_330 (O_330,N_2282,N_2057);
or UO_331 (O_331,N_2623,N_2124);
nand UO_332 (O_332,N_2661,N_2773);
nor UO_333 (O_333,N_2685,N_2330);
and UO_334 (O_334,N_2150,N_2172);
and UO_335 (O_335,N_2404,N_2927);
nand UO_336 (O_336,N_2524,N_2896);
nor UO_337 (O_337,N_2090,N_2149);
or UO_338 (O_338,N_2075,N_2722);
and UO_339 (O_339,N_2290,N_2588);
nand UO_340 (O_340,N_2873,N_2375);
nand UO_341 (O_341,N_2914,N_2701);
or UO_342 (O_342,N_2173,N_2079);
or UO_343 (O_343,N_2841,N_2355);
and UO_344 (O_344,N_2712,N_2656);
nor UO_345 (O_345,N_2536,N_2495);
nor UO_346 (O_346,N_2478,N_2640);
and UO_347 (O_347,N_2241,N_2123);
or UO_348 (O_348,N_2260,N_2723);
and UO_349 (O_349,N_2673,N_2251);
nor UO_350 (O_350,N_2552,N_2888);
nor UO_351 (O_351,N_2549,N_2166);
and UO_352 (O_352,N_2356,N_2530);
nor UO_353 (O_353,N_2065,N_2662);
and UO_354 (O_354,N_2554,N_2597);
or UO_355 (O_355,N_2716,N_2413);
nand UO_356 (O_356,N_2024,N_2209);
nand UO_357 (O_357,N_2944,N_2103);
nand UO_358 (O_358,N_2528,N_2999);
nor UO_359 (O_359,N_2732,N_2248);
nand UO_360 (O_360,N_2368,N_2535);
and UO_361 (O_361,N_2529,N_2595);
or UO_362 (O_362,N_2545,N_2633);
or UO_363 (O_363,N_2592,N_2479);
and UO_364 (O_364,N_2226,N_2519);
nor UO_365 (O_365,N_2556,N_2362);
nand UO_366 (O_366,N_2314,N_2564);
or UO_367 (O_367,N_2650,N_2263);
or UO_368 (O_368,N_2096,N_2031);
or UO_369 (O_369,N_2408,N_2296);
nand UO_370 (O_370,N_2216,N_2285);
nor UO_371 (O_371,N_2064,N_2777);
nor UO_372 (O_372,N_2963,N_2453);
nor UO_373 (O_373,N_2367,N_2407);
nand UO_374 (O_374,N_2657,N_2855);
and UO_375 (O_375,N_2304,N_2969);
nor UO_376 (O_376,N_2229,N_2043);
or UO_377 (O_377,N_2372,N_2534);
nand UO_378 (O_378,N_2801,N_2009);
nor UO_379 (O_379,N_2853,N_2155);
nor UO_380 (O_380,N_2691,N_2758);
nor UO_381 (O_381,N_2848,N_2017);
and UO_382 (O_382,N_2426,N_2987);
and UO_383 (O_383,N_2481,N_2377);
or UO_384 (O_384,N_2110,N_2620);
and UO_385 (O_385,N_2636,N_2157);
nor UO_386 (O_386,N_2558,N_2021);
and UO_387 (O_387,N_2836,N_2480);
and UO_388 (O_388,N_2018,N_2345);
nand UO_389 (O_389,N_2370,N_2729);
nor UO_390 (O_390,N_2205,N_2025);
or UO_391 (O_391,N_2041,N_2425);
or UO_392 (O_392,N_2505,N_2576);
and UO_393 (O_393,N_2780,N_2679);
nand UO_394 (O_394,N_2301,N_2996);
or UO_395 (O_395,N_2038,N_2822);
nand UO_396 (O_396,N_2502,N_2015);
or UO_397 (O_397,N_2921,N_2317);
nor UO_398 (O_398,N_2611,N_2078);
nor UO_399 (O_399,N_2693,N_2765);
or UO_400 (O_400,N_2321,N_2280);
or UO_401 (O_401,N_2489,N_2120);
or UO_402 (O_402,N_2547,N_2371);
and UO_403 (O_403,N_2705,N_2199);
nor UO_404 (O_404,N_2287,N_2013);
or UO_405 (O_405,N_2676,N_2457);
and UO_406 (O_406,N_2794,N_2862);
nand UO_407 (O_407,N_2409,N_2498);
or UO_408 (O_408,N_2222,N_2672);
nand UO_409 (O_409,N_2312,N_2781);
or UO_410 (O_410,N_2587,N_2675);
and UO_411 (O_411,N_2796,N_2807);
nand UO_412 (O_412,N_2365,N_2607);
and UO_413 (O_413,N_2649,N_2499);
nor UO_414 (O_414,N_2134,N_2517);
nand UO_415 (O_415,N_2540,N_2717);
and UO_416 (O_416,N_2922,N_2645);
and UO_417 (O_417,N_2262,N_2419);
nand UO_418 (O_418,N_2214,N_2711);
or UO_419 (O_419,N_2809,N_2297);
and UO_420 (O_420,N_2086,N_2727);
nor UO_421 (O_421,N_2612,N_2336);
and UO_422 (O_422,N_2879,N_2646);
nand UO_423 (O_423,N_2881,N_2217);
and UO_424 (O_424,N_2692,N_2953);
or UO_425 (O_425,N_2450,N_2539);
and UO_426 (O_426,N_2868,N_2351);
or UO_427 (O_427,N_2961,N_2808);
nor UO_428 (O_428,N_2761,N_2320);
nor UO_429 (O_429,N_2104,N_2389);
xor UO_430 (O_430,N_2707,N_2542);
nand UO_431 (O_431,N_2109,N_2568);
nor UO_432 (O_432,N_2050,N_2553);
xor UO_433 (O_433,N_2930,N_2942);
and UO_434 (O_434,N_2983,N_2008);
or UO_435 (O_435,N_2458,N_2752);
nor UO_436 (O_436,N_2071,N_2311);
or UO_437 (O_437,N_2276,N_2463);
and UO_438 (O_438,N_2068,N_2431);
nand UO_439 (O_439,N_2608,N_2412);
nor UO_440 (O_440,N_2570,N_2001);
and UO_441 (O_441,N_2981,N_2181);
or UO_442 (O_442,N_2766,N_2223);
and UO_443 (O_443,N_2083,N_2735);
nor UO_444 (O_444,N_2622,N_2247);
and UO_445 (O_445,N_2503,N_2940);
or UO_446 (O_446,N_2101,N_2358);
or UO_447 (O_447,N_2708,N_2703);
or UO_448 (O_448,N_2894,N_2474);
and UO_449 (O_449,N_2688,N_2560);
and UO_450 (O_450,N_2485,N_2070);
nand UO_451 (O_451,N_2300,N_2580);
or UO_452 (O_452,N_2594,N_2006);
nor UO_453 (O_453,N_2464,N_2783);
or UO_454 (O_454,N_2269,N_2284);
and UO_455 (O_455,N_2525,N_2854);
or UO_456 (O_456,N_2140,N_2393);
nor UO_457 (O_457,N_2077,N_2315);
or UO_458 (O_458,N_2859,N_2027);
and UO_459 (O_459,N_2042,N_2593);
nand UO_460 (O_460,N_2596,N_2730);
xnor UO_461 (O_461,N_2915,N_2674);
nor UO_462 (O_462,N_2219,N_2323);
or UO_463 (O_463,N_2448,N_2193);
or UO_464 (O_464,N_2184,N_2497);
nand UO_465 (O_465,N_2225,N_2252);
and UO_466 (O_466,N_2837,N_2072);
or UO_467 (O_467,N_2313,N_2052);
and UO_468 (O_468,N_2832,N_2445);
or UO_469 (O_469,N_2624,N_2270);
and UO_470 (O_470,N_2228,N_2347);
and UO_471 (O_471,N_2997,N_2741);
and UO_472 (O_472,N_2144,N_2504);
or UO_473 (O_473,N_2923,N_2658);
and UO_474 (O_474,N_2635,N_2697);
or UO_475 (O_475,N_2800,N_2937);
xnor UO_476 (O_476,N_2605,N_2818);
and UO_477 (O_477,N_2238,N_2805);
or UO_478 (O_478,N_2016,N_2088);
nand UO_479 (O_479,N_2965,N_2046);
or UO_480 (O_480,N_2020,N_2105);
nand UO_481 (O_481,N_2383,N_2572);
nor UO_482 (O_482,N_2082,N_2441);
and UO_483 (O_483,N_2302,N_2681);
nand UO_484 (O_484,N_2128,N_2476);
or UO_485 (O_485,N_2843,N_2207);
nor UO_486 (O_486,N_2804,N_2811);
or UO_487 (O_487,N_2904,N_2586);
and UO_488 (O_488,N_2774,N_2694);
or UO_489 (O_489,N_2415,N_2689);
and UO_490 (O_490,N_2484,N_2147);
nor UO_491 (O_491,N_2905,N_2292);
nor UO_492 (O_492,N_2275,N_2218);
and UO_493 (O_493,N_2211,N_2892);
or UO_494 (O_494,N_2893,N_2562);
or UO_495 (O_495,N_2309,N_2949);
and UO_496 (O_496,N_2602,N_2364);
or UO_497 (O_497,N_2427,N_2890);
nand UO_498 (O_498,N_2221,N_2933);
and UO_499 (O_499,N_2452,N_2738);
endmodule