module basic_1500_15000_2000_15_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1145,In_1076);
nand U1 (N_1,In_650,In_582);
nand U2 (N_2,In_665,In_878);
and U3 (N_3,In_1220,In_170);
or U4 (N_4,In_965,In_385);
or U5 (N_5,In_972,In_709);
or U6 (N_6,In_378,In_1128);
nor U7 (N_7,In_1175,In_419);
nand U8 (N_8,In_1137,In_386);
nor U9 (N_9,In_1058,In_375);
nand U10 (N_10,In_106,In_1084);
or U11 (N_11,In_1404,In_1494);
or U12 (N_12,In_417,In_584);
nand U13 (N_13,In_1050,In_169);
and U14 (N_14,In_1386,In_185);
nand U15 (N_15,In_672,In_260);
nand U16 (N_16,In_1185,In_1209);
and U17 (N_17,In_1401,In_432);
nand U18 (N_18,In_610,In_1090);
or U19 (N_19,In_588,In_937);
nand U20 (N_20,In_431,In_873);
nor U21 (N_21,In_1405,In_583);
and U22 (N_22,In_1125,In_59);
and U23 (N_23,In_1206,In_563);
or U24 (N_24,In_805,In_196);
or U25 (N_25,In_90,In_1457);
and U26 (N_26,In_1342,In_1469);
or U27 (N_27,In_1025,In_806);
and U28 (N_28,In_502,In_427);
nor U29 (N_29,In_1049,In_92);
nand U30 (N_30,In_819,In_18);
or U31 (N_31,In_353,In_403);
xor U32 (N_32,In_1416,In_291);
nand U33 (N_33,In_576,In_985);
nand U34 (N_34,In_1020,In_783);
nand U35 (N_35,In_1104,In_1086);
nor U36 (N_36,In_1311,In_737);
nor U37 (N_37,In_430,In_1066);
or U38 (N_38,In_681,In_961);
and U39 (N_39,In_158,In_1451);
nand U40 (N_40,In_578,In_587);
nor U41 (N_41,In_1148,In_405);
and U42 (N_42,In_16,In_296);
nand U43 (N_43,In_590,In_960);
and U44 (N_44,In_705,In_1272);
or U45 (N_45,In_964,In_1171);
and U46 (N_46,In_504,In_199);
nand U47 (N_47,In_1256,In_210);
nand U48 (N_48,In_914,In_597);
or U49 (N_49,In_1307,In_532);
xor U50 (N_50,In_1345,In_861);
and U51 (N_51,In_290,In_855);
or U52 (N_52,In_868,In_990);
nand U53 (N_53,In_1030,In_686);
and U54 (N_54,In_315,In_332);
nor U55 (N_55,In_355,In_1190);
nor U56 (N_56,In_486,In_226);
nand U57 (N_57,In_1078,In_724);
and U58 (N_58,In_903,In_482);
nor U59 (N_59,In_178,In_1458);
and U60 (N_60,In_1394,In_1279);
and U61 (N_61,In_86,In_1268);
nand U62 (N_62,In_358,In_690);
nor U63 (N_63,In_815,In_771);
or U64 (N_64,In_377,In_391);
nand U65 (N_65,In_1036,In_1324);
or U66 (N_66,In_1061,In_768);
or U67 (N_67,In_21,In_182);
nor U68 (N_68,In_693,In_1479);
or U69 (N_69,In_264,In_494);
and U70 (N_70,In_909,In_943);
or U71 (N_71,In_817,In_944);
nand U72 (N_72,In_525,In_1285);
nor U73 (N_73,In_76,In_1046);
nand U74 (N_74,In_1127,In_946);
nor U75 (N_75,In_1444,In_697);
or U76 (N_76,In_956,In_1181);
xor U77 (N_77,In_533,In_1067);
or U78 (N_78,In_850,In_606);
or U79 (N_79,In_623,In_1192);
nand U80 (N_80,In_429,In_320);
nor U81 (N_81,In_269,In_188);
nor U82 (N_82,In_639,In_1143);
and U83 (N_83,In_889,In_1364);
or U84 (N_84,In_495,In_1158);
or U85 (N_85,In_364,In_721);
nand U86 (N_86,In_554,In_97);
or U87 (N_87,In_67,In_428);
nor U88 (N_88,In_1093,In_140);
and U89 (N_89,In_668,In_537);
nand U90 (N_90,In_22,In_1456);
and U91 (N_91,In_785,In_661);
nand U92 (N_92,In_1473,In_1227);
and U93 (N_93,In_1368,In_469);
nand U94 (N_94,In_1026,In_120);
and U95 (N_95,In_1004,In_932);
or U96 (N_96,In_336,In_1480);
nand U97 (N_97,In_401,In_957);
nand U98 (N_98,In_715,In_294);
nand U99 (N_99,In_1033,In_774);
or U100 (N_100,In_52,In_454);
nor U101 (N_101,In_1338,In_833);
or U102 (N_102,In_548,In_841);
or U103 (N_103,In_1083,In_859);
nand U104 (N_104,In_547,In_1297);
and U105 (N_105,In_155,In_1244);
nor U106 (N_106,In_284,In_1400);
nand U107 (N_107,In_297,In_1440);
nor U108 (N_108,In_820,In_238);
nor U109 (N_109,In_1426,In_314);
nor U110 (N_110,In_637,In_176);
nand U111 (N_111,In_995,In_1482);
and U112 (N_112,In_886,In_627);
and U113 (N_113,In_1048,In_232);
or U114 (N_114,In_1197,In_1115);
or U115 (N_115,In_349,In_1402);
or U116 (N_116,In_1374,In_826);
nand U117 (N_117,In_1252,In_477);
and U118 (N_118,In_398,In_986);
nor U119 (N_119,In_1077,In_74);
or U120 (N_120,In_1396,In_1051);
and U121 (N_121,In_1024,In_53);
and U122 (N_122,In_246,In_891);
nand U123 (N_123,In_1159,In_730);
and U124 (N_124,In_271,In_911);
and U125 (N_125,In_757,In_302);
or U126 (N_126,In_784,In_1113);
and U127 (N_127,In_114,In_1210);
nand U128 (N_128,In_1273,In_83);
nor U129 (N_129,In_519,In_1047);
nor U130 (N_130,In_1132,In_1362);
and U131 (N_131,In_950,In_1496);
nor U132 (N_132,In_259,In_234);
nand U133 (N_133,In_838,In_84);
and U134 (N_134,In_435,In_179);
nand U135 (N_135,In_133,In_1350);
or U136 (N_136,In_490,In_604);
or U137 (N_137,In_858,In_272);
or U138 (N_138,In_760,In_871);
nor U139 (N_139,In_94,In_330);
or U140 (N_140,In_483,In_183);
nor U141 (N_141,In_275,In_1208);
and U142 (N_142,In_642,In_1341);
or U143 (N_143,In_982,In_581);
or U144 (N_144,In_1441,In_550);
nand U145 (N_145,In_602,In_1151);
or U146 (N_146,In_892,In_634);
or U147 (N_147,In_1205,In_1277);
or U148 (N_148,In_927,In_1028);
and U149 (N_149,In_465,In_98);
nand U150 (N_150,In_599,In_1261);
nor U151 (N_151,In_1196,In_93);
and U152 (N_152,In_99,In_1382);
nor U153 (N_153,In_162,In_849);
and U154 (N_154,In_569,In_1081);
nand U155 (N_155,In_874,In_773);
and U156 (N_156,In_571,In_794);
and U157 (N_157,In_1359,In_1477);
or U158 (N_158,In_372,In_319);
nand U159 (N_159,In_613,In_3);
nand U160 (N_160,In_896,In_1488);
nor U161 (N_161,In_1318,In_1212);
or U162 (N_162,In_251,In_1353);
or U163 (N_163,In_1008,In_292);
nand U164 (N_164,In_1054,In_7);
or U165 (N_165,In_161,In_60);
nor U166 (N_166,In_68,In_1162);
nor U167 (N_167,In_762,In_632);
or U168 (N_168,In_725,In_1468);
nor U169 (N_169,In_440,In_1089);
or U170 (N_170,In_312,In_611);
nor U171 (N_171,In_1486,In_1329);
nand U172 (N_172,In_173,In_735);
nor U173 (N_173,In_1410,In_1134);
nor U174 (N_174,In_24,In_1327);
and U175 (N_175,In_870,In_1408);
nand U176 (N_176,In_1186,In_553);
nand U177 (N_177,In_1356,In_1021);
nand U178 (N_178,In_126,In_1073);
nand U179 (N_179,In_749,In_575);
and U180 (N_180,In_216,In_1436);
nor U181 (N_181,In_2,In_231);
nor U182 (N_182,In_285,In_603);
and U183 (N_183,In_1462,In_478);
nand U184 (N_184,In_1027,In_273);
and U185 (N_185,In_283,In_148);
nor U186 (N_186,In_1224,In_1225);
or U187 (N_187,In_526,In_729);
nor U188 (N_188,In_1460,In_968);
nor U189 (N_189,In_822,In_1429);
nand U190 (N_190,In_1152,In_952);
nor U191 (N_191,In_306,In_1248);
and U192 (N_192,In_262,In_1012);
nand U193 (N_193,In_100,In_835);
and U194 (N_194,In_840,In_1263);
nor U195 (N_195,In_828,In_712);
or U196 (N_196,In_1161,In_1366);
nand U197 (N_197,In_1249,In_1317);
and U198 (N_198,In_804,In_37);
or U199 (N_199,In_71,In_56);
or U200 (N_200,In_288,In_464);
and U201 (N_201,In_1120,In_1387);
and U202 (N_202,In_1337,In_769);
and U203 (N_203,In_411,In_1393);
and U204 (N_204,In_159,In_1160);
nor U205 (N_205,In_786,In_181);
or U206 (N_206,In_827,In_119);
or U207 (N_207,In_48,In_186);
nand U208 (N_208,In_1465,In_609);
or U209 (N_209,In_782,In_1139);
nor U210 (N_210,In_123,In_1129);
or U211 (N_211,In_667,In_395);
or U212 (N_212,In_1310,In_888);
and U213 (N_213,In_625,In_261);
and U214 (N_214,In_125,In_747);
nand U215 (N_215,In_1322,In_508);
nand U216 (N_216,In_802,In_876);
nor U217 (N_217,In_546,In_540);
nor U218 (N_218,In_605,In_1235);
nand U219 (N_219,In_141,In_118);
nor U220 (N_220,In_363,In_46);
or U221 (N_221,In_880,In_1023);
nor U222 (N_222,In_1278,In_890);
or U223 (N_223,In_751,In_683);
and U224 (N_224,In_542,In_206);
nand U225 (N_225,In_58,In_865);
nor U226 (N_226,In_1,In_39);
nand U227 (N_227,In_1116,In_701);
nor U228 (N_228,In_115,In_474);
nand U229 (N_229,In_1442,In_1122);
nor U230 (N_230,In_414,In_1299);
nand U231 (N_231,In_1424,In_789);
nor U232 (N_232,In_117,In_1022);
nand U233 (N_233,In_561,In_334);
nand U234 (N_234,In_331,In_763);
nor U235 (N_235,In_1379,In_1068);
and U236 (N_236,In_1373,In_1014);
and U237 (N_237,In_1259,In_26);
or U238 (N_238,In_1016,In_1443);
nand U239 (N_239,In_795,In_274);
nor U240 (N_240,In_1371,In_1281);
nor U241 (N_241,In_257,In_921);
or U242 (N_242,In_174,In_1439);
nor U243 (N_243,In_1369,In_1323);
and U244 (N_244,In_493,In_479);
and U245 (N_245,In_416,In_70);
nor U246 (N_246,In_289,In_127);
nor U247 (N_247,In_759,In_1040);
or U248 (N_248,In_351,In_298);
and U249 (N_249,In_679,In_799);
or U250 (N_250,In_452,In_387);
nor U251 (N_251,In_824,In_1301);
nand U252 (N_252,In_1001,In_645);
and U253 (N_253,In_704,In_79);
or U254 (N_254,In_823,In_1094);
and U255 (N_255,In_967,In_1298);
and U256 (N_256,In_433,In_947);
and U257 (N_257,In_212,In_1108);
nand U258 (N_258,In_902,In_406);
nor U259 (N_259,In_505,In_713);
nand U260 (N_260,In_1430,In_574);
nor U261 (N_261,In_139,In_445);
or U262 (N_262,In_359,In_720);
or U263 (N_263,In_1167,In_1293);
or U264 (N_264,In_1126,In_1257);
nor U265 (N_265,In_598,In_233);
or U266 (N_266,In_1111,In_558);
xor U267 (N_267,In_1214,In_191);
and U268 (N_268,In_612,In_1358);
nor U269 (N_269,In_1110,In_1413);
nor U270 (N_270,In_1045,In_1131);
or U271 (N_271,In_205,In_1250);
and U272 (N_272,In_128,In_1392);
nor U273 (N_273,In_566,In_1384);
and U274 (N_274,In_881,In_654);
and U275 (N_275,In_356,In_778);
nand U276 (N_276,In_851,In_116);
and U277 (N_277,In_1072,In_1085);
or U278 (N_278,In_511,In_328);
and U279 (N_279,In_236,In_14);
and U280 (N_280,In_662,In_1437);
nand U281 (N_281,In_136,In_731);
nand U282 (N_282,In_1173,In_1106);
nor U283 (N_283,In_281,In_1388);
and U284 (N_284,In_938,In_893);
nand U285 (N_285,In_1182,In_1464);
or U286 (N_286,In_209,In_1497);
or U287 (N_287,In_644,In_197);
or U288 (N_288,In_339,In_614);
nor U289 (N_289,In_897,In_1280);
and U290 (N_290,In_1255,In_282);
and U291 (N_291,In_1080,In_1476);
nand U292 (N_292,In_1370,In_1253);
nor U293 (N_293,In_481,In_1157);
and U294 (N_294,In_1450,In_211);
nor U295 (N_295,In_168,In_753);
nand U296 (N_296,In_543,In_223);
and U297 (N_297,In_1383,In_696);
nand U298 (N_298,In_253,In_976);
nor U299 (N_299,In_714,In_1150);
nor U300 (N_300,In_676,In_1319);
nor U301 (N_301,In_402,In_577);
nor U302 (N_302,In_919,In_908);
nand U303 (N_303,In_1155,In_468);
nand U304 (N_304,In_863,In_1289);
or U305 (N_305,In_338,In_1215);
and U306 (N_306,In_517,In_258);
nor U307 (N_307,In_1275,In_916);
and U308 (N_308,In_1291,In_1109);
nand U309 (N_309,In_516,In_45);
or U310 (N_310,In_928,In_506);
nor U311 (N_311,In_549,In_245);
nor U312 (N_312,In_1349,In_1245);
or U313 (N_313,In_1467,In_1459);
or U314 (N_314,In_1361,In_163);
and U315 (N_315,In_779,In_1308);
or U316 (N_316,In_974,In_164);
and U317 (N_317,In_448,In_1242);
nor U318 (N_318,In_1236,In_1103);
and U319 (N_319,In_534,In_1487);
nor U320 (N_320,In_572,In_792);
or U321 (N_321,In_1355,In_663);
nor U322 (N_322,In_1455,In_1075);
or U323 (N_323,In_1178,In_180);
and U324 (N_324,In_453,In_772);
or U325 (N_325,In_807,In_1218);
nand U326 (N_326,In_177,In_241);
nand U327 (N_327,In_1052,In_514);
nand U328 (N_328,In_1056,In_963);
or U329 (N_329,In_1112,In_151);
and U330 (N_330,In_423,In_1203);
nor U331 (N_331,In_1217,In_394);
or U332 (N_332,In_224,In_1428);
nor U333 (N_333,In_744,In_203);
nor U334 (N_334,In_781,In_1495);
nor U335 (N_335,In_1414,In_1395);
and U336 (N_336,In_821,In_905);
nand U337 (N_337,In_652,In_9);
and U338 (N_338,In_912,In_1348);
nand U339 (N_339,In_507,In_872);
nand U340 (N_340,In_383,In_631);
and U341 (N_341,In_1309,In_1397);
and U342 (N_342,In_248,In_646);
and U343 (N_343,In_346,In_198);
or U344 (N_344,In_1191,In_501);
and U345 (N_345,In_1062,In_948);
nand U346 (N_346,In_217,In_393);
and U347 (N_347,In_175,In_102);
and U348 (N_348,In_1032,In_635);
and U349 (N_349,In_643,In_616);
nand U350 (N_350,In_521,In_408);
or U351 (N_351,In_201,In_740);
and U352 (N_352,In_955,In_675);
or U353 (N_353,In_329,In_1195);
and U354 (N_354,In_869,In_1042);
or U355 (N_355,In_310,In_237);
nand U356 (N_356,In_1474,In_450);
or U357 (N_357,In_62,In_29);
or U358 (N_358,In_655,In_980);
or U359 (N_359,In_10,In_1069);
nor U360 (N_360,In_702,In_854);
and U361 (N_361,In_787,In_1053);
or U362 (N_362,In_499,In_1452);
nor U363 (N_363,In_28,In_299);
nand U364 (N_364,In_1485,In_1241);
or U365 (N_365,In_293,In_1119);
nor U366 (N_366,In_57,In_410);
nor U367 (N_367,In_1156,In_814);
and U368 (N_368,In_51,In_85);
nor U369 (N_369,In_879,In_1180);
nor U370 (N_370,In_1377,In_682);
and U371 (N_371,In_728,In_997);
nor U372 (N_372,In_1313,In_220);
nand U373 (N_373,In_286,In_1246);
and U374 (N_374,In_1039,In_318);
or U375 (N_375,In_134,In_1340);
nand U376 (N_376,In_108,In_31);
nor U377 (N_377,In_555,In_1211);
nor U378 (N_378,In_1170,In_472);
and U379 (N_379,In_1425,In_1399);
nor U380 (N_380,In_898,In_222);
and U381 (N_381,In_1347,In_1484);
nand U382 (N_382,In_512,In_1326);
or U383 (N_383,In_63,In_620);
and U384 (N_384,In_981,In_930);
nor U385 (N_385,In_1493,In_424);
and U386 (N_386,In_818,In_658);
or U387 (N_387,In_727,In_1071);
nand U388 (N_388,In_137,In_907);
and U389 (N_389,In_716,In_901);
nor U390 (N_390,In_829,In_492);
or U391 (N_391,In_601,In_885);
nand U392 (N_392,In_303,In_848);
nor U393 (N_393,In_834,In_308);
or U394 (N_394,In_1481,In_915);
nand U395 (N_395,In_515,In_1189);
nor U396 (N_396,In_741,In_305);
or U397 (N_397,In_711,In_931);
or U398 (N_398,In_726,In_167);
and U399 (N_399,In_365,In_962);
or U400 (N_400,In_884,In_970);
or U401 (N_401,In_992,In_678);
nand U402 (N_402,In_754,In_1018);
and U403 (N_403,In_689,In_309);
and U404 (N_404,In_129,In_498);
and U405 (N_405,In_1304,In_208);
nor U406 (N_406,In_1124,In_692);
and U407 (N_407,In_1463,In_770);
nor U408 (N_408,In_524,In_500);
or U409 (N_409,In_1184,In_47);
nand U410 (N_410,In_449,In_1019);
or U411 (N_411,In_347,In_1163);
nor U412 (N_412,In_313,In_1146);
nor U413 (N_413,In_1398,In_670);
nor U414 (N_414,In_1409,In_695);
nand U415 (N_415,In_451,In_370);
nor U416 (N_416,In_1063,In_1238);
nand U417 (N_417,In_1375,In_409);
and U418 (N_418,In_791,In_1000);
and U419 (N_419,In_993,In_593);
nand U420 (N_420,In_700,In_766);
nor U421 (N_421,In_81,In_1165);
nor U422 (N_422,In_1312,In_1251);
and U423 (N_423,In_925,In_918);
nand U424 (N_424,In_1445,In_520);
nand U425 (N_425,In_1207,In_1095);
and U426 (N_426,In_69,In_1471);
or U427 (N_427,In_485,In_570);
and U428 (N_428,In_361,In_1449);
nor U429 (N_429,In_926,In_988);
nand U430 (N_430,In_628,In_75);
and U431 (N_431,In_674,In_987);
or U432 (N_432,In_130,In_1390);
nor U433 (N_433,In_883,In_1328);
or U434 (N_434,In_1204,In_1264);
nand U435 (N_435,In_811,In_1117);
nor U436 (N_436,In_382,In_1100);
xnor U437 (N_437,In_641,In_1346);
nand U438 (N_438,In_1079,In_941);
and U439 (N_439,In_1226,In_444);
nor U440 (N_440,In_710,In_1199);
and U441 (N_441,In_311,In_1057);
and U442 (N_442,In_666,In_1176);
and U443 (N_443,In_373,In_1043);
or U444 (N_444,In_1492,In_1188);
nand U445 (N_445,In_187,In_88);
nand U446 (N_446,In_156,In_266);
nand U447 (N_447,In_1360,In_977);
nor U448 (N_448,In_935,In_636);
xnor U449 (N_449,In_552,In_1138);
or U450 (N_450,In_1070,In_1265);
or U451 (N_451,In_812,In_326);
nand U452 (N_452,In_1130,In_559);
nor U453 (N_453,In_121,In_456);
and U454 (N_454,In_1454,In_421);
and U455 (N_455,In_1461,In_708);
or U456 (N_456,In_810,In_743);
nand U457 (N_457,In_40,In_699);
and U458 (N_458,In_1035,In_1006);
and U459 (N_459,In_219,In_752);
and U460 (N_460,In_484,In_1029);
or U461 (N_461,In_202,In_857);
nor U462 (N_462,In_1060,In_1088);
nand U463 (N_463,In_1365,In_1219);
nor U464 (N_464,In_240,In_1201);
and U465 (N_465,In_276,In_160);
and U466 (N_466,In_354,In_23);
and U467 (N_467,In_304,In_1331);
nand U468 (N_468,In_473,In_1343);
nand U469 (N_469,In_418,In_12);
nand U470 (N_470,In_256,In_529);
or U471 (N_471,In_1295,In_415);
nor U472 (N_472,In_287,In_846);
or U473 (N_473,In_573,In_527);
and U474 (N_474,In_594,In_1168);
nor U475 (N_475,In_560,In_638);
or U476 (N_476,In_797,In_213);
or U477 (N_477,In_425,In_1269);
nand U478 (N_478,In_1288,In_470);
nand U479 (N_479,In_1260,In_413);
nor U480 (N_480,In_143,In_44);
or U481 (N_481,In_1417,In_1475);
nor U482 (N_482,In_407,In_476);
nor U483 (N_483,In_1223,In_777);
nand U484 (N_484,In_562,In_882);
or U485 (N_485,In_860,In_669);
and U486 (N_486,In_746,In_321);
nand U487 (N_487,In_30,In_1351);
nor U488 (N_488,In_580,In_89);
and U489 (N_489,In_1101,In_1240);
or U490 (N_490,In_1372,In_255);
nand U491 (N_491,In_564,In_192);
and U492 (N_492,In_32,In_112);
nor U493 (N_493,In_278,In_836);
and U494 (N_494,In_1009,In_11);
and U495 (N_495,In_996,In_979);
nor U496 (N_496,In_971,In_842);
nor U497 (N_497,In_780,In_250);
nor U498 (N_498,In_664,In_487);
nand U499 (N_499,In_1325,In_0);
nor U500 (N_500,In_1011,In_323);
nor U501 (N_501,In_324,In_640);
nor U502 (N_502,In_1284,In_165);
nand U503 (N_503,In_808,In_335);
and U504 (N_504,In_1421,In_913);
nand U505 (N_505,In_270,In_1017);
nand U506 (N_506,In_422,In_719);
nand U507 (N_507,In_390,In_1276);
and U508 (N_508,In_54,In_138);
nand U509 (N_509,In_239,In_1216);
or U510 (N_510,In_940,In_135);
nor U511 (N_511,In_1232,In_837);
or U512 (N_512,In_455,In_1228);
nand U513 (N_513,In_388,In_327);
or U514 (N_514,In_1306,In_556);
or U515 (N_515,In_742,In_325);
and U516 (N_516,In_1147,In_647);
nand U517 (N_517,In_798,In_1169);
and U518 (N_518,In_78,In_1303);
nor U519 (N_519,In_618,In_586);
or U520 (N_520,In_152,In_1332);
and U521 (N_521,In_518,In_371);
nand U522 (N_522,In_366,In_154);
nor U523 (N_523,In_1041,In_687);
nor U524 (N_524,In_1320,In_1490);
nor U525 (N_525,In_190,In_193);
or U526 (N_526,In_252,In_1183);
or U527 (N_527,In_439,In_497);
nor U528 (N_528,In_989,In_242);
or U529 (N_529,In_150,In_1038);
nor U530 (N_530,In_489,In_442);
nor U531 (N_531,In_793,In_43);
nand U532 (N_532,In_1003,In_1007);
nand U533 (N_533,In_959,In_922);
nor U534 (N_534,In_816,In_557);
and U535 (N_535,In_723,In_530);
and U536 (N_536,In_852,In_1098);
nand U537 (N_537,In_934,In_215);
nand U538 (N_538,In_82,In_607);
nand U539 (N_539,In_660,In_171);
and U540 (N_540,In_1380,In_803);
or U541 (N_541,In_1385,In_184);
nor U542 (N_542,In_1415,In_933);
nand U543 (N_543,In_844,In_153);
nand U544 (N_544,In_333,In_579);
nand U545 (N_545,In_839,In_194);
nor U546 (N_546,In_1258,In_1198);
nor U547 (N_547,In_350,In_685);
and U548 (N_548,In_619,In_466);
and U549 (N_549,In_856,In_380);
nand U550 (N_550,In_434,In_756);
and U551 (N_551,In_1002,In_568);
nor U552 (N_552,In_1221,In_1412);
nand U553 (N_553,In_38,In_42);
nor U554 (N_554,In_734,In_953);
or U555 (N_555,In_1321,In_441);
nor U556 (N_556,In_446,In_247);
nor U557 (N_557,In_1407,In_55);
nand U558 (N_558,In_458,In_34);
or U559 (N_559,In_1453,In_671);
and U560 (N_560,In_738,In_8);
xnor U561 (N_561,In_369,In_800);
and U562 (N_562,In_596,In_225);
and U563 (N_563,In_204,In_1031);
or U564 (N_564,In_788,In_345);
and U565 (N_565,In_265,In_301);
or U566 (N_566,In_1064,In_624);
nand U567 (N_567,In_951,In_228);
and U568 (N_568,In_866,In_1433);
xor U569 (N_569,In_389,In_813);
and U570 (N_570,In_1287,In_910);
or U571 (N_571,In_745,In_249);
nor U572 (N_572,In_1107,In_739);
nor U573 (N_573,In_25,In_1334);
nand U574 (N_574,In_1333,In_949);
and U575 (N_575,In_677,In_1123);
xor U576 (N_576,In_1121,In_475);
nor U577 (N_577,In_867,In_622);
or U578 (N_578,In_1427,In_541);
or U579 (N_579,In_733,In_4);
nor U580 (N_580,In_367,In_96);
and U581 (N_581,In_900,In_101);
or U582 (N_582,In_929,In_617);
nand U583 (N_583,In_592,In_6);
nand U584 (N_584,In_457,In_1118);
or U585 (N_585,In_1435,In_35);
and U586 (N_586,In_809,In_999);
nand U587 (N_587,In_142,In_267);
and U588 (N_588,In_91,In_1065);
and U589 (N_589,In_864,In_105);
and U590 (N_590,In_973,In_61);
nand U591 (N_591,In_1213,In_1357);
and U592 (N_592,In_1335,In_1270);
and U593 (N_593,In_1254,In_1294);
and U594 (N_594,In_397,In_923);
nand U595 (N_595,In_1438,In_122);
nand U596 (N_596,In_1286,In_906);
or U597 (N_597,In_1391,In_706);
nand U598 (N_598,In_221,In_1247);
or U599 (N_599,In_467,In_1411);
nand U600 (N_600,In_280,In_1179);
nor U601 (N_601,In_894,In_1172);
nand U602 (N_602,In_945,In_157);
or U603 (N_603,In_887,In_1420);
nand U604 (N_604,In_522,In_404);
nor U605 (N_605,In_942,In_1314);
or U606 (N_606,In_384,In_1447);
nor U607 (N_607,In_368,In_1339);
nor U608 (N_608,In_608,In_1153);
nand U609 (N_609,In_796,In_1352);
or U610 (N_610,In_362,In_830);
and U611 (N_611,In_1133,In_316);
or U612 (N_612,In_1499,In_875);
or U613 (N_613,In_218,In_983);
nor U614 (N_614,In_718,In_994);
and U615 (N_615,In_437,In_899);
nor U616 (N_616,In_936,In_1082);
or U617 (N_617,In_1166,In_1200);
and U618 (N_618,In_775,In_144);
and U619 (N_619,In_459,In_966);
nand U620 (N_620,In_1202,In_147);
or U621 (N_621,In_764,In_924);
nand U622 (N_622,In_1034,In_621);
nor U623 (N_623,In_1418,In_1174);
or U624 (N_624,In_954,In_1194);
nand U625 (N_625,In_322,In_656);
and U626 (N_626,In_1096,In_189);
nor U627 (N_627,In_357,In_13);
nand U628 (N_628,In_615,In_244);
or U629 (N_629,In_1282,In_1367);
or U630 (N_630,In_984,In_491);
or U631 (N_631,In_1091,In_166);
and U632 (N_632,In_761,In_503);
nor U633 (N_633,In_107,In_659);
nand U634 (N_634,In_348,In_254);
nand U635 (N_635,In_1262,In_591);
nor U636 (N_636,In_268,In_567);
or U637 (N_637,In_991,In_649);
nand U638 (N_638,In_400,In_399);
or U639 (N_639,In_1381,In_847);
nor U640 (N_640,In_195,In_72);
or U641 (N_641,In_691,In_132);
xnor U642 (N_642,In_1419,In_1243);
nor U643 (N_643,In_243,In_626);
nand U644 (N_644,In_131,In_703);
nand U645 (N_645,In_230,In_488);
nor U646 (N_646,In_509,In_1274);
nor U647 (N_647,In_27,In_767);
nand U648 (N_648,In_41,In_1378);
and U649 (N_649,In_717,In_460);
nor U650 (N_650,In_300,In_825);
nor U651 (N_651,In_831,In_1431);
or U652 (N_652,In_461,In_1491);
nor U653 (N_653,In_1044,In_633);
or U654 (N_654,In_1292,In_657);
and U655 (N_655,In_531,In_1354);
nand U656 (N_656,In_1013,In_17);
nor U657 (N_657,In_381,In_279);
nand U658 (N_658,In_1144,In_110);
nand U659 (N_659,In_1266,In_688);
and U660 (N_660,In_998,In_673);
nand U661 (N_661,In_1271,In_801);
nor U662 (N_662,In_342,In_392);
nand U663 (N_663,In_600,In_1302);
or U664 (N_664,In_65,In_969);
nand U665 (N_665,In_1315,In_1037);
nor U666 (N_666,In_565,In_109);
and U667 (N_667,In_1105,In_1434);
nor U668 (N_668,In_589,In_1233);
nand U669 (N_669,In_340,In_1403);
or U670 (N_670,In_111,In_104);
and U671 (N_671,In_5,In_344);
nor U672 (N_672,In_1239,In_630);
nor U673 (N_673,In_50,In_1448);
nor U674 (N_674,In_1234,In_651);
nand U675 (N_675,In_975,In_755);
nor U676 (N_676,In_510,In_426);
nor U677 (N_677,In_1283,In_722);
nor U678 (N_678,In_352,In_1154);
or U679 (N_679,In_1055,In_535);
and U680 (N_680,In_146,In_758);
nor U681 (N_681,In_19,In_513);
and U682 (N_682,In_1149,In_832);
nor U683 (N_683,In_420,In_447);
and U684 (N_684,In_480,In_227);
nand U685 (N_685,In_145,In_341);
or U686 (N_686,In_684,In_595);
and U687 (N_687,In_736,In_545);
or U688 (N_688,In_462,In_1290);
nand U689 (N_689,In_1432,In_33);
nand U690 (N_690,In_374,In_1466);
or U691 (N_691,In_412,In_904);
nor U692 (N_692,In_496,In_360);
or U693 (N_693,In_124,In_1330);
nor U694 (N_694,In_528,In_1423);
nand U695 (N_695,In_1230,In_748);
nor U696 (N_696,In_629,In_1114);
nand U697 (N_697,In_750,In_1472);
and U698 (N_698,In_698,In_471);
nand U699 (N_699,In_80,In_732);
nor U700 (N_700,In_1498,In_1422);
or U701 (N_701,In_694,In_1267);
nor U702 (N_702,In_653,In_877);
xor U703 (N_703,In_1136,In_1446);
or U704 (N_704,In_707,In_1097);
or U705 (N_705,In_1229,In_295);
and U706 (N_706,In_523,In_544);
and U707 (N_707,In_1222,In_1489);
or U708 (N_708,In_776,In_538);
nand U709 (N_709,In_1164,In_337);
nand U710 (N_710,In_1005,In_1336);
nor U711 (N_711,In_1015,In_1389);
nand U712 (N_712,In_149,In_680);
nand U713 (N_713,In_443,In_551);
nand U714 (N_714,In_77,In_920);
nor U715 (N_715,In_1142,In_172);
or U716 (N_716,In_66,In_1135);
or U717 (N_717,In_1376,In_1478);
or U718 (N_718,In_229,In_862);
nand U719 (N_719,In_853,In_536);
nand U720 (N_720,In_539,In_36);
nand U721 (N_721,In_1074,In_376);
nor U722 (N_722,In_277,In_585);
or U723 (N_723,In_1010,In_235);
nand U724 (N_724,In_1296,In_1092);
nand U725 (N_725,In_1300,In_1237);
or U726 (N_726,In_1231,In_1099);
nor U727 (N_727,In_1059,In_343);
nor U728 (N_728,In_317,In_1140);
and U729 (N_729,In_436,In_765);
and U730 (N_730,In_978,In_113);
nor U731 (N_731,In_843,In_463);
and U732 (N_732,In_648,In_1363);
and U733 (N_733,In_87,In_1177);
or U734 (N_734,In_1470,In_438);
or U735 (N_735,In_64,In_20);
nand U736 (N_736,In_200,In_1344);
and U737 (N_737,In_379,In_1483);
and U738 (N_738,In_103,In_1193);
nor U739 (N_739,In_958,In_1305);
and U740 (N_740,In_307,In_845);
nand U741 (N_741,In_207,In_1087);
and U742 (N_742,In_939,In_263);
and U743 (N_743,In_1141,In_396);
nor U744 (N_744,In_1187,In_214);
or U745 (N_745,In_1102,In_895);
and U746 (N_746,In_73,In_49);
nor U747 (N_747,In_95,In_790);
nand U748 (N_748,In_15,In_917);
nand U749 (N_749,In_1316,In_1406);
and U750 (N_750,In_256,In_1381);
and U751 (N_751,In_1229,In_1);
nand U752 (N_752,In_745,In_410);
nor U753 (N_753,In_966,In_633);
or U754 (N_754,In_1174,In_254);
and U755 (N_755,In_609,In_720);
nor U756 (N_756,In_1447,In_965);
and U757 (N_757,In_1493,In_107);
nor U758 (N_758,In_400,In_1308);
nand U759 (N_759,In_447,In_1321);
or U760 (N_760,In_611,In_151);
or U761 (N_761,In_140,In_745);
or U762 (N_762,In_322,In_870);
and U763 (N_763,In_892,In_1077);
xnor U764 (N_764,In_269,In_500);
nor U765 (N_765,In_246,In_470);
nor U766 (N_766,In_1499,In_926);
and U767 (N_767,In_361,In_527);
nand U768 (N_768,In_576,In_341);
nor U769 (N_769,In_348,In_527);
nand U770 (N_770,In_1143,In_1338);
or U771 (N_771,In_1362,In_319);
nand U772 (N_772,In_808,In_689);
nand U773 (N_773,In_48,In_308);
or U774 (N_774,In_89,In_1317);
and U775 (N_775,In_814,In_464);
or U776 (N_776,In_913,In_957);
xnor U777 (N_777,In_361,In_857);
or U778 (N_778,In_254,In_122);
and U779 (N_779,In_1212,In_532);
nor U780 (N_780,In_970,In_1122);
nand U781 (N_781,In_561,In_1006);
nand U782 (N_782,In_1153,In_651);
or U783 (N_783,In_240,In_1);
nand U784 (N_784,In_1427,In_45);
and U785 (N_785,In_500,In_726);
and U786 (N_786,In_211,In_364);
or U787 (N_787,In_1084,In_1420);
nor U788 (N_788,In_1425,In_528);
nor U789 (N_789,In_1494,In_827);
nor U790 (N_790,In_596,In_1152);
nor U791 (N_791,In_869,In_359);
or U792 (N_792,In_1001,In_918);
nor U793 (N_793,In_1371,In_914);
or U794 (N_794,In_1025,In_219);
or U795 (N_795,In_239,In_1208);
and U796 (N_796,In_3,In_694);
or U797 (N_797,In_1168,In_724);
or U798 (N_798,In_202,In_783);
nand U799 (N_799,In_1414,In_1078);
or U800 (N_800,In_609,In_712);
or U801 (N_801,In_100,In_700);
or U802 (N_802,In_321,In_1382);
nand U803 (N_803,In_1054,In_1467);
and U804 (N_804,In_351,In_733);
or U805 (N_805,In_41,In_1100);
and U806 (N_806,In_879,In_336);
and U807 (N_807,In_323,In_1415);
nand U808 (N_808,In_80,In_503);
nor U809 (N_809,In_211,In_622);
nor U810 (N_810,In_1032,In_1360);
or U811 (N_811,In_1362,In_782);
and U812 (N_812,In_3,In_984);
and U813 (N_813,In_1189,In_356);
and U814 (N_814,In_1412,In_1076);
or U815 (N_815,In_751,In_623);
nand U816 (N_816,In_148,In_343);
nand U817 (N_817,In_105,In_599);
or U818 (N_818,In_1082,In_542);
and U819 (N_819,In_628,In_805);
and U820 (N_820,In_1039,In_935);
and U821 (N_821,In_582,In_1102);
and U822 (N_822,In_916,In_211);
and U823 (N_823,In_654,In_190);
or U824 (N_824,In_525,In_1213);
and U825 (N_825,In_1417,In_1100);
or U826 (N_826,In_676,In_1245);
and U827 (N_827,In_137,In_699);
xnor U828 (N_828,In_274,In_839);
nor U829 (N_829,In_1059,In_761);
or U830 (N_830,In_1494,In_1457);
or U831 (N_831,In_26,In_313);
and U832 (N_832,In_728,In_979);
and U833 (N_833,In_1020,In_443);
and U834 (N_834,In_23,In_1316);
nand U835 (N_835,In_1259,In_481);
nand U836 (N_836,In_861,In_1410);
nor U837 (N_837,In_37,In_318);
or U838 (N_838,In_396,In_716);
or U839 (N_839,In_1052,In_1147);
and U840 (N_840,In_1210,In_442);
nor U841 (N_841,In_25,In_306);
nor U842 (N_842,In_381,In_200);
nor U843 (N_843,In_937,In_867);
nand U844 (N_844,In_76,In_177);
and U845 (N_845,In_1203,In_1089);
nand U846 (N_846,In_16,In_514);
or U847 (N_847,In_1330,In_450);
nand U848 (N_848,In_1393,In_967);
nand U849 (N_849,In_907,In_637);
and U850 (N_850,In_706,In_1298);
or U851 (N_851,In_184,In_1223);
and U852 (N_852,In_402,In_144);
nand U853 (N_853,In_725,In_821);
or U854 (N_854,In_1490,In_884);
and U855 (N_855,In_655,In_159);
nor U856 (N_856,In_1126,In_401);
and U857 (N_857,In_1039,In_257);
and U858 (N_858,In_1497,In_163);
nand U859 (N_859,In_1487,In_517);
nor U860 (N_860,In_1219,In_1284);
or U861 (N_861,In_1232,In_334);
nand U862 (N_862,In_834,In_198);
nor U863 (N_863,In_1397,In_1432);
nor U864 (N_864,In_367,In_717);
nand U865 (N_865,In_768,In_1260);
nand U866 (N_866,In_1047,In_983);
nor U867 (N_867,In_1466,In_1488);
and U868 (N_868,In_817,In_272);
nor U869 (N_869,In_169,In_455);
or U870 (N_870,In_724,In_103);
and U871 (N_871,In_1058,In_1296);
nor U872 (N_872,In_329,In_199);
nand U873 (N_873,In_1216,In_592);
and U874 (N_874,In_243,In_1493);
nand U875 (N_875,In_1228,In_758);
or U876 (N_876,In_939,In_858);
or U877 (N_877,In_495,In_1453);
or U878 (N_878,In_1083,In_1189);
and U879 (N_879,In_1232,In_654);
nand U880 (N_880,In_980,In_671);
or U881 (N_881,In_397,In_1383);
nand U882 (N_882,In_1283,In_1134);
nand U883 (N_883,In_172,In_1071);
and U884 (N_884,In_1378,In_547);
nand U885 (N_885,In_87,In_757);
and U886 (N_886,In_289,In_1294);
nand U887 (N_887,In_424,In_1328);
nand U888 (N_888,In_906,In_881);
nor U889 (N_889,In_1226,In_837);
nand U890 (N_890,In_97,In_177);
or U891 (N_891,In_765,In_1080);
and U892 (N_892,In_151,In_210);
or U893 (N_893,In_1096,In_268);
or U894 (N_894,In_708,In_434);
and U895 (N_895,In_171,In_1349);
xnor U896 (N_896,In_154,In_195);
and U897 (N_897,In_367,In_255);
xnor U898 (N_898,In_1395,In_900);
nor U899 (N_899,In_1230,In_1244);
nand U900 (N_900,In_1497,In_664);
and U901 (N_901,In_390,In_1423);
and U902 (N_902,In_386,In_205);
and U903 (N_903,In_4,In_1243);
nand U904 (N_904,In_302,In_1310);
or U905 (N_905,In_1287,In_87);
and U906 (N_906,In_1412,In_302);
nand U907 (N_907,In_504,In_1309);
nand U908 (N_908,In_1150,In_92);
nand U909 (N_909,In_151,In_982);
and U910 (N_910,In_1138,In_1096);
nor U911 (N_911,In_347,In_267);
nand U912 (N_912,In_32,In_124);
nand U913 (N_913,In_1218,In_675);
or U914 (N_914,In_382,In_952);
nand U915 (N_915,In_1455,In_96);
nand U916 (N_916,In_1344,In_923);
and U917 (N_917,In_1016,In_563);
nand U918 (N_918,In_19,In_472);
nand U919 (N_919,In_1418,In_700);
or U920 (N_920,In_412,In_88);
or U921 (N_921,In_445,In_909);
or U922 (N_922,In_1238,In_75);
and U923 (N_923,In_981,In_1390);
nand U924 (N_924,In_146,In_632);
nor U925 (N_925,In_414,In_1393);
and U926 (N_926,In_1072,In_395);
nand U927 (N_927,In_722,In_65);
and U928 (N_928,In_1340,In_107);
nand U929 (N_929,In_1258,In_585);
or U930 (N_930,In_118,In_6);
nand U931 (N_931,In_1294,In_618);
nand U932 (N_932,In_158,In_303);
nor U933 (N_933,In_830,In_3);
and U934 (N_934,In_1478,In_1424);
and U935 (N_935,In_1338,In_1253);
nand U936 (N_936,In_229,In_720);
and U937 (N_937,In_448,In_1330);
and U938 (N_938,In_1438,In_199);
or U939 (N_939,In_48,In_422);
and U940 (N_940,In_1079,In_642);
or U941 (N_941,In_69,In_68);
nand U942 (N_942,In_809,In_415);
nand U943 (N_943,In_587,In_557);
and U944 (N_944,In_1325,In_901);
nand U945 (N_945,In_186,In_999);
nand U946 (N_946,In_433,In_672);
nand U947 (N_947,In_1418,In_968);
or U948 (N_948,In_19,In_1423);
or U949 (N_949,In_1296,In_478);
and U950 (N_950,In_381,In_789);
or U951 (N_951,In_125,In_1153);
nor U952 (N_952,In_1268,In_734);
and U953 (N_953,In_1086,In_267);
nor U954 (N_954,In_34,In_173);
and U955 (N_955,In_905,In_471);
nand U956 (N_956,In_658,In_766);
nand U957 (N_957,In_1157,In_626);
or U958 (N_958,In_16,In_628);
nor U959 (N_959,In_601,In_302);
nand U960 (N_960,In_77,In_1187);
nand U961 (N_961,In_385,In_1237);
nor U962 (N_962,In_838,In_186);
nand U963 (N_963,In_548,In_571);
and U964 (N_964,In_1305,In_1420);
and U965 (N_965,In_1218,In_911);
or U966 (N_966,In_333,In_1165);
nor U967 (N_967,In_1023,In_1494);
nand U968 (N_968,In_432,In_1495);
or U969 (N_969,In_789,In_865);
and U970 (N_970,In_388,In_288);
and U971 (N_971,In_291,In_881);
and U972 (N_972,In_1197,In_30);
and U973 (N_973,In_525,In_407);
nor U974 (N_974,In_152,In_618);
and U975 (N_975,In_72,In_124);
or U976 (N_976,In_1321,In_379);
or U977 (N_977,In_740,In_1490);
nor U978 (N_978,In_90,In_607);
and U979 (N_979,In_944,In_1239);
nand U980 (N_980,In_1077,In_495);
nor U981 (N_981,In_333,In_888);
and U982 (N_982,In_736,In_838);
nand U983 (N_983,In_1400,In_152);
nand U984 (N_984,In_494,In_1467);
nor U985 (N_985,In_100,In_619);
or U986 (N_986,In_279,In_545);
or U987 (N_987,In_481,In_484);
nor U988 (N_988,In_1461,In_322);
nor U989 (N_989,In_317,In_800);
or U990 (N_990,In_1034,In_575);
nor U991 (N_991,In_1068,In_298);
and U992 (N_992,In_1486,In_119);
nor U993 (N_993,In_593,In_9);
nor U994 (N_994,In_418,In_733);
or U995 (N_995,In_1423,In_604);
or U996 (N_996,In_408,In_970);
nand U997 (N_997,In_854,In_849);
and U998 (N_998,In_1157,In_472);
or U999 (N_999,In_1238,In_1459);
or U1000 (N_1000,N_522,N_19);
nor U1001 (N_1001,N_952,N_274);
nand U1002 (N_1002,N_345,N_407);
and U1003 (N_1003,N_653,N_256);
or U1004 (N_1004,N_387,N_752);
nand U1005 (N_1005,N_654,N_13);
and U1006 (N_1006,N_816,N_415);
or U1007 (N_1007,N_369,N_129);
nor U1008 (N_1008,N_556,N_83);
nor U1009 (N_1009,N_690,N_416);
nor U1010 (N_1010,N_174,N_319);
or U1011 (N_1011,N_218,N_803);
nand U1012 (N_1012,N_789,N_772);
nor U1013 (N_1013,N_549,N_409);
and U1014 (N_1014,N_465,N_646);
and U1015 (N_1015,N_989,N_843);
nor U1016 (N_1016,N_400,N_657);
and U1017 (N_1017,N_623,N_460);
nor U1018 (N_1018,N_920,N_329);
nand U1019 (N_1019,N_420,N_141);
or U1020 (N_1020,N_406,N_722);
nand U1021 (N_1021,N_709,N_333);
or U1022 (N_1022,N_750,N_717);
and U1023 (N_1023,N_837,N_892);
nand U1024 (N_1024,N_393,N_919);
nor U1025 (N_1025,N_733,N_317);
or U1026 (N_1026,N_427,N_23);
and U1027 (N_1027,N_894,N_878);
and U1028 (N_1028,N_270,N_248);
nand U1029 (N_1029,N_821,N_375);
nor U1030 (N_1030,N_234,N_70);
nand U1031 (N_1031,N_448,N_518);
nand U1032 (N_1032,N_631,N_910);
or U1033 (N_1033,N_179,N_859);
or U1034 (N_1034,N_966,N_201);
nor U1035 (N_1035,N_55,N_413);
or U1036 (N_1036,N_957,N_691);
or U1037 (N_1037,N_969,N_689);
nand U1038 (N_1038,N_147,N_804);
and U1039 (N_1039,N_634,N_109);
and U1040 (N_1040,N_80,N_169);
nand U1041 (N_1041,N_240,N_492);
or U1042 (N_1042,N_110,N_66);
nand U1043 (N_1043,N_189,N_408);
or U1044 (N_1044,N_869,N_73);
nand U1045 (N_1045,N_142,N_106);
nor U1046 (N_1046,N_14,N_753);
and U1047 (N_1047,N_363,N_69);
or U1048 (N_1048,N_632,N_578);
nor U1049 (N_1049,N_356,N_462);
or U1050 (N_1050,N_799,N_216);
and U1051 (N_1051,N_974,N_111);
nand U1052 (N_1052,N_638,N_257);
or U1053 (N_1053,N_673,N_222);
nor U1054 (N_1054,N_644,N_190);
nand U1055 (N_1055,N_504,N_575);
nor U1056 (N_1056,N_891,N_770);
nand U1057 (N_1057,N_811,N_525);
or U1058 (N_1058,N_202,N_585);
nor U1059 (N_1059,N_516,N_624);
nand U1060 (N_1060,N_75,N_498);
and U1061 (N_1061,N_939,N_477);
nand U1062 (N_1062,N_215,N_207);
nor U1063 (N_1063,N_718,N_641);
nand U1064 (N_1064,N_760,N_315);
or U1065 (N_1065,N_383,N_814);
nand U1066 (N_1066,N_245,N_568);
xor U1067 (N_1067,N_873,N_530);
and U1068 (N_1068,N_74,N_990);
nand U1069 (N_1069,N_545,N_376);
nor U1070 (N_1070,N_531,N_22);
nor U1071 (N_1071,N_62,N_312);
nand U1072 (N_1072,N_739,N_671);
or U1073 (N_1073,N_343,N_721);
and U1074 (N_1074,N_981,N_125);
or U1075 (N_1075,N_502,N_64);
nor U1076 (N_1076,N_3,N_205);
nand U1077 (N_1077,N_355,N_359);
or U1078 (N_1078,N_922,N_338);
or U1079 (N_1079,N_337,N_130);
nor U1080 (N_1080,N_506,N_225);
and U1081 (N_1081,N_322,N_209);
and U1082 (N_1082,N_851,N_149);
nor U1083 (N_1083,N_128,N_742);
and U1084 (N_1084,N_609,N_49);
or U1085 (N_1085,N_622,N_348);
and U1086 (N_1086,N_982,N_326);
nand U1087 (N_1087,N_566,N_610);
or U1088 (N_1088,N_135,N_703);
or U1089 (N_1089,N_378,N_801);
and U1090 (N_1090,N_834,N_439);
or U1091 (N_1091,N_674,N_719);
and U1092 (N_1092,N_454,N_954);
and U1093 (N_1093,N_987,N_764);
and U1094 (N_1094,N_133,N_787);
nand U1095 (N_1095,N_395,N_830);
nand U1096 (N_1096,N_479,N_542);
nor U1097 (N_1097,N_441,N_445);
nand U1098 (N_1098,N_267,N_9);
or U1099 (N_1099,N_808,N_436);
and U1100 (N_1100,N_157,N_853);
and U1101 (N_1101,N_204,N_486);
and U1102 (N_1102,N_452,N_405);
and U1103 (N_1103,N_567,N_991);
and U1104 (N_1104,N_451,N_613);
and U1105 (N_1105,N_725,N_265);
nand U1106 (N_1106,N_951,N_306);
or U1107 (N_1107,N_354,N_501);
nand U1108 (N_1108,N_669,N_698);
or U1109 (N_1109,N_18,N_927);
nor U1110 (N_1110,N_170,N_724);
nand U1111 (N_1111,N_94,N_795);
or U1112 (N_1112,N_391,N_438);
nand U1113 (N_1113,N_261,N_797);
nand U1114 (N_1114,N_767,N_140);
nand U1115 (N_1115,N_880,N_308);
nor U1116 (N_1116,N_537,N_586);
or U1117 (N_1117,N_194,N_377);
or U1118 (N_1118,N_561,N_636);
nor U1119 (N_1119,N_771,N_175);
or U1120 (N_1120,N_842,N_574);
and U1121 (N_1121,N_960,N_883);
or U1122 (N_1122,N_693,N_446);
nor U1123 (N_1123,N_361,N_802);
and U1124 (N_1124,N_250,N_12);
or U1125 (N_1125,N_788,N_302);
nand U1126 (N_1126,N_382,N_292);
nor U1127 (N_1127,N_854,N_323);
nand U1128 (N_1128,N_404,N_972);
and U1129 (N_1129,N_325,N_307);
or U1130 (N_1130,N_874,N_210);
and U1131 (N_1131,N_65,N_628);
nand U1132 (N_1132,N_605,N_291);
nor U1133 (N_1133,N_173,N_737);
and U1134 (N_1134,N_857,N_365);
and U1135 (N_1135,N_785,N_212);
nand U1136 (N_1136,N_992,N_712);
or U1137 (N_1137,N_903,N_339);
and U1138 (N_1138,N_444,N_702);
and U1139 (N_1139,N_871,N_579);
nand U1140 (N_1140,N_480,N_794);
and U1141 (N_1141,N_658,N_984);
or U1142 (N_1142,N_134,N_371);
and U1143 (N_1143,N_493,N_227);
and U1144 (N_1144,N_941,N_429);
and U1145 (N_1145,N_652,N_963);
and U1146 (N_1146,N_964,N_380);
and U1147 (N_1147,N_311,N_113);
and U1148 (N_1148,N_226,N_589);
nor U1149 (N_1149,N_366,N_178);
nand U1150 (N_1150,N_560,N_114);
and U1151 (N_1151,N_651,N_546);
and U1152 (N_1152,N_870,N_573);
nor U1153 (N_1153,N_850,N_699);
or U1154 (N_1154,N_642,N_845);
nand U1155 (N_1155,N_98,N_805);
or U1156 (N_1156,N_105,N_81);
or U1157 (N_1157,N_148,N_357);
and U1158 (N_1158,N_995,N_91);
nand U1159 (N_1159,N_158,N_900);
or U1160 (N_1160,N_707,N_513);
nand U1161 (N_1161,N_591,N_428);
nand U1162 (N_1162,N_661,N_188);
and U1163 (N_1163,N_39,N_904);
nor U1164 (N_1164,N_595,N_253);
or U1165 (N_1165,N_385,N_145);
or U1166 (N_1166,N_353,N_263);
nor U1167 (N_1167,N_694,N_24);
nor U1168 (N_1168,N_977,N_784);
and U1169 (N_1169,N_675,N_21);
nor U1170 (N_1170,N_97,N_344);
and U1171 (N_1171,N_119,N_136);
nor U1172 (N_1172,N_536,N_911);
nand U1173 (N_1173,N_303,N_800);
and U1174 (N_1174,N_425,N_749);
or U1175 (N_1175,N_120,N_971);
and U1176 (N_1176,N_381,N_162);
xnor U1177 (N_1177,N_934,N_602);
and U1178 (N_1178,N_379,N_523);
or U1179 (N_1179,N_997,N_540);
nand U1180 (N_1180,N_104,N_96);
and U1181 (N_1181,N_818,N_424);
nor U1182 (N_1182,N_347,N_738);
and U1183 (N_1183,N_47,N_773);
or U1184 (N_1184,N_825,N_778);
or U1185 (N_1185,N_713,N_432);
or U1186 (N_1186,N_763,N_336);
or U1187 (N_1187,N_596,N_466);
and U1188 (N_1188,N_633,N_953);
nor U1189 (N_1189,N_195,N_581);
xnor U1190 (N_1190,N_351,N_213);
xnor U1191 (N_1191,N_84,N_916);
and U1192 (N_1192,N_437,N_824);
or U1193 (N_1193,N_233,N_565);
or U1194 (N_1194,N_933,N_755);
nor U1195 (N_1195,N_876,N_450);
nor U1196 (N_1196,N_423,N_102);
or U1197 (N_1197,N_882,N_386);
or U1198 (N_1198,N_743,N_993);
and U1199 (N_1199,N_362,N_153);
nor U1200 (N_1200,N_676,N_937);
nor U1201 (N_1201,N_751,N_601);
nand U1202 (N_1202,N_67,N_590);
and U1203 (N_1203,N_647,N_171);
and U1204 (N_1204,N_289,N_364);
nor U1205 (N_1205,N_164,N_52);
nand U1206 (N_1206,N_115,N_181);
or U1207 (N_1207,N_761,N_470);
nand U1208 (N_1208,N_687,N_985);
nand U1209 (N_1209,N_783,N_898);
or U1210 (N_1210,N_28,N_714);
or U1211 (N_1211,N_766,N_544);
nand U1212 (N_1212,N_491,N_817);
or U1213 (N_1213,N_48,N_527);
nor U1214 (N_1214,N_123,N_53);
or U1215 (N_1215,N_31,N_731);
nor U1216 (N_1216,N_10,N_367);
and U1217 (N_1217,N_517,N_4);
nor U1218 (N_1218,N_241,N_686);
nand U1219 (N_1219,N_865,N_469);
nor U1220 (N_1220,N_283,N_33);
and U1221 (N_1221,N_756,N_812);
and U1222 (N_1222,N_695,N_666);
nand U1223 (N_1223,N_199,N_45);
or U1224 (N_1224,N_663,N_607);
and U1225 (N_1225,N_417,N_146);
nand U1226 (N_1226,N_776,N_252);
or U1227 (N_1227,N_603,N_598);
nor U1228 (N_1228,N_433,N_979);
and U1229 (N_1229,N_942,N_862);
nor U1230 (N_1230,N_27,N_852);
nor U1231 (N_1231,N_580,N_790);
nor U1232 (N_1232,N_294,N_823);
and U1233 (N_1233,N_727,N_988);
and U1234 (N_1234,N_889,N_112);
nand U1235 (N_1235,N_976,N_374);
and U1236 (N_1236,N_877,N_372);
or U1237 (N_1237,N_606,N_144);
or U1238 (N_1238,N_269,N_685);
and U1239 (N_1239,N_290,N_217);
nand U1240 (N_1240,N_7,N_127);
nor U1241 (N_1241,N_532,N_464);
or U1242 (N_1242,N_100,N_664);
or U1243 (N_1243,N_583,N_863);
nand U1244 (N_1244,N_151,N_611);
or U1245 (N_1245,N_680,N_320);
and U1246 (N_1246,N_926,N_193);
or U1247 (N_1247,N_279,N_499);
nor U1248 (N_1248,N_107,N_422);
nor U1249 (N_1249,N_534,N_798);
nor U1250 (N_1250,N_983,N_500);
or U1251 (N_1251,N_822,N_980);
or U1252 (N_1252,N_288,N_901);
nor U1253 (N_1253,N_779,N_887);
or U1254 (N_1254,N_342,N_529);
and U1255 (N_1255,N_392,N_572);
nor U1256 (N_1256,N_793,N_897);
nor U1257 (N_1257,N_678,N_293);
and U1258 (N_1258,N_961,N_397);
nor U1259 (N_1259,N_160,N_597);
or U1260 (N_1260,N_832,N_5);
nor U1261 (N_1261,N_704,N_736);
nand U1262 (N_1262,N_187,N_373);
and U1263 (N_1263,N_57,N_1);
and U1264 (N_1264,N_543,N_166);
nor U1265 (N_1265,N_72,N_68);
or U1266 (N_1266,N_616,N_440);
and U1267 (N_1267,N_103,N_520);
nand U1268 (N_1268,N_935,N_316);
and U1269 (N_1269,N_280,N_389);
nor U1270 (N_1270,N_515,N_621);
or U1271 (N_1271,N_947,N_258);
nor U1272 (N_1272,N_528,N_973);
nand U1273 (N_1273,N_305,N_820);
nand U1274 (N_1274,N_411,N_124);
and U1275 (N_1275,N_16,N_998);
and U1276 (N_1276,N_925,N_899);
nand U1277 (N_1277,N_324,N_907);
or U1278 (N_1278,N_748,N_708);
and U1279 (N_1279,N_924,N_792);
nor U1280 (N_1280,N_472,N_914);
nand U1281 (N_1281,N_197,N_978);
and U1282 (N_1282,N_370,N_402);
and U1283 (N_1283,N_640,N_885);
nor U1284 (N_1284,N_774,N_399);
nor U1285 (N_1285,N_677,N_893);
nor U1286 (N_1286,N_78,N_777);
nand U1287 (N_1287,N_414,N_223);
nor U1288 (N_1288,N_615,N_861);
nand U1289 (N_1289,N_909,N_273);
and U1290 (N_1290,N_667,N_943);
nor U1291 (N_1291,N_255,N_150);
nor U1292 (N_1292,N_155,N_740);
or U1293 (N_1293,N_582,N_758);
nor U1294 (N_1294,N_512,N_884);
nor U1295 (N_1295,N_327,N_447);
and U1296 (N_1296,N_994,N_430);
and U1297 (N_1297,N_86,N_349);
and U1298 (N_1298,N_34,N_459);
or U1299 (N_1299,N_254,N_36);
nor U1300 (N_1300,N_314,N_945);
nor U1301 (N_1301,N_913,N_99);
nand U1302 (N_1302,N_970,N_905);
and U1303 (N_1303,N_815,N_260);
nor U1304 (N_1304,N_786,N_849);
nor U1305 (N_1305,N_118,N_236);
nor U1306 (N_1306,N_547,N_32);
nand U1307 (N_1307,N_827,N_569);
nor U1308 (N_1308,N_716,N_745);
nor U1309 (N_1309,N_619,N_15);
or U1310 (N_1310,N_780,N_683);
and U1311 (N_1311,N_56,N_95);
and U1312 (N_1312,N_809,N_592);
and U1313 (N_1313,N_59,N_643);
or U1314 (N_1314,N_620,N_588);
and U1315 (N_1315,N_167,N_259);
and U1316 (N_1316,N_866,N_744);
nor U1317 (N_1317,N_846,N_43);
or U1318 (N_1318,N_313,N_475);
nor U1319 (N_1319,N_231,N_192);
or U1320 (N_1320,N_154,N_284);
and U1321 (N_1321,N_38,N_929);
or U1322 (N_1322,N_757,N_729);
or U1323 (N_1323,N_810,N_426);
or U1324 (N_1324,N_285,N_741);
nand U1325 (N_1325,N_828,N_180);
xor U1326 (N_1326,N_948,N_476);
and U1327 (N_1327,N_20,N_858);
nor U1328 (N_1328,N_833,N_487);
nand U1329 (N_1329,N_419,N_630);
nor U1330 (N_1330,N_548,N_266);
or U1331 (N_1331,N_775,N_458);
and U1332 (N_1332,N_50,N_421);
and U1333 (N_1333,N_541,N_54);
nand U1334 (N_1334,N_473,N_896);
or U1335 (N_1335,N_101,N_461);
nand U1336 (N_1336,N_51,N_242);
and U1337 (N_1337,N_728,N_304);
or U1338 (N_1338,N_35,N_697);
nand U1339 (N_1339,N_198,N_635);
nand U1340 (N_1340,N_944,N_553);
nor U1341 (N_1341,N_172,N_844);
or U1342 (N_1342,N_701,N_552);
nor U1343 (N_1343,N_684,N_867);
and U1344 (N_1344,N_649,N_539);
nand U1345 (N_1345,N_625,N_868);
and U1346 (N_1346,N_309,N_453);
nor U1347 (N_1347,N_650,N_116);
and U1348 (N_1348,N_177,N_143);
nor U1349 (N_1349,N_886,N_88);
xnor U1350 (N_1350,N_396,N_272);
nand U1351 (N_1351,N_139,N_490);
nand U1352 (N_1352,N_496,N_29);
and U1353 (N_1353,N_996,N_191);
nor U1354 (N_1354,N_584,N_662);
nand U1355 (N_1355,N_835,N_235);
nand U1356 (N_1356,N_768,N_468);
nand U1357 (N_1357,N_659,N_89);
and U1358 (N_1358,N_958,N_999);
or U1359 (N_1359,N_617,N_554);
or U1360 (N_1360,N_482,N_237);
and U1361 (N_1361,N_390,N_403);
xnor U1362 (N_1362,N_829,N_77);
nand U1363 (N_1363,N_298,N_456);
nand U1364 (N_1364,N_836,N_246);
or U1365 (N_1365,N_219,N_864);
and U1366 (N_1366,N_965,N_940);
and U1367 (N_1367,N_831,N_819);
nand U1368 (N_1368,N_946,N_58);
and U1369 (N_1369,N_271,N_856);
or U1370 (N_1370,N_182,N_524);
xnor U1371 (N_1371,N_521,N_90);
nor U1372 (N_1372,N_847,N_350);
nor U1373 (N_1373,N_551,N_670);
and U1374 (N_1374,N_706,N_986);
nor U1375 (N_1375,N_950,N_495);
nand U1376 (N_1376,N_514,N_30);
nor U1377 (N_1377,N_715,N_519);
and U1378 (N_1378,N_875,N_25);
or U1379 (N_1379,N_478,N_214);
and U1380 (N_1380,N_507,N_185);
and U1381 (N_1381,N_902,N_137);
and U1382 (N_1382,N_681,N_6);
nand U1383 (N_1383,N_442,N_700);
or U1384 (N_1384,N_796,N_682);
and U1385 (N_1385,N_723,N_710);
nor U1386 (N_1386,N_484,N_296);
or U1387 (N_1387,N_557,N_76);
nand U1388 (N_1388,N_108,N_126);
or U1389 (N_1389,N_855,N_570);
nand U1390 (N_1390,N_908,N_17);
or U1391 (N_1391,N_156,N_921);
nand U1392 (N_1392,N_626,N_564);
nand U1393 (N_1393,N_872,N_769);
nand U1394 (N_1394,N_511,N_747);
and U1395 (N_1395,N_224,N_746);
or U1396 (N_1396,N_660,N_587);
or U1397 (N_1397,N_726,N_968);
nand U1398 (N_1398,N_759,N_232);
nor U1399 (N_1399,N_932,N_247);
or U1400 (N_1400,N_330,N_754);
or U1401 (N_1401,N_163,N_959);
or U1402 (N_1402,N_287,N_637);
or U1403 (N_1403,N_394,N_410);
nor U1404 (N_1404,N_938,N_268);
and U1405 (N_1405,N_443,N_879);
or U1406 (N_1406,N_765,N_494);
nor U1407 (N_1407,N_161,N_705);
nand U1408 (N_1408,N_211,N_956);
nor U1409 (N_1409,N_483,N_457);
nand U1410 (N_1410,N_618,N_138);
nor U1411 (N_1411,N_71,N_949);
and U1412 (N_1412,N_229,N_300);
and U1413 (N_1413,N_301,N_340);
or U1414 (N_1414,N_206,N_61);
or U1415 (N_1415,N_917,N_912);
or U1416 (N_1416,N_599,N_826);
or U1417 (N_1417,N_335,N_2);
nor U1418 (N_1418,N_895,N_558);
nand U1419 (N_1419,N_848,N_696);
nand U1420 (N_1420,N_645,N_0);
nor U1421 (N_1421,N_711,N_299);
xor U1422 (N_1422,N_533,N_807);
or U1423 (N_1423,N_967,N_559);
and U1424 (N_1424,N_510,N_321);
xor U1425 (N_1425,N_509,N_200);
or U1426 (N_1426,N_183,N_117);
and U1427 (N_1427,N_40,N_612);
or U1428 (N_1428,N_688,N_434);
nor U1429 (N_1429,N_318,N_276);
nand U1430 (N_1430,N_975,N_526);
nand U1431 (N_1431,N_282,N_593);
nand U1432 (N_1432,N_332,N_388);
or U1433 (N_1433,N_87,N_220);
and U1434 (N_1434,N_412,N_352);
nand U1435 (N_1435,N_485,N_608);
and U1436 (N_1436,N_648,N_131);
nand U1437 (N_1437,N_538,N_221);
nor U1438 (N_1438,N_503,N_79);
or U1439 (N_1439,N_358,N_281);
or U1440 (N_1440,N_840,N_435);
nand U1441 (N_1441,N_629,N_60);
or U1442 (N_1442,N_550,N_243);
nor U1443 (N_1443,N_576,N_46);
nor U1444 (N_1444,N_918,N_806);
nand U1445 (N_1445,N_44,N_735);
nor U1446 (N_1446,N_93,N_449);
or U1447 (N_1447,N_368,N_838);
nor U1448 (N_1448,N_122,N_562);
nand U1449 (N_1449,N_888,N_962);
or U1450 (N_1450,N_781,N_152);
nor U1451 (N_1451,N_535,N_655);
and U1452 (N_1452,N_228,N_594);
nor U1453 (N_1453,N_931,N_782);
nor U1454 (N_1454,N_791,N_604);
or U1455 (N_1455,N_614,N_762);
and U1456 (N_1456,N_627,N_839);
and U1457 (N_1457,N_11,N_813);
nor U1458 (N_1458,N_489,N_82);
and U1459 (N_1459,N_398,N_360);
and U1460 (N_1460,N_577,N_244);
nor U1461 (N_1461,N_600,N_238);
or U1462 (N_1462,N_732,N_656);
nand U1463 (N_1463,N_384,N_692);
or U1464 (N_1464,N_230,N_42);
nor U1465 (N_1465,N_168,N_63);
nand U1466 (N_1466,N_928,N_455);
or U1467 (N_1467,N_346,N_121);
nand U1468 (N_1468,N_331,N_334);
nand U1469 (N_1469,N_159,N_563);
or U1470 (N_1470,N_906,N_474);
nor U1471 (N_1471,N_471,N_41);
nand U1472 (N_1472,N_463,N_930);
nand U1473 (N_1473,N_890,N_505);
nand U1474 (N_1474,N_665,N_341);
and U1475 (N_1475,N_328,N_186);
nand U1476 (N_1476,N_860,N_555);
nor U1477 (N_1477,N_720,N_679);
xnor U1478 (N_1478,N_278,N_639);
or U1479 (N_1479,N_467,N_262);
or U1480 (N_1480,N_8,N_277);
nor U1481 (N_1481,N_668,N_92);
nor U1482 (N_1482,N_881,N_295);
nand U1483 (N_1483,N_26,N_165);
and U1484 (N_1484,N_297,N_730);
nand U1485 (N_1485,N_203,N_401);
nand U1486 (N_1486,N_85,N_915);
nand U1487 (N_1487,N_488,N_481);
nand U1488 (N_1488,N_431,N_571);
and U1489 (N_1489,N_310,N_418);
nor U1490 (N_1490,N_936,N_923);
or U1491 (N_1491,N_955,N_176);
nand U1492 (N_1492,N_249,N_841);
nor U1493 (N_1493,N_184,N_672);
or U1494 (N_1494,N_251,N_37);
nor U1495 (N_1495,N_239,N_264);
and U1496 (N_1496,N_208,N_734);
or U1497 (N_1497,N_497,N_286);
and U1498 (N_1498,N_196,N_132);
or U1499 (N_1499,N_275,N_508);
or U1500 (N_1500,N_375,N_831);
nand U1501 (N_1501,N_227,N_638);
nor U1502 (N_1502,N_468,N_315);
nor U1503 (N_1503,N_875,N_178);
nand U1504 (N_1504,N_815,N_12);
and U1505 (N_1505,N_273,N_202);
or U1506 (N_1506,N_724,N_453);
and U1507 (N_1507,N_136,N_110);
and U1508 (N_1508,N_741,N_966);
and U1509 (N_1509,N_766,N_258);
nand U1510 (N_1510,N_396,N_150);
nor U1511 (N_1511,N_148,N_176);
or U1512 (N_1512,N_591,N_605);
nand U1513 (N_1513,N_103,N_847);
and U1514 (N_1514,N_640,N_563);
nand U1515 (N_1515,N_758,N_190);
and U1516 (N_1516,N_270,N_503);
and U1517 (N_1517,N_337,N_877);
or U1518 (N_1518,N_981,N_24);
nand U1519 (N_1519,N_774,N_448);
nand U1520 (N_1520,N_48,N_296);
or U1521 (N_1521,N_290,N_128);
nand U1522 (N_1522,N_644,N_973);
nor U1523 (N_1523,N_68,N_162);
and U1524 (N_1524,N_99,N_517);
nor U1525 (N_1525,N_431,N_375);
and U1526 (N_1526,N_438,N_623);
nand U1527 (N_1527,N_861,N_631);
and U1528 (N_1528,N_166,N_686);
nor U1529 (N_1529,N_875,N_524);
nand U1530 (N_1530,N_249,N_402);
nor U1531 (N_1531,N_921,N_355);
and U1532 (N_1532,N_1,N_272);
nor U1533 (N_1533,N_880,N_556);
or U1534 (N_1534,N_845,N_428);
nand U1535 (N_1535,N_605,N_486);
xor U1536 (N_1536,N_541,N_124);
and U1537 (N_1537,N_821,N_568);
nor U1538 (N_1538,N_174,N_688);
nor U1539 (N_1539,N_200,N_752);
nor U1540 (N_1540,N_76,N_356);
nor U1541 (N_1541,N_533,N_765);
nor U1542 (N_1542,N_768,N_767);
or U1543 (N_1543,N_878,N_781);
and U1544 (N_1544,N_34,N_982);
or U1545 (N_1545,N_835,N_326);
nor U1546 (N_1546,N_415,N_981);
and U1547 (N_1547,N_316,N_722);
nand U1548 (N_1548,N_824,N_491);
nor U1549 (N_1549,N_418,N_885);
and U1550 (N_1550,N_907,N_157);
and U1551 (N_1551,N_66,N_766);
nor U1552 (N_1552,N_429,N_14);
nand U1553 (N_1553,N_472,N_147);
nor U1554 (N_1554,N_856,N_12);
and U1555 (N_1555,N_61,N_53);
nor U1556 (N_1556,N_960,N_256);
nor U1557 (N_1557,N_557,N_327);
nor U1558 (N_1558,N_349,N_418);
nand U1559 (N_1559,N_120,N_57);
or U1560 (N_1560,N_67,N_517);
nor U1561 (N_1561,N_98,N_687);
or U1562 (N_1562,N_139,N_804);
nand U1563 (N_1563,N_72,N_515);
nor U1564 (N_1564,N_688,N_10);
or U1565 (N_1565,N_521,N_928);
nor U1566 (N_1566,N_583,N_40);
or U1567 (N_1567,N_673,N_26);
and U1568 (N_1568,N_211,N_2);
nand U1569 (N_1569,N_325,N_669);
nor U1570 (N_1570,N_15,N_544);
and U1571 (N_1571,N_166,N_338);
and U1572 (N_1572,N_521,N_870);
nand U1573 (N_1573,N_240,N_961);
nor U1574 (N_1574,N_716,N_117);
xor U1575 (N_1575,N_152,N_173);
nand U1576 (N_1576,N_872,N_698);
and U1577 (N_1577,N_136,N_288);
nor U1578 (N_1578,N_584,N_471);
and U1579 (N_1579,N_600,N_539);
nand U1580 (N_1580,N_228,N_888);
nor U1581 (N_1581,N_133,N_436);
or U1582 (N_1582,N_78,N_786);
nor U1583 (N_1583,N_144,N_225);
nand U1584 (N_1584,N_418,N_685);
or U1585 (N_1585,N_49,N_668);
nor U1586 (N_1586,N_401,N_840);
and U1587 (N_1587,N_733,N_234);
and U1588 (N_1588,N_136,N_230);
or U1589 (N_1589,N_125,N_801);
and U1590 (N_1590,N_815,N_83);
and U1591 (N_1591,N_162,N_673);
nor U1592 (N_1592,N_126,N_522);
and U1593 (N_1593,N_839,N_608);
and U1594 (N_1594,N_265,N_404);
nor U1595 (N_1595,N_897,N_254);
or U1596 (N_1596,N_128,N_504);
or U1597 (N_1597,N_420,N_276);
or U1598 (N_1598,N_761,N_23);
nand U1599 (N_1599,N_512,N_88);
or U1600 (N_1600,N_766,N_822);
or U1601 (N_1601,N_503,N_676);
nor U1602 (N_1602,N_155,N_153);
nor U1603 (N_1603,N_726,N_872);
nand U1604 (N_1604,N_462,N_617);
nand U1605 (N_1605,N_746,N_661);
nand U1606 (N_1606,N_413,N_100);
and U1607 (N_1607,N_342,N_792);
or U1608 (N_1608,N_275,N_35);
or U1609 (N_1609,N_897,N_49);
and U1610 (N_1610,N_774,N_723);
nor U1611 (N_1611,N_784,N_195);
nand U1612 (N_1612,N_249,N_243);
and U1613 (N_1613,N_243,N_207);
nand U1614 (N_1614,N_25,N_448);
and U1615 (N_1615,N_415,N_134);
and U1616 (N_1616,N_871,N_872);
and U1617 (N_1617,N_531,N_960);
nor U1618 (N_1618,N_88,N_697);
nand U1619 (N_1619,N_254,N_946);
nor U1620 (N_1620,N_66,N_197);
or U1621 (N_1621,N_951,N_709);
and U1622 (N_1622,N_709,N_754);
xor U1623 (N_1623,N_716,N_438);
or U1624 (N_1624,N_596,N_272);
nand U1625 (N_1625,N_712,N_140);
nand U1626 (N_1626,N_87,N_171);
nand U1627 (N_1627,N_322,N_733);
nor U1628 (N_1628,N_714,N_493);
or U1629 (N_1629,N_228,N_190);
nor U1630 (N_1630,N_936,N_974);
nand U1631 (N_1631,N_489,N_325);
nand U1632 (N_1632,N_393,N_377);
and U1633 (N_1633,N_603,N_523);
or U1634 (N_1634,N_673,N_671);
nor U1635 (N_1635,N_13,N_341);
and U1636 (N_1636,N_196,N_165);
and U1637 (N_1637,N_593,N_932);
or U1638 (N_1638,N_714,N_69);
and U1639 (N_1639,N_728,N_370);
nand U1640 (N_1640,N_260,N_942);
nor U1641 (N_1641,N_491,N_686);
or U1642 (N_1642,N_445,N_564);
nand U1643 (N_1643,N_612,N_260);
nand U1644 (N_1644,N_170,N_761);
nor U1645 (N_1645,N_469,N_622);
or U1646 (N_1646,N_571,N_253);
or U1647 (N_1647,N_975,N_342);
nor U1648 (N_1648,N_721,N_403);
or U1649 (N_1649,N_956,N_562);
or U1650 (N_1650,N_623,N_909);
nand U1651 (N_1651,N_13,N_460);
or U1652 (N_1652,N_942,N_656);
and U1653 (N_1653,N_951,N_662);
nor U1654 (N_1654,N_133,N_736);
or U1655 (N_1655,N_949,N_364);
nor U1656 (N_1656,N_94,N_421);
nand U1657 (N_1657,N_556,N_158);
nand U1658 (N_1658,N_385,N_486);
and U1659 (N_1659,N_100,N_772);
and U1660 (N_1660,N_71,N_794);
or U1661 (N_1661,N_784,N_843);
nor U1662 (N_1662,N_212,N_293);
or U1663 (N_1663,N_239,N_53);
nand U1664 (N_1664,N_202,N_869);
nor U1665 (N_1665,N_987,N_884);
or U1666 (N_1666,N_424,N_328);
nand U1667 (N_1667,N_526,N_212);
nand U1668 (N_1668,N_804,N_639);
nand U1669 (N_1669,N_206,N_143);
nand U1670 (N_1670,N_544,N_330);
and U1671 (N_1671,N_613,N_305);
and U1672 (N_1672,N_245,N_211);
and U1673 (N_1673,N_173,N_892);
nand U1674 (N_1674,N_159,N_264);
nand U1675 (N_1675,N_572,N_102);
nor U1676 (N_1676,N_364,N_287);
or U1677 (N_1677,N_137,N_866);
and U1678 (N_1678,N_896,N_797);
nor U1679 (N_1679,N_720,N_508);
nand U1680 (N_1680,N_630,N_37);
nor U1681 (N_1681,N_947,N_196);
nor U1682 (N_1682,N_727,N_318);
nand U1683 (N_1683,N_892,N_4);
and U1684 (N_1684,N_777,N_731);
or U1685 (N_1685,N_526,N_610);
nand U1686 (N_1686,N_452,N_14);
nand U1687 (N_1687,N_580,N_399);
and U1688 (N_1688,N_39,N_699);
and U1689 (N_1689,N_117,N_710);
nor U1690 (N_1690,N_626,N_978);
nand U1691 (N_1691,N_680,N_39);
nor U1692 (N_1692,N_958,N_772);
and U1693 (N_1693,N_340,N_944);
nand U1694 (N_1694,N_27,N_118);
or U1695 (N_1695,N_476,N_199);
xnor U1696 (N_1696,N_988,N_888);
nor U1697 (N_1697,N_689,N_23);
nand U1698 (N_1698,N_288,N_735);
nor U1699 (N_1699,N_346,N_677);
nand U1700 (N_1700,N_295,N_934);
and U1701 (N_1701,N_405,N_847);
or U1702 (N_1702,N_586,N_184);
and U1703 (N_1703,N_295,N_87);
nor U1704 (N_1704,N_678,N_769);
nand U1705 (N_1705,N_501,N_293);
or U1706 (N_1706,N_407,N_312);
or U1707 (N_1707,N_257,N_590);
nand U1708 (N_1708,N_195,N_804);
nand U1709 (N_1709,N_44,N_779);
or U1710 (N_1710,N_653,N_439);
or U1711 (N_1711,N_294,N_310);
and U1712 (N_1712,N_593,N_952);
nor U1713 (N_1713,N_971,N_334);
nor U1714 (N_1714,N_298,N_834);
nand U1715 (N_1715,N_998,N_402);
or U1716 (N_1716,N_940,N_772);
or U1717 (N_1717,N_97,N_294);
or U1718 (N_1718,N_170,N_28);
nor U1719 (N_1719,N_295,N_180);
and U1720 (N_1720,N_796,N_460);
nand U1721 (N_1721,N_924,N_379);
nor U1722 (N_1722,N_525,N_487);
or U1723 (N_1723,N_80,N_274);
or U1724 (N_1724,N_826,N_728);
nor U1725 (N_1725,N_621,N_466);
or U1726 (N_1726,N_896,N_520);
and U1727 (N_1727,N_325,N_404);
and U1728 (N_1728,N_906,N_874);
nor U1729 (N_1729,N_39,N_632);
nand U1730 (N_1730,N_837,N_288);
nor U1731 (N_1731,N_347,N_931);
nor U1732 (N_1732,N_928,N_313);
nand U1733 (N_1733,N_420,N_968);
or U1734 (N_1734,N_337,N_910);
or U1735 (N_1735,N_616,N_466);
nor U1736 (N_1736,N_476,N_991);
nor U1737 (N_1737,N_605,N_169);
nand U1738 (N_1738,N_247,N_157);
nand U1739 (N_1739,N_797,N_530);
nor U1740 (N_1740,N_405,N_241);
and U1741 (N_1741,N_542,N_283);
nand U1742 (N_1742,N_816,N_169);
or U1743 (N_1743,N_513,N_326);
and U1744 (N_1744,N_606,N_151);
and U1745 (N_1745,N_680,N_817);
or U1746 (N_1746,N_680,N_344);
and U1747 (N_1747,N_806,N_294);
or U1748 (N_1748,N_899,N_725);
or U1749 (N_1749,N_237,N_532);
nor U1750 (N_1750,N_713,N_416);
nor U1751 (N_1751,N_258,N_281);
nand U1752 (N_1752,N_794,N_38);
or U1753 (N_1753,N_954,N_820);
nor U1754 (N_1754,N_272,N_361);
or U1755 (N_1755,N_485,N_165);
or U1756 (N_1756,N_245,N_322);
nand U1757 (N_1757,N_307,N_584);
and U1758 (N_1758,N_844,N_369);
and U1759 (N_1759,N_82,N_449);
or U1760 (N_1760,N_816,N_230);
and U1761 (N_1761,N_397,N_294);
and U1762 (N_1762,N_472,N_887);
and U1763 (N_1763,N_442,N_495);
nor U1764 (N_1764,N_126,N_925);
or U1765 (N_1765,N_185,N_79);
and U1766 (N_1766,N_744,N_188);
nor U1767 (N_1767,N_941,N_36);
and U1768 (N_1768,N_409,N_348);
and U1769 (N_1769,N_719,N_487);
nand U1770 (N_1770,N_860,N_877);
nor U1771 (N_1771,N_187,N_388);
or U1772 (N_1772,N_329,N_911);
or U1773 (N_1773,N_859,N_145);
nand U1774 (N_1774,N_26,N_397);
nand U1775 (N_1775,N_265,N_61);
or U1776 (N_1776,N_480,N_77);
nand U1777 (N_1777,N_14,N_335);
nor U1778 (N_1778,N_769,N_903);
nor U1779 (N_1779,N_584,N_110);
or U1780 (N_1780,N_477,N_965);
nand U1781 (N_1781,N_769,N_357);
nand U1782 (N_1782,N_110,N_444);
nand U1783 (N_1783,N_792,N_732);
or U1784 (N_1784,N_682,N_592);
nand U1785 (N_1785,N_415,N_176);
and U1786 (N_1786,N_734,N_352);
and U1787 (N_1787,N_801,N_525);
and U1788 (N_1788,N_373,N_530);
or U1789 (N_1789,N_926,N_946);
or U1790 (N_1790,N_864,N_247);
or U1791 (N_1791,N_533,N_894);
nand U1792 (N_1792,N_220,N_389);
or U1793 (N_1793,N_236,N_291);
or U1794 (N_1794,N_230,N_973);
nand U1795 (N_1795,N_956,N_999);
nand U1796 (N_1796,N_706,N_581);
nand U1797 (N_1797,N_640,N_535);
or U1798 (N_1798,N_996,N_472);
or U1799 (N_1799,N_690,N_536);
or U1800 (N_1800,N_354,N_632);
nor U1801 (N_1801,N_857,N_723);
nor U1802 (N_1802,N_210,N_992);
and U1803 (N_1803,N_896,N_815);
or U1804 (N_1804,N_460,N_405);
or U1805 (N_1805,N_598,N_881);
and U1806 (N_1806,N_654,N_273);
nand U1807 (N_1807,N_59,N_257);
nor U1808 (N_1808,N_474,N_540);
and U1809 (N_1809,N_724,N_288);
nor U1810 (N_1810,N_109,N_692);
nand U1811 (N_1811,N_988,N_844);
or U1812 (N_1812,N_859,N_598);
nand U1813 (N_1813,N_575,N_931);
or U1814 (N_1814,N_441,N_897);
or U1815 (N_1815,N_437,N_632);
or U1816 (N_1816,N_21,N_992);
or U1817 (N_1817,N_518,N_647);
nor U1818 (N_1818,N_163,N_956);
or U1819 (N_1819,N_915,N_251);
nand U1820 (N_1820,N_105,N_836);
or U1821 (N_1821,N_660,N_890);
nand U1822 (N_1822,N_294,N_760);
nand U1823 (N_1823,N_750,N_518);
or U1824 (N_1824,N_340,N_856);
nand U1825 (N_1825,N_727,N_665);
or U1826 (N_1826,N_642,N_836);
nor U1827 (N_1827,N_268,N_939);
and U1828 (N_1828,N_659,N_493);
and U1829 (N_1829,N_680,N_159);
nor U1830 (N_1830,N_676,N_229);
or U1831 (N_1831,N_765,N_858);
nand U1832 (N_1832,N_434,N_551);
nand U1833 (N_1833,N_944,N_200);
and U1834 (N_1834,N_497,N_809);
nand U1835 (N_1835,N_332,N_9);
and U1836 (N_1836,N_250,N_122);
and U1837 (N_1837,N_529,N_485);
or U1838 (N_1838,N_755,N_679);
nand U1839 (N_1839,N_557,N_415);
nor U1840 (N_1840,N_701,N_489);
and U1841 (N_1841,N_439,N_274);
nand U1842 (N_1842,N_377,N_619);
xor U1843 (N_1843,N_92,N_920);
nand U1844 (N_1844,N_215,N_71);
and U1845 (N_1845,N_751,N_488);
nor U1846 (N_1846,N_446,N_866);
or U1847 (N_1847,N_962,N_918);
and U1848 (N_1848,N_123,N_990);
or U1849 (N_1849,N_344,N_608);
nor U1850 (N_1850,N_875,N_427);
nor U1851 (N_1851,N_602,N_799);
and U1852 (N_1852,N_794,N_830);
and U1853 (N_1853,N_112,N_334);
or U1854 (N_1854,N_864,N_603);
nand U1855 (N_1855,N_128,N_942);
or U1856 (N_1856,N_799,N_184);
nor U1857 (N_1857,N_283,N_222);
nor U1858 (N_1858,N_488,N_893);
nand U1859 (N_1859,N_63,N_680);
and U1860 (N_1860,N_517,N_981);
or U1861 (N_1861,N_317,N_218);
nor U1862 (N_1862,N_671,N_271);
nor U1863 (N_1863,N_665,N_569);
nor U1864 (N_1864,N_795,N_871);
nor U1865 (N_1865,N_835,N_347);
or U1866 (N_1866,N_339,N_517);
nand U1867 (N_1867,N_471,N_99);
nor U1868 (N_1868,N_814,N_609);
nor U1869 (N_1869,N_475,N_922);
nand U1870 (N_1870,N_390,N_35);
nor U1871 (N_1871,N_233,N_976);
nand U1872 (N_1872,N_448,N_570);
nor U1873 (N_1873,N_42,N_725);
nor U1874 (N_1874,N_311,N_428);
nor U1875 (N_1875,N_184,N_85);
xor U1876 (N_1876,N_930,N_178);
nor U1877 (N_1877,N_484,N_250);
nor U1878 (N_1878,N_647,N_558);
nand U1879 (N_1879,N_738,N_756);
and U1880 (N_1880,N_248,N_338);
nand U1881 (N_1881,N_419,N_756);
nor U1882 (N_1882,N_470,N_251);
nor U1883 (N_1883,N_266,N_993);
nand U1884 (N_1884,N_156,N_143);
and U1885 (N_1885,N_52,N_456);
nand U1886 (N_1886,N_181,N_818);
xnor U1887 (N_1887,N_546,N_311);
nor U1888 (N_1888,N_270,N_42);
nand U1889 (N_1889,N_227,N_708);
or U1890 (N_1890,N_587,N_145);
or U1891 (N_1891,N_524,N_485);
and U1892 (N_1892,N_668,N_510);
or U1893 (N_1893,N_913,N_377);
nand U1894 (N_1894,N_66,N_788);
and U1895 (N_1895,N_297,N_83);
nor U1896 (N_1896,N_600,N_44);
or U1897 (N_1897,N_287,N_832);
nand U1898 (N_1898,N_362,N_669);
nor U1899 (N_1899,N_607,N_139);
or U1900 (N_1900,N_366,N_211);
nor U1901 (N_1901,N_108,N_836);
nor U1902 (N_1902,N_103,N_898);
nor U1903 (N_1903,N_74,N_227);
and U1904 (N_1904,N_429,N_500);
nand U1905 (N_1905,N_633,N_168);
and U1906 (N_1906,N_449,N_788);
or U1907 (N_1907,N_131,N_6);
nand U1908 (N_1908,N_518,N_390);
and U1909 (N_1909,N_932,N_572);
or U1910 (N_1910,N_427,N_111);
or U1911 (N_1911,N_639,N_400);
nor U1912 (N_1912,N_386,N_221);
or U1913 (N_1913,N_867,N_804);
and U1914 (N_1914,N_562,N_713);
nand U1915 (N_1915,N_98,N_678);
or U1916 (N_1916,N_841,N_793);
or U1917 (N_1917,N_161,N_782);
nor U1918 (N_1918,N_44,N_240);
and U1919 (N_1919,N_282,N_359);
or U1920 (N_1920,N_499,N_382);
and U1921 (N_1921,N_387,N_485);
or U1922 (N_1922,N_199,N_707);
nor U1923 (N_1923,N_955,N_713);
nand U1924 (N_1924,N_241,N_109);
or U1925 (N_1925,N_671,N_812);
nor U1926 (N_1926,N_525,N_464);
nor U1927 (N_1927,N_892,N_794);
and U1928 (N_1928,N_997,N_112);
or U1929 (N_1929,N_405,N_408);
nor U1930 (N_1930,N_25,N_534);
and U1931 (N_1931,N_503,N_648);
nand U1932 (N_1932,N_894,N_724);
and U1933 (N_1933,N_971,N_184);
or U1934 (N_1934,N_412,N_785);
or U1935 (N_1935,N_181,N_441);
nand U1936 (N_1936,N_536,N_299);
and U1937 (N_1937,N_220,N_969);
nor U1938 (N_1938,N_323,N_538);
or U1939 (N_1939,N_463,N_152);
or U1940 (N_1940,N_249,N_421);
and U1941 (N_1941,N_616,N_865);
or U1942 (N_1942,N_697,N_973);
and U1943 (N_1943,N_291,N_247);
nor U1944 (N_1944,N_352,N_255);
or U1945 (N_1945,N_905,N_403);
or U1946 (N_1946,N_885,N_429);
nor U1947 (N_1947,N_227,N_812);
and U1948 (N_1948,N_743,N_72);
nor U1949 (N_1949,N_611,N_389);
or U1950 (N_1950,N_217,N_398);
nor U1951 (N_1951,N_483,N_391);
and U1952 (N_1952,N_463,N_481);
or U1953 (N_1953,N_57,N_182);
or U1954 (N_1954,N_236,N_303);
and U1955 (N_1955,N_80,N_258);
nor U1956 (N_1956,N_336,N_461);
nand U1957 (N_1957,N_824,N_27);
nor U1958 (N_1958,N_183,N_338);
nand U1959 (N_1959,N_621,N_55);
xor U1960 (N_1960,N_638,N_419);
or U1961 (N_1961,N_960,N_961);
nand U1962 (N_1962,N_961,N_905);
or U1963 (N_1963,N_619,N_227);
nand U1964 (N_1964,N_13,N_306);
or U1965 (N_1965,N_973,N_139);
and U1966 (N_1966,N_299,N_485);
or U1967 (N_1967,N_823,N_795);
nand U1968 (N_1968,N_448,N_820);
nor U1969 (N_1969,N_784,N_454);
nand U1970 (N_1970,N_526,N_701);
and U1971 (N_1971,N_89,N_433);
nand U1972 (N_1972,N_579,N_837);
and U1973 (N_1973,N_307,N_417);
and U1974 (N_1974,N_539,N_105);
nand U1975 (N_1975,N_573,N_434);
or U1976 (N_1976,N_922,N_10);
nand U1977 (N_1977,N_983,N_841);
and U1978 (N_1978,N_565,N_71);
nand U1979 (N_1979,N_144,N_162);
and U1980 (N_1980,N_137,N_535);
nand U1981 (N_1981,N_979,N_108);
nor U1982 (N_1982,N_614,N_793);
and U1983 (N_1983,N_836,N_887);
nor U1984 (N_1984,N_768,N_593);
or U1985 (N_1985,N_60,N_102);
or U1986 (N_1986,N_595,N_567);
nor U1987 (N_1987,N_325,N_153);
nor U1988 (N_1988,N_992,N_829);
nand U1989 (N_1989,N_439,N_202);
nor U1990 (N_1990,N_736,N_539);
and U1991 (N_1991,N_550,N_767);
xor U1992 (N_1992,N_272,N_113);
nor U1993 (N_1993,N_845,N_858);
or U1994 (N_1994,N_486,N_60);
nor U1995 (N_1995,N_231,N_789);
nor U1996 (N_1996,N_150,N_279);
nand U1997 (N_1997,N_960,N_746);
nor U1998 (N_1998,N_510,N_84);
and U1999 (N_1999,N_319,N_32);
nand U2000 (N_2000,N_1202,N_1158);
nand U2001 (N_2001,N_1298,N_1626);
and U2002 (N_2002,N_1361,N_1805);
or U2003 (N_2003,N_1827,N_1146);
or U2004 (N_2004,N_1223,N_1166);
nor U2005 (N_2005,N_1544,N_1157);
nand U2006 (N_2006,N_1501,N_1760);
nand U2007 (N_2007,N_1715,N_1155);
or U2008 (N_2008,N_1232,N_1914);
nand U2009 (N_2009,N_1791,N_1987);
and U2010 (N_2010,N_1034,N_1741);
or U2011 (N_2011,N_1488,N_1210);
nand U2012 (N_2012,N_1005,N_1369);
and U2013 (N_2013,N_1968,N_1356);
and U2014 (N_2014,N_1265,N_1239);
nor U2015 (N_2015,N_1422,N_1958);
nand U2016 (N_2016,N_1830,N_1907);
or U2017 (N_2017,N_1744,N_1056);
and U2018 (N_2018,N_1342,N_1818);
nor U2019 (N_2019,N_1185,N_1776);
or U2020 (N_2020,N_1716,N_1226);
nand U2021 (N_2021,N_1974,N_1785);
and U2022 (N_2022,N_1217,N_1855);
nand U2023 (N_2023,N_1296,N_1896);
or U2024 (N_2024,N_1929,N_1343);
and U2025 (N_2025,N_1534,N_1360);
and U2026 (N_2026,N_1559,N_1992);
and U2027 (N_2027,N_1708,N_1611);
nand U2028 (N_2028,N_1364,N_1581);
or U2029 (N_2029,N_1172,N_1551);
and U2030 (N_2030,N_1315,N_1354);
or U2031 (N_2031,N_1413,N_1850);
or U2032 (N_2032,N_1114,N_1746);
and U2033 (N_2033,N_1765,N_1464);
nor U2034 (N_2034,N_1523,N_1379);
nand U2035 (N_2035,N_1200,N_1740);
or U2036 (N_2036,N_1527,N_1206);
and U2037 (N_2037,N_1717,N_1510);
nand U2038 (N_2038,N_1045,N_1489);
nor U2039 (N_2039,N_1171,N_1231);
and U2040 (N_2040,N_1757,N_1605);
nor U2041 (N_2041,N_1684,N_1745);
nor U2042 (N_2042,N_1869,N_1181);
nor U2043 (N_2043,N_1552,N_1937);
and U2044 (N_2044,N_1040,N_1083);
or U2045 (N_2045,N_1766,N_1951);
nor U2046 (N_2046,N_1052,N_1648);
or U2047 (N_2047,N_1486,N_1883);
nor U2048 (N_2048,N_1313,N_1060);
nand U2049 (N_2049,N_1505,N_1508);
nor U2050 (N_2050,N_1945,N_1768);
and U2051 (N_2051,N_1152,N_1407);
and U2052 (N_2052,N_1685,N_1906);
nor U2053 (N_2053,N_1334,N_1917);
or U2054 (N_2054,N_1008,N_1738);
nor U2055 (N_2055,N_1997,N_1899);
and U2056 (N_2056,N_1151,N_1509);
nor U2057 (N_2057,N_1310,N_1555);
or U2058 (N_2058,N_1779,N_1991);
nand U2059 (N_2059,N_1507,N_1292);
and U2060 (N_2060,N_1366,N_1935);
nand U2061 (N_2061,N_1886,N_1731);
nor U2062 (N_2062,N_1936,N_1515);
or U2063 (N_2063,N_1299,N_1859);
nand U2064 (N_2064,N_1763,N_1520);
nand U2065 (N_2065,N_1112,N_1681);
nor U2066 (N_2066,N_1032,N_1982);
or U2067 (N_2067,N_1088,N_1759);
or U2068 (N_2068,N_1405,N_1988);
xor U2069 (N_2069,N_1687,N_1624);
nand U2070 (N_2070,N_1260,N_1482);
nand U2071 (N_2071,N_1538,N_1621);
nor U2072 (N_2072,N_1102,N_1294);
or U2073 (N_2073,N_1762,N_1126);
nand U2074 (N_2074,N_1353,N_1182);
nand U2075 (N_2075,N_1129,N_1915);
or U2076 (N_2076,N_1381,N_1051);
nand U2077 (N_2077,N_1363,N_1625);
and U2078 (N_2078,N_1068,N_1478);
nand U2079 (N_2079,N_1355,N_1093);
or U2080 (N_2080,N_1638,N_1054);
or U2081 (N_2081,N_1016,N_1517);
or U2082 (N_2082,N_1655,N_1100);
nand U2083 (N_2083,N_1325,N_1187);
nor U2084 (N_2084,N_1807,N_1575);
nor U2085 (N_2085,N_1007,N_1604);
and U2086 (N_2086,N_1404,N_1423);
and U2087 (N_2087,N_1536,N_1341);
nand U2088 (N_2088,N_1673,N_1639);
nor U2089 (N_2089,N_1878,N_1911);
nor U2090 (N_2090,N_1814,N_1709);
nand U2091 (N_2091,N_1980,N_1011);
or U2092 (N_2092,N_1944,N_1468);
or U2093 (N_2093,N_1280,N_1029);
nor U2094 (N_2094,N_1981,N_1970);
nand U2095 (N_2095,N_1619,N_1679);
nor U2096 (N_2096,N_1594,N_1872);
and U2097 (N_2097,N_1309,N_1119);
nor U2098 (N_2098,N_1756,N_1730);
or U2099 (N_2099,N_1326,N_1149);
nand U2100 (N_2100,N_1449,N_1487);
xnor U2101 (N_2101,N_1824,N_1108);
xor U2102 (N_2102,N_1408,N_1771);
nor U2103 (N_2103,N_1380,N_1703);
nand U2104 (N_2104,N_1868,N_1925);
and U2105 (N_2105,N_1454,N_1021);
nand U2106 (N_2106,N_1680,N_1165);
or U2107 (N_2107,N_1026,N_1793);
nand U2108 (N_2108,N_1522,N_1122);
and U2109 (N_2109,N_1645,N_1257);
or U2110 (N_2110,N_1456,N_1316);
or U2111 (N_2111,N_1751,N_1568);
and U2112 (N_2112,N_1263,N_1349);
and U2113 (N_2113,N_1173,N_1601);
nor U2114 (N_2114,N_1588,N_1537);
nor U2115 (N_2115,N_1030,N_1599);
nand U2116 (N_2116,N_1177,N_1993);
or U2117 (N_2117,N_1526,N_1547);
or U2118 (N_2118,N_1311,N_1339);
or U2119 (N_2119,N_1632,N_1983);
nor U2120 (N_2120,N_1403,N_1127);
or U2121 (N_2121,N_1495,N_1590);
nand U2122 (N_2122,N_1261,N_1038);
nand U2123 (N_2123,N_1873,N_1284);
or U2124 (N_2124,N_1041,N_1887);
or U2125 (N_2125,N_1282,N_1840);
nor U2126 (N_2126,N_1367,N_1233);
nand U2127 (N_2127,N_1305,N_1193);
nand U2128 (N_2128,N_1434,N_1195);
nand U2129 (N_2129,N_1365,N_1490);
nor U2130 (N_2130,N_1163,N_1711);
and U2131 (N_2131,N_1714,N_1994);
and U2132 (N_2132,N_1373,N_1104);
or U2133 (N_2133,N_1203,N_1494);
nor U2134 (N_2134,N_1137,N_1235);
and U2135 (N_2135,N_1596,N_1909);
and U2136 (N_2136,N_1159,N_1053);
or U2137 (N_2137,N_1270,N_1323);
and U2138 (N_2138,N_1246,N_1216);
nor U2139 (N_2139,N_1739,N_1245);
nand U2140 (N_2140,N_1875,N_1242);
and U2141 (N_2141,N_1585,N_1975);
and U2142 (N_2142,N_1044,N_1389);
nor U2143 (N_2143,N_1258,N_1902);
nand U2144 (N_2144,N_1368,N_1212);
xnor U2145 (N_2145,N_1276,N_1941);
or U2146 (N_2146,N_1701,N_1147);
and U2147 (N_2147,N_1448,N_1416);
or U2148 (N_2148,N_1497,N_1699);
or U2149 (N_2149,N_1096,N_1782);
nor U2150 (N_2150,N_1792,N_1479);
nor U2151 (N_2151,N_1065,N_1786);
nor U2152 (N_2152,N_1848,N_1672);
and U2153 (N_2153,N_1773,N_1338);
nor U2154 (N_2154,N_1787,N_1291);
nand U2155 (N_2155,N_1635,N_1075);
xor U2156 (N_2156,N_1682,N_1653);
nand U2157 (N_2157,N_1721,N_1283);
and U2158 (N_2158,N_1586,N_1560);
nor U2159 (N_2159,N_1188,N_1806);
nand U2160 (N_2160,N_1749,N_1607);
nor U2161 (N_2161,N_1074,N_1098);
nor U2162 (N_2162,N_1058,N_1895);
and U2163 (N_2163,N_1199,N_1308);
nor U2164 (N_2164,N_1804,N_1829);
xnor U2165 (N_2165,N_1161,N_1406);
nand U2166 (N_2166,N_1928,N_1014);
or U2167 (N_2167,N_1630,N_1566);
nand U2168 (N_2168,N_1640,N_1080);
nand U2169 (N_2169,N_1811,N_1402);
and U2170 (N_2170,N_1301,N_1481);
or U2171 (N_2171,N_1399,N_1854);
nor U2172 (N_2172,N_1207,N_1750);
nor U2173 (N_2173,N_1264,N_1634);
nand U2174 (N_2174,N_1472,N_1591);
nand U2175 (N_2175,N_1861,N_1857);
nor U2176 (N_2176,N_1908,N_1947);
nor U2177 (N_2177,N_1437,N_1595);
or U2178 (N_2178,N_1965,N_1251);
nand U2179 (N_2179,N_1531,N_1557);
nand U2180 (N_2180,N_1105,N_1447);
nor U2181 (N_2181,N_1256,N_1274);
nand U2182 (N_2182,N_1345,N_1015);
or U2183 (N_2183,N_1962,N_1237);
nor U2184 (N_2184,N_1204,N_1898);
nand U2185 (N_2185,N_1115,N_1860);
nand U2186 (N_2186,N_1395,N_1241);
or U2187 (N_2187,N_1583,N_1775);
and U2188 (N_2188,N_1894,N_1225);
nor U2189 (N_2189,N_1117,N_1485);
and U2190 (N_2190,N_1278,N_1304);
nand U2191 (N_2191,N_1977,N_1229);
and U2192 (N_2192,N_1162,N_1694);
and U2193 (N_2193,N_1042,N_1973);
or U2194 (N_2194,N_1417,N_1372);
and U2195 (N_2195,N_1238,N_1192);
and U2196 (N_2196,N_1781,N_1702);
or U2197 (N_2197,N_1332,N_1135);
nor U2198 (N_2198,N_1259,N_1059);
and U2199 (N_2199,N_1445,N_1144);
nand U2200 (N_2200,N_1153,N_1427);
nor U2201 (N_2201,N_1674,N_1921);
nor U2202 (N_2202,N_1003,N_1443);
nand U2203 (N_2203,N_1118,N_1211);
or U2204 (N_2204,N_1397,N_1213);
and U2205 (N_2205,N_1543,N_1101);
or U2206 (N_2206,N_1580,N_1451);
and U2207 (N_2207,N_1039,N_1574);
nor U2208 (N_2208,N_1554,N_1004);
or U2209 (N_2209,N_1669,N_1504);
or U2210 (N_2210,N_1132,N_1984);
or U2211 (N_2211,N_1167,N_1371);
and U2212 (N_2212,N_1772,N_1518);
or U2213 (N_2213,N_1348,N_1067);
nor U2214 (N_2214,N_1589,N_1441);
nor U2215 (N_2215,N_1573,N_1459);
and U2216 (N_2216,N_1475,N_1664);
and U2217 (N_2217,N_1603,N_1963);
and U2218 (N_2218,N_1277,N_1808);
nand U2219 (N_2219,N_1866,N_1424);
nor U2220 (N_2220,N_1871,N_1484);
or U2221 (N_2221,N_1198,N_1795);
nor U2222 (N_2222,N_1946,N_1374);
nand U2223 (N_2223,N_1327,N_1724);
or U2224 (N_2224,N_1483,N_1667);
and U2225 (N_2225,N_1753,N_1440);
nor U2226 (N_2226,N_1950,N_1500);
or U2227 (N_2227,N_1357,N_1387);
nor U2228 (N_2228,N_1613,N_1439);
nor U2229 (N_2229,N_1659,N_1577);
or U2230 (N_2230,N_1512,N_1697);
or U2231 (N_2231,N_1706,N_1723);
nand U2232 (N_2232,N_1492,N_1470);
nor U2233 (N_2233,N_1436,N_1670);
or U2234 (N_2234,N_1932,N_1428);
xor U2235 (N_2235,N_1764,N_1183);
or U2236 (N_2236,N_1879,N_1430);
nand U2237 (N_2237,N_1136,N_1617);
nor U2238 (N_2238,N_1322,N_1453);
nand U2239 (N_2239,N_1817,N_1650);
or U2240 (N_2240,N_1462,N_1734);
and U2241 (N_2241,N_1948,N_1598);
nor U2242 (N_2242,N_1143,N_1156);
or U2243 (N_2243,N_1446,N_1286);
or U2244 (N_2244,N_1769,N_1471);
xnor U2245 (N_2245,N_1657,N_1934);
or U2246 (N_2246,N_1602,N_1689);
and U2247 (N_2247,N_1073,N_1031);
or U2248 (N_2248,N_1838,N_1333);
and U2249 (N_2249,N_1018,N_1966);
nor U2250 (N_2250,N_1839,N_1912);
or U2251 (N_2251,N_1616,N_1415);
or U2252 (N_2252,N_1180,N_1215);
nor U2253 (N_2253,N_1396,N_1972);
nand U2254 (N_2254,N_1091,N_1425);
or U2255 (N_2255,N_1747,N_1656);
or U2256 (N_2256,N_1230,N_1567);
nand U2257 (N_2257,N_1019,N_1922);
nor U2258 (N_2258,N_1995,N_1778);
nand U2259 (N_2259,N_1275,N_1633);
nand U2260 (N_2260,N_1642,N_1130);
and U2261 (N_2261,N_1438,N_1222);
nand U2262 (N_2262,N_1240,N_1465);
nand U2263 (N_2263,N_1877,N_1208);
nand U2264 (N_2264,N_1797,N_1600);
xnor U2265 (N_2265,N_1272,N_1777);
and U2266 (N_2266,N_1606,N_1513);
or U2267 (N_2267,N_1178,N_1477);
nand U2268 (N_2268,N_1224,N_1758);
or U2269 (N_2269,N_1248,N_1087);
and U2270 (N_2270,N_1710,N_1281);
and U2271 (N_2271,N_1111,N_1964);
and U2272 (N_2272,N_1141,N_1578);
nor U2273 (N_2273,N_1347,N_1300);
and U2274 (N_2274,N_1287,N_1418);
or U2275 (N_2275,N_1466,N_1062);
or U2276 (N_2276,N_1884,N_1535);
nand U2277 (N_2277,N_1770,N_1121);
nand U2278 (N_2278,N_1939,N_1061);
and U2279 (N_2279,N_1521,N_1097);
or U2280 (N_2280,N_1138,N_1893);
nand U2281 (N_2281,N_1079,N_1221);
or U2282 (N_2282,N_1214,N_1996);
nand U2283 (N_2283,N_1120,N_1089);
nand U2284 (N_2284,N_1641,N_1849);
and U2285 (N_2285,N_1463,N_1072);
or U2286 (N_2286,N_1092,N_1285);
nor U2287 (N_2287,N_1103,N_1558);
nand U2288 (N_2288,N_1978,N_1442);
or U2289 (N_2289,N_1385,N_1823);
nand U2290 (N_2290,N_1023,N_1954);
nand U2291 (N_2291,N_1289,N_1306);
and U2292 (N_2292,N_1433,N_1913);
xor U2293 (N_2293,N_1450,N_1660);
and U2294 (N_2294,N_1796,N_1570);
nor U2295 (N_2295,N_1190,N_1812);
nand U2296 (N_2296,N_1125,N_1870);
nor U2297 (N_2297,N_1903,N_1094);
nand U2298 (N_2298,N_1789,N_1057);
nand U2299 (N_2299,N_1048,N_1351);
nand U2300 (N_2300,N_1476,N_1455);
and U2301 (N_2301,N_1234,N_1002);
nor U2302 (N_2302,N_1761,N_1754);
nor U2303 (N_2303,N_1295,N_1401);
or U2304 (N_2304,N_1540,N_1525);
nor U2305 (N_2305,N_1228,N_1565);
nor U2306 (N_2306,N_1362,N_1627);
or U2307 (N_2307,N_1196,N_1790);
nand U2308 (N_2308,N_1064,N_1001);
xor U2309 (N_2309,N_1955,N_1688);
and U2310 (N_2310,N_1006,N_1255);
and U2311 (N_2311,N_1891,N_1546);
and U2312 (N_2312,N_1961,N_1169);
nor U2313 (N_2313,N_1267,N_1279);
nand U2314 (N_2314,N_1086,N_1736);
and U2315 (N_2315,N_1391,N_1825);
and U2316 (N_2316,N_1841,N_1429);
or U2317 (N_2317,N_1545,N_1550);
nand U2318 (N_2318,N_1113,N_1249);
nor U2319 (N_2319,N_1250,N_1035);
or U2320 (N_2320,N_1020,N_1133);
nand U2321 (N_2321,N_1923,N_1931);
nand U2322 (N_2322,N_1317,N_1506);
and U2323 (N_2323,N_1665,N_1066);
or U2324 (N_2324,N_1563,N_1219);
nand U2325 (N_2325,N_1095,N_1375);
nand U2326 (N_2326,N_1678,N_1957);
nor U2327 (N_2327,N_1220,N_1106);
nor U2328 (N_2328,N_1847,N_1358);
or U2329 (N_2329,N_1022,N_1432);
nand U2330 (N_2330,N_1168,N_1370);
nand U2331 (N_2331,N_1646,N_1880);
and U2332 (N_2332,N_1910,N_1969);
nand U2333 (N_2333,N_1856,N_1392);
nor U2334 (N_2334,N_1046,N_1346);
nand U2335 (N_2335,N_1986,N_1658);
or U2336 (N_2336,N_1549,N_1302);
nor U2337 (N_2337,N_1253,N_1556);
nor U2338 (N_2338,N_1890,N_1844);
nand U2339 (N_2339,N_1836,N_1989);
or U2340 (N_2340,N_1191,N_1835);
or U2341 (N_2341,N_1400,N_1393);
nor U2342 (N_2342,N_1078,N_1107);
nor U2343 (N_2343,N_1900,N_1542);
or U2344 (N_2344,N_1410,N_1131);
nand U2345 (N_2345,N_1904,N_1612);
and U2346 (N_2346,N_1533,N_1853);
and U2347 (N_2347,N_1767,N_1189);
and U2348 (N_2348,N_1718,N_1644);
nor U2349 (N_2349,N_1254,N_1412);
or U2350 (N_2350,N_1201,N_1288);
or U2351 (N_2351,N_1597,N_1938);
nand U2352 (N_2352,N_1524,N_1124);
nor U2353 (N_2353,N_1328,N_1319);
nor U2354 (N_2354,N_1729,N_1394);
or U2355 (N_2355,N_1419,N_1918);
nor U2356 (N_2356,N_1892,N_1452);
and U2357 (N_2357,N_1378,N_1426);
nor U2358 (N_2358,N_1676,N_1318);
and U2359 (N_2359,N_1919,N_1331);
nor U2360 (N_2360,N_1979,N_1649);
or U2361 (N_2361,N_1218,N_1514);
or U2362 (N_2362,N_1809,N_1592);
nand U2363 (N_2363,N_1615,N_1541);
nor U2364 (N_2364,N_1852,N_1502);
nor U2365 (N_2365,N_1735,N_1109);
and U2366 (N_2366,N_1637,N_1321);
nand U2367 (N_2367,N_1608,N_1082);
nor U2368 (N_2368,N_1435,N_1268);
nand U2369 (N_2369,N_1695,N_1561);
nor U2370 (N_2370,N_1050,N_1047);
and U2371 (N_2371,N_1942,N_1949);
nand U2372 (N_2372,N_1794,N_1384);
or U2373 (N_2373,N_1874,N_1421);
xnor U2374 (N_2374,N_1473,N_1071);
or U2375 (N_2375,N_1273,N_1352);
nor U2376 (N_2376,N_1828,N_1085);
or U2377 (N_2377,N_1142,N_1614);
or U2378 (N_2378,N_1532,N_1376);
nor U2379 (N_2379,N_1247,N_1150);
nor U2380 (N_2380,N_1139,N_1810);
xnor U2381 (N_2381,N_1564,N_1084);
nand U2382 (N_2382,N_1314,N_1123);
nor U2383 (N_2383,N_1713,N_1335);
or U2384 (N_2384,N_1174,N_1388);
and U2385 (N_2385,N_1845,N_1290);
and U2386 (N_2386,N_1553,N_1293);
nor U2387 (N_2387,N_1755,N_1926);
or U2388 (N_2388,N_1788,N_1145);
and U2389 (N_2389,N_1693,N_1010);
nor U2390 (N_2390,N_1712,N_1800);
nand U2391 (N_2391,N_1186,N_1076);
nor U2392 (N_2392,N_1832,N_1460);
nand U2393 (N_2393,N_1227,N_1269);
nor U2394 (N_2394,N_1843,N_1205);
nor U2395 (N_2395,N_1266,N_1737);
nand U2396 (N_2396,N_1698,N_1519);
or U2397 (N_2397,N_1742,N_1028);
or U2398 (N_2398,N_1069,N_1834);
nand U2399 (N_2399,N_1569,N_1528);
nand U2400 (N_2400,N_1382,N_1386);
nor U2401 (N_2401,N_1511,N_1831);
nand U2402 (N_2402,N_1865,N_1628);
or U2403 (N_2403,N_1197,N_1833);
or U2404 (N_2404,N_1726,N_1622);
and U2405 (N_2405,N_1036,N_1176);
nand U2406 (N_2406,N_1683,N_1976);
nand U2407 (N_2407,N_1572,N_1236);
and U2408 (N_2408,N_1055,N_1889);
or U2409 (N_2409,N_1390,N_1692);
and U2410 (N_2410,N_1337,N_1705);
or U2411 (N_2411,N_1457,N_1803);
and U2412 (N_2412,N_1691,N_1733);
or U2413 (N_2413,N_1467,N_1184);
nand U2414 (N_2414,N_1043,N_1728);
nand U2415 (N_2415,N_1330,N_1013);
and U2416 (N_2416,N_1398,N_1815);
or U2417 (N_2417,N_1732,N_1774);
nand U2418 (N_2418,N_1480,N_1303);
nor U2419 (N_2419,N_1539,N_1491);
nand U2420 (N_2420,N_1798,N_1312);
nor U2421 (N_2421,N_1668,N_1444);
or U2422 (N_2422,N_1933,N_1110);
nor U2423 (N_2423,N_1985,N_1858);
and U2424 (N_2424,N_1643,N_1820);
nand U2425 (N_2425,N_1340,N_1881);
nor U2426 (N_2426,N_1920,N_1458);
nand U2427 (N_2427,N_1888,N_1671);
nand U2428 (N_2428,N_1722,N_1516);
nor U2429 (N_2429,N_1905,N_1719);
or U2430 (N_2430,N_1837,N_1179);
and U2431 (N_2431,N_1952,N_1324);
nand U2432 (N_2432,N_1049,N_1474);
nand U2433 (N_2433,N_1846,N_1647);
nor U2434 (N_2434,N_1307,N_1027);
nand U2435 (N_2435,N_1209,N_1576);
and U2436 (N_2436,N_1940,N_1725);
nor U2437 (N_2437,N_1009,N_1675);
and U2438 (N_2438,N_1562,N_1999);
nand U2439 (N_2439,N_1953,N_1593);
and U2440 (N_2440,N_1037,N_1024);
nor U2441 (N_2441,N_1461,N_1727);
nand U2442 (N_2442,N_1243,N_1496);
or U2443 (N_2443,N_1377,N_1498);
or U2444 (N_2444,N_1863,N_1700);
nor U2445 (N_2445,N_1099,N_1529);
nand U2446 (N_2446,N_1677,N_1956);
xor U2447 (N_2447,N_1587,N_1017);
or U2448 (N_2448,N_1662,N_1943);
nor U2449 (N_2449,N_1784,N_1081);
nor U2450 (N_2450,N_1194,N_1244);
or U2451 (N_2451,N_1148,N_1383);
nand U2452 (N_2452,N_1897,N_1707);
nor U2453 (N_2453,N_1164,N_1609);
nor U2454 (N_2454,N_1025,N_1651);
xnor U2455 (N_2455,N_1901,N_1420);
nor U2456 (N_2456,N_1320,N_1629);
nand U2457 (N_2457,N_1620,N_1801);
and U2458 (N_2458,N_1431,N_1990);
and U2459 (N_2459,N_1499,N_1652);
nand U2460 (N_2460,N_1134,N_1160);
nand U2461 (N_2461,N_1584,N_1864);
nor U2462 (N_2462,N_1170,N_1821);
nor U2463 (N_2463,N_1618,N_1867);
and U2464 (N_2464,N_1816,N_1359);
nor U2465 (N_2465,N_1012,N_1579);
or U2466 (N_2466,N_1882,N_1876);
nor U2467 (N_2467,N_1262,N_1623);
and U2468 (N_2468,N_1885,N_1690);
nand U2469 (N_2469,N_1927,N_1631);
or U2470 (N_2470,N_1924,N_1411);
nor U2471 (N_2471,N_1822,N_1154);
or U2472 (N_2472,N_1826,N_1297);
and U2473 (N_2473,N_1503,N_1813);
nor U2474 (N_2474,N_1571,N_1842);
and U2475 (N_2475,N_1271,N_1252);
and U2476 (N_2476,N_1128,N_1802);
and U2477 (N_2477,N_1851,N_1654);
and U2478 (N_2478,N_1063,N_1530);
nand U2479 (N_2479,N_1819,N_1998);
nor U2480 (N_2480,N_1033,N_1960);
or U2481 (N_2481,N_1661,N_1862);
and U2482 (N_2482,N_1090,N_1582);
and U2483 (N_2483,N_1548,N_1663);
and U2484 (N_2484,N_1783,N_1967);
or U2485 (N_2485,N_1175,N_1666);
nor U2486 (N_2486,N_1140,N_1344);
or U2487 (N_2487,N_1077,N_1414);
nor U2488 (N_2488,N_1329,N_1636);
xor U2489 (N_2489,N_1959,N_1000);
and U2490 (N_2490,N_1780,N_1752);
nor U2491 (N_2491,N_1469,N_1799);
and U2492 (N_2492,N_1743,N_1930);
or U2493 (N_2493,N_1704,N_1350);
nand U2494 (N_2494,N_1493,N_1971);
nand U2495 (N_2495,N_1336,N_1070);
or U2496 (N_2496,N_1686,N_1748);
and U2497 (N_2497,N_1610,N_1916);
nor U2498 (N_2498,N_1720,N_1409);
nor U2499 (N_2499,N_1696,N_1116);
nor U2500 (N_2500,N_1836,N_1300);
or U2501 (N_2501,N_1121,N_1908);
nor U2502 (N_2502,N_1087,N_1712);
or U2503 (N_2503,N_1130,N_1330);
nand U2504 (N_2504,N_1982,N_1348);
nand U2505 (N_2505,N_1657,N_1360);
xor U2506 (N_2506,N_1086,N_1151);
nor U2507 (N_2507,N_1639,N_1148);
or U2508 (N_2508,N_1875,N_1889);
nor U2509 (N_2509,N_1770,N_1288);
nor U2510 (N_2510,N_1658,N_1283);
or U2511 (N_2511,N_1054,N_1335);
or U2512 (N_2512,N_1943,N_1186);
and U2513 (N_2513,N_1259,N_1465);
nand U2514 (N_2514,N_1764,N_1935);
nand U2515 (N_2515,N_1161,N_1555);
and U2516 (N_2516,N_1095,N_1505);
and U2517 (N_2517,N_1055,N_1565);
nor U2518 (N_2518,N_1493,N_1899);
or U2519 (N_2519,N_1857,N_1196);
or U2520 (N_2520,N_1102,N_1370);
nor U2521 (N_2521,N_1817,N_1616);
nor U2522 (N_2522,N_1551,N_1134);
nor U2523 (N_2523,N_1199,N_1875);
or U2524 (N_2524,N_1133,N_1855);
and U2525 (N_2525,N_1507,N_1442);
nand U2526 (N_2526,N_1972,N_1682);
and U2527 (N_2527,N_1765,N_1370);
or U2528 (N_2528,N_1144,N_1000);
nor U2529 (N_2529,N_1882,N_1379);
and U2530 (N_2530,N_1505,N_1567);
or U2531 (N_2531,N_1613,N_1106);
nand U2532 (N_2532,N_1293,N_1051);
nand U2533 (N_2533,N_1683,N_1838);
and U2534 (N_2534,N_1613,N_1737);
or U2535 (N_2535,N_1277,N_1460);
nor U2536 (N_2536,N_1820,N_1968);
xnor U2537 (N_2537,N_1205,N_1224);
nor U2538 (N_2538,N_1280,N_1500);
or U2539 (N_2539,N_1655,N_1592);
or U2540 (N_2540,N_1040,N_1567);
or U2541 (N_2541,N_1162,N_1081);
nand U2542 (N_2542,N_1126,N_1024);
nor U2543 (N_2543,N_1014,N_1792);
nor U2544 (N_2544,N_1548,N_1649);
and U2545 (N_2545,N_1180,N_1593);
nand U2546 (N_2546,N_1371,N_1383);
xor U2547 (N_2547,N_1711,N_1810);
nand U2548 (N_2548,N_1361,N_1968);
nand U2549 (N_2549,N_1839,N_1745);
or U2550 (N_2550,N_1420,N_1229);
or U2551 (N_2551,N_1330,N_1053);
nand U2552 (N_2552,N_1650,N_1000);
nand U2553 (N_2553,N_1971,N_1991);
or U2554 (N_2554,N_1443,N_1927);
nor U2555 (N_2555,N_1813,N_1465);
or U2556 (N_2556,N_1919,N_1323);
and U2557 (N_2557,N_1287,N_1769);
and U2558 (N_2558,N_1726,N_1254);
and U2559 (N_2559,N_1939,N_1677);
or U2560 (N_2560,N_1450,N_1390);
nor U2561 (N_2561,N_1067,N_1309);
nand U2562 (N_2562,N_1036,N_1983);
or U2563 (N_2563,N_1094,N_1397);
nand U2564 (N_2564,N_1868,N_1908);
nand U2565 (N_2565,N_1628,N_1428);
nand U2566 (N_2566,N_1147,N_1170);
and U2567 (N_2567,N_1618,N_1248);
nor U2568 (N_2568,N_1338,N_1532);
nor U2569 (N_2569,N_1913,N_1593);
and U2570 (N_2570,N_1805,N_1231);
nand U2571 (N_2571,N_1007,N_1991);
nand U2572 (N_2572,N_1662,N_1163);
nand U2573 (N_2573,N_1864,N_1078);
nand U2574 (N_2574,N_1602,N_1017);
nor U2575 (N_2575,N_1405,N_1896);
nand U2576 (N_2576,N_1043,N_1192);
nand U2577 (N_2577,N_1477,N_1200);
nand U2578 (N_2578,N_1239,N_1121);
nor U2579 (N_2579,N_1712,N_1161);
or U2580 (N_2580,N_1044,N_1080);
and U2581 (N_2581,N_1287,N_1397);
nand U2582 (N_2582,N_1829,N_1992);
nor U2583 (N_2583,N_1858,N_1418);
and U2584 (N_2584,N_1905,N_1909);
nand U2585 (N_2585,N_1284,N_1821);
nand U2586 (N_2586,N_1475,N_1920);
nand U2587 (N_2587,N_1461,N_1820);
and U2588 (N_2588,N_1161,N_1834);
or U2589 (N_2589,N_1402,N_1327);
nor U2590 (N_2590,N_1229,N_1893);
nor U2591 (N_2591,N_1660,N_1233);
nor U2592 (N_2592,N_1443,N_1694);
and U2593 (N_2593,N_1784,N_1604);
and U2594 (N_2594,N_1720,N_1775);
nor U2595 (N_2595,N_1520,N_1986);
nand U2596 (N_2596,N_1126,N_1858);
and U2597 (N_2597,N_1587,N_1577);
nand U2598 (N_2598,N_1008,N_1367);
nor U2599 (N_2599,N_1396,N_1288);
or U2600 (N_2600,N_1509,N_1341);
nor U2601 (N_2601,N_1271,N_1647);
or U2602 (N_2602,N_1679,N_1536);
or U2603 (N_2603,N_1422,N_1294);
nor U2604 (N_2604,N_1435,N_1385);
and U2605 (N_2605,N_1343,N_1706);
nand U2606 (N_2606,N_1592,N_1488);
or U2607 (N_2607,N_1067,N_1837);
and U2608 (N_2608,N_1812,N_1612);
and U2609 (N_2609,N_1740,N_1119);
nand U2610 (N_2610,N_1722,N_1021);
and U2611 (N_2611,N_1128,N_1901);
nor U2612 (N_2612,N_1626,N_1194);
or U2613 (N_2613,N_1392,N_1540);
and U2614 (N_2614,N_1831,N_1343);
and U2615 (N_2615,N_1703,N_1089);
or U2616 (N_2616,N_1137,N_1569);
and U2617 (N_2617,N_1702,N_1040);
nand U2618 (N_2618,N_1659,N_1019);
nor U2619 (N_2619,N_1703,N_1595);
and U2620 (N_2620,N_1703,N_1850);
or U2621 (N_2621,N_1389,N_1656);
nor U2622 (N_2622,N_1330,N_1965);
and U2623 (N_2623,N_1478,N_1865);
nand U2624 (N_2624,N_1855,N_1860);
and U2625 (N_2625,N_1901,N_1501);
or U2626 (N_2626,N_1183,N_1581);
nand U2627 (N_2627,N_1217,N_1596);
nor U2628 (N_2628,N_1224,N_1404);
nor U2629 (N_2629,N_1349,N_1273);
nand U2630 (N_2630,N_1139,N_1435);
and U2631 (N_2631,N_1421,N_1935);
nand U2632 (N_2632,N_1169,N_1059);
and U2633 (N_2633,N_1086,N_1728);
nor U2634 (N_2634,N_1027,N_1124);
nand U2635 (N_2635,N_1747,N_1207);
and U2636 (N_2636,N_1758,N_1196);
nand U2637 (N_2637,N_1278,N_1842);
nand U2638 (N_2638,N_1488,N_1476);
nand U2639 (N_2639,N_1400,N_1315);
and U2640 (N_2640,N_1432,N_1876);
or U2641 (N_2641,N_1992,N_1923);
and U2642 (N_2642,N_1065,N_1149);
or U2643 (N_2643,N_1885,N_1915);
and U2644 (N_2644,N_1587,N_1449);
and U2645 (N_2645,N_1972,N_1534);
nor U2646 (N_2646,N_1602,N_1311);
nand U2647 (N_2647,N_1234,N_1034);
or U2648 (N_2648,N_1802,N_1675);
and U2649 (N_2649,N_1376,N_1388);
and U2650 (N_2650,N_1547,N_1424);
nor U2651 (N_2651,N_1215,N_1735);
nor U2652 (N_2652,N_1601,N_1270);
or U2653 (N_2653,N_1615,N_1660);
and U2654 (N_2654,N_1237,N_1020);
nor U2655 (N_2655,N_1590,N_1957);
or U2656 (N_2656,N_1829,N_1283);
nand U2657 (N_2657,N_1357,N_1052);
and U2658 (N_2658,N_1772,N_1789);
nand U2659 (N_2659,N_1030,N_1584);
nand U2660 (N_2660,N_1157,N_1250);
or U2661 (N_2661,N_1207,N_1084);
or U2662 (N_2662,N_1751,N_1514);
nor U2663 (N_2663,N_1052,N_1381);
nand U2664 (N_2664,N_1721,N_1831);
or U2665 (N_2665,N_1935,N_1024);
or U2666 (N_2666,N_1669,N_1271);
and U2667 (N_2667,N_1320,N_1011);
and U2668 (N_2668,N_1474,N_1479);
nand U2669 (N_2669,N_1813,N_1765);
nor U2670 (N_2670,N_1277,N_1991);
nand U2671 (N_2671,N_1388,N_1851);
nor U2672 (N_2672,N_1422,N_1863);
nor U2673 (N_2673,N_1191,N_1991);
nor U2674 (N_2674,N_1171,N_1470);
nand U2675 (N_2675,N_1056,N_1417);
and U2676 (N_2676,N_1981,N_1600);
nand U2677 (N_2677,N_1594,N_1091);
nor U2678 (N_2678,N_1380,N_1706);
and U2679 (N_2679,N_1132,N_1054);
nor U2680 (N_2680,N_1924,N_1805);
nor U2681 (N_2681,N_1112,N_1457);
and U2682 (N_2682,N_1504,N_1529);
and U2683 (N_2683,N_1802,N_1760);
nand U2684 (N_2684,N_1921,N_1837);
nor U2685 (N_2685,N_1943,N_1152);
nor U2686 (N_2686,N_1018,N_1388);
or U2687 (N_2687,N_1384,N_1357);
and U2688 (N_2688,N_1247,N_1988);
nand U2689 (N_2689,N_1343,N_1999);
nor U2690 (N_2690,N_1808,N_1381);
nor U2691 (N_2691,N_1538,N_1598);
nand U2692 (N_2692,N_1691,N_1590);
and U2693 (N_2693,N_1066,N_1507);
and U2694 (N_2694,N_1199,N_1055);
nand U2695 (N_2695,N_1280,N_1771);
or U2696 (N_2696,N_1669,N_1280);
nor U2697 (N_2697,N_1037,N_1237);
nand U2698 (N_2698,N_1870,N_1314);
or U2699 (N_2699,N_1615,N_1585);
or U2700 (N_2700,N_1282,N_1878);
nand U2701 (N_2701,N_1345,N_1146);
nor U2702 (N_2702,N_1892,N_1645);
nor U2703 (N_2703,N_1109,N_1722);
nor U2704 (N_2704,N_1133,N_1001);
nor U2705 (N_2705,N_1834,N_1372);
nand U2706 (N_2706,N_1794,N_1851);
or U2707 (N_2707,N_1159,N_1005);
nor U2708 (N_2708,N_1099,N_1104);
nor U2709 (N_2709,N_1799,N_1572);
nand U2710 (N_2710,N_1215,N_1253);
or U2711 (N_2711,N_1856,N_1209);
nand U2712 (N_2712,N_1744,N_1965);
and U2713 (N_2713,N_1106,N_1147);
nand U2714 (N_2714,N_1807,N_1708);
and U2715 (N_2715,N_1610,N_1150);
nor U2716 (N_2716,N_1534,N_1570);
or U2717 (N_2717,N_1669,N_1916);
nand U2718 (N_2718,N_1059,N_1461);
nand U2719 (N_2719,N_1792,N_1491);
nor U2720 (N_2720,N_1865,N_1011);
and U2721 (N_2721,N_1985,N_1057);
and U2722 (N_2722,N_1053,N_1604);
nand U2723 (N_2723,N_1149,N_1324);
nand U2724 (N_2724,N_1150,N_1323);
nand U2725 (N_2725,N_1914,N_1566);
nand U2726 (N_2726,N_1864,N_1134);
nand U2727 (N_2727,N_1426,N_1438);
nor U2728 (N_2728,N_1760,N_1693);
and U2729 (N_2729,N_1046,N_1075);
nand U2730 (N_2730,N_1553,N_1051);
or U2731 (N_2731,N_1828,N_1877);
or U2732 (N_2732,N_1042,N_1358);
and U2733 (N_2733,N_1892,N_1924);
xor U2734 (N_2734,N_1343,N_1032);
nor U2735 (N_2735,N_1750,N_1483);
and U2736 (N_2736,N_1434,N_1288);
or U2737 (N_2737,N_1633,N_1201);
nand U2738 (N_2738,N_1706,N_1807);
nand U2739 (N_2739,N_1711,N_1745);
xor U2740 (N_2740,N_1674,N_1158);
nand U2741 (N_2741,N_1733,N_1443);
or U2742 (N_2742,N_1359,N_1808);
nand U2743 (N_2743,N_1555,N_1305);
nor U2744 (N_2744,N_1003,N_1706);
nand U2745 (N_2745,N_1158,N_1118);
and U2746 (N_2746,N_1705,N_1596);
and U2747 (N_2747,N_1562,N_1666);
nor U2748 (N_2748,N_1294,N_1863);
and U2749 (N_2749,N_1661,N_1605);
and U2750 (N_2750,N_1088,N_1647);
and U2751 (N_2751,N_1681,N_1316);
nor U2752 (N_2752,N_1293,N_1208);
nand U2753 (N_2753,N_1508,N_1502);
and U2754 (N_2754,N_1380,N_1294);
and U2755 (N_2755,N_1218,N_1386);
and U2756 (N_2756,N_1969,N_1904);
nor U2757 (N_2757,N_1297,N_1922);
nand U2758 (N_2758,N_1242,N_1587);
and U2759 (N_2759,N_1145,N_1407);
or U2760 (N_2760,N_1307,N_1846);
and U2761 (N_2761,N_1053,N_1656);
and U2762 (N_2762,N_1659,N_1314);
nor U2763 (N_2763,N_1639,N_1134);
or U2764 (N_2764,N_1225,N_1447);
nor U2765 (N_2765,N_1548,N_1713);
xor U2766 (N_2766,N_1264,N_1443);
and U2767 (N_2767,N_1969,N_1559);
or U2768 (N_2768,N_1642,N_1350);
nand U2769 (N_2769,N_1478,N_1212);
or U2770 (N_2770,N_1109,N_1071);
nor U2771 (N_2771,N_1400,N_1568);
nor U2772 (N_2772,N_1563,N_1804);
nor U2773 (N_2773,N_1215,N_1047);
and U2774 (N_2774,N_1630,N_1236);
nand U2775 (N_2775,N_1164,N_1038);
or U2776 (N_2776,N_1548,N_1959);
nor U2777 (N_2777,N_1832,N_1397);
or U2778 (N_2778,N_1862,N_1257);
and U2779 (N_2779,N_1394,N_1737);
nor U2780 (N_2780,N_1518,N_1900);
nor U2781 (N_2781,N_1766,N_1633);
nor U2782 (N_2782,N_1310,N_1732);
or U2783 (N_2783,N_1910,N_1026);
nand U2784 (N_2784,N_1518,N_1547);
nand U2785 (N_2785,N_1753,N_1602);
nor U2786 (N_2786,N_1165,N_1783);
or U2787 (N_2787,N_1012,N_1165);
nand U2788 (N_2788,N_1362,N_1998);
nand U2789 (N_2789,N_1891,N_1567);
nand U2790 (N_2790,N_1340,N_1193);
and U2791 (N_2791,N_1803,N_1463);
nand U2792 (N_2792,N_1257,N_1485);
and U2793 (N_2793,N_1113,N_1594);
nor U2794 (N_2794,N_1911,N_1072);
nand U2795 (N_2795,N_1243,N_1785);
or U2796 (N_2796,N_1873,N_1560);
or U2797 (N_2797,N_1982,N_1955);
or U2798 (N_2798,N_1567,N_1352);
or U2799 (N_2799,N_1635,N_1129);
and U2800 (N_2800,N_1692,N_1246);
and U2801 (N_2801,N_1382,N_1049);
or U2802 (N_2802,N_1599,N_1430);
nor U2803 (N_2803,N_1093,N_1915);
or U2804 (N_2804,N_1188,N_1082);
nand U2805 (N_2805,N_1298,N_1194);
or U2806 (N_2806,N_1355,N_1856);
nand U2807 (N_2807,N_1431,N_1627);
or U2808 (N_2808,N_1203,N_1192);
nor U2809 (N_2809,N_1822,N_1916);
and U2810 (N_2810,N_1604,N_1838);
or U2811 (N_2811,N_1468,N_1891);
and U2812 (N_2812,N_1988,N_1010);
nand U2813 (N_2813,N_1468,N_1108);
and U2814 (N_2814,N_1446,N_1898);
or U2815 (N_2815,N_1902,N_1092);
nor U2816 (N_2816,N_1561,N_1669);
or U2817 (N_2817,N_1203,N_1467);
nor U2818 (N_2818,N_1198,N_1342);
and U2819 (N_2819,N_1631,N_1612);
nand U2820 (N_2820,N_1735,N_1892);
nor U2821 (N_2821,N_1969,N_1800);
nor U2822 (N_2822,N_1007,N_1270);
nand U2823 (N_2823,N_1718,N_1296);
nand U2824 (N_2824,N_1333,N_1476);
nor U2825 (N_2825,N_1328,N_1099);
nand U2826 (N_2826,N_1942,N_1314);
and U2827 (N_2827,N_1797,N_1961);
and U2828 (N_2828,N_1239,N_1048);
xor U2829 (N_2829,N_1139,N_1127);
and U2830 (N_2830,N_1256,N_1515);
or U2831 (N_2831,N_1492,N_1602);
or U2832 (N_2832,N_1361,N_1287);
and U2833 (N_2833,N_1000,N_1397);
nand U2834 (N_2834,N_1272,N_1519);
or U2835 (N_2835,N_1613,N_1063);
nor U2836 (N_2836,N_1889,N_1651);
nand U2837 (N_2837,N_1162,N_1070);
and U2838 (N_2838,N_1134,N_1455);
or U2839 (N_2839,N_1744,N_1019);
nor U2840 (N_2840,N_1319,N_1468);
and U2841 (N_2841,N_1171,N_1526);
nor U2842 (N_2842,N_1289,N_1496);
nor U2843 (N_2843,N_1873,N_1738);
and U2844 (N_2844,N_1924,N_1755);
and U2845 (N_2845,N_1126,N_1950);
nand U2846 (N_2846,N_1263,N_1706);
or U2847 (N_2847,N_1290,N_1959);
nand U2848 (N_2848,N_1779,N_1132);
nor U2849 (N_2849,N_1036,N_1773);
or U2850 (N_2850,N_1053,N_1996);
nor U2851 (N_2851,N_1371,N_1287);
nand U2852 (N_2852,N_1189,N_1521);
nor U2853 (N_2853,N_1642,N_1327);
or U2854 (N_2854,N_1839,N_1131);
nor U2855 (N_2855,N_1474,N_1686);
or U2856 (N_2856,N_1895,N_1073);
and U2857 (N_2857,N_1152,N_1905);
nor U2858 (N_2858,N_1545,N_1527);
nand U2859 (N_2859,N_1400,N_1254);
or U2860 (N_2860,N_1785,N_1982);
nor U2861 (N_2861,N_1438,N_1229);
nor U2862 (N_2862,N_1918,N_1167);
xnor U2863 (N_2863,N_1441,N_1590);
nor U2864 (N_2864,N_1714,N_1105);
or U2865 (N_2865,N_1508,N_1980);
or U2866 (N_2866,N_1828,N_1057);
nand U2867 (N_2867,N_1093,N_1601);
nand U2868 (N_2868,N_1351,N_1855);
nor U2869 (N_2869,N_1402,N_1578);
nand U2870 (N_2870,N_1495,N_1761);
nor U2871 (N_2871,N_1631,N_1031);
or U2872 (N_2872,N_1323,N_1598);
and U2873 (N_2873,N_1830,N_1459);
and U2874 (N_2874,N_1645,N_1751);
nor U2875 (N_2875,N_1767,N_1367);
nor U2876 (N_2876,N_1729,N_1485);
or U2877 (N_2877,N_1323,N_1837);
nor U2878 (N_2878,N_1946,N_1024);
nand U2879 (N_2879,N_1648,N_1261);
nor U2880 (N_2880,N_1881,N_1808);
nor U2881 (N_2881,N_1730,N_1480);
nor U2882 (N_2882,N_1706,N_1262);
nand U2883 (N_2883,N_1656,N_1566);
nor U2884 (N_2884,N_1314,N_1099);
nor U2885 (N_2885,N_1429,N_1590);
nor U2886 (N_2886,N_1024,N_1767);
nor U2887 (N_2887,N_1977,N_1766);
nand U2888 (N_2888,N_1180,N_1398);
and U2889 (N_2889,N_1370,N_1780);
or U2890 (N_2890,N_1329,N_1000);
and U2891 (N_2891,N_1098,N_1737);
or U2892 (N_2892,N_1371,N_1805);
xnor U2893 (N_2893,N_1471,N_1582);
nand U2894 (N_2894,N_1119,N_1090);
nand U2895 (N_2895,N_1323,N_1588);
and U2896 (N_2896,N_1019,N_1562);
nor U2897 (N_2897,N_1856,N_1352);
nand U2898 (N_2898,N_1233,N_1422);
nand U2899 (N_2899,N_1582,N_1038);
and U2900 (N_2900,N_1973,N_1670);
nand U2901 (N_2901,N_1258,N_1335);
or U2902 (N_2902,N_1392,N_1846);
or U2903 (N_2903,N_1422,N_1600);
nand U2904 (N_2904,N_1797,N_1935);
and U2905 (N_2905,N_1744,N_1282);
nor U2906 (N_2906,N_1615,N_1624);
or U2907 (N_2907,N_1650,N_1027);
or U2908 (N_2908,N_1059,N_1093);
nor U2909 (N_2909,N_1194,N_1993);
and U2910 (N_2910,N_1207,N_1924);
nand U2911 (N_2911,N_1485,N_1934);
or U2912 (N_2912,N_1053,N_1738);
nand U2913 (N_2913,N_1268,N_1973);
and U2914 (N_2914,N_1096,N_1505);
or U2915 (N_2915,N_1044,N_1494);
nand U2916 (N_2916,N_1669,N_1737);
or U2917 (N_2917,N_1390,N_1212);
or U2918 (N_2918,N_1042,N_1272);
or U2919 (N_2919,N_1739,N_1794);
and U2920 (N_2920,N_1456,N_1610);
nand U2921 (N_2921,N_1873,N_1590);
nand U2922 (N_2922,N_1274,N_1208);
xor U2923 (N_2923,N_1916,N_1825);
or U2924 (N_2924,N_1769,N_1961);
nand U2925 (N_2925,N_1079,N_1547);
nor U2926 (N_2926,N_1434,N_1989);
or U2927 (N_2927,N_1678,N_1956);
nand U2928 (N_2928,N_1396,N_1473);
nor U2929 (N_2929,N_1939,N_1521);
or U2930 (N_2930,N_1833,N_1644);
and U2931 (N_2931,N_1475,N_1703);
and U2932 (N_2932,N_1592,N_1822);
nor U2933 (N_2933,N_1543,N_1696);
and U2934 (N_2934,N_1919,N_1963);
nand U2935 (N_2935,N_1464,N_1456);
and U2936 (N_2936,N_1989,N_1765);
nor U2937 (N_2937,N_1323,N_1001);
or U2938 (N_2938,N_1107,N_1132);
and U2939 (N_2939,N_1479,N_1569);
and U2940 (N_2940,N_1395,N_1189);
or U2941 (N_2941,N_1207,N_1653);
nor U2942 (N_2942,N_1486,N_1109);
or U2943 (N_2943,N_1507,N_1135);
nor U2944 (N_2944,N_1822,N_1750);
and U2945 (N_2945,N_1059,N_1668);
or U2946 (N_2946,N_1031,N_1796);
nand U2947 (N_2947,N_1956,N_1135);
or U2948 (N_2948,N_1507,N_1549);
nor U2949 (N_2949,N_1545,N_1981);
and U2950 (N_2950,N_1909,N_1672);
or U2951 (N_2951,N_1677,N_1405);
nand U2952 (N_2952,N_1704,N_1613);
nand U2953 (N_2953,N_1130,N_1652);
or U2954 (N_2954,N_1303,N_1538);
and U2955 (N_2955,N_1187,N_1729);
nand U2956 (N_2956,N_1977,N_1098);
and U2957 (N_2957,N_1614,N_1435);
nor U2958 (N_2958,N_1402,N_1571);
and U2959 (N_2959,N_1059,N_1466);
or U2960 (N_2960,N_1253,N_1042);
or U2961 (N_2961,N_1752,N_1206);
or U2962 (N_2962,N_1872,N_1194);
or U2963 (N_2963,N_1524,N_1173);
and U2964 (N_2964,N_1978,N_1401);
nand U2965 (N_2965,N_1337,N_1715);
nor U2966 (N_2966,N_1925,N_1289);
nor U2967 (N_2967,N_1720,N_1155);
or U2968 (N_2968,N_1576,N_1724);
or U2969 (N_2969,N_1022,N_1664);
or U2970 (N_2970,N_1070,N_1235);
and U2971 (N_2971,N_1181,N_1072);
nor U2972 (N_2972,N_1117,N_1381);
and U2973 (N_2973,N_1090,N_1347);
and U2974 (N_2974,N_1498,N_1075);
or U2975 (N_2975,N_1886,N_1827);
and U2976 (N_2976,N_1075,N_1982);
nand U2977 (N_2977,N_1992,N_1707);
and U2978 (N_2978,N_1124,N_1223);
and U2979 (N_2979,N_1728,N_1638);
nand U2980 (N_2980,N_1080,N_1094);
and U2981 (N_2981,N_1971,N_1375);
and U2982 (N_2982,N_1555,N_1522);
nand U2983 (N_2983,N_1031,N_1299);
nor U2984 (N_2984,N_1024,N_1047);
or U2985 (N_2985,N_1730,N_1064);
nor U2986 (N_2986,N_1462,N_1273);
or U2987 (N_2987,N_1021,N_1511);
or U2988 (N_2988,N_1239,N_1322);
nor U2989 (N_2989,N_1862,N_1554);
or U2990 (N_2990,N_1393,N_1485);
and U2991 (N_2991,N_1607,N_1283);
nor U2992 (N_2992,N_1775,N_1166);
nand U2993 (N_2993,N_1559,N_1198);
nor U2994 (N_2994,N_1095,N_1899);
or U2995 (N_2995,N_1741,N_1185);
and U2996 (N_2996,N_1727,N_1545);
nor U2997 (N_2997,N_1731,N_1996);
or U2998 (N_2998,N_1102,N_1809);
nand U2999 (N_2999,N_1793,N_1375);
nand U3000 (N_3000,N_2921,N_2509);
or U3001 (N_3001,N_2021,N_2725);
and U3002 (N_3002,N_2825,N_2307);
or U3003 (N_3003,N_2263,N_2269);
nor U3004 (N_3004,N_2848,N_2150);
nor U3005 (N_3005,N_2650,N_2272);
nand U3006 (N_3006,N_2333,N_2931);
nor U3007 (N_3007,N_2399,N_2197);
and U3008 (N_3008,N_2194,N_2732);
nor U3009 (N_3009,N_2506,N_2571);
nand U3010 (N_3010,N_2053,N_2047);
nand U3011 (N_3011,N_2028,N_2225);
and U3012 (N_3012,N_2934,N_2964);
and U3013 (N_3013,N_2359,N_2039);
and U3014 (N_3014,N_2956,N_2790);
nor U3015 (N_3015,N_2688,N_2190);
or U3016 (N_3016,N_2629,N_2530);
and U3017 (N_3017,N_2349,N_2829);
nor U3018 (N_3018,N_2670,N_2497);
and U3019 (N_3019,N_2122,N_2946);
and U3020 (N_3020,N_2974,N_2920);
or U3021 (N_3021,N_2412,N_2116);
or U3022 (N_3022,N_2246,N_2797);
nor U3023 (N_3023,N_2351,N_2988);
nor U3024 (N_3024,N_2483,N_2198);
and U3025 (N_3025,N_2250,N_2710);
or U3026 (N_3026,N_2409,N_2214);
nand U3027 (N_3027,N_2299,N_2220);
nor U3028 (N_3028,N_2281,N_2109);
or U3029 (N_3029,N_2885,N_2646);
and U3030 (N_3030,N_2756,N_2437);
or U3031 (N_3031,N_2998,N_2906);
and U3032 (N_3032,N_2827,N_2100);
and U3033 (N_3033,N_2037,N_2556);
and U3034 (N_3034,N_2619,N_2199);
and U3035 (N_3035,N_2529,N_2522);
nor U3036 (N_3036,N_2467,N_2612);
and U3037 (N_3037,N_2961,N_2420);
and U3038 (N_3038,N_2962,N_2933);
and U3039 (N_3039,N_2006,N_2130);
nand U3040 (N_3040,N_2842,N_2032);
nand U3041 (N_3041,N_2415,N_2490);
or U3042 (N_3042,N_2864,N_2027);
nor U3043 (N_3043,N_2751,N_2630);
and U3044 (N_3044,N_2652,N_2965);
or U3045 (N_3045,N_2381,N_2115);
and U3046 (N_3046,N_2915,N_2636);
and U3047 (N_3047,N_2748,N_2063);
or U3048 (N_3048,N_2777,N_2254);
nand U3049 (N_3049,N_2236,N_2152);
nor U3050 (N_3050,N_2749,N_2262);
nor U3051 (N_3051,N_2408,N_2248);
and U3052 (N_3052,N_2810,N_2304);
nor U3053 (N_3053,N_2653,N_2905);
or U3054 (N_3054,N_2091,N_2118);
nand U3055 (N_3055,N_2332,N_2428);
and U3056 (N_3056,N_2702,N_2955);
nor U3057 (N_3057,N_2193,N_2338);
nor U3058 (N_3058,N_2442,N_2891);
or U3059 (N_3059,N_2256,N_2231);
nor U3060 (N_3060,N_2999,N_2947);
or U3061 (N_3061,N_2243,N_2106);
and U3062 (N_3062,N_2648,N_2136);
nor U3063 (N_3063,N_2877,N_2580);
and U3064 (N_3064,N_2685,N_2210);
or U3065 (N_3065,N_2012,N_2561);
nor U3066 (N_3066,N_2681,N_2387);
or U3067 (N_3067,N_2835,N_2633);
nor U3068 (N_3068,N_2696,N_2910);
and U3069 (N_3069,N_2919,N_2523);
nor U3070 (N_3070,N_2493,N_2200);
or U3071 (N_3071,N_2083,N_2609);
and U3072 (N_3072,N_2585,N_2917);
and U3073 (N_3073,N_2794,N_2870);
nor U3074 (N_3074,N_2557,N_2061);
nor U3075 (N_3075,N_2867,N_2623);
or U3076 (N_3076,N_2142,N_2881);
nand U3077 (N_3077,N_2573,N_2785);
nand U3078 (N_3078,N_2948,N_2520);
nor U3079 (N_3079,N_2731,N_2882);
nand U3080 (N_3080,N_2977,N_2172);
nand U3081 (N_3081,N_2570,N_2085);
nand U3082 (N_3082,N_2103,N_2291);
nor U3083 (N_3083,N_2496,N_2798);
nand U3084 (N_3084,N_2218,N_2383);
and U3085 (N_3085,N_2659,N_2159);
nand U3086 (N_3086,N_2701,N_2903);
or U3087 (N_3087,N_2153,N_2958);
and U3088 (N_3088,N_2241,N_2158);
nor U3089 (N_3089,N_2562,N_2382);
nand U3090 (N_3090,N_2173,N_2235);
nand U3091 (N_3091,N_2292,N_2872);
and U3092 (N_3092,N_2188,N_2875);
nor U3093 (N_3093,N_2936,N_2823);
and U3094 (N_3094,N_2967,N_2238);
or U3095 (N_3095,N_2993,N_2795);
nor U3096 (N_3096,N_2691,N_2591);
or U3097 (N_3097,N_2322,N_2449);
nand U3098 (N_3098,N_2501,N_2365);
and U3099 (N_3099,N_2282,N_2357);
nor U3100 (N_3100,N_2995,N_2097);
nand U3101 (N_3101,N_2337,N_2957);
nor U3102 (N_3102,N_2900,N_2041);
and U3103 (N_3103,N_2505,N_2229);
or U3104 (N_3104,N_2760,N_2727);
or U3105 (N_3105,N_2963,N_2985);
nor U3106 (N_3106,N_2853,N_2156);
nor U3107 (N_3107,N_2287,N_2930);
nand U3108 (N_3108,N_2604,N_2233);
nor U3109 (N_3109,N_2464,N_2558);
or U3110 (N_3110,N_2356,N_2026);
nor U3111 (N_3111,N_2471,N_2617);
and U3112 (N_3112,N_2576,N_2801);
nor U3113 (N_3113,N_2997,N_2878);
and U3114 (N_3114,N_2073,N_2697);
and U3115 (N_3115,N_2279,N_2347);
and U3116 (N_3116,N_2439,N_2462);
nand U3117 (N_3117,N_2384,N_2452);
and U3118 (N_3118,N_2326,N_2285);
and U3119 (N_3119,N_2622,N_2743);
nand U3120 (N_3120,N_2703,N_2278);
nand U3121 (N_3121,N_2478,N_2966);
and U3122 (N_3122,N_2157,N_2082);
nand U3123 (N_3123,N_2839,N_2475);
or U3124 (N_3124,N_2911,N_2215);
and U3125 (N_3125,N_2232,N_2127);
and U3126 (N_3126,N_2178,N_2302);
nand U3127 (N_3127,N_2513,N_2717);
and U3128 (N_3128,N_2160,N_2042);
and U3129 (N_3129,N_2539,N_2773);
and U3130 (N_3130,N_2744,N_2613);
nand U3131 (N_3131,N_2857,N_2016);
or U3132 (N_3132,N_2597,N_2112);
nor U3133 (N_3133,N_2972,N_2588);
nand U3134 (N_3134,N_2147,N_2712);
or U3135 (N_3135,N_2267,N_2336);
nor U3136 (N_3136,N_2371,N_2473);
or U3137 (N_3137,N_2874,N_2472);
or U3138 (N_3138,N_2540,N_2444);
and U3139 (N_3139,N_2148,N_2805);
or U3140 (N_3140,N_2058,N_2252);
or U3141 (N_3141,N_2763,N_2455);
or U3142 (N_3142,N_2072,N_2960);
and U3143 (N_3143,N_2192,N_2895);
or U3144 (N_3144,N_2799,N_2355);
nand U3145 (N_3145,N_2525,N_2901);
and U3146 (N_3146,N_2672,N_2907);
nand U3147 (N_3147,N_2855,N_2312);
and U3148 (N_3148,N_2404,N_2902);
and U3149 (N_3149,N_2802,N_2854);
or U3150 (N_3150,N_2459,N_2055);
or U3151 (N_3151,N_2768,N_2542);
and U3152 (N_3152,N_2577,N_2364);
or U3153 (N_3153,N_2244,N_2013);
nand U3154 (N_3154,N_2837,N_2165);
or U3155 (N_3155,N_2692,N_2675);
or U3156 (N_3156,N_2821,N_2264);
nor U3157 (N_3157,N_2660,N_2319);
nor U3158 (N_3158,N_2943,N_2203);
nor U3159 (N_3159,N_2488,N_2954);
nand U3160 (N_3160,N_2071,N_2929);
nand U3161 (N_3161,N_2549,N_2020);
or U3162 (N_3162,N_2531,N_2888);
and U3163 (N_3163,N_2873,N_2078);
nor U3164 (N_3164,N_2563,N_2677);
or U3165 (N_3165,N_2125,N_2694);
nand U3166 (N_3166,N_2851,N_2313);
nor U3167 (N_3167,N_2368,N_2753);
or U3168 (N_3168,N_2145,N_2253);
or U3169 (N_3169,N_2626,N_2879);
nand U3170 (N_3170,N_2693,N_2024);
and U3171 (N_3171,N_2524,N_2820);
or U3172 (N_3172,N_2782,N_2804);
and U3173 (N_3173,N_2275,N_2300);
and U3174 (N_3174,N_2031,N_2186);
nor U3175 (N_3175,N_2819,N_2719);
nand U3176 (N_3176,N_2240,N_2335);
and U3177 (N_3177,N_2952,N_2423);
or U3178 (N_3178,N_2087,N_2162);
or U3179 (N_3179,N_2003,N_2987);
nor U3180 (N_3180,N_2639,N_2228);
or U3181 (N_3181,N_2137,N_2057);
nor U3182 (N_3182,N_2863,N_2611);
or U3183 (N_3183,N_2463,N_2434);
nor U3184 (N_3184,N_2069,N_2308);
nor U3185 (N_3185,N_2414,N_2504);
or U3186 (N_3186,N_2447,N_2108);
and U3187 (N_3187,N_2352,N_2126);
or U3188 (N_3188,N_2117,N_2286);
nor U3189 (N_3189,N_2986,N_2034);
nor U3190 (N_3190,N_2984,N_2981);
or U3191 (N_3191,N_2537,N_2724);
nor U3192 (N_3192,N_2080,N_2551);
xor U3193 (N_3193,N_2209,N_2315);
nand U3194 (N_3194,N_2655,N_2750);
or U3195 (N_3195,N_2913,N_2051);
and U3196 (N_3196,N_2800,N_2305);
nor U3197 (N_3197,N_2765,N_2594);
and U3198 (N_3198,N_2486,N_2323);
nor U3199 (N_3199,N_2832,N_2762);
nand U3200 (N_3200,N_2219,N_2916);
and U3201 (N_3201,N_2926,N_2280);
nor U3202 (N_3202,N_2969,N_2747);
and U3203 (N_3203,N_2084,N_2850);
nor U3204 (N_3204,N_2043,N_2124);
and U3205 (N_3205,N_2318,N_2195);
or U3206 (N_3206,N_2840,N_2081);
and U3207 (N_3207,N_2251,N_2339);
nand U3208 (N_3208,N_2089,N_2369);
and U3209 (N_3209,N_2861,N_2757);
nand U3210 (N_3210,N_2179,N_2389);
or U3211 (N_3211,N_2038,N_2184);
nor U3212 (N_3212,N_2858,N_2425);
nand U3213 (N_3213,N_2424,N_2699);
nor U3214 (N_3214,N_2975,N_2092);
nor U3215 (N_3215,N_2255,N_2481);
nand U3216 (N_3216,N_2128,N_2469);
nor U3217 (N_3217,N_2945,N_2880);
xor U3218 (N_3218,N_2884,N_2499);
or U3219 (N_3219,N_2990,N_2546);
nand U3220 (N_3220,N_2970,N_2890);
and U3221 (N_3221,N_2064,N_2163);
or U3222 (N_3222,N_2535,N_2706);
and U3223 (N_3223,N_2457,N_2651);
nand U3224 (N_3224,N_2859,N_2018);
nand U3225 (N_3225,N_2908,N_2207);
or U3226 (N_3226,N_2213,N_2134);
and U3227 (N_3227,N_2758,N_2949);
and U3228 (N_3228,N_2470,N_2010);
nor U3229 (N_3229,N_2616,N_2040);
or U3230 (N_3230,N_2224,N_2528);
and U3231 (N_3231,N_2796,N_2932);
or U3232 (N_3232,N_2569,N_2595);
nand U3233 (N_3233,N_2397,N_2909);
nand U3234 (N_3234,N_2321,N_2599);
nand U3235 (N_3235,N_2270,N_2979);
or U3236 (N_3236,N_2690,N_2781);
nand U3237 (N_3237,N_2632,N_2568);
and U3238 (N_3238,N_2477,N_2410);
and U3239 (N_3239,N_2713,N_2334);
or U3240 (N_3240,N_2367,N_2489);
nand U3241 (N_3241,N_2893,N_2432);
or U3242 (N_3242,N_2771,N_2366);
nand U3243 (N_3243,N_2788,N_2474);
or U3244 (N_3244,N_2258,N_2348);
nand U3245 (N_3245,N_2944,N_2327);
or U3246 (N_3246,N_2564,N_2803);
and U3247 (N_3247,N_2450,N_2146);
or U3248 (N_3248,N_2754,N_2941);
or U3249 (N_3249,N_2283,N_2668);
nand U3250 (N_3250,N_2191,N_2086);
nand U3251 (N_3251,N_2306,N_2548);
or U3252 (N_3252,N_2868,N_2579);
nor U3253 (N_3253,N_2606,N_2590);
and U3254 (N_3254,N_2787,N_2761);
nor U3255 (N_3255,N_2683,N_2634);
and U3256 (N_3256,N_2353,N_2733);
nor U3257 (N_3257,N_2290,N_2922);
nand U3258 (N_3258,N_2673,N_2614);
nor U3259 (N_3259,N_2316,N_2918);
nand U3260 (N_3260,N_2992,N_2608);
or U3261 (N_3261,N_2543,N_2716);
and U3262 (N_3262,N_2674,N_2996);
nand U3263 (N_3263,N_2741,N_2730);
nor U3264 (N_3264,N_2023,N_2793);
or U3265 (N_3265,N_2989,N_2645);
and U3266 (N_3266,N_2400,N_2422);
or U3267 (N_3267,N_2871,N_2119);
and U3268 (N_3268,N_2360,N_2418);
nor U3269 (N_3269,N_2401,N_2566);
or U3270 (N_3270,N_2700,N_2492);
or U3271 (N_3271,N_2638,N_2405);
nor U3272 (N_3272,N_2680,N_2887);
or U3273 (N_3273,N_2096,N_2904);
nand U3274 (N_3274,N_2860,N_2665);
and U3275 (N_3275,N_2077,N_2076);
or U3276 (N_3276,N_2170,N_2752);
nand U3277 (N_3277,N_2536,N_2094);
nand U3278 (N_3278,N_2216,N_2138);
xnor U3279 (N_3279,N_2598,N_2704);
xnor U3280 (N_3280,N_2155,N_2030);
nor U3281 (N_3281,N_2000,N_2324);
nand U3282 (N_3282,N_2066,N_2484);
and U3283 (N_3283,N_2206,N_2846);
and U3284 (N_3284,N_2586,N_2377);
nand U3285 (N_3285,N_2684,N_2005);
nor U3286 (N_3286,N_2249,N_2721);
nand U3287 (N_3287,N_2789,N_2247);
or U3288 (N_3288,N_2237,N_2779);
nand U3289 (N_3289,N_2547,N_2056);
nand U3290 (N_3290,N_2667,N_2132);
and U3291 (N_3291,N_2074,N_2011);
nand U3292 (N_3292,N_2971,N_2784);
nor U3293 (N_3293,N_2592,N_2661);
xnor U3294 (N_3294,N_2242,N_2664);
nand U3295 (N_3295,N_2705,N_2458);
or U3296 (N_3296,N_2847,N_2897);
and U3297 (N_3297,N_2627,N_2927);
nand U3298 (N_3298,N_2385,N_2806);
nand U3299 (N_3299,N_2643,N_2378);
nand U3300 (N_3300,N_2380,N_2445);
or U3301 (N_3301,N_2429,N_2105);
nor U3302 (N_3302,N_2375,N_2654);
nor U3303 (N_3303,N_2376,N_2487);
and U3304 (N_3304,N_2177,N_2642);
and U3305 (N_3305,N_2396,N_2894);
nand U3306 (N_3306,N_2766,N_2565);
nand U3307 (N_3307,N_2682,N_2476);
and U3308 (N_3308,N_2976,N_2968);
nor U3309 (N_3309,N_2658,N_2391);
or U3310 (N_3310,N_2303,N_2663);
nor U3311 (N_3311,N_2838,N_2245);
or U3312 (N_3312,N_2959,N_2494);
or U3313 (N_3313,N_2786,N_2541);
xnor U3314 (N_3314,N_2849,N_2273);
nor U3315 (N_3315,N_2676,N_2780);
nor U3316 (N_3316,N_2644,N_2774);
and U3317 (N_3317,N_2104,N_2002);
or U3318 (N_3318,N_2869,N_2048);
and U3319 (N_3319,N_2831,N_2886);
nor U3320 (N_3320,N_2394,N_2257);
and U3321 (N_3321,N_2809,N_2695);
and U3322 (N_3322,N_2271,N_2435);
nand U3323 (N_3323,N_2393,N_2346);
nand U3324 (N_3324,N_2482,N_2640);
and U3325 (N_3325,N_2552,N_2554);
nand U3326 (N_3326,N_2519,N_2413);
nand U3327 (N_3327,N_2709,N_2912);
nand U3328 (N_3328,N_2739,N_2102);
nand U3329 (N_3329,N_2465,N_2289);
and U3330 (N_3330,N_2161,N_2268);
or U3331 (N_3331,N_2411,N_2657);
and U3332 (N_3332,N_2807,N_2892);
nor U3333 (N_3333,N_2527,N_2631);
and U3334 (N_3334,N_2007,N_2582);
nand U3335 (N_3335,N_2154,N_2507);
or U3336 (N_3336,N_2764,N_2735);
or U3337 (N_3337,N_2711,N_2679);
and U3338 (N_3338,N_2274,N_2615);
and U3339 (N_3339,N_2973,N_2534);
nor U3340 (N_3340,N_2379,N_2852);
nor U3341 (N_3341,N_2828,N_2817);
or U3342 (N_3342,N_2440,N_2553);
and U3343 (N_3343,N_2044,N_2373);
or U3344 (N_3344,N_2196,N_2468);
and U3345 (N_3345,N_2398,N_2671);
nand U3346 (N_3346,N_2171,N_2433);
or U3347 (N_3347,N_2620,N_2362);
nand U3348 (N_3348,N_2426,N_2395);
or U3349 (N_3349,N_2637,N_2815);
or U3350 (N_3350,N_2386,N_2431);
nor U3351 (N_3351,N_2451,N_2180);
nand U3352 (N_3352,N_2816,N_2239);
and U3353 (N_3353,N_2980,N_2572);
or U3354 (N_3354,N_2792,N_2123);
or U3355 (N_3355,N_2578,N_2601);
nor U3356 (N_3356,N_2075,N_2830);
nand U3357 (N_3357,N_2009,N_2940);
nand U3358 (N_3358,N_2416,N_2361);
or U3359 (N_3359,N_2288,N_2480);
nand U3360 (N_3360,N_2978,N_2176);
nor U3361 (N_3361,N_2737,N_2350);
nor U3362 (N_3362,N_2707,N_2098);
and U3363 (N_3363,N_2625,N_2419);
or U3364 (N_3364,N_2298,N_2844);
and U3365 (N_3365,N_2149,N_2372);
or U3366 (N_3366,N_2341,N_2205);
nand U3367 (N_3367,N_2698,N_2441);
nor U3368 (N_3368,N_2746,N_2610);
nor U3369 (N_3369,N_2330,N_2456);
and U3370 (N_3370,N_2755,N_2515);
or U3371 (N_3371,N_2046,N_2508);
nand U3372 (N_3372,N_2769,N_2182);
nor U3373 (N_3373,N_2221,N_2928);
or U3374 (N_3374,N_2358,N_2814);
and U3375 (N_3375,N_2720,N_2421);
and U3376 (N_3376,N_2151,N_2924);
xor U3377 (N_3377,N_2417,N_2516);
nand U3378 (N_3378,N_2550,N_2059);
or U3379 (N_3379,N_2589,N_2669);
nand U3380 (N_3380,N_2320,N_2001);
and U3381 (N_3381,N_2718,N_2466);
xnor U3382 (N_3382,N_2185,N_2227);
nor U3383 (N_3383,N_2461,N_2994);
nor U3384 (N_3384,N_2628,N_2230);
or U3385 (N_3385,N_2222,N_2656);
nand U3386 (N_3386,N_2938,N_2596);
nor U3387 (N_3387,N_2354,N_2982);
nand U3388 (N_3388,N_2783,N_2204);
nand U3389 (N_3389,N_2942,N_2107);
nand U3390 (N_3390,N_2736,N_2343);
nand U3391 (N_3391,N_2164,N_2297);
or U3392 (N_3392,N_2953,N_2110);
or U3393 (N_3393,N_2485,N_2495);
or U3394 (N_3394,N_2544,N_2388);
and U3395 (N_3395,N_2175,N_2143);
nor U3396 (N_3396,N_2772,N_2402);
or U3397 (N_3397,N_2939,N_2647);
nor U3398 (N_3398,N_2454,N_2277);
or U3399 (N_3399,N_2131,N_2951);
or U3400 (N_3400,N_2723,N_2574);
or U3401 (N_3401,N_2033,N_2896);
nand U3402 (N_3402,N_2050,N_2935);
nand U3403 (N_3403,N_2166,N_2883);
and U3404 (N_3404,N_2070,N_2045);
and U3405 (N_3405,N_2641,N_2446);
or U3406 (N_3406,N_2301,N_2635);
and U3407 (N_3407,N_2062,N_2135);
and U3408 (N_3408,N_2845,N_2778);
and U3409 (N_3409,N_2088,N_2649);
or U3410 (N_3410,N_2726,N_2022);
xnor U3411 (N_3411,N_2407,N_2168);
or U3412 (N_3412,N_2602,N_2189);
nand U3413 (N_3413,N_2065,N_2004);
or U3414 (N_3414,N_2517,N_2114);
and U3415 (N_3415,N_2687,N_2511);
nand U3416 (N_3416,N_2775,N_2008);
nand U3417 (N_3417,N_2605,N_2510);
nor U3418 (N_3418,N_2049,N_2923);
nand U3419 (N_3419,N_2503,N_2403);
nor U3420 (N_3420,N_2406,N_2866);
nand U3421 (N_3421,N_2317,N_2448);
nor U3422 (N_3422,N_2822,N_2309);
nand U3423 (N_3423,N_2223,N_2438);
or U3424 (N_3424,N_2526,N_2502);
xor U3425 (N_3425,N_2791,N_2101);
nor U3426 (N_3426,N_2211,N_2689);
or U3427 (N_3427,N_2133,N_2841);
and U3428 (N_3428,N_2035,N_2618);
nand U3429 (N_3429,N_2460,N_2436);
nor U3430 (N_3430,N_2555,N_2090);
nor U3431 (N_3431,N_2276,N_2139);
nand U3432 (N_3432,N_2583,N_2093);
nor U3433 (N_3433,N_2311,N_2111);
and U3434 (N_3434,N_2714,N_2374);
and U3435 (N_3435,N_2603,N_2068);
or U3436 (N_3436,N_2036,N_2141);
xnor U3437 (N_3437,N_2167,N_2331);
nand U3438 (N_3438,N_2686,N_2812);
nor U3439 (N_3439,N_2261,N_2767);
or U3440 (N_3440,N_2843,N_2865);
nand U3441 (N_3441,N_2808,N_2325);
nand U3442 (N_3442,N_2824,N_2342);
nor U3443 (N_3443,N_2740,N_2293);
and U3444 (N_3444,N_2738,N_2836);
nand U3445 (N_3445,N_2226,N_2479);
nor U3446 (N_3446,N_2745,N_2587);
nor U3447 (N_3447,N_2925,N_2314);
nor U3448 (N_3448,N_2512,N_2060);
and U3449 (N_3449,N_2937,N_2734);
nand U3450 (N_3450,N_2532,N_2581);
or U3451 (N_3451,N_2329,N_2593);
nor U3452 (N_3452,N_2491,N_2140);
or U3453 (N_3453,N_2430,N_2328);
and U3454 (N_3454,N_2560,N_2174);
or U3455 (N_3455,N_2500,N_2518);
nor U3456 (N_3456,N_2834,N_2678);
and U3457 (N_3457,N_2183,N_2811);
or U3458 (N_3458,N_2538,N_2453);
and U3459 (N_3459,N_2559,N_2856);
nor U3460 (N_3460,N_2129,N_2521);
or U3461 (N_3461,N_2759,N_2095);
nand U3462 (N_3462,N_2427,N_2054);
and U3463 (N_3463,N_2624,N_2722);
nor U3464 (N_3464,N_2284,N_2019);
nand U3465 (N_3465,N_2545,N_2708);
and U3466 (N_3466,N_2370,N_2567);
nand U3467 (N_3467,N_2295,N_2607);
nand U3468 (N_3468,N_2120,N_2208);
or U3469 (N_3469,N_2344,N_2584);
nor U3470 (N_3470,N_2898,N_2212);
nand U3471 (N_3471,N_2294,N_2234);
nor U3472 (N_3472,N_2014,N_2169);
nor U3473 (N_3473,N_2296,N_2729);
xnor U3474 (N_3474,N_2121,N_2575);
nor U3475 (N_3475,N_2029,N_2265);
nand U3476 (N_3476,N_2025,N_2662);
nand U3477 (N_3477,N_2181,N_2363);
or U3478 (N_3478,N_2666,N_2187);
nor U3479 (N_3479,N_2345,N_2015);
and U3480 (N_3480,N_2728,N_2813);
and U3481 (N_3481,N_2833,N_2201);
nand U3482 (N_3482,N_2260,N_2113);
and U3483 (N_3483,N_2392,N_2621);
and U3484 (N_3484,N_2202,N_2144);
nand U3485 (N_3485,N_2266,N_2862);
and U3486 (N_3486,N_2217,N_2876);
nand U3487 (N_3487,N_2818,N_2310);
and U3488 (N_3488,N_2950,N_2340);
nand U3489 (N_3489,N_2259,N_2099);
nand U3490 (N_3490,N_2600,N_2533);
nor U3491 (N_3491,N_2826,N_2742);
and U3492 (N_3492,N_2770,N_2017);
nor U3493 (N_3493,N_2514,N_2991);
and U3494 (N_3494,N_2079,N_2914);
or U3495 (N_3495,N_2889,N_2983);
xor U3496 (N_3496,N_2899,N_2390);
nand U3497 (N_3497,N_2067,N_2715);
nand U3498 (N_3498,N_2776,N_2052);
and U3499 (N_3499,N_2498,N_2443);
nand U3500 (N_3500,N_2046,N_2318);
and U3501 (N_3501,N_2220,N_2509);
or U3502 (N_3502,N_2651,N_2145);
nand U3503 (N_3503,N_2629,N_2032);
and U3504 (N_3504,N_2801,N_2119);
nand U3505 (N_3505,N_2350,N_2316);
and U3506 (N_3506,N_2339,N_2302);
and U3507 (N_3507,N_2902,N_2292);
nor U3508 (N_3508,N_2817,N_2166);
nor U3509 (N_3509,N_2787,N_2757);
nand U3510 (N_3510,N_2164,N_2738);
nor U3511 (N_3511,N_2665,N_2788);
and U3512 (N_3512,N_2557,N_2080);
nor U3513 (N_3513,N_2520,N_2826);
nor U3514 (N_3514,N_2198,N_2099);
or U3515 (N_3515,N_2915,N_2740);
nand U3516 (N_3516,N_2254,N_2548);
or U3517 (N_3517,N_2538,N_2497);
and U3518 (N_3518,N_2365,N_2725);
and U3519 (N_3519,N_2916,N_2065);
nand U3520 (N_3520,N_2953,N_2178);
or U3521 (N_3521,N_2216,N_2286);
nand U3522 (N_3522,N_2573,N_2261);
nor U3523 (N_3523,N_2717,N_2249);
nor U3524 (N_3524,N_2477,N_2149);
nand U3525 (N_3525,N_2005,N_2639);
or U3526 (N_3526,N_2588,N_2140);
nand U3527 (N_3527,N_2350,N_2627);
or U3528 (N_3528,N_2238,N_2353);
and U3529 (N_3529,N_2071,N_2651);
nor U3530 (N_3530,N_2064,N_2383);
and U3531 (N_3531,N_2922,N_2676);
nor U3532 (N_3532,N_2016,N_2307);
and U3533 (N_3533,N_2239,N_2898);
nand U3534 (N_3534,N_2727,N_2273);
or U3535 (N_3535,N_2939,N_2598);
nand U3536 (N_3536,N_2942,N_2266);
and U3537 (N_3537,N_2030,N_2498);
nor U3538 (N_3538,N_2497,N_2205);
or U3539 (N_3539,N_2346,N_2208);
and U3540 (N_3540,N_2516,N_2876);
and U3541 (N_3541,N_2714,N_2882);
nand U3542 (N_3542,N_2987,N_2540);
or U3543 (N_3543,N_2152,N_2140);
nand U3544 (N_3544,N_2159,N_2543);
nand U3545 (N_3545,N_2360,N_2093);
nand U3546 (N_3546,N_2416,N_2499);
and U3547 (N_3547,N_2566,N_2190);
or U3548 (N_3548,N_2067,N_2163);
nand U3549 (N_3549,N_2601,N_2486);
nand U3550 (N_3550,N_2354,N_2348);
xor U3551 (N_3551,N_2450,N_2209);
or U3552 (N_3552,N_2550,N_2453);
nand U3553 (N_3553,N_2748,N_2918);
nor U3554 (N_3554,N_2984,N_2481);
nor U3555 (N_3555,N_2988,N_2569);
and U3556 (N_3556,N_2088,N_2650);
nor U3557 (N_3557,N_2110,N_2474);
nand U3558 (N_3558,N_2138,N_2207);
nor U3559 (N_3559,N_2504,N_2314);
nand U3560 (N_3560,N_2708,N_2006);
and U3561 (N_3561,N_2064,N_2761);
nor U3562 (N_3562,N_2932,N_2485);
nor U3563 (N_3563,N_2718,N_2569);
and U3564 (N_3564,N_2296,N_2255);
or U3565 (N_3565,N_2865,N_2404);
and U3566 (N_3566,N_2083,N_2464);
and U3567 (N_3567,N_2631,N_2010);
nor U3568 (N_3568,N_2570,N_2384);
and U3569 (N_3569,N_2551,N_2212);
and U3570 (N_3570,N_2039,N_2046);
nand U3571 (N_3571,N_2352,N_2372);
nand U3572 (N_3572,N_2121,N_2896);
and U3573 (N_3573,N_2027,N_2345);
or U3574 (N_3574,N_2736,N_2588);
nor U3575 (N_3575,N_2755,N_2454);
or U3576 (N_3576,N_2171,N_2220);
or U3577 (N_3577,N_2507,N_2661);
nand U3578 (N_3578,N_2553,N_2354);
and U3579 (N_3579,N_2761,N_2617);
or U3580 (N_3580,N_2345,N_2131);
or U3581 (N_3581,N_2833,N_2398);
and U3582 (N_3582,N_2659,N_2783);
and U3583 (N_3583,N_2141,N_2079);
and U3584 (N_3584,N_2068,N_2301);
nand U3585 (N_3585,N_2248,N_2494);
nand U3586 (N_3586,N_2622,N_2275);
or U3587 (N_3587,N_2528,N_2269);
and U3588 (N_3588,N_2405,N_2485);
and U3589 (N_3589,N_2525,N_2791);
or U3590 (N_3590,N_2743,N_2373);
and U3591 (N_3591,N_2775,N_2301);
nand U3592 (N_3592,N_2678,N_2045);
nor U3593 (N_3593,N_2774,N_2238);
nor U3594 (N_3594,N_2743,N_2884);
and U3595 (N_3595,N_2716,N_2179);
or U3596 (N_3596,N_2276,N_2503);
xnor U3597 (N_3597,N_2243,N_2747);
nand U3598 (N_3598,N_2901,N_2543);
or U3599 (N_3599,N_2773,N_2842);
or U3600 (N_3600,N_2745,N_2282);
nand U3601 (N_3601,N_2261,N_2586);
xnor U3602 (N_3602,N_2199,N_2162);
nand U3603 (N_3603,N_2299,N_2653);
nand U3604 (N_3604,N_2388,N_2810);
and U3605 (N_3605,N_2211,N_2069);
nand U3606 (N_3606,N_2011,N_2095);
and U3607 (N_3607,N_2114,N_2948);
and U3608 (N_3608,N_2243,N_2170);
nor U3609 (N_3609,N_2170,N_2910);
nor U3610 (N_3610,N_2327,N_2526);
and U3611 (N_3611,N_2656,N_2885);
and U3612 (N_3612,N_2645,N_2711);
or U3613 (N_3613,N_2521,N_2417);
and U3614 (N_3614,N_2514,N_2841);
nor U3615 (N_3615,N_2945,N_2658);
xor U3616 (N_3616,N_2249,N_2264);
and U3617 (N_3617,N_2941,N_2813);
nand U3618 (N_3618,N_2178,N_2673);
and U3619 (N_3619,N_2576,N_2159);
and U3620 (N_3620,N_2748,N_2009);
nand U3621 (N_3621,N_2684,N_2785);
or U3622 (N_3622,N_2985,N_2966);
and U3623 (N_3623,N_2617,N_2071);
nor U3624 (N_3624,N_2604,N_2967);
xnor U3625 (N_3625,N_2677,N_2938);
or U3626 (N_3626,N_2438,N_2263);
nand U3627 (N_3627,N_2557,N_2589);
nand U3628 (N_3628,N_2849,N_2921);
nor U3629 (N_3629,N_2758,N_2565);
nor U3630 (N_3630,N_2269,N_2191);
nor U3631 (N_3631,N_2905,N_2762);
nand U3632 (N_3632,N_2436,N_2190);
or U3633 (N_3633,N_2303,N_2422);
or U3634 (N_3634,N_2945,N_2819);
xor U3635 (N_3635,N_2598,N_2838);
or U3636 (N_3636,N_2696,N_2918);
nor U3637 (N_3637,N_2944,N_2728);
nor U3638 (N_3638,N_2678,N_2913);
nor U3639 (N_3639,N_2104,N_2130);
nor U3640 (N_3640,N_2583,N_2924);
or U3641 (N_3641,N_2625,N_2741);
nand U3642 (N_3642,N_2390,N_2745);
nor U3643 (N_3643,N_2414,N_2279);
nor U3644 (N_3644,N_2124,N_2641);
or U3645 (N_3645,N_2513,N_2463);
nand U3646 (N_3646,N_2894,N_2227);
nor U3647 (N_3647,N_2087,N_2049);
and U3648 (N_3648,N_2910,N_2906);
or U3649 (N_3649,N_2102,N_2571);
and U3650 (N_3650,N_2958,N_2648);
nand U3651 (N_3651,N_2369,N_2393);
nand U3652 (N_3652,N_2505,N_2990);
nand U3653 (N_3653,N_2447,N_2602);
nor U3654 (N_3654,N_2077,N_2453);
nor U3655 (N_3655,N_2168,N_2290);
and U3656 (N_3656,N_2700,N_2772);
nand U3657 (N_3657,N_2410,N_2511);
and U3658 (N_3658,N_2757,N_2537);
and U3659 (N_3659,N_2515,N_2100);
or U3660 (N_3660,N_2996,N_2185);
or U3661 (N_3661,N_2753,N_2468);
nor U3662 (N_3662,N_2632,N_2188);
and U3663 (N_3663,N_2155,N_2210);
nand U3664 (N_3664,N_2745,N_2622);
nand U3665 (N_3665,N_2562,N_2700);
and U3666 (N_3666,N_2375,N_2327);
or U3667 (N_3667,N_2748,N_2181);
and U3668 (N_3668,N_2830,N_2113);
nor U3669 (N_3669,N_2011,N_2382);
and U3670 (N_3670,N_2915,N_2592);
nor U3671 (N_3671,N_2947,N_2113);
and U3672 (N_3672,N_2065,N_2802);
nand U3673 (N_3673,N_2447,N_2620);
nor U3674 (N_3674,N_2730,N_2922);
and U3675 (N_3675,N_2968,N_2261);
nor U3676 (N_3676,N_2192,N_2269);
nand U3677 (N_3677,N_2413,N_2432);
or U3678 (N_3678,N_2602,N_2728);
and U3679 (N_3679,N_2519,N_2593);
nor U3680 (N_3680,N_2616,N_2351);
nand U3681 (N_3681,N_2731,N_2426);
and U3682 (N_3682,N_2441,N_2958);
nor U3683 (N_3683,N_2712,N_2485);
nand U3684 (N_3684,N_2643,N_2962);
or U3685 (N_3685,N_2205,N_2944);
nor U3686 (N_3686,N_2741,N_2628);
and U3687 (N_3687,N_2142,N_2544);
and U3688 (N_3688,N_2904,N_2568);
nor U3689 (N_3689,N_2965,N_2430);
and U3690 (N_3690,N_2645,N_2801);
nand U3691 (N_3691,N_2107,N_2159);
and U3692 (N_3692,N_2789,N_2694);
and U3693 (N_3693,N_2593,N_2701);
or U3694 (N_3694,N_2127,N_2655);
or U3695 (N_3695,N_2106,N_2993);
nand U3696 (N_3696,N_2688,N_2344);
nand U3697 (N_3697,N_2843,N_2765);
and U3698 (N_3698,N_2722,N_2474);
and U3699 (N_3699,N_2651,N_2747);
nor U3700 (N_3700,N_2831,N_2020);
nand U3701 (N_3701,N_2622,N_2051);
and U3702 (N_3702,N_2075,N_2920);
or U3703 (N_3703,N_2261,N_2376);
nand U3704 (N_3704,N_2165,N_2253);
nand U3705 (N_3705,N_2153,N_2549);
or U3706 (N_3706,N_2051,N_2400);
nand U3707 (N_3707,N_2997,N_2839);
nor U3708 (N_3708,N_2215,N_2386);
nand U3709 (N_3709,N_2241,N_2948);
nor U3710 (N_3710,N_2655,N_2088);
and U3711 (N_3711,N_2550,N_2557);
and U3712 (N_3712,N_2571,N_2539);
or U3713 (N_3713,N_2527,N_2124);
nor U3714 (N_3714,N_2500,N_2050);
nand U3715 (N_3715,N_2866,N_2321);
nor U3716 (N_3716,N_2445,N_2970);
nor U3717 (N_3717,N_2502,N_2059);
and U3718 (N_3718,N_2414,N_2031);
nand U3719 (N_3719,N_2903,N_2714);
nor U3720 (N_3720,N_2267,N_2222);
nor U3721 (N_3721,N_2556,N_2250);
nand U3722 (N_3722,N_2376,N_2412);
nor U3723 (N_3723,N_2502,N_2229);
or U3724 (N_3724,N_2762,N_2252);
nor U3725 (N_3725,N_2660,N_2474);
or U3726 (N_3726,N_2870,N_2354);
or U3727 (N_3727,N_2670,N_2486);
and U3728 (N_3728,N_2640,N_2301);
nor U3729 (N_3729,N_2899,N_2219);
nand U3730 (N_3730,N_2447,N_2499);
nor U3731 (N_3731,N_2080,N_2031);
or U3732 (N_3732,N_2468,N_2924);
and U3733 (N_3733,N_2962,N_2572);
and U3734 (N_3734,N_2011,N_2231);
nand U3735 (N_3735,N_2569,N_2488);
nor U3736 (N_3736,N_2775,N_2045);
nand U3737 (N_3737,N_2124,N_2155);
nand U3738 (N_3738,N_2347,N_2641);
nor U3739 (N_3739,N_2723,N_2219);
or U3740 (N_3740,N_2410,N_2980);
nor U3741 (N_3741,N_2617,N_2200);
nand U3742 (N_3742,N_2130,N_2066);
or U3743 (N_3743,N_2674,N_2708);
nor U3744 (N_3744,N_2892,N_2904);
nand U3745 (N_3745,N_2976,N_2462);
nand U3746 (N_3746,N_2967,N_2233);
or U3747 (N_3747,N_2309,N_2494);
nor U3748 (N_3748,N_2975,N_2336);
nand U3749 (N_3749,N_2285,N_2744);
or U3750 (N_3750,N_2197,N_2763);
nor U3751 (N_3751,N_2401,N_2801);
nand U3752 (N_3752,N_2488,N_2800);
nor U3753 (N_3753,N_2321,N_2260);
nor U3754 (N_3754,N_2178,N_2919);
nor U3755 (N_3755,N_2963,N_2535);
and U3756 (N_3756,N_2171,N_2096);
and U3757 (N_3757,N_2924,N_2633);
nand U3758 (N_3758,N_2826,N_2023);
and U3759 (N_3759,N_2429,N_2341);
nand U3760 (N_3760,N_2772,N_2140);
or U3761 (N_3761,N_2083,N_2856);
nor U3762 (N_3762,N_2216,N_2154);
nand U3763 (N_3763,N_2189,N_2580);
and U3764 (N_3764,N_2336,N_2450);
nor U3765 (N_3765,N_2301,N_2845);
nor U3766 (N_3766,N_2948,N_2816);
nor U3767 (N_3767,N_2930,N_2753);
and U3768 (N_3768,N_2888,N_2574);
nor U3769 (N_3769,N_2299,N_2474);
or U3770 (N_3770,N_2139,N_2082);
and U3771 (N_3771,N_2694,N_2962);
or U3772 (N_3772,N_2687,N_2601);
nor U3773 (N_3773,N_2345,N_2967);
nand U3774 (N_3774,N_2374,N_2938);
nor U3775 (N_3775,N_2645,N_2623);
nand U3776 (N_3776,N_2252,N_2432);
or U3777 (N_3777,N_2432,N_2848);
or U3778 (N_3778,N_2152,N_2789);
or U3779 (N_3779,N_2676,N_2458);
and U3780 (N_3780,N_2227,N_2019);
and U3781 (N_3781,N_2745,N_2288);
or U3782 (N_3782,N_2015,N_2393);
nand U3783 (N_3783,N_2049,N_2033);
and U3784 (N_3784,N_2809,N_2620);
nand U3785 (N_3785,N_2892,N_2255);
nor U3786 (N_3786,N_2568,N_2175);
or U3787 (N_3787,N_2811,N_2982);
nand U3788 (N_3788,N_2189,N_2828);
and U3789 (N_3789,N_2500,N_2991);
nor U3790 (N_3790,N_2293,N_2737);
or U3791 (N_3791,N_2435,N_2647);
and U3792 (N_3792,N_2213,N_2389);
and U3793 (N_3793,N_2164,N_2299);
and U3794 (N_3794,N_2806,N_2198);
nor U3795 (N_3795,N_2474,N_2141);
or U3796 (N_3796,N_2096,N_2273);
nor U3797 (N_3797,N_2363,N_2558);
nor U3798 (N_3798,N_2098,N_2471);
nand U3799 (N_3799,N_2864,N_2313);
nand U3800 (N_3800,N_2171,N_2750);
and U3801 (N_3801,N_2302,N_2935);
or U3802 (N_3802,N_2412,N_2159);
or U3803 (N_3803,N_2645,N_2991);
nand U3804 (N_3804,N_2859,N_2373);
nor U3805 (N_3805,N_2803,N_2880);
and U3806 (N_3806,N_2099,N_2030);
nand U3807 (N_3807,N_2097,N_2691);
and U3808 (N_3808,N_2849,N_2576);
or U3809 (N_3809,N_2778,N_2626);
nor U3810 (N_3810,N_2272,N_2303);
or U3811 (N_3811,N_2706,N_2731);
and U3812 (N_3812,N_2318,N_2689);
and U3813 (N_3813,N_2372,N_2389);
or U3814 (N_3814,N_2774,N_2089);
nor U3815 (N_3815,N_2635,N_2011);
nand U3816 (N_3816,N_2933,N_2763);
or U3817 (N_3817,N_2311,N_2121);
nor U3818 (N_3818,N_2184,N_2266);
nor U3819 (N_3819,N_2982,N_2130);
and U3820 (N_3820,N_2148,N_2827);
nor U3821 (N_3821,N_2775,N_2935);
nand U3822 (N_3822,N_2119,N_2979);
nor U3823 (N_3823,N_2826,N_2958);
or U3824 (N_3824,N_2273,N_2226);
nor U3825 (N_3825,N_2386,N_2027);
nor U3826 (N_3826,N_2962,N_2632);
nand U3827 (N_3827,N_2018,N_2374);
nor U3828 (N_3828,N_2698,N_2231);
nor U3829 (N_3829,N_2833,N_2789);
nand U3830 (N_3830,N_2528,N_2204);
or U3831 (N_3831,N_2393,N_2046);
nand U3832 (N_3832,N_2294,N_2492);
and U3833 (N_3833,N_2337,N_2221);
nand U3834 (N_3834,N_2212,N_2246);
or U3835 (N_3835,N_2019,N_2846);
nor U3836 (N_3836,N_2767,N_2418);
nor U3837 (N_3837,N_2877,N_2077);
or U3838 (N_3838,N_2620,N_2098);
xor U3839 (N_3839,N_2489,N_2263);
nor U3840 (N_3840,N_2371,N_2583);
and U3841 (N_3841,N_2570,N_2654);
and U3842 (N_3842,N_2171,N_2261);
or U3843 (N_3843,N_2089,N_2809);
nand U3844 (N_3844,N_2776,N_2686);
nand U3845 (N_3845,N_2904,N_2130);
and U3846 (N_3846,N_2277,N_2762);
and U3847 (N_3847,N_2495,N_2982);
nor U3848 (N_3848,N_2271,N_2235);
or U3849 (N_3849,N_2747,N_2610);
nand U3850 (N_3850,N_2102,N_2217);
or U3851 (N_3851,N_2285,N_2843);
nand U3852 (N_3852,N_2891,N_2716);
nand U3853 (N_3853,N_2028,N_2754);
and U3854 (N_3854,N_2447,N_2278);
or U3855 (N_3855,N_2634,N_2742);
and U3856 (N_3856,N_2271,N_2840);
nand U3857 (N_3857,N_2550,N_2684);
nor U3858 (N_3858,N_2156,N_2851);
and U3859 (N_3859,N_2906,N_2026);
nand U3860 (N_3860,N_2697,N_2329);
nor U3861 (N_3861,N_2891,N_2433);
or U3862 (N_3862,N_2316,N_2430);
and U3863 (N_3863,N_2160,N_2722);
nand U3864 (N_3864,N_2955,N_2047);
nor U3865 (N_3865,N_2688,N_2078);
nor U3866 (N_3866,N_2245,N_2994);
nor U3867 (N_3867,N_2364,N_2941);
nand U3868 (N_3868,N_2353,N_2646);
nor U3869 (N_3869,N_2744,N_2596);
or U3870 (N_3870,N_2902,N_2580);
or U3871 (N_3871,N_2474,N_2843);
or U3872 (N_3872,N_2847,N_2238);
and U3873 (N_3873,N_2142,N_2241);
nand U3874 (N_3874,N_2466,N_2966);
and U3875 (N_3875,N_2125,N_2742);
or U3876 (N_3876,N_2411,N_2718);
and U3877 (N_3877,N_2567,N_2004);
and U3878 (N_3878,N_2237,N_2719);
nor U3879 (N_3879,N_2083,N_2052);
nor U3880 (N_3880,N_2081,N_2694);
nand U3881 (N_3881,N_2764,N_2170);
or U3882 (N_3882,N_2685,N_2527);
and U3883 (N_3883,N_2407,N_2555);
and U3884 (N_3884,N_2083,N_2292);
or U3885 (N_3885,N_2766,N_2581);
or U3886 (N_3886,N_2340,N_2762);
and U3887 (N_3887,N_2787,N_2771);
nor U3888 (N_3888,N_2937,N_2577);
nor U3889 (N_3889,N_2561,N_2942);
or U3890 (N_3890,N_2178,N_2757);
and U3891 (N_3891,N_2873,N_2353);
and U3892 (N_3892,N_2886,N_2055);
nor U3893 (N_3893,N_2052,N_2965);
and U3894 (N_3894,N_2429,N_2548);
or U3895 (N_3895,N_2447,N_2716);
nand U3896 (N_3896,N_2971,N_2657);
and U3897 (N_3897,N_2025,N_2006);
or U3898 (N_3898,N_2134,N_2305);
nor U3899 (N_3899,N_2094,N_2417);
and U3900 (N_3900,N_2347,N_2208);
and U3901 (N_3901,N_2543,N_2040);
nand U3902 (N_3902,N_2440,N_2236);
and U3903 (N_3903,N_2126,N_2769);
nand U3904 (N_3904,N_2489,N_2744);
nor U3905 (N_3905,N_2784,N_2979);
and U3906 (N_3906,N_2578,N_2754);
nor U3907 (N_3907,N_2212,N_2409);
nand U3908 (N_3908,N_2546,N_2660);
and U3909 (N_3909,N_2268,N_2988);
nor U3910 (N_3910,N_2920,N_2926);
nand U3911 (N_3911,N_2249,N_2609);
or U3912 (N_3912,N_2995,N_2239);
or U3913 (N_3913,N_2107,N_2764);
nand U3914 (N_3914,N_2023,N_2908);
nand U3915 (N_3915,N_2703,N_2776);
and U3916 (N_3916,N_2531,N_2820);
and U3917 (N_3917,N_2847,N_2160);
nor U3918 (N_3918,N_2343,N_2469);
and U3919 (N_3919,N_2227,N_2900);
nor U3920 (N_3920,N_2455,N_2747);
nor U3921 (N_3921,N_2668,N_2453);
and U3922 (N_3922,N_2363,N_2505);
nor U3923 (N_3923,N_2620,N_2680);
nand U3924 (N_3924,N_2202,N_2672);
nand U3925 (N_3925,N_2775,N_2137);
and U3926 (N_3926,N_2680,N_2131);
or U3927 (N_3927,N_2964,N_2140);
or U3928 (N_3928,N_2155,N_2374);
nor U3929 (N_3929,N_2860,N_2609);
and U3930 (N_3930,N_2673,N_2634);
and U3931 (N_3931,N_2980,N_2737);
or U3932 (N_3932,N_2303,N_2346);
nand U3933 (N_3933,N_2145,N_2569);
nand U3934 (N_3934,N_2110,N_2372);
nor U3935 (N_3935,N_2583,N_2334);
nor U3936 (N_3936,N_2937,N_2738);
nor U3937 (N_3937,N_2054,N_2742);
and U3938 (N_3938,N_2262,N_2563);
and U3939 (N_3939,N_2018,N_2029);
or U3940 (N_3940,N_2410,N_2442);
nor U3941 (N_3941,N_2732,N_2928);
nand U3942 (N_3942,N_2014,N_2069);
and U3943 (N_3943,N_2178,N_2268);
nand U3944 (N_3944,N_2329,N_2957);
or U3945 (N_3945,N_2153,N_2258);
nor U3946 (N_3946,N_2530,N_2249);
nand U3947 (N_3947,N_2571,N_2706);
nand U3948 (N_3948,N_2111,N_2823);
nand U3949 (N_3949,N_2785,N_2815);
or U3950 (N_3950,N_2422,N_2935);
nand U3951 (N_3951,N_2726,N_2522);
and U3952 (N_3952,N_2606,N_2071);
nor U3953 (N_3953,N_2372,N_2198);
nor U3954 (N_3954,N_2432,N_2446);
nor U3955 (N_3955,N_2276,N_2642);
xnor U3956 (N_3956,N_2262,N_2350);
or U3957 (N_3957,N_2440,N_2893);
nor U3958 (N_3958,N_2368,N_2711);
or U3959 (N_3959,N_2817,N_2553);
nand U3960 (N_3960,N_2556,N_2148);
nand U3961 (N_3961,N_2283,N_2690);
nand U3962 (N_3962,N_2716,N_2239);
and U3963 (N_3963,N_2427,N_2599);
or U3964 (N_3964,N_2535,N_2207);
and U3965 (N_3965,N_2950,N_2201);
nor U3966 (N_3966,N_2239,N_2736);
and U3967 (N_3967,N_2557,N_2011);
and U3968 (N_3968,N_2801,N_2259);
or U3969 (N_3969,N_2834,N_2797);
and U3970 (N_3970,N_2149,N_2546);
and U3971 (N_3971,N_2839,N_2209);
and U3972 (N_3972,N_2583,N_2453);
nand U3973 (N_3973,N_2005,N_2786);
nand U3974 (N_3974,N_2499,N_2137);
nor U3975 (N_3975,N_2145,N_2287);
nor U3976 (N_3976,N_2975,N_2087);
nand U3977 (N_3977,N_2469,N_2000);
nand U3978 (N_3978,N_2017,N_2303);
nand U3979 (N_3979,N_2067,N_2148);
nor U3980 (N_3980,N_2900,N_2174);
and U3981 (N_3981,N_2095,N_2948);
nor U3982 (N_3982,N_2636,N_2613);
and U3983 (N_3983,N_2822,N_2987);
or U3984 (N_3984,N_2412,N_2607);
nand U3985 (N_3985,N_2994,N_2145);
nand U3986 (N_3986,N_2045,N_2674);
or U3987 (N_3987,N_2832,N_2711);
nand U3988 (N_3988,N_2019,N_2173);
nor U3989 (N_3989,N_2797,N_2224);
or U3990 (N_3990,N_2165,N_2891);
and U3991 (N_3991,N_2403,N_2739);
and U3992 (N_3992,N_2039,N_2307);
or U3993 (N_3993,N_2600,N_2669);
nand U3994 (N_3994,N_2364,N_2107);
nand U3995 (N_3995,N_2887,N_2690);
and U3996 (N_3996,N_2566,N_2679);
or U3997 (N_3997,N_2001,N_2490);
or U3998 (N_3998,N_2315,N_2879);
nor U3999 (N_3999,N_2448,N_2445);
nor U4000 (N_4000,N_3273,N_3266);
and U4001 (N_4001,N_3896,N_3921);
nand U4002 (N_4002,N_3474,N_3036);
nand U4003 (N_4003,N_3932,N_3803);
nand U4004 (N_4004,N_3115,N_3804);
nand U4005 (N_4005,N_3145,N_3869);
nor U4006 (N_4006,N_3245,N_3829);
nand U4007 (N_4007,N_3868,N_3898);
and U4008 (N_4008,N_3989,N_3355);
and U4009 (N_4009,N_3359,N_3949);
nand U4010 (N_4010,N_3909,N_3040);
or U4011 (N_4011,N_3992,N_3608);
nor U4012 (N_4012,N_3322,N_3328);
nor U4013 (N_4013,N_3690,N_3627);
and U4014 (N_4014,N_3200,N_3546);
nand U4015 (N_4015,N_3089,N_3060);
nand U4016 (N_4016,N_3802,N_3498);
and U4017 (N_4017,N_3648,N_3346);
nand U4018 (N_4018,N_3053,N_3764);
nor U4019 (N_4019,N_3864,N_3001);
nor U4020 (N_4020,N_3570,N_3470);
or U4021 (N_4021,N_3042,N_3452);
nor U4022 (N_4022,N_3796,N_3335);
nand U4023 (N_4023,N_3344,N_3997);
nand U4024 (N_4024,N_3289,N_3173);
and U4025 (N_4025,N_3126,N_3084);
nand U4026 (N_4026,N_3419,N_3483);
nor U4027 (N_4027,N_3268,N_3315);
nor U4028 (N_4028,N_3025,N_3068);
nor U4029 (N_4029,N_3103,N_3774);
or U4030 (N_4030,N_3890,N_3778);
and U4031 (N_4031,N_3426,N_3882);
nor U4032 (N_4032,N_3101,N_3350);
and U4033 (N_4033,N_3855,N_3611);
or U4034 (N_4034,N_3842,N_3505);
and U4035 (N_4035,N_3279,N_3747);
nor U4036 (N_4036,N_3693,N_3100);
xnor U4037 (N_4037,N_3277,N_3584);
xnor U4038 (N_4038,N_3246,N_3565);
and U4039 (N_4039,N_3554,N_3749);
and U4040 (N_4040,N_3230,N_3338);
and U4041 (N_4041,N_3791,N_3991);
and U4042 (N_4042,N_3724,N_3961);
nor U4043 (N_4043,N_3951,N_3574);
or U4044 (N_4044,N_3139,N_3159);
and U4045 (N_4045,N_3889,N_3895);
nand U4046 (N_4046,N_3244,N_3821);
and U4047 (N_4047,N_3027,N_3958);
or U4048 (N_4048,N_3886,N_3447);
nand U4049 (N_4049,N_3336,N_3538);
nor U4050 (N_4050,N_3500,N_3734);
nor U4051 (N_4051,N_3222,N_3286);
or U4052 (N_4052,N_3475,N_3697);
nor U4053 (N_4053,N_3105,N_3699);
nor U4054 (N_4054,N_3398,N_3317);
and U4055 (N_4055,N_3768,N_3963);
nor U4056 (N_4056,N_3742,N_3823);
or U4057 (N_4057,N_3748,N_3850);
or U4058 (N_4058,N_3014,N_3861);
or U4059 (N_4059,N_3463,N_3352);
and U4060 (N_4060,N_3662,N_3930);
and U4061 (N_4061,N_3226,N_3251);
and U4062 (N_4062,N_3950,N_3467);
and U4063 (N_4063,N_3123,N_3037);
or U4064 (N_4064,N_3739,N_3518);
nand U4065 (N_4065,N_3225,N_3333);
and U4066 (N_4066,N_3603,N_3309);
and U4067 (N_4067,N_3334,N_3032);
or U4068 (N_4068,N_3642,N_3598);
nand U4069 (N_4069,N_3982,N_3920);
or U4070 (N_4070,N_3468,N_3947);
nor U4071 (N_4071,N_3516,N_3329);
or U4072 (N_4072,N_3704,N_3425);
nor U4073 (N_4073,N_3388,N_3087);
nor U4074 (N_4074,N_3683,N_3806);
nor U4075 (N_4075,N_3323,N_3576);
xor U4076 (N_4076,N_3255,N_3210);
nor U4077 (N_4077,N_3363,N_3128);
or U4078 (N_4078,N_3853,N_3149);
or U4079 (N_4079,N_3974,N_3685);
nor U4080 (N_4080,N_3540,N_3472);
or U4081 (N_4081,N_3617,N_3296);
and U4082 (N_4082,N_3899,N_3741);
or U4083 (N_4083,N_3075,N_3833);
and U4084 (N_4084,N_3239,N_3867);
nand U4085 (N_4085,N_3863,N_3763);
nor U4086 (N_4086,N_3029,N_3519);
nand U4087 (N_4087,N_3043,N_3348);
nand U4088 (N_4088,N_3637,N_3848);
and U4089 (N_4089,N_3368,N_3097);
nand U4090 (N_4090,N_3142,N_3085);
or U4091 (N_4091,N_3612,N_3714);
nand U4092 (N_4092,N_3917,N_3428);
and U4093 (N_4093,N_3358,N_3736);
and U4094 (N_4094,N_3187,N_3526);
nand U4095 (N_4095,N_3914,N_3031);
and U4096 (N_4096,N_3413,N_3487);
nor U4097 (N_4097,N_3249,N_3202);
nor U4098 (N_4098,N_3347,N_3373);
nand U4099 (N_4099,N_3086,N_3223);
and U4100 (N_4100,N_3935,N_3593);
and U4101 (N_4101,N_3504,N_3872);
and U4102 (N_4102,N_3532,N_3525);
nor U4103 (N_4103,N_3826,N_3232);
or U4104 (N_4104,N_3253,N_3773);
nor U4105 (N_4105,N_3401,N_3229);
nand U4106 (N_4106,N_3651,N_3883);
or U4107 (N_4107,N_3012,N_3281);
nand U4108 (N_4108,N_3915,N_3464);
and U4109 (N_4109,N_3479,N_3288);
and U4110 (N_4110,N_3605,N_3018);
nor U4111 (N_4111,N_3726,N_3473);
or U4112 (N_4112,N_3046,N_3619);
or U4113 (N_4113,N_3929,N_3759);
nand U4114 (N_4114,N_3687,N_3894);
nor U4115 (N_4115,N_3050,N_3843);
or U4116 (N_4116,N_3160,N_3181);
nor U4117 (N_4117,N_3962,N_3865);
and U4118 (N_4118,N_3379,N_3201);
nor U4119 (N_4119,N_3258,N_3108);
or U4120 (N_4120,N_3730,N_3874);
or U4121 (N_4121,N_3357,N_3583);
nor U4122 (N_4122,N_3313,N_3389);
or U4123 (N_4123,N_3321,N_3717);
nand U4124 (N_4124,N_3820,N_3545);
and U4125 (N_4125,N_3204,N_3190);
or U4126 (N_4126,N_3019,N_3632);
nor U4127 (N_4127,N_3420,N_3035);
and U4128 (N_4128,N_3134,N_3297);
and U4129 (N_4129,N_3137,N_3020);
or U4130 (N_4130,N_3613,N_3553);
or U4131 (N_4131,N_3713,N_3711);
and U4132 (N_4132,N_3393,N_3331);
or U4133 (N_4133,N_3444,N_3660);
or U4134 (N_4134,N_3503,N_3146);
nor U4135 (N_4135,N_3870,N_3852);
nand U4136 (N_4136,N_3508,N_3440);
or U4137 (N_4137,N_3096,N_3410);
and U4138 (N_4138,N_3625,N_3912);
nor U4139 (N_4139,N_3016,N_3345);
or U4140 (N_4140,N_3445,N_3725);
and U4141 (N_4141,N_3509,N_3620);
or U4142 (N_4142,N_3606,N_3955);
and U4143 (N_4143,N_3234,N_3924);
nand U4144 (N_4144,N_3892,N_3885);
nand U4145 (N_4145,N_3933,N_3422);
and U4146 (N_4146,N_3825,N_3117);
or U4147 (N_4147,N_3477,N_3589);
and U4148 (N_4148,N_3536,N_3495);
nand U4149 (N_4149,N_3460,N_3983);
or U4150 (N_4150,N_3969,N_3877);
nor U4151 (N_4151,N_3623,N_3878);
and U4152 (N_4152,N_3788,N_3291);
nand U4153 (N_4153,N_3158,N_3506);
or U4154 (N_4154,N_3985,N_3166);
nand U4155 (N_4155,N_3026,N_3702);
nor U4156 (N_4156,N_3607,N_3417);
nand U4157 (N_4157,N_3165,N_3072);
nor U4158 (N_4158,N_3716,N_3143);
or U4159 (N_4159,N_3111,N_3340);
or U4160 (N_4160,N_3925,N_3396);
or U4161 (N_4161,N_3757,N_3649);
and U4162 (N_4162,N_3275,N_3449);
nand U4163 (N_4163,N_3937,N_3265);
nor U4164 (N_4164,N_3446,N_3399);
or U4165 (N_4165,N_3911,N_3384);
nand U4166 (N_4166,N_3127,N_3926);
nand U4167 (N_4167,N_3183,N_3065);
and U4168 (N_4168,N_3125,N_3318);
nand U4169 (N_4169,N_3070,N_3694);
nor U4170 (N_4170,N_3762,N_3793);
and U4171 (N_4171,N_3539,N_3119);
or U4172 (N_4172,N_3847,N_3339);
or U4173 (N_4173,N_3209,N_3481);
or U4174 (N_4174,N_3535,N_3161);
or U4175 (N_4175,N_3575,N_3164);
nor U4176 (N_4176,N_3840,N_3723);
or U4177 (N_4177,N_3988,N_3186);
nand U4178 (N_4178,N_3354,N_3695);
or U4179 (N_4179,N_3615,N_3799);
and U4180 (N_4180,N_3585,N_3549);
or U4181 (N_4181,N_3008,N_3370);
and U4182 (N_4182,N_3692,N_3755);
and U4183 (N_4183,N_3066,N_3228);
nor U4184 (N_4184,N_3372,N_3942);
nor U4185 (N_4185,N_3681,N_3062);
nand U4186 (N_4186,N_3858,N_3174);
or U4187 (N_4187,N_3436,N_3626);
or U4188 (N_4188,N_3217,N_3691);
nor U4189 (N_4189,N_3720,N_3324);
and U4190 (N_4190,N_3392,N_3800);
or U4191 (N_4191,N_3601,N_3064);
and U4192 (N_4192,N_3953,N_3492);
nor U4193 (N_4193,N_3657,N_3835);
nor U4194 (N_4194,N_3750,N_3709);
xor U4195 (N_4195,N_3990,N_3088);
nor U4196 (N_4196,N_3740,N_3079);
nor U4197 (N_4197,N_3529,N_3300);
nand U4198 (N_4198,N_3592,N_3795);
or U4199 (N_4199,N_3458,N_3466);
nor U4200 (N_4200,N_3203,N_3644);
nor U4201 (N_4201,N_3394,N_3729);
nand U4202 (N_4202,N_3367,N_3023);
and U4203 (N_4203,N_3423,N_3490);
and U4204 (N_4204,N_3743,N_3561);
or U4205 (N_4205,N_3563,N_3298);
or U4206 (N_4206,N_3786,N_3150);
and U4207 (N_4207,N_3587,N_3718);
nand U4208 (N_4208,N_3378,N_3941);
nand U4209 (N_4209,N_3319,N_3881);
and U4210 (N_4210,N_3443,N_3973);
nand U4211 (N_4211,N_3531,N_3812);
nand U4212 (N_4212,N_3212,N_3414);
xor U4213 (N_4213,N_3261,N_3674);
and U4214 (N_4214,N_3185,N_3263);
or U4215 (N_4215,N_3433,N_3283);
or U4216 (N_4216,N_3307,N_3964);
nor U4217 (N_4217,N_3517,N_3302);
nand U4218 (N_4218,N_3559,N_3332);
or U4219 (N_4219,N_3664,N_3006);
nor U4220 (N_4220,N_3844,N_3430);
nor U4221 (N_4221,N_3024,N_3972);
or U4222 (N_4222,N_3956,N_3555);
or U4223 (N_4223,N_3661,N_3513);
or U4224 (N_4224,N_3993,N_3003);
nor U4225 (N_4225,N_3597,N_3952);
and U4226 (N_4226,N_3269,N_3405);
and U4227 (N_4227,N_3815,N_3510);
nand U4228 (N_4228,N_3327,N_3011);
or U4229 (N_4229,N_3916,N_3507);
and U4230 (N_4230,N_3659,N_3670);
and U4231 (N_4231,N_3779,N_3049);
or U4232 (N_4232,N_3501,N_3193);
nand U4233 (N_4233,N_3775,N_3397);
nand U4234 (N_4234,N_3044,N_3987);
and U4235 (N_4235,N_3910,N_3631);
and U4236 (N_4236,N_3010,N_3696);
and U4237 (N_4237,N_3654,N_3927);
or U4238 (N_4238,N_3282,N_3560);
and U4239 (N_4239,N_3904,N_3280);
and U4240 (N_4240,N_3364,N_3866);
nor U4241 (N_4241,N_3454,N_3184);
nand U4242 (N_4242,N_3262,N_3076);
or U4243 (N_4243,N_3052,N_3073);
or U4244 (N_4244,N_3469,N_3996);
or U4245 (N_4245,N_3290,N_3579);
or U4246 (N_4246,N_3241,N_3577);
or U4247 (N_4247,N_3544,N_3240);
and U4248 (N_4248,N_3624,N_3442);
and U4249 (N_4249,N_3299,N_3270);
and U4250 (N_4250,N_3429,N_3248);
nand U4251 (N_4251,N_3219,N_3094);
or U4252 (N_4252,N_3017,N_3353);
and U4253 (N_4253,N_3977,N_3056);
nor U4254 (N_4254,N_3330,N_3004);
or U4255 (N_4255,N_3254,N_3527);
nor U4256 (N_4256,N_3873,N_3058);
nor U4257 (N_4257,N_3640,N_3152);
and U4258 (N_4258,N_3144,N_3580);
and U4259 (N_4259,N_3995,N_3453);
or U4260 (N_4260,N_3198,N_3682);
nand U4261 (N_4261,N_3839,N_3267);
and U4262 (N_4262,N_3633,N_3550);
nor U4263 (N_4263,N_3635,N_3737);
or U4264 (N_4264,N_3566,N_3938);
and U4265 (N_4265,N_3807,N_3294);
nor U4266 (N_4266,N_3178,N_3636);
nor U4267 (N_4267,N_3689,N_3744);
or U4268 (N_4268,N_3171,N_3845);
and U4269 (N_4269,N_3409,N_3761);
nor U4270 (N_4270,N_3292,N_3502);
and U4271 (N_4271,N_3213,N_3189);
nor U4272 (N_4272,N_3528,N_3622);
or U4273 (N_4273,N_3385,N_3887);
nor U4274 (N_4274,N_3197,N_3706);
nor U4275 (N_4275,N_3902,N_3599);
or U4276 (N_4276,N_3135,N_3721);
or U4277 (N_4277,N_3569,N_3922);
and U4278 (N_4278,N_3156,N_3207);
and U4279 (N_4279,N_3216,N_3805);
or U4280 (N_4280,N_3907,N_3939);
and U4281 (N_4281,N_3686,N_3421);
and U4282 (N_4282,N_3256,N_3424);
nand U4283 (N_4283,N_3325,N_3499);
or U4284 (N_4284,N_3221,N_3541);
nand U4285 (N_4285,N_3168,N_3703);
and U4286 (N_4286,N_3782,N_3968);
nor U4287 (N_4287,N_3512,N_3628);
nor U4288 (N_4288,N_3630,N_3391);
nor U4289 (N_4289,N_3471,N_3998);
and U4290 (N_4290,N_3196,N_3252);
nand U4291 (N_4291,N_3638,N_3028);
or U4292 (N_4292,N_3320,N_3387);
nand U4293 (N_4293,N_3979,N_3588);
or U4294 (N_4294,N_3784,N_3752);
nand U4295 (N_4295,N_3130,N_3705);
and U4296 (N_4296,N_3960,N_3403);
nor U4297 (N_4297,N_3356,N_3090);
or U4298 (N_4298,N_3754,N_3067);
nand U4299 (N_4299,N_3081,N_3530);
and U4300 (N_4300,N_3057,N_3792);
nor U4301 (N_4301,N_3667,N_3179);
and U4302 (N_4302,N_3522,N_3602);
and U4303 (N_4303,N_3641,N_3177);
or U4304 (N_4304,N_3365,N_3383);
and U4305 (N_4305,N_3643,N_3303);
and U4306 (N_4306,N_3860,N_3816);
nor U4307 (N_4307,N_3341,N_3071);
nand U4308 (N_4308,N_3722,N_3830);
nor U4309 (N_4309,N_3945,N_3155);
and U4310 (N_4310,N_3836,N_3074);
and U4311 (N_4311,N_3293,N_3944);
or U4312 (N_4312,N_3811,N_3129);
nand U4313 (N_4313,N_3063,N_3000);
xnor U4314 (N_4314,N_3231,N_3295);
and U4315 (N_4315,N_3250,N_3157);
and U4316 (N_4316,N_3059,N_3936);
nand U4317 (N_4317,N_3665,N_3954);
nand U4318 (N_4318,N_3854,N_3562);
or U4319 (N_4319,N_3571,N_3191);
nor U4320 (N_4320,N_3272,N_3680);
and U4321 (N_4321,N_3366,N_3243);
and U4322 (N_4322,N_3287,N_3647);
nor U4323 (N_4323,N_3653,N_3908);
or U4324 (N_4324,N_3822,N_3832);
and U4325 (N_4325,N_3769,N_3880);
nor U4326 (N_4326,N_3871,N_3316);
or U4327 (N_4327,N_3999,N_3375);
or U4328 (N_4328,N_3175,N_3376);
nand U4329 (N_4329,N_3192,N_3543);
and U4330 (N_4330,N_3113,N_3215);
nand U4331 (N_4331,N_3514,N_3451);
and U4332 (N_4332,N_3572,N_3491);
nor U4333 (N_4333,N_3311,N_3118);
nand U4334 (N_4334,N_3986,N_3114);
or U4335 (N_4335,N_3439,N_3061);
nand U4336 (N_4336,N_3797,N_3520);
or U4337 (N_4337,N_3274,N_3099);
and U4338 (N_4338,N_3913,N_3578);
nand U4339 (N_4339,N_3609,N_3182);
and U4340 (N_4340,N_3489,N_3900);
and U4341 (N_4341,N_3038,N_3511);
or U4342 (N_4342,N_3227,N_3879);
nand U4343 (N_4343,N_3080,N_3051);
nor U4344 (N_4344,N_3808,N_3151);
nor U4345 (N_4345,N_3484,N_3102);
nor U4346 (N_4346,N_3819,N_3362);
and U4347 (N_4347,N_3970,N_3594);
and U4348 (N_4348,N_3095,N_3668);
nor U4349 (N_4349,N_3596,N_3351);
nand U4350 (N_4350,N_3172,N_3039);
nand U4351 (N_4351,N_3776,N_3257);
nor U4352 (N_4352,N_3818,N_3783);
xnor U4353 (N_4353,N_3437,N_3701);
or U4354 (N_4354,N_3715,N_3618);
and U4355 (N_4355,N_3054,N_3971);
nand U4356 (N_4356,N_3814,N_3482);
nand U4357 (N_4357,N_3194,N_3582);
nand U4358 (N_4358,N_3790,N_3573);
nand U4359 (N_4359,N_3888,N_3548);
and U4360 (N_4360,N_3523,N_3147);
nand U4361 (N_4361,N_3259,N_3493);
nand U4362 (N_4362,N_3918,N_3310);
and U4363 (N_4363,N_3745,N_3542);
nor U4364 (N_4364,N_3903,N_3707);
or U4365 (N_4365,N_3305,N_3719);
and U4366 (N_4366,N_3634,N_3337);
or U4367 (N_4367,N_3556,N_3478);
nand U4368 (N_4368,N_3361,N_3106);
or U4369 (N_4369,N_3116,N_3837);
nor U4370 (N_4370,N_3673,N_3284);
and U4371 (N_4371,N_3712,N_3906);
nor U4372 (N_4372,N_3756,N_3343);
or U4373 (N_4373,N_3733,N_3948);
nor U4374 (N_4374,N_3676,N_3678);
or U4375 (N_4375,N_3461,N_3154);
and U4376 (N_4376,N_3663,N_3371);
or U4377 (N_4377,N_3236,N_3276);
nand U4378 (N_4378,N_3672,N_3496);
and U4379 (N_4379,N_3264,N_3271);
and U4380 (N_4380,N_3377,N_3893);
and U4381 (N_4381,N_3285,N_3838);
nand U4382 (N_4382,N_3136,N_3374);
nand U4383 (N_4383,N_3153,N_3002);
nand U4384 (N_4384,N_3777,N_3801);
or U4385 (N_4385,N_3199,N_3308);
and U4386 (N_4386,N_3732,N_3034);
nand U4387 (N_4387,N_3533,N_3557);
or U4388 (N_4388,N_3176,N_3859);
or U4389 (N_4389,N_3655,N_3940);
or U4390 (N_4390,N_3170,N_3132);
or U4391 (N_4391,N_3946,N_3669);
or U4392 (N_4392,N_3188,N_3304);
nor U4393 (N_4393,N_3476,N_3408);
nor U4394 (N_4394,N_3772,N_3923);
nand U4395 (N_4395,N_3901,N_3404);
or U4396 (N_4396,N_3238,N_3984);
nand U4397 (N_4397,N_3224,N_3005);
and U4398 (N_4398,N_3301,N_3567);
and U4399 (N_4399,N_3235,N_3810);
and U4400 (N_4400,N_3746,N_3834);
or U4401 (N_4401,N_3486,N_3122);
nand U4402 (N_4402,N_3975,N_3069);
or U4403 (N_4403,N_3104,N_3537);
nor U4404 (N_4404,N_3978,N_3427);
nand U4405 (N_4405,N_3798,N_3586);
and U4406 (N_4406,N_3698,N_3456);
or U4407 (N_4407,N_3411,N_3862);
and U4408 (N_4408,N_3934,N_3218);
nor U4409 (N_4409,N_3415,N_3395);
and U4410 (N_4410,N_3163,N_3846);
and U4411 (N_4411,N_3919,N_3831);
nand U4412 (N_4412,N_3547,N_3380);
or U4413 (N_4413,N_3030,N_3459);
nor U4414 (N_4414,N_3614,N_3434);
nand U4415 (N_4415,N_3206,N_3679);
nand U4416 (N_4416,N_3813,N_3214);
and U4417 (N_4417,N_3098,N_3959);
nand U4418 (N_4418,N_3767,N_3590);
nor U4419 (N_4419,N_3827,N_3432);
nor U4420 (N_4420,N_3360,N_3208);
or U4421 (N_4421,N_3233,N_3817);
nand U4422 (N_4422,N_3450,N_3457);
nor U4423 (N_4423,N_3078,N_3278);
nand U4424 (N_4424,N_3242,N_3581);
nand U4425 (N_4425,N_3112,N_3688);
and U4426 (N_4426,N_3728,N_3684);
nor U4427 (N_4427,N_3306,N_3671);
nand U4428 (N_4428,N_3994,N_3621);
nor U4429 (N_4429,N_3981,N_3015);
nor U4430 (N_4430,N_3211,N_3789);
nor U4431 (N_4431,N_3013,N_3794);
nor U4432 (N_4432,N_3237,N_3131);
and U4433 (N_4433,N_3857,N_3438);
nand U4434 (N_4434,N_3708,N_3406);
or U4435 (N_4435,N_3021,N_3342);
xor U4436 (N_4436,N_3677,N_3326);
and U4437 (N_4437,N_3124,N_3604);
or U4438 (N_4438,N_3650,N_3093);
nor U4439 (N_4439,N_3600,N_3760);
nor U4440 (N_4440,N_3133,N_3897);
or U4441 (N_4441,N_3407,N_3480);
or U4442 (N_4442,N_3735,N_3416);
and U4443 (N_4443,N_3418,N_3435);
nor U4444 (N_4444,N_3083,N_3652);
and U4445 (N_4445,N_3656,N_3876);
nor U4446 (N_4446,N_3727,N_3041);
nand U4447 (N_4447,N_3645,N_3082);
or U4448 (N_4448,N_3260,N_3666);
nand U4449 (N_4449,N_3465,N_3851);
and U4450 (N_4450,N_3314,N_3928);
nor U4451 (N_4451,N_3824,N_3180);
and U4452 (N_4452,N_3386,N_3770);
nand U4453 (N_4453,N_3700,N_3891);
or U4454 (N_4454,N_3765,N_3441);
nor U4455 (N_4455,N_3485,N_3966);
nand U4456 (N_4456,N_3521,N_3140);
or U4457 (N_4457,N_3167,N_3675);
nand U4458 (N_4458,N_3841,N_3884);
nand U4459 (N_4459,N_3787,N_3055);
nor U4460 (N_4460,N_3220,N_3077);
nand U4461 (N_4461,N_3091,N_3766);
or U4462 (N_4462,N_3488,N_3148);
or U4463 (N_4463,N_3048,N_3110);
nand U4464 (N_4464,N_3771,N_3107);
nor U4465 (N_4465,N_3120,N_3639);
nand U4466 (N_4466,N_3007,N_3738);
nor U4467 (N_4467,N_3616,N_3109);
nand U4468 (N_4468,N_3809,N_3534);
and U4469 (N_4469,N_3349,N_3009);
nand U4470 (N_4470,N_3448,N_3494);
nor U4471 (N_4471,N_3967,N_3205);
nor U4472 (N_4472,N_3957,N_3431);
and U4473 (N_4473,N_3564,N_3758);
nand U4474 (N_4474,N_3658,N_3856);
and U4475 (N_4475,N_3568,N_3595);
or U4476 (N_4476,N_3141,N_3195);
nor U4477 (N_4477,N_3710,N_3169);
nand U4478 (N_4478,N_3781,N_3731);
nand U4479 (N_4479,N_3515,N_3247);
and U4480 (N_4480,N_3931,N_3875);
nand U4481 (N_4481,N_3905,N_3558);
and U4482 (N_4482,N_3785,N_3753);
nor U4483 (N_4483,N_3033,N_3976);
and U4484 (N_4484,N_3980,N_3092);
or U4485 (N_4485,N_3780,N_3965);
nor U4486 (N_4486,N_3629,N_3121);
nand U4487 (N_4487,N_3162,N_3312);
or U4488 (N_4488,N_3390,N_3138);
or U4489 (N_4489,N_3849,N_3412);
nand U4490 (N_4490,N_3369,N_3552);
nor U4491 (N_4491,N_3402,N_3382);
nor U4492 (N_4492,N_3943,N_3381);
and U4493 (N_4493,N_3400,N_3524);
nor U4494 (N_4494,N_3022,N_3646);
nor U4495 (N_4495,N_3047,N_3551);
and U4496 (N_4496,N_3828,N_3497);
nand U4497 (N_4497,N_3591,N_3610);
nor U4498 (N_4498,N_3045,N_3462);
nand U4499 (N_4499,N_3751,N_3455);
or U4500 (N_4500,N_3187,N_3818);
and U4501 (N_4501,N_3061,N_3450);
or U4502 (N_4502,N_3581,N_3408);
nor U4503 (N_4503,N_3783,N_3393);
nor U4504 (N_4504,N_3752,N_3366);
nor U4505 (N_4505,N_3664,N_3361);
or U4506 (N_4506,N_3510,N_3762);
nor U4507 (N_4507,N_3908,N_3723);
nand U4508 (N_4508,N_3615,N_3217);
and U4509 (N_4509,N_3164,N_3742);
nor U4510 (N_4510,N_3579,N_3089);
nor U4511 (N_4511,N_3301,N_3777);
or U4512 (N_4512,N_3769,N_3331);
nor U4513 (N_4513,N_3506,N_3278);
nor U4514 (N_4514,N_3767,N_3760);
or U4515 (N_4515,N_3279,N_3187);
or U4516 (N_4516,N_3167,N_3158);
nor U4517 (N_4517,N_3748,N_3650);
nor U4518 (N_4518,N_3842,N_3212);
nor U4519 (N_4519,N_3572,N_3265);
nand U4520 (N_4520,N_3876,N_3366);
nor U4521 (N_4521,N_3628,N_3827);
and U4522 (N_4522,N_3434,N_3773);
nor U4523 (N_4523,N_3503,N_3245);
and U4524 (N_4524,N_3287,N_3263);
or U4525 (N_4525,N_3428,N_3687);
nand U4526 (N_4526,N_3447,N_3651);
nor U4527 (N_4527,N_3984,N_3500);
nand U4528 (N_4528,N_3817,N_3970);
or U4529 (N_4529,N_3781,N_3280);
and U4530 (N_4530,N_3104,N_3101);
and U4531 (N_4531,N_3961,N_3097);
or U4532 (N_4532,N_3024,N_3844);
and U4533 (N_4533,N_3738,N_3250);
or U4534 (N_4534,N_3668,N_3468);
or U4535 (N_4535,N_3925,N_3880);
or U4536 (N_4536,N_3137,N_3071);
or U4537 (N_4537,N_3408,N_3460);
or U4538 (N_4538,N_3302,N_3376);
nand U4539 (N_4539,N_3027,N_3689);
or U4540 (N_4540,N_3020,N_3239);
or U4541 (N_4541,N_3007,N_3606);
nand U4542 (N_4542,N_3300,N_3920);
nor U4543 (N_4543,N_3689,N_3018);
nand U4544 (N_4544,N_3786,N_3569);
nand U4545 (N_4545,N_3136,N_3478);
nand U4546 (N_4546,N_3127,N_3559);
nor U4547 (N_4547,N_3790,N_3137);
nand U4548 (N_4548,N_3387,N_3158);
nor U4549 (N_4549,N_3296,N_3066);
nand U4550 (N_4550,N_3907,N_3216);
nand U4551 (N_4551,N_3655,N_3632);
nor U4552 (N_4552,N_3545,N_3000);
nor U4553 (N_4553,N_3437,N_3990);
nand U4554 (N_4554,N_3103,N_3877);
or U4555 (N_4555,N_3232,N_3587);
and U4556 (N_4556,N_3275,N_3891);
and U4557 (N_4557,N_3816,N_3470);
and U4558 (N_4558,N_3887,N_3917);
nor U4559 (N_4559,N_3839,N_3354);
nand U4560 (N_4560,N_3589,N_3670);
nor U4561 (N_4561,N_3508,N_3937);
or U4562 (N_4562,N_3475,N_3064);
nor U4563 (N_4563,N_3099,N_3744);
and U4564 (N_4564,N_3780,N_3711);
or U4565 (N_4565,N_3272,N_3971);
or U4566 (N_4566,N_3224,N_3733);
and U4567 (N_4567,N_3571,N_3897);
nand U4568 (N_4568,N_3313,N_3662);
or U4569 (N_4569,N_3162,N_3013);
and U4570 (N_4570,N_3350,N_3390);
and U4571 (N_4571,N_3978,N_3063);
and U4572 (N_4572,N_3283,N_3175);
and U4573 (N_4573,N_3683,N_3257);
nand U4574 (N_4574,N_3715,N_3021);
nand U4575 (N_4575,N_3678,N_3310);
nor U4576 (N_4576,N_3989,N_3736);
and U4577 (N_4577,N_3648,N_3154);
or U4578 (N_4578,N_3417,N_3247);
or U4579 (N_4579,N_3935,N_3866);
nor U4580 (N_4580,N_3098,N_3061);
and U4581 (N_4581,N_3803,N_3928);
nor U4582 (N_4582,N_3258,N_3121);
and U4583 (N_4583,N_3444,N_3467);
and U4584 (N_4584,N_3138,N_3168);
nor U4585 (N_4585,N_3736,N_3294);
nor U4586 (N_4586,N_3128,N_3611);
nand U4587 (N_4587,N_3107,N_3749);
nand U4588 (N_4588,N_3842,N_3715);
xor U4589 (N_4589,N_3743,N_3672);
and U4590 (N_4590,N_3926,N_3435);
or U4591 (N_4591,N_3477,N_3892);
and U4592 (N_4592,N_3000,N_3002);
nand U4593 (N_4593,N_3137,N_3553);
and U4594 (N_4594,N_3861,N_3723);
and U4595 (N_4595,N_3755,N_3981);
xor U4596 (N_4596,N_3871,N_3235);
or U4597 (N_4597,N_3954,N_3349);
or U4598 (N_4598,N_3005,N_3420);
nand U4599 (N_4599,N_3310,N_3500);
or U4600 (N_4600,N_3021,N_3028);
and U4601 (N_4601,N_3669,N_3608);
nor U4602 (N_4602,N_3321,N_3059);
xnor U4603 (N_4603,N_3773,N_3025);
and U4604 (N_4604,N_3000,N_3787);
nand U4605 (N_4605,N_3450,N_3576);
or U4606 (N_4606,N_3671,N_3221);
or U4607 (N_4607,N_3403,N_3310);
and U4608 (N_4608,N_3126,N_3218);
and U4609 (N_4609,N_3910,N_3058);
or U4610 (N_4610,N_3912,N_3616);
nor U4611 (N_4611,N_3868,N_3343);
nor U4612 (N_4612,N_3961,N_3449);
or U4613 (N_4613,N_3283,N_3769);
or U4614 (N_4614,N_3617,N_3359);
or U4615 (N_4615,N_3263,N_3795);
or U4616 (N_4616,N_3998,N_3754);
xor U4617 (N_4617,N_3975,N_3862);
or U4618 (N_4618,N_3146,N_3106);
and U4619 (N_4619,N_3405,N_3119);
nand U4620 (N_4620,N_3674,N_3101);
or U4621 (N_4621,N_3363,N_3217);
or U4622 (N_4622,N_3533,N_3852);
and U4623 (N_4623,N_3477,N_3662);
or U4624 (N_4624,N_3444,N_3818);
nand U4625 (N_4625,N_3370,N_3753);
or U4626 (N_4626,N_3653,N_3516);
and U4627 (N_4627,N_3095,N_3796);
nor U4628 (N_4628,N_3184,N_3351);
nand U4629 (N_4629,N_3947,N_3819);
and U4630 (N_4630,N_3930,N_3407);
and U4631 (N_4631,N_3425,N_3249);
nor U4632 (N_4632,N_3538,N_3781);
or U4633 (N_4633,N_3308,N_3461);
nand U4634 (N_4634,N_3745,N_3362);
or U4635 (N_4635,N_3960,N_3971);
nand U4636 (N_4636,N_3739,N_3825);
and U4637 (N_4637,N_3833,N_3615);
or U4638 (N_4638,N_3068,N_3160);
and U4639 (N_4639,N_3013,N_3316);
or U4640 (N_4640,N_3883,N_3079);
nand U4641 (N_4641,N_3002,N_3031);
and U4642 (N_4642,N_3631,N_3657);
nand U4643 (N_4643,N_3760,N_3398);
nand U4644 (N_4644,N_3917,N_3337);
nor U4645 (N_4645,N_3510,N_3495);
nor U4646 (N_4646,N_3611,N_3794);
and U4647 (N_4647,N_3451,N_3566);
or U4648 (N_4648,N_3629,N_3589);
nor U4649 (N_4649,N_3084,N_3501);
nor U4650 (N_4650,N_3344,N_3386);
nand U4651 (N_4651,N_3008,N_3649);
nor U4652 (N_4652,N_3737,N_3141);
nand U4653 (N_4653,N_3935,N_3061);
and U4654 (N_4654,N_3280,N_3902);
nor U4655 (N_4655,N_3798,N_3852);
or U4656 (N_4656,N_3362,N_3759);
nand U4657 (N_4657,N_3476,N_3712);
nand U4658 (N_4658,N_3841,N_3463);
nor U4659 (N_4659,N_3470,N_3292);
nor U4660 (N_4660,N_3849,N_3231);
nand U4661 (N_4661,N_3791,N_3724);
or U4662 (N_4662,N_3422,N_3689);
nor U4663 (N_4663,N_3683,N_3161);
xnor U4664 (N_4664,N_3882,N_3639);
nor U4665 (N_4665,N_3582,N_3986);
nand U4666 (N_4666,N_3379,N_3294);
nand U4667 (N_4667,N_3005,N_3466);
or U4668 (N_4668,N_3391,N_3966);
nor U4669 (N_4669,N_3416,N_3405);
and U4670 (N_4670,N_3192,N_3501);
or U4671 (N_4671,N_3094,N_3977);
xor U4672 (N_4672,N_3493,N_3970);
nor U4673 (N_4673,N_3147,N_3878);
and U4674 (N_4674,N_3978,N_3489);
nor U4675 (N_4675,N_3238,N_3481);
and U4676 (N_4676,N_3314,N_3441);
and U4677 (N_4677,N_3319,N_3803);
and U4678 (N_4678,N_3231,N_3707);
nor U4679 (N_4679,N_3273,N_3224);
nor U4680 (N_4680,N_3223,N_3174);
nand U4681 (N_4681,N_3381,N_3554);
nor U4682 (N_4682,N_3780,N_3798);
or U4683 (N_4683,N_3595,N_3118);
nand U4684 (N_4684,N_3002,N_3321);
nand U4685 (N_4685,N_3827,N_3612);
and U4686 (N_4686,N_3141,N_3033);
nor U4687 (N_4687,N_3563,N_3726);
or U4688 (N_4688,N_3840,N_3207);
and U4689 (N_4689,N_3444,N_3999);
nand U4690 (N_4690,N_3946,N_3598);
nor U4691 (N_4691,N_3028,N_3123);
or U4692 (N_4692,N_3830,N_3861);
and U4693 (N_4693,N_3610,N_3705);
nor U4694 (N_4694,N_3179,N_3828);
and U4695 (N_4695,N_3552,N_3018);
nor U4696 (N_4696,N_3389,N_3087);
or U4697 (N_4697,N_3556,N_3490);
nand U4698 (N_4698,N_3195,N_3500);
nand U4699 (N_4699,N_3739,N_3596);
or U4700 (N_4700,N_3369,N_3669);
nor U4701 (N_4701,N_3724,N_3409);
nand U4702 (N_4702,N_3902,N_3652);
nor U4703 (N_4703,N_3001,N_3097);
and U4704 (N_4704,N_3088,N_3110);
and U4705 (N_4705,N_3600,N_3432);
and U4706 (N_4706,N_3652,N_3630);
or U4707 (N_4707,N_3995,N_3087);
nand U4708 (N_4708,N_3689,N_3561);
or U4709 (N_4709,N_3678,N_3513);
nand U4710 (N_4710,N_3224,N_3790);
or U4711 (N_4711,N_3208,N_3943);
and U4712 (N_4712,N_3491,N_3160);
nand U4713 (N_4713,N_3411,N_3640);
nand U4714 (N_4714,N_3578,N_3629);
nand U4715 (N_4715,N_3077,N_3117);
xor U4716 (N_4716,N_3972,N_3407);
and U4717 (N_4717,N_3814,N_3515);
nor U4718 (N_4718,N_3042,N_3322);
or U4719 (N_4719,N_3791,N_3498);
or U4720 (N_4720,N_3737,N_3543);
nand U4721 (N_4721,N_3497,N_3450);
and U4722 (N_4722,N_3804,N_3063);
nor U4723 (N_4723,N_3856,N_3481);
nand U4724 (N_4724,N_3237,N_3789);
xnor U4725 (N_4725,N_3917,N_3969);
and U4726 (N_4726,N_3526,N_3091);
nand U4727 (N_4727,N_3392,N_3757);
and U4728 (N_4728,N_3220,N_3414);
or U4729 (N_4729,N_3189,N_3562);
or U4730 (N_4730,N_3689,N_3956);
or U4731 (N_4731,N_3009,N_3363);
nor U4732 (N_4732,N_3087,N_3589);
nand U4733 (N_4733,N_3254,N_3225);
nand U4734 (N_4734,N_3008,N_3813);
and U4735 (N_4735,N_3378,N_3344);
nand U4736 (N_4736,N_3290,N_3755);
or U4737 (N_4737,N_3410,N_3493);
or U4738 (N_4738,N_3095,N_3945);
and U4739 (N_4739,N_3266,N_3864);
xnor U4740 (N_4740,N_3084,N_3469);
and U4741 (N_4741,N_3261,N_3427);
nand U4742 (N_4742,N_3989,N_3434);
nor U4743 (N_4743,N_3120,N_3660);
nor U4744 (N_4744,N_3892,N_3279);
and U4745 (N_4745,N_3704,N_3238);
and U4746 (N_4746,N_3589,N_3137);
or U4747 (N_4747,N_3225,N_3557);
or U4748 (N_4748,N_3817,N_3975);
nand U4749 (N_4749,N_3770,N_3534);
nor U4750 (N_4750,N_3939,N_3348);
nor U4751 (N_4751,N_3670,N_3514);
and U4752 (N_4752,N_3938,N_3488);
nand U4753 (N_4753,N_3354,N_3657);
and U4754 (N_4754,N_3687,N_3728);
or U4755 (N_4755,N_3955,N_3518);
or U4756 (N_4756,N_3150,N_3157);
and U4757 (N_4757,N_3556,N_3955);
or U4758 (N_4758,N_3156,N_3841);
and U4759 (N_4759,N_3154,N_3760);
nand U4760 (N_4760,N_3787,N_3823);
nand U4761 (N_4761,N_3854,N_3114);
nor U4762 (N_4762,N_3491,N_3303);
nor U4763 (N_4763,N_3135,N_3864);
and U4764 (N_4764,N_3151,N_3589);
nand U4765 (N_4765,N_3419,N_3205);
nor U4766 (N_4766,N_3411,N_3873);
xnor U4767 (N_4767,N_3697,N_3016);
nand U4768 (N_4768,N_3829,N_3404);
nor U4769 (N_4769,N_3581,N_3329);
and U4770 (N_4770,N_3903,N_3220);
nand U4771 (N_4771,N_3579,N_3527);
nand U4772 (N_4772,N_3508,N_3105);
or U4773 (N_4773,N_3482,N_3615);
and U4774 (N_4774,N_3160,N_3744);
nand U4775 (N_4775,N_3603,N_3626);
and U4776 (N_4776,N_3361,N_3091);
nand U4777 (N_4777,N_3066,N_3224);
nand U4778 (N_4778,N_3933,N_3696);
nand U4779 (N_4779,N_3945,N_3566);
and U4780 (N_4780,N_3178,N_3990);
or U4781 (N_4781,N_3124,N_3693);
nor U4782 (N_4782,N_3670,N_3055);
or U4783 (N_4783,N_3790,N_3647);
or U4784 (N_4784,N_3298,N_3086);
nand U4785 (N_4785,N_3724,N_3834);
nor U4786 (N_4786,N_3986,N_3308);
or U4787 (N_4787,N_3340,N_3614);
nand U4788 (N_4788,N_3615,N_3078);
and U4789 (N_4789,N_3594,N_3735);
or U4790 (N_4790,N_3808,N_3939);
nor U4791 (N_4791,N_3580,N_3936);
nand U4792 (N_4792,N_3676,N_3670);
and U4793 (N_4793,N_3003,N_3243);
or U4794 (N_4794,N_3679,N_3936);
nand U4795 (N_4795,N_3938,N_3212);
nand U4796 (N_4796,N_3531,N_3565);
nand U4797 (N_4797,N_3308,N_3059);
and U4798 (N_4798,N_3576,N_3852);
or U4799 (N_4799,N_3759,N_3078);
nor U4800 (N_4800,N_3792,N_3576);
nand U4801 (N_4801,N_3191,N_3709);
nand U4802 (N_4802,N_3065,N_3310);
nor U4803 (N_4803,N_3936,N_3106);
or U4804 (N_4804,N_3814,N_3454);
nor U4805 (N_4805,N_3297,N_3838);
and U4806 (N_4806,N_3764,N_3616);
and U4807 (N_4807,N_3404,N_3719);
nand U4808 (N_4808,N_3421,N_3602);
nand U4809 (N_4809,N_3841,N_3433);
nor U4810 (N_4810,N_3023,N_3664);
nand U4811 (N_4811,N_3234,N_3814);
nand U4812 (N_4812,N_3888,N_3810);
nor U4813 (N_4813,N_3719,N_3320);
or U4814 (N_4814,N_3890,N_3282);
nand U4815 (N_4815,N_3270,N_3242);
and U4816 (N_4816,N_3700,N_3825);
nand U4817 (N_4817,N_3426,N_3786);
nand U4818 (N_4818,N_3755,N_3302);
and U4819 (N_4819,N_3571,N_3232);
or U4820 (N_4820,N_3277,N_3449);
and U4821 (N_4821,N_3215,N_3070);
nor U4822 (N_4822,N_3660,N_3049);
or U4823 (N_4823,N_3074,N_3347);
or U4824 (N_4824,N_3831,N_3606);
nand U4825 (N_4825,N_3898,N_3975);
and U4826 (N_4826,N_3584,N_3675);
nor U4827 (N_4827,N_3351,N_3271);
nor U4828 (N_4828,N_3927,N_3846);
and U4829 (N_4829,N_3772,N_3765);
nor U4830 (N_4830,N_3006,N_3497);
nand U4831 (N_4831,N_3524,N_3407);
nor U4832 (N_4832,N_3640,N_3187);
xnor U4833 (N_4833,N_3079,N_3058);
and U4834 (N_4834,N_3813,N_3445);
xor U4835 (N_4835,N_3165,N_3029);
and U4836 (N_4836,N_3959,N_3049);
or U4837 (N_4837,N_3099,N_3000);
nand U4838 (N_4838,N_3734,N_3853);
or U4839 (N_4839,N_3602,N_3269);
or U4840 (N_4840,N_3090,N_3625);
nor U4841 (N_4841,N_3436,N_3057);
nand U4842 (N_4842,N_3762,N_3672);
nor U4843 (N_4843,N_3522,N_3927);
nand U4844 (N_4844,N_3683,N_3390);
or U4845 (N_4845,N_3958,N_3598);
and U4846 (N_4846,N_3212,N_3975);
and U4847 (N_4847,N_3120,N_3725);
nor U4848 (N_4848,N_3939,N_3565);
nor U4849 (N_4849,N_3368,N_3718);
and U4850 (N_4850,N_3644,N_3120);
and U4851 (N_4851,N_3725,N_3834);
and U4852 (N_4852,N_3701,N_3760);
nand U4853 (N_4853,N_3971,N_3515);
nor U4854 (N_4854,N_3959,N_3512);
and U4855 (N_4855,N_3036,N_3609);
or U4856 (N_4856,N_3353,N_3990);
nand U4857 (N_4857,N_3832,N_3522);
nor U4858 (N_4858,N_3500,N_3550);
or U4859 (N_4859,N_3640,N_3033);
nor U4860 (N_4860,N_3170,N_3898);
nor U4861 (N_4861,N_3567,N_3032);
nor U4862 (N_4862,N_3417,N_3087);
nor U4863 (N_4863,N_3302,N_3136);
and U4864 (N_4864,N_3062,N_3680);
nand U4865 (N_4865,N_3784,N_3173);
and U4866 (N_4866,N_3144,N_3675);
nor U4867 (N_4867,N_3214,N_3424);
nand U4868 (N_4868,N_3057,N_3427);
or U4869 (N_4869,N_3840,N_3663);
or U4870 (N_4870,N_3686,N_3413);
nand U4871 (N_4871,N_3497,N_3951);
nor U4872 (N_4872,N_3555,N_3536);
or U4873 (N_4873,N_3607,N_3883);
nand U4874 (N_4874,N_3423,N_3927);
and U4875 (N_4875,N_3218,N_3920);
nand U4876 (N_4876,N_3405,N_3617);
and U4877 (N_4877,N_3901,N_3452);
nand U4878 (N_4878,N_3907,N_3366);
or U4879 (N_4879,N_3319,N_3900);
nor U4880 (N_4880,N_3571,N_3017);
or U4881 (N_4881,N_3391,N_3893);
nor U4882 (N_4882,N_3040,N_3586);
nor U4883 (N_4883,N_3665,N_3790);
and U4884 (N_4884,N_3016,N_3977);
nor U4885 (N_4885,N_3239,N_3983);
nor U4886 (N_4886,N_3342,N_3955);
nor U4887 (N_4887,N_3312,N_3587);
nand U4888 (N_4888,N_3603,N_3206);
nand U4889 (N_4889,N_3136,N_3077);
or U4890 (N_4890,N_3249,N_3486);
or U4891 (N_4891,N_3314,N_3437);
nor U4892 (N_4892,N_3973,N_3187);
and U4893 (N_4893,N_3843,N_3761);
nand U4894 (N_4894,N_3360,N_3832);
and U4895 (N_4895,N_3743,N_3922);
xor U4896 (N_4896,N_3796,N_3445);
or U4897 (N_4897,N_3917,N_3257);
nand U4898 (N_4898,N_3313,N_3693);
or U4899 (N_4899,N_3390,N_3499);
nor U4900 (N_4900,N_3550,N_3544);
and U4901 (N_4901,N_3844,N_3728);
nand U4902 (N_4902,N_3960,N_3671);
or U4903 (N_4903,N_3981,N_3598);
nor U4904 (N_4904,N_3307,N_3637);
and U4905 (N_4905,N_3596,N_3421);
nand U4906 (N_4906,N_3016,N_3952);
nand U4907 (N_4907,N_3880,N_3863);
nand U4908 (N_4908,N_3976,N_3721);
and U4909 (N_4909,N_3883,N_3593);
nand U4910 (N_4910,N_3002,N_3334);
or U4911 (N_4911,N_3038,N_3450);
nand U4912 (N_4912,N_3365,N_3512);
or U4913 (N_4913,N_3868,N_3988);
or U4914 (N_4914,N_3891,N_3673);
nor U4915 (N_4915,N_3580,N_3290);
nor U4916 (N_4916,N_3350,N_3863);
nor U4917 (N_4917,N_3357,N_3706);
or U4918 (N_4918,N_3583,N_3912);
or U4919 (N_4919,N_3918,N_3113);
and U4920 (N_4920,N_3241,N_3306);
nand U4921 (N_4921,N_3019,N_3247);
nand U4922 (N_4922,N_3761,N_3488);
and U4923 (N_4923,N_3261,N_3271);
and U4924 (N_4924,N_3579,N_3151);
or U4925 (N_4925,N_3388,N_3309);
or U4926 (N_4926,N_3998,N_3344);
or U4927 (N_4927,N_3017,N_3198);
and U4928 (N_4928,N_3529,N_3639);
and U4929 (N_4929,N_3730,N_3348);
nand U4930 (N_4930,N_3563,N_3091);
or U4931 (N_4931,N_3298,N_3990);
nor U4932 (N_4932,N_3213,N_3731);
or U4933 (N_4933,N_3063,N_3977);
or U4934 (N_4934,N_3472,N_3710);
or U4935 (N_4935,N_3924,N_3769);
and U4936 (N_4936,N_3625,N_3870);
nand U4937 (N_4937,N_3779,N_3882);
xnor U4938 (N_4938,N_3703,N_3701);
or U4939 (N_4939,N_3621,N_3202);
or U4940 (N_4940,N_3948,N_3381);
nand U4941 (N_4941,N_3211,N_3671);
nand U4942 (N_4942,N_3725,N_3074);
and U4943 (N_4943,N_3307,N_3130);
nand U4944 (N_4944,N_3369,N_3167);
nand U4945 (N_4945,N_3888,N_3113);
or U4946 (N_4946,N_3004,N_3301);
and U4947 (N_4947,N_3114,N_3588);
or U4948 (N_4948,N_3300,N_3521);
and U4949 (N_4949,N_3454,N_3986);
nor U4950 (N_4950,N_3436,N_3034);
nand U4951 (N_4951,N_3705,N_3305);
or U4952 (N_4952,N_3257,N_3945);
or U4953 (N_4953,N_3531,N_3614);
or U4954 (N_4954,N_3058,N_3149);
nand U4955 (N_4955,N_3484,N_3517);
nor U4956 (N_4956,N_3986,N_3779);
nand U4957 (N_4957,N_3288,N_3187);
and U4958 (N_4958,N_3656,N_3949);
nand U4959 (N_4959,N_3904,N_3590);
nor U4960 (N_4960,N_3482,N_3725);
and U4961 (N_4961,N_3430,N_3616);
and U4962 (N_4962,N_3859,N_3644);
nand U4963 (N_4963,N_3138,N_3915);
or U4964 (N_4964,N_3835,N_3699);
and U4965 (N_4965,N_3298,N_3325);
or U4966 (N_4966,N_3004,N_3382);
or U4967 (N_4967,N_3276,N_3230);
and U4968 (N_4968,N_3405,N_3218);
and U4969 (N_4969,N_3146,N_3489);
nor U4970 (N_4970,N_3828,N_3506);
or U4971 (N_4971,N_3303,N_3317);
nand U4972 (N_4972,N_3884,N_3976);
nor U4973 (N_4973,N_3991,N_3182);
or U4974 (N_4974,N_3369,N_3765);
nor U4975 (N_4975,N_3054,N_3379);
nor U4976 (N_4976,N_3462,N_3149);
or U4977 (N_4977,N_3814,N_3474);
nand U4978 (N_4978,N_3856,N_3371);
nand U4979 (N_4979,N_3145,N_3372);
or U4980 (N_4980,N_3060,N_3274);
nand U4981 (N_4981,N_3290,N_3570);
or U4982 (N_4982,N_3952,N_3541);
and U4983 (N_4983,N_3336,N_3576);
nand U4984 (N_4984,N_3952,N_3454);
or U4985 (N_4985,N_3643,N_3513);
nor U4986 (N_4986,N_3825,N_3194);
or U4987 (N_4987,N_3831,N_3410);
or U4988 (N_4988,N_3014,N_3349);
and U4989 (N_4989,N_3987,N_3048);
and U4990 (N_4990,N_3088,N_3283);
and U4991 (N_4991,N_3792,N_3072);
nand U4992 (N_4992,N_3294,N_3571);
and U4993 (N_4993,N_3948,N_3413);
nand U4994 (N_4994,N_3512,N_3159);
nor U4995 (N_4995,N_3113,N_3611);
and U4996 (N_4996,N_3509,N_3091);
and U4997 (N_4997,N_3541,N_3171);
nor U4998 (N_4998,N_3722,N_3392);
nor U4999 (N_4999,N_3387,N_3360);
nand U5000 (N_5000,N_4206,N_4706);
and U5001 (N_5001,N_4750,N_4988);
nor U5002 (N_5002,N_4529,N_4942);
and U5003 (N_5003,N_4082,N_4471);
or U5004 (N_5004,N_4943,N_4397);
nand U5005 (N_5005,N_4044,N_4455);
nor U5006 (N_5006,N_4899,N_4910);
or U5007 (N_5007,N_4317,N_4609);
and U5008 (N_5008,N_4945,N_4782);
nand U5009 (N_5009,N_4733,N_4885);
nand U5010 (N_5010,N_4353,N_4540);
nand U5011 (N_5011,N_4081,N_4032);
and U5012 (N_5012,N_4647,N_4523);
xor U5013 (N_5013,N_4475,N_4739);
or U5014 (N_5014,N_4230,N_4664);
or U5015 (N_5015,N_4777,N_4967);
or U5016 (N_5016,N_4846,N_4793);
nor U5017 (N_5017,N_4993,N_4510);
and U5018 (N_5018,N_4209,N_4274);
or U5019 (N_5019,N_4221,N_4096);
and U5020 (N_5020,N_4227,N_4610);
and U5021 (N_5021,N_4045,N_4040);
nor U5022 (N_5022,N_4173,N_4662);
nand U5023 (N_5023,N_4047,N_4603);
or U5024 (N_5024,N_4421,N_4524);
or U5025 (N_5025,N_4054,N_4228);
and U5026 (N_5026,N_4727,N_4002);
or U5027 (N_5027,N_4550,N_4406);
or U5028 (N_5028,N_4607,N_4242);
nand U5029 (N_5029,N_4426,N_4888);
and U5030 (N_5030,N_4407,N_4290);
nor U5031 (N_5031,N_4578,N_4494);
nand U5032 (N_5032,N_4181,N_4629);
nor U5033 (N_5033,N_4011,N_4861);
nor U5034 (N_5034,N_4215,N_4346);
nor U5035 (N_5035,N_4724,N_4157);
nand U5036 (N_5036,N_4229,N_4222);
or U5037 (N_5037,N_4612,N_4763);
and U5038 (N_5038,N_4464,N_4369);
nor U5039 (N_5039,N_4370,N_4050);
and U5040 (N_5040,N_4863,N_4444);
nand U5041 (N_5041,N_4994,N_4488);
and U5042 (N_5042,N_4218,N_4594);
nor U5043 (N_5043,N_4087,N_4357);
nand U5044 (N_5044,N_4907,N_4768);
nand U5045 (N_5045,N_4261,N_4252);
nor U5046 (N_5046,N_4666,N_4984);
nor U5047 (N_5047,N_4283,N_4693);
or U5048 (N_5048,N_4841,N_4869);
and U5049 (N_5049,N_4920,N_4364);
nor U5050 (N_5050,N_4122,N_4792);
nand U5051 (N_5051,N_4385,N_4311);
and U5052 (N_5052,N_4915,N_4095);
and U5053 (N_5053,N_4005,N_4536);
nor U5054 (N_5054,N_4534,N_4022);
nor U5055 (N_5055,N_4258,N_4403);
or U5056 (N_5056,N_4618,N_4198);
or U5057 (N_5057,N_4580,N_4518);
nand U5058 (N_5058,N_4485,N_4375);
nor U5059 (N_5059,N_4889,N_4966);
nor U5060 (N_5060,N_4744,N_4960);
nand U5061 (N_5061,N_4249,N_4587);
and U5062 (N_5062,N_4619,N_4756);
or U5063 (N_5063,N_4731,N_4588);
nand U5064 (N_5064,N_4884,N_4527);
or U5065 (N_5065,N_4279,N_4876);
and U5066 (N_5066,N_4093,N_4710);
nand U5067 (N_5067,N_4663,N_4977);
nor U5068 (N_5068,N_4162,N_4103);
and U5069 (N_5069,N_4320,N_4288);
and U5070 (N_5070,N_4097,N_4453);
nand U5071 (N_5071,N_4965,N_4018);
or U5072 (N_5072,N_4029,N_4199);
and U5073 (N_5073,N_4454,N_4189);
nor U5074 (N_5074,N_4027,N_4037);
nand U5075 (N_5075,N_4718,N_4380);
nand U5076 (N_5076,N_4055,N_4246);
nor U5077 (N_5077,N_4061,N_4735);
or U5078 (N_5078,N_4428,N_4312);
nor U5079 (N_5079,N_4676,N_4887);
nor U5080 (N_5080,N_4979,N_4091);
nand U5081 (N_5081,N_4741,N_4234);
or U5082 (N_5082,N_4668,N_4470);
nand U5083 (N_5083,N_4056,N_4952);
nor U5084 (N_5084,N_4650,N_4682);
or U5085 (N_5085,N_4345,N_4704);
and U5086 (N_5086,N_4220,N_4784);
nand U5087 (N_5087,N_4197,N_4009);
nand U5088 (N_5088,N_4975,N_4113);
nand U5089 (N_5089,N_4673,N_4694);
nor U5090 (N_5090,N_4467,N_4561);
nor U5091 (N_5091,N_4131,N_4275);
and U5092 (N_5092,N_4382,N_4900);
nand U5093 (N_5093,N_4505,N_4543);
or U5094 (N_5094,N_4124,N_4719);
nor U5095 (N_5095,N_4203,N_4882);
nand U5096 (N_5096,N_4867,N_4812);
and U5097 (N_5097,N_4086,N_4277);
xor U5098 (N_5098,N_4624,N_4962);
or U5099 (N_5099,N_4526,N_4504);
and U5100 (N_5100,N_4049,N_4384);
or U5101 (N_5101,N_4102,N_4716);
and U5102 (N_5102,N_4310,N_4796);
or U5103 (N_5103,N_4707,N_4123);
or U5104 (N_5104,N_4502,N_4946);
nor U5105 (N_5105,N_4099,N_4699);
nand U5106 (N_5106,N_4951,N_4469);
nand U5107 (N_5107,N_4630,N_4348);
or U5108 (N_5108,N_4150,N_4373);
nand U5109 (N_5109,N_4649,N_4094);
nand U5110 (N_5110,N_4964,N_4268);
nand U5111 (N_5111,N_4155,N_4287);
nand U5112 (N_5112,N_4438,N_4423);
xnor U5113 (N_5113,N_4387,N_4414);
nand U5114 (N_5114,N_4970,N_4680);
and U5115 (N_5115,N_4713,N_4922);
and U5116 (N_5116,N_4341,N_4466);
or U5117 (N_5117,N_4273,N_4686);
nor U5118 (N_5118,N_4814,N_4521);
nor U5119 (N_5119,N_4519,N_4323);
nor U5120 (N_5120,N_4795,N_4271);
nor U5121 (N_5121,N_4765,N_4759);
and U5122 (N_5122,N_4703,N_4245);
nand U5123 (N_5123,N_4877,N_4826);
nand U5124 (N_5124,N_4358,N_4180);
and U5125 (N_5125,N_4642,N_4685);
nor U5126 (N_5126,N_4304,N_4168);
or U5127 (N_5127,N_4278,N_4210);
and U5128 (N_5128,N_4544,N_4016);
xor U5129 (N_5129,N_4672,N_4657);
nor U5130 (N_5130,N_4963,N_4762);
or U5131 (N_5131,N_4798,N_4591);
or U5132 (N_5132,N_4912,N_4169);
nor U5133 (N_5133,N_4042,N_4194);
nor U5134 (N_5134,N_4506,N_4794);
nor U5135 (N_5135,N_4282,N_4146);
or U5136 (N_5136,N_4003,N_4939);
nor U5137 (N_5137,N_4542,N_4462);
or U5138 (N_5138,N_4441,N_4213);
nand U5139 (N_5139,N_4626,N_4625);
and U5140 (N_5140,N_4916,N_4377);
or U5141 (N_5141,N_4605,N_4092);
nor U5142 (N_5142,N_4669,N_4190);
nand U5143 (N_5143,N_4745,N_4247);
or U5144 (N_5144,N_4257,N_4381);
or U5145 (N_5145,N_4886,N_4151);
and U5146 (N_5146,N_4412,N_4995);
and U5147 (N_5147,N_4742,N_4868);
and U5148 (N_5148,N_4374,N_4390);
and U5149 (N_5149,N_4422,N_4065);
nor U5150 (N_5150,N_4319,N_4827);
nor U5151 (N_5151,N_4138,N_4493);
and U5152 (N_5152,N_4064,N_4976);
or U5153 (N_5153,N_4949,N_4060);
and U5154 (N_5154,N_4262,N_4959);
nand U5155 (N_5155,N_4326,N_4844);
and U5156 (N_5156,N_4001,N_4328);
and U5157 (N_5157,N_4327,N_4557);
xor U5158 (N_5158,N_4145,N_4191);
nand U5159 (N_5159,N_4276,N_4058);
or U5160 (N_5160,N_4108,N_4458);
and U5161 (N_5161,N_4683,N_4452);
nand U5162 (N_5162,N_4919,N_4817);
nand U5163 (N_5163,N_4950,N_4986);
nand U5164 (N_5164,N_4871,N_4205);
nand U5165 (N_5165,N_4646,N_4280);
or U5166 (N_5166,N_4818,N_4532);
or U5167 (N_5167,N_4007,N_4971);
nor U5168 (N_5168,N_4039,N_4985);
nand U5169 (N_5169,N_4581,N_4656);
nand U5170 (N_5170,N_4072,N_4350);
nor U5171 (N_5171,N_4803,N_4677);
and U5172 (N_5172,N_4417,N_4116);
or U5173 (N_5173,N_4243,N_4398);
and U5174 (N_5174,N_4926,N_4335);
nor U5175 (N_5175,N_4324,N_4478);
or U5176 (N_5176,N_4315,N_4297);
and U5177 (N_5177,N_4204,N_4430);
or U5178 (N_5178,N_4434,N_4017);
and U5179 (N_5179,N_4879,N_4689);
and U5180 (N_5180,N_4235,N_4025);
nor U5181 (N_5181,N_4165,N_4176);
nor U5182 (N_5182,N_4780,N_4259);
nand U5183 (N_5183,N_4309,N_4331);
and U5184 (N_5184,N_4779,N_4063);
nand U5185 (N_5185,N_4177,N_4495);
nand U5186 (N_5186,N_4643,N_4752);
or U5187 (N_5187,N_4034,N_4142);
and U5188 (N_5188,N_4820,N_4823);
nand U5189 (N_5189,N_4300,N_4582);
and U5190 (N_5190,N_4256,N_4171);
or U5191 (N_5191,N_4507,N_4313);
nand U5192 (N_5192,N_4571,N_4559);
or U5193 (N_5193,N_4847,N_4289);
or U5194 (N_5194,N_4109,N_4957);
nand U5195 (N_5195,N_4244,N_4723);
and U5196 (N_5196,N_4130,N_4178);
or U5197 (N_5197,N_4264,N_4447);
nor U5198 (N_5198,N_4681,N_4404);
or U5199 (N_5199,N_4816,N_4878);
and U5200 (N_5200,N_4248,N_4751);
nand U5201 (N_5201,N_4314,N_4562);
or U5202 (N_5202,N_4875,N_4574);
or U5203 (N_5203,N_4365,N_4084);
nor U5204 (N_5204,N_4254,N_4648);
nor U5205 (N_5205,N_4567,N_4391);
nand U5206 (N_5206,N_4355,N_4940);
and U5207 (N_5207,N_4321,N_4590);
and U5208 (N_5208,N_4987,N_4859);
nor U5209 (N_5209,N_4435,N_4400);
nor U5210 (N_5210,N_4183,N_4698);
or U5211 (N_5211,N_4990,N_4267);
nand U5212 (N_5212,N_4708,N_4896);
or U5213 (N_5213,N_4376,N_4476);
or U5214 (N_5214,N_4424,N_4316);
or U5215 (N_5215,N_4132,N_4338);
and U5216 (N_5216,N_4974,N_4790);
and U5217 (N_5217,N_4738,N_4757);
and U5218 (N_5218,N_4905,N_4644);
or U5219 (N_5219,N_4748,N_4651);
or U5220 (N_5220,N_4163,N_4051);
nand U5221 (N_5221,N_4490,N_4786);
or U5222 (N_5222,N_4208,N_4645);
nand U5223 (N_5223,N_4457,N_4831);
or U5224 (N_5224,N_4613,N_4783);
and U5225 (N_5225,N_4773,N_4539);
nor U5226 (N_5226,N_4491,N_4127);
and U5227 (N_5227,N_4969,N_4764);
nor U5228 (N_5228,N_4860,N_4895);
and U5229 (N_5229,N_4356,N_4849);
and U5230 (N_5230,N_4460,N_4118);
or U5231 (N_5231,N_4632,N_4892);
and U5232 (N_5232,N_4968,N_4568);
and U5233 (N_5233,N_4909,N_4941);
nor U5234 (N_5234,N_4448,N_4715);
and U5235 (N_5235,N_4620,N_4720);
nand U5236 (N_5236,N_4921,N_4137);
nor U5237 (N_5237,N_4269,N_4822);
nor U5238 (N_5238,N_4425,N_4069);
and U5239 (N_5239,N_4658,N_4956);
and U5240 (N_5240,N_4351,N_4639);
nor U5241 (N_5241,N_4484,N_4486);
and U5242 (N_5242,N_4272,N_4537);
and U5243 (N_5243,N_4419,N_4545);
nor U5244 (N_5244,N_4325,N_4894);
nor U5245 (N_5245,N_4563,N_4201);
nand U5246 (N_5246,N_4931,N_4501);
nand U5247 (N_5247,N_4980,N_4927);
or U5248 (N_5248,N_4347,N_4429);
or U5249 (N_5249,N_4890,N_4083);
and U5250 (N_5250,N_4797,N_4695);
and U5251 (N_5251,N_4004,N_4548);
and U5252 (N_5252,N_4405,N_4824);
or U5253 (N_5253,N_4932,N_4013);
and U5254 (N_5254,N_4936,N_4667);
or U5255 (N_5255,N_4641,N_4593);
nand U5256 (N_5256,N_4866,N_4726);
nand U5257 (N_5257,N_4378,N_4174);
nor U5258 (N_5258,N_4498,N_4697);
nor U5259 (N_5259,N_4600,N_4508);
nand U5260 (N_5260,N_4547,N_4730);
nor U5261 (N_5261,N_4874,N_4306);
or U5262 (N_5262,N_4046,N_4813);
nand U5263 (N_5263,N_4688,N_4333);
and U5264 (N_5264,N_4788,N_4520);
nor U5265 (N_5265,N_4660,N_4217);
or U5266 (N_5266,N_4253,N_4829);
or U5267 (N_5267,N_4802,N_4074);
nor U5268 (N_5268,N_4608,N_4237);
and U5269 (N_5269,N_4166,N_4515);
nor U5270 (N_5270,N_4158,N_4010);
nor U5271 (N_5271,N_4621,N_4184);
nor U5272 (N_5272,N_4477,N_4635);
nand U5273 (N_5273,N_4395,N_4778);
nand U5274 (N_5274,N_4791,N_4251);
nor U5275 (N_5275,N_4599,N_4839);
or U5276 (N_5276,N_4804,N_4755);
and U5277 (N_5277,N_4585,N_4000);
nand U5278 (N_5278,N_4020,N_4615);
nand U5279 (N_5279,N_4893,N_4767);
nand U5280 (N_5280,N_4935,N_4053);
nor U5281 (N_5281,N_4120,N_4821);
and U5282 (N_5282,N_4800,N_4554);
nor U5283 (N_5283,N_4512,N_4579);
or U5284 (N_5284,N_4517,N_4904);
nor U5285 (N_5285,N_4670,N_4690);
nand U5286 (N_5286,N_4308,N_4700);
and U5287 (N_5287,N_4442,N_4528);
or U5288 (N_5288,N_4701,N_4570);
and U5289 (N_5289,N_4807,N_4024);
nand U5290 (N_5290,N_4775,N_4446);
nor U5291 (N_5291,N_4451,N_4634);
and U5292 (N_5292,N_4908,N_4611);
nor U5293 (N_5293,N_4903,N_4129);
and U5294 (N_5294,N_4553,N_4100);
nand U5295 (N_5295,N_4292,N_4073);
or U5296 (N_5296,N_4255,N_4622);
nand U5297 (N_5297,N_4911,N_4115);
nor U5298 (N_5298,N_4972,N_4617);
nand U5299 (N_5299,N_4872,N_4787);
or U5300 (N_5300,N_4810,N_4705);
nand U5301 (N_5301,N_4164,N_4367);
nor U5302 (N_5302,N_4525,N_4891);
nor U5303 (N_5303,N_4427,N_4147);
and U5304 (N_5304,N_4339,N_4873);
nand U5305 (N_5305,N_4354,N_4396);
nor U5306 (N_5306,N_4696,N_4898);
and U5307 (N_5307,N_4152,N_4533);
and U5308 (N_5308,N_4068,N_4728);
and U5309 (N_5309,N_4575,N_4709);
and U5310 (N_5310,N_4363,N_4474);
or U5311 (N_5311,N_4433,N_4413);
nor U5312 (N_5312,N_4006,N_4989);
nor U5313 (N_5313,N_4322,N_4743);
or U5314 (N_5314,N_4776,N_4855);
nor U5315 (N_5315,N_4125,N_4144);
or U5316 (N_5316,N_4854,N_4233);
or U5317 (N_5317,N_4106,N_4602);
or U5318 (N_5318,N_4489,N_4981);
nand U5319 (N_5319,N_4806,N_4296);
nand U5320 (N_5320,N_4511,N_4436);
nor U5321 (N_5321,N_4577,N_4241);
nand U5322 (N_5322,N_4026,N_4437);
or U5323 (N_5323,N_4606,N_4837);
and U5324 (N_5324,N_4295,N_4172);
and U5325 (N_5325,N_4461,N_4573);
or U5326 (N_5326,N_4937,N_4953);
nand U5327 (N_5327,N_4389,N_4415);
and U5328 (N_5328,N_4535,N_4850);
nand U5329 (N_5329,N_4134,N_4770);
or U5330 (N_5330,N_4913,N_4736);
and U5331 (N_5331,N_4598,N_4117);
nand U5332 (N_5332,N_4114,N_4352);
or U5333 (N_5333,N_4028,N_4923);
or U5334 (N_5334,N_4361,N_4133);
nor U5335 (N_5335,N_4684,N_4263);
and U5336 (N_5336,N_4774,N_4088);
nand U5337 (N_5337,N_4388,N_4769);
nor U5338 (N_5338,N_4303,N_4362);
and U5339 (N_5339,N_4809,N_4307);
or U5340 (N_5340,N_4075,N_4604);
nor U5341 (N_5341,N_4214,N_4572);
nand U5342 (N_5342,N_4336,N_4500);
nand U5343 (N_5343,N_4048,N_4465);
or U5344 (N_5344,N_4149,N_4678);
nor U5345 (N_5345,N_4182,N_4071);
nor U5346 (N_5346,N_4337,N_4958);
nand U5347 (N_5347,N_4298,N_4401);
nor U5348 (N_5348,N_4631,N_4196);
or U5349 (N_5349,N_4586,N_4140);
nand U5350 (N_5350,N_4418,N_4250);
nand U5351 (N_5351,N_4193,N_4239);
and U5352 (N_5352,N_4819,N_4760);
nand U5353 (N_5353,N_4785,N_4556);
nand U5354 (N_5354,N_4749,N_4012);
and U5355 (N_5355,N_4443,N_4514);
and U5356 (N_5356,N_4293,N_4111);
or U5357 (N_5357,N_4973,N_4754);
or U5358 (N_5358,N_4030,N_4901);
nand U5359 (N_5359,N_4496,N_4240);
nor U5360 (N_5360,N_4232,N_4432);
nand U5361 (N_5361,N_4212,N_4070);
or U5362 (N_5362,N_4549,N_4772);
or U5363 (N_5363,N_4179,N_4789);
nand U5364 (N_5364,N_4035,N_4801);
nand U5365 (N_5365,N_4623,N_4207);
nor U5366 (N_5366,N_4136,N_4799);
and U5367 (N_5367,N_4480,N_4483);
nor U5368 (N_5368,N_4948,N_4153);
nor U5369 (N_5369,N_4997,N_4566);
nand U5370 (N_5370,N_4954,N_4052);
or U5371 (N_5371,N_4286,N_4638);
nor U5372 (N_5372,N_4552,N_4342);
and U5373 (N_5373,N_4815,N_4654);
and U5374 (N_5374,N_4947,N_4747);
nor U5375 (N_5375,N_4918,N_4104);
nand U5376 (N_5376,N_4781,N_4080);
nand U5377 (N_5377,N_4360,N_4349);
nand U5378 (N_5378,N_4692,N_4862);
and U5379 (N_5379,N_4019,N_4226);
nor U5380 (N_5380,N_4301,N_4479);
nand U5381 (N_5381,N_4126,N_4858);
nor U5382 (N_5382,N_4712,N_4408);
nor U5383 (N_5383,N_4564,N_4085);
and U5384 (N_5384,N_4597,N_4431);
nor U5385 (N_5385,N_4661,N_4961);
nand U5386 (N_5386,N_4805,N_4679);
and U5387 (N_5387,N_4729,N_4601);
and U5388 (N_5388,N_4595,N_4031);
nand U5389 (N_5389,N_4238,N_4934);
and U5390 (N_5390,N_4659,N_4671);
nand U5391 (N_5391,N_4231,N_4291);
nor U5392 (N_5392,N_4456,N_4546);
and U5393 (N_5393,N_4721,N_4655);
nand U5394 (N_5394,N_4864,N_4897);
nor U5395 (N_5395,N_4033,N_4192);
and U5396 (N_5396,N_4285,N_4038);
xnor U5397 (N_5397,N_4516,N_4852);
or U5398 (N_5398,N_4522,N_4833);
nor U5399 (N_5399,N_4420,N_4691);
nor U5400 (N_5400,N_4170,N_4856);
nand U5401 (N_5401,N_4021,N_4996);
and U5402 (N_5402,N_4383,N_4284);
or U5403 (N_5403,N_4834,N_4265);
nor U5404 (N_5404,N_4141,N_4260);
nand U5405 (N_5405,N_4737,N_4808);
and U5406 (N_5406,N_4848,N_4998);
and U5407 (N_5407,N_4880,N_4687);
or U5408 (N_5408,N_4513,N_4665);
nor U5409 (N_5409,N_4497,N_4105);
and U5410 (N_5410,N_4386,N_4371);
nand U5411 (N_5411,N_4637,N_4583);
or U5412 (N_5412,N_4825,N_4991);
or U5413 (N_5413,N_4565,N_4343);
nor U5414 (N_5414,N_4299,N_4740);
nor U5415 (N_5415,N_4558,N_4023);
and U5416 (N_5416,N_4098,N_4481);
or U5417 (N_5417,N_4128,N_4368);
nand U5418 (N_5418,N_4938,N_4175);
or U5419 (N_5419,N_4928,N_4392);
or U5420 (N_5420,N_4836,N_4186);
or U5421 (N_5421,N_4394,N_4714);
nor U5422 (N_5422,N_4416,N_4592);
or U5423 (N_5423,N_4236,N_4902);
and U5424 (N_5424,N_4154,N_4842);
or U5425 (N_5425,N_4090,N_4541);
nor U5426 (N_5426,N_4076,N_4211);
and U5427 (N_5427,N_4223,N_4062);
nand U5428 (N_5428,N_4857,N_4627);
nor U5429 (N_5429,N_4982,N_4569);
nand U5430 (N_5430,N_4944,N_4924);
nor U5431 (N_5431,N_4851,N_4294);
nor U5432 (N_5432,N_4077,N_4187);
and U5433 (N_5433,N_4188,N_4161);
nor U5434 (N_5434,N_4036,N_4402);
or U5435 (N_5435,N_4459,N_4933);
nand U5436 (N_5436,N_4761,N_4576);
nor U5437 (N_5437,N_4066,N_4992);
or U5438 (N_5438,N_4616,N_4143);
or U5439 (N_5439,N_4318,N_4482);
and U5440 (N_5440,N_4633,N_4393);
nand U5441 (N_5441,N_4121,N_4925);
nor U5442 (N_5442,N_4359,N_4509);
nor U5443 (N_5443,N_4445,N_4119);
or U5444 (N_5444,N_4200,N_4135);
or U5445 (N_5445,N_4725,N_4555);
nand U5446 (N_5446,N_4881,N_4159);
and U5447 (N_5447,N_4139,N_4530);
or U5448 (N_5448,N_4266,N_4487);
nor U5449 (N_5449,N_4840,N_4379);
and U5450 (N_5450,N_4057,N_4409);
nor U5451 (N_5451,N_4440,N_4329);
nor U5452 (N_5452,N_4828,N_4883);
and U5453 (N_5453,N_4472,N_4766);
and U5454 (N_5454,N_4835,N_4185);
nor U5455 (N_5455,N_4195,N_4281);
and U5456 (N_5456,N_4499,N_4732);
and U5457 (N_5457,N_4929,N_4640);
nor U5458 (N_5458,N_4399,N_4584);
nor U5459 (N_5459,N_4302,N_4830);
and U5460 (N_5460,N_4439,N_4330);
nor U5461 (N_5461,N_4079,N_4372);
nand U5462 (N_5462,N_4332,N_4219);
nand U5463 (N_5463,N_4473,N_4628);
and U5464 (N_5464,N_4838,N_4110);
or U5465 (N_5465,N_4845,N_4078);
or U5466 (N_5466,N_4334,N_4832);
or U5467 (N_5467,N_4955,N_4156);
or U5468 (N_5468,N_4717,N_4450);
nand U5469 (N_5469,N_4906,N_4538);
and U5470 (N_5470,N_4652,N_4043);
or U5471 (N_5471,N_4059,N_4224);
or U5472 (N_5472,N_4216,N_4107);
or U5473 (N_5473,N_4148,N_4589);
or U5474 (N_5474,N_4674,N_4914);
or U5475 (N_5475,N_4999,N_4225);
nand U5476 (N_5476,N_4853,N_4089);
nand U5477 (N_5477,N_4160,N_4411);
nand U5478 (N_5478,N_4410,N_4983);
or U5479 (N_5479,N_4978,N_4917);
and U5480 (N_5480,N_4008,N_4758);
and U5481 (N_5481,N_4112,N_4653);
and U5482 (N_5482,N_4041,N_4101);
and U5483 (N_5483,N_4843,N_4865);
nor U5484 (N_5484,N_4551,N_4531);
nand U5485 (N_5485,N_4870,N_4636);
or U5486 (N_5486,N_4305,N_4202);
nand U5487 (N_5487,N_4930,N_4614);
or U5488 (N_5488,N_4702,N_4463);
nor U5489 (N_5489,N_4015,N_4492);
nand U5490 (N_5490,N_4468,N_4734);
nand U5491 (N_5491,N_4067,N_4449);
and U5492 (N_5492,N_4675,N_4811);
nor U5493 (N_5493,N_4503,N_4753);
or U5494 (N_5494,N_4270,N_4596);
or U5495 (N_5495,N_4711,N_4560);
nor U5496 (N_5496,N_4344,N_4167);
or U5497 (N_5497,N_4722,N_4746);
and U5498 (N_5498,N_4014,N_4340);
or U5499 (N_5499,N_4366,N_4771);
nor U5500 (N_5500,N_4843,N_4270);
nand U5501 (N_5501,N_4145,N_4690);
and U5502 (N_5502,N_4151,N_4235);
or U5503 (N_5503,N_4914,N_4448);
nand U5504 (N_5504,N_4827,N_4167);
and U5505 (N_5505,N_4409,N_4461);
and U5506 (N_5506,N_4967,N_4077);
nor U5507 (N_5507,N_4421,N_4158);
xor U5508 (N_5508,N_4616,N_4523);
or U5509 (N_5509,N_4886,N_4281);
or U5510 (N_5510,N_4763,N_4657);
and U5511 (N_5511,N_4880,N_4104);
and U5512 (N_5512,N_4087,N_4052);
and U5513 (N_5513,N_4849,N_4450);
nand U5514 (N_5514,N_4146,N_4254);
nand U5515 (N_5515,N_4863,N_4517);
or U5516 (N_5516,N_4587,N_4151);
nor U5517 (N_5517,N_4417,N_4235);
and U5518 (N_5518,N_4723,N_4183);
or U5519 (N_5519,N_4994,N_4071);
nor U5520 (N_5520,N_4138,N_4715);
nor U5521 (N_5521,N_4146,N_4907);
nor U5522 (N_5522,N_4656,N_4174);
nand U5523 (N_5523,N_4906,N_4748);
or U5524 (N_5524,N_4334,N_4765);
or U5525 (N_5525,N_4761,N_4307);
and U5526 (N_5526,N_4082,N_4877);
nor U5527 (N_5527,N_4377,N_4487);
nand U5528 (N_5528,N_4560,N_4940);
or U5529 (N_5529,N_4625,N_4531);
or U5530 (N_5530,N_4464,N_4043);
or U5531 (N_5531,N_4639,N_4902);
nor U5532 (N_5532,N_4067,N_4804);
or U5533 (N_5533,N_4135,N_4024);
and U5534 (N_5534,N_4439,N_4889);
nor U5535 (N_5535,N_4120,N_4125);
and U5536 (N_5536,N_4991,N_4364);
and U5537 (N_5537,N_4779,N_4524);
nand U5538 (N_5538,N_4331,N_4274);
nor U5539 (N_5539,N_4051,N_4892);
or U5540 (N_5540,N_4785,N_4234);
or U5541 (N_5541,N_4696,N_4799);
nor U5542 (N_5542,N_4119,N_4816);
or U5543 (N_5543,N_4159,N_4201);
and U5544 (N_5544,N_4092,N_4837);
or U5545 (N_5545,N_4578,N_4473);
and U5546 (N_5546,N_4575,N_4181);
and U5547 (N_5547,N_4193,N_4634);
nor U5548 (N_5548,N_4735,N_4901);
or U5549 (N_5549,N_4380,N_4965);
nor U5550 (N_5550,N_4750,N_4079);
and U5551 (N_5551,N_4921,N_4327);
and U5552 (N_5552,N_4680,N_4600);
and U5553 (N_5553,N_4562,N_4446);
nor U5554 (N_5554,N_4439,N_4847);
nor U5555 (N_5555,N_4644,N_4810);
nor U5556 (N_5556,N_4736,N_4512);
and U5557 (N_5557,N_4352,N_4081);
or U5558 (N_5558,N_4538,N_4059);
and U5559 (N_5559,N_4367,N_4748);
and U5560 (N_5560,N_4590,N_4633);
nor U5561 (N_5561,N_4699,N_4718);
nor U5562 (N_5562,N_4181,N_4983);
nand U5563 (N_5563,N_4199,N_4930);
nand U5564 (N_5564,N_4525,N_4263);
nand U5565 (N_5565,N_4956,N_4423);
and U5566 (N_5566,N_4737,N_4335);
or U5567 (N_5567,N_4245,N_4293);
or U5568 (N_5568,N_4491,N_4072);
nor U5569 (N_5569,N_4859,N_4206);
nor U5570 (N_5570,N_4050,N_4085);
nand U5571 (N_5571,N_4726,N_4350);
nor U5572 (N_5572,N_4786,N_4992);
nand U5573 (N_5573,N_4501,N_4508);
nor U5574 (N_5574,N_4462,N_4560);
and U5575 (N_5575,N_4357,N_4441);
nand U5576 (N_5576,N_4484,N_4946);
and U5577 (N_5577,N_4731,N_4958);
and U5578 (N_5578,N_4858,N_4992);
and U5579 (N_5579,N_4192,N_4358);
nand U5580 (N_5580,N_4077,N_4043);
nor U5581 (N_5581,N_4830,N_4185);
or U5582 (N_5582,N_4174,N_4925);
and U5583 (N_5583,N_4468,N_4934);
nor U5584 (N_5584,N_4970,N_4451);
and U5585 (N_5585,N_4710,N_4815);
nor U5586 (N_5586,N_4194,N_4157);
or U5587 (N_5587,N_4176,N_4216);
nand U5588 (N_5588,N_4652,N_4878);
or U5589 (N_5589,N_4341,N_4975);
nor U5590 (N_5590,N_4453,N_4037);
nand U5591 (N_5591,N_4162,N_4688);
nand U5592 (N_5592,N_4651,N_4148);
and U5593 (N_5593,N_4392,N_4043);
or U5594 (N_5594,N_4538,N_4851);
nand U5595 (N_5595,N_4155,N_4980);
nand U5596 (N_5596,N_4293,N_4373);
or U5597 (N_5597,N_4410,N_4671);
nand U5598 (N_5598,N_4220,N_4753);
nor U5599 (N_5599,N_4307,N_4385);
nor U5600 (N_5600,N_4651,N_4928);
nand U5601 (N_5601,N_4534,N_4685);
and U5602 (N_5602,N_4692,N_4670);
nor U5603 (N_5603,N_4521,N_4286);
or U5604 (N_5604,N_4449,N_4778);
nand U5605 (N_5605,N_4346,N_4411);
nand U5606 (N_5606,N_4937,N_4588);
or U5607 (N_5607,N_4674,N_4152);
nor U5608 (N_5608,N_4266,N_4317);
nand U5609 (N_5609,N_4997,N_4789);
nor U5610 (N_5610,N_4293,N_4916);
nor U5611 (N_5611,N_4746,N_4204);
nor U5612 (N_5612,N_4531,N_4142);
or U5613 (N_5613,N_4377,N_4008);
nor U5614 (N_5614,N_4485,N_4926);
and U5615 (N_5615,N_4386,N_4841);
nor U5616 (N_5616,N_4144,N_4070);
and U5617 (N_5617,N_4594,N_4452);
or U5618 (N_5618,N_4257,N_4338);
and U5619 (N_5619,N_4648,N_4101);
nand U5620 (N_5620,N_4943,N_4571);
and U5621 (N_5621,N_4230,N_4073);
or U5622 (N_5622,N_4212,N_4053);
nor U5623 (N_5623,N_4860,N_4304);
or U5624 (N_5624,N_4822,N_4198);
or U5625 (N_5625,N_4817,N_4956);
nor U5626 (N_5626,N_4800,N_4750);
nor U5627 (N_5627,N_4339,N_4782);
nor U5628 (N_5628,N_4480,N_4797);
and U5629 (N_5629,N_4092,N_4068);
and U5630 (N_5630,N_4068,N_4146);
or U5631 (N_5631,N_4832,N_4695);
nor U5632 (N_5632,N_4032,N_4255);
nor U5633 (N_5633,N_4661,N_4253);
and U5634 (N_5634,N_4248,N_4312);
or U5635 (N_5635,N_4662,N_4674);
nor U5636 (N_5636,N_4539,N_4909);
and U5637 (N_5637,N_4852,N_4033);
and U5638 (N_5638,N_4675,N_4301);
nand U5639 (N_5639,N_4464,N_4091);
nor U5640 (N_5640,N_4408,N_4744);
nand U5641 (N_5641,N_4341,N_4981);
nor U5642 (N_5642,N_4163,N_4626);
nor U5643 (N_5643,N_4938,N_4643);
nand U5644 (N_5644,N_4763,N_4407);
and U5645 (N_5645,N_4754,N_4550);
or U5646 (N_5646,N_4547,N_4321);
nor U5647 (N_5647,N_4721,N_4378);
nand U5648 (N_5648,N_4046,N_4755);
nor U5649 (N_5649,N_4871,N_4129);
nand U5650 (N_5650,N_4666,N_4588);
or U5651 (N_5651,N_4836,N_4592);
and U5652 (N_5652,N_4322,N_4548);
or U5653 (N_5653,N_4947,N_4578);
nor U5654 (N_5654,N_4874,N_4579);
or U5655 (N_5655,N_4167,N_4553);
nor U5656 (N_5656,N_4630,N_4993);
and U5657 (N_5657,N_4303,N_4549);
or U5658 (N_5658,N_4537,N_4656);
nand U5659 (N_5659,N_4806,N_4083);
nand U5660 (N_5660,N_4970,N_4078);
nand U5661 (N_5661,N_4125,N_4463);
and U5662 (N_5662,N_4073,N_4777);
nor U5663 (N_5663,N_4260,N_4591);
nand U5664 (N_5664,N_4937,N_4041);
or U5665 (N_5665,N_4133,N_4308);
and U5666 (N_5666,N_4990,N_4158);
and U5667 (N_5667,N_4849,N_4741);
nand U5668 (N_5668,N_4445,N_4942);
and U5669 (N_5669,N_4864,N_4942);
or U5670 (N_5670,N_4047,N_4596);
nor U5671 (N_5671,N_4847,N_4923);
nand U5672 (N_5672,N_4713,N_4266);
nand U5673 (N_5673,N_4435,N_4888);
nand U5674 (N_5674,N_4569,N_4697);
xnor U5675 (N_5675,N_4046,N_4220);
and U5676 (N_5676,N_4971,N_4795);
nand U5677 (N_5677,N_4423,N_4271);
or U5678 (N_5678,N_4842,N_4386);
and U5679 (N_5679,N_4292,N_4962);
and U5680 (N_5680,N_4356,N_4765);
and U5681 (N_5681,N_4645,N_4649);
or U5682 (N_5682,N_4420,N_4793);
nand U5683 (N_5683,N_4529,N_4741);
or U5684 (N_5684,N_4409,N_4758);
nand U5685 (N_5685,N_4178,N_4318);
or U5686 (N_5686,N_4830,N_4809);
nand U5687 (N_5687,N_4002,N_4968);
nand U5688 (N_5688,N_4856,N_4956);
or U5689 (N_5689,N_4651,N_4920);
or U5690 (N_5690,N_4961,N_4906);
nand U5691 (N_5691,N_4117,N_4651);
or U5692 (N_5692,N_4291,N_4856);
nand U5693 (N_5693,N_4224,N_4099);
nor U5694 (N_5694,N_4861,N_4333);
nand U5695 (N_5695,N_4775,N_4800);
nor U5696 (N_5696,N_4008,N_4178);
or U5697 (N_5697,N_4206,N_4634);
and U5698 (N_5698,N_4203,N_4876);
or U5699 (N_5699,N_4091,N_4189);
and U5700 (N_5700,N_4180,N_4704);
and U5701 (N_5701,N_4274,N_4609);
nor U5702 (N_5702,N_4592,N_4771);
nor U5703 (N_5703,N_4401,N_4752);
nand U5704 (N_5704,N_4724,N_4495);
and U5705 (N_5705,N_4690,N_4938);
or U5706 (N_5706,N_4917,N_4599);
or U5707 (N_5707,N_4428,N_4918);
nand U5708 (N_5708,N_4164,N_4441);
and U5709 (N_5709,N_4929,N_4363);
nand U5710 (N_5710,N_4126,N_4887);
nand U5711 (N_5711,N_4941,N_4288);
and U5712 (N_5712,N_4194,N_4152);
nor U5713 (N_5713,N_4620,N_4637);
nor U5714 (N_5714,N_4362,N_4673);
nand U5715 (N_5715,N_4967,N_4430);
and U5716 (N_5716,N_4572,N_4281);
xnor U5717 (N_5717,N_4839,N_4912);
nor U5718 (N_5718,N_4803,N_4217);
nor U5719 (N_5719,N_4871,N_4657);
nor U5720 (N_5720,N_4407,N_4946);
nor U5721 (N_5721,N_4209,N_4392);
nor U5722 (N_5722,N_4814,N_4417);
or U5723 (N_5723,N_4347,N_4405);
nor U5724 (N_5724,N_4535,N_4033);
and U5725 (N_5725,N_4952,N_4226);
and U5726 (N_5726,N_4926,N_4015);
and U5727 (N_5727,N_4134,N_4346);
nor U5728 (N_5728,N_4719,N_4341);
or U5729 (N_5729,N_4657,N_4981);
and U5730 (N_5730,N_4497,N_4932);
nor U5731 (N_5731,N_4882,N_4172);
nand U5732 (N_5732,N_4494,N_4330);
nor U5733 (N_5733,N_4862,N_4713);
nand U5734 (N_5734,N_4404,N_4053);
or U5735 (N_5735,N_4646,N_4835);
or U5736 (N_5736,N_4058,N_4839);
and U5737 (N_5737,N_4301,N_4166);
and U5738 (N_5738,N_4510,N_4432);
or U5739 (N_5739,N_4923,N_4767);
or U5740 (N_5740,N_4487,N_4698);
nand U5741 (N_5741,N_4598,N_4571);
and U5742 (N_5742,N_4362,N_4217);
or U5743 (N_5743,N_4877,N_4830);
nor U5744 (N_5744,N_4034,N_4315);
nor U5745 (N_5745,N_4559,N_4804);
nor U5746 (N_5746,N_4972,N_4712);
and U5747 (N_5747,N_4153,N_4425);
nor U5748 (N_5748,N_4525,N_4316);
nor U5749 (N_5749,N_4512,N_4642);
nand U5750 (N_5750,N_4918,N_4702);
and U5751 (N_5751,N_4661,N_4660);
nor U5752 (N_5752,N_4877,N_4226);
nor U5753 (N_5753,N_4855,N_4725);
nor U5754 (N_5754,N_4093,N_4798);
nor U5755 (N_5755,N_4646,N_4505);
and U5756 (N_5756,N_4123,N_4851);
and U5757 (N_5757,N_4626,N_4437);
nand U5758 (N_5758,N_4706,N_4951);
nor U5759 (N_5759,N_4164,N_4186);
nor U5760 (N_5760,N_4045,N_4274);
nand U5761 (N_5761,N_4618,N_4588);
or U5762 (N_5762,N_4022,N_4880);
and U5763 (N_5763,N_4450,N_4804);
and U5764 (N_5764,N_4791,N_4694);
nor U5765 (N_5765,N_4284,N_4456);
nor U5766 (N_5766,N_4666,N_4380);
nand U5767 (N_5767,N_4676,N_4830);
nor U5768 (N_5768,N_4668,N_4949);
or U5769 (N_5769,N_4757,N_4957);
nor U5770 (N_5770,N_4356,N_4446);
or U5771 (N_5771,N_4411,N_4317);
nor U5772 (N_5772,N_4789,N_4534);
nor U5773 (N_5773,N_4970,N_4763);
and U5774 (N_5774,N_4481,N_4492);
and U5775 (N_5775,N_4651,N_4324);
nor U5776 (N_5776,N_4997,N_4758);
nand U5777 (N_5777,N_4005,N_4355);
nand U5778 (N_5778,N_4845,N_4335);
and U5779 (N_5779,N_4625,N_4234);
or U5780 (N_5780,N_4782,N_4419);
nand U5781 (N_5781,N_4311,N_4258);
nand U5782 (N_5782,N_4268,N_4936);
and U5783 (N_5783,N_4797,N_4824);
or U5784 (N_5784,N_4462,N_4312);
and U5785 (N_5785,N_4213,N_4336);
nor U5786 (N_5786,N_4327,N_4379);
nor U5787 (N_5787,N_4041,N_4856);
nand U5788 (N_5788,N_4036,N_4077);
nor U5789 (N_5789,N_4233,N_4324);
or U5790 (N_5790,N_4599,N_4995);
and U5791 (N_5791,N_4667,N_4796);
nor U5792 (N_5792,N_4298,N_4756);
nand U5793 (N_5793,N_4658,N_4886);
nand U5794 (N_5794,N_4641,N_4190);
nand U5795 (N_5795,N_4977,N_4414);
xor U5796 (N_5796,N_4235,N_4419);
nand U5797 (N_5797,N_4691,N_4577);
and U5798 (N_5798,N_4281,N_4349);
or U5799 (N_5799,N_4749,N_4180);
nor U5800 (N_5800,N_4755,N_4359);
nor U5801 (N_5801,N_4547,N_4989);
nand U5802 (N_5802,N_4390,N_4363);
nand U5803 (N_5803,N_4906,N_4014);
nor U5804 (N_5804,N_4555,N_4497);
or U5805 (N_5805,N_4330,N_4561);
nand U5806 (N_5806,N_4175,N_4498);
and U5807 (N_5807,N_4937,N_4548);
and U5808 (N_5808,N_4564,N_4715);
nand U5809 (N_5809,N_4481,N_4027);
nand U5810 (N_5810,N_4108,N_4666);
nor U5811 (N_5811,N_4227,N_4707);
nand U5812 (N_5812,N_4699,N_4028);
nor U5813 (N_5813,N_4618,N_4703);
nand U5814 (N_5814,N_4032,N_4339);
nor U5815 (N_5815,N_4362,N_4265);
and U5816 (N_5816,N_4461,N_4649);
or U5817 (N_5817,N_4335,N_4603);
nand U5818 (N_5818,N_4764,N_4292);
and U5819 (N_5819,N_4202,N_4078);
nand U5820 (N_5820,N_4393,N_4205);
nor U5821 (N_5821,N_4647,N_4331);
nor U5822 (N_5822,N_4526,N_4088);
nand U5823 (N_5823,N_4311,N_4504);
nand U5824 (N_5824,N_4372,N_4185);
or U5825 (N_5825,N_4783,N_4265);
nand U5826 (N_5826,N_4203,N_4182);
nand U5827 (N_5827,N_4489,N_4236);
and U5828 (N_5828,N_4337,N_4194);
and U5829 (N_5829,N_4029,N_4059);
or U5830 (N_5830,N_4635,N_4670);
xnor U5831 (N_5831,N_4040,N_4116);
and U5832 (N_5832,N_4182,N_4168);
nor U5833 (N_5833,N_4618,N_4405);
or U5834 (N_5834,N_4491,N_4560);
and U5835 (N_5835,N_4421,N_4366);
nand U5836 (N_5836,N_4481,N_4710);
or U5837 (N_5837,N_4286,N_4249);
or U5838 (N_5838,N_4677,N_4648);
nand U5839 (N_5839,N_4102,N_4985);
or U5840 (N_5840,N_4156,N_4487);
nand U5841 (N_5841,N_4443,N_4269);
nor U5842 (N_5842,N_4705,N_4415);
or U5843 (N_5843,N_4664,N_4580);
or U5844 (N_5844,N_4524,N_4623);
nor U5845 (N_5845,N_4171,N_4799);
nand U5846 (N_5846,N_4513,N_4271);
and U5847 (N_5847,N_4709,N_4555);
nand U5848 (N_5848,N_4267,N_4483);
or U5849 (N_5849,N_4425,N_4841);
nand U5850 (N_5850,N_4434,N_4856);
nor U5851 (N_5851,N_4503,N_4584);
nor U5852 (N_5852,N_4062,N_4783);
nor U5853 (N_5853,N_4424,N_4307);
or U5854 (N_5854,N_4177,N_4458);
nor U5855 (N_5855,N_4659,N_4150);
or U5856 (N_5856,N_4632,N_4272);
and U5857 (N_5857,N_4446,N_4746);
nor U5858 (N_5858,N_4210,N_4664);
nor U5859 (N_5859,N_4169,N_4298);
nand U5860 (N_5860,N_4869,N_4146);
and U5861 (N_5861,N_4445,N_4795);
or U5862 (N_5862,N_4405,N_4600);
or U5863 (N_5863,N_4570,N_4954);
and U5864 (N_5864,N_4898,N_4859);
nand U5865 (N_5865,N_4305,N_4178);
and U5866 (N_5866,N_4462,N_4072);
and U5867 (N_5867,N_4628,N_4501);
or U5868 (N_5868,N_4735,N_4290);
and U5869 (N_5869,N_4405,N_4525);
and U5870 (N_5870,N_4573,N_4487);
nand U5871 (N_5871,N_4773,N_4219);
nand U5872 (N_5872,N_4328,N_4469);
and U5873 (N_5873,N_4374,N_4874);
nor U5874 (N_5874,N_4070,N_4295);
and U5875 (N_5875,N_4539,N_4574);
nand U5876 (N_5876,N_4160,N_4322);
nand U5877 (N_5877,N_4686,N_4736);
nand U5878 (N_5878,N_4663,N_4399);
nand U5879 (N_5879,N_4637,N_4767);
nand U5880 (N_5880,N_4157,N_4637);
nand U5881 (N_5881,N_4348,N_4227);
nand U5882 (N_5882,N_4030,N_4207);
nor U5883 (N_5883,N_4957,N_4479);
nand U5884 (N_5884,N_4400,N_4004);
nor U5885 (N_5885,N_4457,N_4486);
nor U5886 (N_5886,N_4431,N_4717);
nand U5887 (N_5887,N_4859,N_4481);
nand U5888 (N_5888,N_4953,N_4711);
nor U5889 (N_5889,N_4214,N_4267);
nand U5890 (N_5890,N_4672,N_4280);
or U5891 (N_5891,N_4602,N_4337);
nand U5892 (N_5892,N_4699,N_4156);
xor U5893 (N_5893,N_4933,N_4080);
nand U5894 (N_5894,N_4306,N_4001);
nor U5895 (N_5895,N_4583,N_4440);
nand U5896 (N_5896,N_4848,N_4302);
and U5897 (N_5897,N_4057,N_4728);
nor U5898 (N_5898,N_4266,N_4192);
nand U5899 (N_5899,N_4086,N_4258);
nor U5900 (N_5900,N_4870,N_4442);
or U5901 (N_5901,N_4672,N_4736);
nor U5902 (N_5902,N_4117,N_4278);
nand U5903 (N_5903,N_4599,N_4224);
nand U5904 (N_5904,N_4307,N_4263);
and U5905 (N_5905,N_4699,N_4914);
and U5906 (N_5906,N_4945,N_4919);
or U5907 (N_5907,N_4115,N_4461);
and U5908 (N_5908,N_4162,N_4825);
and U5909 (N_5909,N_4387,N_4793);
and U5910 (N_5910,N_4366,N_4794);
nand U5911 (N_5911,N_4228,N_4834);
nand U5912 (N_5912,N_4164,N_4655);
and U5913 (N_5913,N_4740,N_4855);
nand U5914 (N_5914,N_4190,N_4790);
nor U5915 (N_5915,N_4799,N_4166);
nand U5916 (N_5916,N_4802,N_4851);
nor U5917 (N_5917,N_4767,N_4689);
nand U5918 (N_5918,N_4865,N_4560);
and U5919 (N_5919,N_4778,N_4643);
and U5920 (N_5920,N_4263,N_4047);
and U5921 (N_5921,N_4607,N_4058);
nand U5922 (N_5922,N_4834,N_4778);
nor U5923 (N_5923,N_4429,N_4099);
nand U5924 (N_5924,N_4870,N_4679);
nor U5925 (N_5925,N_4674,N_4653);
and U5926 (N_5926,N_4403,N_4417);
and U5927 (N_5927,N_4526,N_4319);
and U5928 (N_5928,N_4596,N_4009);
and U5929 (N_5929,N_4987,N_4334);
nand U5930 (N_5930,N_4285,N_4161);
nor U5931 (N_5931,N_4512,N_4544);
nand U5932 (N_5932,N_4203,N_4041);
or U5933 (N_5933,N_4530,N_4075);
and U5934 (N_5934,N_4718,N_4580);
nor U5935 (N_5935,N_4461,N_4503);
nor U5936 (N_5936,N_4309,N_4827);
or U5937 (N_5937,N_4442,N_4851);
nand U5938 (N_5938,N_4232,N_4430);
and U5939 (N_5939,N_4235,N_4888);
nor U5940 (N_5940,N_4110,N_4709);
nor U5941 (N_5941,N_4493,N_4496);
nor U5942 (N_5942,N_4729,N_4310);
nor U5943 (N_5943,N_4892,N_4252);
nor U5944 (N_5944,N_4423,N_4042);
or U5945 (N_5945,N_4826,N_4441);
and U5946 (N_5946,N_4695,N_4295);
or U5947 (N_5947,N_4057,N_4989);
or U5948 (N_5948,N_4517,N_4258);
or U5949 (N_5949,N_4926,N_4937);
and U5950 (N_5950,N_4629,N_4045);
nand U5951 (N_5951,N_4969,N_4721);
or U5952 (N_5952,N_4584,N_4144);
or U5953 (N_5953,N_4335,N_4566);
or U5954 (N_5954,N_4551,N_4698);
or U5955 (N_5955,N_4952,N_4971);
or U5956 (N_5956,N_4925,N_4784);
nand U5957 (N_5957,N_4553,N_4894);
and U5958 (N_5958,N_4822,N_4013);
and U5959 (N_5959,N_4060,N_4847);
nand U5960 (N_5960,N_4378,N_4546);
nor U5961 (N_5961,N_4586,N_4194);
or U5962 (N_5962,N_4868,N_4535);
nand U5963 (N_5963,N_4253,N_4642);
nand U5964 (N_5964,N_4324,N_4038);
nor U5965 (N_5965,N_4595,N_4248);
nor U5966 (N_5966,N_4601,N_4528);
nor U5967 (N_5967,N_4216,N_4180);
or U5968 (N_5968,N_4089,N_4778);
or U5969 (N_5969,N_4261,N_4144);
and U5970 (N_5970,N_4732,N_4353);
or U5971 (N_5971,N_4697,N_4469);
nand U5972 (N_5972,N_4678,N_4920);
nor U5973 (N_5973,N_4420,N_4888);
nand U5974 (N_5974,N_4759,N_4906);
nand U5975 (N_5975,N_4444,N_4416);
or U5976 (N_5976,N_4516,N_4074);
nand U5977 (N_5977,N_4961,N_4753);
and U5978 (N_5978,N_4277,N_4222);
or U5979 (N_5979,N_4839,N_4796);
nand U5980 (N_5980,N_4179,N_4371);
and U5981 (N_5981,N_4274,N_4311);
or U5982 (N_5982,N_4047,N_4839);
nand U5983 (N_5983,N_4591,N_4278);
and U5984 (N_5984,N_4138,N_4353);
nor U5985 (N_5985,N_4314,N_4689);
nor U5986 (N_5986,N_4720,N_4264);
and U5987 (N_5987,N_4219,N_4996);
and U5988 (N_5988,N_4032,N_4688);
nand U5989 (N_5989,N_4884,N_4168);
and U5990 (N_5990,N_4864,N_4138);
and U5991 (N_5991,N_4699,N_4230);
nor U5992 (N_5992,N_4258,N_4796);
and U5993 (N_5993,N_4748,N_4160);
nand U5994 (N_5994,N_4233,N_4487);
and U5995 (N_5995,N_4202,N_4609);
and U5996 (N_5996,N_4130,N_4237);
and U5997 (N_5997,N_4607,N_4881);
or U5998 (N_5998,N_4261,N_4507);
nor U5999 (N_5999,N_4662,N_4444);
nand U6000 (N_6000,N_5778,N_5356);
or U6001 (N_6001,N_5655,N_5779);
and U6002 (N_6002,N_5208,N_5569);
nand U6003 (N_6003,N_5621,N_5534);
and U6004 (N_6004,N_5211,N_5343);
nor U6005 (N_6005,N_5338,N_5003);
or U6006 (N_6006,N_5784,N_5846);
nor U6007 (N_6007,N_5931,N_5812);
nand U6008 (N_6008,N_5600,N_5457);
or U6009 (N_6009,N_5976,N_5149);
and U6010 (N_6010,N_5521,N_5496);
and U6011 (N_6011,N_5929,N_5664);
nand U6012 (N_6012,N_5644,N_5725);
and U6013 (N_6013,N_5366,N_5728);
nand U6014 (N_6014,N_5167,N_5809);
and U6015 (N_6015,N_5394,N_5877);
or U6016 (N_6016,N_5363,N_5265);
nand U6017 (N_6017,N_5783,N_5381);
or U6018 (N_6018,N_5468,N_5276);
and U6019 (N_6019,N_5067,N_5515);
and U6020 (N_6020,N_5874,N_5080);
nand U6021 (N_6021,N_5190,N_5432);
or U6022 (N_6022,N_5486,N_5843);
xor U6023 (N_6023,N_5004,N_5596);
and U6024 (N_6024,N_5082,N_5593);
and U6025 (N_6025,N_5707,N_5449);
nor U6026 (N_6026,N_5665,N_5757);
and U6027 (N_6027,N_5337,N_5044);
or U6028 (N_6028,N_5415,N_5505);
nor U6029 (N_6029,N_5267,N_5735);
nor U6030 (N_6030,N_5698,N_5667);
and U6031 (N_6031,N_5446,N_5478);
nand U6032 (N_6032,N_5053,N_5632);
and U6033 (N_6033,N_5403,N_5856);
nand U6034 (N_6034,N_5933,N_5290);
or U6035 (N_6035,N_5409,N_5001);
nor U6036 (N_6036,N_5994,N_5558);
nor U6037 (N_6037,N_5300,N_5891);
nor U6038 (N_6038,N_5260,N_5752);
nor U6039 (N_6039,N_5225,N_5886);
and U6040 (N_6040,N_5477,N_5463);
and U6041 (N_6041,N_5304,N_5016);
and U6042 (N_6042,N_5714,N_5743);
nand U6043 (N_6043,N_5557,N_5883);
nand U6044 (N_6044,N_5148,N_5283);
nor U6045 (N_6045,N_5934,N_5209);
and U6046 (N_6046,N_5266,N_5835);
nor U6047 (N_6047,N_5199,N_5636);
or U6048 (N_6048,N_5316,N_5749);
or U6049 (N_6049,N_5972,N_5187);
nand U6050 (N_6050,N_5746,N_5969);
or U6051 (N_6051,N_5805,N_5269);
or U6052 (N_6052,N_5335,N_5135);
and U6053 (N_6053,N_5470,N_5639);
and U6054 (N_6054,N_5777,N_5120);
nor U6055 (N_6055,N_5516,N_5163);
or U6056 (N_6056,N_5560,N_5367);
nand U6057 (N_6057,N_5464,N_5890);
or U6058 (N_6058,N_5117,N_5832);
and U6059 (N_6059,N_5501,N_5045);
nor U6060 (N_6060,N_5176,N_5368);
nor U6061 (N_6061,N_5935,N_5207);
nor U6062 (N_6062,N_5105,N_5800);
nor U6063 (N_6063,N_5833,N_5005);
nor U6064 (N_6064,N_5303,N_5110);
nor U6065 (N_6065,N_5041,N_5906);
or U6066 (N_6066,N_5706,N_5022);
nand U6067 (N_6067,N_5161,N_5955);
or U6068 (N_6068,N_5490,N_5693);
or U6069 (N_6069,N_5370,N_5765);
or U6070 (N_6070,N_5766,N_5776);
nand U6071 (N_6071,N_5151,N_5197);
nand U6072 (N_6072,N_5093,N_5322);
nand U6073 (N_6073,N_5548,N_5499);
nor U6074 (N_6074,N_5503,N_5523);
or U6075 (N_6075,N_5459,N_5063);
and U6076 (N_6076,N_5851,N_5722);
nor U6077 (N_6077,N_5861,N_5084);
nor U6078 (N_6078,N_5065,N_5305);
and U6079 (N_6079,N_5658,N_5050);
or U6080 (N_6080,N_5231,N_5362);
and U6081 (N_6081,N_5940,N_5100);
or U6082 (N_6082,N_5221,N_5000);
nor U6083 (N_6083,N_5518,N_5307);
and U6084 (N_6084,N_5991,N_5302);
nand U6085 (N_6085,N_5326,N_5491);
or U6086 (N_6086,N_5237,N_5913);
nor U6087 (N_6087,N_5359,N_5530);
and U6088 (N_6088,N_5963,N_5713);
or U6089 (N_6089,N_5287,N_5150);
and U6090 (N_6090,N_5118,N_5026);
nand U6091 (N_6091,N_5819,N_5545);
nor U6092 (N_6092,N_5130,N_5182);
and U6093 (N_6093,N_5637,N_5426);
nor U6094 (N_6094,N_5971,N_5447);
nand U6095 (N_6095,N_5369,N_5576);
and U6096 (N_6096,N_5180,N_5660);
nor U6097 (N_6097,N_5482,N_5159);
nor U6098 (N_6098,N_5411,N_5358);
nor U6099 (N_6099,N_5919,N_5719);
or U6100 (N_6100,N_5618,N_5871);
nor U6101 (N_6101,N_5453,N_5932);
or U6102 (N_6102,N_5519,N_5444);
or U6103 (N_6103,N_5824,N_5382);
and U6104 (N_6104,N_5494,N_5755);
nor U6105 (N_6105,N_5248,N_5780);
or U6106 (N_6106,N_5608,N_5385);
or U6107 (N_6107,N_5537,N_5200);
nor U6108 (N_6108,N_5522,N_5051);
nor U6109 (N_6109,N_5244,N_5634);
nor U6110 (N_6110,N_5679,N_5448);
or U6111 (N_6111,N_5483,N_5028);
or U6112 (N_6112,N_5928,N_5690);
or U6113 (N_6113,N_5075,N_5256);
or U6114 (N_6114,N_5295,N_5320);
or U6115 (N_6115,N_5333,N_5625);
nor U6116 (N_6116,N_5195,N_5953);
or U6117 (N_6117,N_5344,N_5346);
and U6118 (N_6118,N_5327,N_5222);
nand U6119 (N_6119,N_5046,N_5823);
nor U6120 (N_6120,N_5708,N_5175);
nor U6121 (N_6121,N_5952,N_5774);
nor U6122 (N_6122,N_5592,N_5254);
nand U6123 (N_6123,N_5709,N_5471);
or U6124 (N_6124,N_5002,N_5628);
nor U6125 (N_6125,N_5853,N_5827);
nand U6126 (N_6126,N_5351,N_5390);
nor U6127 (N_6127,N_5830,N_5204);
and U6128 (N_6128,N_5021,N_5035);
and U6129 (N_6129,N_5297,N_5253);
or U6130 (N_6130,N_5443,N_5330);
nor U6131 (N_6131,N_5629,N_5810);
nor U6132 (N_6132,N_5980,N_5416);
xnor U6133 (N_6133,N_5506,N_5088);
or U6134 (N_6134,N_5631,N_5410);
nor U6135 (N_6135,N_5109,N_5252);
or U6136 (N_6136,N_5387,N_5349);
nor U6137 (N_6137,N_5179,N_5687);
nand U6138 (N_6138,N_5480,N_5122);
nand U6139 (N_6139,N_5077,N_5795);
or U6140 (N_6140,N_5609,N_5588);
and U6141 (N_6141,N_5828,N_5941);
nand U6142 (N_6142,N_5694,N_5087);
nand U6143 (N_6143,N_5060,N_5597);
and U6144 (N_6144,N_5128,N_5526);
nand U6145 (N_6145,N_5820,N_5651);
nor U6146 (N_6146,N_5570,N_5272);
and U6147 (N_6147,N_5845,N_5578);
and U6148 (N_6148,N_5927,N_5773);
or U6149 (N_6149,N_5884,N_5427);
nand U6150 (N_6150,N_5481,N_5691);
or U6151 (N_6151,N_5879,N_5170);
or U6152 (N_6152,N_5909,N_5900);
nand U6153 (N_6153,N_5603,N_5663);
and U6154 (N_6154,N_5323,N_5126);
or U6155 (N_6155,N_5798,N_5689);
and U6156 (N_6156,N_5371,N_5720);
or U6157 (N_6157,N_5716,N_5153);
or U6158 (N_6158,N_5852,N_5250);
or U6159 (N_6159,N_5177,N_5703);
and U6160 (N_6160,N_5113,N_5364);
xor U6161 (N_6161,N_5648,N_5699);
and U6162 (N_6162,N_5057,N_5577);
nor U6163 (N_6163,N_5069,N_5354);
and U6164 (N_6164,N_5990,N_5347);
nand U6165 (N_6165,N_5400,N_5575);
nand U6166 (N_6166,N_5702,N_5974);
nand U6167 (N_6167,N_5284,N_5194);
nand U6168 (N_6168,N_5997,N_5977);
nor U6169 (N_6169,N_5042,N_5393);
or U6170 (N_6170,N_5677,N_5676);
and U6171 (N_6171,N_5081,N_5762);
or U6172 (N_6172,N_5450,N_5073);
nand U6173 (N_6173,N_5383,N_5811);
and U6174 (N_6174,N_5642,N_5152);
nor U6175 (N_6175,N_5585,N_5350);
nand U6176 (N_6176,N_5924,N_5511);
nand U6177 (N_6177,N_5419,N_5888);
nand U6178 (N_6178,N_5988,N_5864);
or U6179 (N_6179,N_5547,N_5842);
or U6180 (N_6180,N_5581,N_5355);
or U6181 (N_6181,N_5684,N_5649);
nor U6182 (N_6182,N_5311,N_5761);
nor U6183 (N_6183,N_5860,N_5185);
nor U6184 (N_6184,N_5103,N_5285);
and U6185 (N_6185,N_5626,N_5544);
and U6186 (N_6186,N_5897,N_5227);
and U6187 (N_6187,N_5123,N_5034);
nor U6188 (N_6188,N_5741,N_5551);
nand U6189 (N_6189,N_5525,N_5907);
nand U6190 (N_6190,N_5959,N_5321);
and U6191 (N_6191,N_5580,N_5696);
nand U6192 (N_6192,N_5460,N_5881);
nor U6193 (N_6193,N_5198,N_5917);
nand U6194 (N_6194,N_5683,N_5561);
or U6195 (N_6195,N_5378,N_5859);
nor U6196 (N_6196,N_5492,N_5294);
nand U6197 (N_6197,N_5296,N_5033);
or U6198 (N_6198,N_5956,N_5674);
and U6199 (N_6199,N_5309,N_5498);
and U6200 (N_6200,N_5771,N_5539);
nor U6201 (N_6201,N_5858,N_5574);
nor U6202 (N_6202,N_5158,N_5524);
nand U6203 (N_6203,N_5220,N_5196);
nand U6204 (N_6204,N_5745,N_5388);
nand U6205 (N_6205,N_5174,N_5764);
nand U6206 (N_6206,N_5937,N_5226);
and U6207 (N_6207,N_5425,N_5454);
nor U6208 (N_6208,N_5509,N_5389);
xnor U6209 (N_6209,N_5587,N_5738);
and U6210 (N_6210,N_5873,N_5566);
and U6211 (N_6211,N_5930,N_5816);
nor U6212 (N_6212,N_5101,N_5132);
and U6213 (N_6213,N_5704,N_5062);
nand U6214 (N_6214,N_5656,N_5318);
or U6215 (N_6215,N_5939,N_5601);
nand U6216 (N_6216,N_5657,N_5513);
nand U6217 (N_6217,N_5882,N_5353);
and U6218 (N_6218,N_5280,N_5205);
or U6219 (N_6219,N_5943,N_5680);
and U6220 (N_6220,N_5815,N_5666);
nor U6221 (N_6221,N_5517,N_5301);
and U6222 (N_6222,N_5412,N_5633);
and U6223 (N_6223,N_5573,N_5386);
nor U6224 (N_6224,N_5023,N_5549);
and U6225 (N_6225,N_5408,N_5914);
nand U6226 (N_6226,N_5586,N_5831);
nand U6227 (N_6227,N_5944,N_5079);
nor U6228 (N_6228,N_5672,N_5405);
or U6229 (N_6229,N_5993,N_5155);
and U6230 (N_6230,N_5854,N_5512);
and U6231 (N_6231,N_5872,N_5781);
or U6232 (N_6232,N_5345,N_5214);
nand U6233 (N_6233,N_5989,N_5039);
xor U6234 (N_6234,N_5822,N_5911);
or U6235 (N_6235,N_5068,N_5992);
nand U6236 (N_6236,N_5291,N_5896);
or U6237 (N_6237,N_5750,N_5686);
nand U6238 (N_6238,N_5982,N_5893);
or U6239 (N_6239,N_5701,N_5133);
and U6240 (N_6240,N_5747,N_5869);
or U6241 (N_6241,N_5638,N_5726);
nand U6242 (N_6242,N_5641,N_5485);
and U6243 (N_6243,N_5475,N_5379);
nor U6244 (N_6244,N_5230,N_5406);
nand U6245 (N_6245,N_5685,N_5186);
nand U6246 (N_6246,N_5748,N_5462);
nor U6247 (N_6247,N_5908,N_5985);
or U6248 (N_6248,N_5712,N_5546);
or U6249 (N_6249,N_5912,N_5440);
nor U6250 (N_6250,N_5352,N_5404);
nor U6251 (N_6251,N_5692,N_5488);
and U6252 (N_6252,N_5098,N_5071);
nand U6253 (N_6253,N_5365,N_5675);
nor U6254 (N_6254,N_5834,N_5315);
nor U6255 (N_6255,N_5423,N_5792);
nor U6256 (N_6256,N_5754,N_5235);
nor U6257 (N_6257,N_5737,N_5555);
nand U6258 (N_6258,N_5863,N_5605);
and U6259 (N_6259,N_5620,N_5559);
and U6260 (N_6260,N_5962,N_5239);
nor U6261 (N_6261,N_5401,N_5553);
and U6262 (N_6262,N_5966,N_5849);
nor U6263 (N_6263,N_5348,N_5164);
or U6264 (N_6264,N_5829,N_5188);
or U6265 (N_6265,N_5855,N_5027);
or U6266 (N_6266,N_5430,N_5236);
nand U6267 (N_6267,N_5407,N_5903);
and U6268 (N_6268,N_5438,N_5115);
nor U6269 (N_6269,N_5247,N_5514);
nand U6270 (N_6270,N_5865,N_5589);
nor U6271 (N_6271,N_5808,N_5995);
nor U6272 (N_6272,N_5541,N_5172);
or U6273 (N_6273,N_5623,N_5616);
or U6274 (N_6274,N_5682,N_5157);
nor U6275 (N_6275,N_5329,N_5178);
nor U6276 (N_6276,N_5238,N_5218);
nor U6277 (N_6277,N_5528,N_5536);
xnor U6278 (N_6278,N_5251,N_5090);
nor U6279 (N_6279,N_5332,N_5504);
and U6280 (N_6280,N_5146,N_5759);
or U6281 (N_6281,N_5889,N_5261);
and U6282 (N_6282,N_5949,N_5718);
and U6283 (N_6283,N_5095,N_5184);
and U6284 (N_6284,N_5461,N_5905);
nand U6285 (N_6285,N_5210,N_5421);
and U6286 (N_6286,N_5019,N_5840);
or U6287 (N_6287,N_5607,N_5775);
nor U6288 (N_6288,N_5740,N_5173);
nor U6289 (N_6289,N_5769,N_5610);
or U6290 (N_6290,N_5978,N_5613);
and U6291 (N_6291,N_5328,N_5141);
nand U6292 (N_6292,N_5009,N_5011);
nor U6293 (N_6293,N_5531,N_5710);
nand U6294 (N_6294,N_5788,N_5466);
or U6295 (N_6295,N_5377,N_5627);
and U6296 (N_6296,N_5241,N_5880);
nand U6297 (N_6297,N_5894,N_5476);
and U6298 (N_6298,N_5850,N_5950);
nand U6299 (N_6299,N_5192,N_5552);
and U6300 (N_6300,N_5724,N_5671);
or U6301 (N_6301,N_5507,N_5030);
and U6302 (N_6302,N_5439,N_5617);
and U6303 (N_6303,N_5751,N_5271);
nand U6304 (N_6304,N_5255,N_5681);
nand U6305 (N_6305,N_5987,N_5233);
xor U6306 (N_6306,N_5313,N_5916);
nand U6307 (N_6307,N_5036,N_5785);
nor U6308 (N_6308,N_5138,N_5008);
or U6309 (N_6309,N_5437,N_5938);
and U6310 (N_6310,N_5054,N_5479);
and U6311 (N_6311,N_5422,N_5398);
nand U6312 (N_6312,N_5124,N_5020);
and U6313 (N_6313,N_5040,N_5533);
or U6314 (N_6314,N_5262,N_5467);
and U6315 (N_6315,N_5223,N_5535);
and U6316 (N_6316,N_5878,N_5844);
nor U6317 (N_6317,N_5331,N_5567);
and U6318 (N_6318,N_5431,N_5892);
nor U6319 (N_6319,N_5614,N_5787);
xor U6320 (N_6320,N_5540,N_5234);
nand U6321 (N_6321,N_5374,N_5984);
nand U6322 (N_6322,N_5837,N_5836);
nand U6323 (N_6323,N_5116,N_5797);
and U6324 (N_6324,N_5181,N_5038);
nand U6325 (N_6325,N_5274,N_5814);
and U6326 (N_6326,N_5670,N_5742);
nand U6327 (N_6327,N_5550,N_5895);
nand U6328 (N_6328,N_5455,N_5612);
or U6329 (N_6329,N_5145,N_5465);
or U6330 (N_6330,N_5538,N_5257);
nor U6331 (N_6331,N_5089,N_5495);
nor U6332 (N_6332,N_5072,N_5817);
nand U6333 (N_6333,N_5543,N_5286);
xnor U6334 (N_6334,N_5794,N_5074);
or U6335 (N_6335,N_5136,N_5862);
or U6336 (N_6336,N_5782,N_5695);
or U6337 (N_6337,N_5730,N_5076);
nor U6338 (N_6338,N_5583,N_5564);
and U6339 (N_6339,N_5847,N_5622);
nor U6340 (N_6340,N_5542,N_5424);
and U6341 (N_6341,N_5414,N_5242);
and U6342 (N_6342,N_5804,N_5213);
or U6343 (N_6343,N_5119,N_5868);
nand U6344 (N_6344,N_5129,N_5114);
nand U6345 (N_6345,N_5563,N_5012);
nand U6346 (N_6346,N_5606,N_5936);
and U6347 (N_6347,N_5434,N_5032);
nand U6348 (N_6348,N_5918,N_5973);
nor U6349 (N_6349,N_5014,N_5598);
or U6350 (N_6350,N_5711,N_5954);
nand U6351 (N_6351,N_5796,N_5996);
or U6352 (N_6352,N_5277,N_5529);
nand U6353 (N_6353,N_5314,N_5052);
nand U6354 (N_6354,N_5066,N_5139);
nor U6355 (N_6355,N_5160,N_5768);
or U6356 (N_6356,N_5127,N_5154);
nand U6357 (N_6357,N_5922,N_5733);
or U6358 (N_6358,N_5216,N_5212);
nor U6359 (N_6359,N_5169,N_5452);
and U6360 (N_6360,N_5336,N_5281);
or U6361 (N_6361,N_5981,N_5246);
and U6362 (N_6362,N_5380,N_5640);
nor U6363 (N_6363,N_5965,N_5224);
nor U6364 (N_6364,N_5571,N_5111);
or U6365 (N_6365,N_5064,N_5970);
nand U6366 (N_6366,N_5435,N_5801);
nor U6367 (N_6367,N_5920,N_5772);
nor U6368 (N_6368,N_5165,N_5968);
or U6369 (N_6369,N_5147,N_5334);
and U6370 (N_6370,N_5317,N_5442);
or U6371 (N_6371,N_5958,N_5556);
nor U6372 (N_6372,N_5156,N_5085);
and U6373 (N_6373,N_5292,N_5268);
or U6374 (N_6374,N_5899,N_5999);
and U6375 (N_6375,N_5669,N_5493);
and U6376 (N_6376,N_5700,N_5289);
nand U6377 (N_6377,N_5086,N_5018);
nor U6378 (N_6378,N_5705,N_5361);
or U6379 (N_6379,N_5029,N_5131);
nand U6380 (N_6380,N_5166,N_5789);
nor U6381 (N_6381,N_5373,N_5144);
nand U6382 (N_6382,N_5049,N_5191);
nand U6383 (N_6383,N_5125,N_5678);
nand U6384 (N_6384,N_5572,N_5715);
and U6385 (N_6385,N_5721,N_5661);
nand U6386 (N_6386,N_5171,N_5875);
and U6387 (N_6387,N_5595,N_5668);
nor U6388 (N_6388,N_5376,N_5697);
nor U6389 (N_6389,N_5484,N_5469);
or U6390 (N_6390,N_5565,N_5392);
or U6391 (N_6391,N_5372,N_5786);
and U6392 (N_6392,N_5078,N_5734);
or U6393 (N_6393,N_5399,N_5445);
and U6394 (N_6394,N_5961,N_5803);
and U6395 (N_6395,N_5510,N_5717);
or U6396 (N_6396,N_5998,N_5500);
nor U6397 (N_6397,N_5568,N_5635);
nor U6398 (N_6398,N_5839,N_5308);
nor U6399 (N_6399,N_5472,N_5967);
or U6400 (N_6400,N_5688,N_5357);
nor U6401 (N_6401,N_5288,N_5312);
nor U6402 (N_6402,N_5278,N_5031);
and U6403 (N_6403,N_5240,N_5731);
nor U6404 (N_6404,N_5898,N_5942);
nor U6405 (N_6405,N_5418,N_5790);
and U6406 (N_6406,N_5094,N_5143);
nand U6407 (N_6407,N_5653,N_5611);
or U6408 (N_6408,N_5857,N_5429);
nand U6409 (N_6409,N_5645,N_5402);
and U6410 (N_6410,N_5433,N_5092);
nand U6411 (N_6411,N_5168,N_5739);
nand U6412 (N_6412,N_5582,N_5986);
nand U6413 (N_6413,N_5727,N_5017);
nand U6414 (N_6414,N_5791,N_5202);
or U6415 (N_6415,N_5921,N_5902);
or U6416 (N_6416,N_5428,N_5591);
nand U6417 (N_6417,N_5043,N_5901);
nand U6418 (N_6418,N_5306,N_5474);
nand U6419 (N_6419,N_5189,N_5947);
nand U6420 (N_6420,N_5243,N_5599);
or U6421 (N_6421,N_5979,N_5489);
nand U6422 (N_6422,N_5520,N_5245);
or U6423 (N_6423,N_5083,N_5102);
or U6424 (N_6424,N_5983,N_5630);
nand U6425 (N_6425,N_5015,N_5048);
or U6426 (N_6426,N_5826,N_5887);
nor U6427 (N_6427,N_5013,N_5923);
nor U6428 (N_6428,N_5813,N_5584);
or U6429 (N_6429,N_5059,N_5391);
nand U6430 (N_6430,N_5108,N_5298);
or U6431 (N_6431,N_5232,N_5807);
nor U6432 (N_6432,N_5107,N_5770);
and U6433 (N_6433,N_5228,N_5723);
nor U6434 (N_6434,N_5193,N_5763);
nand U6435 (N_6435,N_5793,N_5293);
nand U6436 (N_6436,N_5736,N_5342);
or U6437 (N_6437,N_5112,N_5659);
and U6438 (N_6438,N_5818,N_5643);
or U6439 (N_6439,N_5061,N_5867);
nand U6440 (N_6440,N_5957,N_5904);
nor U6441 (N_6441,N_5926,N_5183);
and U6442 (N_6442,N_5341,N_5652);
nor U6443 (N_6443,N_5456,N_5451);
nor U6444 (N_6444,N_5647,N_5885);
nor U6445 (N_6445,N_5602,N_5134);
nand U6446 (N_6446,N_5104,N_5099);
nand U6447 (N_6447,N_5876,N_5910);
and U6448 (N_6448,N_5436,N_5217);
nor U6449 (N_6449,N_5413,N_5324);
nor U6450 (N_6450,N_5758,N_5870);
or U6451 (N_6451,N_5753,N_5673);
nand U6452 (N_6452,N_5508,N_5219);
nand U6453 (N_6453,N_5091,N_5502);
or U6454 (N_6454,N_5579,N_5487);
nor U6455 (N_6455,N_5058,N_5760);
nand U6456 (N_6456,N_5756,N_5946);
and U6457 (N_6457,N_5396,N_5848);
and U6458 (N_6458,N_5273,N_5258);
nor U6459 (N_6459,N_5615,N_5825);
and U6460 (N_6460,N_5201,N_5654);
nand U6461 (N_6461,N_5096,N_5554);
nand U6462 (N_6462,N_5744,N_5106);
or U6463 (N_6463,N_5732,N_5767);
or U6464 (N_6464,N_5838,N_5270);
or U6465 (N_6465,N_5604,N_5594);
or U6466 (N_6466,N_5037,N_5325);
and U6467 (N_6467,N_5441,N_5951);
nand U6468 (N_6468,N_5006,N_5562);
nor U6469 (N_6469,N_5319,N_5025);
nand U6470 (N_6470,N_5473,N_5249);
or U6471 (N_6471,N_5360,N_5821);
or U6472 (N_6472,N_5010,N_5384);
or U6473 (N_6473,N_5263,N_5527);
nor U6474 (N_6474,N_5140,N_5121);
or U6475 (N_6475,N_5458,N_5137);
nand U6476 (N_6476,N_5420,N_5945);
nor U6477 (N_6477,N_5806,N_5229);
nand U6478 (N_6478,N_5299,N_5264);
nor U6479 (N_6479,N_5799,N_5162);
and U6480 (N_6480,N_5206,N_5279);
nor U6481 (N_6481,N_5275,N_5960);
nor U6482 (N_6482,N_5964,N_5259);
nor U6483 (N_6483,N_5142,N_5070);
and U6484 (N_6484,N_5497,N_5925);
or U6485 (N_6485,N_5047,N_5395);
and U6486 (N_6486,N_5729,N_5915);
nor U6487 (N_6487,N_5841,N_5340);
nor U6488 (N_6488,N_5802,N_5056);
nand U6489 (N_6489,N_5282,N_5375);
nor U6490 (N_6490,N_5975,N_5397);
and U6491 (N_6491,N_5203,N_5339);
or U6492 (N_6492,N_5662,N_5310);
nor U6493 (N_6493,N_5532,N_5055);
or U6494 (N_6494,N_5097,N_5417);
nand U6495 (N_6495,N_5215,N_5024);
nand U6496 (N_6496,N_5866,N_5007);
or U6497 (N_6497,N_5650,N_5590);
nand U6498 (N_6498,N_5948,N_5619);
nor U6499 (N_6499,N_5624,N_5646);
nand U6500 (N_6500,N_5244,N_5874);
and U6501 (N_6501,N_5349,N_5599);
and U6502 (N_6502,N_5604,N_5657);
nand U6503 (N_6503,N_5805,N_5457);
nor U6504 (N_6504,N_5046,N_5352);
or U6505 (N_6505,N_5192,N_5633);
nand U6506 (N_6506,N_5831,N_5599);
nor U6507 (N_6507,N_5592,N_5967);
and U6508 (N_6508,N_5294,N_5679);
nand U6509 (N_6509,N_5379,N_5925);
or U6510 (N_6510,N_5194,N_5090);
or U6511 (N_6511,N_5382,N_5942);
or U6512 (N_6512,N_5780,N_5525);
and U6513 (N_6513,N_5880,N_5533);
nand U6514 (N_6514,N_5717,N_5520);
nand U6515 (N_6515,N_5309,N_5028);
or U6516 (N_6516,N_5248,N_5825);
nand U6517 (N_6517,N_5526,N_5734);
nand U6518 (N_6518,N_5836,N_5053);
nand U6519 (N_6519,N_5687,N_5343);
nor U6520 (N_6520,N_5814,N_5910);
and U6521 (N_6521,N_5925,N_5134);
and U6522 (N_6522,N_5679,N_5495);
xnor U6523 (N_6523,N_5987,N_5359);
nor U6524 (N_6524,N_5644,N_5812);
or U6525 (N_6525,N_5767,N_5261);
and U6526 (N_6526,N_5856,N_5937);
and U6527 (N_6527,N_5049,N_5674);
or U6528 (N_6528,N_5324,N_5098);
nor U6529 (N_6529,N_5976,N_5326);
and U6530 (N_6530,N_5533,N_5191);
nor U6531 (N_6531,N_5615,N_5226);
nor U6532 (N_6532,N_5275,N_5513);
nand U6533 (N_6533,N_5715,N_5639);
and U6534 (N_6534,N_5076,N_5717);
or U6535 (N_6535,N_5133,N_5670);
nor U6536 (N_6536,N_5147,N_5173);
and U6537 (N_6537,N_5908,N_5609);
and U6538 (N_6538,N_5155,N_5271);
nor U6539 (N_6539,N_5814,N_5499);
and U6540 (N_6540,N_5755,N_5125);
nand U6541 (N_6541,N_5223,N_5145);
or U6542 (N_6542,N_5502,N_5421);
or U6543 (N_6543,N_5212,N_5856);
or U6544 (N_6544,N_5174,N_5523);
and U6545 (N_6545,N_5947,N_5775);
or U6546 (N_6546,N_5887,N_5601);
and U6547 (N_6547,N_5919,N_5893);
nand U6548 (N_6548,N_5428,N_5932);
and U6549 (N_6549,N_5981,N_5215);
nor U6550 (N_6550,N_5348,N_5717);
and U6551 (N_6551,N_5306,N_5573);
and U6552 (N_6552,N_5949,N_5240);
nor U6553 (N_6553,N_5110,N_5165);
nor U6554 (N_6554,N_5318,N_5473);
or U6555 (N_6555,N_5684,N_5800);
and U6556 (N_6556,N_5578,N_5951);
nand U6557 (N_6557,N_5815,N_5927);
nor U6558 (N_6558,N_5484,N_5594);
and U6559 (N_6559,N_5340,N_5031);
or U6560 (N_6560,N_5224,N_5498);
nor U6561 (N_6561,N_5292,N_5421);
and U6562 (N_6562,N_5680,N_5794);
or U6563 (N_6563,N_5775,N_5657);
nand U6564 (N_6564,N_5191,N_5108);
or U6565 (N_6565,N_5437,N_5276);
or U6566 (N_6566,N_5594,N_5467);
nor U6567 (N_6567,N_5562,N_5930);
or U6568 (N_6568,N_5728,N_5875);
nand U6569 (N_6569,N_5809,N_5386);
or U6570 (N_6570,N_5043,N_5923);
or U6571 (N_6571,N_5113,N_5093);
or U6572 (N_6572,N_5671,N_5987);
nand U6573 (N_6573,N_5755,N_5220);
nor U6574 (N_6574,N_5337,N_5867);
and U6575 (N_6575,N_5588,N_5970);
or U6576 (N_6576,N_5038,N_5719);
nand U6577 (N_6577,N_5687,N_5785);
nand U6578 (N_6578,N_5737,N_5440);
nand U6579 (N_6579,N_5883,N_5819);
xor U6580 (N_6580,N_5899,N_5595);
nor U6581 (N_6581,N_5622,N_5055);
or U6582 (N_6582,N_5078,N_5593);
or U6583 (N_6583,N_5122,N_5371);
nand U6584 (N_6584,N_5214,N_5125);
or U6585 (N_6585,N_5398,N_5634);
or U6586 (N_6586,N_5882,N_5453);
or U6587 (N_6587,N_5201,N_5058);
or U6588 (N_6588,N_5493,N_5605);
nor U6589 (N_6589,N_5797,N_5388);
or U6590 (N_6590,N_5236,N_5050);
and U6591 (N_6591,N_5671,N_5006);
and U6592 (N_6592,N_5315,N_5161);
and U6593 (N_6593,N_5343,N_5318);
xor U6594 (N_6594,N_5337,N_5531);
or U6595 (N_6595,N_5456,N_5661);
or U6596 (N_6596,N_5089,N_5472);
and U6597 (N_6597,N_5705,N_5899);
or U6598 (N_6598,N_5647,N_5465);
nand U6599 (N_6599,N_5983,N_5282);
and U6600 (N_6600,N_5575,N_5959);
and U6601 (N_6601,N_5368,N_5346);
nand U6602 (N_6602,N_5350,N_5567);
or U6603 (N_6603,N_5407,N_5711);
nor U6604 (N_6604,N_5453,N_5653);
and U6605 (N_6605,N_5971,N_5288);
nor U6606 (N_6606,N_5158,N_5012);
and U6607 (N_6607,N_5464,N_5263);
nor U6608 (N_6608,N_5453,N_5954);
nand U6609 (N_6609,N_5902,N_5165);
nand U6610 (N_6610,N_5740,N_5041);
nor U6611 (N_6611,N_5413,N_5625);
and U6612 (N_6612,N_5815,N_5052);
nor U6613 (N_6613,N_5886,N_5070);
nor U6614 (N_6614,N_5993,N_5212);
and U6615 (N_6615,N_5519,N_5825);
nor U6616 (N_6616,N_5036,N_5007);
nand U6617 (N_6617,N_5467,N_5051);
and U6618 (N_6618,N_5075,N_5008);
nor U6619 (N_6619,N_5640,N_5859);
or U6620 (N_6620,N_5828,N_5092);
nor U6621 (N_6621,N_5988,N_5622);
nand U6622 (N_6622,N_5523,N_5838);
and U6623 (N_6623,N_5566,N_5293);
nand U6624 (N_6624,N_5234,N_5005);
and U6625 (N_6625,N_5984,N_5690);
or U6626 (N_6626,N_5772,N_5109);
and U6627 (N_6627,N_5459,N_5620);
and U6628 (N_6628,N_5647,N_5127);
nor U6629 (N_6629,N_5664,N_5747);
and U6630 (N_6630,N_5033,N_5793);
and U6631 (N_6631,N_5539,N_5142);
nor U6632 (N_6632,N_5730,N_5631);
nand U6633 (N_6633,N_5166,N_5798);
and U6634 (N_6634,N_5825,N_5973);
or U6635 (N_6635,N_5890,N_5191);
nor U6636 (N_6636,N_5144,N_5467);
nor U6637 (N_6637,N_5377,N_5406);
or U6638 (N_6638,N_5939,N_5195);
nor U6639 (N_6639,N_5473,N_5356);
or U6640 (N_6640,N_5229,N_5765);
or U6641 (N_6641,N_5814,N_5055);
nand U6642 (N_6642,N_5298,N_5416);
and U6643 (N_6643,N_5666,N_5886);
or U6644 (N_6644,N_5318,N_5260);
nand U6645 (N_6645,N_5690,N_5492);
or U6646 (N_6646,N_5624,N_5181);
and U6647 (N_6647,N_5085,N_5846);
and U6648 (N_6648,N_5991,N_5260);
nand U6649 (N_6649,N_5933,N_5638);
or U6650 (N_6650,N_5031,N_5249);
nand U6651 (N_6651,N_5518,N_5767);
nand U6652 (N_6652,N_5957,N_5837);
nand U6653 (N_6653,N_5339,N_5124);
or U6654 (N_6654,N_5434,N_5765);
or U6655 (N_6655,N_5181,N_5679);
nor U6656 (N_6656,N_5203,N_5439);
or U6657 (N_6657,N_5121,N_5246);
or U6658 (N_6658,N_5108,N_5885);
nor U6659 (N_6659,N_5415,N_5786);
and U6660 (N_6660,N_5689,N_5679);
and U6661 (N_6661,N_5248,N_5941);
and U6662 (N_6662,N_5943,N_5970);
nor U6663 (N_6663,N_5427,N_5213);
and U6664 (N_6664,N_5530,N_5209);
nand U6665 (N_6665,N_5545,N_5259);
nor U6666 (N_6666,N_5909,N_5366);
or U6667 (N_6667,N_5016,N_5391);
or U6668 (N_6668,N_5762,N_5940);
nor U6669 (N_6669,N_5359,N_5639);
nor U6670 (N_6670,N_5309,N_5724);
nand U6671 (N_6671,N_5103,N_5140);
nand U6672 (N_6672,N_5909,N_5715);
and U6673 (N_6673,N_5121,N_5086);
and U6674 (N_6674,N_5985,N_5235);
nor U6675 (N_6675,N_5232,N_5755);
and U6676 (N_6676,N_5600,N_5274);
or U6677 (N_6677,N_5812,N_5264);
and U6678 (N_6678,N_5777,N_5952);
nand U6679 (N_6679,N_5644,N_5228);
nor U6680 (N_6680,N_5402,N_5918);
and U6681 (N_6681,N_5306,N_5005);
or U6682 (N_6682,N_5913,N_5661);
nand U6683 (N_6683,N_5426,N_5668);
nor U6684 (N_6684,N_5121,N_5633);
nor U6685 (N_6685,N_5956,N_5396);
nand U6686 (N_6686,N_5049,N_5636);
or U6687 (N_6687,N_5496,N_5500);
or U6688 (N_6688,N_5153,N_5805);
nand U6689 (N_6689,N_5573,N_5121);
and U6690 (N_6690,N_5794,N_5017);
nor U6691 (N_6691,N_5101,N_5689);
or U6692 (N_6692,N_5466,N_5929);
and U6693 (N_6693,N_5655,N_5448);
nor U6694 (N_6694,N_5555,N_5332);
or U6695 (N_6695,N_5843,N_5572);
and U6696 (N_6696,N_5767,N_5158);
nand U6697 (N_6697,N_5991,N_5885);
and U6698 (N_6698,N_5067,N_5774);
nor U6699 (N_6699,N_5192,N_5271);
nand U6700 (N_6700,N_5367,N_5033);
nor U6701 (N_6701,N_5678,N_5976);
and U6702 (N_6702,N_5448,N_5788);
nand U6703 (N_6703,N_5749,N_5233);
nor U6704 (N_6704,N_5897,N_5170);
and U6705 (N_6705,N_5679,N_5135);
nand U6706 (N_6706,N_5468,N_5484);
nor U6707 (N_6707,N_5990,N_5253);
or U6708 (N_6708,N_5496,N_5412);
or U6709 (N_6709,N_5075,N_5598);
and U6710 (N_6710,N_5392,N_5740);
nor U6711 (N_6711,N_5945,N_5418);
nand U6712 (N_6712,N_5688,N_5757);
and U6713 (N_6713,N_5236,N_5168);
or U6714 (N_6714,N_5607,N_5641);
and U6715 (N_6715,N_5048,N_5340);
nor U6716 (N_6716,N_5376,N_5978);
nor U6717 (N_6717,N_5327,N_5627);
and U6718 (N_6718,N_5442,N_5118);
or U6719 (N_6719,N_5567,N_5066);
and U6720 (N_6720,N_5549,N_5383);
or U6721 (N_6721,N_5365,N_5823);
nand U6722 (N_6722,N_5358,N_5865);
and U6723 (N_6723,N_5465,N_5928);
nand U6724 (N_6724,N_5228,N_5298);
or U6725 (N_6725,N_5061,N_5637);
and U6726 (N_6726,N_5149,N_5694);
nand U6727 (N_6727,N_5008,N_5846);
and U6728 (N_6728,N_5902,N_5766);
and U6729 (N_6729,N_5406,N_5961);
and U6730 (N_6730,N_5537,N_5093);
nand U6731 (N_6731,N_5638,N_5313);
or U6732 (N_6732,N_5758,N_5863);
and U6733 (N_6733,N_5075,N_5738);
nor U6734 (N_6734,N_5506,N_5059);
nor U6735 (N_6735,N_5965,N_5194);
nand U6736 (N_6736,N_5184,N_5536);
xnor U6737 (N_6737,N_5467,N_5654);
or U6738 (N_6738,N_5388,N_5537);
nand U6739 (N_6739,N_5114,N_5347);
or U6740 (N_6740,N_5887,N_5299);
nor U6741 (N_6741,N_5216,N_5242);
nand U6742 (N_6742,N_5636,N_5098);
nor U6743 (N_6743,N_5656,N_5499);
nor U6744 (N_6744,N_5532,N_5371);
nor U6745 (N_6745,N_5959,N_5814);
nand U6746 (N_6746,N_5983,N_5504);
and U6747 (N_6747,N_5335,N_5143);
nand U6748 (N_6748,N_5851,N_5792);
xor U6749 (N_6749,N_5757,N_5165);
nor U6750 (N_6750,N_5332,N_5483);
nand U6751 (N_6751,N_5875,N_5760);
nor U6752 (N_6752,N_5911,N_5377);
and U6753 (N_6753,N_5804,N_5976);
and U6754 (N_6754,N_5565,N_5199);
nor U6755 (N_6755,N_5411,N_5495);
nand U6756 (N_6756,N_5353,N_5997);
or U6757 (N_6757,N_5322,N_5488);
or U6758 (N_6758,N_5306,N_5873);
nand U6759 (N_6759,N_5432,N_5414);
and U6760 (N_6760,N_5555,N_5220);
and U6761 (N_6761,N_5249,N_5094);
nor U6762 (N_6762,N_5004,N_5316);
nor U6763 (N_6763,N_5268,N_5211);
nand U6764 (N_6764,N_5095,N_5835);
and U6765 (N_6765,N_5896,N_5557);
nand U6766 (N_6766,N_5870,N_5283);
nand U6767 (N_6767,N_5937,N_5303);
and U6768 (N_6768,N_5925,N_5217);
or U6769 (N_6769,N_5611,N_5533);
and U6770 (N_6770,N_5050,N_5404);
or U6771 (N_6771,N_5370,N_5869);
nand U6772 (N_6772,N_5163,N_5333);
and U6773 (N_6773,N_5324,N_5998);
or U6774 (N_6774,N_5963,N_5422);
or U6775 (N_6775,N_5824,N_5112);
or U6776 (N_6776,N_5514,N_5562);
nand U6777 (N_6777,N_5815,N_5626);
or U6778 (N_6778,N_5126,N_5789);
or U6779 (N_6779,N_5223,N_5902);
xnor U6780 (N_6780,N_5225,N_5308);
nand U6781 (N_6781,N_5064,N_5877);
nor U6782 (N_6782,N_5036,N_5146);
nor U6783 (N_6783,N_5372,N_5231);
and U6784 (N_6784,N_5240,N_5195);
nand U6785 (N_6785,N_5350,N_5839);
nand U6786 (N_6786,N_5577,N_5648);
nor U6787 (N_6787,N_5427,N_5433);
nand U6788 (N_6788,N_5049,N_5718);
or U6789 (N_6789,N_5946,N_5067);
and U6790 (N_6790,N_5022,N_5070);
nand U6791 (N_6791,N_5772,N_5993);
and U6792 (N_6792,N_5711,N_5258);
nor U6793 (N_6793,N_5678,N_5159);
nand U6794 (N_6794,N_5064,N_5571);
and U6795 (N_6795,N_5325,N_5393);
and U6796 (N_6796,N_5376,N_5969);
nand U6797 (N_6797,N_5454,N_5763);
and U6798 (N_6798,N_5735,N_5445);
nand U6799 (N_6799,N_5070,N_5516);
and U6800 (N_6800,N_5670,N_5935);
nand U6801 (N_6801,N_5249,N_5779);
or U6802 (N_6802,N_5981,N_5356);
nand U6803 (N_6803,N_5987,N_5402);
nor U6804 (N_6804,N_5879,N_5826);
and U6805 (N_6805,N_5952,N_5453);
nand U6806 (N_6806,N_5526,N_5098);
nor U6807 (N_6807,N_5834,N_5153);
nand U6808 (N_6808,N_5944,N_5971);
and U6809 (N_6809,N_5175,N_5207);
nor U6810 (N_6810,N_5625,N_5763);
and U6811 (N_6811,N_5202,N_5093);
or U6812 (N_6812,N_5831,N_5354);
and U6813 (N_6813,N_5109,N_5376);
and U6814 (N_6814,N_5879,N_5600);
nand U6815 (N_6815,N_5969,N_5623);
nand U6816 (N_6816,N_5877,N_5767);
xnor U6817 (N_6817,N_5408,N_5040);
nor U6818 (N_6818,N_5538,N_5486);
and U6819 (N_6819,N_5636,N_5746);
or U6820 (N_6820,N_5350,N_5273);
nand U6821 (N_6821,N_5006,N_5725);
nand U6822 (N_6822,N_5599,N_5310);
or U6823 (N_6823,N_5118,N_5572);
and U6824 (N_6824,N_5701,N_5973);
or U6825 (N_6825,N_5527,N_5001);
nand U6826 (N_6826,N_5357,N_5601);
nand U6827 (N_6827,N_5604,N_5774);
or U6828 (N_6828,N_5747,N_5002);
nor U6829 (N_6829,N_5202,N_5520);
nor U6830 (N_6830,N_5707,N_5090);
nand U6831 (N_6831,N_5853,N_5318);
nor U6832 (N_6832,N_5097,N_5093);
or U6833 (N_6833,N_5441,N_5649);
or U6834 (N_6834,N_5037,N_5218);
and U6835 (N_6835,N_5880,N_5014);
nor U6836 (N_6836,N_5851,N_5176);
nand U6837 (N_6837,N_5959,N_5431);
or U6838 (N_6838,N_5572,N_5635);
nand U6839 (N_6839,N_5482,N_5185);
and U6840 (N_6840,N_5881,N_5800);
or U6841 (N_6841,N_5109,N_5995);
or U6842 (N_6842,N_5941,N_5327);
or U6843 (N_6843,N_5594,N_5853);
nand U6844 (N_6844,N_5548,N_5510);
nand U6845 (N_6845,N_5898,N_5193);
nand U6846 (N_6846,N_5624,N_5004);
and U6847 (N_6847,N_5367,N_5309);
nand U6848 (N_6848,N_5418,N_5732);
nor U6849 (N_6849,N_5023,N_5114);
nor U6850 (N_6850,N_5968,N_5365);
nor U6851 (N_6851,N_5801,N_5278);
nand U6852 (N_6852,N_5472,N_5012);
nand U6853 (N_6853,N_5151,N_5818);
and U6854 (N_6854,N_5924,N_5320);
nor U6855 (N_6855,N_5032,N_5045);
nor U6856 (N_6856,N_5117,N_5250);
nand U6857 (N_6857,N_5427,N_5040);
or U6858 (N_6858,N_5595,N_5066);
and U6859 (N_6859,N_5383,N_5704);
nand U6860 (N_6860,N_5393,N_5123);
or U6861 (N_6861,N_5207,N_5398);
or U6862 (N_6862,N_5987,N_5639);
nand U6863 (N_6863,N_5962,N_5691);
or U6864 (N_6864,N_5304,N_5358);
nand U6865 (N_6865,N_5221,N_5076);
or U6866 (N_6866,N_5590,N_5749);
nand U6867 (N_6867,N_5172,N_5512);
xor U6868 (N_6868,N_5329,N_5862);
and U6869 (N_6869,N_5471,N_5822);
nand U6870 (N_6870,N_5457,N_5803);
nand U6871 (N_6871,N_5022,N_5515);
nor U6872 (N_6872,N_5152,N_5242);
and U6873 (N_6873,N_5556,N_5899);
or U6874 (N_6874,N_5697,N_5186);
nand U6875 (N_6875,N_5917,N_5620);
and U6876 (N_6876,N_5754,N_5226);
nor U6877 (N_6877,N_5069,N_5724);
nor U6878 (N_6878,N_5280,N_5259);
or U6879 (N_6879,N_5520,N_5434);
and U6880 (N_6880,N_5354,N_5490);
or U6881 (N_6881,N_5034,N_5629);
and U6882 (N_6882,N_5873,N_5488);
nand U6883 (N_6883,N_5117,N_5640);
nor U6884 (N_6884,N_5222,N_5815);
nand U6885 (N_6885,N_5484,N_5136);
and U6886 (N_6886,N_5920,N_5510);
nor U6887 (N_6887,N_5631,N_5662);
nor U6888 (N_6888,N_5580,N_5485);
and U6889 (N_6889,N_5288,N_5916);
nor U6890 (N_6890,N_5742,N_5920);
nor U6891 (N_6891,N_5510,N_5307);
nand U6892 (N_6892,N_5878,N_5963);
nor U6893 (N_6893,N_5293,N_5811);
and U6894 (N_6894,N_5060,N_5008);
nor U6895 (N_6895,N_5518,N_5198);
nor U6896 (N_6896,N_5395,N_5018);
nor U6897 (N_6897,N_5919,N_5384);
and U6898 (N_6898,N_5787,N_5677);
nand U6899 (N_6899,N_5713,N_5042);
nor U6900 (N_6900,N_5803,N_5544);
nand U6901 (N_6901,N_5396,N_5728);
nand U6902 (N_6902,N_5068,N_5429);
or U6903 (N_6903,N_5558,N_5766);
nor U6904 (N_6904,N_5930,N_5635);
nand U6905 (N_6905,N_5735,N_5865);
nor U6906 (N_6906,N_5195,N_5433);
or U6907 (N_6907,N_5685,N_5486);
and U6908 (N_6908,N_5232,N_5470);
nor U6909 (N_6909,N_5861,N_5660);
nand U6910 (N_6910,N_5816,N_5460);
nor U6911 (N_6911,N_5175,N_5574);
and U6912 (N_6912,N_5897,N_5939);
nor U6913 (N_6913,N_5048,N_5053);
nor U6914 (N_6914,N_5253,N_5208);
and U6915 (N_6915,N_5103,N_5222);
and U6916 (N_6916,N_5715,N_5954);
nand U6917 (N_6917,N_5025,N_5437);
and U6918 (N_6918,N_5301,N_5238);
or U6919 (N_6919,N_5553,N_5116);
or U6920 (N_6920,N_5501,N_5968);
nor U6921 (N_6921,N_5073,N_5863);
nand U6922 (N_6922,N_5224,N_5250);
nand U6923 (N_6923,N_5377,N_5958);
and U6924 (N_6924,N_5023,N_5542);
nand U6925 (N_6925,N_5566,N_5973);
or U6926 (N_6926,N_5088,N_5306);
or U6927 (N_6927,N_5762,N_5075);
nand U6928 (N_6928,N_5446,N_5555);
nand U6929 (N_6929,N_5252,N_5581);
or U6930 (N_6930,N_5210,N_5881);
or U6931 (N_6931,N_5669,N_5161);
or U6932 (N_6932,N_5631,N_5479);
nor U6933 (N_6933,N_5237,N_5452);
nor U6934 (N_6934,N_5858,N_5737);
and U6935 (N_6935,N_5190,N_5281);
or U6936 (N_6936,N_5610,N_5981);
or U6937 (N_6937,N_5222,N_5581);
or U6938 (N_6938,N_5718,N_5938);
nand U6939 (N_6939,N_5110,N_5017);
nand U6940 (N_6940,N_5804,N_5230);
and U6941 (N_6941,N_5703,N_5280);
nand U6942 (N_6942,N_5289,N_5007);
nand U6943 (N_6943,N_5953,N_5838);
or U6944 (N_6944,N_5840,N_5170);
or U6945 (N_6945,N_5532,N_5451);
nor U6946 (N_6946,N_5055,N_5243);
nand U6947 (N_6947,N_5925,N_5625);
nor U6948 (N_6948,N_5378,N_5597);
and U6949 (N_6949,N_5949,N_5477);
nor U6950 (N_6950,N_5025,N_5850);
nor U6951 (N_6951,N_5766,N_5734);
nor U6952 (N_6952,N_5375,N_5362);
xor U6953 (N_6953,N_5832,N_5946);
nor U6954 (N_6954,N_5229,N_5284);
and U6955 (N_6955,N_5101,N_5368);
nand U6956 (N_6956,N_5701,N_5873);
nor U6957 (N_6957,N_5655,N_5773);
nor U6958 (N_6958,N_5568,N_5542);
and U6959 (N_6959,N_5775,N_5902);
and U6960 (N_6960,N_5696,N_5938);
nor U6961 (N_6961,N_5132,N_5242);
or U6962 (N_6962,N_5875,N_5822);
or U6963 (N_6963,N_5463,N_5123);
nand U6964 (N_6964,N_5350,N_5580);
nor U6965 (N_6965,N_5104,N_5692);
nand U6966 (N_6966,N_5110,N_5446);
nand U6967 (N_6967,N_5892,N_5691);
or U6968 (N_6968,N_5702,N_5453);
nor U6969 (N_6969,N_5291,N_5662);
or U6970 (N_6970,N_5974,N_5303);
and U6971 (N_6971,N_5821,N_5126);
nand U6972 (N_6972,N_5798,N_5199);
nor U6973 (N_6973,N_5244,N_5687);
nand U6974 (N_6974,N_5287,N_5363);
nor U6975 (N_6975,N_5840,N_5965);
and U6976 (N_6976,N_5552,N_5938);
and U6977 (N_6977,N_5369,N_5567);
and U6978 (N_6978,N_5707,N_5277);
nor U6979 (N_6979,N_5934,N_5336);
or U6980 (N_6980,N_5867,N_5959);
or U6981 (N_6981,N_5583,N_5786);
or U6982 (N_6982,N_5229,N_5238);
nor U6983 (N_6983,N_5062,N_5022);
and U6984 (N_6984,N_5253,N_5794);
and U6985 (N_6985,N_5218,N_5330);
or U6986 (N_6986,N_5910,N_5891);
or U6987 (N_6987,N_5697,N_5693);
nand U6988 (N_6988,N_5952,N_5307);
nand U6989 (N_6989,N_5784,N_5749);
or U6990 (N_6990,N_5616,N_5271);
nor U6991 (N_6991,N_5546,N_5807);
nand U6992 (N_6992,N_5359,N_5298);
nor U6993 (N_6993,N_5559,N_5818);
nand U6994 (N_6994,N_5328,N_5094);
nand U6995 (N_6995,N_5360,N_5785);
nand U6996 (N_6996,N_5617,N_5340);
or U6997 (N_6997,N_5933,N_5410);
nand U6998 (N_6998,N_5413,N_5111);
nor U6999 (N_6999,N_5692,N_5509);
and U7000 (N_7000,N_6368,N_6210);
and U7001 (N_7001,N_6899,N_6299);
nor U7002 (N_7002,N_6016,N_6557);
and U7003 (N_7003,N_6204,N_6052);
nand U7004 (N_7004,N_6571,N_6115);
nand U7005 (N_7005,N_6757,N_6582);
and U7006 (N_7006,N_6732,N_6618);
nor U7007 (N_7007,N_6507,N_6638);
and U7008 (N_7008,N_6498,N_6238);
or U7009 (N_7009,N_6673,N_6942);
nand U7010 (N_7010,N_6463,N_6734);
or U7011 (N_7011,N_6758,N_6107);
and U7012 (N_7012,N_6380,N_6400);
nor U7013 (N_7013,N_6137,N_6147);
nand U7014 (N_7014,N_6139,N_6303);
and U7015 (N_7015,N_6510,N_6004);
nor U7016 (N_7016,N_6670,N_6185);
and U7017 (N_7017,N_6288,N_6837);
nor U7018 (N_7018,N_6241,N_6202);
and U7019 (N_7019,N_6746,N_6259);
nor U7020 (N_7020,N_6026,N_6982);
and U7021 (N_7021,N_6116,N_6071);
or U7022 (N_7022,N_6782,N_6079);
and U7023 (N_7023,N_6347,N_6583);
and U7024 (N_7024,N_6540,N_6991);
or U7025 (N_7025,N_6114,N_6033);
nor U7026 (N_7026,N_6740,N_6058);
and U7027 (N_7027,N_6785,N_6705);
or U7028 (N_7028,N_6146,N_6756);
and U7029 (N_7029,N_6887,N_6577);
nand U7030 (N_7030,N_6654,N_6766);
and U7031 (N_7031,N_6012,N_6057);
and U7032 (N_7032,N_6459,N_6763);
nand U7033 (N_7033,N_6983,N_6993);
nor U7034 (N_7034,N_6775,N_6417);
or U7035 (N_7035,N_6936,N_6219);
nand U7036 (N_7036,N_6244,N_6932);
nand U7037 (N_7037,N_6410,N_6869);
or U7038 (N_7038,N_6614,N_6158);
and U7039 (N_7039,N_6729,N_6579);
nor U7040 (N_7040,N_6726,N_6119);
or U7041 (N_7041,N_6945,N_6234);
nand U7042 (N_7042,N_6500,N_6858);
nor U7043 (N_7043,N_6327,N_6904);
or U7044 (N_7044,N_6255,N_6990);
and U7045 (N_7045,N_6431,N_6143);
nand U7046 (N_7046,N_6915,N_6964);
nor U7047 (N_7047,N_6326,N_6632);
or U7048 (N_7048,N_6674,N_6329);
nor U7049 (N_7049,N_6002,N_6061);
or U7050 (N_7050,N_6753,N_6651);
or U7051 (N_7051,N_6446,N_6434);
or U7052 (N_7052,N_6132,N_6968);
and U7053 (N_7053,N_6230,N_6166);
nor U7054 (N_7054,N_6124,N_6967);
nand U7055 (N_7055,N_6669,N_6903);
and U7056 (N_7056,N_6502,N_6205);
or U7057 (N_7057,N_6625,N_6831);
or U7058 (N_7058,N_6642,N_6416);
or U7059 (N_7059,N_6499,N_6679);
nor U7060 (N_7060,N_6795,N_6351);
or U7061 (N_7061,N_6037,N_6925);
or U7062 (N_7062,N_6515,N_6661);
or U7063 (N_7063,N_6769,N_6695);
nand U7064 (N_7064,N_6650,N_6429);
nor U7065 (N_7065,N_6573,N_6055);
nor U7066 (N_7066,N_6145,N_6163);
nor U7067 (N_7067,N_6880,N_6509);
or U7068 (N_7068,N_6840,N_6193);
nand U7069 (N_7069,N_6867,N_6525);
nand U7070 (N_7070,N_6387,N_6598);
and U7071 (N_7071,N_6554,N_6284);
or U7072 (N_7072,N_6118,N_6229);
and U7073 (N_7073,N_6767,N_6045);
or U7074 (N_7074,N_6042,N_6112);
nand U7075 (N_7075,N_6710,N_6896);
or U7076 (N_7076,N_6454,N_6104);
nor U7077 (N_7077,N_6103,N_6847);
nand U7078 (N_7078,N_6195,N_6129);
nand U7079 (N_7079,N_6302,N_6276);
and U7080 (N_7080,N_6580,N_6863);
or U7081 (N_7081,N_6138,N_6452);
nor U7082 (N_7082,N_6881,N_6736);
and U7083 (N_7083,N_6414,N_6585);
and U7084 (N_7084,N_6728,N_6181);
nand U7085 (N_7085,N_6700,N_6965);
xor U7086 (N_7086,N_6517,N_6804);
nor U7087 (N_7087,N_6701,N_6271);
and U7088 (N_7088,N_6290,N_6605);
or U7089 (N_7089,N_6047,N_6802);
and U7090 (N_7090,N_6151,N_6253);
nand U7091 (N_7091,N_6972,N_6934);
or U7092 (N_7092,N_6349,N_6369);
or U7093 (N_7093,N_6636,N_6018);
or U7094 (N_7094,N_6824,N_6487);
or U7095 (N_7095,N_6225,N_6168);
nor U7096 (N_7096,N_6312,N_6176);
or U7097 (N_7097,N_6875,N_6059);
or U7098 (N_7098,N_6631,N_6162);
nand U7099 (N_7099,N_6864,N_6978);
and U7100 (N_7100,N_6707,N_6960);
nand U7101 (N_7101,N_6572,N_6218);
nand U7102 (N_7102,N_6656,N_6992);
nand U7103 (N_7103,N_6551,N_6826);
nor U7104 (N_7104,N_6095,N_6280);
or U7105 (N_7105,N_6346,N_6818);
and U7106 (N_7106,N_6727,N_6739);
nor U7107 (N_7107,N_6134,N_6536);
nor U7108 (N_7108,N_6086,N_6981);
and U7109 (N_7109,N_6783,N_6492);
and U7110 (N_7110,N_6626,N_6196);
nor U7111 (N_7111,N_6444,N_6366);
nor U7112 (N_7112,N_6422,N_6220);
or U7113 (N_7113,N_6286,N_6954);
nor U7114 (N_7114,N_6297,N_6791);
or U7115 (N_7115,N_6628,N_6997);
or U7116 (N_7116,N_6512,N_6741);
or U7117 (N_7117,N_6479,N_6556);
or U7118 (N_7118,N_6278,N_6722);
nand U7119 (N_7119,N_6472,N_6592);
and U7120 (N_7120,N_6878,N_6174);
nand U7121 (N_7121,N_6566,N_6647);
or U7122 (N_7122,N_6017,N_6015);
nand U7123 (N_7123,N_6248,N_6040);
nor U7124 (N_7124,N_6078,N_6325);
nand U7125 (N_7125,N_6443,N_6064);
or U7126 (N_7126,N_6501,N_6352);
and U7127 (N_7127,N_6738,N_6730);
nand U7128 (N_7128,N_6148,N_6603);
nor U7129 (N_7129,N_6568,N_6039);
and U7130 (N_7130,N_6950,N_6610);
nand U7131 (N_7131,N_6305,N_6888);
nor U7132 (N_7132,N_6135,N_6923);
nand U7133 (N_7133,N_6706,N_6339);
nand U7134 (N_7134,N_6426,N_6399);
or U7135 (N_7135,N_6354,N_6270);
nor U7136 (N_7136,N_6165,N_6000);
and U7137 (N_7137,N_6609,N_6643);
nor U7138 (N_7138,N_6296,N_6341);
nor U7139 (N_7139,N_6180,N_6486);
nor U7140 (N_7140,N_6066,N_6121);
and U7141 (N_7141,N_6937,N_6406);
nor U7142 (N_7142,N_6687,N_6298);
nand U7143 (N_7143,N_6910,N_6876);
nor U7144 (N_7144,N_6591,N_6250);
and U7145 (N_7145,N_6697,N_6587);
and U7146 (N_7146,N_6357,N_6093);
nor U7147 (N_7147,N_6986,N_6488);
or U7148 (N_7148,N_6192,N_6083);
or U7149 (N_7149,N_6908,N_6633);
or U7150 (N_7150,N_6489,N_6513);
and U7151 (N_7151,N_6274,N_6649);
nand U7152 (N_7152,N_6608,N_6914);
nand U7153 (N_7153,N_6862,N_6313);
or U7154 (N_7154,N_6519,N_6279);
or U7155 (N_7155,N_6224,N_6081);
or U7156 (N_7156,N_6806,N_6413);
nand U7157 (N_7157,N_6569,N_6301);
nand U7158 (N_7158,N_6419,N_6835);
or U7159 (N_7159,N_6521,N_6594);
and U7160 (N_7160,N_6029,N_6949);
nor U7161 (N_7161,N_6987,N_6825);
or U7162 (N_7162,N_6542,N_6704);
nand U7163 (N_7163,N_6362,N_6761);
or U7164 (N_7164,N_6764,N_6593);
nor U7165 (N_7165,N_6090,N_6214);
nand U7166 (N_7166,N_6323,N_6317);
nand U7167 (N_7167,N_6639,N_6264);
nand U7168 (N_7168,N_6531,N_6751);
and U7169 (N_7169,N_6389,N_6013);
and U7170 (N_7170,N_6433,N_6772);
nor U7171 (N_7171,N_6401,N_6784);
nor U7172 (N_7172,N_6141,N_6179);
nand U7173 (N_7173,N_6088,N_6810);
and U7174 (N_7174,N_6544,N_6379);
or U7175 (N_7175,N_6754,N_6561);
nor U7176 (N_7176,N_6518,N_6645);
and U7177 (N_7177,N_6172,N_6690);
nand U7178 (N_7178,N_6073,N_6657);
nand U7179 (N_7179,N_6886,N_6282);
or U7180 (N_7180,N_6998,N_6342);
nand U7181 (N_7181,N_6617,N_6249);
nand U7182 (N_7182,N_6503,N_6939);
or U7183 (N_7183,N_6160,N_6957);
or U7184 (N_7184,N_6044,N_6331);
nand U7185 (N_7185,N_6091,N_6456);
and U7186 (N_7186,N_6333,N_6318);
nor U7187 (N_7187,N_6630,N_6283);
or U7188 (N_7188,N_6708,N_6381);
nor U7189 (N_7189,N_6439,N_6916);
or U7190 (N_7190,N_6269,N_6606);
nor U7191 (N_7191,N_6808,N_6130);
xor U7192 (N_7192,N_6336,N_6604);
and U7193 (N_7193,N_6909,N_6493);
and U7194 (N_7194,N_6021,N_6760);
and U7195 (N_7195,N_6799,N_6685);
and U7196 (N_7196,N_6830,N_6872);
nand U7197 (N_7197,N_6197,N_6584);
xnor U7198 (N_7198,N_6227,N_6098);
or U7199 (N_7199,N_6043,N_6467);
nor U7200 (N_7200,N_6156,N_6921);
nor U7201 (N_7201,N_6050,N_6745);
or U7202 (N_7202,N_6527,N_6948);
nor U7203 (N_7203,N_6848,N_6719);
nor U7204 (N_7204,N_6892,N_6611);
and U7205 (N_7205,N_6069,N_6874);
or U7206 (N_7206,N_6335,N_6524);
or U7207 (N_7207,N_6947,N_6721);
and U7208 (N_7208,N_6184,N_6574);
and U7209 (N_7209,N_6613,N_6311);
and U7210 (N_7210,N_6917,N_6984);
or U7211 (N_7211,N_6407,N_6348);
nor U7212 (N_7212,N_6843,N_6842);
xnor U7213 (N_7213,N_6355,N_6711);
nand U7214 (N_7214,N_6820,N_6516);
or U7215 (N_7215,N_6702,N_6671);
nand U7216 (N_7216,N_6668,N_6662);
nand U7217 (N_7217,N_6003,N_6023);
nand U7218 (N_7218,N_6200,N_6849);
nand U7219 (N_7219,N_6844,N_6226);
nor U7220 (N_7220,N_6251,N_6222);
nand U7221 (N_7221,N_6567,N_6750);
or U7222 (N_7222,N_6770,N_6683);
nor U7223 (N_7223,N_6712,N_6664);
or U7224 (N_7224,N_6126,N_6749);
nor U7225 (N_7225,N_6075,N_6599);
nor U7226 (N_7226,N_6217,N_6962);
or U7227 (N_7227,N_6694,N_6581);
nor U7228 (N_7228,N_6667,N_6242);
nor U7229 (N_7229,N_6666,N_6365);
nand U7230 (N_7230,N_6142,N_6080);
nand U7231 (N_7231,N_6438,N_6684);
nor U7232 (N_7232,N_6320,N_6113);
and U7233 (N_7233,N_6007,N_6575);
nor U7234 (N_7234,N_6788,N_6879);
and U7235 (N_7235,N_6010,N_6056);
and U7236 (N_7236,N_6032,N_6319);
nor U7237 (N_7237,N_6966,N_6063);
nand U7238 (N_7238,N_6999,N_6367);
nor U7239 (N_7239,N_6691,N_6263);
or U7240 (N_7240,N_6337,N_6272);
nor U7241 (N_7241,N_6236,N_6309);
nand U7242 (N_7242,N_6239,N_6257);
nand U7243 (N_7243,N_6123,N_6445);
nand U7244 (N_7244,N_6240,N_6857);
nand U7245 (N_7245,N_6310,N_6304);
nand U7246 (N_7246,N_6530,N_6852);
or U7247 (N_7247,N_6807,N_6550);
or U7248 (N_7248,N_6877,N_6839);
and U7249 (N_7249,N_6441,N_6001);
or U7250 (N_7250,N_6590,N_6070);
nor U7251 (N_7251,N_6332,N_6228);
nor U7252 (N_7252,N_6128,N_6461);
or U7253 (N_7253,N_6779,N_6829);
nand U7254 (N_7254,N_6562,N_6482);
or U7255 (N_7255,N_6053,N_6637);
and U7256 (N_7256,N_6906,N_6555);
nand U7257 (N_7257,N_6635,N_6612);
and U7258 (N_7258,N_6316,N_6405);
nand U7259 (N_7259,N_6797,N_6122);
nand U7260 (N_7260,N_6212,N_6131);
and U7261 (N_7261,N_6776,N_6928);
nor U7262 (N_7262,N_6895,N_6930);
nand U7263 (N_7263,N_6552,N_6321);
and U7264 (N_7264,N_6773,N_6087);
nand U7265 (N_7265,N_6440,N_6468);
and U7266 (N_7266,N_6287,N_6315);
or U7267 (N_7267,N_6005,N_6538);
or U7268 (N_7268,N_6809,N_6723);
nand U7269 (N_7269,N_6989,N_6774);
nor U7270 (N_7270,N_6344,N_6496);
and U7271 (N_7271,N_6988,N_6660);
nand U7272 (N_7272,N_6940,N_6485);
nand U7273 (N_7273,N_6101,N_6973);
nor U7274 (N_7274,N_6520,N_6768);
or U7275 (N_7275,N_6450,N_6935);
xnor U7276 (N_7276,N_6725,N_6164);
and U7277 (N_7277,N_6415,N_6159);
nand U7278 (N_7278,N_6827,N_6644);
nand U7279 (N_7279,N_6359,N_6698);
and U7280 (N_7280,N_6762,N_6565);
nand U7281 (N_7281,N_6623,N_6979);
and U7282 (N_7282,N_6109,N_6360);
nor U7283 (N_7283,N_6289,N_6437);
and U7284 (N_7284,N_6832,N_6363);
and U7285 (N_7285,N_6871,N_6523);
or U7286 (N_7286,N_6514,N_6815);
or U7287 (N_7287,N_6851,N_6996);
nand U7288 (N_7288,N_6085,N_6428);
and U7289 (N_7289,N_6024,N_6386);
nand U7290 (N_7290,N_6334,N_6621);
and U7291 (N_7291,N_6790,N_6006);
and U7292 (N_7292,N_6595,N_6777);
nand U7293 (N_7293,N_6374,N_6744);
nand U7294 (N_7294,N_6927,N_6752);
or U7295 (N_7295,N_6281,N_6385);
nor U7296 (N_7296,N_6794,N_6068);
and U7297 (N_7297,N_6466,N_6976);
and U7298 (N_7298,N_6716,N_6813);
or U7299 (N_7299,N_6850,N_6448);
nand U7300 (N_7300,N_6009,N_6682);
nand U7301 (N_7301,N_6285,N_6511);
or U7302 (N_7302,N_6860,N_6314);
and U7303 (N_7303,N_6823,N_6529);
and U7304 (N_7304,N_6120,N_6977);
nand U7305 (N_7305,N_6933,N_6108);
and U7306 (N_7306,N_6350,N_6060);
or U7307 (N_7307,N_6092,N_6534);
nor U7308 (N_7308,N_6918,N_6207);
nand U7309 (N_7309,N_6046,N_6570);
nand U7310 (N_7310,N_6586,N_6364);
nor U7311 (N_7311,N_6019,N_6789);
nor U7312 (N_7312,N_6640,N_6924);
and U7313 (N_7313,N_6911,N_6803);
xor U7314 (N_7314,N_6854,N_6372);
and U7315 (N_7315,N_6549,N_6041);
or U7316 (N_7316,N_6865,N_6898);
nand U7317 (N_7317,N_6475,N_6490);
and U7318 (N_7318,N_6796,N_6247);
nor U7319 (N_7319,N_6971,N_6233);
nand U7320 (N_7320,N_6755,N_6149);
and U7321 (N_7321,N_6476,N_6853);
and U7322 (N_7322,N_6470,N_6034);
nor U7323 (N_7323,N_6483,N_6970);
or U7324 (N_7324,N_6048,N_6338);
nand U7325 (N_7325,N_6397,N_6627);
or U7326 (N_7326,N_6235,N_6816);
nand U7327 (N_7327,N_6919,N_6084);
nand U7328 (N_7328,N_6717,N_6961);
or U7329 (N_7329,N_6600,N_6330);
nor U7330 (N_7330,N_6469,N_6607);
nor U7331 (N_7331,N_6678,N_6480);
nor U7332 (N_7332,N_6931,N_6328);
and U7333 (N_7333,N_6624,N_6901);
nor U7334 (N_7334,N_6491,N_6713);
nand U7335 (N_7335,N_6956,N_6402);
or U7336 (N_7336,N_6177,N_6038);
and U7337 (N_7337,N_6343,N_6051);
and U7338 (N_7338,N_6457,N_6273);
and U7339 (N_7339,N_6140,N_6735);
or U7340 (N_7340,N_6462,N_6306);
or U7341 (N_7341,N_6356,N_6508);
or U7342 (N_7342,N_6646,N_6194);
and U7343 (N_7343,N_6245,N_6846);
and U7344 (N_7344,N_6696,N_6008);
nor U7345 (N_7345,N_6481,N_6912);
and U7346 (N_7346,N_6543,N_6453);
or U7347 (N_7347,N_6619,N_6424);
nand U7348 (N_7348,N_6541,N_6375);
and U7349 (N_7349,N_6054,N_6792);
and U7350 (N_7350,N_6099,N_6747);
or U7351 (N_7351,N_6020,N_6748);
and U7352 (N_7352,N_6277,N_6153);
or U7353 (N_7353,N_6267,N_6724);
nand U7354 (N_7354,N_6294,N_6836);
nor U7355 (N_7355,N_6648,N_6464);
nor U7356 (N_7356,N_6199,N_6946);
or U7357 (N_7357,N_6035,N_6377);
nand U7358 (N_7358,N_6855,N_6620);
nor U7359 (N_7359,N_6111,N_6819);
xor U7360 (N_7360,N_6778,N_6822);
and U7361 (N_7361,N_6206,N_6564);
and U7362 (N_7362,N_6237,N_6256);
or U7363 (N_7363,N_6532,N_6834);
or U7364 (N_7364,N_6558,N_6067);
and U7365 (N_7365,N_6022,N_6963);
nor U7366 (N_7366,N_6065,N_6187);
and U7367 (N_7367,N_6188,N_6262);
xnor U7368 (N_7368,N_6526,N_6944);
and U7369 (N_7369,N_6025,N_6345);
nand U7370 (N_7370,N_6216,N_6152);
or U7371 (N_7371,N_6127,N_6588);
nor U7372 (N_7372,N_6036,N_6560);
or U7373 (N_7373,N_6689,N_6393);
nor U7374 (N_7374,N_6897,N_6412);
nor U7375 (N_7375,N_6293,N_6471);
or U7376 (N_7376,N_6985,N_6699);
nand U7377 (N_7377,N_6391,N_6442);
nand U7378 (N_7378,N_6223,N_6658);
nand U7379 (N_7379,N_6382,N_6014);
nand U7380 (N_7380,N_6292,N_6894);
nand U7381 (N_7381,N_6680,N_6266);
or U7382 (N_7382,N_6186,N_6845);
or U7383 (N_7383,N_6929,N_6432);
nand U7384 (N_7384,N_6893,N_6828);
nand U7385 (N_7385,N_6408,N_6157);
and U7386 (N_7386,N_6378,N_6535);
nor U7387 (N_7387,N_6506,N_6873);
and U7388 (N_7388,N_6952,N_6252);
nand U7389 (N_7389,N_6615,N_6975);
and U7390 (N_7390,N_6404,N_6089);
and U7391 (N_7391,N_6686,N_6907);
or U7392 (N_7392,N_6420,N_6136);
and U7393 (N_7393,N_6905,N_6943);
nand U7394 (N_7394,N_6601,N_6465);
xor U7395 (N_7395,N_6161,N_6801);
nor U7396 (N_7396,N_6074,N_6522);
or U7397 (N_7397,N_6629,N_6173);
or U7398 (N_7398,N_6505,N_6602);
nor U7399 (N_7399,N_6798,N_6616);
nor U7400 (N_7400,N_6793,N_6677);
nand U7401 (N_7401,N_6926,N_6028);
nand U7402 (N_7402,N_6353,N_6484);
and U7403 (N_7403,N_6548,N_6714);
or U7404 (N_7404,N_6681,N_6547);
and U7405 (N_7405,N_6733,N_6409);
nand U7406 (N_7406,N_6882,N_6436);
nand U7407 (N_7407,N_6418,N_6100);
nand U7408 (N_7408,N_6994,N_6451);
nand U7409 (N_7409,N_6995,N_6675);
or U7410 (N_7410,N_6150,N_6170);
nand U7411 (N_7411,N_6641,N_6383);
nand U7412 (N_7412,N_6105,N_6155);
xnor U7413 (N_7413,N_6403,N_6358);
and U7414 (N_7414,N_6838,N_6295);
and U7415 (N_7415,N_6821,N_6497);
nand U7416 (N_7416,N_6737,N_6211);
nand U7417 (N_7417,N_6361,N_6902);
nor U7418 (N_7418,N_6183,N_6027);
nor U7419 (N_7419,N_6388,N_6787);
nor U7420 (N_7420,N_6261,N_6900);
nand U7421 (N_7421,N_6913,N_6076);
nor U7422 (N_7422,N_6421,N_6395);
nand U7423 (N_7423,N_6477,N_6731);
and U7424 (N_7424,N_6889,N_6665);
nand U7425 (N_7425,N_6455,N_6265);
and U7426 (N_7426,N_6423,N_6692);
nand U7427 (N_7427,N_6715,N_6563);
nor U7428 (N_7428,N_6082,N_6528);
nor U7429 (N_7429,N_6841,N_6167);
and U7430 (N_7430,N_6144,N_6031);
or U7431 (N_7431,N_6676,N_6110);
nand U7432 (N_7432,N_6232,N_6545);
or U7433 (N_7433,N_6133,N_6655);
xor U7434 (N_7434,N_6049,N_6953);
nand U7435 (N_7435,N_6883,N_6300);
or U7436 (N_7436,N_6322,N_6425);
nand U7437 (N_7437,N_6030,N_6576);
or U7438 (N_7438,N_6652,N_6938);
and U7439 (N_7439,N_6473,N_6371);
nor U7440 (N_7440,N_6198,N_6494);
nand U7441 (N_7441,N_6659,N_6203);
nor U7442 (N_7442,N_6324,N_6861);
and U7443 (N_7443,N_6072,N_6922);
or U7444 (N_7444,N_6688,N_6718);
or U7445 (N_7445,N_6191,N_6275);
nor U7446 (N_7446,N_6663,N_6969);
or U7447 (N_7447,N_6759,N_6106);
and U7448 (N_7448,N_6182,N_6578);
nor U7449 (N_7449,N_6394,N_6743);
nand U7450 (N_7450,N_6478,N_6062);
or U7451 (N_7451,N_6125,N_6833);
nor U7452 (N_7452,N_6427,N_6537);
nor U7453 (N_7453,N_6622,N_6077);
nand U7454 (N_7454,N_6765,N_6384);
and U7455 (N_7455,N_6546,N_6097);
or U7456 (N_7456,N_6458,N_6742);
or U7457 (N_7457,N_6866,N_6589);
or U7458 (N_7458,N_6959,N_6246);
and U7459 (N_7459,N_6221,N_6171);
and U7460 (N_7460,N_6460,N_6398);
nand U7461 (N_7461,N_6597,N_6447);
or U7462 (N_7462,N_6553,N_6254);
or U7463 (N_7463,N_6096,N_6449);
and U7464 (N_7464,N_6094,N_6781);
nand U7465 (N_7465,N_6780,N_6307);
xnor U7466 (N_7466,N_6291,N_6856);
nor U7467 (N_7467,N_6396,N_6260);
or U7468 (N_7468,N_6805,N_6208);
and U7469 (N_7469,N_6884,N_6811);
and U7470 (N_7470,N_6308,N_6920);
nand U7471 (N_7471,N_6539,N_6411);
and U7472 (N_7472,N_6231,N_6885);
nor U7473 (N_7473,N_6201,N_6951);
nor U7474 (N_7474,N_6213,N_6258);
nand U7475 (N_7475,N_6955,N_6504);
nor U7476 (N_7476,N_6814,N_6559);
nor U7477 (N_7477,N_6495,N_6974);
nand U7478 (N_7478,N_6890,N_6011);
or U7479 (N_7479,N_6474,N_6154);
or U7480 (N_7480,N_6817,N_6268);
or U7481 (N_7481,N_6243,N_6390);
nand U7482 (N_7482,N_6859,N_6693);
and U7483 (N_7483,N_6958,N_6430);
and U7484 (N_7484,N_6175,N_6102);
nand U7485 (N_7485,N_6868,N_6117);
nor U7486 (N_7486,N_6190,N_6169);
and U7487 (N_7487,N_6709,N_6980);
nor U7488 (N_7488,N_6800,N_6178);
xor U7489 (N_7489,N_6340,N_6634);
or U7490 (N_7490,N_6533,N_6653);
or U7491 (N_7491,N_6370,N_6891);
and U7492 (N_7492,N_6771,N_6703);
or U7493 (N_7493,N_6786,N_6720);
nor U7494 (N_7494,N_6870,N_6596);
nand U7495 (N_7495,N_6672,N_6435);
or U7496 (N_7496,N_6376,N_6812);
or U7497 (N_7497,N_6392,N_6209);
or U7498 (N_7498,N_6215,N_6373);
or U7499 (N_7499,N_6189,N_6941);
nor U7500 (N_7500,N_6868,N_6772);
nor U7501 (N_7501,N_6307,N_6911);
or U7502 (N_7502,N_6220,N_6089);
nand U7503 (N_7503,N_6460,N_6447);
nand U7504 (N_7504,N_6919,N_6738);
or U7505 (N_7505,N_6660,N_6791);
nor U7506 (N_7506,N_6241,N_6289);
nor U7507 (N_7507,N_6144,N_6958);
nand U7508 (N_7508,N_6293,N_6677);
and U7509 (N_7509,N_6847,N_6087);
nand U7510 (N_7510,N_6338,N_6381);
or U7511 (N_7511,N_6520,N_6659);
nor U7512 (N_7512,N_6762,N_6275);
and U7513 (N_7513,N_6815,N_6026);
nand U7514 (N_7514,N_6581,N_6807);
and U7515 (N_7515,N_6835,N_6163);
nor U7516 (N_7516,N_6968,N_6278);
or U7517 (N_7517,N_6874,N_6584);
or U7518 (N_7518,N_6177,N_6991);
or U7519 (N_7519,N_6022,N_6096);
and U7520 (N_7520,N_6822,N_6889);
or U7521 (N_7521,N_6019,N_6560);
nor U7522 (N_7522,N_6432,N_6622);
nand U7523 (N_7523,N_6033,N_6085);
or U7524 (N_7524,N_6061,N_6552);
xnor U7525 (N_7525,N_6687,N_6574);
and U7526 (N_7526,N_6004,N_6831);
or U7527 (N_7527,N_6692,N_6682);
nor U7528 (N_7528,N_6953,N_6846);
and U7529 (N_7529,N_6047,N_6561);
and U7530 (N_7530,N_6289,N_6454);
nor U7531 (N_7531,N_6361,N_6210);
or U7532 (N_7532,N_6286,N_6963);
nand U7533 (N_7533,N_6964,N_6822);
nand U7534 (N_7534,N_6418,N_6715);
and U7535 (N_7535,N_6042,N_6249);
and U7536 (N_7536,N_6174,N_6782);
or U7537 (N_7537,N_6750,N_6662);
or U7538 (N_7538,N_6040,N_6074);
or U7539 (N_7539,N_6872,N_6309);
or U7540 (N_7540,N_6167,N_6331);
or U7541 (N_7541,N_6297,N_6754);
nor U7542 (N_7542,N_6856,N_6795);
or U7543 (N_7543,N_6190,N_6597);
and U7544 (N_7544,N_6947,N_6809);
nor U7545 (N_7545,N_6451,N_6940);
and U7546 (N_7546,N_6375,N_6856);
nor U7547 (N_7547,N_6608,N_6920);
nor U7548 (N_7548,N_6607,N_6790);
nor U7549 (N_7549,N_6480,N_6222);
nor U7550 (N_7550,N_6015,N_6780);
or U7551 (N_7551,N_6556,N_6249);
nand U7552 (N_7552,N_6536,N_6723);
and U7553 (N_7553,N_6743,N_6900);
nand U7554 (N_7554,N_6498,N_6455);
or U7555 (N_7555,N_6857,N_6973);
nor U7556 (N_7556,N_6093,N_6540);
nor U7557 (N_7557,N_6891,N_6271);
and U7558 (N_7558,N_6952,N_6652);
nand U7559 (N_7559,N_6548,N_6590);
and U7560 (N_7560,N_6766,N_6734);
nand U7561 (N_7561,N_6361,N_6950);
and U7562 (N_7562,N_6493,N_6284);
nand U7563 (N_7563,N_6081,N_6219);
nor U7564 (N_7564,N_6264,N_6977);
and U7565 (N_7565,N_6166,N_6364);
nand U7566 (N_7566,N_6811,N_6890);
nand U7567 (N_7567,N_6937,N_6875);
or U7568 (N_7568,N_6329,N_6495);
nor U7569 (N_7569,N_6055,N_6309);
and U7570 (N_7570,N_6667,N_6001);
and U7571 (N_7571,N_6691,N_6272);
or U7572 (N_7572,N_6245,N_6237);
or U7573 (N_7573,N_6360,N_6086);
nand U7574 (N_7574,N_6917,N_6002);
and U7575 (N_7575,N_6695,N_6728);
nand U7576 (N_7576,N_6275,N_6367);
or U7577 (N_7577,N_6525,N_6024);
nand U7578 (N_7578,N_6321,N_6754);
nor U7579 (N_7579,N_6641,N_6460);
nor U7580 (N_7580,N_6144,N_6362);
or U7581 (N_7581,N_6353,N_6895);
nor U7582 (N_7582,N_6695,N_6648);
or U7583 (N_7583,N_6546,N_6800);
and U7584 (N_7584,N_6183,N_6578);
or U7585 (N_7585,N_6802,N_6847);
and U7586 (N_7586,N_6282,N_6702);
and U7587 (N_7587,N_6494,N_6646);
nor U7588 (N_7588,N_6927,N_6126);
and U7589 (N_7589,N_6980,N_6433);
and U7590 (N_7590,N_6929,N_6643);
nand U7591 (N_7591,N_6889,N_6810);
nand U7592 (N_7592,N_6247,N_6058);
nor U7593 (N_7593,N_6393,N_6130);
and U7594 (N_7594,N_6378,N_6526);
nor U7595 (N_7595,N_6673,N_6793);
nor U7596 (N_7596,N_6460,N_6807);
xor U7597 (N_7597,N_6169,N_6159);
nand U7598 (N_7598,N_6381,N_6594);
and U7599 (N_7599,N_6591,N_6395);
or U7600 (N_7600,N_6902,N_6084);
nand U7601 (N_7601,N_6132,N_6362);
or U7602 (N_7602,N_6635,N_6258);
and U7603 (N_7603,N_6537,N_6687);
or U7604 (N_7604,N_6078,N_6547);
nor U7605 (N_7605,N_6301,N_6106);
or U7606 (N_7606,N_6902,N_6147);
or U7607 (N_7607,N_6701,N_6470);
nor U7608 (N_7608,N_6229,N_6300);
nand U7609 (N_7609,N_6857,N_6400);
nand U7610 (N_7610,N_6239,N_6940);
nor U7611 (N_7611,N_6293,N_6619);
nand U7612 (N_7612,N_6869,N_6864);
nor U7613 (N_7613,N_6195,N_6092);
and U7614 (N_7614,N_6867,N_6613);
nand U7615 (N_7615,N_6753,N_6154);
nand U7616 (N_7616,N_6274,N_6096);
nor U7617 (N_7617,N_6188,N_6222);
or U7618 (N_7618,N_6466,N_6105);
nor U7619 (N_7619,N_6031,N_6638);
or U7620 (N_7620,N_6840,N_6407);
nor U7621 (N_7621,N_6879,N_6489);
and U7622 (N_7622,N_6090,N_6921);
or U7623 (N_7623,N_6004,N_6578);
nand U7624 (N_7624,N_6263,N_6820);
nor U7625 (N_7625,N_6048,N_6502);
and U7626 (N_7626,N_6997,N_6952);
or U7627 (N_7627,N_6161,N_6134);
nand U7628 (N_7628,N_6727,N_6410);
and U7629 (N_7629,N_6621,N_6141);
nand U7630 (N_7630,N_6831,N_6457);
nor U7631 (N_7631,N_6806,N_6209);
or U7632 (N_7632,N_6951,N_6613);
or U7633 (N_7633,N_6829,N_6987);
nand U7634 (N_7634,N_6834,N_6598);
or U7635 (N_7635,N_6482,N_6074);
or U7636 (N_7636,N_6561,N_6142);
nor U7637 (N_7637,N_6970,N_6417);
or U7638 (N_7638,N_6338,N_6502);
and U7639 (N_7639,N_6687,N_6201);
nand U7640 (N_7640,N_6599,N_6794);
or U7641 (N_7641,N_6859,N_6476);
nand U7642 (N_7642,N_6257,N_6845);
nand U7643 (N_7643,N_6376,N_6019);
nor U7644 (N_7644,N_6620,N_6859);
and U7645 (N_7645,N_6214,N_6589);
nand U7646 (N_7646,N_6776,N_6915);
xor U7647 (N_7647,N_6457,N_6204);
and U7648 (N_7648,N_6980,N_6559);
or U7649 (N_7649,N_6797,N_6409);
nor U7650 (N_7650,N_6290,N_6332);
nand U7651 (N_7651,N_6649,N_6293);
nand U7652 (N_7652,N_6414,N_6799);
nand U7653 (N_7653,N_6278,N_6551);
or U7654 (N_7654,N_6081,N_6089);
or U7655 (N_7655,N_6260,N_6835);
nand U7656 (N_7656,N_6810,N_6778);
xnor U7657 (N_7657,N_6638,N_6006);
nand U7658 (N_7658,N_6384,N_6842);
nand U7659 (N_7659,N_6972,N_6459);
nor U7660 (N_7660,N_6741,N_6467);
or U7661 (N_7661,N_6287,N_6676);
nor U7662 (N_7662,N_6349,N_6539);
and U7663 (N_7663,N_6424,N_6660);
nand U7664 (N_7664,N_6479,N_6835);
and U7665 (N_7665,N_6260,N_6395);
nor U7666 (N_7666,N_6712,N_6844);
nand U7667 (N_7667,N_6740,N_6343);
nor U7668 (N_7668,N_6885,N_6826);
and U7669 (N_7669,N_6393,N_6631);
nand U7670 (N_7670,N_6830,N_6813);
nor U7671 (N_7671,N_6828,N_6894);
or U7672 (N_7672,N_6931,N_6106);
nand U7673 (N_7673,N_6162,N_6466);
or U7674 (N_7674,N_6478,N_6066);
or U7675 (N_7675,N_6054,N_6317);
or U7676 (N_7676,N_6982,N_6704);
and U7677 (N_7677,N_6110,N_6770);
nand U7678 (N_7678,N_6257,N_6881);
and U7679 (N_7679,N_6203,N_6109);
nand U7680 (N_7680,N_6765,N_6169);
and U7681 (N_7681,N_6923,N_6782);
nor U7682 (N_7682,N_6893,N_6536);
and U7683 (N_7683,N_6622,N_6066);
nor U7684 (N_7684,N_6482,N_6346);
or U7685 (N_7685,N_6333,N_6182);
or U7686 (N_7686,N_6472,N_6278);
and U7687 (N_7687,N_6902,N_6194);
nand U7688 (N_7688,N_6660,N_6783);
or U7689 (N_7689,N_6904,N_6529);
and U7690 (N_7690,N_6443,N_6868);
and U7691 (N_7691,N_6122,N_6975);
nor U7692 (N_7692,N_6624,N_6401);
nor U7693 (N_7693,N_6506,N_6104);
or U7694 (N_7694,N_6912,N_6038);
and U7695 (N_7695,N_6892,N_6612);
and U7696 (N_7696,N_6692,N_6768);
and U7697 (N_7697,N_6417,N_6926);
nand U7698 (N_7698,N_6776,N_6177);
or U7699 (N_7699,N_6349,N_6696);
or U7700 (N_7700,N_6188,N_6116);
and U7701 (N_7701,N_6490,N_6941);
nand U7702 (N_7702,N_6454,N_6207);
or U7703 (N_7703,N_6140,N_6345);
nand U7704 (N_7704,N_6594,N_6703);
nand U7705 (N_7705,N_6263,N_6447);
nor U7706 (N_7706,N_6175,N_6208);
and U7707 (N_7707,N_6692,N_6741);
nand U7708 (N_7708,N_6023,N_6158);
and U7709 (N_7709,N_6043,N_6910);
and U7710 (N_7710,N_6207,N_6809);
and U7711 (N_7711,N_6148,N_6099);
or U7712 (N_7712,N_6423,N_6377);
or U7713 (N_7713,N_6302,N_6703);
and U7714 (N_7714,N_6836,N_6899);
nor U7715 (N_7715,N_6717,N_6955);
or U7716 (N_7716,N_6301,N_6413);
xor U7717 (N_7717,N_6758,N_6691);
nor U7718 (N_7718,N_6201,N_6177);
or U7719 (N_7719,N_6306,N_6381);
nand U7720 (N_7720,N_6005,N_6527);
nand U7721 (N_7721,N_6270,N_6463);
nor U7722 (N_7722,N_6158,N_6263);
and U7723 (N_7723,N_6047,N_6929);
nor U7724 (N_7724,N_6780,N_6270);
or U7725 (N_7725,N_6907,N_6429);
or U7726 (N_7726,N_6185,N_6415);
or U7727 (N_7727,N_6455,N_6509);
and U7728 (N_7728,N_6772,N_6715);
or U7729 (N_7729,N_6886,N_6819);
nand U7730 (N_7730,N_6124,N_6150);
or U7731 (N_7731,N_6787,N_6363);
or U7732 (N_7732,N_6766,N_6662);
and U7733 (N_7733,N_6115,N_6009);
or U7734 (N_7734,N_6268,N_6621);
nor U7735 (N_7735,N_6423,N_6293);
nand U7736 (N_7736,N_6596,N_6903);
or U7737 (N_7737,N_6325,N_6416);
nor U7738 (N_7738,N_6487,N_6213);
and U7739 (N_7739,N_6206,N_6312);
and U7740 (N_7740,N_6352,N_6677);
nand U7741 (N_7741,N_6437,N_6490);
nor U7742 (N_7742,N_6930,N_6766);
and U7743 (N_7743,N_6268,N_6987);
nand U7744 (N_7744,N_6722,N_6491);
nand U7745 (N_7745,N_6706,N_6788);
nand U7746 (N_7746,N_6007,N_6954);
and U7747 (N_7747,N_6669,N_6583);
nand U7748 (N_7748,N_6811,N_6777);
and U7749 (N_7749,N_6292,N_6305);
nand U7750 (N_7750,N_6997,N_6833);
nand U7751 (N_7751,N_6352,N_6159);
nand U7752 (N_7752,N_6746,N_6439);
and U7753 (N_7753,N_6116,N_6593);
and U7754 (N_7754,N_6353,N_6864);
nor U7755 (N_7755,N_6305,N_6991);
and U7756 (N_7756,N_6778,N_6099);
nor U7757 (N_7757,N_6167,N_6415);
or U7758 (N_7758,N_6006,N_6673);
nor U7759 (N_7759,N_6390,N_6043);
nor U7760 (N_7760,N_6096,N_6060);
or U7761 (N_7761,N_6655,N_6683);
and U7762 (N_7762,N_6386,N_6226);
and U7763 (N_7763,N_6866,N_6015);
nand U7764 (N_7764,N_6807,N_6604);
nor U7765 (N_7765,N_6672,N_6866);
nor U7766 (N_7766,N_6415,N_6206);
xor U7767 (N_7767,N_6804,N_6246);
or U7768 (N_7768,N_6812,N_6655);
and U7769 (N_7769,N_6621,N_6792);
nand U7770 (N_7770,N_6743,N_6539);
or U7771 (N_7771,N_6315,N_6004);
and U7772 (N_7772,N_6860,N_6312);
or U7773 (N_7773,N_6339,N_6381);
or U7774 (N_7774,N_6384,N_6768);
nor U7775 (N_7775,N_6155,N_6553);
and U7776 (N_7776,N_6086,N_6084);
or U7777 (N_7777,N_6931,N_6630);
nand U7778 (N_7778,N_6507,N_6939);
or U7779 (N_7779,N_6702,N_6183);
nand U7780 (N_7780,N_6143,N_6004);
nand U7781 (N_7781,N_6428,N_6670);
nand U7782 (N_7782,N_6725,N_6325);
or U7783 (N_7783,N_6087,N_6964);
and U7784 (N_7784,N_6375,N_6975);
nand U7785 (N_7785,N_6649,N_6067);
or U7786 (N_7786,N_6541,N_6568);
or U7787 (N_7787,N_6179,N_6724);
nand U7788 (N_7788,N_6614,N_6147);
nor U7789 (N_7789,N_6525,N_6537);
nand U7790 (N_7790,N_6904,N_6836);
nor U7791 (N_7791,N_6931,N_6225);
nand U7792 (N_7792,N_6310,N_6433);
or U7793 (N_7793,N_6655,N_6312);
and U7794 (N_7794,N_6559,N_6533);
nor U7795 (N_7795,N_6855,N_6358);
nor U7796 (N_7796,N_6014,N_6910);
nand U7797 (N_7797,N_6139,N_6572);
nand U7798 (N_7798,N_6853,N_6675);
nor U7799 (N_7799,N_6059,N_6231);
nand U7800 (N_7800,N_6515,N_6586);
nor U7801 (N_7801,N_6049,N_6006);
and U7802 (N_7802,N_6552,N_6343);
or U7803 (N_7803,N_6345,N_6083);
or U7804 (N_7804,N_6225,N_6420);
or U7805 (N_7805,N_6358,N_6613);
or U7806 (N_7806,N_6771,N_6370);
nand U7807 (N_7807,N_6310,N_6319);
xnor U7808 (N_7808,N_6843,N_6090);
and U7809 (N_7809,N_6514,N_6167);
and U7810 (N_7810,N_6669,N_6388);
or U7811 (N_7811,N_6980,N_6921);
nand U7812 (N_7812,N_6338,N_6624);
nand U7813 (N_7813,N_6153,N_6628);
nand U7814 (N_7814,N_6545,N_6554);
nor U7815 (N_7815,N_6180,N_6757);
or U7816 (N_7816,N_6904,N_6739);
and U7817 (N_7817,N_6525,N_6926);
or U7818 (N_7818,N_6363,N_6726);
nand U7819 (N_7819,N_6026,N_6868);
and U7820 (N_7820,N_6264,N_6689);
or U7821 (N_7821,N_6126,N_6407);
or U7822 (N_7822,N_6024,N_6495);
nand U7823 (N_7823,N_6879,N_6311);
and U7824 (N_7824,N_6451,N_6258);
or U7825 (N_7825,N_6393,N_6176);
nand U7826 (N_7826,N_6853,N_6218);
nand U7827 (N_7827,N_6086,N_6990);
or U7828 (N_7828,N_6794,N_6506);
and U7829 (N_7829,N_6003,N_6157);
nand U7830 (N_7830,N_6323,N_6223);
nand U7831 (N_7831,N_6267,N_6177);
nand U7832 (N_7832,N_6527,N_6393);
and U7833 (N_7833,N_6976,N_6160);
nand U7834 (N_7834,N_6480,N_6463);
or U7835 (N_7835,N_6885,N_6388);
and U7836 (N_7836,N_6597,N_6188);
or U7837 (N_7837,N_6722,N_6855);
and U7838 (N_7838,N_6297,N_6286);
and U7839 (N_7839,N_6396,N_6994);
nand U7840 (N_7840,N_6823,N_6897);
xnor U7841 (N_7841,N_6748,N_6205);
or U7842 (N_7842,N_6766,N_6141);
and U7843 (N_7843,N_6613,N_6161);
nand U7844 (N_7844,N_6320,N_6472);
and U7845 (N_7845,N_6047,N_6805);
and U7846 (N_7846,N_6136,N_6659);
or U7847 (N_7847,N_6546,N_6658);
and U7848 (N_7848,N_6641,N_6044);
or U7849 (N_7849,N_6938,N_6962);
or U7850 (N_7850,N_6618,N_6961);
nand U7851 (N_7851,N_6271,N_6389);
nand U7852 (N_7852,N_6588,N_6221);
nand U7853 (N_7853,N_6284,N_6652);
nand U7854 (N_7854,N_6513,N_6502);
nor U7855 (N_7855,N_6033,N_6496);
or U7856 (N_7856,N_6896,N_6511);
or U7857 (N_7857,N_6624,N_6008);
nand U7858 (N_7858,N_6971,N_6544);
nor U7859 (N_7859,N_6419,N_6901);
and U7860 (N_7860,N_6929,N_6642);
or U7861 (N_7861,N_6607,N_6152);
or U7862 (N_7862,N_6767,N_6952);
and U7863 (N_7863,N_6874,N_6005);
and U7864 (N_7864,N_6445,N_6281);
nor U7865 (N_7865,N_6835,N_6104);
xnor U7866 (N_7866,N_6317,N_6097);
or U7867 (N_7867,N_6010,N_6260);
nand U7868 (N_7868,N_6676,N_6592);
nand U7869 (N_7869,N_6470,N_6529);
and U7870 (N_7870,N_6463,N_6894);
and U7871 (N_7871,N_6669,N_6774);
and U7872 (N_7872,N_6766,N_6243);
nor U7873 (N_7873,N_6874,N_6305);
nor U7874 (N_7874,N_6199,N_6064);
nand U7875 (N_7875,N_6478,N_6751);
nor U7876 (N_7876,N_6564,N_6718);
or U7877 (N_7877,N_6502,N_6817);
nand U7878 (N_7878,N_6586,N_6311);
nand U7879 (N_7879,N_6516,N_6897);
nor U7880 (N_7880,N_6534,N_6087);
and U7881 (N_7881,N_6031,N_6403);
nor U7882 (N_7882,N_6907,N_6490);
nand U7883 (N_7883,N_6187,N_6000);
and U7884 (N_7884,N_6349,N_6809);
or U7885 (N_7885,N_6171,N_6063);
nor U7886 (N_7886,N_6396,N_6543);
nor U7887 (N_7887,N_6761,N_6358);
or U7888 (N_7888,N_6642,N_6065);
nor U7889 (N_7889,N_6453,N_6947);
or U7890 (N_7890,N_6964,N_6370);
and U7891 (N_7891,N_6961,N_6583);
nand U7892 (N_7892,N_6653,N_6569);
nor U7893 (N_7893,N_6232,N_6099);
nor U7894 (N_7894,N_6860,N_6157);
or U7895 (N_7895,N_6569,N_6709);
nor U7896 (N_7896,N_6558,N_6396);
and U7897 (N_7897,N_6786,N_6459);
nor U7898 (N_7898,N_6836,N_6507);
nor U7899 (N_7899,N_6380,N_6555);
and U7900 (N_7900,N_6806,N_6384);
nand U7901 (N_7901,N_6654,N_6326);
or U7902 (N_7902,N_6388,N_6527);
nor U7903 (N_7903,N_6083,N_6579);
and U7904 (N_7904,N_6347,N_6338);
nand U7905 (N_7905,N_6153,N_6727);
nand U7906 (N_7906,N_6194,N_6082);
nand U7907 (N_7907,N_6131,N_6034);
nand U7908 (N_7908,N_6832,N_6395);
nor U7909 (N_7909,N_6865,N_6303);
or U7910 (N_7910,N_6076,N_6255);
nor U7911 (N_7911,N_6564,N_6926);
nor U7912 (N_7912,N_6206,N_6685);
or U7913 (N_7913,N_6627,N_6076);
or U7914 (N_7914,N_6879,N_6138);
and U7915 (N_7915,N_6275,N_6769);
nor U7916 (N_7916,N_6837,N_6383);
and U7917 (N_7917,N_6420,N_6564);
and U7918 (N_7918,N_6163,N_6700);
nor U7919 (N_7919,N_6208,N_6800);
or U7920 (N_7920,N_6472,N_6160);
or U7921 (N_7921,N_6877,N_6866);
nor U7922 (N_7922,N_6429,N_6998);
or U7923 (N_7923,N_6228,N_6884);
nor U7924 (N_7924,N_6801,N_6420);
nand U7925 (N_7925,N_6589,N_6181);
and U7926 (N_7926,N_6375,N_6621);
nor U7927 (N_7927,N_6325,N_6912);
and U7928 (N_7928,N_6961,N_6535);
nor U7929 (N_7929,N_6024,N_6433);
nor U7930 (N_7930,N_6253,N_6738);
nor U7931 (N_7931,N_6649,N_6504);
and U7932 (N_7932,N_6932,N_6739);
or U7933 (N_7933,N_6129,N_6610);
or U7934 (N_7934,N_6907,N_6090);
or U7935 (N_7935,N_6328,N_6899);
and U7936 (N_7936,N_6534,N_6426);
and U7937 (N_7937,N_6731,N_6724);
nand U7938 (N_7938,N_6791,N_6438);
and U7939 (N_7939,N_6973,N_6685);
or U7940 (N_7940,N_6094,N_6293);
xnor U7941 (N_7941,N_6898,N_6385);
xor U7942 (N_7942,N_6827,N_6278);
and U7943 (N_7943,N_6183,N_6637);
nor U7944 (N_7944,N_6185,N_6864);
and U7945 (N_7945,N_6410,N_6044);
nor U7946 (N_7946,N_6963,N_6096);
and U7947 (N_7947,N_6400,N_6016);
xor U7948 (N_7948,N_6974,N_6878);
or U7949 (N_7949,N_6932,N_6418);
or U7950 (N_7950,N_6031,N_6708);
and U7951 (N_7951,N_6380,N_6468);
nand U7952 (N_7952,N_6408,N_6276);
nand U7953 (N_7953,N_6260,N_6414);
nand U7954 (N_7954,N_6330,N_6364);
nor U7955 (N_7955,N_6720,N_6420);
nor U7956 (N_7956,N_6119,N_6584);
xor U7957 (N_7957,N_6903,N_6384);
nand U7958 (N_7958,N_6013,N_6848);
nand U7959 (N_7959,N_6451,N_6416);
xor U7960 (N_7960,N_6036,N_6125);
nor U7961 (N_7961,N_6398,N_6465);
or U7962 (N_7962,N_6732,N_6121);
nand U7963 (N_7963,N_6587,N_6981);
and U7964 (N_7964,N_6556,N_6131);
nand U7965 (N_7965,N_6087,N_6930);
and U7966 (N_7966,N_6099,N_6390);
and U7967 (N_7967,N_6440,N_6892);
or U7968 (N_7968,N_6398,N_6836);
and U7969 (N_7969,N_6153,N_6109);
or U7970 (N_7970,N_6169,N_6048);
or U7971 (N_7971,N_6924,N_6789);
or U7972 (N_7972,N_6621,N_6710);
and U7973 (N_7973,N_6401,N_6034);
nand U7974 (N_7974,N_6719,N_6096);
nand U7975 (N_7975,N_6437,N_6745);
or U7976 (N_7976,N_6766,N_6332);
nor U7977 (N_7977,N_6050,N_6940);
nor U7978 (N_7978,N_6313,N_6708);
or U7979 (N_7979,N_6000,N_6166);
nand U7980 (N_7980,N_6309,N_6075);
or U7981 (N_7981,N_6801,N_6910);
and U7982 (N_7982,N_6616,N_6899);
and U7983 (N_7983,N_6539,N_6556);
nand U7984 (N_7984,N_6325,N_6373);
nor U7985 (N_7985,N_6949,N_6805);
nand U7986 (N_7986,N_6282,N_6332);
nand U7987 (N_7987,N_6745,N_6402);
nand U7988 (N_7988,N_6359,N_6149);
and U7989 (N_7989,N_6237,N_6470);
and U7990 (N_7990,N_6232,N_6856);
or U7991 (N_7991,N_6242,N_6597);
or U7992 (N_7992,N_6965,N_6552);
and U7993 (N_7993,N_6871,N_6020);
nor U7994 (N_7994,N_6017,N_6668);
nor U7995 (N_7995,N_6843,N_6928);
nand U7996 (N_7996,N_6249,N_6402);
or U7997 (N_7997,N_6618,N_6585);
nand U7998 (N_7998,N_6919,N_6895);
or U7999 (N_7999,N_6514,N_6202);
and U8000 (N_8000,N_7851,N_7827);
nor U8001 (N_8001,N_7937,N_7835);
and U8002 (N_8002,N_7706,N_7503);
and U8003 (N_8003,N_7923,N_7408);
nand U8004 (N_8004,N_7523,N_7529);
or U8005 (N_8005,N_7838,N_7443);
nor U8006 (N_8006,N_7048,N_7386);
and U8007 (N_8007,N_7362,N_7670);
nand U8008 (N_8008,N_7546,N_7277);
and U8009 (N_8009,N_7571,N_7493);
nor U8010 (N_8010,N_7820,N_7289);
nor U8011 (N_8011,N_7790,N_7601);
nand U8012 (N_8012,N_7707,N_7662);
nor U8013 (N_8013,N_7795,N_7187);
nand U8014 (N_8014,N_7673,N_7936);
nand U8015 (N_8015,N_7957,N_7946);
nor U8016 (N_8016,N_7919,N_7881);
xor U8017 (N_8017,N_7448,N_7489);
nor U8018 (N_8018,N_7251,N_7532);
nor U8019 (N_8019,N_7732,N_7243);
nor U8020 (N_8020,N_7276,N_7176);
and U8021 (N_8021,N_7792,N_7294);
or U8022 (N_8022,N_7457,N_7093);
and U8023 (N_8023,N_7070,N_7181);
and U8024 (N_8024,N_7085,N_7623);
or U8025 (N_8025,N_7814,N_7422);
nor U8026 (N_8026,N_7863,N_7885);
nand U8027 (N_8027,N_7679,N_7620);
nand U8028 (N_8028,N_7803,N_7375);
nand U8029 (N_8029,N_7752,N_7001);
nand U8030 (N_8030,N_7029,N_7495);
and U8031 (N_8031,N_7008,N_7369);
and U8032 (N_8032,N_7855,N_7105);
or U8033 (N_8033,N_7870,N_7753);
and U8034 (N_8034,N_7607,N_7904);
and U8035 (N_8035,N_7939,N_7500);
nor U8036 (N_8036,N_7134,N_7877);
or U8037 (N_8037,N_7406,N_7960);
nor U8038 (N_8038,N_7226,N_7565);
nand U8039 (N_8039,N_7195,N_7638);
nor U8040 (N_8040,N_7608,N_7157);
and U8041 (N_8041,N_7050,N_7247);
and U8042 (N_8042,N_7568,N_7393);
nor U8043 (N_8043,N_7983,N_7279);
nand U8044 (N_8044,N_7480,N_7065);
nand U8045 (N_8045,N_7127,N_7669);
and U8046 (N_8046,N_7668,N_7124);
nor U8047 (N_8047,N_7179,N_7521);
nand U8048 (N_8048,N_7793,N_7929);
or U8049 (N_8049,N_7367,N_7190);
and U8050 (N_8050,N_7522,N_7817);
or U8051 (N_8051,N_7713,N_7501);
or U8052 (N_8052,N_7206,N_7297);
or U8053 (N_8053,N_7321,N_7429);
nor U8054 (N_8054,N_7789,N_7990);
nor U8055 (N_8055,N_7126,N_7976);
and U8056 (N_8056,N_7117,N_7557);
and U8057 (N_8057,N_7802,N_7760);
nand U8058 (N_8058,N_7116,N_7841);
nor U8059 (N_8059,N_7512,N_7016);
nor U8060 (N_8060,N_7705,N_7524);
or U8061 (N_8061,N_7862,N_7384);
and U8062 (N_8062,N_7040,N_7428);
nor U8063 (N_8063,N_7007,N_7371);
or U8064 (N_8064,N_7080,N_7824);
nor U8065 (N_8065,N_7242,N_7472);
nor U8066 (N_8066,N_7028,N_7166);
and U8067 (N_8067,N_7373,N_7858);
and U8068 (N_8068,N_7951,N_7041);
or U8069 (N_8069,N_7423,N_7054);
or U8070 (N_8070,N_7777,N_7746);
nand U8071 (N_8071,N_7391,N_7685);
or U8072 (N_8072,N_7628,N_7142);
or U8073 (N_8073,N_7376,N_7515);
nand U8074 (N_8074,N_7214,N_7337);
xnor U8075 (N_8075,N_7053,N_7101);
nor U8076 (N_8076,N_7823,N_7184);
and U8077 (N_8077,N_7551,N_7119);
nor U8078 (N_8078,N_7261,N_7811);
nand U8079 (N_8079,N_7916,N_7306);
nand U8080 (N_8080,N_7934,N_7970);
nand U8081 (N_8081,N_7043,N_7879);
or U8082 (N_8082,N_7924,N_7664);
or U8083 (N_8083,N_7897,N_7785);
or U8084 (N_8084,N_7398,N_7316);
nand U8085 (N_8085,N_7766,N_7025);
nand U8086 (N_8086,N_7816,N_7368);
or U8087 (N_8087,N_7658,N_7599);
nand U8088 (N_8088,N_7971,N_7490);
nand U8089 (N_8089,N_7241,N_7612);
nand U8090 (N_8090,N_7891,N_7107);
nand U8091 (N_8091,N_7477,N_7909);
xor U8092 (N_8092,N_7992,N_7009);
or U8093 (N_8093,N_7458,N_7562);
or U8094 (N_8094,N_7921,N_7901);
or U8095 (N_8095,N_7530,N_7852);
or U8096 (N_8096,N_7847,N_7868);
nand U8097 (N_8097,N_7483,N_7436);
nand U8098 (N_8098,N_7697,N_7613);
nand U8099 (N_8099,N_7572,N_7022);
or U8100 (N_8100,N_7060,N_7010);
and U8101 (N_8101,N_7514,N_7587);
or U8102 (N_8102,N_7889,N_7660);
nor U8103 (N_8103,N_7087,N_7118);
and U8104 (N_8104,N_7584,N_7412);
nor U8105 (N_8105,N_7162,N_7736);
nand U8106 (N_8106,N_7420,N_7636);
and U8107 (N_8107,N_7558,N_7005);
nor U8108 (N_8108,N_7191,N_7433);
nor U8109 (N_8109,N_7577,N_7606);
nand U8110 (N_8110,N_7950,N_7164);
nor U8111 (N_8111,N_7399,N_7594);
xor U8112 (N_8112,N_7309,N_7357);
nor U8113 (N_8113,N_7273,N_7459);
nand U8114 (N_8114,N_7938,N_7940);
nand U8115 (N_8115,N_7567,N_7962);
nor U8116 (N_8116,N_7517,N_7447);
and U8117 (N_8117,N_7775,N_7439);
and U8118 (N_8118,N_7017,N_7890);
nand U8119 (N_8119,N_7570,N_7254);
and U8120 (N_8120,N_7407,N_7026);
nor U8121 (N_8121,N_7583,N_7544);
or U8122 (N_8122,N_7298,N_7268);
nor U8123 (N_8123,N_7895,N_7278);
nor U8124 (N_8124,N_7350,N_7286);
and U8125 (N_8125,N_7073,N_7002);
and U8126 (N_8126,N_7536,N_7339);
nor U8127 (N_8127,N_7061,N_7066);
and U8128 (N_8128,N_7762,N_7663);
nor U8129 (N_8129,N_7138,N_7171);
nor U8130 (N_8130,N_7013,N_7351);
nand U8131 (N_8131,N_7382,N_7682);
and U8132 (N_8132,N_7733,N_7481);
or U8133 (N_8133,N_7759,N_7322);
xor U8134 (N_8134,N_7100,N_7131);
and U8135 (N_8135,N_7989,N_7588);
and U8136 (N_8136,N_7293,N_7011);
and U8137 (N_8137,N_7945,N_7084);
nand U8138 (N_8138,N_7069,N_7036);
or U8139 (N_8139,N_7754,N_7857);
and U8140 (N_8140,N_7200,N_7192);
or U8141 (N_8141,N_7262,N_7220);
and U8142 (N_8142,N_7353,N_7019);
nand U8143 (N_8143,N_7692,N_7260);
and U8144 (N_8144,N_7738,N_7215);
nand U8145 (N_8145,N_7888,N_7642);
or U8146 (N_8146,N_7854,N_7747);
or U8147 (N_8147,N_7083,N_7499);
nor U8148 (N_8148,N_7987,N_7378);
nor U8149 (N_8149,N_7604,N_7056);
nand U8150 (N_8150,N_7963,N_7426);
nand U8151 (N_8151,N_7033,N_7155);
or U8152 (N_8152,N_7829,N_7074);
nor U8153 (N_8153,N_7462,N_7504);
and U8154 (N_8154,N_7358,N_7218);
or U8155 (N_8155,N_7227,N_7198);
nand U8156 (N_8156,N_7819,N_7641);
nor U8157 (N_8157,N_7973,N_7235);
and U8158 (N_8158,N_7619,N_7264);
nand U8159 (N_8159,N_7096,N_7898);
or U8160 (N_8160,N_7640,N_7566);
and U8161 (N_8161,N_7874,N_7534);
nand U8162 (N_8162,N_7219,N_7645);
and U8163 (N_8163,N_7346,N_7609);
or U8164 (N_8164,N_7781,N_7552);
xnor U8165 (N_8165,N_7094,N_7072);
nand U8166 (N_8166,N_7238,N_7441);
and U8167 (N_8167,N_7849,N_7912);
nor U8168 (N_8168,N_7341,N_7304);
nand U8169 (N_8169,N_7637,N_7284);
nand U8170 (N_8170,N_7834,N_7977);
nand U8171 (N_8171,N_7632,N_7086);
nand U8172 (N_8172,N_7123,N_7867);
or U8173 (N_8173,N_7463,N_7768);
nor U8174 (N_8174,N_7130,N_7342);
or U8175 (N_8175,N_7751,N_7804);
nand U8176 (N_8176,N_7696,N_7914);
nor U8177 (N_8177,N_7366,N_7108);
or U8178 (N_8178,N_7161,N_7794);
or U8179 (N_8179,N_7791,N_7699);
nand U8180 (N_8180,N_7224,N_7132);
nor U8181 (N_8181,N_7401,N_7385);
and U8182 (N_8182,N_7216,N_7797);
nor U8183 (N_8183,N_7338,N_7694);
nor U8184 (N_8184,N_7465,N_7869);
nand U8185 (N_8185,N_7763,N_7943);
or U8186 (N_8186,N_7000,N_7389);
nand U8187 (N_8187,N_7466,N_7853);
and U8188 (N_8188,N_7948,N_7639);
or U8189 (N_8189,N_7556,N_7656);
nor U8190 (N_8190,N_7303,N_7807);
nor U8191 (N_8191,N_7347,N_7249);
or U8192 (N_8192,N_7431,N_7169);
and U8193 (N_8193,N_7875,N_7240);
or U8194 (N_8194,N_7605,N_7329);
or U8195 (N_8195,N_7246,N_7614);
and U8196 (N_8196,N_7941,N_7442);
or U8197 (N_8197,N_7896,N_7648);
and U8198 (N_8198,N_7248,N_7310);
nand U8199 (N_8199,N_7984,N_7404);
or U8200 (N_8200,N_7545,N_7295);
and U8201 (N_8201,N_7880,N_7933);
or U8202 (N_8202,N_7674,N_7892);
xnor U8203 (N_8203,N_7727,N_7438);
nand U8204 (N_8204,N_7182,N_7801);
nor U8205 (N_8205,N_7311,N_7030);
and U8206 (N_8206,N_7403,N_7947);
or U8207 (N_8207,N_7655,N_7413);
or U8208 (N_8208,N_7830,N_7505);
nand U8209 (N_8209,N_7742,N_7223);
and U8210 (N_8210,N_7654,N_7905);
and U8211 (N_8211,N_7764,N_7773);
xnor U8212 (N_8212,N_7509,N_7245);
nor U8213 (N_8213,N_7721,N_7460);
and U8214 (N_8214,N_7396,N_7133);
or U8215 (N_8215,N_7475,N_7954);
nor U8216 (N_8216,N_7405,N_7313);
and U8217 (N_8217,N_7272,N_7774);
nand U8218 (N_8218,N_7917,N_7174);
nand U8219 (N_8219,N_7724,N_7569);
and U8220 (N_8220,N_7837,N_7708);
nand U8221 (N_8221,N_7221,N_7045);
nor U8222 (N_8222,N_7267,N_7996);
xnor U8223 (N_8223,N_7319,N_7856);
nand U8224 (N_8224,N_7831,N_7330);
nor U8225 (N_8225,N_7893,N_7709);
or U8226 (N_8226,N_7952,N_7815);
and U8227 (N_8227,N_7003,N_7213);
or U8228 (N_8228,N_7550,N_7843);
and U8229 (N_8229,N_7488,N_7497);
and U8230 (N_8230,N_7666,N_7236);
and U8231 (N_8231,N_7553,N_7149);
nand U8232 (N_8232,N_7334,N_7519);
or U8233 (N_8233,N_7111,N_7474);
or U8234 (N_8234,N_7626,N_7986);
nand U8235 (N_8235,N_7826,N_7145);
or U8236 (N_8236,N_7031,N_7998);
nand U8237 (N_8237,N_7115,N_7361);
and U8238 (N_8238,N_7450,N_7095);
and U8239 (N_8239,N_7578,N_7547);
nand U8240 (N_8240,N_7427,N_7180);
nor U8241 (N_8241,N_7994,N_7717);
or U8242 (N_8242,N_7381,N_7210);
nor U8243 (N_8243,N_7106,N_7675);
nor U8244 (N_8244,N_7435,N_7528);
or U8245 (N_8245,N_7091,N_7907);
nand U8246 (N_8246,N_7549,N_7209);
or U8247 (N_8247,N_7078,N_7445);
and U8248 (N_8248,N_7315,N_7822);
nand U8249 (N_8249,N_7740,N_7365);
nor U8250 (N_8250,N_7518,N_7038);
or U8251 (N_8251,N_7006,N_7769);
nand U8252 (N_8252,N_7370,N_7643);
nor U8253 (N_8253,N_7991,N_7538);
and U8254 (N_8254,N_7920,N_7222);
nor U8255 (N_8255,N_7300,N_7424);
or U8256 (N_8256,N_7308,N_7484);
nor U8257 (N_8257,N_7354,N_7743);
nand U8258 (N_8258,N_7592,N_7511);
nor U8259 (N_8259,N_7531,N_7148);
xnor U8260 (N_8260,N_7416,N_7114);
and U8261 (N_8261,N_7681,N_7395);
nand U8262 (N_8262,N_7652,N_7884);
nand U8263 (N_8263,N_7756,N_7507);
nand U8264 (N_8264,N_7363,N_7098);
nor U8265 (N_8265,N_7141,N_7014);
nor U8266 (N_8266,N_7324,N_7312);
nor U8267 (N_8267,N_7502,N_7980);
and U8268 (N_8268,N_7906,N_7902);
nor U8269 (N_8269,N_7335,N_7748);
nor U8270 (N_8270,N_7672,N_7799);
nand U8271 (N_8271,N_7492,N_7352);
and U8272 (N_8272,N_7023,N_7621);
nand U8273 (N_8273,N_7812,N_7104);
nand U8274 (N_8274,N_7355,N_7018);
and U8275 (N_8275,N_7199,N_7320);
or U8276 (N_8276,N_7788,N_7051);
nor U8277 (N_8277,N_7899,N_7269);
or U8278 (N_8278,N_7274,N_7446);
nor U8279 (N_8279,N_7090,N_7786);
nor U8280 (N_8280,N_7318,N_7903);
or U8281 (N_8281,N_7972,N_7156);
and U8282 (N_8282,N_7876,N_7981);
nand U8283 (N_8283,N_7735,N_7964);
or U8284 (N_8284,N_7930,N_7110);
or U8285 (N_8285,N_7478,N_7861);
nand U8286 (N_8286,N_7471,N_7581);
nand U8287 (N_8287,N_7927,N_7202);
or U8288 (N_8288,N_7539,N_7633);
or U8289 (N_8289,N_7122,N_7932);
or U8290 (N_8290,N_7183,N_7228);
and U8291 (N_8291,N_7715,N_7402);
or U8292 (N_8292,N_7167,N_7840);
nor U8293 (N_8293,N_7301,N_7255);
and U8294 (N_8294,N_7741,N_7582);
nor U8295 (N_8295,N_7667,N_7808);
nor U8296 (N_8296,N_7173,N_7886);
nand U8297 (N_8297,N_7392,N_7653);
nand U8298 (N_8298,N_7757,N_7437);
nor U8299 (N_8299,N_7958,N_7288);
nand U8300 (N_8300,N_7783,N_7170);
or U8301 (N_8301,N_7575,N_7409);
and U8302 (N_8302,N_7676,N_7340);
nand U8303 (N_8303,N_7453,N_7510);
nor U8304 (N_8304,N_7800,N_7969);
or U8305 (N_8305,N_7178,N_7563);
nand U8306 (N_8306,N_7139,N_7356);
nor U8307 (N_8307,N_7470,N_7772);
nor U8308 (N_8308,N_7535,N_7151);
nand U8309 (N_8309,N_7417,N_7469);
nand U8310 (N_8310,N_7845,N_7237);
nor U8311 (N_8311,N_7059,N_7314);
or U8312 (N_8312,N_7635,N_7864);
nand U8313 (N_8313,N_7419,N_7387);
nand U8314 (N_8314,N_7928,N_7491);
nand U8315 (N_8315,N_7143,N_7135);
or U8316 (N_8316,N_7252,N_7610);
nor U8317 (N_8317,N_7418,N_7878);
nand U8318 (N_8318,N_7729,N_7076);
and U8319 (N_8319,N_7196,N_7617);
nor U8320 (N_8320,N_7825,N_7344);
or U8321 (N_8321,N_7476,N_7624);
or U8322 (N_8322,N_7266,N_7750);
or U8323 (N_8323,N_7555,N_7828);
and U8324 (N_8324,N_7516,N_7873);
nand U8325 (N_8325,N_7331,N_7755);
nand U8326 (N_8326,N_7968,N_7720);
nor U8327 (N_8327,N_7136,N_7999);
or U8328 (N_8328,N_7348,N_7440);
and U8329 (N_8329,N_7302,N_7649);
and U8330 (N_8330,N_7533,N_7140);
nor U8331 (N_8331,N_7911,N_7374);
and U8332 (N_8332,N_7580,N_7410);
or U8333 (N_8333,N_7452,N_7739);
or U8334 (N_8334,N_7573,N_7872);
or U8335 (N_8335,N_7559,N_7871);
nand U8336 (N_8336,N_7978,N_7383);
nor U8337 (N_8337,N_7965,N_7691);
nor U8338 (N_8338,N_7281,N_7918);
and U8339 (N_8339,N_7291,N_7922);
or U8340 (N_8340,N_7454,N_7296);
nor U8341 (N_8341,N_7686,N_7726);
nand U8342 (N_8342,N_7798,N_7688);
and U8343 (N_8343,N_7818,N_7703);
or U8344 (N_8344,N_7081,N_7125);
and U8345 (N_8345,N_7730,N_7714);
and U8346 (N_8346,N_7586,N_7597);
xor U8347 (N_8347,N_7024,N_7684);
nor U8348 (N_8348,N_7778,N_7627);
or U8349 (N_8349,N_7629,N_7359);
nor U8350 (N_8350,N_7548,N_7044);
or U8351 (N_8351,N_7833,N_7813);
nor U8352 (N_8352,N_7064,N_7576);
or U8353 (N_8353,N_7887,N_7305);
nor U8354 (N_8354,N_7844,N_7900);
or U8355 (N_8355,N_7109,N_7482);
nor U8356 (N_8356,N_7239,N_7165);
and U8357 (N_8357,N_7647,N_7035);
nor U8358 (N_8358,N_7527,N_7702);
or U8359 (N_8359,N_7959,N_7217);
nand U8360 (N_8360,N_7722,N_7388);
or U8361 (N_8361,N_7832,N_7787);
and U8362 (N_8362,N_7015,N_7718);
and U8363 (N_8363,N_7935,N_7467);
nand U8364 (N_8364,N_7486,N_7665);
nand U8365 (N_8365,N_7079,N_7737);
nand U8366 (N_8366,N_7865,N_7479);
nand U8367 (N_8367,N_7651,N_7942);
or U8368 (N_8368,N_7400,N_7485);
and U8369 (N_8369,N_7377,N_7343);
or U8370 (N_8370,N_7695,N_7103);
nand U8371 (N_8371,N_7961,N_7229);
nor U8372 (N_8372,N_7077,N_7711);
and U8373 (N_8373,N_7644,N_7129);
and U8374 (N_8374,N_7710,N_7526);
nand U8375 (N_8375,N_7208,N_7283);
nor U8376 (N_8376,N_7997,N_7317);
or U8377 (N_8377,N_7603,N_7915);
or U8378 (N_8378,N_7543,N_7256);
nand U8379 (N_8379,N_7197,N_7290);
nand U8380 (N_8380,N_7646,N_7771);
nor U8381 (N_8381,N_7456,N_7498);
and U8382 (N_8382,N_7250,N_7542);
and U8383 (N_8383,N_7967,N_7693);
nand U8384 (N_8384,N_7683,N_7541);
nand U8385 (N_8385,N_7204,N_7770);
nand U8386 (N_8386,N_7455,N_7846);
nor U8387 (N_8387,N_7671,N_7327);
or U8388 (N_8388,N_7979,N_7779);
or U8389 (N_8389,N_7230,N_7554);
nor U8390 (N_8390,N_7415,N_7860);
nor U8391 (N_8391,N_7451,N_7842);
nand U8392 (N_8392,N_7449,N_7767);
nand U8393 (N_8393,N_7175,N_7468);
nor U8394 (N_8394,N_7848,N_7150);
and U8395 (N_8395,N_7379,N_7432);
nand U8396 (N_8396,N_7995,N_7461);
nor U8397 (N_8397,N_7956,N_7021);
nand U8398 (N_8398,N_7414,N_7698);
and U8399 (N_8399,N_7650,N_7520);
or U8400 (N_8400,N_7177,N_7953);
or U8401 (N_8401,N_7689,N_7257);
and U8402 (N_8402,N_7231,N_7944);
or U8403 (N_8403,N_7211,N_7537);
and U8404 (N_8404,N_7168,N_7931);
and U8405 (N_8405,N_7780,N_7839);
nand U8406 (N_8406,N_7244,N_7212);
nor U8407 (N_8407,N_7836,N_7444);
nand U8408 (N_8408,N_7147,N_7364);
nor U8409 (N_8409,N_7850,N_7745);
and U8410 (N_8410,N_7796,N_7285);
and U8411 (N_8411,N_7047,N_7068);
nand U8412 (N_8412,N_7152,N_7595);
and U8413 (N_8413,N_7113,N_7719);
and U8414 (N_8414,N_7593,N_7307);
and U8415 (N_8415,N_7776,N_7725);
and U8416 (N_8416,N_7622,N_7020);
or U8417 (N_8417,N_7806,N_7102);
xor U8418 (N_8418,N_7188,N_7280);
nor U8419 (N_8419,N_7194,N_7004);
nand U8420 (N_8420,N_7411,N_7883);
and U8421 (N_8421,N_7275,N_7496);
and U8422 (N_8422,N_7602,N_7039);
and U8423 (N_8423,N_7282,N_7193);
or U8424 (N_8424,N_7513,N_7046);
nor U8425 (N_8425,N_7634,N_7160);
nor U8426 (N_8426,N_7525,N_7349);
xor U8427 (N_8427,N_7232,N_7680);
nand U8428 (N_8428,N_7089,N_7042);
nor U8429 (N_8429,N_7380,N_7265);
nor U8430 (N_8430,N_7128,N_7585);
nand U8431 (N_8431,N_7225,N_7866);
and U8432 (N_8432,N_7333,N_7390);
nand U8433 (N_8433,N_7966,N_7678);
nor U8434 (N_8434,N_7271,N_7332);
or U8435 (N_8435,N_7723,N_7661);
nor U8436 (N_8436,N_7590,N_7434);
or U8437 (N_8437,N_7146,N_7630);
or U8438 (N_8438,N_7596,N_7487);
nand U8439 (N_8439,N_7974,N_7234);
or U8440 (N_8440,N_7473,N_7600);
nor U8441 (N_8441,N_7201,N_7882);
or U8442 (N_8442,N_7805,N_7579);
nor U8443 (N_8443,N_7425,N_7032);
nor U8444 (N_8444,N_7092,N_7062);
nor U8445 (N_8445,N_7203,N_7659);
nor U8446 (N_8446,N_7421,N_7716);
and U8447 (N_8447,N_7494,N_7299);
nor U8448 (N_8448,N_7611,N_7012);
nor U8449 (N_8449,N_7207,N_7027);
nor U8450 (N_8450,N_7993,N_7120);
or U8451 (N_8451,N_7326,N_7761);
nor U8452 (N_8452,N_7057,N_7894);
or U8453 (N_8453,N_7055,N_7657);
nor U8454 (N_8454,N_7591,N_7058);
nor U8455 (N_8455,N_7589,N_7063);
or U8456 (N_8456,N_7263,N_7082);
nand U8457 (N_8457,N_7172,N_7728);
nor U8458 (N_8458,N_7144,N_7186);
nor U8459 (N_8459,N_7949,N_7397);
nor U8460 (N_8460,N_7758,N_7052);
or U8461 (N_8461,N_7809,N_7325);
nor U8462 (N_8462,N_7067,N_7618);
or U8463 (N_8463,N_7925,N_7616);
nor U8464 (N_8464,N_7259,N_7859);
or U8465 (N_8465,N_7508,N_7372);
or U8466 (N_8466,N_7345,N_7205);
and U8467 (N_8467,N_7985,N_7323);
and U8468 (N_8468,N_7394,N_7071);
xor U8469 (N_8469,N_7574,N_7185);
or U8470 (N_8470,N_7926,N_7782);
nor U8471 (N_8471,N_7163,N_7701);
nor U8472 (N_8472,N_7336,N_7464);
nor U8473 (N_8473,N_7233,N_7561);
or U8474 (N_8474,N_7784,N_7988);
or U8475 (N_8475,N_7121,N_7049);
and U8476 (N_8476,N_7258,N_7744);
and U8477 (N_8477,N_7153,N_7821);
or U8478 (N_8478,N_7690,N_7955);
nor U8479 (N_8479,N_7687,N_7037);
nand U8480 (N_8480,N_7360,N_7112);
and U8481 (N_8481,N_7910,N_7328);
and U8482 (N_8482,N_7159,N_7598);
nand U8483 (N_8483,N_7712,N_7704);
and U8484 (N_8484,N_7765,N_7137);
nor U8485 (N_8485,N_7292,N_7075);
nor U8486 (N_8486,N_7731,N_7099);
or U8487 (N_8487,N_7631,N_7270);
nor U8488 (N_8488,N_7253,N_7506);
nor U8489 (N_8489,N_7625,N_7615);
or U8490 (N_8490,N_7189,N_7560);
nand U8491 (N_8491,N_7908,N_7287);
and U8492 (N_8492,N_7975,N_7097);
and U8493 (N_8493,N_7154,N_7810);
and U8494 (N_8494,N_7564,N_7700);
or U8495 (N_8495,N_7540,N_7088);
nor U8496 (N_8496,N_7749,N_7982);
or U8497 (N_8497,N_7158,N_7913);
nand U8498 (N_8498,N_7677,N_7430);
nand U8499 (N_8499,N_7034,N_7734);
nand U8500 (N_8500,N_7950,N_7844);
and U8501 (N_8501,N_7845,N_7023);
nand U8502 (N_8502,N_7018,N_7614);
nor U8503 (N_8503,N_7889,N_7633);
nand U8504 (N_8504,N_7300,N_7488);
and U8505 (N_8505,N_7513,N_7550);
or U8506 (N_8506,N_7604,N_7147);
nor U8507 (N_8507,N_7701,N_7273);
nor U8508 (N_8508,N_7960,N_7105);
and U8509 (N_8509,N_7508,N_7462);
or U8510 (N_8510,N_7619,N_7693);
nand U8511 (N_8511,N_7211,N_7913);
and U8512 (N_8512,N_7167,N_7418);
nor U8513 (N_8513,N_7105,N_7154);
and U8514 (N_8514,N_7749,N_7232);
nor U8515 (N_8515,N_7548,N_7769);
and U8516 (N_8516,N_7744,N_7824);
and U8517 (N_8517,N_7418,N_7208);
or U8518 (N_8518,N_7405,N_7630);
nor U8519 (N_8519,N_7445,N_7870);
or U8520 (N_8520,N_7023,N_7467);
xnor U8521 (N_8521,N_7290,N_7075);
and U8522 (N_8522,N_7698,N_7672);
nor U8523 (N_8523,N_7448,N_7659);
nor U8524 (N_8524,N_7452,N_7974);
nand U8525 (N_8525,N_7622,N_7408);
and U8526 (N_8526,N_7278,N_7970);
or U8527 (N_8527,N_7073,N_7187);
or U8528 (N_8528,N_7319,N_7282);
nor U8529 (N_8529,N_7297,N_7110);
nor U8530 (N_8530,N_7050,N_7576);
and U8531 (N_8531,N_7158,N_7214);
or U8532 (N_8532,N_7049,N_7707);
nand U8533 (N_8533,N_7333,N_7897);
nor U8534 (N_8534,N_7327,N_7708);
and U8535 (N_8535,N_7799,N_7338);
nor U8536 (N_8536,N_7718,N_7487);
and U8537 (N_8537,N_7381,N_7832);
nor U8538 (N_8538,N_7426,N_7234);
or U8539 (N_8539,N_7494,N_7686);
or U8540 (N_8540,N_7706,N_7916);
nand U8541 (N_8541,N_7080,N_7720);
nor U8542 (N_8542,N_7085,N_7508);
nor U8543 (N_8543,N_7143,N_7965);
nor U8544 (N_8544,N_7136,N_7063);
nand U8545 (N_8545,N_7299,N_7922);
or U8546 (N_8546,N_7999,N_7255);
nand U8547 (N_8547,N_7558,N_7788);
or U8548 (N_8548,N_7732,N_7599);
and U8549 (N_8549,N_7588,N_7887);
nor U8550 (N_8550,N_7747,N_7794);
or U8551 (N_8551,N_7754,N_7149);
nand U8552 (N_8552,N_7056,N_7480);
nand U8553 (N_8553,N_7866,N_7026);
and U8554 (N_8554,N_7231,N_7109);
nand U8555 (N_8555,N_7577,N_7134);
nand U8556 (N_8556,N_7280,N_7622);
nor U8557 (N_8557,N_7574,N_7730);
nand U8558 (N_8558,N_7468,N_7934);
nor U8559 (N_8559,N_7904,N_7834);
nand U8560 (N_8560,N_7457,N_7605);
or U8561 (N_8561,N_7763,N_7553);
nor U8562 (N_8562,N_7016,N_7881);
nand U8563 (N_8563,N_7319,N_7985);
and U8564 (N_8564,N_7413,N_7560);
nand U8565 (N_8565,N_7788,N_7652);
or U8566 (N_8566,N_7319,N_7714);
and U8567 (N_8567,N_7127,N_7416);
nor U8568 (N_8568,N_7741,N_7373);
or U8569 (N_8569,N_7931,N_7389);
and U8570 (N_8570,N_7909,N_7738);
and U8571 (N_8571,N_7127,N_7404);
nand U8572 (N_8572,N_7218,N_7654);
nor U8573 (N_8573,N_7411,N_7069);
or U8574 (N_8574,N_7379,N_7173);
or U8575 (N_8575,N_7968,N_7773);
nand U8576 (N_8576,N_7093,N_7479);
nand U8577 (N_8577,N_7040,N_7767);
or U8578 (N_8578,N_7907,N_7152);
and U8579 (N_8579,N_7496,N_7717);
and U8580 (N_8580,N_7426,N_7774);
or U8581 (N_8581,N_7436,N_7937);
nand U8582 (N_8582,N_7865,N_7793);
and U8583 (N_8583,N_7324,N_7856);
or U8584 (N_8584,N_7136,N_7510);
or U8585 (N_8585,N_7316,N_7639);
nor U8586 (N_8586,N_7632,N_7171);
and U8587 (N_8587,N_7255,N_7517);
and U8588 (N_8588,N_7548,N_7302);
nor U8589 (N_8589,N_7188,N_7128);
nand U8590 (N_8590,N_7068,N_7226);
and U8591 (N_8591,N_7194,N_7512);
nor U8592 (N_8592,N_7764,N_7074);
nor U8593 (N_8593,N_7427,N_7007);
nor U8594 (N_8594,N_7559,N_7421);
and U8595 (N_8595,N_7753,N_7152);
nand U8596 (N_8596,N_7259,N_7926);
nand U8597 (N_8597,N_7362,N_7562);
nand U8598 (N_8598,N_7290,N_7240);
and U8599 (N_8599,N_7289,N_7911);
nand U8600 (N_8600,N_7088,N_7327);
nand U8601 (N_8601,N_7448,N_7407);
nand U8602 (N_8602,N_7600,N_7082);
or U8603 (N_8603,N_7183,N_7966);
nand U8604 (N_8604,N_7317,N_7846);
nand U8605 (N_8605,N_7142,N_7333);
nor U8606 (N_8606,N_7338,N_7421);
or U8607 (N_8607,N_7839,N_7225);
nor U8608 (N_8608,N_7066,N_7986);
nand U8609 (N_8609,N_7440,N_7232);
nand U8610 (N_8610,N_7924,N_7437);
nor U8611 (N_8611,N_7963,N_7919);
nand U8612 (N_8612,N_7465,N_7056);
or U8613 (N_8613,N_7603,N_7998);
nor U8614 (N_8614,N_7865,N_7334);
nor U8615 (N_8615,N_7699,N_7967);
or U8616 (N_8616,N_7617,N_7647);
and U8617 (N_8617,N_7929,N_7203);
or U8618 (N_8618,N_7064,N_7706);
nand U8619 (N_8619,N_7799,N_7747);
or U8620 (N_8620,N_7390,N_7036);
and U8621 (N_8621,N_7906,N_7718);
nor U8622 (N_8622,N_7755,N_7137);
and U8623 (N_8623,N_7956,N_7484);
nor U8624 (N_8624,N_7590,N_7881);
or U8625 (N_8625,N_7690,N_7845);
or U8626 (N_8626,N_7800,N_7034);
or U8627 (N_8627,N_7237,N_7517);
nand U8628 (N_8628,N_7137,N_7564);
and U8629 (N_8629,N_7686,N_7522);
nor U8630 (N_8630,N_7191,N_7830);
nand U8631 (N_8631,N_7536,N_7616);
or U8632 (N_8632,N_7690,N_7200);
nor U8633 (N_8633,N_7498,N_7122);
nor U8634 (N_8634,N_7357,N_7119);
nand U8635 (N_8635,N_7213,N_7429);
or U8636 (N_8636,N_7827,N_7167);
and U8637 (N_8637,N_7653,N_7011);
nor U8638 (N_8638,N_7485,N_7508);
nand U8639 (N_8639,N_7619,N_7360);
nand U8640 (N_8640,N_7408,N_7437);
and U8641 (N_8641,N_7790,N_7148);
or U8642 (N_8642,N_7965,N_7174);
nor U8643 (N_8643,N_7003,N_7708);
and U8644 (N_8644,N_7863,N_7827);
and U8645 (N_8645,N_7668,N_7191);
nor U8646 (N_8646,N_7198,N_7235);
nand U8647 (N_8647,N_7800,N_7403);
or U8648 (N_8648,N_7009,N_7087);
or U8649 (N_8649,N_7580,N_7090);
or U8650 (N_8650,N_7060,N_7445);
or U8651 (N_8651,N_7190,N_7593);
and U8652 (N_8652,N_7328,N_7010);
or U8653 (N_8653,N_7049,N_7069);
nor U8654 (N_8654,N_7440,N_7222);
nor U8655 (N_8655,N_7438,N_7986);
or U8656 (N_8656,N_7558,N_7931);
and U8657 (N_8657,N_7629,N_7623);
nand U8658 (N_8658,N_7213,N_7855);
and U8659 (N_8659,N_7821,N_7887);
and U8660 (N_8660,N_7027,N_7642);
or U8661 (N_8661,N_7229,N_7447);
nand U8662 (N_8662,N_7448,N_7160);
nand U8663 (N_8663,N_7483,N_7877);
nor U8664 (N_8664,N_7251,N_7085);
or U8665 (N_8665,N_7560,N_7492);
nand U8666 (N_8666,N_7495,N_7289);
nor U8667 (N_8667,N_7659,N_7757);
and U8668 (N_8668,N_7861,N_7352);
and U8669 (N_8669,N_7062,N_7600);
and U8670 (N_8670,N_7378,N_7960);
nor U8671 (N_8671,N_7140,N_7482);
or U8672 (N_8672,N_7316,N_7808);
nor U8673 (N_8673,N_7827,N_7285);
nand U8674 (N_8674,N_7466,N_7242);
and U8675 (N_8675,N_7130,N_7477);
and U8676 (N_8676,N_7781,N_7583);
and U8677 (N_8677,N_7646,N_7360);
nor U8678 (N_8678,N_7817,N_7300);
nand U8679 (N_8679,N_7180,N_7610);
or U8680 (N_8680,N_7735,N_7341);
or U8681 (N_8681,N_7535,N_7145);
or U8682 (N_8682,N_7501,N_7623);
nor U8683 (N_8683,N_7355,N_7784);
nor U8684 (N_8684,N_7413,N_7337);
nand U8685 (N_8685,N_7857,N_7882);
nor U8686 (N_8686,N_7628,N_7302);
nor U8687 (N_8687,N_7984,N_7953);
nand U8688 (N_8688,N_7876,N_7497);
nand U8689 (N_8689,N_7417,N_7813);
nand U8690 (N_8690,N_7202,N_7682);
nand U8691 (N_8691,N_7446,N_7173);
and U8692 (N_8692,N_7059,N_7813);
or U8693 (N_8693,N_7932,N_7098);
and U8694 (N_8694,N_7363,N_7086);
and U8695 (N_8695,N_7709,N_7941);
or U8696 (N_8696,N_7492,N_7215);
or U8697 (N_8697,N_7395,N_7550);
nand U8698 (N_8698,N_7723,N_7785);
nand U8699 (N_8699,N_7629,N_7342);
and U8700 (N_8700,N_7867,N_7789);
or U8701 (N_8701,N_7115,N_7301);
or U8702 (N_8702,N_7275,N_7648);
or U8703 (N_8703,N_7671,N_7244);
xor U8704 (N_8704,N_7306,N_7702);
or U8705 (N_8705,N_7245,N_7163);
and U8706 (N_8706,N_7806,N_7566);
and U8707 (N_8707,N_7308,N_7018);
nor U8708 (N_8708,N_7834,N_7082);
nand U8709 (N_8709,N_7953,N_7906);
nand U8710 (N_8710,N_7037,N_7326);
xor U8711 (N_8711,N_7863,N_7497);
or U8712 (N_8712,N_7475,N_7134);
or U8713 (N_8713,N_7926,N_7214);
and U8714 (N_8714,N_7052,N_7624);
and U8715 (N_8715,N_7489,N_7844);
nand U8716 (N_8716,N_7410,N_7612);
nor U8717 (N_8717,N_7573,N_7440);
or U8718 (N_8718,N_7548,N_7599);
nand U8719 (N_8719,N_7775,N_7327);
nand U8720 (N_8720,N_7970,N_7043);
nand U8721 (N_8721,N_7698,N_7909);
nand U8722 (N_8722,N_7553,N_7251);
nand U8723 (N_8723,N_7224,N_7753);
and U8724 (N_8724,N_7651,N_7410);
nand U8725 (N_8725,N_7578,N_7816);
nand U8726 (N_8726,N_7335,N_7410);
nor U8727 (N_8727,N_7516,N_7021);
nor U8728 (N_8728,N_7253,N_7569);
nand U8729 (N_8729,N_7954,N_7192);
nand U8730 (N_8730,N_7613,N_7810);
and U8731 (N_8731,N_7280,N_7015);
or U8732 (N_8732,N_7941,N_7701);
nand U8733 (N_8733,N_7938,N_7727);
nor U8734 (N_8734,N_7301,N_7367);
nand U8735 (N_8735,N_7865,N_7131);
or U8736 (N_8736,N_7980,N_7707);
or U8737 (N_8737,N_7797,N_7775);
and U8738 (N_8738,N_7848,N_7505);
nor U8739 (N_8739,N_7871,N_7214);
nor U8740 (N_8740,N_7682,N_7976);
and U8741 (N_8741,N_7712,N_7967);
nand U8742 (N_8742,N_7022,N_7672);
nand U8743 (N_8743,N_7123,N_7048);
nand U8744 (N_8744,N_7347,N_7018);
nand U8745 (N_8745,N_7739,N_7463);
nor U8746 (N_8746,N_7862,N_7494);
and U8747 (N_8747,N_7224,N_7930);
or U8748 (N_8748,N_7369,N_7484);
nor U8749 (N_8749,N_7319,N_7944);
nor U8750 (N_8750,N_7420,N_7526);
xor U8751 (N_8751,N_7162,N_7174);
or U8752 (N_8752,N_7075,N_7253);
or U8753 (N_8753,N_7339,N_7587);
or U8754 (N_8754,N_7895,N_7926);
nand U8755 (N_8755,N_7477,N_7911);
and U8756 (N_8756,N_7043,N_7727);
and U8757 (N_8757,N_7740,N_7552);
nor U8758 (N_8758,N_7634,N_7951);
and U8759 (N_8759,N_7998,N_7085);
and U8760 (N_8760,N_7799,N_7762);
and U8761 (N_8761,N_7351,N_7192);
and U8762 (N_8762,N_7679,N_7661);
nand U8763 (N_8763,N_7549,N_7164);
nor U8764 (N_8764,N_7731,N_7656);
nand U8765 (N_8765,N_7709,N_7745);
or U8766 (N_8766,N_7479,N_7918);
nor U8767 (N_8767,N_7022,N_7497);
nand U8768 (N_8768,N_7199,N_7060);
and U8769 (N_8769,N_7253,N_7454);
nor U8770 (N_8770,N_7712,N_7604);
or U8771 (N_8771,N_7393,N_7659);
nand U8772 (N_8772,N_7951,N_7169);
and U8773 (N_8773,N_7439,N_7006);
nor U8774 (N_8774,N_7519,N_7103);
and U8775 (N_8775,N_7033,N_7899);
nand U8776 (N_8776,N_7264,N_7111);
or U8777 (N_8777,N_7423,N_7565);
and U8778 (N_8778,N_7649,N_7089);
and U8779 (N_8779,N_7995,N_7777);
or U8780 (N_8780,N_7130,N_7354);
nor U8781 (N_8781,N_7866,N_7270);
nor U8782 (N_8782,N_7466,N_7568);
nand U8783 (N_8783,N_7882,N_7358);
nand U8784 (N_8784,N_7047,N_7179);
or U8785 (N_8785,N_7540,N_7765);
or U8786 (N_8786,N_7602,N_7674);
nor U8787 (N_8787,N_7681,N_7791);
and U8788 (N_8788,N_7572,N_7857);
nand U8789 (N_8789,N_7208,N_7596);
nand U8790 (N_8790,N_7196,N_7378);
nand U8791 (N_8791,N_7422,N_7164);
or U8792 (N_8792,N_7096,N_7242);
or U8793 (N_8793,N_7661,N_7607);
nand U8794 (N_8794,N_7758,N_7348);
or U8795 (N_8795,N_7776,N_7215);
nand U8796 (N_8796,N_7109,N_7153);
and U8797 (N_8797,N_7790,N_7192);
and U8798 (N_8798,N_7036,N_7394);
or U8799 (N_8799,N_7703,N_7312);
and U8800 (N_8800,N_7793,N_7348);
or U8801 (N_8801,N_7874,N_7968);
or U8802 (N_8802,N_7179,N_7881);
or U8803 (N_8803,N_7113,N_7581);
nand U8804 (N_8804,N_7996,N_7462);
or U8805 (N_8805,N_7167,N_7931);
or U8806 (N_8806,N_7948,N_7321);
nand U8807 (N_8807,N_7422,N_7428);
nor U8808 (N_8808,N_7822,N_7367);
or U8809 (N_8809,N_7033,N_7602);
and U8810 (N_8810,N_7228,N_7769);
xor U8811 (N_8811,N_7824,N_7798);
and U8812 (N_8812,N_7456,N_7774);
and U8813 (N_8813,N_7254,N_7205);
and U8814 (N_8814,N_7719,N_7790);
nand U8815 (N_8815,N_7104,N_7288);
or U8816 (N_8816,N_7914,N_7333);
nand U8817 (N_8817,N_7445,N_7823);
or U8818 (N_8818,N_7679,N_7550);
or U8819 (N_8819,N_7486,N_7277);
and U8820 (N_8820,N_7634,N_7729);
or U8821 (N_8821,N_7295,N_7943);
nand U8822 (N_8822,N_7403,N_7259);
and U8823 (N_8823,N_7001,N_7061);
or U8824 (N_8824,N_7220,N_7668);
or U8825 (N_8825,N_7085,N_7279);
or U8826 (N_8826,N_7974,N_7834);
and U8827 (N_8827,N_7924,N_7224);
nor U8828 (N_8828,N_7763,N_7376);
nand U8829 (N_8829,N_7858,N_7685);
nor U8830 (N_8830,N_7182,N_7473);
and U8831 (N_8831,N_7527,N_7056);
and U8832 (N_8832,N_7703,N_7773);
nand U8833 (N_8833,N_7251,N_7828);
nand U8834 (N_8834,N_7153,N_7404);
nand U8835 (N_8835,N_7162,N_7289);
and U8836 (N_8836,N_7018,N_7649);
nand U8837 (N_8837,N_7898,N_7818);
nor U8838 (N_8838,N_7783,N_7798);
nand U8839 (N_8839,N_7561,N_7907);
and U8840 (N_8840,N_7085,N_7486);
and U8841 (N_8841,N_7854,N_7445);
nand U8842 (N_8842,N_7150,N_7610);
and U8843 (N_8843,N_7087,N_7159);
and U8844 (N_8844,N_7194,N_7369);
nor U8845 (N_8845,N_7734,N_7478);
and U8846 (N_8846,N_7675,N_7678);
nor U8847 (N_8847,N_7594,N_7905);
or U8848 (N_8848,N_7401,N_7405);
or U8849 (N_8849,N_7918,N_7038);
or U8850 (N_8850,N_7458,N_7183);
nor U8851 (N_8851,N_7435,N_7326);
nor U8852 (N_8852,N_7591,N_7138);
or U8853 (N_8853,N_7577,N_7548);
and U8854 (N_8854,N_7881,N_7627);
or U8855 (N_8855,N_7563,N_7353);
or U8856 (N_8856,N_7305,N_7464);
nand U8857 (N_8857,N_7581,N_7508);
or U8858 (N_8858,N_7911,N_7265);
nor U8859 (N_8859,N_7754,N_7860);
nor U8860 (N_8860,N_7536,N_7407);
or U8861 (N_8861,N_7822,N_7957);
and U8862 (N_8862,N_7111,N_7741);
nand U8863 (N_8863,N_7720,N_7168);
and U8864 (N_8864,N_7789,N_7233);
nand U8865 (N_8865,N_7628,N_7346);
nand U8866 (N_8866,N_7453,N_7461);
nor U8867 (N_8867,N_7516,N_7117);
nand U8868 (N_8868,N_7927,N_7496);
nor U8869 (N_8869,N_7969,N_7660);
and U8870 (N_8870,N_7001,N_7538);
and U8871 (N_8871,N_7779,N_7752);
and U8872 (N_8872,N_7416,N_7059);
nand U8873 (N_8873,N_7911,N_7000);
nand U8874 (N_8874,N_7873,N_7272);
and U8875 (N_8875,N_7229,N_7993);
and U8876 (N_8876,N_7310,N_7971);
nand U8877 (N_8877,N_7428,N_7806);
nand U8878 (N_8878,N_7915,N_7768);
nor U8879 (N_8879,N_7684,N_7142);
nand U8880 (N_8880,N_7237,N_7838);
and U8881 (N_8881,N_7587,N_7245);
nand U8882 (N_8882,N_7861,N_7446);
or U8883 (N_8883,N_7361,N_7906);
nand U8884 (N_8884,N_7816,N_7233);
or U8885 (N_8885,N_7519,N_7178);
nor U8886 (N_8886,N_7401,N_7781);
and U8887 (N_8887,N_7463,N_7257);
nor U8888 (N_8888,N_7016,N_7250);
nand U8889 (N_8889,N_7502,N_7123);
or U8890 (N_8890,N_7577,N_7041);
nor U8891 (N_8891,N_7552,N_7192);
and U8892 (N_8892,N_7420,N_7933);
nand U8893 (N_8893,N_7395,N_7425);
or U8894 (N_8894,N_7615,N_7152);
and U8895 (N_8895,N_7117,N_7881);
or U8896 (N_8896,N_7649,N_7189);
nand U8897 (N_8897,N_7868,N_7387);
or U8898 (N_8898,N_7039,N_7283);
nand U8899 (N_8899,N_7959,N_7285);
nand U8900 (N_8900,N_7135,N_7630);
nor U8901 (N_8901,N_7203,N_7285);
and U8902 (N_8902,N_7524,N_7518);
or U8903 (N_8903,N_7004,N_7035);
nand U8904 (N_8904,N_7160,N_7979);
nand U8905 (N_8905,N_7905,N_7620);
xor U8906 (N_8906,N_7071,N_7778);
or U8907 (N_8907,N_7873,N_7367);
or U8908 (N_8908,N_7935,N_7886);
and U8909 (N_8909,N_7872,N_7501);
and U8910 (N_8910,N_7817,N_7607);
nor U8911 (N_8911,N_7284,N_7201);
nand U8912 (N_8912,N_7548,N_7357);
and U8913 (N_8913,N_7572,N_7766);
nor U8914 (N_8914,N_7299,N_7778);
nand U8915 (N_8915,N_7591,N_7319);
and U8916 (N_8916,N_7449,N_7845);
nor U8917 (N_8917,N_7897,N_7405);
nand U8918 (N_8918,N_7630,N_7941);
and U8919 (N_8919,N_7237,N_7320);
and U8920 (N_8920,N_7750,N_7913);
or U8921 (N_8921,N_7852,N_7258);
or U8922 (N_8922,N_7108,N_7993);
or U8923 (N_8923,N_7423,N_7080);
nor U8924 (N_8924,N_7960,N_7585);
or U8925 (N_8925,N_7624,N_7111);
nand U8926 (N_8926,N_7925,N_7201);
and U8927 (N_8927,N_7290,N_7385);
nor U8928 (N_8928,N_7436,N_7395);
nand U8929 (N_8929,N_7496,N_7077);
nor U8930 (N_8930,N_7774,N_7116);
nand U8931 (N_8931,N_7620,N_7391);
or U8932 (N_8932,N_7286,N_7213);
nor U8933 (N_8933,N_7436,N_7912);
or U8934 (N_8934,N_7694,N_7366);
nor U8935 (N_8935,N_7641,N_7823);
and U8936 (N_8936,N_7756,N_7477);
and U8937 (N_8937,N_7678,N_7157);
or U8938 (N_8938,N_7069,N_7867);
or U8939 (N_8939,N_7824,N_7426);
and U8940 (N_8940,N_7913,N_7381);
or U8941 (N_8941,N_7787,N_7469);
nand U8942 (N_8942,N_7321,N_7594);
or U8943 (N_8943,N_7376,N_7981);
nand U8944 (N_8944,N_7863,N_7201);
or U8945 (N_8945,N_7021,N_7165);
nand U8946 (N_8946,N_7629,N_7554);
and U8947 (N_8947,N_7933,N_7516);
or U8948 (N_8948,N_7197,N_7422);
and U8949 (N_8949,N_7749,N_7178);
or U8950 (N_8950,N_7240,N_7886);
and U8951 (N_8951,N_7701,N_7614);
and U8952 (N_8952,N_7309,N_7902);
and U8953 (N_8953,N_7578,N_7534);
nor U8954 (N_8954,N_7041,N_7260);
nand U8955 (N_8955,N_7605,N_7351);
and U8956 (N_8956,N_7377,N_7157);
and U8957 (N_8957,N_7719,N_7923);
or U8958 (N_8958,N_7093,N_7349);
nand U8959 (N_8959,N_7773,N_7803);
and U8960 (N_8960,N_7794,N_7965);
or U8961 (N_8961,N_7549,N_7234);
nand U8962 (N_8962,N_7404,N_7867);
and U8963 (N_8963,N_7082,N_7871);
xor U8964 (N_8964,N_7518,N_7814);
nor U8965 (N_8965,N_7133,N_7935);
nor U8966 (N_8966,N_7028,N_7246);
nor U8967 (N_8967,N_7044,N_7639);
nand U8968 (N_8968,N_7721,N_7120);
and U8969 (N_8969,N_7041,N_7918);
nand U8970 (N_8970,N_7096,N_7763);
nand U8971 (N_8971,N_7028,N_7560);
or U8972 (N_8972,N_7436,N_7346);
nand U8973 (N_8973,N_7351,N_7380);
or U8974 (N_8974,N_7614,N_7534);
nand U8975 (N_8975,N_7413,N_7442);
nor U8976 (N_8976,N_7312,N_7314);
or U8977 (N_8977,N_7291,N_7306);
and U8978 (N_8978,N_7035,N_7713);
nor U8979 (N_8979,N_7618,N_7641);
nand U8980 (N_8980,N_7323,N_7492);
and U8981 (N_8981,N_7230,N_7396);
or U8982 (N_8982,N_7402,N_7562);
nor U8983 (N_8983,N_7423,N_7737);
and U8984 (N_8984,N_7201,N_7469);
or U8985 (N_8985,N_7584,N_7380);
nand U8986 (N_8986,N_7352,N_7081);
or U8987 (N_8987,N_7114,N_7583);
and U8988 (N_8988,N_7606,N_7032);
or U8989 (N_8989,N_7930,N_7602);
and U8990 (N_8990,N_7487,N_7355);
and U8991 (N_8991,N_7269,N_7716);
nand U8992 (N_8992,N_7309,N_7149);
or U8993 (N_8993,N_7913,N_7879);
or U8994 (N_8994,N_7579,N_7743);
nand U8995 (N_8995,N_7914,N_7387);
nand U8996 (N_8996,N_7401,N_7289);
or U8997 (N_8997,N_7491,N_7297);
and U8998 (N_8998,N_7479,N_7703);
or U8999 (N_8999,N_7024,N_7942);
nand U9000 (N_9000,N_8969,N_8424);
and U9001 (N_9001,N_8551,N_8224);
and U9002 (N_9002,N_8060,N_8243);
or U9003 (N_9003,N_8235,N_8766);
nor U9004 (N_9004,N_8359,N_8640);
nor U9005 (N_9005,N_8286,N_8271);
or U9006 (N_9006,N_8309,N_8694);
nand U9007 (N_9007,N_8530,N_8390);
nand U9008 (N_9008,N_8531,N_8478);
nor U9009 (N_9009,N_8036,N_8542);
and U9010 (N_9010,N_8804,N_8084);
nand U9011 (N_9011,N_8067,N_8693);
and U9012 (N_9012,N_8041,N_8737);
nor U9013 (N_9013,N_8805,N_8559);
and U9014 (N_9014,N_8610,N_8690);
nand U9015 (N_9015,N_8656,N_8715);
xor U9016 (N_9016,N_8139,N_8381);
nor U9017 (N_9017,N_8046,N_8516);
or U9018 (N_9018,N_8782,N_8460);
or U9019 (N_9019,N_8176,N_8898);
nand U9020 (N_9020,N_8903,N_8502);
or U9021 (N_9021,N_8170,N_8221);
nor U9022 (N_9022,N_8863,N_8131);
or U9023 (N_9023,N_8042,N_8930);
or U9024 (N_9024,N_8733,N_8957);
nand U9025 (N_9025,N_8261,N_8312);
and U9026 (N_9026,N_8966,N_8540);
nor U9027 (N_9027,N_8707,N_8403);
and U9028 (N_9028,N_8661,N_8807);
nand U9029 (N_9029,N_8239,N_8480);
or U9030 (N_9030,N_8518,N_8498);
nor U9031 (N_9031,N_8052,N_8616);
nand U9032 (N_9032,N_8878,N_8982);
or U9033 (N_9033,N_8816,N_8301);
or U9034 (N_9034,N_8653,N_8713);
nor U9035 (N_9035,N_8488,N_8014);
nor U9036 (N_9036,N_8647,N_8706);
and U9037 (N_9037,N_8682,N_8337);
nor U9038 (N_9038,N_8035,N_8007);
or U9039 (N_9039,N_8907,N_8228);
and U9040 (N_9040,N_8742,N_8254);
nor U9041 (N_9041,N_8075,N_8011);
nor U9042 (N_9042,N_8560,N_8673);
nand U9043 (N_9043,N_8865,N_8435);
nand U9044 (N_9044,N_8281,N_8943);
nand U9045 (N_9045,N_8140,N_8624);
and U9046 (N_9046,N_8776,N_8008);
nor U9047 (N_9047,N_8797,N_8576);
nor U9048 (N_9048,N_8380,N_8636);
nor U9049 (N_9049,N_8377,N_8853);
and U9050 (N_9050,N_8732,N_8596);
nor U9051 (N_9051,N_8545,N_8701);
nor U9052 (N_9052,N_8563,N_8099);
or U9053 (N_9053,N_8144,N_8473);
or U9054 (N_9054,N_8592,N_8984);
nand U9055 (N_9055,N_8942,N_8843);
and U9056 (N_9056,N_8594,N_8976);
nand U9057 (N_9057,N_8794,N_8323);
and U9058 (N_9058,N_8882,N_8894);
nand U9059 (N_9059,N_8220,N_8638);
and U9060 (N_9060,N_8810,N_8864);
and U9061 (N_9061,N_8858,N_8961);
nand U9062 (N_9062,N_8096,N_8280);
nand U9063 (N_9063,N_8072,N_8040);
nand U9064 (N_9064,N_8983,N_8463);
and U9065 (N_9065,N_8829,N_8155);
and U9066 (N_9066,N_8423,N_8465);
nand U9067 (N_9067,N_8136,N_8289);
nand U9068 (N_9068,N_8141,N_8826);
or U9069 (N_9069,N_8857,N_8253);
nor U9070 (N_9070,N_8368,N_8762);
and U9071 (N_9071,N_8487,N_8991);
nand U9072 (N_9072,N_8953,N_8043);
and U9073 (N_9073,N_8836,N_8106);
or U9074 (N_9074,N_8555,N_8348);
or U9075 (N_9075,N_8058,N_8727);
nand U9076 (N_9076,N_8366,N_8455);
or U9077 (N_9077,N_8407,N_8291);
or U9078 (N_9078,N_8497,N_8845);
and U9079 (N_9079,N_8840,N_8834);
or U9080 (N_9080,N_8595,N_8108);
nand U9081 (N_9081,N_8338,N_8973);
or U9082 (N_9082,N_8102,N_8247);
and U9083 (N_9083,N_8893,N_8955);
or U9084 (N_9084,N_8097,N_8468);
nand U9085 (N_9085,N_8978,N_8436);
or U9086 (N_9086,N_8245,N_8785);
or U9087 (N_9087,N_8669,N_8087);
and U9088 (N_9088,N_8216,N_8318);
and U9089 (N_9089,N_8924,N_8607);
and U9090 (N_9090,N_8900,N_8946);
and U9091 (N_9091,N_8929,N_8507);
nand U9092 (N_9092,N_8584,N_8244);
xnor U9093 (N_9093,N_8406,N_8045);
and U9094 (N_9094,N_8740,N_8928);
and U9095 (N_9095,N_8009,N_8609);
or U9096 (N_9096,N_8920,N_8404);
nor U9097 (N_9097,N_8288,N_8699);
or U9098 (N_9098,N_8529,N_8203);
and U9099 (N_9099,N_8909,N_8501);
nand U9100 (N_9100,N_8362,N_8416);
nor U9101 (N_9101,N_8428,N_8723);
nor U9102 (N_9102,N_8830,N_8241);
nand U9103 (N_9103,N_8586,N_8562);
nor U9104 (N_9104,N_8887,N_8789);
and U9105 (N_9105,N_8971,N_8490);
or U9106 (N_9106,N_8815,N_8996);
nand U9107 (N_9107,N_8225,N_8324);
and U9108 (N_9108,N_8189,N_8968);
or U9109 (N_9109,N_8258,N_8837);
or U9110 (N_9110,N_8462,N_8208);
nand U9111 (N_9111,N_8438,N_8933);
nand U9112 (N_9112,N_8588,N_8371);
nor U9113 (N_9113,N_8457,N_8904);
nor U9114 (N_9114,N_8877,N_8828);
nand U9115 (N_9115,N_8307,N_8617);
nand U9116 (N_9116,N_8772,N_8374);
or U9117 (N_9117,N_8524,N_8979);
and U9118 (N_9118,N_8447,N_8913);
nor U9119 (N_9119,N_8384,N_8070);
nand U9120 (N_9120,N_8160,N_8965);
nand U9121 (N_9121,N_8506,N_8902);
and U9122 (N_9122,N_8652,N_8484);
nor U9123 (N_9123,N_8206,N_8477);
and U9124 (N_9124,N_8875,N_8604);
nand U9125 (N_9125,N_8015,N_8059);
and U9126 (N_9126,N_8411,N_8410);
and U9127 (N_9127,N_8093,N_8730);
and U9128 (N_9128,N_8449,N_8747);
and U9129 (N_9129,N_8284,N_8495);
and U9130 (N_9130,N_8535,N_8358);
or U9131 (N_9131,N_8944,N_8485);
or U9132 (N_9132,N_8593,N_8055);
or U9133 (N_9133,N_8811,N_8728);
or U9134 (N_9134,N_8489,N_8214);
and U9135 (N_9135,N_8899,N_8212);
xnor U9136 (N_9136,N_8739,N_8382);
and U9137 (N_9137,N_8549,N_8166);
nor U9138 (N_9138,N_8252,N_8431);
or U9139 (N_9139,N_8975,N_8251);
nand U9140 (N_9140,N_8743,N_8546);
and U9141 (N_9141,N_8325,N_8023);
nand U9142 (N_9142,N_8672,N_8614);
or U9143 (N_9143,N_8022,N_8082);
nand U9144 (N_9144,N_8685,N_8111);
nor U9145 (N_9145,N_8660,N_8866);
or U9146 (N_9146,N_8020,N_8705);
nand U9147 (N_9147,N_8453,N_8990);
nand U9148 (N_9148,N_8658,N_8057);
nor U9149 (N_9149,N_8736,N_8197);
or U9150 (N_9150,N_8226,N_8885);
or U9151 (N_9151,N_8077,N_8849);
nor U9152 (N_9152,N_8134,N_8038);
or U9153 (N_9153,N_8951,N_8080);
nand U9154 (N_9154,N_8612,N_8575);
or U9155 (N_9155,N_8839,N_8724);
nand U9156 (N_9156,N_8912,N_8405);
nor U9157 (N_9157,N_8151,N_8343);
nand U9158 (N_9158,N_8687,N_8356);
nor U9159 (N_9159,N_8599,N_8491);
nand U9160 (N_9160,N_8964,N_8376);
and U9161 (N_9161,N_8110,N_8388);
and U9162 (N_9162,N_8282,N_8421);
or U9163 (N_9163,N_8475,N_8981);
and U9164 (N_9164,N_8364,N_8700);
and U9165 (N_9165,N_8391,N_8958);
nor U9166 (N_9166,N_8026,N_8886);
or U9167 (N_9167,N_8222,N_8056);
and U9168 (N_9168,N_8665,N_8033);
and U9169 (N_9169,N_8274,N_8856);
and U9170 (N_9170,N_8873,N_8319);
xor U9171 (N_9171,N_8623,N_8167);
nor U9172 (N_9172,N_8444,N_8127);
and U9173 (N_9173,N_8925,N_8795);
and U9174 (N_9174,N_8426,N_8165);
nand U9175 (N_9175,N_8063,N_8149);
or U9176 (N_9176,N_8517,N_8526);
nor U9177 (N_9177,N_8051,N_8544);
or U9178 (N_9178,N_8211,N_8628);
nor U9179 (N_9179,N_8445,N_8750);
or U9180 (N_9180,N_8527,N_8948);
or U9181 (N_9181,N_8392,N_8613);
or U9182 (N_9182,N_8788,N_8105);
nor U9183 (N_9183,N_8980,N_8564);
nand U9184 (N_9184,N_8351,N_8691);
nor U9185 (N_9185,N_8128,N_8717);
and U9186 (N_9186,N_8499,N_8704);
nand U9187 (N_9187,N_8164,N_8369);
or U9188 (N_9188,N_8570,N_8117);
or U9189 (N_9189,N_8771,N_8327);
and U9190 (N_9190,N_8360,N_8010);
nand U9191 (N_9191,N_8365,N_8914);
nand U9192 (N_9192,N_8315,N_8012);
and U9193 (N_9193,N_8270,N_8272);
and U9194 (N_9194,N_8994,N_8352);
nand U9195 (N_9195,N_8896,N_8357);
nand U9196 (N_9196,N_8967,N_8764);
nand U9197 (N_9197,N_8671,N_8071);
nor U9198 (N_9198,N_8825,N_8006);
xnor U9199 (N_9199,N_8910,N_8585);
nor U9200 (N_9200,N_8088,N_8814);
nand U9201 (N_9201,N_8695,N_8722);
and U9202 (N_9202,N_8784,N_8999);
nand U9203 (N_9203,N_8630,N_8657);
nand U9204 (N_9204,N_8154,N_8440);
or U9205 (N_9205,N_8299,N_8977);
and U9206 (N_9206,N_8278,N_8400);
or U9207 (N_9207,N_8279,N_8079);
nor U9208 (N_9208,N_8760,N_8918);
or U9209 (N_9209,N_8321,N_8459);
nand U9210 (N_9210,N_8275,N_8970);
nand U9211 (N_9211,N_8684,N_8726);
nand U9212 (N_9212,N_8582,N_8565);
nor U9213 (N_9213,N_8703,N_8314);
and U9214 (N_9214,N_8567,N_8231);
and U9215 (N_9215,N_8751,N_8842);
or U9216 (N_9216,N_8800,N_8114);
nand U9217 (N_9217,N_8210,N_8787);
and U9218 (N_9218,N_8399,N_8632);
or U9219 (N_9219,N_8068,N_8611);
nand U9220 (N_9220,N_8417,N_8121);
nand U9221 (N_9221,N_8854,N_8135);
and U9222 (N_9222,N_8443,N_8408);
and U9223 (N_9223,N_8791,N_8827);
nor U9224 (N_9224,N_8073,N_8092);
or U9225 (N_9225,N_8494,N_8735);
and U9226 (N_9226,N_8474,N_8193);
and U9227 (N_9227,N_8115,N_8832);
nand U9228 (N_9228,N_8777,N_8960);
nand U9229 (N_9229,N_8393,N_8897);
nor U9230 (N_9230,N_8932,N_8870);
and U9231 (N_9231,N_8763,N_8219);
and U9232 (N_9232,N_8859,N_8074);
or U9233 (N_9233,N_8892,N_8395);
and U9234 (N_9234,N_8086,N_8752);
nor U9235 (N_9235,N_8163,N_8643);
and U9236 (N_9236,N_8525,N_8838);
nor U9237 (N_9237,N_8808,N_8822);
or U9238 (N_9238,N_8332,N_8234);
or U9239 (N_9239,N_8622,N_8770);
and U9240 (N_9240,N_8028,N_8541);
nor U9241 (N_9241,N_8619,N_8126);
nor U9242 (N_9242,N_8744,N_8013);
and U9243 (N_9243,N_8940,N_8341);
nor U9244 (N_9244,N_8150,N_8504);
nor U9245 (N_9245,N_8016,N_8688);
or U9246 (N_9246,N_8831,N_8880);
nand U9247 (N_9247,N_8238,N_8620);
nor U9248 (N_9248,N_8152,N_8945);
or U9249 (N_9249,N_8179,N_8786);
nand U9250 (N_9250,N_8668,N_8230);
and U9251 (N_9251,N_8361,N_8508);
nor U9252 (N_9252,N_8601,N_8353);
or U9253 (N_9253,N_8533,N_8186);
nand U9254 (N_9254,N_8402,N_8302);
nand U9255 (N_9255,N_8861,N_8047);
or U9256 (N_9256,N_8850,N_8846);
nor U9257 (N_9257,N_8452,N_8470);
or U9258 (N_9258,N_8881,N_8566);
nand U9259 (N_9259,N_8681,N_8686);
and U9260 (N_9260,N_8019,N_8989);
nor U9261 (N_9261,N_8265,N_8482);
or U9262 (N_9262,N_8202,N_8579);
or U9263 (N_9263,N_8153,N_8386);
and U9264 (N_9264,N_8574,N_8716);
and U9265 (N_9265,N_8534,N_8833);
and U9266 (N_9266,N_8064,N_8862);
or U9267 (N_9267,N_8118,N_8554);
nand U9268 (N_9268,N_8890,N_8333);
or U9269 (N_9269,N_8646,N_8821);
or U9270 (N_9270,N_8187,N_8448);
nand U9271 (N_9271,N_8532,N_8439);
nor U9272 (N_9272,N_8335,N_8195);
nor U9273 (N_9273,N_8769,N_8293);
or U9274 (N_9274,N_8401,N_8227);
nand U9275 (N_9275,N_8577,N_8956);
or U9276 (N_9276,N_8005,N_8156);
or U9277 (N_9277,N_8626,N_8146);
and U9278 (N_9278,N_8027,N_8874);
or U9279 (N_9279,N_8655,N_8602);
nor U9280 (N_9280,N_8172,N_8169);
nand U9281 (N_9281,N_8848,N_8383);
nor U9282 (N_9282,N_8458,N_8032);
and U9283 (N_9283,N_8679,N_8683);
nand U9284 (N_9284,N_8414,N_8773);
nand U9285 (N_9285,N_8062,N_8483);
xnor U9286 (N_9286,N_8180,N_8412);
or U9287 (N_9287,N_8952,N_8556);
or U9288 (N_9288,N_8519,N_8606);
or U9289 (N_9289,N_8420,N_8528);
and U9290 (N_9290,N_8986,N_8198);
nor U9291 (N_9291,N_8394,N_8915);
or U9292 (N_9292,N_8342,N_8547);
and U9293 (N_9293,N_8631,N_8514);
nand U9294 (N_9294,N_8844,N_8793);
or U9295 (N_9295,N_8992,N_8132);
nor U9296 (N_9296,N_8017,N_8250);
or U9297 (N_9297,N_8138,N_8761);
or U9298 (N_9298,N_8905,N_8583);
or U9299 (N_9299,N_8486,N_8629);
nor U9300 (N_9300,N_8213,N_8756);
and U9301 (N_9301,N_8031,N_8851);
and U9302 (N_9302,N_8988,N_8954);
and U9303 (N_9303,N_8133,N_8003);
and U9304 (N_9304,N_8702,N_8290);
and U9305 (N_9305,N_8917,N_8720);
nor U9306 (N_9306,N_8397,N_8550);
nand U9307 (N_9307,N_8322,N_8446);
or U9308 (N_9308,N_8678,N_8817);
nand U9309 (N_9309,N_8109,N_8300);
nor U9310 (N_9310,N_8171,N_8974);
and U9311 (N_9311,N_8199,N_8911);
nor U9312 (N_9312,N_8137,N_8888);
xor U9313 (N_9313,N_8512,N_8159);
and U9314 (N_9314,N_8568,N_8696);
or U9315 (N_9315,N_8259,N_8835);
or U9316 (N_9316,N_8367,N_8581);
or U9317 (N_9317,N_8513,N_8260);
or U9318 (N_9318,N_8561,N_8758);
and U9319 (N_9319,N_8158,N_8884);
nor U9320 (N_9320,N_8000,N_8759);
and U9321 (N_9321,N_8065,N_8263);
nor U9322 (N_9322,N_8142,N_8266);
nand U9323 (N_9323,N_8240,N_8799);
and U9324 (N_9324,N_8370,N_8441);
or U9325 (N_9325,N_8124,N_8476);
and U9326 (N_9326,N_8451,N_8895);
or U9327 (N_9327,N_8190,N_8675);
or U9328 (N_9328,N_8178,N_8269);
nand U9329 (N_9329,N_8125,N_8605);
and U9330 (N_9330,N_8711,N_8454);
nand U9331 (N_9331,N_8608,N_8995);
nand U9332 (N_9332,N_8340,N_8298);
xnor U9333 (N_9333,N_8801,N_8147);
and U9334 (N_9334,N_8091,N_8303);
nor U9335 (N_9335,N_8157,N_8676);
nand U9336 (N_9336,N_8456,N_8634);
or U9337 (N_9337,N_8698,N_8419);
nand U9338 (N_9338,N_8871,N_8292);
and U9339 (N_9339,N_8089,N_8373);
and U9340 (N_9340,N_8308,N_8783);
nor U9341 (N_9341,N_8387,N_8818);
or U9342 (N_9342,N_8409,N_8824);
or U9343 (N_9343,N_8218,N_8641);
nand U9344 (N_9344,N_8589,N_8191);
nand U9345 (N_9345,N_8328,N_8237);
nand U9346 (N_9346,N_8037,N_8174);
nor U9347 (N_9347,N_8578,N_8347);
nand U9348 (N_9348,N_8637,N_8709);
and U9349 (N_9349,N_8883,N_8201);
or U9350 (N_9350,N_8642,N_8537);
nor U9351 (N_9351,N_8354,N_8719);
nor U9352 (N_9352,N_8908,N_8223);
or U9353 (N_9353,N_8867,N_8746);
nor U9354 (N_9354,N_8796,N_8648);
or U9355 (N_9355,N_8615,N_8923);
or U9356 (N_9356,N_8030,N_8745);
or U9357 (N_9357,N_8813,N_8034);
and U9358 (N_9358,N_8569,N_8442);
or U9359 (N_9359,N_8116,N_8129);
or U9360 (N_9360,N_8069,N_8538);
nand U9361 (N_9361,N_8748,N_8767);
or U9362 (N_9362,N_8083,N_8331);
nor U9363 (N_9363,N_8644,N_8217);
nor U9364 (N_9364,N_8183,N_8820);
nor U9365 (N_9365,N_8204,N_8479);
or U9366 (N_9366,N_8363,N_8078);
nor U9367 (N_9367,N_8916,N_8714);
and U9368 (N_9368,N_8076,N_8779);
or U9369 (N_9369,N_8081,N_8493);
nand U9370 (N_9370,N_8249,N_8667);
nand U9371 (N_9371,N_8339,N_8434);
or U9372 (N_9372,N_8464,N_8103);
and U9373 (N_9373,N_8649,N_8625);
nand U9374 (N_9374,N_8185,N_8768);
or U9375 (N_9375,N_8509,N_8757);
nor U9376 (N_9376,N_8054,N_8855);
or U9377 (N_9377,N_8635,N_8018);
nor U9378 (N_9378,N_8432,N_8385);
nand U9379 (N_9379,N_8122,N_8847);
or U9380 (N_9380,N_8734,N_8329);
nor U9381 (N_9381,N_8295,N_8048);
and U9382 (N_9382,N_8304,N_8044);
nand U9383 (N_9383,N_8334,N_8543);
nand U9384 (N_9384,N_8868,N_8515);
and U9385 (N_9385,N_8674,N_8173);
or U9386 (N_9386,N_8998,N_8264);
and U9387 (N_9387,N_8194,N_8936);
or U9388 (N_9388,N_8860,N_8107);
and U9389 (N_9389,N_8598,N_8100);
or U9390 (N_9390,N_8511,N_8841);
or U9391 (N_9391,N_8389,N_8311);
or U9392 (N_9392,N_8677,N_8350);
or U9393 (N_9393,N_8781,N_8242);
or U9394 (N_9394,N_8085,N_8061);
and U9395 (N_9395,N_8765,N_8774);
nand U9396 (N_9396,N_8066,N_8901);
and U9397 (N_9397,N_8778,N_8294);
nor U9398 (N_9398,N_8651,N_8196);
nor U9399 (N_9399,N_8375,N_8130);
nor U9400 (N_9400,N_8947,N_8466);
nor U9401 (N_9401,N_8320,N_8267);
nor U9402 (N_9402,N_8664,N_8654);
or U9403 (N_9403,N_8277,N_8120);
nand U9404 (N_9404,N_8305,N_8580);
and U9405 (N_9405,N_8257,N_8573);
nor U9406 (N_9406,N_8852,N_8162);
or U9407 (N_9407,N_8963,N_8104);
and U9408 (N_9408,N_8938,N_8729);
nor U9409 (N_9409,N_8557,N_8558);
nor U9410 (N_9410,N_8879,N_8236);
nor U9411 (N_9411,N_8819,N_8520);
nor U9412 (N_9412,N_8712,N_8987);
nand U9413 (N_9413,N_8603,N_8906);
nand U9414 (N_9414,N_8467,N_8572);
or U9415 (N_9415,N_8627,N_8993);
or U9416 (N_9416,N_8024,N_8548);
nand U9417 (N_9417,N_8869,N_8738);
nand U9418 (N_9418,N_8919,N_8510);
and U9419 (N_9419,N_8143,N_8181);
nor U9420 (N_9420,N_8823,N_8168);
or U9421 (N_9421,N_8433,N_8809);
and U9422 (N_9422,N_8553,N_8256);
or U9423 (N_9423,N_8207,N_8429);
or U9424 (N_9424,N_8276,N_8184);
or U9425 (N_9425,N_8378,N_8306);
and U9426 (N_9426,N_8934,N_8316);
nor U9427 (N_9427,N_8001,N_8755);
and U9428 (N_9428,N_8689,N_8413);
and U9429 (N_9429,N_8496,N_8937);
or U9430 (N_9430,N_8792,N_8552);
nor U9431 (N_9431,N_8721,N_8050);
nor U9432 (N_9432,N_8725,N_8317);
and U9433 (N_9433,N_8505,N_8113);
and U9434 (N_9434,N_8002,N_8021);
nor U9435 (N_9435,N_8025,N_8876);
and U9436 (N_9436,N_8273,N_8398);
and U9437 (N_9437,N_8188,N_8330);
and U9438 (N_9438,N_8425,N_8029);
and U9439 (N_9439,N_8663,N_8004);
or U9440 (N_9440,N_8095,N_8539);
nand U9441 (N_9441,N_8396,N_8469);
and U9442 (N_9442,N_8205,N_8255);
or U9443 (N_9443,N_8939,N_8621);
or U9444 (N_9444,N_8492,N_8461);
or U9445 (N_9445,N_8336,N_8680);
or U9446 (N_9446,N_8536,N_8098);
or U9447 (N_9447,N_8039,N_8941);
or U9448 (N_9448,N_8645,N_8430);
nand U9449 (N_9449,N_8692,N_8962);
and U9450 (N_9450,N_8798,N_8522);
or U9451 (N_9451,N_8889,N_8803);
and U9452 (N_9452,N_8659,N_8297);
or U9453 (N_9453,N_8618,N_8285);
nand U9454 (N_9454,N_8215,N_8248);
or U9455 (N_9455,N_8600,N_8345);
nand U9456 (N_9456,N_8422,N_8112);
xnor U9457 (N_9457,N_8521,N_8471);
nor U9458 (N_9458,N_8229,N_8500);
nor U9459 (N_9459,N_8959,N_8283);
nor U9460 (N_9460,N_8472,N_8891);
and U9461 (N_9461,N_8597,N_8935);
nand U9462 (N_9462,N_8145,N_8346);
nor U9463 (N_9463,N_8209,N_8175);
nor U9464 (N_9464,N_8775,N_8326);
or U9465 (N_9465,N_8872,N_8780);
nor U9466 (N_9466,N_8148,N_8931);
and U9467 (N_9467,N_8503,N_8571);
nand U9468 (N_9468,N_8650,N_8741);
nor U9469 (N_9469,N_8262,N_8749);
nand U9470 (N_9470,N_8710,N_8587);
nor U9471 (N_9471,N_8927,N_8481);
nor U9472 (N_9472,N_8662,N_8090);
nor U9473 (N_9473,N_8182,N_8177);
or U9474 (N_9474,N_8697,N_8349);
or U9475 (N_9475,N_8344,N_8094);
and U9476 (N_9476,N_8437,N_8731);
or U9477 (N_9477,N_8718,N_8119);
nor U9478 (N_9478,N_8926,N_8790);
and U9479 (N_9479,N_8450,N_8949);
nor U9480 (N_9480,N_8192,N_8590);
nor U9481 (N_9481,N_8233,N_8427);
nand U9482 (N_9482,N_8922,N_8049);
and U9483 (N_9483,N_8753,N_8287);
and U9484 (N_9484,N_8200,N_8161);
nor U9485 (N_9485,N_8123,N_8523);
or U9486 (N_9486,N_8997,N_8310);
or U9487 (N_9487,N_8950,N_8296);
or U9488 (N_9488,N_8268,N_8379);
and U9489 (N_9489,N_8355,N_8313);
nor U9490 (N_9490,N_8985,N_8972);
nand U9491 (N_9491,N_8101,N_8670);
and U9492 (N_9492,N_8666,N_8633);
nor U9493 (N_9493,N_8921,N_8418);
and U9494 (N_9494,N_8232,N_8053);
nand U9495 (N_9495,N_8806,N_8802);
xnor U9496 (N_9496,N_8708,N_8591);
nor U9497 (N_9497,N_8812,N_8754);
or U9498 (N_9498,N_8246,N_8639);
and U9499 (N_9499,N_8415,N_8372);
nand U9500 (N_9500,N_8744,N_8300);
or U9501 (N_9501,N_8697,N_8206);
nand U9502 (N_9502,N_8664,N_8789);
and U9503 (N_9503,N_8081,N_8576);
and U9504 (N_9504,N_8930,N_8280);
nor U9505 (N_9505,N_8248,N_8433);
or U9506 (N_9506,N_8606,N_8749);
or U9507 (N_9507,N_8689,N_8896);
and U9508 (N_9508,N_8866,N_8847);
and U9509 (N_9509,N_8004,N_8338);
nand U9510 (N_9510,N_8163,N_8753);
and U9511 (N_9511,N_8731,N_8247);
or U9512 (N_9512,N_8692,N_8064);
or U9513 (N_9513,N_8601,N_8906);
or U9514 (N_9514,N_8399,N_8756);
xnor U9515 (N_9515,N_8699,N_8367);
nor U9516 (N_9516,N_8606,N_8433);
or U9517 (N_9517,N_8699,N_8900);
and U9518 (N_9518,N_8989,N_8278);
nand U9519 (N_9519,N_8493,N_8316);
and U9520 (N_9520,N_8747,N_8332);
xnor U9521 (N_9521,N_8843,N_8012);
nand U9522 (N_9522,N_8924,N_8105);
and U9523 (N_9523,N_8866,N_8812);
and U9524 (N_9524,N_8537,N_8310);
nor U9525 (N_9525,N_8249,N_8662);
or U9526 (N_9526,N_8561,N_8152);
or U9527 (N_9527,N_8641,N_8053);
and U9528 (N_9528,N_8701,N_8695);
and U9529 (N_9529,N_8259,N_8566);
nand U9530 (N_9530,N_8663,N_8215);
or U9531 (N_9531,N_8023,N_8671);
nand U9532 (N_9532,N_8818,N_8726);
and U9533 (N_9533,N_8094,N_8777);
nor U9534 (N_9534,N_8036,N_8682);
nand U9535 (N_9535,N_8548,N_8341);
nor U9536 (N_9536,N_8077,N_8151);
and U9537 (N_9537,N_8103,N_8300);
nor U9538 (N_9538,N_8100,N_8734);
nand U9539 (N_9539,N_8765,N_8854);
and U9540 (N_9540,N_8936,N_8478);
or U9541 (N_9541,N_8850,N_8780);
nor U9542 (N_9542,N_8404,N_8904);
nand U9543 (N_9543,N_8116,N_8686);
and U9544 (N_9544,N_8043,N_8880);
nor U9545 (N_9545,N_8103,N_8225);
nand U9546 (N_9546,N_8451,N_8622);
or U9547 (N_9547,N_8990,N_8620);
nor U9548 (N_9548,N_8967,N_8852);
or U9549 (N_9549,N_8624,N_8365);
nand U9550 (N_9550,N_8526,N_8595);
and U9551 (N_9551,N_8749,N_8052);
nor U9552 (N_9552,N_8323,N_8774);
nor U9553 (N_9553,N_8967,N_8214);
or U9554 (N_9554,N_8250,N_8887);
and U9555 (N_9555,N_8915,N_8045);
nor U9556 (N_9556,N_8161,N_8941);
or U9557 (N_9557,N_8778,N_8617);
nor U9558 (N_9558,N_8401,N_8637);
and U9559 (N_9559,N_8832,N_8580);
nor U9560 (N_9560,N_8058,N_8703);
nor U9561 (N_9561,N_8866,N_8005);
and U9562 (N_9562,N_8128,N_8025);
nor U9563 (N_9563,N_8976,N_8655);
nor U9564 (N_9564,N_8354,N_8762);
or U9565 (N_9565,N_8294,N_8923);
or U9566 (N_9566,N_8853,N_8671);
and U9567 (N_9567,N_8385,N_8850);
and U9568 (N_9568,N_8039,N_8432);
nand U9569 (N_9569,N_8524,N_8387);
and U9570 (N_9570,N_8688,N_8827);
or U9571 (N_9571,N_8803,N_8535);
nand U9572 (N_9572,N_8412,N_8677);
or U9573 (N_9573,N_8179,N_8442);
or U9574 (N_9574,N_8477,N_8098);
xor U9575 (N_9575,N_8683,N_8929);
and U9576 (N_9576,N_8611,N_8572);
or U9577 (N_9577,N_8248,N_8883);
and U9578 (N_9578,N_8716,N_8943);
or U9579 (N_9579,N_8757,N_8827);
nand U9580 (N_9580,N_8540,N_8158);
nor U9581 (N_9581,N_8624,N_8041);
nand U9582 (N_9582,N_8782,N_8338);
and U9583 (N_9583,N_8448,N_8467);
nor U9584 (N_9584,N_8268,N_8101);
nand U9585 (N_9585,N_8791,N_8813);
nor U9586 (N_9586,N_8013,N_8918);
nor U9587 (N_9587,N_8610,N_8020);
and U9588 (N_9588,N_8039,N_8348);
nand U9589 (N_9589,N_8698,N_8870);
and U9590 (N_9590,N_8132,N_8417);
nor U9591 (N_9591,N_8217,N_8846);
nor U9592 (N_9592,N_8472,N_8105);
nand U9593 (N_9593,N_8528,N_8386);
and U9594 (N_9594,N_8316,N_8993);
nand U9595 (N_9595,N_8135,N_8719);
and U9596 (N_9596,N_8134,N_8847);
or U9597 (N_9597,N_8413,N_8795);
nand U9598 (N_9598,N_8876,N_8920);
or U9599 (N_9599,N_8004,N_8330);
and U9600 (N_9600,N_8466,N_8671);
and U9601 (N_9601,N_8218,N_8875);
nor U9602 (N_9602,N_8484,N_8263);
or U9603 (N_9603,N_8350,N_8263);
and U9604 (N_9604,N_8736,N_8358);
nor U9605 (N_9605,N_8295,N_8827);
nand U9606 (N_9606,N_8420,N_8577);
or U9607 (N_9607,N_8681,N_8434);
and U9608 (N_9608,N_8127,N_8407);
or U9609 (N_9609,N_8454,N_8697);
or U9610 (N_9610,N_8610,N_8316);
nor U9611 (N_9611,N_8813,N_8208);
nor U9612 (N_9612,N_8274,N_8135);
or U9613 (N_9613,N_8952,N_8151);
and U9614 (N_9614,N_8186,N_8289);
or U9615 (N_9615,N_8193,N_8016);
nor U9616 (N_9616,N_8018,N_8951);
nand U9617 (N_9617,N_8226,N_8703);
and U9618 (N_9618,N_8295,N_8299);
nand U9619 (N_9619,N_8049,N_8010);
or U9620 (N_9620,N_8752,N_8135);
and U9621 (N_9621,N_8117,N_8770);
and U9622 (N_9622,N_8641,N_8788);
nand U9623 (N_9623,N_8162,N_8342);
and U9624 (N_9624,N_8215,N_8093);
nand U9625 (N_9625,N_8405,N_8392);
and U9626 (N_9626,N_8983,N_8078);
nor U9627 (N_9627,N_8601,N_8606);
nor U9628 (N_9628,N_8916,N_8939);
and U9629 (N_9629,N_8818,N_8839);
nand U9630 (N_9630,N_8759,N_8468);
and U9631 (N_9631,N_8126,N_8365);
or U9632 (N_9632,N_8738,N_8149);
nand U9633 (N_9633,N_8823,N_8268);
and U9634 (N_9634,N_8673,N_8395);
nor U9635 (N_9635,N_8541,N_8082);
or U9636 (N_9636,N_8216,N_8590);
nor U9637 (N_9637,N_8367,N_8006);
nand U9638 (N_9638,N_8585,N_8095);
or U9639 (N_9639,N_8601,N_8654);
or U9640 (N_9640,N_8726,N_8416);
or U9641 (N_9641,N_8733,N_8446);
nor U9642 (N_9642,N_8808,N_8678);
and U9643 (N_9643,N_8837,N_8610);
or U9644 (N_9644,N_8565,N_8966);
nor U9645 (N_9645,N_8176,N_8439);
nand U9646 (N_9646,N_8533,N_8733);
or U9647 (N_9647,N_8650,N_8050);
and U9648 (N_9648,N_8077,N_8476);
or U9649 (N_9649,N_8372,N_8685);
and U9650 (N_9650,N_8736,N_8426);
xor U9651 (N_9651,N_8282,N_8639);
nand U9652 (N_9652,N_8780,N_8089);
nor U9653 (N_9653,N_8488,N_8230);
nor U9654 (N_9654,N_8291,N_8849);
and U9655 (N_9655,N_8084,N_8653);
and U9656 (N_9656,N_8756,N_8445);
or U9657 (N_9657,N_8705,N_8683);
or U9658 (N_9658,N_8535,N_8955);
and U9659 (N_9659,N_8832,N_8535);
and U9660 (N_9660,N_8532,N_8795);
and U9661 (N_9661,N_8683,N_8347);
nand U9662 (N_9662,N_8496,N_8278);
nor U9663 (N_9663,N_8925,N_8585);
nand U9664 (N_9664,N_8738,N_8727);
or U9665 (N_9665,N_8300,N_8056);
or U9666 (N_9666,N_8589,N_8241);
nand U9667 (N_9667,N_8039,N_8524);
nor U9668 (N_9668,N_8490,N_8131);
and U9669 (N_9669,N_8316,N_8181);
nand U9670 (N_9670,N_8801,N_8078);
and U9671 (N_9671,N_8855,N_8472);
or U9672 (N_9672,N_8751,N_8825);
or U9673 (N_9673,N_8249,N_8996);
or U9674 (N_9674,N_8725,N_8083);
or U9675 (N_9675,N_8290,N_8308);
or U9676 (N_9676,N_8718,N_8595);
nor U9677 (N_9677,N_8245,N_8610);
and U9678 (N_9678,N_8380,N_8315);
nor U9679 (N_9679,N_8016,N_8135);
or U9680 (N_9680,N_8982,N_8952);
nand U9681 (N_9681,N_8770,N_8718);
and U9682 (N_9682,N_8952,N_8098);
and U9683 (N_9683,N_8771,N_8100);
nand U9684 (N_9684,N_8571,N_8526);
nor U9685 (N_9685,N_8244,N_8549);
and U9686 (N_9686,N_8109,N_8127);
nand U9687 (N_9687,N_8250,N_8884);
nor U9688 (N_9688,N_8268,N_8359);
and U9689 (N_9689,N_8674,N_8177);
and U9690 (N_9690,N_8917,N_8518);
or U9691 (N_9691,N_8232,N_8054);
nand U9692 (N_9692,N_8298,N_8958);
nor U9693 (N_9693,N_8074,N_8142);
nor U9694 (N_9694,N_8329,N_8706);
or U9695 (N_9695,N_8462,N_8354);
nor U9696 (N_9696,N_8101,N_8199);
nor U9697 (N_9697,N_8146,N_8505);
or U9698 (N_9698,N_8005,N_8692);
and U9699 (N_9699,N_8431,N_8528);
and U9700 (N_9700,N_8967,N_8062);
and U9701 (N_9701,N_8140,N_8963);
and U9702 (N_9702,N_8106,N_8864);
or U9703 (N_9703,N_8168,N_8563);
or U9704 (N_9704,N_8315,N_8704);
or U9705 (N_9705,N_8287,N_8719);
nor U9706 (N_9706,N_8290,N_8483);
and U9707 (N_9707,N_8655,N_8100);
nor U9708 (N_9708,N_8001,N_8703);
and U9709 (N_9709,N_8075,N_8247);
or U9710 (N_9710,N_8512,N_8155);
nand U9711 (N_9711,N_8387,N_8518);
and U9712 (N_9712,N_8517,N_8285);
nor U9713 (N_9713,N_8412,N_8578);
nor U9714 (N_9714,N_8307,N_8093);
or U9715 (N_9715,N_8362,N_8816);
and U9716 (N_9716,N_8469,N_8151);
nand U9717 (N_9717,N_8950,N_8366);
xor U9718 (N_9718,N_8155,N_8571);
nor U9719 (N_9719,N_8612,N_8849);
and U9720 (N_9720,N_8851,N_8209);
or U9721 (N_9721,N_8801,N_8900);
nor U9722 (N_9722,N_8856,N_8812);
and U9723 (N_9723,N_8630,N_8746);
and U9724 (N_9724,N_8271,N_8771);
nor U9725 (N_9725,N_8569,N_8243);
nor U9726 (N_9726,N_8293,N_8204);
or U9727 (N_9727,N_8921,N_8667);
nand U9728 (N_9728,N_8506,N_8218);
and U9729 (N_9729,N_8736,N_8075);
nand U9730 (N_9730,N_8714,N_8760);
or U9731 (N_9731,N_8006,N_8782);
nand U9732 (N_9732,N_8702,N_8912);
nand U9733 (N_9733,N_8849,N_8628);
and U9734 (N_9734,N_8806,N_8624);
nor U9735 (N_9735,N_8853,N_8348);
and U9736 (N_9736,N_8568,N_8677);
nand U9737 (N_9737,N_8359,N_8385);
and U9738 (N_9738,N_8588,N_8913);
nand U9739 (N_9739,N_8928,N_8705);
nand U9740 (N_9740,N_8917,N_8043);
nor U9741 (N_9741,N_8718,N_8204);
or U9742 (N_9742,N_8013,N_8130);
and U9743 (N_9743,N_8491,N_8719);
nor U9744 (N_9744,N_8881,N_8430);
and U9745 (N_9745,N_8477,N_8227);
nor U9746 (N_9746,N_8800,N_8656);
nor U9747 (N_9747,N_8889,N_8380);
or U9748 (N_9748,N_8411,N_8402);
nor U9749 (N_9749,N_8261,N_8225);
or U9750 (N_9750,N_8464,N_8403);
or U9751 (N_9751,N_8929,N_8319);
and U9752 (N_9752,N_8918,N_8997);
or U9753 (N_9753,N_8263,N_8288);
and U9754 (N_9754,N_8402,N_8901);
nand U9755 (N_9755,N_8746,N_8261);
and U9756 (N_9756,N_8095,N_8369);
and U9757 (N_9757,N_8974,N_8385);
nor U9758 (N_9758,N_8324,N_8673);
and U9759 (N_9759,N_8169,N_8391);
and U9760 (N_9760,N_8810,N_8141);
nor U9761 (N_9761,N_8769,N_8002);
and U9762 (N_9762,N_8548,N_8338);
and U9763 (N_9763,N_8559,N_8882);
or U9764 (N_9764,N_8353,N_8530);
nor U9765 (N_9765,N_8545,N_8992);
nand U9766 (N_9766,N_8075,N_8307);
nand U9767 (N_9767,N_8395,N_8645);
or U9768 (N_9768,N_8329,N_8615);
nand U9769 (N_9769,N_8516,N_8418);
nor U9770 (N_9770,N_8619,N_8513);
nor U9771 (N_9771,N_8933,N_8494);
nand U9772 (N_9772,N_8824,N_8965);
nand U9773 (N_9773,N_8592,N_8796);
or U9774 (N_9774,N_8803,N_8279);
nor U9775 (N_9775,N_8064,N_8962);
nand U9776 (N_9776,N_8600,N_8626);
or U9777 (N_9777,N_8301,N_8090);
nand U9778 (N_9778,N_8075,N_8096);
and U9779 (N_9779,N_8603,N_8397);
nor U9780 (N_9780,N_8345,N_8708);
nand U9781 (N_9781,N_8901,N_8149);
and U9782 (N_9782,N_8078,N_8273);
nor U9783 (N_9783,N_8892,N_8152);
or U9784 (N_9784,N_8420,N_8473);
nand U9785 (N_9785,N_8837,N_8691);
or U9786 (N_9786,N_8800,N_8890);
nor U9787 (N_9787,N_8497,N_8178);
and U9788 (N_9788,N_8699,N_8671);
or U9789 (N_9789,N_8157,N_8880);
nor U9790 (N_9790,N_8500,N_8460);
or U9791 (N_9791,N_8850,N_8065);
nor U9792 (N_9792,N_8400,N_8749);
and U9793 (N_9793,N_8761,N_8974);
nor U9794 (N_9794,N_8999,N_8869);
nand U9795 (N_9795,N_8203,N_8476);
or U9796 (N_9796,N_8517,N_8477);
nor U9797 (N_9797,N_8900,N_8169);
and U9798 (N_9798,N_8059,N_8443);
and U9799 (N_9799,N_8363,N_8620);
and U9800 (N_9800,N_8615,N_8577);
nand U9801 (N_9801,N_8589,N_8027);
nand U9802 (N_9802,N_8536,N_8838);
or U9803 (N_9803,N_8971,N_8289);
nand U9804 (N_9804,N_8239,N_8861);
or U9805 (N_9805,N_8788,N_8454);
or U9806 (N_9806,N_8233,N_8607);
or U9807 (N_9807,N_8602,N_8671);
and U9808 (N_9808,N_8241,N_8767);
or U9809 (N_9809,N_8834,N_8403);
and U9810 (N_9810,N_8269,N_8621);
and U9811 (N_9811,N_8264,N_8401);
or U9812 (N_9812,N_8230,N_8106);
and U9813 (N_9813,N_8144,N_8522);
nand U9814 (N_9814,N_8653,N_8616);
nand U9815 (N_9815,N_8943,N_8360);
or U9816 (N_9816,N_8848,N_8291);
and U9817 (N_9817,N_8587,N_8354);
or U9818 (N_9818,N_8454,N_8468);
or U9819 (N_9819,N_8274,N_8870);
nor U9820 (N_9820,N_8425,N_8699);
and U9821 (N_9821,N_8083,N_8912);
nand U9822 (N_9822,N_8406,N_8694);
and U9823 (N_9823,N_8426,N_8212);
and U9824 (N_9824,N_8849,N_8737);
nand U9825 (N_9825,N_8933,N_8983);
and U9826 (N_9826,N_8336,N_8740);
xnor U9827 (N_9827,N_8236,N_8560);
and U9828 (N_9828,N_8345,N_8573);
nor U9829 (N_9829,N_8054,N_8007);
and U9830 (N_9830,N_8215,N_8249);
nor U9831 (N_9831,N_8049,N_8409);
nor U9832 (N_9832,N_8454,N_8036);
nor U9833 (N_9833,N_8105,N_8821);
xor U9834 (N_9834,N_8492,N_8416);
nand U9835 (N_9835,N_8595,N_8696);
nand U9836 (N_9836,N_8370,N_8857);
and U9837 (N_9837,N_8531,N_8059);
or U9838 (N_9838,N_8073,N_8342);
nor U9839 (N_9839,N_8070,N_8978);
nand U9840 (N_9840,N_8501,N_8868);
and U9841 (N_9841,N_8617,N_8276);
or U9842 (N_9842,N_8104,N_8208);
and U9843 (N_9843,N_8350,N_8007);
or U9844 (N_9844,N_8139,N_8238);
nand U9845 (N_9845,N_8811,N_8063);
nor U9846 (N_9846,N_8737,N_8987);
nor U9847 (N_9847,N_8696,N_8508);
nand U9848 (N_9848,N_8450,N_8813);
nor U9849 (N_9849,N_8409,N_8025);
or U9850 (N_9850,N_8578,N_8793);
or U9851 (N_9851,N_8149,N_8539);
nand U9852 (N_9852,N_8539,N_8598);
or U9853 (N_9853,N_8375,N_8119);
or U9854 (N_9854,N_8761,N_8796);
nand U9855 (N_9855,N_8164,N_8994);
and U9856 (N_9856,N_8576,N_8031);
or U9857 (N_9857,N_8480,N_8687);
and U9858 (N_9858,N_8494,N_8771);
and U9859 (N_9859,N_8323,N_8417);
or U9860 (N_9860,N_8949,N_8584);
nand U9861 (N_9861,N_8148,N_8770);
nand U9862 (N_9862,N_8948,N_8737);
or U9863 (N_9863,N_8036,N_8523);
and U9864 (N_9864,N_8915,N_8654);
and U9865 (N_9865,N_8607,N_8990);
and U9866 (N_9866,N_8522,N_8834);
nor U9867 (N_9867,N_8993,N_8132);
nand U9868 (N_9868,N_8944,N_8389);
nand U9869 (N_9869,N_8487,N_8029);
nor U9870 (N_9870,N_8424,N_8149);
or U9871 (N_9871,N_8671,N_8406);
nand U9872 (N_9872,N_8267,N_8058);
nor U9873 (N_9873,N_8537,N_8114);
or U9874 (N_9874,N_8018,N_8510);
or U9875 (N_9875,N_8518,N_8107);
nand U9876 (N_9876,N_8597,N_8426);
nand U9877 (N_9877,N_8402,N_8994);
nand U9878 (N_9878,N_8659,N_8879);
nor U9879 (N_9879,N_8360,N_8188);
nor U9880 (N_9880,N_8506,N_8289);
or U9881 (N_9881,N_8080,N_8259);
nor U9882 (N_9882,N_8489,N_8805);
nor U9883 (N_9883,N_8731,N_8608);
nor U9884 (N_9884,N_8023,N_8167);
and U9885 (N_9885,N_8516,N_8345);
or U9886 (N_9886,N_8597,N_8438);
or U9887 (N_9887,N_8232,N_8070);
nand U9888 (N_9888,N_8427,N_8760);
and U9889 (N_9889,N_8632,N_8764);
and U9890 (N_9890,N_8710,N_8367);
nor U9891 (N_9891,N_8751,N_8369);
nor U9892 (N_9892,N_8934,N_8203);
nor U9893 (N_9893,N_8660,N_8421);
nor U9894 (N_9894,N_8458,N_8941);
nor U9895 (N_9895,N_8289,N_8453);
nand U9896 (N_9896,N_8567,N_8863);
nand U9897 (N_9897,N_8942,N_8600);
and U9898 (N_9898,N_8743,N_8022);
nor U9899 (N_9899,N_8588,N_8490);
nor U9900 (N_9900,N_8163,N_8281);
xnor U9901 (N_9901,N_8615,N_8021);
and U9902 (N_9902,N_8204,N_8687);
or U9903 (N_9903,N_8774,N_8145);
nor U9904 (N_9904,N_8330,N_8860);
and U9905 (N_9905,N_8848,N_8851);
and U9906 (N_9906,N_8689,N_8102);
nand U9907 (N_9907,N_8650,N_8641);
nor U9908 (N_9908,N_8096,N_8011);
and U9909 (N_9909,N_8561,N_8053);
or U9910 (N_9910,N_8755,N_8683);
nor U9911 (N_9911,N_8158,N_8268);
nand U9912 (N_9912,N_8172,N_8675);
nor U9913 (N_9913,N_8314,N_8587);
nor U9914 (N_9914,N_8737,N_8844);
nand U9915 (N_9915,N_8660,N_8785);
and U9916 (N_9916,N_8979,N_8400);
nor U9917 (N_9917,N_8623,N_8045);
and U9918 (N_9918,N_8034,N_8032);
or U9919 (N_9919,N_8937,N_8463);
nand U9920 (N_9920,N_8080,N_8096);
or U9921 (N_9921,N_8869,N_8748);
or U9922 (N_9922,N_8801,N_8752);
nand U9923 (N_9923,N_8180,N_8471);
or U9924 (N_9924,N_8978,N_8331);
or U9925 (N_9925,N_8934,N_8213);
and U9926 (N_9926,N_8229,N_8713);
nand U9927 (N_9927,N_8315,N_8868);
and U9928 (N_9928,N_8521,N_8831);
nor U9929 (N_9929,N_8579,N_8186);
and U9930 (N_9930,N_8193,N_8355);
nand U9931 (N_9931,N_8436,N_8690);
nand U9932 (N_9932,N_8345,N_8458);
nand U9933 (N_9933,N_8029,N_8537);
or U9934 (N_9934,N_8910,N_8634);
nor U9935 (N_9935,N_8057,N_8191);
nand U9936 (N_9936,N_8002,N_8512);
or U9937 (N_9937,N_8553,N_8235);
nand U9938 (N_9938,N_8145,N_8197);
or U9939 (N_9939,N_8024,N_8176);
and U9940 (N_9940,N_8293,N_8615);
and U9941 (N_9941,N_8290,N_8148);
or U9942 (N_9942,N_8918,N_8793);
nand U9943 (N_9943,N_8228,N_8372);
nor U9944 (N_9944,N_8821,N_8006);
or U9945 (N_9945,N_8782,N_8075);
and U9946 (N_9946,N_8191,N_8901);
nand U9947 (N_9947,N_8730,N_8372);
nand U9948 (N_9948,N_8775,N_8455);
nor U9949 (N_9949,N_8159,N_8973);
and U9950 (N_9950,N_8171,N_8908);
and U9951 (N_9951,N_8722,N_8410);
nand U9952 (N_9952,N_8978,N_8397);
nor U9953 (N_9953,N_8039,N_8019);
and U9954 (N_9954,N_8410,N_8919);
nand U9955 (N_9955,N_8150,N_8995);
nand U9956 (N_9956,N_8731,N_8226);
nand U9957 (N_9957,N_8550,N_8147);
and U9958 (N_9958,N_8426,N_8302);
nor U9959 (N_9959,N_8463,N_8732);
nand U9960 (N_9960,N_8730,N_8775);
and U9961 (N_9961,N_8773,N_8389);
nor U9962 (N_9962,N_8823,N_8735);
and U9963 (N_9963,N_8367,N_8484);
nand U9964 (N_9964,N_8234,N_8651);
nand U9965 (N_9965,N_8555,N_8214);
xor U9966 (N_9966,N_8281,N_8912);
nor U9967 (N_9967,N_8161,N_8375);
or U9968 (N_9968,N_8100,N_8795);
or U9969 (N_9969,N_8848,N_8237);
nor U9970 (N_9970,N_8629,N_8116);
or U9971 (N_9971,N_8532,N_8160);
nor U9972 (N_9972,N_8984,N_8762);
and U9973 (N_9973,N_8332,N_8270);
and U9974 (N_9974,N_8215,N_8930);
nor U9975 (N_9975,N_8447,N_8699);
nand U9976 (N_9976,N_8101,N_8997);
nor U9977 (N_9977,N_8991,N_8850);
nand U9978 (N_9978,N_8772,N_8820);
nand U9979 (N_9979,N_8166,N_8977);
nand U9980 (N_9980,N_8258,N_8916);
nor U9981 (N_9981,N_8724,N_8377);
nand U9982 (N_9982,N_8571,N_8429);
or U9983 (N_9983,N_8964,N_8505);
nand U9984 (N_9984,N_8309,N_8979);
nand U9985 (N_9985,N_8702,N_8919);
nand U9986 (N_9986,N_8243,N_8108);
nor U9987 (N_9987,N_8593,N_8267);
and U9988 (N_9988,N_8663,N_8001);
or U9989 (N_9989,N_8576,N_8324);
and U9990 (N_9990,N_8059,N_8022);
nor U9991 (N_9991,N_8199,N_8204);
or U9992 (N_9992,N_8523,N_8466);
or U9993 (N_9993,N_8993,N_8185);
or U9994 (N_9994,N_8708,N_8265);
nand U9995 (N_9995,N_8566,N_8500);
or U9996 (N_9996,N_8267,N_8719);
nand U9997 (N_9997,N_8688,N_8476);
nor U9998 (N_9998,N_8495,N_8357);
and U9999 (N_9999,N_8923,N_8253);
nand U10000 (N_10000,N_9565,N_9177);
nor U10001 (N_10001,N_9933,N_9663);
xor U10002 (N_10002,N_9907,N_9976);
nand U10003 (N_10003,N_9748,N_9382);
nor U10004 (N_10004,N_9231,N_9316);
and U10005 (N_10005,N_9846,N_9902);
nor U10006 (N_10006,N_9474,N_9550);
or U10007 (N_10007,N_9359,N_9242);
or U10008 (N_10008,N_9763,N_9900);
and U10009 (N_10009,N_9878,N_9221);
nor U10010 (N_10010,N_9125,N_9817);
or U10011 (N_10011,N_9313,N_9455);
or U10012 (N_10012,N_9969,N_9584);
or U10013 (N_10013,N_9533,N_9184);
nand U10014 (N_10014,N_9349,N_9091);
and U10015 (N_10015,N_9200,N_9682);
and U10016 (N_10016,N_9440,N_9097);
nor U10017 (N_10017,N_9758,N_9771);
and U10018 (N_10018,N_9942,N_9258);
nor U10019 (N_10019,N_9409,N_9241);
and U10020 (N_10020,N_9862,N_9454);
and U10021 (N_10021,N_9496,N_9248);
nand U10022 (N_10022,N_9710,N_9483);
or U10023 (N_10023,N_9290,N_9443);
nor U10024 (N_10024,N_9583,N_9743);
nor U10025 (N_10025,N_9800,N_9792);
and U10026 (N_10026,N_9595,N_9538);
nand U10027 (N_10027,N_9661,N_9752);
and U10028 (N_10028,N_9611,N_9946);
or U10029 (N_10029,N_9259,N_9963);
or U10030 (N_10030,N_9145,N_9022);
and U10031 (N_10031,N_9340,N_9903);
nor U10032 (N_10032,N_9066,N_9686);
and U10033 (N_10033,N_9732,N_9670);
nor U10034 (N_10034,N_9726,N_9169);
or U10035 (N_10035,N_9618,N_9815);
nand U10036 (N_10036,N_9772,N_9322);
and U10037 (N_10037,N_9479,N_9343);
or U10038 (N_10038,N_9502,N_9991);
nor U10039 (N_10039,N_9674,N_9228);
nand U10040 (N_10040,N_9109,N_9396);
and U10041 (N_10041,N_9196,N_9139);
nand U10042 (N_10042,N_9117,N_9769);
and U10043 (N_10043,N_9958,N_9744);
nor U10044 (N_10044,N_9971,N_9999);
and U10045 (N_10045,N_9959,N_9143);
or U10046 (N_10046,N_9041,N_9943);
and U10047 (N_10047,N_9233,N_9503);
nand U10048 (N_10048,N_9014,N_9548);
or U10049 (N_10049,N_9968,N_9468);
and U10050 (N_10050,N_9446,N_9577);
or U10051 (N_10051,N_9337,N_9941);
or U10052 (N_10052,N_9362,N_9456);
and U10053 (N_10053,N_9694,N_9247);
nand U10054 (N_10054,N_9069,N_9168);
or U10055 (N_10055,N_9731,N_9688);
nor U10056 (N_10056,N_9605,N_9552);
nor U10057 (N_10057,N_9499,N_9011);
nor U10058 (N_10058,N_9534,N_9255);
nor U10059 (N_10059,N_9910,N_9784);
and U10060 (N_10060,N_9957,N_9882);
or U10061 (N_10061,N_9916,N_9111);
or U10062 (N_10062,N_9972,N_9647);
or U10063 (N_10063,N_9436,N_9394);
or U10064 (N_10064,N_9803,N_9016);
nand U10065 (N_10065,N_9852,N_9819);
and U10066 (N_10066,N_9604,N_9720);
and U10067 (N_10067,N_9914,N_9851);
or U10068 (N_10068,N_9315,N_9360);
nor U10069 (N_10069,N_9229,N_9628);
and U10070 (N_10070,N_9045,N_9966);
nand U10071 (N_10071,N_9240,N_9642);
nor U10072 (N_10072,N_9660,N_9201);
and U10073 (N_10073,N_9459,N_9312);
or U10074 (N_10074,N_9094,N_9325);
or U10075 (N_10075,N_9600,N_9239);
nor U10076 (N_10076,N_9765,N_9853);
nor U10077 (N_10077,N_9634,N_9980);
and U10078 (N_10078,N_9612,N_9385);
nor U10079 (N_10079,N_9261,N_9149);
and U10080 (N_10080,N_9133,N_9112);
nand U10081 (N_10081,N_9932,N_9633);
or U10082 (N_10082,N_9896,N_9831);
nor U10083 (N_10083,N_9469,N_9345);
nor U10084 (N_10084,N_9064,N_9392);
nor U10085 (N_10085,N_9764,N_9774);
nand U10086 (N_10086,N_9408,N_9141);
nand U10087 (N_10087,N_9637,N_9861);
or U10088 (N_10088,N_9281,N_9063);
and U10089 (N_10089,N_9323,N_9842);
nand U10090 (N_10090,N_9737,N_9414);
nand U10091 (N_10091,N_9830,N_9378);
nor U10092 (N_10092,N_9400,N_9371);
xnor U10093 (N_10093,N_9978,N_9926);
nor U10094 (N_10094,N_9442,N_9755);
nand U10095 (N_10095,N_9954,N_9477);
or U10096 (N_10096,N_9529,N_9592);
and U10097 (N_10097,N_9568,N_9101);
and U10098 (N_10098,N_9614,N_9865);
nor U10099 (N_10099,N_9386,N_9104);
nor U10100 (N_10100,N_9730,N_9489);
or U10101 (N_10101,N_9844,N_9977);
nand U10102 (N_10102,N_9825,N_9357);
nand U10103 (N_10103,N_9286,N_9399);
nand U10104 (N_10104,N_9300,N_9164);
and U10105 (N_10105,N_9782,N_9249);
and U10106 (N_10106,N_9673,N_9656);
nor U10107 (N_10107,N_9301,N_9823);
nor U10108 (N_10108,N_9330,N_9582);
or U10109 (N_10109,N_9662,N_9197);
nand U10110 (N_10110,N_9355,N_9307);
nand U10111 (N_10111,N_9993,N_9339);
nand U10112 (N_10112,N_9348,N_9713);
or U10113 (N_10113,N_9571,N_9645);
or U10114 (N_10114,N_9036,N_9346);
nor U10115 (N_10115,N_9146,N_9653);
and U10116 (N_10116,N_9873,N_9018);
nor U10117 (N_10117,N_9812,N_9756);
nand U10118 (N_10118,N_9155,N_9027);
nor U10119 (N_10119,N_9945,N_9938);
nand U10120 (N_10120,N_9344,N_9911);
nand U10121 (N_10121,N_9198,N_9319);
nand U10122 (N_10122,N_9585,N_9947);
nor U10123 (N_10123,N_9975,N_9162);
nand U10124 (N_10124,N_9740,N_9147);
nor U10125 (N_10125,N_9875,N_9078);
nand U10126 (N_10126,N_9292,N_9203);
and U10127 (N_10127,N_9361,N_9305);
nand U10128 (N_10128,N_9212,N_9033);
nand U10129 (N_10129,N_9423,N_9789);
nand U10130 (N_10130,N_9032,N_9961);
nand U10131 (N_10131,N_9106,N_9519);
and U10132 (N_10132,N_9920,N_9025);
nor U10133 (N_10133,N_9620,N_9320);
nor U10134 (N_10134,N_9699,N_9126);
and U10135 (N_10135,N_9801,N_9510);
nand U10136 (N_10136,N_9780,N_9257);
nor U10137 (N_10137,N_9759,N_9836);
nor U10138 (N_10138,N_9543,N_9490);
nand U10139 (N_10139,N_9722,N_9799);
or U10140 (N_10140,N_9088,N_9981);
or U10141 (N_10141,N_9296,N_9718);
or U10142 (N_10142,N_9567,N_9291);
nand U10143 (N_10143,N_9429,N_9283);
xnor U10144 (N_10144,N_9691,N_9912);
or U10145 (N_10145,N_9679,N_9165);
nand U10146 (N_10146,N_9504,N_9302);
nor U10147 (N_10147,N_9492,N_9821);
nor U10148 (N_10148,N_9625,N_9497);
nor U10149 (N_10149,N_9950,N_9042);
or U10150 (N_10150,N_9608,N_9988);
and U10151 (N_10151,N_9219,N_9705);
nand U10152 (N_10152,N_9708,N_9176);
nand U10153 (N_10153,N_9530,N_9935);
nand U10154 (N_10154,N_9452,N_9683);
or U10155 (N_10155,N_9603,N_9796);
and U10156 (N_10156,N_9901,N_9967);
nand U10157 (N_10157,N_9835,N_9086);
nand U10158 (N_10158,N_9849,N_9578);
or U10159 (N_10159,N_9401,N_9639);
nand U10160 (N_10160,N_9199,N_9928);
nor U10161 (N_10161,N_9788,N_9115);
nand U10162 (N_10162,N_9453,N_9505);
and U10163 (N_10163,N_9013,N_9417);
nand U10164 (N_10164,N_9557,N_9905);
nand U10165 (N_10165,N_9881,N_9411);
and U10166 (N_10166,N_9513,N_9692);
and U10167 (N_10167,N_9338,N_9331);
or U10168 (N_10168,N_9160,N_9648);
nand U10169 (N_10169,N_9186,N_9246);
nand U10170 (N_10170,N_9471,N_9406);
and U10171 (N_10171,N_9695,N_9965);
or U10172 (N_10172,N_9553,N_9341);
nor U10173 (N_10173,N_9277,N_9668);
nor U10174 (N_10174,N_9706,N_9138);
nand U10175 (N_10175,N_9890,N_9298);
and U10176 (N_10176,N_9591,N_9517);
nand U10177 (N_10177,N_9278,N_9579);
or U10178 (N_10178,N_9480,N_9880);
and U10179 (N_10179,N_9868,N_9264);
and U10180 (N_10180,N_9797,N_9949);
nand U10181 (N_10181,N_9224,N_9093);
and U10182 (N_10182,N_9657,N_9811);
nor U10183 (N_10183,N_9897,N_9824);
nand U10184 (N_10184,N_9217,N_9478);
or U10185 (N_10185,N_9631,N_9092);
nor U10186 (N_10186,N_9415,N_9282);
and U10187 (N_10187,N_9118,N_9791);
and U10188 (N_10188,N_9222,N_9314);
nor U10189 (N_10189,N_9876,N_9883);
nor U10190 (N_10190,N_9485,N_9391);
and U10191 (N_10191,N_9056,N_9745);
or U10192 (N_10192,N_9077,N_9108);
nor U10193 (N_10193,N_9923,N_9623);
xnor U10194 (N_10194,N_9643,N_9974);
or U10195 (N_10195,N_9716,N_9606);
nand U10196 (N_10196,N_9570,N_9472);
nand U10197 (N_10197,N_9098,N_9243);
nor U10198 (N_10198,N_9986,N_9617);
nor U10199 (N_10199,N_9132,N_9735);
nor U10200 (N_10200,N_9170,N_9019);
nand U10201 (N_10201,N_9171,N_9151);
nand U10202 (N_10202,N_9630,N_9488);
and U10203 (N_10203,N_9377,N_9952);
nand U10204 (N_10204,N_9003,N_9150);
nor U10205 (N_10205,N_9253,N_9860);
or U10206 (N_10206,N_9226,N_9757);
nand U10207 (N_10207,N_9798,N_9012);
or U10208 (N_10208,N_9616,N_9421);
nand U10209 (N_10209,N_9924,N_9393);
nor U10210 (N_10210,N_9299,N_9058);
and U10211 (N_10211,N_9736,N_9641);
and U10212 (N_10212,N_9029,N_9794);
nand U10213 (N_10213,N_9651,N_9351);
and U10214 (N_10214,N_9712,N_9665);
and U10215 (N_10215,N_9274,N_9114);
nor U10216 (N_10216,N_9425,N_9754);
and U10217 (N_10217,N_9805,N_9742);
and U10218 (N_10218,N_9137,N_9829);
nand U10219 (N_10219,N_9157,N_9515);
nand U10220 (N_10220,N_9540,N_9163);
or U10221 (N_10221,N_9470,N_9659);
nand U10222 (N_10222,N_9609,N_9894);
xnor U10223 (N_10223,N_9702,N_9367);
nor U10224 (N_10224,N_9580,N_9887);
or U10225 (N_10225,N_9675,N_9318);
nand U10226 (N_10226,N_9514,N_9328);
nand U10227 (N_10227,N_9687,N_9384);
and U10228 (N_10228,N_9287,N_9937);
nand U10229 (N_10229,N_9619,N_9070);
and U10230 (N_10230,N_9061,N_9395);
and U10231 (N_10231,N_9256,N_9021);
nand U10232 (N_10232,N_9684,N_9715);
nand U10233 (N_10233,N_9227,N_9711);
nor U10234 (N_10234,N_9956,N_9899);
nand U10235 (N_10235,N_9563,N_9273);
nand U10236 (N_10236,N_9463,N_9918);
and U10237 (N_10237,N_9105,N_9590);
nand U10238 (N_10238,N_9481,N_9840);
and U10239 (N_10239,N_9867,N_9407);
or U10240 (N_10240,N_9962,N_9336);
nor U10241 (N_10241,N_9096,N_9549);
or U10242 (N_10242,N_9953,N_9216);
or U10243 (N_10243,N_9944,N_9927);
nand U10244 (N_10244,N_9809,N_9048);
or U10245 (N_10245,N_9770,N_9664);
or U10246 (N_10246,N_9741,N_9178);
or U10247 (N_10247,N_9329,N_9102);
or U10248 (N_10248,N_9363,N_9572);
or U10249 (N_10249,N_9215,N_9704);
or U10250 (N_10250,N_9768,N_9116);
and U10251 (N_10251,N_9484,N_9778);
and U10252 (N_10252,N_9060,N_9214);
nand U10253 (N_10253,N_9297,N_9627);
and U10254 (N_10254,N_9521,N_9095);
or U10255 (N_10255,N_9413,N_9326);
or U10256 (N_10256,N_9593,N_9269);
and U10257 (N_10257,N_9564,N_9026);
or U10258 (N_10258,N_9099,N_9158);
or U10259 (N_10259,N_9375,N_9508);
nand U10260 (N_10260,N_9308,N_9156);
and U10261 (N_10261,N_9276,N_9885);
nor U10262 (N_10262,N_9075,N_9775);
or U10263 (N_10263,N_9310,N_9327);
and U10264 (N_10264,N_9154,N_9934);
and U10265 (N_10265,N_9955,N_9655);
or U10266 (N_10266,N_9826,N_9939);
and U10267 (N_10267,N_9839,N_9244);
or U10268 (N_10268,N_9640,N_9005);
and U10269 (N_10269,N_9236,N_9527);
and U10270 (N_10270,N_9404,N_9051);
and U10271 (N_10271,N_9390,N_9152);
nand U10272 (N_10272,N_9467,N_9250);
nand U10273 (N_10273,N_9810,N_9676);
nor U10274 (N_10274,N_9110,N_9693);
nand U10275 (N_10275,N_9723,N_9951);
and U10276 (N_10276,N_9410,N_9071);
nand U10277 (N_10277,N_9379,N_9816);
nor U10278 (N_10278,N_9002,N_9895);
nor U10279 (N_10279,N_9220,N_9268);
or U10280 (N_10280,N_9893,N_9856);
and U10281 (N_10281,N_9294,N_9696);
or U10282 (N_10282,N_9520,N_9173);
nand U10283 (N_10283,N_9419,N_9245);
or U10284 (N_10284,N_9304,N_9223);
and U10285 (N_10285,N_9350,N_9587);
nor U10286 (N_10286,N_9424,N_9898);
and U10287 (N_10287,N_9669,N_9418);
or U10288 (N_10288,N_9841,N_9877);
nor U10289 (N_10289,N_9370,N_9435);
or U10290 (N_10290,N_9365,N_9008);
or U10291 (N_10291,N_9444,N_9654);
or U10292 (N_10292,N_9272,N_9891);
nor U10293 (N_10293,N_9987,N_9525);
nor U10294 (N_10294,N_9131,N_9624);
and U10295 (N_10295,N_9437,N_9622);
and U10296 (N_10296,N_9059,N_9804);
and U10297 (N_10297,N_9889,N_9028);
or U10298 (N_10298,N_9166,N_9677);
nand U10299 (N_10299,N_9389,N_9597);
and U10300 (N_10300,N_9030,N_9834);
or U10301 (N_10301,N_9303,N_9082);
and U10302 (N_10302,N_9621,N_9858);
nor U10303 (N_10303,N_9855,N_9439);
nand U10304 (N_10304,N_9293,N_9306);
nand U10305 (N_10305,N_9746,N_9122);
nand U10306 (N_10306,N_9596,N_9031);
and U10307 (N_10307,N_9964,N_9536);
nor U10308 (N_10308,N_9973,N_9428);
or U10309 (N_10309,N_9140,N_9172);
and U10310 (N_10310,N_9495,N_9434);
nand U10311 (N_10311,N_9284,N_9506);
nand U10312 (N_10312,N_9050,N_9930);
or U10313 (N_10313,N_9888,N_9646);
nand U10314 (N_10314,N_9235,N_9234);
or U10315 (N_10315,N_9000,N_9120);
nor U10316 (N_10316,N_9103,N_9380);
nor U10317 (N_10317,N_9067,N_9369);
and U10318 (N_10318,N_9501,N_9083);
nor U10319 (N_10319,N_9180,N_9204);
nor U10320 (N_10320,N_9491,N_9984);
nor U10321 (N_10321,N_9864,N_9448);
nand U10322 (N_10322,N_9807,N_9594);
nor U10323 (N_10323,N_9919,N_9317);
xor U10324 (N_10324,N_9561,N_9874);
and U10325 (N_10325,N_9017,N_9279);
nor U10326 (N_10326,N_9832,N_9445);
and U10327 (N_10327,N_9689,N_9649);
nand U10328 (N_10328,N_9678,N_9790);
and U10329 (N_10329,N_9194,N_9827);
nand U10330 (N_10330,N_9144,N_9087);
nand U10331 (N_10331,N_9509,N_9921);
nand U10332 (N_10332,N_9422,N_9431);
or U10333 (N_10333,N_9569,N_9982);
and U10334 (N_10334,N_9680,N_9430);
and U10335 (N_10335,N_9124,N_9667);
nor U10336 (N_10336,N_9024,N_9260);
and U10337 (N_10337,N_9733,N_9813);
or U10338 (N_10338,N_9209,N_9554);
and U10339 (N_10339,N_9522,N_9475);
and U10340 (N_10340,N_9703,N_9237);
or U10341 (N_10341,N_9004,N_9205);
or U10342 (N_10342,N_9588,N_9466);
and U10343 (N_10343,N_9857,N_9929);
and U10344 (N_10344,N_9191,N_9808);
nor U10345 (N_10345,N_9739,N_9206);
or U10346 (N_10346,N_9321,N_9848);
and U10347 (N_10347,N_9034,N_9523);
and U10348 (N_10348,N_9866,N_9761);
or U10349 (N_10349,N_9053,N_9751);
and U10350 (N_10350,N_9188,N_9650);
nor U10351 (N_10351,N_9906,N_9498);
or U10352 (N_10352,N_9979,N_9432);
and U10353 (N_10353,N_9546,N_9107);
xnor U10354 (N_10354,N_9265,N_9698);
or U10355 (N_10355,N_9925,N_9334);
nand U10356 (N_10356,N_9035,N_9054);
and U10357 (N_10357,N_9332,N_9208);
and U10358 (N_10358,N_9535,N_9179);
nor U10359 (N_10359,N_9010,N_9581);
or U10360 (N_10360,N_9562,N_9438);
nand U10361 (N_10361,N_9528,N_9773);
nor U10362 (N_10362,N_9997,N_9190);
nand U10363 (N_10363,N_9983,N_9936);
or U10364 (N_10364,N_9507,N_9181);
nand U10365 (N_10365,N_9374,N_9052);
or U10366 (N_10366,N_9601,N_9762);
and U10367 (N_10367,N_9948,N_9904);
nor U10368 (N_10368,N_9412,N_9285);
and U10369 (N_10369,N_9405,N_9420);
nor U10370 (N_10370,N_9613,N_9129);
nor U10371 (N_10371,N_9749,N_9366);
nor U10372 (N_10372,N_9566,N_9555);
and U10373 (N_10373,N_9252,N_9015);
nor U10374 (N_10374,N_9289,N_9023);
nor U10375 (N_10375,N_9922,N_9725);
nand U10376 (N_10376,N_9068,N_9072);
or U10377 (N_10377,N_9079,N_9074);
nor U10378 (N_10378,N_9065,N_9960);
or U10379 (N_10379,N_9055,N_9863);
or U10380 (N_10380,N_9447,N_9451);
nand U10381 (N_10381,N_9473,N_9822);
nor U10382 (N_10382,N_9460,N_9192);
nand U10383 (N_10383,N_9558,N_9970);
nor U10384 (N_10384,N_9009,N_9892);
nor U10385 (N_10385,N_9161,N_9311);
or U10386 (N_10386,N_9275,N_9576);
nand U10387 (N_10387,N_9006,N_9130);
nand U10388 (N_10388,N_9020,N_9602);
nor U10389 (N_10389,N_9270,N_9870);
and U10390 (N_10390,N_9043,N_9747);
and U10391 (N_10391,N_9869,N_9262);
nor U10392 (N_10392,N_9556,N_9182);
nand U10393 (N_10393,N_9403,N_9714);
nor U10394 (N_10394,N_9493,N_9547);
or U10395 (N_10395,N_9352,N_9781);
and U10396 (N_10396,N_9884,N_9793);
nand U10397 (N_10397,N_9335,N_9760);
nand U10398 (N_10398,N_9787,N_9001);
nor U10399 (N_10399,N_9148,N_9465);
nand U10400 (N_10400,N_9786,N_9128);
nand U10401 (N_10401,N_9402,N_9537);
nand U10402 (N_10402,N_9776,N_9038);
or U10403 (N_10403,N_9607,N_9802);
nand U10404 (N_10404,N_9777,N_9599);
nand U10405 (N_10405,N_9127,N_9090);
or U10406 (N_10406,N_9397,N_9076);
nand U10407 (N_10407,N_9719,N_9511);
or U10408 (N_10408,N_9464,N_9037);
nor U10409 (N_10409,N_9845,N_9398);
and U10410 (N_10410,N_9347,N_9383);
nand U10411 (N_10411,N_9635,N_9218);
nor U10412 (N_10412,N_9872,N_9457);
and U10413 (N_10413,N_9994,N_9724);
and U10414 (N_10414,N_9785,N_9871);
nor U10415 (N_10415,N_9238,N_9193);
and U10416 (N_10416,N_9046,N_9159);
and U10417 (N_10417,N_9427,N_9985);
or U10418 (N_10418,N_9057,N_9820);
and U10419 (N_10419,N_9598,N_9998);
and U10420 (N_10420,N_9462,N_9288);
and U10421 (N_10421,N_9586,N_9119);
and U10422 (N_10422,N_9230,N_9544);
or U10423 (N_10423,N_9610,N_9175);
nand U10424 (N_10424,N_9135,N_9990);
nand U10425 (N_10425,N_9727,N_9734);
nand U10426 (N_10426,N_9142,N_9859);
nand U10427 (N_10427,N_9461,N_9806);
nand U10428 (N_10428,N_9615,N_9373);
nand U10429 (N_10429,N_9263,N_9494);
nor U10430 (N_10430,N_9039,N_9372);
or U10431 (N_10431,N_9211,N_9123);
nand U10432 (N_10432,N_9353,N_9766);
nor U10433 (N_10433,N_9271,N_9526);
or U10434 (N_10434,N_9685,N_9280);
nand U10435 (N_10435,N_9047,N_9915);
nand U10436 (N_10436,N_9189,N_9837);
and U10437 (N_10437,N_9251,N_9210);
and U10438 (N_10438,N_9551,N_9085);
or U10439 (N_10439,N_9658,N_9195);
or U10440 (N_10440,N_9100,N_9167);
or U10441 (N_10441,N_9940,N_9207);
nor U10442 (N_10442,N_9482,N_9795);
or U10443 (N_10443,N_9681,N_9545);
nor U10444 (N_10444,N_9995,N_9376);
nor U10445 (N_10445,N_9254,N_9854);
xnor U10446 (N_10446,N_9458,N_9487);
nand U10447 (N_10447,N_9559,N_9652);
and U10448 (N_10448,N_9381,N_9153);
or U10449 (N_10449,N_9202,N_9574);
or U10450 (N_10450,N_9416,N_9666);
or U10451 (N_10451,N_9783,N_9629);
and U10452 (N_10452,N_9185,N_9542);
nor U10453 (N_10453,N_9886,N_9516);
nand U10454 (N_10454,N_9049,N_9358);
nor U10455 (N_10455,N_9364,N_9518);
nand U10456 (N_10456,N_9931,N_9267);
nor U10457 (N_10457,N_9843,N_9387);
or U10458 (N_10458,N_9136,N_9531);
nand U10459 (N_10459,N_9814,N_9187);
and U10460 (N_10460,N_9709,N_9721);
and U10461 (N_10461,N_9632,N_9589);
or U10462 (N_10462,N_9486,N_9838);
nor U10463 (N_10463,N_9174,N_9909);
and U10464 (N_10464,N_9062,N_9309);
and U10465 (N_10465,N_9626,N_9913);
or U10466 (N_10466,N_9908,N_9992);
nand U10467 (N_10467,N_9750,N_9575);
nor U10468 (N_10468,N_9450,N_9368);
or U10469 (N_10469,N_9539,N_9084);
nand U10470 (N_10470,N_9779,N_9040);
or U10471 (N_10471,N_9644,N_9728);
nor U10472 (N_10472,N_9500,N_9671);
nand U10473 (N_10473,N_9701,N_9818);
or U10474 (N_10474,N_9707,N_9044);
and U10475 (N_10475,N_9532,N_9573);
or U10476 (N_10476,N_9080,N_9638);
and U10477 (N_10477,N_9388,N_9356);
or U10478 (N_10478,N_9636,N_9753);
nand U10479 (N_10479,N_9354,N_9081);
or U10480 (N_10480,N_9996,N_9121);
nand U10481 (N_10481,N_9441,N_9700);
or U10482 (N_10482,N_9828,N_9089);
nor U10483 (N_10483,N_9007,N_9433);
or U10484 (N_10484,N_9476,N_9847);
nand U10485 (N_10485,N_9690,N_9426);
or U10486 (N_10486,N_9113,N_9295);
and U10487 (N_10487,N_9324,N_9183);
nor U10488 (N_10488,N_9225,N_9134);
nand U10489 (N_10489,N_9449,N_9266);
nor U10490 (N_10490,N_9512,N_9541);
nand U10491 (N_10491,N_9333,N_9850);
nand U10492 (N_10492,N_9672,N_9989);
nand U10493 (N_10493,N_9917,N_9073);
or U10494 (N_10494,N_9213,N_9767);
nand U10495 (N_10495,N_9717,N_9697);
nor U10496 (N_10496,N_9879,N_9342);
nand U10497 (N_10497,N_9524,N_9738);
nand U10498 (N_10498,N_9560,N_9833);
or U10499 (N_10499,N_9729,N_9232);
nand U10500 (N_10500,N_9952,N_9178);
or U10501 (N_10501,N_9737,N_9226);
or U10502 (N_10502,N_9378,N_9287);
and U10503 (N_10503,N_9236,N_9825);
and U10504 (N_10504,N_9556,N_9676);
nor U10505 (N_10505,N_9587,N_9220);
nor U10506 (N_10506,N_9704,N_9220);
or U10507 (N_10507,N_9417,N_9556);
or U10508 (N_10508,N_9576,N_9900);
and U10509 (N_10509,N_9262,N_9129);
and U10510 (N_10510,N_9162,N_9789);
nor U10511 (N_10511,N_9619,N_9577);
and U10512 (N_10512,N_9270,N_9160);
or U10513 (N_10513,N_9059,N_9689);
nor U10514 (N_10514,N_9001,N_9197);
or U10515 (N_10515,N_9579,N_9218);
nor U10516 (N_10516,N_9413,N_9545);
nand U10517 (N_10517,N_9733,N_9533);
and U10518 (N_10518,N_9762,N_9171);
nand U10519 (N_10519,N_9383,N_9479);
nand U10520 (N_10520,N_9942,N_9545);
or U10521 (N_10521,N_9120,N_9954);
and U10522 (N_10522,N_9509,N_9698);
and U10523 (N_10523,N_9137,N_9504);
nand U10524 (N_10524,N_9321,N_9392);
nand U10525 (N_10525,N_9073,N_9613);
nand U10526 (N_10526,N_9945,N_9841);
or U10527 (N_10527,N_9382,N_9839);
or U10528 (N_10528,N_9121,N_9910);
or U10529 (N_10529,N_9190,N_9620);
or U10530 (N_10530,N_9212,N_9352);
and U10531 (N_10531,N_9809,N_9039);
and U10532 (N_10532,N_9016,N_9508);
nor U10533 (N_10533,N_9517,N_9749);
nor U10534 (N_10534,N_9903,N_9942);
nor U10535 (N_10535,N_9514,N_9414);
and U10536 (N_10536,N_9776,N_9703);
nor U10537 (N_10537,N_9060,N_9413);
and U10538 (N_10538,N_9751,N_9718);
and U10539 (N_10539,N_9451,N_9762);
or U10540 (N_10540,N_9214,N_9088);
nor U10541 (N_10541,N_9263,N_9772);
and U10542 (N_10542,N_9499,N_9187);
nor U10543 (N_10543,N_9745,N_9947);
nand U10544 (N_10544,N_9063,N_9029);
or U10545 (N_10545,N_9621,N_9899);
or U10546 (N_10546,N_9591,N_9823);
nand U10547 (N_10547,N_9912,N_9237);
nand U10548 (N_10548,N_9348,N_9217);
nand U10549 (N_10549,N_9348,N_9396);
nand U10550 (N_10550,N_9056,N_9160);
nand U10551 (N_10551,N_9404,N_9386);
nand U10552 (N_10552,N_9427,N_9840);
nor U10553 (N_10553,N_9196,N_9016);
nor U10554 (N_10554,N_9704,N_9316);
nand U10555 (N_10555,N_9128,N_9294);
or U10556 (N_10556,N_9562,N_9522);
nand U10557 (N_10557,N_9042,N_9681);
and U10558 (N_10558,N_9705,N_9949);
or U10559 (N_10559,N_9076,N_9626);
and U10560 (N_10560,N_9362,N_9054);
or U10561 (N_10561,N_9193,N_9654);
nor U10562 (N_10562,N_9669,N_9746);
and U10563 (N_10563,N_9906,N_9904);
and U10564 (N_10564,N_9519,N_9362);
nor U10565 (N_10565,N_9167,N_9653);
or U10566 (N_10566,N_9382,N_9667);
or U10567 (N_10567,N_9266,N_9582);
nand U10568 (N_10568,N_9321,N_9991);
nand U10569 (N_10569,N_9462,N_9099);
or U10570 (N_10570,N_9527,N_9053);
or U10571 (N_10571,N_9651,N_9319);
or U10572 (N_10572,N_9759,N_9600);
nand U10573 (N_10573,N_9038,N_9683);
and U10574 (N_10574,N_9807,N_9954);
and U10575 (N_10575,N_9966,N_9169);
nand U10576 (N_10576,N_9757,N_9723);
or U10577 (N_10577,N_9683,N_9988);
and U10578 (N_10578,N_9407,N_9669);
and U10579 (N_10579,N_9698,N_9161);
or U10580 (N_10580,N_9311,N_9652);
and U10581 (N_10581,N_9851,N_9725);
and U10582 (N_10582,N_9074,N_9730);
and U10583 (N_10583,N_9957,N_9157);
nor U10584 (N_10584,N_9271,N_9628);
nor U10585 (N_10585,N_9992,N_9400);
nand U10586 (N_10586,N_9459,N_9984);
and U10587 (N_10587,N_9852,N_9104);
or U10588 (N_10588,N_9748,N_9184);
nand U10589 (N_10589,N_9592,N_9145);
and U10590 (N_10590,N_9572,N_9088);
or U10591 (N_10591,N_9848,N_9196);
nand U10592 (N_10592,N_9369,N_9082);
or U10593 (N_10593,N_9029,N_9702);
and U10594 (N_10594,N_9065,N_9273);
nor U10595 (N_10595,N_9255,N_9063);
nand U10596 (N_10596,N_9187,N_9803);
or U10597 (N_10597,N_9479,N_9411);
and U10598 (N_10598,N_9394,N_9198);
nor U10599 (N_10599,N_9321,N_9045);
nand U10600 (N_10600,N_9650,N_9285);
nand U10601 (N_10601,N_9968,N_9852);
or U10602 (N_10602,N_9745,N_9338);
nor U10603 (N_10603,N_9175,N_9394);
or U10604 (N_10604,N_9731,N_9873);
nor U10605 (N_10605,N_9518,N_9983);
nand U10606 (N_10606,N_9808,N_9290);
and U10607 (N_10607,N_9538,N_9833);
and U10608 (N_10608,N_9602,N_9515);
and U10609 (N_10609,N_9734,N_9519);
nor U10610 (N_10610,N_9286,N_9784);
nor U10611 (N_10611,N_9094,N_9645);
nor U10612 (N_10612,N_9769,N_9395);
nand U10613 (N_10613,N_9110,N_9495);
nand U10614 (N_10614,N_9056,N_9429);
nor U10615 (N_10615,N_9286,N_9807);
nor U10616 (N_10616,N_9930,N_9041);
nor U10617 (N_10617,N_9602,N_9060);
nand U10618 (N_10618,N_9966,N_9858);
nor U10619 (N_10619,N_9658,N_9469);
and U10620 (N_10620,N_9876,N_9328);
nor U10621 (N_10621,N_9176,N_9057);
nand U10622 (N_10622,N_9702,N_9103);
xnor U10623 (N_10623,N_9601,N_9346);
nand U10624 (N_10624,N_9304,N_9748);
nand U10625 (N_10625,N_9264,N_9973);
or U10626 (N_10626,N_9128,N_9530);
or U10627 (N_10627,N_9649,N_9140);
xnor U10628 (N_10628,N_9547,N_9650);
nor U10629 (N_10629,N_9572,N_9438);
and U10630 (N_10630,N_9924,N_9907);
nor U10631 (N_10631,N_9588,N_9943);
xnor U10632 (N_10632,N_9099,N_9020);
and U10633 (N_10633,N_9214,N_9631);
nand U10634 (N_10634,N_9507,N_9503);
and U10635 (N_10635,N_9896,N_9676);
nor U10636 (N_10636,N_9403,N_9145);
or U10637 (N_10637,N_9327,N_9368);
xnor U10638 (N_10638,N_9209,N_9142);
or U10639 (N_10639,N_9888,N_9608);
and U10640 (N_10640,N_9119,N_9548);
nor U10641 (N_10641,N_9560,N_9848);
or U10642 (N_10642,N_9703,N_9988);
nor U10643 (N_10643,N_9998,N_9761);
nand U10644 (N_10644,N_9243,N_9537);
or U10645 (N_10645,N_9667,N_9770);
nand U10646 (N_10646,N_9527,N_9570);
and U10647 (N_10647,N_9551,N_9199);
and U10648 (N_10648,N_9092,N_9635);
and U10649 (N_10649,N_9911,N_9249);
nand U10650 (N_10650,N_9403,N_9212);
xor U10651 (N_10651,N_9240,N_9019);
nor U10652 (N_10652,N_9777,N_9239);
or U10653 (N_10653,N_9241,N_9427);
nand U10654 (N_10654,N_9218,N_9061);
nor U10655 (N_10655,N_9462,N_9592);
nor U10656 (N_10656,N_9901,N_9510);
nor U10657 (N_10657,N_9132,N_9985);
or U10658 (N_10658,N_9097,N_9858);
nor U10659 (N_10659,N_9017,N_9011);
nor U10660 (N_10660,N_9474,N_9738);
and U10661 (N_10661,N_9453,N_9060);
and U10662 (N_10662,N_9786,N_9772);
nor U10663 (N_10663,N_9911,N_9623);
and U10664 (N_10664,N_9593,N_9849);
or U10665 (N_10665,N_9241,N_9117);
and U10666 (N_10666,N_9989,N_9700);
and U10667 (N_10667,N_9847,N_9199);
and U10668 (N_10668,N_9901,N_9861);
xnor U10669 (N_10669,N_9020,N_9090);
and U10670 (N_10670,N_9133,N_9374);
nor U10671 (N_10671,N_9481,N_9382);
and U10672 (N_10672,N_9576,N_9393);
nand U10673 (N_10673,N_9949,N_9445);
nand U10674 (N_10674,N_9580,N_9750);
nor U10675 (N_10675,N_9714,N_9716);
or U10676 (N_10676,N_9458,N_9191);
nand U10677 (N_10677,N_9495,N_9230);
nor U10678 (N_10678,N_9073,N_9021);
nor U10679 (N_10679,N_9493,N_9177);
or U10680 (N_10680,N_9140,N_9452);
nor U10681 (N_10681,N_9540,N_9791);
nor U10682 (N_10682,N_9658,N_9997);
and U10683 (N_10683,N_9989,N_9059);
nand U10684 (N_10684,N_9635,N_9877);
nor U10685 (N_10685,N_9339,N_9128);
and U10686 (N_10686,N_9149,N_9654);
nand U10687 (N_10687,N_9678,N_9483);
or U10688 (N_10688,N_9880,N_9941);
and U10689 (N_10689,N_9895,N_9458);
or U10690 (N_10690,N_9743,N_9898);
nor U10691 (N_10691,N_9402,N_9448);
nand U10692 (N_10692,N_9370,N_9111);
nor U10693 (N_10693,N_9229,N_9419);
or U10694 (N_10694,N_9980,N_9424);
or U10695 (N_10695,N_9731,N_9211);
and U10696 (N_10696,N_9702,N_9143);
and U10697 (N_10697,N_9320,N_9884);
and U10698 (N_10698,N_9300,N_9342);
and U10699 (N_10699,N_9696,N_9027);
and U10700 (N_10700,N_9122,N_9794);
nor U10701 (N_10701,N_9662,N_9388);
and U10702 (N_10702,N_9846,N_9579);
nand U10703 (N_10703,N_9469,N_9012);
and U10704 (N_10704,N_9840,N_9805);
nand U10705 (N_10705,N_9657,N_9223);
and U10706 (N_10706,N_9215,N_9076);
nand U10707 (N_10707,N_9501,N_9065);
nand U10708 (N_10708,N_9678,N_9397);
and U10709 (N_10709,N_9182,N_9393);
or U10710 (N_10710,N_9057,N_9469);
nor U10711 (N_10711,N_9668,N_9763);
or U10712 (N_10712,N_9110,N_9481);
nand U10713 (N_10713,N_9828,N_9751);
nand U10714 (N_10714,N_9084,N_9151);
nor U10715 (N_10715,N_9965,N_9321);
nor U10716 (N_10716,N_9863,N_9296);
nand U10717 (N_10717,N_9758,N_9720);
and U10718 (N_10718,N_9360,N_9600);
nor U10719 (N_10719,N_9240,N_9167);
nor U10720 (N_10720,N_9873,N_9517);
nor U10721 (N_10721,N_9701,N_9217);
or U10722 (N_10722,N_9292,N_9213);
and U10723 (N_10723,N_9170,N_9427);
nor U10724 (N_10724,N_9982,N_9345);
nor U10725 (N_10725,N_9500,N_9709);
nand U10726 (N_10726,N_9685,N_9655);
nor U10727 (N_10727,N_9313,N_9020);
nor U10728 (N_10728,N_9980,N_9104);
or U10729 (N_10729,N_9651,N_9111);
and U10730 (N_10730,N_9417,N_9464);
xor U10731 (N_10731,N_9973,N_9347);
nor U10732 (N_10732,N_9000,N_9577);
nor U10733 (N_10733,N_9209,N_9246);
nand U10734 (N_10734,N_9911,N_9682);
xor U10735 (N_10735,N_9420,N_9248);
xnor U10736 (N_10736,N_9358,N_9678);
and U10737 (N_10737,N_9631,N_9750);
and U10738 (N_10738,N_9664,N_9647);
nor U10739 (N_10739,N_9066,N_9763);
nand U10740 (N_10740,N_9377,N_9228);
nand U10741 (N_10741,N_9757,N_9828);
and U10742 (N_10742,N_9618,N_9710);
nand U10743 (N_10743,N_9199,N_9588);
nand U10744 (N_10744,N_9916,N_9082);
nor U10745 (N_10745,N_9360,N_9297);
and U10746 (N_10746,N_9567,N_9413);
and U10747 (N_10747,N_9923,N_9399);
and U10748 (N_10748,N_9231,N_9450);
nor U10749 (N_10749,N_9762,N_9650);
nor U10750 (N_10750,N_9541,N_9456);
and U10751 (N_10751,N_9655,N_9152);
or U10752 (N_10752,N_9603,N_9026);
and U10753 (N_10753,N_9914,N_9877);
and U10754 (N_10754,N_9130,N_9188);
and U10755 (N_10755,N_9127,N_9623);
and U10756 (N_10756,N_9692,N_9398);
or U10757 (N_10757,N_9051,N_9131);
nand U10758 (N_10758,N_9660,N_9394);
or U10759 (N_10759,N_9585,N_9101);
and U10760 (N_10760,N_9793,N_9320);
and U10761 (N_10761,N_9225,N_9322);
nor U10762 (N_10762,N_9768,N_9071);
nand U10763 (N_10763,N_9673,N_9396);
nor U10764 (N_10764,N_9893,N_9726);
nor U10765 (N_10765,N_9778,N_9081);
nand U10766 (N_10766,N_9989,N_9113);
or U10767 (N_10767,N_9038,N_9384);
and U10768 (N_10768,N_9643,N_9855);
nor U10769 (N_10769,N_9603,N_9014);
and U10770 (N_10770,N_9681,N_9174);
nor U10771 (N_10771,N_9217,N_9155);
nand U10772 (N_10772,N_9306,N_9587);
nand U10773 (N_10773,N_9721,N_9975);
nor U10774 (N_10774,N_9568,N_9655);
nor U10775 (N_10775,N_9458,N_9462);
nand U10776 (N_10776,N_9564,N_9789);
or U10777 (N_10777,N_9104,N_9256);
nand U10778 (N_10778,N_9697,N_9204);
and U10779 (N_10779,N_9845,N_9970);
nor U10780 (N_10780,N_9556,N_9221);
nor U10781 (N_10781,N_9983,N_9034);
nand U10782 (N_10782,N_9019,N_9586);
nand U10783 (N_10783,N_9252,N_9959);
nand U10784 (N_10784,N_9640,N_9986);
nor U10785 (N_10785,N_9705,N_9935);
nand U10786 (N_10786,N_9635,N_9475);
or U10787 (N_10787,N_9421,N_9487);
nand U10788 (N_10788,N_9724,N_9613);
nand U10789 (N_10789,N_9342,N_9997);
nand U10790 (N_10790,N_9888,N_9881);
nor U10791 (N_10791,N_9375,N_9356);
or U10792 (N_10792,N_9115,N_9748);
or U10793 (N_10793,N_9238,N_9723);
nor U10794 (N_10794,N_9629,N_9676);
nand U10795 (N_10795,N_9058,N_9237);
nor U10796 (N_10796,N_9940,N_9674);
nand U10797 (N_10797,N_9346,N_9132);
xor U10798 (N_10798,N_9948,N_9574);
nand U10799 (N_10799,N_9377,N_9513);
nand U10800 (N_10800,N_9453,N_9969);
or U10801 (N_10801,N_9079,N_9298);
nor U10802 (N_10802,N_9904,N_9887);
nor U10803 (N_10803,N_9562,N_9219);
or U10804 (N_10804,N_9913,N_9878);
nor U10805 (N_10805,N_9354,N_9708);
nor U10806 (N_10806,N_9855,N_9809);
and U10807 (N_10807,N_9611,N_9490);
nand U10808 (N_10808,N_9320,N_9207);
nor U10809 (N_10809,N_9679,N_9046);
or U10810 (N_10810,N_9942,N_9298);
or U10811 (N_10811,N_9538,N_9088);
nor U10812 (N_10812,N_9762,N_9140);
and U10813 (N_10813,N_9621,N_9507);
or U10814 (N_10814,N_9850,N_9023);
xor U10815 (N_10815,N_9195,N_9979);
nor U10816 (N_10816,N_9599,N_9218);
nand U10817 (N_10817,N_9203,N_9043);
and U10818 (N_10818,N_9162,N_9202);
and U10819 (N_10819,N_9694,N_9492);
and U10820 (N_10820,N_9710,N_9976);
nand U10821 (N_10821,N_9334,N_9744);
nand U10822 (N_10822,N_9339,N_9711);
nor U10823 (N_10823,N_9974,N_9269);
and U10824 (N_10824,N_9920,N_9331);
nand U10825 (N_10825,N_9476,N_9601);
nand U10826 (N_10826,N_9937,N_9095);
or U10827 (N_10827,N_9803,N_9920);
nor U10828 (N_10828,N_9850,N_9780);
and U10829 (N_10829,N_9294,N_9689);
or U10830 (N_10830,N_9702,N_9111);
nand U10831 (N_10831,N_9534,N_9233);
or U10832 (N_10832,N_9554,N_9019);
nor U10833 (N_10833,N_9923,N_9024);
or U10834 (N_10834,N_9136,N_9649);
and U10835 (N_10835,N_9990,N_9832);
nor U10836 (N_10836,N_9560,N_9921);
nand U10837 (N_10837,N_9331,N_9339);
nor U10838 (N_10838,N_9286,N_9580);
or U10839 (N_10839,N_9469,N_9008);
nor U10840 (N_10840,N_9522,N_9929);
nand U10841 (N_10841,N_9114,N_9115);
and U10842 (N_10842,N_9225,N_9645);
xnor U10843 (N_10843,N_9147,N_9105);
nand U10844 (N_10844,N_9911,N_9987);
and U10845 (N_10845,N_9297,N_9549);
and U10846 (N_10846,N_9810,N_9092);
nor U10847 (N_10847,N_9969,N_9622);
and U10848 (N_10848,N_9413,N_9435);
nand U10849 (N_10849,N_9059,N_9364);
nor U10850 (N_10850,N_9226,N_9625);
xnor U10851 (N_10851,N_9691,N_9964);
nor U10852 (N_10852,N_9950,N_9231);
and U10853 (N_10853,N_9232,N_9168);
nor U10854 (N_10854,N_9896,N_9993);
and U10855 (N_10855,N_9634,N_9517);
nand U10856 (N_10856,N_9507,N_9106);
nor U10857 (N_10857,N_9315,N_9861);
or U10858 (N_10858,N_9918,N_9032);
nor U10859 (N_10859,N_9064,N_9153);
nor U10860 (N_10860,N_9801,N_9010);
or U10861 (N_10861,N_9561,N_9528);
and U10862 (N_10862,N_9723,N_9008);
nand U10863 (N_10863,N_9224,N_9362);
nor U10864 (N_10864,N_9858,N_9546);
nor U10865 (N_10865,N_9421,N_9469);
and U10866 (N_10866,N_9892,N_9113);
nand U10867 (N_10867,N_9897,N_9545);
and U10868 (N_10868,N_9568,N_9038);
or U10869 (N_10869,N_9481,N_9364);
or U10870 (N_10870,N_9243,N_9601);
nor U10871 (N_10871,N_9618,N_9505);
or U10872 (N_10872,N_9320,N_9984);
or U10873 (N_10873,N_9684,N_9123);
or U10874 (N_10874,N_9560,N_9631);
or U10875 (N_10875,N_9306,N_9927);
or U10876 (N_10876,N_9381,N_9130);
or U10877 (N_10877,N_9603,N_9223);
or U10878 (N_10878,N_9987,N_9660);
nand U10879 (N_10879,N_9184,N_9964);
nor U10880 (N_10880,N_9479,N_9184);
and U10881 (N_10881,N_9651,N_9658);
nand U10882 (N_10882,N_9507,N_9481);
or U10883 (N_10883,N_9975,N_9994);
and U10884 (N_10884,N_9165,N_9341);
and U10885 (N_10885,N_9185,N_9822);
nand U10886 (N_10886,N_9912,N_9884);
nand U10887 (N_10887,N_9689,N_9008);
nor U10888 (N_10888,N_9196,N_9137);
nand U10889 (N_10889,N_9855,N_9896);
nor U10890 (N_10890,N_9446,N_9357);
nand U10891 (N_10891,N_9474,N_9100);
nand U10892 (N_10892,N_9614,N_9054);
and U10893 (N_10893,N_9801,N_9490);
nand U10894 (N_10894,N_9683,N_9270);
nand U10895 (N_10895,N_9497,N_9785);
nand U10896 (N_10896,N_9018,N_9117);
and U10897 (N_10897,N_9345,N_9915);
and U10898 (N_10898,N_9750,N_9841);
or U10899 (N_10899,N_9722,N_9503);
nand U10900 (N_10900,N_9831,N_9057);
nor U10901 (N_10901,N_9648,N_9288);
nor U10902 (N_10902,N_9041,N_9671);
and U10903 (N_10903,N_9026,N_9501);
or U10904 (N_10904,N_9460,N_9501);
and U10905 (N_10905,N_9497,N_9208);
nor U10906 (N_10906,N_9102,N_9743);
nand U10907 (N_10907,N_9243,N_9541);
or U10908 (N_10908,N_9032,N_9707);
or U10909 (N_10909,N_9732,N_9796);
and U10910 (N_10910,N_9015,N_9316);
nand U10911 (N_10911,N_9886,N_9646);
nor U10912 (N_10912,N_9348,N_9554);
nand U10913 (N_10913,N_9027,N_9665);
or U10914 (N_10914,N_9662,N_9275);
nand U10915 (N_10915,N_9126,N_9636);
and U10916 (N_10916,N_9473,N_9594);
or U10917 (N_10917,N_9766,N_9905);
and U10918 (N_10918,N_9782,N_9944);
and U10919 (N_10919,N_9258,N_9923);
and U10920 (N_10920,N_9471,N_9650);
and U10921 (N_10921,N_9149,N_9426);
nand U10922 (N_10922,N_9952,N_9315);
and U10923 (N_10923,N_9340,N_9066);
or U10924 (N_10924,N_9381,N_9345);
nor U10925 (N_10925,N_9182,N_9117);
or U10926 (N_10926,N_9327,N_9828);
and U10927 (N_10927,N_9166,N_9576);
or U10928 (N_10928,N_9197,N_9042);
or U10929 (N_10929,N_9163,N_9754);
nand U10930 (N_10930,N_9698,N_9164);
nor U10931 (N_10931,N_9197,N_9048);
nor U10932 (N_10932,N_9438,N_9984);
nor U10933 (N_10933,N_9352,N_9013);
nor U10934 (N_10934,N_9020,N_9241);
nor U10935 (N_10935,N_9164,N_9811);
or U10936 (N_10936,N_9222,N_9584);
and U10937 (N_10937,N_9654,N_9726);
nand U10938 (N_10938,N_9158,N_9828);
or U10939 (N_10939,N_9923,N_9537);
or U10940 (N_10940,N_9513,N_9770);
or U10941 (N_10941,N_9291,N_9304);
nand U10942 (N_10942,N_9788,N_9042);
or U10943 (N_10943,N_9875,N_9131);
nor U10944 (N_10944,N_9740,N_9987);
and U10945 (N_10945,N_9340,N_9130);
or U10946 (N_10946,N_9140,N_9201);
nand U10947 (N_10947,N_9670,N_9297);
nor U10948 (N_10948,N_9946,N_9745);
nand U10949 (N_10949,N_9271,N_9598);
nand U10950 (N_10950,N_9994,N_9657);
and U10951 (N_10951,N_9670,N_9004);
nor U10952 (N_10952,N_9997,N_9430);
nor U10953 (N_10953,N_9792,N_9562);
nor U10954 (N_10954,N_9911,N_9566);
nor U10955 (N_10955,N_9230,N_9886);
or U10956 (N_10956,N_9180,N_9771);
or U10957 (N_10957,N_9849,N_9398);
nor U10958 (N_10958,N_9339,N_9682);
nor U10959 (N_10959,N_9476,N_9013);
and U10960 (N_10960,N_9470,N_9140);
nor U10961 (N_10961,N_9989,N_9798);
and U10962 (N_10962,N_9556,N_9247);
or U10963 (N_10963,N_9213,N_9921);
and U10964 (N_10964,N_9113,N_9567);
or U10965 (N_10965,N_9255,N_9799);
nand U10966 (N_10966,N_9372,N_9766);
nor U10967 (N_10967,N_9079,N_9536);
and U10968 (N_10968,N_9796,N_9937);
nor U10969 (N_10969,N_9304,N_9641);
and U10970 (N_10970,N_9077,N_9422);
and U10971 (N_10971,N_9912,N_9110);
nor U10972 (N_10972,N_9641,N_9905);
nand U10973 (N_10973,N_9089,N_9088);
and U10974 (N_10974,N_9711,N_9822);
or U10975 (N_10975,N_9953,N_9889);
and U10976 (N_10976,N_9809,N_9754);
nand U10977 (N_10977,N_9977,N_9267);
or U10978 (N_10978,N_9292,N_9826);
and U10979 (N_10979,N_9239,N_9513);
or U10980 (N_10980,N_9710,N_9218);
or U10981 (N_10981,N_9515,N_9544);
nor U10982 (N_10982,N_9901,N_9190);
and U10983 (N_10983,N_9827,N_9527);
and U10984 (N_10984,N_9108,N_9795);
nor U10985 (N_10985,N_9144,N_9190);
or U10986 (N_10986,N_9246,N_9135);
nor U10987 (N_10987,N_9459,N_9856);
nor U10988 (N_10988,N_9415,N_9399);
nand U10989 (N_10989,N_9075,N_9058);
nand U10990 (N_10990,N_9410,N_9196);
nand U10991 (N_10991,N_9890,N_9265);
nor U10992 (N_10992,N_9131,N_9279);
nor U10993 (N_10993,N_9445,N_9468);
or U10994 (N_10994,N_9745,N_9573);
xnor U10995 (N_10995,N_9803,N_9854);
or U10996 (N_10996,N_9574,N_9497);
and U10997 (N_10997,N_9846,N_9092);
nand U10998 (N_10998,N_9493,N_9454);
xnor U10999 (N_10999,N_9488,N_9491);
and U11000 (N_11000,N_10425,N_10929);
or U11001 (N_11001,N_10277,N_10309);
nand U11002 (N_11002,N_10751,N_10257);
nand U11003 (N_11003,N_10680,N_10305);
nand U11004 (N_11004,N_10820,N_10593);
nor U11005 (N_11005,N_10823,N_10069);
or U11006 (N_11006,N_10448,N_10082);
or U11007 (N_11007,N_10832,N_10387);
or U11008 (N_11008,N_10895,N_10958);
and U11009 (N_11009,N_10123,N_10652);
or U11010 (N_11010,N_10273,N_10172);
nand U11011 (N_11011,N_10466,N_10226);
nor U11012 (N_11012,N_10383,N_10406);
and U11013 (N_11013,N_10570,N_10013);
nand U11014 (N_11014,N_10645,N_10436);
and U11015 (N_11015,N_10946,N_10221);
nand U11016 (N_11016,N_10312,N_10608);
nor U11017 (N_11017,N_10026,N_10083);
nor U11018 (N_11018,N_10749,N_10396);
nand U11019 (N_11019,N_10010,N_10977);
nor U11020 (N_11020,N_10419,N_10216);
and U11021 (N_11021,N_10214,N_10508);
or U11022 (N_11022,N_10354,N_10066);
and U11023 (N_11023,N_10871,N_10594);
nand U11024 (N_11024,N_10367,N_10587);
nor U11025 (N_11025,N_10036,N_10971);
or U11026 (N_11026,N_10404,N_10099);
nand U11027 (N_11027,N_10524,N_10317);
nand U11028 (N_11028,N_10428,N_10442);
and U11029 (N_11029,N_10539,N_10073);
or U11030 (N_11030,N_10794,N_10389);
nand U11031 (N_11031,N_10759,N_10825);
nand U11032 (N_11032,N_10999,N_10154);
or U11033 (N_11033,N_10050,N_10950);
or U11034 (N_11034,N_10515,N_10654);
nor U11035 (N_11035,N_10206,N_10330);
nand U11036 (N_11036,N_10027,N_10502);
and U11037 (N_11037,N_10271,N_10527);
and U11038 (N_11038,N_10045,N_10709);
or U11039 (N_11039,N_10876,N_10571);
nand U11040 (N_11040,N_10056,N_10243);
or U11041 (N_11041,N_10705,N_10846);
nor U11042 (N_11042,N_10266,N_10673);
nor U11043 (N_11043,N_10995,N_10016);
nor U11044 (N_11044,N_10969,N_10345);
nor U11045 (N_11045,N_10880,N_10166);
nor U11046 (N_11046,N_10248,N_10219);
nor U11047 (N_11047,N_10694,N_10476);
nor U11048 (N_11048,N_10774,N_10504);
nand U11049 (N_11049,N_10197,N_10132);
nand U11050 (N_11050,N_10331,N_10105);
or U11051 (N_11051,N_10429,N_10440);
or U11052 (N_11052,N_10636,N_10807);
and U11053 (N_11053,N_10110,N_10019);
or U11054 (N_11054,N_10778,N_10664);
or U11055 (N_11055,N_10981,N_10472);
nand U11056 (N_11056,N_10042,N_10230);
and U11057 (N_11057,N_10407,N_10638);
nand U11058 (N_11058,N_10282,N_10731);
or U11059 (N_11059,N_10691,N_10304);
nor U11060 (N_11060,N_10937,N_10015);
and U11061 (N_11061,N_10746,N_10438);
and U11062 (N_11062,N_10585,N_10366);
nand U11063 (N_11063,N_10382,N_10677);
nor U11064 (N_11064,N_10355,N_10433);
nand U11065 (N_11065,N_10810,N_10191);
nand U11066 (N_11066,N_10421,N_10058);
nor U11067 (N_11067,N_10035,N_10919);
or U11068 (N_11068,N_10564,N_10048);
or U11069 (N_11069,N_10333,N_10402);
and U11070 (N_11070,N_10097,N_10588);
nand U11071 (N_11071,N_10041,N_10475);
or U11072 (N_11072,N_10306,N_10431);
and U11073 (N_11073,N_10684,N_10343);
nand U11074 (N_11074,N_10454,N_10102);
or U11075 (N_11075,N_10095,N_10228);
nand U11076 (N_11076,N_10573,N_10894);
or U11077 (N_11077,N_10557,N_10905);
nand U11078 (N_11078,N_10827,N_10093);
nand U11079 (N_11079,N_10193,N_10092);
or U11080 (N_11080,N_10081,N_10992);
and U11081 (N_11081,N_10457,N_10761);
and U11082 (N_11082,N_10922,N_10898);
nand U11083 (N_11083,N_10857,N_10190);
or U11084 (N_11084,N_10183,N_10967);
nor U11085 (N_11085,N_10822,N_10965);
nor U11086 (N_11086,N_10443,N_10264);
nor U11087 (N_11087,N_10000,N_10662);
nor U11088 (N_11088,N_10916,N_10757);
and U11089 (N_11089,N_10234,N_10043);
and U11090 (N_11090,N_10959,N_10004);
nor U11091 (N_11091,N_10742,N_10784);
nor U11092 (N_11092,N_10704,N_10499);
and U11093 (N_11093,N_10868,N_10314);
and U11094 (N_11094,N_10113,N_10427);
and U11095 (N_11095,N_10743,N_10416);
and U11096 (N_11096,N_10802,N_10061);
and U11097 (N_11097,N_10131,N_10915);
or U11098 (N_11098,N_10816,N_10686);
or U11099 (N_11099,N_10773,N_10633);
nor U11100 (N_11100,N_10543,N_10459);
and U11101 (N_11101,N_10115,N_10232);
nor U11102 (N_11102,N_10414,N_10768);
nand U11103 (N_11103,N_10982,N_10644);
nand U11104 (N_11104,N_10639,N_10159);
nor U11105 (N_11105,N_10853,N_10568);
nand U11106 (N_11106,N_10521,N_10405);
nand U11107 (N_11107,N_10994,N_10783);
nor U11108 (N_11108,N_10575,N_10213);
nor U11109 (N_11109,N_10562,N_10702);
nor U11110 (N_11110,N_10386,N_10390);
nand U11111 (N_11111,N_10149,N_10653);
nor U11112 (N_11112,N_10323,N_10065);
nor U11113 (N_11113,N_10201,N_10837);
nor U11114 (N_11114,N_10711,N_10690);
or U11115 (N_11115,N_10031,N_10423);
nand U11116 (N_11116,N_10782,N_10998);
nand U11117 (N_11117,N_10723,N_10186);
xor U11118 (N_11118,N_10302,N_10514);
nand U11119 (N_11119,N_10618,N_10077);
or U11120 (N_11120,N_10603,N_10732);
nand U11121 (N_11121,N_10252,N_10523);
nand U11122 (N_11122,N_10362,N_10260);
and U11123 (N_11123,N_10579,N_10801);
and U11124 (N_11124,N_10787,N_10493);
nor U11125 (N_11125,N_10556,N_10391);
or U11126 (N_11126,N_10849,N_10393);
and U11127 (N_11127,N_10621,N_10484);
nor U11128 (N_11128,N_10003,N_10326);
nand U11129 (N_11129,N_10296,N_10430);
nor U11130 (N_11130,N_10278,N_10545);
or U11131 (N_11131,N_10780,N_10974);
or U11132 (N_11132,N_10164,N_10175);
nand U11133 (N_11133,N_10225,N_10688);
xnor U11134 (N_11134,N_10991,N_10954);
nor U11135 (N_11135,N_10920,N_10318);
nor U11136 (N_11136,N_10046,N_10879);
nor U11137 (N_11137,N_10675,N_10637);
nand U11138 (N_11138,N_10152,N_10829);
or U11139 (N_11139,N_10174,N_10265);
or U11140 (N_11140,N_10291,N_10032);
nor U11141 (N_11141,N_10119,N_10666);
nor U11142 (N_11142,N_10388,N_10049);
nand U11143 (N_11143,N_10805,N_10187);
xor U11144 (N_11144,N_10712,N_10057);
and U11145 (N_11145,N_10755,N_10384);
or U11146 (N_11146,N_10199,N_10855);
nand U11147 (N_11147,N_10486,N_10926);
or U11148 (N_11148,N_10566,N_10841);
and U11149 (N_11149,N_10506,N_10250);
nand U11150 (N_11150,N_10833,N_10192);
and U11151 (N_11151,N_10669,N_10939);
or U11152 (N_11152,N_10434,N_10553);
nor U11153 (N_11153,N_10750,N_10215);
nor U11154 (N_11154,N_10945,N_10426);
nand U11155 (N_11155,N_10329,N_10394);
nor U11156 (N_11156,N_10660,N_10874);
or U11157 (N_11157,N_10293,N_10203);
nand U11158 (N_11158,N_10128,N_10311);
or U11159 (N_11159,N_10209,N_10490);
nor U11160 (N_11160,N_10933,N_10964);
nand U11161 (N_11161,N_10733,N_10944);
and U11162 (N_11162,N_10520,N_10699);
nor U11163 (N_11163,N_10210,N_10068);
nor U11164 (N_11164,N_10158,N_10589);
nand U11165 (N_11165,N_10665,N_10717);
or U11166 (N_11166,N_10301,N_10947);
nand U11167 (N_11167,N_10075,N_10104);
and U11168 (N_11168,N_10903,N_10904);
nand U11169 (N_11169,N_10772,N_10245);
nor U11170 (N_11170,N_10814,N_10489);
and U11171 (N_11171,N_10600,N_10285);
nand U11172 (N_11172,N_10581,N_10361);
or U11173 (N_11173,N_10283,N_10925);
nor U11174 (N_11174,N_10351,N_10526);
or U11175 (N_11175,N_10308,N_10558);
nor U11176 (N_11176,N_10718,N_10830);
or U11177 (N_11177,N_10122,N_10622);
xnor U11178 (N_11178,N_10635,N_10655);
nand U11179 (N_11179,N_10125,N_10909);
or U11180 (N_11180,N_10497,N_10332);
or U11181 (N_11181,N_10307,N_10327);
nand U11182 (N_11182,N_10085,N_10471);
or U11183 (N_11183,N_10349,N_10021);
and U11184 (N_11184,N_10927,N_10029);
nor U11185 (N_11185,N_10348,N_10646);
or U11186 (N_11186,N_10107,N_10697);
nand U11187 (N_11187,N_10628,N_10978);
nand U11188 (N_11188,N_10181,N_10074);
or U11189 (N_11189,N_10725,N_10184);
nor U11190 (N_11190,N_10151,N_10340);
and U11191 (N_11191,N_10202,N_10873);
and U11192 (N_11192,N_10272,N_10500);
nand U11193 (N_11193,N_10747,N_10530);
or U11194 (N_11194,N_10313,N_10888);
nor U11195 (N_11195,N_10576,N_10990);
nor U11196 (N_11196,N_10398,N_10133);
nor U11197 (N_11197,N_10872,N_10844);
nor U11198 (N_11198,N_10692,N_10851);
nand U11199 (N_11199,N_10739,N_10465);
nor U11200 (N_11200,N_10336,N_10033);
or U11201 (N_11201,N_10987,N_10403);
nand U11202 (N_11202,N_10949,N_10578);
nand U11203 (N_11203,N_10094,N_10136);
and U11204 (N_11204,N_10790,N_10258);
or U11205 (N_11205,N_10605,N_10613);
nand U11206 (N_11206,N_10224,N_10847);
or U11207 (N_11207,N_10509,N_10631);
and U11208 (N_11208,N_10634,N_10617);
or U11209 (N_11209,N_10240,N_10063);
xor U11210 (N_11210,N_10494,N_10452);
nor U11211 (N_11211,N_10522,N_10217);
or U11212 (N_11212,N_10775,N_10337);
nand U11213 (N_11213,N_10208,N_10900);
nand U11214 (N_11214,N_10720,N_10678);
and U11215 (N_11215,N_10072,N_10834);
and U11216 (N_11216,N_10098,N_10059);
or U11217 (N_11217,N_10795,N_10713);
nor U11218 (N_11218,N_10207,N_10116);
nor U11219 (N_11219,N_10357,N_10339);
and U11220 (N_11220,N_10547,N_10862);
nand U11221 (N_11221,N_10346,N_10111);
and U11222 (N_11222,N_10037,N_10195);
or U11223 (N_11223,N_10320,N_10651);
and U11224 (N_11224,N_10267,N_10319);
and U11225 (N_11225,N_10194,N_10657);
or U11226 (N_11226,N_10086,N_10134);
xnor U11227 (N_11227,N_10567,N_10860);
or U11228 (N_11228,N_10884,N_10610);
and U11229 (N_11229,N_10812,N_10084);
nand U11230 (N_11230,N_10112,N_10650);
nor U11231 (N_11231,N_10124,N_10445);
nor U11232 (N_11232,N_10663,N_10024);
or U11233 (N_11233,N_10381,N_10079);
or U11234 (N_11234,N_10117,N_10815);
and U11235 (N_11235,N_10565,N_10932);
or U11236 (N_11236,N_10769,N_10292);
or U11237 (N_11237,N_10413,N_10276);
and U11238 (N_11238,N_10754,N_10441);
nand U11239 (N_11239,N_10231,N_10512);
or U11240 (N_11240,N_10185,N_10218);
nand U11241 (N_11241,N_10917,N_10334);
nand U11242 (N_11242,N_10546,N_10253);
or U11243 (N_11243,N_10196,N_10598);
or U11244 (N_11244,N_10410,N_10885);
or U11245 (N_11245,N_10719,N_10563);
and U11246 (N_11246,N_10912,N_10931);
nor U11247 (N_11247,N_10316,N_10420);
or U11248 (N_11248,N_10352,N_10039);
and U11249 (N_11249,N_10765,N_10979);
or U11250 (N_11250,N_10785,N_10627);
nand U11251 (N_11251,N_10776,N_10344);
or U11252 (N_11252,N_10474,N_10503);
and U11253 (N_11253,N_10656,N_10062);
nand U11254 (N_11254,N_10511,N_10325);
nand U11255 (N_11255,N_10242,N_10800);
or U11256 (N_11256,N_10997,N_10055);
or U11257 (N_11257,N_10649,N_10268);
nor U11258 (N_11258,N_10461,N_10890);
nor U11259 (N_11259,N_10941,N_10752);
nor U11260 (N_11260,N_10850,N_10411);
nand U11261 (N_11261,N_10590,N_10706);
or U11262 (N_11262,N_10727,N_10087);
or U11263 (N_11263,N_10896,N_10241);
and U11264 (N_11264,N_10447,N_10446);
nand U11265 (N_11265,N_10624,N_10714);
or U11266 (N_11266,N_10288,N_10412);
nor U11267 (N_11267,N_10030,N_10060);
or U11268 (N_11268,N_10993,N_10014);
nand U11269 (N_11269,N_10818,N_10914);
nand U11270 (N_11270,N_10940,N_10467);
and U11271 (N_11271,N_10685,N_10477);
nor U11272 (N_11272,N_10744,N_10683);
and U11273 (N_11273,N_10821,N_10372);
and U11274 (N_11274,N_10843,N_10067);
nor U11275 (N_11275,N_10806,N_10321);
nor U11276 (N_11276,N_10803,N_10948);
or U11277 (N_11277,N_10487,N_10517);
or U11278 (N_11278,N_10882,N_10147);
and U11279 (N_11279,N_10145,N_10659);
and U11280 (N_11280,N_10179,N_10473);
or U11281 (N_11281,N_10962,N_10549);
nand U11282 (N_11282,N_10672,N_10369);
and U11283 (N_11283,N_10458,N_10040);
nor U11284 (N_11284,N_10148,N_10485);
nand U11285 (N_11285,N_10642,N_10350);
nand U11286 (N_11286,N_10729,N_10342);
and U11287 (N_11287,N_10583,N_10237);
or U11288 (N_11288,N_10163,N_10938);
nor U11289 (N_11289,N_10848,N_10020);
nor U11290 (N_11290,N_10592,N_10178);
nand U11291 (N_11291,N_10364,N_10956);
or U11292 (N_11292,N_10138,N_10828);
or U11293 (N_11293,N_10771,N_10619);
and U11294 (N_11294,N_10137,N_10541);
nand U11295 (N_11295,N_10670,N_10096);
nand U11296 (N_11296,N_10943,N_10510);
nor U11297 (N_11297,N_10883,N_10470);
xnor U11298 (N_11298,N_10797,N_10298);
and U11299 (N_11299,N_10375,N_10923);
nor U11300 (N_11300,N_10373,N_10501);
or U11301 (N_11301,N_10047,N_10409);
nor U11302 (N_11302,N_10574,N_10865);
and U11303 (N_11303,N_10518,N_10781);
and U11304 (N_11304,N_10824,N_10715);
or U11305 (N_11305,N_10599,N_10255);
and U11306 (N_11306,N_10881,N_10328);
or U11307 (N_11307,N_10435,N_10831);
and U11308 (N_11308,N_10701,N_10295);
or U11309 (N_11309,N_10845,N_10052);
nor U11310 (N_11310,N_10363,N_10368);
or U11311 (N_11311,N_10798,N_10970);
nand U11312 (N_11312,N_10756,N_10341);
nor U11313 (N_11313,N_10985,N_10239);
and U11314 (N_11314,N_10989,N_10170);
nor U11315 (N_11315,N_10616,N_10141);
nand U11316 (N_11316,N_10674,N_10643);
nand U11317 (N_11317,N_10380,N_10463);
and U11318 (N_11318,N_10211,N_10017);
or U11319 (N_11319,N_10988,N_10222);
or U11320 (N_11320,N_10893,N_10205);
nor U11321 (N_11321,N_10089,N_10469);
or U11322 (N_11322,N_10960,N_10764);
and U11323 (N_11323,N_10708,N_10836);
or U11324 (N_11324,N_10495,N_10840);
and U11325 (N_11325,N_10819,N_10233);
and U11326 (N_11326,N_10813,N_10235);
or U11327 (N_11327,N_10548,N_10401);
nand U11328 (N_11328,N_10177,N_10569);
and U11329 (N_11329,N_10921,N_10281);
nor U11330 (N_11330,N_10127,N_10753);
or U11331 (N_11331,N_10299,N_10101);
and U11332 (N_11332,N_10360,N_10051);
and U11333 (N_11333,N_10609,N_10005);
or U11334 (N_11334,N_10864,N_10737);
and U11335 (N_11335,N_10863,N_10748);
or U11336 (N_11336,N_10424,N_10934);
and U11337 (N_11337,N_10130,N_10379);
or U11338 (N_11338,N_10952,N_10607);
and U11339 (N_11339,N_10290,N_10796);
or U11340 (N_11340,N_10595,N_10724);
nand U11341 (N_11341,N_10577,N_10262);
nor U11342 (N_11342,N_10601,N_10176);
nand U11343 (N_11343,N_10906,N_10745);
and U11344 (N_11344,N_10852,N_10076);
nor U11345 (N_11345,N_10826,N_10513);
and U11346 (N_11346,N_10156,N_10220);
nand U11347 (N_11347,N_10418,N_10399);
and U11348 (N_11348,N_10973,N_10996);
and U11349 (N_11349,N_10165,N_10584);
nand U11350 (N_11350,N_10162,N_10012);
nor U11351 (N_11351,N_10707,N_10189);
and U11352 (N_11352,N_10687,N_10786);
or U11353 (N_11353,N_10070,N_10335);
and U11354 (N_11354,N_10789,N_10682);
or U11355 (N_11355,N_10792,N_10908);
nand U11356 (N_11356,N_10018,N_10365);
and U11357 (N_11357,N_10910,N_10450);
and U11358 (N_11358,N_10171,N_10247);
and U11359 (N_11359,N_10735,N_10377);
nor U11360 (N_11360,N_10359,N_10038);
and U11361 (N_11361,N_10808,N_10155);
nor U11362 (N_11362,N_10198,N_10641);
and U11363 (N_11363,N_10263,N_10693);
or U11364 (N_11364,N_10779,N_10322);
nor U11365 (N_11365,N_10839,N_10550);
and U11366 (N_11366,N_10835,N_10280);
nor U11367 (N_11367,N_10953,N_10294);
or U11368 (N_11368,N_10400,N_10054);
or U11369 (N_11369,N_10227,N_10432);
nor U11370 (N_11370,N_10975,N_10212);
nor U11371 (N_11371,N_10626,N_10173);
nand U11372 (N_11372,N_10561,N_10555);
nand U11373 (N_11373,N_10544,N_10870);
nand U11374 (N_11374,N_10417,N_10867);
and U11375 (N_11375,N_10611,N_10453);
nor U11376 (N_11376,N_10274,N_10942);
or U11377 (N_11377,N_10736,N_10090);
nor U11378 (N_11378,N_10572,N_10261);
or U11379 (N_11379,N_10488,N_10415);
or U11380 (N_11380,N_10728,N_10540);
nand U11381 (N_11381,N_10236,N_10044);
and U11382 (N_11382,N_10606,N_10385);
nand U11383 (N_11383,N_10150,N_10586);
nor U11384 (N_11384,N_10703,N_10793);
nand U11385 (N_11385,N_10891,N_10596);
or U11386 (N_11386,N_10554,N_10951);
or U11387 (N_11387,N_10455,N_10482);
or U11388 (N_11388,N_10632,N_10002);
and U11389 (N_11389,N_10114,N_10249);
nand U11390 (N_11390,N_10439,N_10135);
nor U11391 (N_11391,N_10877,N_10552);
nand U11392 (N_11392,N_10791,N_10028);
or U11393 (N_11393,N_10408,N_10788);
nand U11394 (N_11394,N_10300,N_10740);
nand U11395 (N_11395,N_10961,N_10696);
nor U11396 (N_11396,N_10286,N_10315);
or U11397 (N_11397,N_10244,N_10287);
nand U11398 (N_11398,N_10139,N_10491);
nor U11399 (N_11399,N_10809,N_10804);
nand U11400 (N_11400,N_10551,N_10532);
and U11401 (N_11401,N_10758,N_10395);
nand U11402 (N_11402,N_10620,N_10188);
nor U11403 (N_11403,N_10721,N_10918);
and U11404 (N_11404,N_10126,N_10615);
nor U11405 (N_11405,N_10935,N_10143);
nor U11406 (N_11406,N_10695,N_10770);
or U11407 (N_11407,N_10538,N_10861);
and U11408 (N_11408,N_10121,N_10422);
and U11409 (N_11409,N_10913,N_10525);
and U11410 (N_11410,N_10930,N_10007);
or U11411 (N_11411,N_10681,N_10106);
nand U11412 (N_11412,N_10980,N_10338);
and U11413 (N_11413,N_10760,N_10505);
and U11414 (N_11414,N_10397,N_10460);
nand U11415 (N_11415,N_10902,N_10279);
and U11416 (N_11416,N_10025,N_10671);
and U11417 (N_11417,N_10256,N_10580);
nor U11418 (N_11418,N_10088,N_10023);
nand U11419 (N_11419,N_10766,N_10928);
nand U11420 (N_11420,N_10738,N_10534);
or U11421 (N_11421,N_10668,N_10464);
nand U11422 (N_11422,N_10180,N_10071);
nand U11423 (N_11423,N_10838,N_10392);
nand U11424 (N_11424,N_10378,N_10109);
nor U11425 (N_11425,N_10957,N_10437);
nand U11426 (N_11426,N_10667,N_10859);
or U11427 (N_11427,N_10182,N_10034);
nor U11428 (N_11428,N_10661,N_10936);
nand U11429 (N_11429,N_10591,N_10972);
nor U11430 (N_11430,N_10444,N_10456);
nor U11431 (N_11431,N_10648,N_10157);
or U11432 (N_11432,N_10889,N_10080);
or U11433 (N_11433,N_10078,N_10966);
and U11434 (N_11434,N_10623,N_10011);
nand U11435 (N_11435,N_10371,N_10238);
xnor U11436 (N_11436,N_10899,N_10542);
or U11437 (N_11437,N_10963,N_10376);
and U11438 (N_11438,N_10767,N_10842);
nand U11439 (N_11439,N_10516,N_10100);
or U11440 (N_11440,N_10146,N_10854);
and U11441 (N_11441,N_10144,N_10533);
nor U11442 (N_11442,N_10161,N_10223);
nor U11443 (N_11443,N_10478,N_10856);
nor U11444 (N_11444,N_10142,N_10531);
or U11445 (N_11445,N_10878,N_10480);
or U11446 (N_11446,N_10604,N_10289);
or U11447 (N_11447,N_10108,N_10559);
nor U11448 (N_11448,N_10886,N_10887);
and U11449 (N_11449,N_10153,N_10911);
nor U11450 (N_11450,N_10762,N_10251);
or U11451 (N_11451,N_10022,N_10630);
and U11452 (N_11452,N_10496,N_10507);
and U11453 (N_11453,N_10356,N_10679);
nand U11454 (N_11454,N_10519,N_10892);
and U11455 (N_11455,N_10536,N_10614);
and U11456 (N_11456,N_10763,N_10700);
and U11457 (N_11457,N_10924,N_10730);
nor U11458 (N_11458,N_10897,N_10347);
or U11459 (N_11459,N_10468,N_10103);
or U11460 (N_11460,N_10799,N_10229);
nor U11461 (N_11461,N_10284,N_10270);
and U11462 (N_11462,N_10498,N_10869);
and U11463 (N_11463,N_10374,N_10275);
nor U11464 (N_11464,N_10976,N_10118);
nor U11465 (N_11465,N_10875,N_10640);
nor U11466 (N_11466,N_10204,N_10167);
or U11467 (N_11467,N_10907,N_10528);
nand U11468 (N_11468,N_10716,N_10492);
nand U11469 (N_11469,N_10658,N_10168);
nand U11470 (N_11470,N_10858,N_10698);
and U11471 (N_11471,N_10726,N_10254);
and U11472 (N_11472,N_10535,N_10612);
or U11473 (N_11473,N_10324,N_10529);
nand U11474 (N_11474,N_10734,N_10358);
nand U11475 (N_11475,N_10160,N_10091);
nor U11476 (N_11476,N_10984,N_10560);
or U11477 (N_11477,N_10741,N_10710);
and U11478 (N_11478,N_10817,N_10169);
nand U11479 (N_11479,N_10968,N_10310);
nand U11480 (N_11480,N_10297,N_10537);
and U11481 (N_11481,N_10629,N_10353);
and U11482 (N_11482,N_10722,N_10479);
and U11483 (N_11483,N_10064,N_10901);
or U11484 (N_11484,N_10582,N_10462);
and U11485 (N_11485,N_10370,N_10676);
and U11486 (N_11486,N_10001,N_10602);
or U11487 (N_11487,N_10259,N_10597);
nand U11488 (N_11488,N_10483,N_10303);
or U11489 (N_11489,N_10246,N_10008);
nor U11490 (N_11490,N_10200,N_10053);
nand U11491 (N_11491,N_10811,N_10983);
and U11492 (N_11492,N_10866,N_10481);
or U11493 (N_11493,N_10777,N_10269);
nand U11494 (N_11494,N_10006,N_10647);
or U11495 (N_11495,N_10120,N_10625);
or U11496 (N_11496,N_10009,N_10451);
nand U11497 (N_11497,N_10129,N_10986);
nand U11498 (N_11498,N_10449,N_10140);
or U11499 (N_11499,N_10689,N_10955);
nor U11500 (N_11500,N_10937,N_10640);
nor U11501 (N_11501,N_10317,N_10875);
and U11502 (N_11502,N_10902,N_10380);
nor U11503 (N_11503,N_10878,N_10069);
and U11504 (N_11504,N_10953,N_10527);
or U11505 (N_11505,N_10505,N_10509);
nor U11506 (N_11506,N_10324,N_10381);
or U11507 (N_11507,N_10647,N_10639);
or U11508 (N_11508,N_10688,N_10482);
or U11509 (N_11509,N_10507,N_10757);
and U11510 (N_11510,N_10824,N_10360);
nand U11511 (N_11511,N_10652,N_10229);
or U11512 (N_11512,N_10226,N_10572);
and U11513 (N_11513,N_10503,N_10719);
and U11514 (N_11514,N_10273,N_10361);
or U11515 (N_11515,N_10726,N_10354);
or U11516 (N_11516,N_10040,N_10656);
nor U11517 (N_11517,N_10797,N_10198);
nor U11518 (N_11518,N_10994,N_10055);
and U11519 (N_11519,N_10671,N_10447);
nand U11520 (N_11520,N_10940,N_10140);
nor U11521 (N_11521,N_10984,N_10605);
or U11522 (N_11522,N_10906,N_10234);
or U11523 (N_11523,N_10375,N_10283);
nand U11524 (N_11524,N_10575,N_10445);
nor U11525 (N_11525,N_10420,N_10415);
nand U11526 (N_11526,N_10331,N_10368);
nand U11527 (N_11527,N_10435,N_10907);
and U11528 (N_11528,N_10631,N_10012);
and U11529 (N_11529,N_10216,N_10794);
nor U11530 (N_11530,N_10713,N_10428);
nand U11531 (N_11531,N_10541,N_10210);
nand U11532 (N_11532,N_10715,N_10489);
or U11533 (N_11533,N_10473,N_10219);
and U11534 (N_11534,N_10095,N_10193);
nor U11535 (N_11535,N_10074,N_10551);
and U11536 (N_11536,N_10612,N_10278);
and U11537 (N_11537,N_10690,N_10346);
or U11538 (N_11538,N_10526,N_10576);
nand U11539 (N_11539,N_10193,N_10688);
or U11540 (N_11540,N_10142,N_10018);
or U11541 (N_11541,N_10933,N_10327);
or U11542 (N_11542,N_10440,N_10124);
and U11543 (N_11543,N_10613,N_10031);
or U11544 (N_11544,N_10851,N_10170);
nand U11545 (N_11545,N_10545,N_10725);
or U11546 (N_11546,N_10366,N_10750);
and U11547 (N_11547,N_10732,N_10341);
or U11548 (N_11548,N_10833,N_10995);
or U11549 (N_11549,N_10754,N_10339);
nand U11550 (N_11550,N_10359,N_10288);
or U11551 (N_11551,N_10780,N_10255);
nor U11552 (N_11552,N_10214,N_10354);
nor U11553 (N_11553,N_10647,N_10427);
or U11554 (N_11554,N_10507,N_10244);
nand U11555 (N_11555,N_10445,N_10414);
and U11556 (N_11556,N_10034,N_10857);
nor U11557 (N_11557,N_10439,N_10591);
and U11558 (N_11558,N_10293,N_10448);
and U11559 (N_11559,N_10859,N_10489);
and U11560 (N_11560,N_10806,N_10358);
or U11561 (N_11561,N_10616,N_10845);
nor U11562 (N_11562,N_10834,N_10704);
nand U11563 (N_11563,N_10310,N_10488);
and U11564 (N_11564,N_10194,N_10882);
nor U11565 (N_11565,N_10894,N_10578);
nand U11566 (N_11566,N_10732,N_10059);
nand U11567 (N_11567,N_10967,N_10809);
nand U11568 (N_11568,N_10916,N_10903);
nor U11569 (N_11569,N_10783,N_10955);
nand U11570 (N_11570,N_10682,N_10337);
or U11571 (N_11571,N_10114,N_10794);
nor U11572 (N_11572,N_10088,N_10296);
nand U11573 (N_11573,N_10000,N_10263);
or U11574 (N_11574,N_10470,N_10098);
and U11575 (N_11575,N_10336,N_10118);
and U11576 (N_11576,N_10999,N_10342);
nand U11577 (N_11577,N_10711,N_10390);
nor U11578 (N_11578,N_10323,N_10653);
and U11579 (N_11579,N_10778,N_10299);
and U11580 (N_11580,N_10021,N_10087);
nor U11581 (N_11581,N_10123,N_10575);
nand U11582 (N_11582,N_10136,N_10135);
nor U11583 (N_11583,N_10152,N_10091);
nand U11584 (N_11584,N_10924,N_10012);
and U11585 (N_11585,N_10577,N_10301);
nor U11586 (N_11586,N_10168,N_10751);
nand U11587 (N_11587,N_10933,N_10679);
nand U11588 (N_11588,N_10210,N_10235);
nor U11589 (N_11589,N_10452,N_10587);
nor U11590 (N_11590,N_10207,N_10221);
nand U11591 (N_11591,N_10417,N_10673);
or U11592 (N_11592,N_10755,N_10146);
and U11593 (N_11593,N_10593,N_10421);
and U11594 (N_11594,N_10033,N_10127);
or U11595 (N_11595,N_10775,N_10950);
and U11596 (N_11596,N_10272,N_10054);
and U11597 (N_11597,N_10271,N_10220);
nor U11598 (N_11598,N_10737,N_10419);
nor U11599 (N_11599,N_10824,N_10546);
nor U11600 (N_11600,N_10074,N_10791);
or U11601 (N_11601,N_10056,N_10743);
nor U11602 (N_11602,N_10839,N_10613);
or U11603 (N_11603,N_10197,N_10805);
and U11604 (N_11604,N_10721,N_10177);
nor U11605 (N_11605,N_10960,N_10824);
and U11606 (N_11606,N_10786,N_10377);
nor U11607 (N_11607,N_10491,N_10848);
and U11608 (N_11608,N_10222,N_10409);
or U11609 (N_11609,N_10198,N_10019);
nor U11610 (N_11610,N_10807,N_10799);
nand U11611 (N_11611,N_10122,N_10083);
nand U11612 (N_11612,N_10106,N_10127);
and U11613 (N_11613,N_10751,N_10194);
or U11614 (N_11614,N_10747,N_10106);
nor U11615 (N_11615,N_10090,N_10236);
nor U11616 (N_11616,N_10535,N_10385);
nand U11617 (N_11617,N_10767,N_10825);
nor U11618 (N_11618,N_10027,N_10218);
nor U11619 (N_11619,N_10449,N_10843);
or U11620 (N_11620,N_10653,N_10284);
or U11621 (N_11621,N_10937,N_10856);
or U11622 (N_11622,N_10331,N_10159);
and U11623 (N_11623,N_10840,N_10269);
nor U11624 (N_11624,N_10184,N_10496);
nor U11625 (N_11625,N_10327,N_10342);
nand U11626 (N_11626,N_10677,N_10347);
or U11627 (N_11627,N_10557,N_10888);
or U11628 (N_11628,N_10410,N_10761);
nor U11629 (N_11629,N_10826,N_10927);
or U11630 (N_11630,N_10499,N_10706);
and U11631 (N_11631,N_10032,N_10458);
or U11632 (N_11632,N_10736,N_10240);
nand U11633 (N_11633,N_10848,N_10063);
and U11634 (N_11634,N_10033,N_10585);
or U11635 (N_11635,N_10197,N_10732);
and U11636 (N_11636,N_10332,N_10891);
and U11637 (N_11637,N_10360,N_10908);
nand U11638 (N_11638,N_10755,N_10268);
nor U11639 (N_11639,N_10957,N_10730);
nand U11640 (N_11640,N_10137,N_10951);
or U11641 (N_11641,N_10660,N_10763);
nor U11642 (N_11642,N_10415,N_10862);
or U11643 (N_11643,N_10371,N_10761);
or U11644 (N_11644,N_10019,N_10135);
nand U11645 (N_11645,N_10415,N_10104);
and U11646 (N_11646,N_10715,N_10607);
nand U11647 (N_11647,N_10556,N_10495);
and U11648 (N_11648,N_10205,N_10768);
nor U11649 (N_11649,N_10326,N_10916);
and U11650 (N_11650,N_10757,N_10976);
nand U11651 (N_11651,N_10078,N_10667);
nand U11652 (N_11652,N_10415,N_10620);
nand U11653 (N_11653,N_10043,N_10844);
and U11654 (N_11654,N_10585,N_10541);
and U11655 (N_11655,N_10873,N_10813);
nand U11656 (N_11656,N_10926,N_10345);
nand U11657 (N_11657,N_10739,N_10818);
and U11658 (N_11658,N_10638,N_10583);
nand U11659 (N_11659,N_10989,N_10877);
and U11660 (N_11660,N_10307,N_10421);
nor U11661 (N_11661,N_10079,N_10898);
nand U11662 (N_11662,N_10799,N_10802);
or U11663 (N_11663,N_10248,N_10433);
and U11664 (N_11664,N_10180,N_10593);
and U11665 (N_11665,N_10092,N_10528);
and U11666 (N_11666,N_10905,N_10238);
nand U11667 (N_11667,N_10118,N_10684);
nor U11668 (N_11668,N_10783,N_10801);
or U11669 (N_11669,N_10531,N_10011);
nand U11670 (N_11670,N_10830,N_10344);
or U11671 (N_11671,N_10868,N_10288);
nand U11672 (N_11672,N_10859,N_10816);
or U11673 (N_11673,N_10393,N_10092);
and U11674 (N_11674,N_10432,N_10429);
and U11675 (N_11675,N_10464,N_10019);
nor U11676 (N_11676,N_10438,N_10975);
nand U11677 (N_11677,N_10331,N_10689);
and U11678 (N_11678,N_10076,N_10271);
nor U11679 (N_11679,N_10803,N_10010);
nand U11680 (N_11680,N_10253,N_10328);
and U11681 (N_11681,N_10751,N_10710);
and U11682 (N_11682,N_10593,N_10090);
or U11683 (N_11683,N_10491,N_10385);
and U11684 (N_11684,N_10697,N_10490);
and U11685 (N_11685,N_10417,N_10080);
nor U11686 (N_11686,N_10764,N_10252);
nand U11687 (N_11687,N_10065,N_10332);
or U11688 (N_11688,N_10941,N_10735);
nand U11689 (N_11689,N_10195,N_10116);
or U11690 (N_11690,N_10426,N_10031);
or U11691 (N_11691,N_10298,N_10334);
nor U11692 (N_11692,N_10024,N_10948);
nor U11693 (N_11693,N_10849,N_10065);
nor U11694 (N_11694,N_10782,N_10198);
and U11695 (N_11695,N_10134,N_10823);
nand U11696 (N_11696,N_10798,N_10207);
or U11697 (N_11697,N_10847,N_10557);
and U11698 (N_11698,N_10256,N_10005);
and U11699 (N_11699,N_10501,N_10253);
nor U11700 (N_11700,N_10173,N_10843);
nand U11701 (N_11701,N_10282,N_10099);
nand U11702 (N_11702,N_10065,N_10396);
xnor U11703 (N_11703,N_10947,N_10950);
and U11704 (N_11704,N_10916,N_10015);
or U11705 (N_11705,N_10544,N_10708);
or U11706 (N_11706,N_10026,N_10288);
nand U11707 (N_11707,N_10250,N_10835);
nand U11708 (N_11708,N_10317,N_10977);
nand U11709 (N_11709,N_10304,N_10318);
nor U11710 (N_11710,N_10324,N_10311);
nand U11711 (N_11711,N_10200,N_10275);
nor U11712 (N_11712,N_10384,N_10883);
nand U11713 (N_11713,N_10851,N_10090);
nor U11714 (N_11714,N_10799,N_10101);
or U11715 (N_11715,N_10857,N_10413);
or U11716 (N_11716,N_10767,N_10579);
and U11717 (N_11717,N_10967,N_10987);
or U11718 (N_11718,N_10573,N_10118);
and U11719 (N_11719,N_10084,N_10487);
nor U11720 (N_11720,N_10900,N_10227);
or U11721 (N_11721,N_10325,N_10216);
or U11722 (N_11722,N_10614,N_10230);
and U11723 (N_11723,N_10523,N_10861);
nor U11724 (N_11724,N_10408,N_10967);
and U11725 (N_11725,N_10607,N_10435);
nand U11726 (N_11726,N_10626,N_10346);
and U11727 (N_11727,N_10080,N_10803);
nor U11728 (N_11728,N_10626,N_10457);
nor U11729 (N_11729,N_10074,N_10068);
nor U11730 (N_11730,N_10550,N_10576);
or U11731 (N_11731,N_10740,N_10866);
nand U11732 (N_11732,N_10029,N_10325);
nor U11733 (N_11733,N_10409,N_10365);
nor U11734 (N_11734,N_10992,N_10748);
nand U11735 (N_11735,N_10712,N_10777);
or U11736 (N_11736,N_10581,N_10936);
nor U11737 (N_11737,N_10611,N_10898);
nand U11738 (N_11738,N_10922,N_10579);
nand U11739 (N_11739,N_10849,N_10536);
or U11740 (N_11740,N_10141,N_10404);
and U11741 (N_11741,N_10809,N_10141);
and U11742 (N_11742,N_10654,N_10095);
and U11743 (N_11743,N_10649,N_10562);
nand U11744 (N_11744,N_10556,N_10328);
nand U11745 (N_11745,N_10699,N_10167);
nand U11746 (N_11746,N_10313,N_10123);
nand U11747 (N_11747,N_10980,N_10822);
nand U11748 (N_11748,N_10206,N_10765);
or U11749 (N_11749,N_10117,N_10641);
nor U11750 (N_11750,N_10006,N_10886);
or U11751 (N_11751,N_10430,N_10146);
nor U11752 (N_11752,N_10886,N_10755);
and U11753 (N_11753,N_10353,N_10598);
nor U11754 (N_11754,N_10069,N_10492);
nor U11755 (N_11755,N_10060,N_10751);
nand U11756 (N_11756,N_10032,N_10594);
and U11757 (N_11757,N_10604,N_10766);
nor U11758 (N_11758,N_10039,N_10316);
nand U11759 (N_11759,N_10406,N_10757);
nor U11760 (N_11760,N_10184,N_10531);
and U11761 (N_11761,N_10819,N_10411);
or U11762 (N_11762,N_10665,N_10845);
nor U11763 (N_11763,N_10960,N_10831);
or U11764 (N_11764,N_10596,N_10634);
nor U11765 (N_11765,N_10599,N_10704);
nand U11766 (N_11766,N_10804,N_10738);
and U11767 (N_11767,N_10508,N_10227);
or U11768 (N_11768,N_10023,N_10623);
nand U11769 (N_11769,N_10335,N_10549);
nand U11770 (N_11770,N_10082,N_10370);
and U11771 (N_11771,N_10117,N_10014);
nand U11772 (N_11772,N_10557,N_10425);
and U11773 (N_11773,N_10993,N_10436);
nor U11774 (N_11774,N_10651,N_10323);
nor U11775 (N_11775,N_10436,N_10202);
nand U11776 (N_11776,N_10699,N_10565);
and U11777 (N_11777,N_10683,N_10628);
nor U11778 (N_11778,N_10230,N_10482);
nor U11779 (N_11779,N_10732,N_10207);
nor U11780 (N_11780,N_10071,N_10513);
xnor U11781 (N_11781,N_10509,N_10487);
nor U11782 (N_11782,N_10004,N_10907);
nand U11783 (N_11783,N_10507,N_10918);
nor U11784 (N_11784,N_10415,N_10726);
nor U11785 (N_11785,N_10928,N_10513);
or U11786 (N_11786,N_10114,N_10990);
or U11787 (N_11787,N_10888,N_10239);
nor U11788 (N_11788,N_10650,N_10602);
and U11789 (N_11789,N_10707,N_10333);
nor U11790 (N_11790,N_10360,N_10411);
or U11791 (N_11791,N_10872,N_10612);
or U11792 (N_11792,N_10322,N_10178);
nand U11793 (N_11793,N_10133,N_10536);
nand U11794 (N_11794,N_10943,N_10476);
xor U11795 (N_11795,N_10051,N_10408);
and U11796 (N_11796,N_10430,N_10173);
nand U11797 (N_11797,N_10476,N_10612);
nand U11798 (N_11798,N_10762,N_10565);
nand U11799 (N_11799,N_10614,N_10023);
nor U11800 (N_11800,N_10089,N_10620);
or U11801 (N_11801,N_10004,N_10371);
nor U11802 (N_11802,N_10066,N_10297);
and U11803 (N_11803,N_10211,N_10755);
and U11804 (N_11804,N_10594,N_10952);
nand U11805 (N_11805,N_10587,N_10561);
nor U11806 (N_11806,N_10505,N_10018);
nand U11807 (N_11807,N_10132,N_10700);
and U11808 (N_11808,N_10272,N_10184);
xor U11809 (N_11809,N_10404,N_10567);
nand U11810 (N_11810,N_10488,N_10704);
nand U11811 (N_11811,N_10760,N_10748);
nand U11812 (N_11812,N_10882,N_10412);
nor U11813 (N_11813,N_10534,N_10774);
and U11814 (N_11814,N_10094,N_10243);
nand U11815 (N_11815,N_10981,N_10421);
nand U11816 (N_11816,N_10513,N_10325);
or U11817 (N_11817,N_10790,N_10039);
nor U11818 (N_11818,N_10667,N_10203);
or U11819 (N_11819,N_10789,N_10156);
or U11820 (N_11820,N_10083,N_10809);
nor U11821 (N_11821,N_10045,N_10452);
and U11822 (N_11822,N_10421,N_10699);
nand U11823 (N_11823,N_10388,N_10716);
or U11824 (N_11824,N_10790,N_10031);
nand U11825 (N_11825,N_10291,N_10902);
and U11826 (N_11826,N_10904,N_10525);
or U11827 (N_11827,N_10861,N_10422);
and U11828 (N_11828,N_10231,N_10387);
or U11829 (N_11829,N_10570,N_10617);
and U11830 (N_11830,N_10235,N_10556);
or U11831 (N_11831,N_10902,N_10241);
or U11832 (N_11832,N_10502,N_10186);
nand U11833 (N_11833,N_10294,N_10311);
or U11834 (N_11834,N_10968,N_10532);
and U11835 (N_11835,N_10745,N_10605);
or U11836 (N_11836,N_10078,N_10732);
nor U11837 (N_11837,N_10027,N_10326);
nand U11838 (N_11838,N_10427,N_10755);
and U11839 (N_11839,N_10428,N_10516);
and U11840 (N_11840,N_10563,N_10903);
and U11841 (N_11841,N_10647,N_10727);
nand U11842 (N_11842,N_10340,N_10591);
and U11843 (N_11843,N_10908,N_10366);
or U11844 (N_11844,N_10584,N_10643);
nor U11845 (N_11845,N_10074,N_10194);
or U11846 (N_11846,N_10202,N_10475);
or U11847 (N_11847,N_10705,N_10683);
nand U11848 (N_11848,N_10559,N_10254);
nor U11849 (N_11849,N_10248,N_10846);
nand U11850 (N_11850,N_10754,N_10516);
and U11851 (N_11851,N_10696,N_10453);
or U11852 (N_11852,N_10113,N_10680);
and U11853 (N_11853,N_10939,N_10333);
nor U11854 (N_11854,N_10667,N_10427);
and U11855 (N_11855,N_10782,N_10335);
or U11856 (N_11856,N_10330,N_10592);
nand U11857 (N_11857,N_10508,N_10706);
and U11858 (N_11858,N_10201,N_10564);
nor U11859 (N_11859,N_10055,N_10273);
nor U11860 (N_11860,N_10008,N_10814);
and U11861 (N_11861,N_10386,N_10770);
and U11862 (N_11862,N_10619,N_10303);
xnor U11863 (N_11863,N_10518,N_10223);
nand U11864 (N_11864,N_10479,N_10632);
and U11865 (N_11865,N_10917,N_10548);
or U11866 (N_11866,N_10141,N_10390);
nor U11867 (N_11867,N_10143,N_10903);
nand U11868 (N_11868,N_10004,N_10559);
nand U11869 (N_11869,N_10627,N_10537);
or U11870 (N_11870,N_10056,N_10395);
or U11871 (N_11871,N_10365,N_10600);
nand U11872 (N_11872,N_10158,N_10605);
or U11873 (N_11873,N_10873,N_10937);
nor U11874 (N_11874,N_10224,N_10580);
nor U11875 (N_11875,N_10341,N_10337);
and U11876 (N_11876,N_10252,N_10349);
or U11877 (N_11877,N_10403,N_10126);
or U11878 (N_11878,N_10501,N_10533);
nor U11879 (N_11879,N_10134,N_10048);
and U11880 (N_11880,N_10984,N_10728);
or U11881 (N_11881,N_10281,N_10013);
nand U11882 (N_11882,N_10873,N_10004);
and U11883 (N_11883,N_10978,N_10324);
and U11884 (N_11884,N_10621,N_10395);
nor U11885 (N_11885,N_10754,N_10707);
nor U11886 (N_11886,N_10787,N_10274);
nor U11887 (N_11887,N_10139,N_10057);
and U11888 (N_11888,N_10781,N_10236);
nor U11889 (N_11889,N_10480,N_10014);
and U11890 (N_11890,N_10319,N_10402);
nor U11891 (N_11891,N_10083,N_10079);
and U11892 (N_11892,N_10616,N_10539);
nand U11893 (N_11893,N_10623,N_10079);
nor U11894 (N_11894,N_10042,N_10914);
nor U11895 (N_11895,N_10041,N_10704);
and U11896 (N_11896,N_10891,N_10908);
nand U11897 (N_11897,N_10750,N_10626);
nor U11898 (N_11898,N_10978,N_10164);
or U11899 (N_11899,N_10211,N_10697);
nor U11900 (N_11900,N_10369,N_10954);
and U11901 (N_11901,N_10295,N_10847);
nand U11902 (N_11902,N_10795,N_10802);
and U11903 (N_11903,N_10400,N_10474);
nor U11904 (N_11904,N_10337,N_10665);
or U11905 (N_11905,N_10182,N_10110);
or U11906 (N_11906,N_10335,N_10552);
nor U11907 (N_11907,N_10887,N_10251);
or U11908 (N_11908,N_10537,N_10644);
or U11909 (N_11909,N_10510,N_10531);
nand U11910 (N_11910,N_10204,N_10737);
nand U11911 (N_11911,N_10195,N_10074);
nor U11912 (N_11912,N_10860,N_10821);
nand U11913 (N_11913,N_10318,N_10575);
nor U11914 (N_11914,N_10849,N_10818);
nand U11915 (N_11915,N_10821,N_10610);
and U11916 (N_11916,N_10304,N_10481);
nor U11917 (N_11917,N_10052,N_10962);
nor U11918 (N_11918,N_10130,N_10449);
xor U11919 (N_11919,N_10364,N_10568);
or U11920 (N_11920,N_10848,N_10975);
or U11921 (N_11921,N_10490,N_10971);
nor U11922 (N_11922,N_10821,N_10873);
nand U11923 (N_11923,N_10156,N_10066);
nor U11924 (N_11924,N_10515,N_10067);
nor U11925 (N_11925,N_10395,N_10882);
and U11926 (N_11926,N_10425,N_10724);
nand U11927 (N_11927,N_10681,N_10960);
nor U11928 (N_11928,N_10145,N_10080);
nor U11929 (N_11929,N_10856,N_10240);
or U11930 (N_11930,N_10914,N_10916);
or U11931 (N_11931,N_10838,N_10041);
and U11932 (N_11932,N_10616,N_10528);
or U11933 (N_11933,N_10085,N_10926);
or U11934 (N_11934,N_10043,N_10211);
nand U11935 (N_11935,N_10006,N_10032);
and U11936 (N_11936,N_10231,N_10164);
nand U11937 (N_11937,N_10483,N_10525);
or U11938 (N_11938,N_10143,N_10826);
nor U11939 (N_11939,N_10272,N_10623);
nand U11940 (N_11940,N_10693,N_10318);
nand U11941 (N_11941,N_10090,N_10267);
nand U11942 (N_11942,N_10300,N_10577);
nand U11943 (N_11943,N_10467,N_10792);
and U11944 (N_11944,N_10508,N_10205);
nand U11945 (N_11945,N_10431,N_10878);
nand U11946 (N_11946,N_10968,N_10309);
or U11947 (N_11947,N_10618,N_10386);
and U11948 (N_11948,N_10350,N_10376);
and U11949 (N_11949,N_10174,N_10442);
or U11950 (N_11950,N_10611,N_10487);
nand U11951 (N_11951,N_10524,N_10665);
nor U11952 (N_11952,N_10574,N_10139);
nor U11953 (N_11953,N_10843,N_10440);
and U11954 (N_11954,N_10467,N_10053);
and U11955 (N_11955,N_10580,N_10701);
nor U11956 (N_11956,N_10503,N_10874);
nor U11957 (N_11957,N_10676,N_10155);
and U11958 (N_11958,N_10318,N_10694);
nand U11959 (N_11959,N_10546,N_10191);
and U11960 (N_11960,N_10227,N_10062);
and U11961 (N_11961,N_10101,N_10363);
nor U11962 (N_11962,N_10712,N_10591);
nor U11963 (N_11963,N_10797,N_10680);
or U11964 (N_11964,N_10518,N_10091);
nand U11965 (N_11965,N_10187,N_10835);
or U11966 (N_11966,N_10362,N_10950);
nor U11967 (N_11967,N_10612,N_10266);
and U11968 (N_11968,N_10171,N_10736);
or U11969 (N_11969,N_10687,N_10168);
nand U11970 (N_11970,N_10685,N_10465);
or U11971 (N_11971,N_10872,N_10743);
nand U11972 (N_11972,N_10902,N_10006);
nor U11973 (N_11973,N_10965,N_10248);
nand U11974 (N_11974,N_10186,N_10345);
nand U11975 (N_11975,N_10224,N_10293);
nor U11976 (N_11976,N_10669,N_10535);
nand U11977 (N_11977,N_10869,N_10247);
nand U11978 (N_11978,N_10557,N_10933);
or U11979 (N_11979,N_10785,N_10051);
nor U11980 (N_11980,N_10084,N_10964);
and U11981 (N_11981,N_10690,N_10101);
nor U11982 (N_11982,N_10588,N_10532);
or U11983 (N_11983,N_10616,N_10136);
nand U11984 (N_11984,N_10280,N_10797);
or U11985 (N_11985,N_10911,N_10934);
and U11986 (N_11986,N_10745,N_10950);
nor U11987 (N_11987,N_10961,N_10056);
nand U11988 (N_11988,N_10179,N_10491);
or U11989 (N_11989,N_10957,N_10413);
and U11990 (N_11990,N_10989,N_10064);
and U11991 (N_11991,N_10431,N_10106);
nand U11992 (N_11992,N_10924,N_10831);
nor U11993 (N_11993,N_10580,N_10544);
or U11994 (N_11994,N_10241,N_10908);
nand U11995 (N_11995,N_10000,N_10150);
nor U11996 (N_11996,N_10566,N_10214);
or U11997 (N_11997,N_10307,N_10353);
or U11998 (N_11998,N_10596,N_10897);
and U11999 (N_11999,N_10973,N_10556);
nor U12000 (N_12000,N_11116,N_11942);
or U12001 (N_12001,N_11084,N_11809);
or U12002 (N_12002,N_11453,N_11724);
nand U12003 (N_12003,N_11923,N_11940);
nand U12004 (N_12004,N_11554,N_11027);
nand U12005 (N_12005,N_11450,N_11402);
and U12006 (N_12006,N_11862,N_11120);
nor U12007 (N_12007,N_11593,N_11657);
or U12008 (N_12008,N_11331,N_11845);
nor U12009 (N_12009,N_11600,N_11935);
or U12010 (N_12010,N_11165,N_11231);
nand U12011 (N_12011,N_11547,N_11031);
nor U12012 (N_12012,N_11028,N_11322);
nor U12013 (N_12013,N_11202,N_11772);
and U12014 (N_12014,N_11316,N_11083);
and U12015 (N_12015,N_11236,N_11254);
nand U12016 (N_12016,N_11419,N_11278);
and U12017 (N_12017,N_11005,N_11753);
and U12018 (N_12018,N_11454,N_11505);
nand U12019 (N_12019,N_11650,N_11915);
and U12020 (N_12020,N_11251,N_11150);
nand U12021 (N_12021,N_11598,N_11566);
nor U12022 (N_12022,N_11426,N_11726);
and U12023 (N_12023,N_11892,N_11347);
and U12024 (N_12024,N_11571,N_11436);
and U12025 (N_12025,N_11752,N_11981);
nor U12026 (N_12026,N_11445,N_11523);
nor U12027 (N_12027,N_11449,N_11335);
nand U12028 (N_12028,N_11570,N_11574);
or U12029 (N_12029,N_11379,N_11536);
nand U12030 (N_12030,N_11243,N_11813);
or U12031 (N_12031,N_11766,N_11645);
nand U12032 (N_12032,N_11023,N_11765);
nor U12033 (N_12033,N_11176,N_11821);
or U12034 (N_12034,N_11201,N_11599);
and U12035 (N_12035,N_11431,N_11851);
and U12036 (N_12036,N_11149,N_11049);
and U12037 (N_12037,N_11115,N_11587);
or U12038 (N_12038,N_11016,N_11706);
and U12039 (N_12039,N_11998,N_11467);
nand U12040 (N_12040,N_11485,N_11954);
nand U12041 (N_12041,N_11708,N_11052);
nand U12042 (N_12042,N_11489,N_11070);
nand U12043 (N_12043,N_11819,N_11302);
nor U12044 (N_12044,N_11518,N_11076);
or U12045 (N_12045,N_11994,N_11349);
nor U12046 (N_12046,N_11498,N_11939);
nor U12047 (N_12047,N_11517,N_11350);
and U12048 (N_12048,N_11656,N_11672);
or U12049 (N_12049,N_11741,N_11546);
nor U12050 (N_12050,N_11849,N_11143);
or U12051 (N_12051,N_11397,N_11261);
and U12052 (N_12052,N_11369,N_11474);
and U12053 (N_12053,N_11738,N_11889);
nand U12054 (N_12054,N_11913,N_11673);
nor U12055 (N_12055,N_11004,N_11705);
or U12056 (N_12056,N_11992,N_11987);
nand U12057 (N_12057,N_11240,N_11944);
nor U12058 (N_12058,N_11875,N_11100);
or U12059 (N_12059,N_11924,N_11929);
or U12060 (N_12060,N_11811,N_11011);
nor U12061 (N_12061,N_11400,N_11962);
and U12062 (N_12062,N_11660,N_11647);
or U12063 (N_12063,N_11510,N_11702);
nand U12064 (N_12064,N_11095,N_11793);
nor U12065 (N_12065,N_11636,N_11443);
or U12066 (N_12066,N_11947,N_11687);
nor U12067 (N_12067,N_11665,N_11334);
nor U12068 (N_12068,N_11319,N_11899);
or U12069 (N_12069,N_11978,N_11195);
and U12070 (N_12070,N_11662,N_11373);
nand U12071 (N_12071,N_11325,N_11293);
or U12072 (N_12072,N_11385,N_11843);
nor U12073 (N_12073,N_11001,N_11966);
and U12074 (N_12074,N_11663,N_11241);
nand U12075 (N_12075,N_11042,N_11785);
and U12076 (N_12076,N_11631,N_11117);
nor U12077 (N_12077,N_11689,N_11879);
or U12078 (N_12078,N_11051,N_11317);
and U12079 (N_12079,N_11473,N_11310);
or U12080 (N_12080,N_11842,N_11520);
nand U12081 (N_12081,N_11792,N_11747);
nand U12082 (N_12082,N_11368,N_11465);
nand U12083 (N_12083,N_11728,N_11207);
or U12084 (N_12084,N_11912,N_11774);
or U12085 (N_12085,N_11957,N_11769);
or U12086 (N_12086,N_11700,N_11054);
nor U12087 (N_12087,N_11602,N_11839);
and U12088 (N_12088,N_11579,N_11305);
nand U12089 (N_12089,N_11896,N_11482);
or U12090 (N_12090,N_11595,N_11079);
nor U12091 (N_12091,N_11914,N_11577);
or U12092 (N_12092,N_11122,N_11210);
and U12093 (N_12093,N_11416,N_11346);
nand U12094 (N_12094,N_11737,N_11945);
and U12095 (N_12095,N_11556,N_11246);
and U12096 (N_12096,N_11275,N_11492);
or U12097 (N_12097,N_11794,N_11736);
nor U12098 (N_12098,N_11628,N_11418);
or U12099 (N_12099,N_11890,N_11191);
and U12100 (N_12100,N_11098,N_11442);
nor U12101 (N_12101,N_11539,N_11357);
nand U12102 (N_12102,N_11363,N_11804);
or U12103 (N_12103,N_11818,N_11999);
nand U12104 (N_12104,N_11290,N_11757);
nand U12105 (N_12105,N_11003,N_11641);
or U12106 (N_12106,N_11615,N_11755);
or U12107 (N_12107,N_11208,N_11718);
nand U12108 (N_12108,N_11131,N_11775);
and U12109 (N_12109,N_11424,N_11730);
nand U12110 (N_12110,N_11918,N_11986);
nor U12111 (N_12111,N_11040,N_11676);
or U12112 (N_12112,N_11487,N_11974);
or U12113 (N_12113,N_11903,N_11359);
nor U12114 (N_12114,N_11220,N_11959);
and U12115 (N_12115,N_11965,N_11835);
and U12116 (N_12116,N_11211,N_11941);
nand U12117 (N_12117,N_11611,N_11073);
nand U12118 (N_12118,N_11614,N_11980);
nor U12119 (N_12119,N_11691,N_11438);
or U12120 (N_12120,N_11114,N_11332);
nor U12121 (N_12121,N_11770,N_11277);
and U12122 (N_12122,N_11366,N_11723);
nor U12123 (N_12123,N_11783,N_11074);
nor U12124 (N_12124,N_11107,N_11789);
nor U12125 (N_12125,N_11434,N_11938);
nor U12126 (N_12126,N_11681,N_11483);
and U12127 (N_12127,N_11716,N_11091);
nor U12128 (N_12128,N_11597,N_11573);
or U12129 (N_12129,N_11226,N_11499);
nand U12130 (N_12130,N_11285,N_11298);
or U12131 (N_12131,N_11104,N_11612);
nor U12132 (N_12132,N_11704,N_11739);
and U12133 (N_12133,N_11190,N_11734);
nor U12134 (N_12134,N_11435,N_11745);
and U12135 (N_12135,N_11856,N_11698);
nor U12136 (N_12136,N_11067,N_11948);
nor U12137 (N_12137,N_11559,N_11633);
or U12138 (N_12138,N_11232,N_11670);
nand U12139 (N_12139,N_11015,N_11626);
or U12140 (N_12140,N_11427,N_11197);
or U12141 (N_12141,N_11922,N_11946);
or U12142 (N_12142,N_11420,N_11163);
nor U12143 (N_12143,N_11183,N_11853);
nor U12144 (N_12144,N_11399,N_11292);
nor U12145 (N_12145,N_11549,N_11330);
nand U12146 (N_12146,N_11963,N_11223);
and U12147 (N_12147,N_11508,N_11072);
or U12148 (N_12148,N_11652,N_11224);
nand U12149 (N_12149,N_11830,N_11158);
and U12150 (N_12150,N_11428,N_11287);
nand U12151 (N_12151,N_11022,N_11297);
and U12152 (N_12152,N_11627,N_11867);
and U12153 (N_12153,N_11280,N_11413);
and U12154 (N_12154,N_11196,N_11970);
or U12155 (N_12155,N_11021,N_11129);
nand U12156 (N_12156,N_11527,N_11898);
nand U12157 (N_12157,N_11175,N_11250);
nand U12158 (N_12158,N_11266,N_11490);
and U12159 (N_12159,N_11771,N_11356);
and U12160 (N_12160,N_11823,N_11475);
nand U12161 (N_12161,N_11113,N_11586);
nor U12162 (N_12162,N_11184,N_11919);
nand U12163 (N_12163,N_11460,N_11082);
nor U12164 (N_12164,N_11758,N_11264);
or U12165 (N_12165,N_11217,N_11168);
nand U12166 (N_12166,N_11256,N_11638);
and U12167 (N_12167,N_11212,N_11282);
and U12168 (N_12168,N_11905,N_11410);
xnor U12169 (N_12169,N_11964,N_11674);
nor U12170 (N_12170,N_11136,N_11563);
nand U12171 (N_12171,N_11119,N_11312);
or U12172 (N_12172,N_11582,N_11625);
nand U12173 (N_12173,N_11058,N_11642);
or U12174 (N_12174,N_11046,N_11699);
nor U12175 (N_12175,N_11388,N_11019);
or U12176 (N_12176,N_11484,N_11390);
and U12177 (N_12177,N_11404,N_11541);
and U12178 (N_12178,N_11105,N_11050);
or U12179 (N_12179,N_11927,N_11459);
or U12180 (N_12180,N_11315,N_11081);
and U12181 (N_12181,N_11881,N_11291);
nand U12182 (N_12182,N_11815,N_11542);
nor U12183 (N_12183,N_11463,N_11384);
and U12184 (N_12184,N_11043,N_11895);
nor U12185 (N_12185,N_11784,N_11760);
and U12186 (N_12186,N_11786,N_11407);
nor U12187 (N_12187,N_11365,N_11761);
and U12188 (N_12188,N_11893,N_11778);
nand U12189 (N_12189,N_11267,N_11382);
nor U12190 (N_12190,N_11683,N_11692);
or U12191 (N_12191,N_11500,N_11213);
nand U12192 (N_12192,N_11863,N_11167);
nor U12193 (N_12193,N_11949,N_11861);
xor U12194 (N_12194,N_11985,N_11956);
or U12195 (N_12195,N_11584,N_11677);
and U12196 (N_12196,N_11328,N_11776);
or U12197 (N_12197,N_11480,N_11429);
or U12198 (N_12198,N_11558,N_11376);
nor U12199 (N_12199,N_11478,N_11130);
nand U12200 (N_12200,N_11118,N_11873);
nor U12201 (N_12201,N_11838,N_11621);
and U12202 (N_12202,N_11060,N_11069);
nand U12203 (N_12203,N_11779,N_11528);
or U12204 (N_12204,N_11958,N_11353);
nor U12205 (N_12205,N_11086,N_11930);
nand U12206 (N_12206,N_11870,N_11010);
nand U12207 (N_12207,N_11911,N_11807);
nand U12208 (N_12208,N_11777,N_11173);
nor U12209 (N_12209,N_11780,N_11925);
nand U12210 (N_12210,N_11354,N_11617);
or U12211 (N_12211,N_11170,N_11560);
nor U12212 (N_12212,N_11455,N_11697);
nand U12213 (N_12213,N_11068,N_11448);
and U12214 (N_12214,N_11472,N_11844);
or U12215 (N_12215,N_11592,N_11178);
xnor U12216 (N_12216,N_11321,N_11502);
nand U12217 (N_12217,N_11034,N_11995);
nand U12218 (N_12218,N_11147,N_11378);
nor U12219 (N_12219,N_11580,N_11111);
nor U12220 (N_12220,N_11591,N_11880);
and U12221 (N_12221,N_11491,N_11979);
nand U12222 (N_12222,N_11768,N_11565);
nor U12223 (N_12223,N_11693,N_11237);
nand U12224 (N_12224,N_11869,N_11507);
or U12225 (N_12225,N_11790,N_11715);
nor U12226 (N_12226,N_11061,N_11516);
or U12227 (N_12227,N_11537,N_11375);
nor U12228 (N_12228,N_11216,N_11194);
or U12229 (N_12229,N_11634,N_11294);
nand U12230 (N_12230,N_11831,N_11470);
or U12231 (N_12231,N_11495,N_11743);
and U12232 (N_12232,N_11406,N_11457);
nand U12233 (N_12233,N_11193,N_11872);
and U12234 (N_12234,N_11464,N_11253);
or U12235 (N_12235,N_11396,N_11719);
nor U12236 (N_12236,N_11504,N_11742);
nand U12237 (N_12237,N_11198,N_11658);
or U12238 (N_12238,N_11572,N_11910);
nand U12239 (N_12239,N_11125,N_11740);
or U12240 (N_12240,N_11169,N_11735);
and U12241 (N_12241,N_11497,N_11336);
nor U12242 (N_12242,N_11530,N_11206);
and U12243 (N_12243,N_11444,N_11000);
nor U12244 (N_12244,N_11952,N_11340);
or U12245 (N_12245,N_11127,N_11901);
and U12246 (N_12246,N_11616,N_11605);
nor U12247 (N_12247,N_11533,N_11540);
nor U12248 (N_12248,N_11447,N_11437);
nor U12249 (N_12249,N_11188,N_11555);
nor U12250 (N_12250,N_11265,N_11848);
and U12251 (N_12251,N_11764,N_11812);
nor U12252 (N_12252,N_11171,N_11931);
nor U12253 (N_12253,N_11675,N_11065);
or U12254 (N_12254,N_11415,N_11306);
and U12255 (N_12255,N_11215,N_11393);
nand U12256 (N_12256,N_11270,N_11466);
nor U12257 (N_12257,N_11151,N_11020);
nand U12258 (N_12258,N_11064,N_11679);
nor U12259 (N_12259,N_11759,N_11684);
nand U12260 (N_12260,N_11531,N_11274);
nand U12261 (N_12261,N_11339,N_11829);
and U12262 (N_12262,N_11341,N_11525);
nor U12263 (N_12263,N_11623,N_11874);
and U12264 (N_12264,N_11351,N_11865);
or U12265 (N_12265,N_11653,N_11799);
nand U12266 (N_12266,N_11696,N_11797);
or U12267 (N_12267,N_11686,N_11134);
nand U12268 (N_12268,N_11878,N_11097);
nor U12269 (N_12269,N_11661,N_11668);
or U12270 (N_12270,N_11493,N_11891);
nand U12271 (N_12271,N_11141,N_11648);
nor U12272 (N_12272,N_11486,N_11229);
nor U12273 (N_12273,N_11313,N_11303);
nand U12274 (N_12274,N_11383,N_11386);
and U12275 (N_12275,N_11900,N_11707);
nor U12276 (N_12276,N_11284,N_11909);
nor U12277 (N_12277,N_11128,N_11701);
or U12278 (N_12278,N_11477,N_11245);
or U12279 (N_12279,N_11036,N_11209);
nand U12280 (N_12280,N_11479,N_11047);
or U12281 (N_12281,N_11221,N_11088);
nand U12282 (N_12282,N_11132,N_11904);
xnor U12283 (N_12283,N_11259,N_11551);
nand U12284 (N_12284,N_11808,N_11791);
and U12285 (N_12285,N_11834,N_11272);
nand U12286 (N_12286,N_11468,N_11989);
nor U12287 (N_12287,N_11235,N_11972);
nand U12288 (N_12288,N_11545,N_11519);
and U12289 (N_12289,N_11717,N_11894);
and U12290 (N_12290,N_11532,N_11446);
xor U12291 (N_12291,N_11943,N_11816);
nand U12292 (N_12292,N_11488,N_11973);
nand U12293 (N_12293,N_11884,N_11968);
or U12294 (N_12294,N_11014,N_11389);
or U12295 (N_12295,N_11581,N_11967);
nor U12296 (N_12296,N_11133,N_11139);
nor U12297 (N_12297,N_11348,N_11227);
nor U12298 (N_12298,N_11921,N_11888);
nor U12299 (N_12299,N_11961,N_11762);
nor U12300 (N_12300,N_11934,N_11535);
and U12301 (N_12301,N_11417,N_11377);
or U12302 (N_12302,N_11090,N_11108);
and U12303 (N_12303,N_11897,N_11344);
nor U12304 (N_12304,N_11576,N_11917);
nor U12305 (N_12305,N_11337,N_11859);
nand U12306 (N_12306,N_11976,N_11620);
or U12307 (N_12307,N_11564,N_11077);
nor U12308 (N_12308,N_11039,N_11515);
and U12309 (N_12309,N_11059,N_11864);
nor U12310 (N_12310,N_11123,N_11550);
nor U12311 (N_12311,N_11982,N_11822);
or U12312 (N_12312,N_11087,N_11476);
or U12313 (N_12313,N_11756,N_11326);
and U12314 (N_12314,N_11012,N_11110);
nand U12315 (N_12315,N_11398,N_11876);
nor U12316 (N_12316,N_11725,N_11360);
nand U12317 (N_12317,N_11273,N_11695);
nor U12318 (N_12318,N_11990,N_11607);
nor U12319 (N_12319,N_11886,N_11561);
and U12320 (N_12320,N_11364,N_11361);
nor U12321 (N_12321,N_11618,N_11342);
nor U12322 (N_12322,N_11569,N_11824);
and U12323 (N_12323,N_11112,N_11481);
nor U12324 (N_12324,N_11932,N_11920);
nor U12325 (N_12325,N_11260,N_11374);
or U12326 (N_12326,N_11380,N_11187);
nand U12327 (N_12327,N_11055,N_11802);
and U12328 (N_12328,N_11013,N_11255);
and U12329 (N_12329,N_11056,N_11439);
and U12330 (N_12330,N_11732,N_11093);
or U12331 (N_12331,N_11145,N_11174);
and U12332 (N_12332,N_11276,N_11640);
nor U12333 (N_12333,N_11680,N_11412);
nor U12334 (N_12334,N_11283,N_11846);
nor U12335 (N_12335,N_11782,N_11309);
nor U12336 (N_12336,N_11234,N_11629);
and U12337 (N_12337,N_11109,N_11529);
or U12338 (N_12338,N_11907,N_11308);
nor U12339 (N_12339,N_11749,N_11401);
or U12340 (N_12340,N_11506,N_11295);
and U12341 (N_12341,N_11137,N_11805);
and U12342 (N_12342,N_11144,N_11578);
nand U12343 (N_12343,N_11304,N_11075);
nor U12344 (N_12344,N_11440,N_11601);
nand U12345 (N_12345,N_11690,N_11078);
nand U12346 (N_12346,N_11199,N_11557);
nand U12347 (N_12347,N_11583,N_11152);
nor U12348 (N_12348,N_11214,N_11162);
or U12349 (N_12349,N_11159,N_11422);
or U12350 (N_12350,N_11751,N_11841);
and U12351 (N_12351,N_11955,N_11156);
and U12352 (N_12352,N_11562,N_11832);
and U12353 (N_12353,N_11358,N_11180);
nor U12354 (N_12354,N_11244,N_11323);
nor U12355 (N_12355,N_11024,N_11637);
nor U12356 (N_12356,N_11710,N_11902);
nand U12357 (N_12357,N_11370,N_11269);
or U12358 (N_12358,N_11544,N_11062);
and U12359 (N_12359,N_11763,N_11063);
nand U12360 (N_12360,N_11327,N_11588);
and U12361 (N_12361,N_11318,N_11635);
nand U12362 (N_12362,N_11836,N_11750);
and U12363 (N_12363,N_11575,N_11639);
xnor U12364 (N_12364,N_11858,N_11659);
nor U12365 (N_12365,N_11514,N_11852);
nor U12366 (N_12366,N_11936,N_11263);
nor U12367 (N_12367,N_11085,N_11126);
and U12368 (N_12368,N_11709,N_11320);
nand U12369 (N_12369,N_11367,N_11604);
or U12370 (N_12370,N_11271,N_11606);
or U12371 (N_12371,N_11703,N_11803);
or U12372 (N_12372,N_11773,N_11568);
nand U12373 (N_12373,N_11646,N_11857);
nand U12374 (N_12374,N_11182,N_11017);
nor U12375 (N_12375,N_11458,N_11928);
and U12376 (N_12376,N_11387,N_11155);
or U12377 (N_12377,N_11146,N_11185);
nand U12378 (N_12378,N_11722,N_11984);
or U12379 (N_12379,N_11177,N_11509);
or U12380 (N_12380,N_11613,N_11733);
and U12381 (N_12381,N_11712,N_11589);
nand U12382 (N_12382,N_11664,N_11247);
and U12383 (N_12383,N_11553,N_11008);
nor U12384 (N_12384,N_11311,N_11307);
and U12385 (N_12385,N_11820,N_11372);
and U12386 (N_12386,N_11038,N_11788);
nor U12387 (N_12387,N_11099,N_11007);
and U12388 (N_12388,N_11871,N_11833);
nand U12389 (N_12389,N_11524,N_11101);
or U12390 (N_12390,N_11975,N_11219);
nor U12391 (N_12391,N_11160,N_11603);
and U12392 (N_12392,N_11826,N_11814);
nor U12393 (N_12393,N_11685,N_11996);
or U12394 (N_12394,N_11452,N_11969);
or U12395 (N_12395,N_11721,N_11189);
nand U12396 (N_12396,N_11409,N_11585);
and U12397 (N_12397,N_11071,N_11644);
or U12398 (N_12398,N_11333,N_11837);
and U12399 (N_12399,N_11461,N_11157);
nor U12400 (N_12400,N_11140,N_11825);
nand U12401 (N_12401,N_11522,N_11025);
or U12402 (N_12402,N_11106,N_11142);
nor U12403 (N_12403,N_11230,N_11391);
nand U12404 (N_12404,N_11887,N_11590);
nor U12405 (N_12405,N_11186,N_11496);
and U12406 (N_12406,N_11882,N_11030);
nand U12407 (N_12407,N_11352,N_11154);
and U12408 (N_12408,N_11619,N_11314);
nor U12409 (N_12409,N_11355,N_11854);
nand U12410 (N_12410,N_11866,N_11033);
nor U12411 (N_12411,N_11937,N_11471);
nand U12412 (N_12412,N_11225,N_11800);
or U12413 (N_12413,N_11711,N_11268);
and U12414 (N_12414,N_11667,N_11655);
nor U12415 (N_12415,N_11430,N_11649);
nor U12416 (N_12416,N_11289,N_11503);
nand U12417 (N_12417,N_11624,N_11172);
and U12418 (N_12418,N_11138,N_11026);
nor U12419 (N_12419,N_11096,N_11469);
or U12420 (N_12420,N_11009,N_11767);
nor U12421 (N_12421,N_11511,N_11997);
nor U12422 (N_12422,N_11092,N_11192);
nor U12423 (N_12423,N_11299,N_11827);
xor U12424 (N_12424,N_11850,N_11727);
nor U12425 (N_12425,N_11257,N_11552);
nand U12426 (N_12426,N_11281,N_11433);
and U12427 (N_12427,N_11423,N_11729);
and U12428 (N_12428,N_11610,N_11181);
nor U12429 (N_12429,N_11787,N_11501);
and U12430 (N_12430,N_11045,N_11103);
or U12431 (N_12431,N_11204,N_11029);
or U12432 (N_12432,N_11166,N_11682);
and U12433 (N_12433,N_11411,N_11094);
nand U12434 (N_12434,N_11153,N_11991);
nand U12435 (N_12435,N_11748,N_11993);
nor U12436 (N_12436,N_11885,N_11300);
nor U12437 (N_12437,N_11630,N_11301);
nor U12438 (N_12438,N_11381,N_11526);
nor U12439 (N_12439,N_11249,N_11248);
or U12440 (N_12440,N_11731,N_11608);
and U12441 (N_12441,N_11288,N_11262);
nor U12442 (N_12442,N_11035,N_11037);
nor U12443 (N_12443,N_11988,N_11494);
nor U12444 (N_12444,N_11960,N_11286);
nand U12445 (N_12445,N_11258,N_11746);
nor U12446 (N_12446,N_11983,N_11694);
nor U12447 (N_12447,N_11643,N_11102);
nor U12448 (N_12448,N_11161,N_11951);
or U12449 (N_12449,N_11041,N_11950);
nand U12450 (N_12450,N_11622,N_11044);
and U12451 (N_12451,N_11798,N_11080);
nand U12452 (N_12452,N_11296,N_11203);
nand U12453 (N_12453,N_11343,N_11002);
nand U12454 (N_12454,N_11855,N_11324);
or U12455 (N_12455,N_11164,N_11933);
and U12456 (N_12456,N_11414,N_11394);
or U12457 (N_12457,N_11953,N_11441);
nand U12458 (N_12458,N_11048,N_11926);
or U12459 (N_12459,N_11548,N_11200);
nand U12460 (N_12460,N_11392,N_11408);
and U12461 (N_12461,N_11432,N_11908);
nand U12462 (N_12462,N_11720,N_11860);
nor U12463 (N_12463,N_11252,N_11847);
and U12464 (N_12464,N_11512,N_11688);
nor U12465 (N_12465,N_11395,N_11654);
nor U12466 (N_12466,N_11238,N_11817);
and U12467 (N_12467,N_11279,N_11754);
and U12468 (N_12468,N_11066,N_11877);
and U12469 (N_12469,N_11521,N_11124);
nand U12470 (N_12470,N_11089,N_11538);
nor U12471 (N_12471,N_11371,N_11513);
nand U12472 (N_12472,N_11218,N_11795);
and U12473 (N_12473,N_11713,N_11810);
or U12474 (N_12474,N_11971,N_11148);
and U12475 (N_12475,N_11462,N_11632);
and U12476 (N_12476,N_11669,N_11714);
or U12477 (N_12477,N_11451,N_11594);
or U12478 (N_12478,N_11678,N_11006);
and U12479 (N_12479,N_11840,N_11242);
or U12480 (N_12480,N_11239,N_11906);
nand U12481 (N_12481,N_11228,N_11977);
or U12482 (N_12482,N_11609,N_11828);
nand U12483 (N_12483,N_11671,N_11205);
and U12484 (N_12484,N_11801,N_11222);
and U12485 (N_12485,N_11806,N_11421);
nand U12486 (N_12486,N_11032,N_11233);
nor U12487 (N_12487,N_11179,N_11135);
nor U12488 (N_12488,N_11567,N_11868);
nand U12489 (N_12489,N_11345,N_11916);
nor U12490 (N_12490,N_11329,N_11883);
nor U12491 (N_12491,N_11121,N_11596);
nand U12492 (N_12492,N_11057,N_11796);
nand U12493 (N_12493,N_11651,N_11053);
and U12494 (N_12494,N_11403,N_11338);
nor U12495 (N_12495,N_11405,N_11781);
nand U12496 (N_12496,N_11425,N_11534);
nor U12497 (N_12497,N_11744,N_11362);
and U12498 (N_12498,N_11456,N_11018);
or U12499 (N_12499,N_11543,N_11666);
nor U12500 (N_12500,N_11831,N_11190);
nand U12501 (N_12501,N_11894,N_11228);
nor U12502 (N_12502,N_11371,N_11768);
nor U12503 (N_12503,N_11413,N_11870);
nor U12504 (N_12504,N_11121,N_11930);
nand U12505 (N_12505,N_11660,N_11865);
nand U12506 (N_12506,N_11412,N_11600);
or U12507 (N_12507,N_11348,N_11221);
nand U12508 (N_12508,N_11289,N_11747);
and U12509 (N_12509,N_11374,N_11043);
and U12510 (N_12510,N_11270,N_11360);
nand U12511 (N_12511,N_11978,N_11155);
nor U12512 (N_12512,N_11350,N_11292);
and U12513 (N_12513,N_11967,N_11711);
nor U12514 (N_12514,N_11545,N_11855);
xnor U12515 (N_12515,N_11878,N_11289);
nor U12516 (N_12516,N_11179,N_11251);
and U12517 (N_12517,N_11191,N_11143);
nand U12518 (N_12518,N_11909,N_11716);
nor U12519 (N_12519,N_11876,N_11200);
nand U12520 (N_12520,N_11236,N_11310);
or U12521 (N_12521,N_11423,N_11099);
nor U12522 (N_12522,N_11013,N_11586);
nor U12523 (N_12523,N_11870,N_11485);
or U12524 (N_12524,N_11274,N_11042);
xor U12525 (N_12525,N_11701,N_11510);
nor U12526 (N_12526,N_11505,N_11726);
nor U12527 (N_12527,N_11575,N_11921);
or U12528 (N_12528,N_11651,N_11710);
and U12529 (N_12529,N_11493,N_11924);
nand U12530 (N_12530,N_11904,N_11632);
nand U12531 (N_12531,N_11229,N_11135);
nand U12532 (N_12532,N_11428,N_11366);
nor U12533 (N_12533,N_11414,N_11995);
nand U12534 (N_12534,N_11713,N_11648);
nor U12535 (N_12535,N_11535,N_11828);
or U12536 (N_12536,N_11960,N_11378);
nand U12537 (N_12537,N_11494,N_11654);
nor U12538 (N_12538,N_11637,N_11982);
nand U12539 (N_12539,N_11901,N_11601);
nand U12540 (N_12540,N_11325,N_11924);
nor U12541 (N_12541,N_11606,N_11017);
nor U12542 (N_12542,N_11612,N_11216);
and U12543 (N_12543,N_11041,N_11212);
or U12544 (N_12544,N_11050,N_11462);
nand U12545 (N_12545,N_11675,N_11907);
or U12546 (N_12546,N_11979,N_11085);
nand U12547 (N_12547,N_11351,N_11377);
nand U12548 (N_12548,N_11597,N_11425);
and U12549 (N_12549,N_11420,N_11805);
or U12550 (N_12550,N_11508,N_11966);
nor U12551 (N_12551,N_11606,N_11077);
or U12552 (N_12552,N_11066,N_11401);
or U12553 (N_12553,N_11595,N_11133);
nor U12554 (N_12554,N_11703,N_11892);
or U12555 (N_12555,N_11313,N_11765);
and U12556 (N_12556,N_11164,N_11839);
or U12557 (N_12557,N_11213,N_11628);
nor U12558 (N_12558,N_11081,N_11287);
or U12559 (N_12559,N_11902,N_11105);
nor U12560 (N_12560,N_11871,N_11244);
or U12561 (N_12561,N_11272,N_11228);
nor U12562 (N_12562,N_11782,N_11726);
nor U12563 (N_12563,N_11894,N_11438);
and U12564 (N_12564,N_11865,N_11566);
and U12565 (N_12565,N_11916,N_11020);
and U12566 (N_12566,N_11618,N_11629);
nand U12567 (N_12567,N_11916,N_11474);
and U12568 (N_12568,N_11021,N_11448);
nand U12569 (N_12569,N_11799,N_11204);
and U12570 (N_12570,N_11541,N_11105);
and U12571 (N_12571,N_11364,N_11573);
nor U12572 (N_12572,N_11378,N_11984);
or U12573 (N_12573,N_11609,N_11483);
nand U12574 (N_12574,N_11104,N_11040);
and U12575 (N_12575,N_11222,N_11764);
nor U12576 (N_12576,N_11788,N_11576);
or U12577 (N_12577,N_11107,N_11272);
and U12578 (N_12578,N_11719,N_11203);
nor U12579 (N_12579,N_11718,N_11037);
nor U12580 (N_12580,N_11162,N_11258);
nand U12581 (N_12581,N_11828,N_11862);
or U12582 (N_12582,N_11417,N_11994);
nand U12583 (N_12583,N_11325,N_11609);
and U12584 (N_12584,N_11866,N_11905);
nand U12585 (N_12585,N_11844,N_11122);
nor U12586 (N_12586,N_11890,N_11719);
and U12587 (N_12587,N_11627,N_11708);
nand U12588 (N_12588,N_11132,N_11310);
and U12589 (N_12589,N_11062,N_11347);
or U12590 (N_12590,N_11513,N_11672);
nor U12591 (N_12591,N_11666,N_11704);
nand U12592 (N_12592,N_11407,N_11755);
nand U12593 (N_12593,N_11774,N_11257);
nor U12594 (N_12594,N_11978,N_11892);
or U12595 (N_12595,N_11900,N_11295);
and U12596 (N_12596,N_11065,N_11924);
nor U12597 (N_12597,N_11263,N_11875);
nor U12598 (N_12598,N_11108,N_11577);
and U12599 (N_12599,N_11092,N_11590);
nand U12600 (N_12600,N_11043,N_11382);
nand U12601 (N_12601,N_11997,N_11409);
nand U12602 (N_12602,N_11461,N_11306);
and U12603 (N_12603,N_11680,N_11054);
or U12604 (N_12604,N_11389,N_11898);
nor U12605 (N_12605,N_11593,N_11877);
and U12606 (N_12606,N_11614,N_11696);
nor U12607 (N_12607,N_11830,N_11707);
and U12608 (N_12608,N_11374,N_11830);
nand U12609 (N_12609,N_11901,N_11142);
or U12610 (N_12610,N_11247,N_11398);
nand U12611 (N_12611,N_11291,N_11790);
and U12612 (N_12612,N_11764,N_11659);
nand U12613 (N_12613,N_11614,N_11375);
nor U12614 (N_12614,N_11949,N_11871);
and U12615 (N_12615,N_11250,N_11502);
or U12616 (N_12616,N_11299,N_11459);
nand U12617 (N_12617,N_11143,N_11828);
nor U12618 (N_12618,N_11694,N_11704);
nand U12619 (N_12619,N_11031,N_11959);
nand U12620 (N_12620,N_11281,N_11109);
nand U12621 (N_12621,N_11629,N_11650);
nor U12622 (N_12622,N_11242,N_11127);
or U12623 (N_12623,N_11213,N_11040);
nand U12624 (N_12624,N_11261,N_11434);
and U12625 (N_12625,N_11242,N_11064);
or U12626 (N_12626,N_11106,N_11999);
nor U12627 (N_12627,N_11407,N_11441);
nand U12628 (N_12628,N_11403,N_11860);
nor U12629 (N_12629,N_11233,N_11487);
and U12630 (N_12630,N_11257,N_11147);
and U12631 (N_12631,N_11147,N_11042);
or U12632 (N_12632,N_11394,N_11566);
nor U12633 (N_12633,N_11359,N_11047);
and U12634 (N_12634,N_11677,N_11003);
nor U12635 (N_12635,N_11090,N_11309);
or U12636 (N_12636,N_11959,N_11866);
and U12637 (N_12637,N_11636,N_11812);
nand U12638 (N_12638,N_11498,N_11682);
nor U12639 (N_12639,N_11504,N_11204);
or U12640 (N_12640,N_11328,N_11796);
nor U12641 (N_12641,N_11388,N_11479);
nand U12642 (N_12642,N_11614,N_11582);
or U12643 (N_12643,N_11919,N_11170);
nand U12644 (N_12644,N_11015,N_11421);
nand U12645 (N_12645,N_11859,N_11502);
or U12646 (N_12646,N_11035,N_11329);
nand U12647 (N_12647,N_11511,N_11954);
nor U12648 (N_12648,N_11825,N_11830);
nor U12649 (N_12649,N_11528,N_11403);
and U12650 (N_12650,N_11154,N_11491);
nand U12651 (N_12651,N_11979,N_11486);
nor U12652 (N_12652,N_11372,N_11137);
nand U12653 (N_12653,N_11234,N_11611);
and U12654 (N_12654,N_11936,N_11352);
nor U12655 (N_12655,N_11756,N_11383);
or U12656 (N_12656,N_11845,N_11144);
nor U12657 (N_12657,N_11663,N_11155);
and U12658 (N_12658,N_11571,N_11481);
nand U12659 (N_12659,N_11808,N_11843);
nor U12660 (N_12660,N_11474,N_11472);
nor U12661 (N_12661,N_11057,N_11686);
and U12662 (N_12662,N_11232,N_11956);
and U12663 (N_12663,N_11809,N_11334);
and U12664 (N_12664,N_11391,N_11468);
nand U12665 (N_12665,N_11869,N_11384);
nor U12666 (N_12666,N_11443,N_11585);
nand U12667 (N_12667,N_11673,N_11973);
nand U12668 (N_12668,N_11537,N_11461);
or U12669 (N_12669,N_11179,N_11014);
nand U12670 (N_12670,N_11666,N_11356);
or U12671 (N_12671,N_11023,N_11083);
and U12672 (N_12672,N_11907,N_11897);
and U12673 (N_12673,N_11224,N_11657);
nand U12674 (N_12674,N_11606,N_11086);
xnor U12675 (N_12675,N_11119,N_11956);
and U12676 (N_12676,N_11379,N_11936);
nor U12677 (N_12677,N_11535,N_11064);
and U12678 (N_12678,N_11301,N_11790);
nor U12679 (N_12679,N_11202,N_11624);
or U12680 (N_12680,N_11274,N_11031);
nor U12681 (N_12681,N_11301,N_11858);
nor U12682 (N_12682,N_11202,N_11890);
and U12683 (N_12683,N_11018,N_11768);
and U12684 (N_12684,N_11739,N_11120);
or U12685 (N_12685,N_11376,N_11945);
nand U12686 (N_12686,N_11521,N_11917);
and U12687 (N_12687,N_11801,N_11349);
nand U12688 (N_12688,N_11171,N_11747);
and U12689 (N_12689,N_11203,N_11168);
or U12690 (N_12690,N_11204,N_11495);
nand U12691 (N_12691,N_11757,N_11875);
nor U12692 (N_12692,N_11326,N_11238);
or U12693 (N_12693,N_11594,N_11478);
nand U12694 (N_12694,N_11827,N_11630);
nor U12695 (N_12695,N_11688,N_11236);
nor U12696 (N_12696,N_11280,N_11222);
nor U12697 (N_12697,N_11479,N_11761);
and U12698 (N_12698,N_11888,N_11702);
nand U12699 (N_12699,N_11781,N_11579);
nor U12700 (N_12700,N_11693,N_11984);
xor U12701 (N_12701,N_11284,N_11775);
and U12702 (N_12702,N_11424,N_11791);
or U12703 (N_12703,N_11077,N_11797);
nor U12704 (N_12704,N_11310,N_11841);
or U12705 (N_12705,N_11193,N_11976);
or U12706 (N_12706,N_11185,N_11450);
or U12707 (N_12707,N_11070,N_11864);
nand U12708 (N_12708,N_11549,N_11597);
or U12709 (N_12709,N_11893,N_11102);
or U12710 (N_12710,N_11555,N_11783);
or U12711 (N_12711,N_11563,N_11903);
nand U12712 (N_12712,N_11770,N_11298);
nand U12713 (N_12713,N_11522,N_11219);
nand U12714 (N_12714,N_11375,N_11090);
nor U12715 (N_12715,N_11658,N_11143);
nand U12716 (N_12716,N_11006,N_11042);
and U12717 (N_12717,N_11490,N_11860);
or U12718 (N_12718,N_11968,N_11020);
nor U12719 (N_12719,N_11172,N_11357);
nor U12720 (N_12720,N_11202,N_11583);
nor U12721 (N_12721,N_11616,N_11534);
and U12722 (N_12722,N_11042,N_11957);
nand U12723 (N_12723,N_11041,N_11598);
or U12724 (N_12724,N_11990,N_11478);
and U12725 (N_12725,N_11055,N_11835);
nor U12726 (N_12726,N_11686,N_11951);
nand U12727 (N_12727,N_11873,N_11528);
nor U12728 (N_12728,N_11058,N_11364);
nand U12729 (N_12729,N_11507,N_11892);
and U12730 (N_12730,N_11981,N_11179);
nand U12731 (N_12731,N_11853,N_11567);
and U12732 (N_12732,N_11808,N_11756);
or U12733 (N_12733,N_11196,N_11023);
and U12734 (N_12734,N_11723,N_11088);
or U12735 (N_12735,N_11377,N_11531);
nor U12736 (N_12736,N_11685,N_11406);
or U12737 (N_12737,N_11988,N_11394);
nor U12738 (N_12738,N_11338,N_11666);
and U12739 (N_12739,N_11808,N_11540);
nor U12740 (N_12740,N_11626,N_11599);
and U12741 (N_12741,N_11484,N_11360);
nor U12742 (N_12742,N_11382,N_11371);
xnor U12743 (N_12743,N_11615,N_11702);
or U12744 (N_12744,N_11977,N_11564);
nand U12745 (N_12745,N_11818,N_11627);
or U12746 (N_12746,N_11855,N_11829);
nor U12747 (N_12747,N_11313,N_11825);
or U12748 (N_12748,N_11050,N_11107);
nor U12749 (N_12749,N_11938,N_11298);
or U12750 (N_12750,N_11783,N_11945);
or U12751 (N_12751,N_11266,N_11244);
nand U12752 (N_12752,N_11015,N_11678);
or U12753 (N_12753,N_11683,N_11418);
nand U12754 (N_12754,N_11382,N_11673);
nand U12755 (N_12755,N_11173,N_11859);
or U12756 (N_12756,N_11917,N_11431);
and U12757 (N_12757,N_11527,N_11584);
nand U12758 (N_12758,N_11747,N_11996);
nand U12759 (N_12759,N_11740,N_11988);
nor U12760 (N_12760,N_11549,N_11813);
nand U12761 (N_12761,N_11758,N_11933);
or U12762 (N_12762,N_11525,N_11100);
and U12763 (N_12763,N_11316,N_11936);
and U12764 (N_12764,N_11311,N_11177);
nor U12765 (N_12765,N_11977,N_11036);
and U12766 (N_12766,N_11879,N_11699);
or U12767 (N_12767,N_11362,N_11411);
nand U12768 (N_12768,N_11941,N_11094);
nand U12769 (N_12769,N_11616,N_11953);
or U12770 (N_12770,N_11641,N_11095);
nand U12771 (N_12771,N_11409,N_11636);
nand U12772 (N_12772,N_11296,N_11327);
nor U12773 (N_12773,N_11094,N_11821);
and U12774 (N_12774,N_11808,N_11600);
nor U12775 (N_12775,N_11586,N_11116);
nand U12776 (N_12776,N_11212,N_11721);
nand U12777 (N_12777,N_11344,N_11565);
nor U12778 (N_12778,N_11018,N_11070);
nor U12779 (N_12779,N_11806,N_11487);
nand U12780 (N_12780,N_11242,N_11784);
xnor U12781 (N_12781,N_11281,N_11074);
nor U12782 (N_12782,N_11733,N_11115);
nand U12783 (N_12783,N_11546,N_11508);
nand U12784 (N_12784,N_11083,N_11094);
nand U12785 (N_12785,N_11338,N_11772);
nor U12786 (N_12786,N_11678,N_11244);
nor U12787 (N_12787,N_11965,N_11928);
and U12788 (N_12788,N_11571,N_11838);
nand U12789 (N_12789,N_11212,N_11315);
and U12790 (N_12790,N_11278,N_11867);
or U12791 (N_12791,N_11092,N_11979);
nand U12792 (N_12792,N_11067,N_11459);
and U12793 (N_12793,N_11347,N_11752);
and U12794 (N_12794,N_11538,N_11015);
or U12795 (N_12795,N_11440,N_11839);
or U12796 (N_12796,N_11078,N_11037);
and U12797 (N_12797,N_11618,N_11045);
nand U12798 (N_12798,N_11248,N_11207);
and U12799 (N_12799,N_11040,N_11485);
nand U12800 (N_12800,N_11021,N_11085);
or U12801 (N_12801,N_11597,N_11635);
or U12802 (N_12802,N_11735,N_11189);
nand U12803 (N_12803,N_11708,N_11203);
or U12804 (N_12804,N_11563,N_11785);
or U12805 (N_12805,N_11858,N_11981);
nand U12806 (N_12806,N_11765,N_11919);
nor U12807 (N_12807,N_11148,N_11077);
nor U12808 (N_12808,N_11657,N_11839);
nand U12809 (N_12809,N_11740,N_11653);
nor U12810 (N_12810,N_11033,N_11054);
and U12811 (N_12811,N_11458,N_11171);
nor U12812 (N_12812,N_11882,N_11134);
nand U12813 (N_12813,N_11451,N_11586);
and U12814 (N_12814,N_11209,N_11212);
and U12815 (N_12815,N_11811,N_11364);
nand U12816 (N_12816,N_11314,N_11137);
nor U12817 (N_12817,N_11641,N_11694);
nand U12818 (N_12818,N_11685,N_11014);
nand U12819 (N_12819,N_11727,N_11004);
nand U12820 (N_12820,N_11252,N_11709);
nand U12821 (N_12821,N_11513,N_11096);
and U12822 (N_12822,N_11093,N_11182);
or U12823 (N_12823,N_11893,N_11848);
nor U12824 (N_12824,N_11547,N_11074);
and U12825 (N_12825,N_11815,N_11942);
nor U12826 (N_12826,N_11846,N_11384);
nand U12827 (N_12827,N_11206,N_11997);
nand U12828 (N_12828,N_11477,N_11550);
nand U12829 (N_12829,N_11624,N_11472);
nor U12830 (N_12830,N_11190,N_11622);
and U12831 (N_12831,N_11581,N_11393);
or U12832 (N_12832,N_11568,N_11886);
or U12833 (N_12833,N_11697,N_11774);
and U12834 (N_12834,N_11605,N_11191);
or U12835 (N_12835,N_11351,N_11800);
and U12836 (N_12836,N_11933,N_11905);
and U12837 (N_12837,N_11316,N_11874);
and U12838 (N_12838,N_11704,N_11103);
or U12839 (N_12839,N_11032,N_11793);
nand U12840 (N_12840,N_11599,N_11888);
nor U12841 (N_12841,N_11200,N_11178);
and U12842 (N_12842,N_11723,N_11704);
or U12843 (N_12843,N_11419,N_11519);
and U12844 (N_12844,N_11724,N_11526);
nand U12845 (N_12845,N_11871,N_11465);
nor U12846 (N_12846,N_11333,N_11529);
nand U12847 (N_12847,N_11935,N_11651);
nor U12848 (N_12848,N_11285,N_11784);
and U12849 (N_12849,N_11902,N_11116);
or U12850 (N_12850,N_11650,N_11804);
or U12851 (N_12851,N_11192,N_11964);
nor U12852 (N_12852,N_11854,N_11165);
nor U12853 (N_12853,N_11219,N_11340);
and U12854 (N_12854,N_11586,N_11944);
nor U12855 (N_12855,N_11145,N_11093);
nor U12856 (N_12856,N_11241,N_11526);
nand U12857 (N_12857,N_11679,N_11643);
nand U12858 (N_12858,N_11620,N_11846);
nand U12859 (N_12859,N_11733,N_11417);
nand U12860 (N_12860,N_11178,N_11674);
or U12861 (N_12861,N_11588,N_11452);
or U12862 (N_12862,N_11869,N_11945);
nor U12863 (N_12863,N_11408,N_11433);
or U12864 (N_12864,N_11603,N_11693);
and U12865 (N_12865,N_11863,N_11345);
and U12866 (N_12866,N_11475,N_11157);
and U12867 (N_12867,N_11285,N_11081);
or U12868 (N_12868,N_11234,N_11422);
or U12869 (N_12869,N_11887,N_11385);
or U12870 (N_12870,N_11438,N_11841);
or U12871 (N_12871,N_11935,N_11646);
and U12872 (N_12872,N_11824,N_11285);
nor U12873 (N_12873,N_11081,N_11877);
nor U12874 (N_12874,N_11139,N_11290);
and U12875 (N_12875,N_11427,N_11008);
and U12876 (N_12876,N_11694,N_11919);
and U12877 (N_12877,N_11246,N_11711);
nand U12878 (N_12878,N_11878,N_11554);
and U12879 (N_12879,N_11970,N_11247);
and U12880 (N_12880,N_11360,N_11615);
nand U12881 (N_12881,N_11139,N_11042);
nor U12882 (N_12882,N_11465,N_11584);
or U12883 (N_12883,N_11091,N_11230);
and U12884 (N_12884,N_11476,N_11234);
or U12885 (N_12885,N_11421,N_11046);
nand U12886 (N_12886,N_11261,N_11946);
or U12887 (N_12887,N_11361,N_11600);
and U12888 (N_12888,N_11729,N_11523);
and U12889 (N_12889,N_11209,N_11422);
nand U12890 (N_12890,N_11424,N_11743);
nand U12891 (N_12891,N_11884,N_11545);
or U12892 (N_12892,N_11994,N_11038);
nor U12893 (N_12893,N_11894,N_11962);
nand U12894 (N_12894,N_11106,N_11226);
and U12895 (N_12895,N_11131,N_11685);
nor U12896 (N_12896,N_11509,N_11325);
and U12897 (N_12897,N_11827,N_11194);
nor U12898 (N_12898,N_11349,N_11646);
or U12899 (N_12899,N_11301,N_11970);
or U12900 (N_12900,N_11061,N_11560);
xor U12901 (N_12901,N_11758,N_11250);
nand U12902 (N_12902,N_11380,N_11622);
nand U12903 (N_12903,N_11319,N_11401);
and U12904 (N_12904,N_11749,N_11032);
nand U12905 (N_12905,N_11882,N_11190);
and U12906 (N_12906,N_11279,N_11830);
nor U12907 (N_12907,N_11159,N_11904);
and U12908 (N_12908,N_11653,N_11845);
and U12909 (N_12909,N_11570,N_11463);
nand U12910 (N_12910,N_11173,N_11724);
or U12911 (N_12911,N_11899,N_11102);
or U12912 (N_12912,N_11937,N_11764);
nand U12913 (N_12913,N_11150,N_11470);
and U12914 (N_12914,N_11450,N_11273);
nor U12915 (N_12915,N_11311,N_11039);
nor U12916 (N_12916,N_11990,N_11002);
nand U12917 (N_12917,N_11406,N_11897);
or U12918 (N_12918,N_11275,N_11666);
nor U12919 (N_12919,N_11984,N_11109);
and U12920 (N_12920,N_11758,N_11762);
and U12921 (N_12921,N_11767,N_11855);
and U12922 (N_12922,N_11210,N_11330);
nand U12923 (N_12923,N_11201,N_11898);
and U12924 (N_12924,N_11294,N_11014);
or U12925 (N_12925,N_11321,N_11102);
nor U12926 (N_12926,N_11637,N_11415);
nand U12927 (N_12927,N_11225,N_11744);
nor U12928 (N_12928,N_11474,N_11792);
or U12929 (N_12929,N_11050,N_11898);
or U12930 (N_12930,N_11842,N_11382);
or U12931 (N_12931,N_11701,N_11595);
and U12932 (N_12932,N_11357,N_11296);
and U12933 (N_12933,N_11445,N_11746);
nor U12934 (N_12934,N_11727,N_11994);
nor U12935 (N_12935,N_11705,N_11853);
or U12936 (N_12936,N_11350,N_11125);
nand U12937 (N_12937,N_11888,N_11812);
or U12938 (N_12938,N_11997,N_11332);
nand U12939 (N_12939,N_11083,N_11727);
or U12940 (N_12940,N_11960,N_11260);
nand U12941 (N_12941,N_11947,N_11593);
nand U12942 (N_12942,N_11070,N_11926);
nand U12943 (N_12943,N_11949,N_11554);
nand U12944 (N_12944,N_11750,N_11386);
nand U12945 (N_12945,N_11093,N_11715);
xor U12946 (N_12946,N_11029,N_11855);
and U12947 (N_12947,N_11255,N_11879);
nand U12948 (N_12948,N_11117,N_11080);
or U12949 (N_12949,N_11571,N_11194);
nand U12950 (N_12950,N_11262,N_11258);
or U12951 (N_12951,N_11916,N_11783);
and U12952 (N_12952,N_11063,N_11426);
and U12953 (N_12953,N_11122,N_11905);
and U12954 (N_12954,N_11943,N_11255);
nand U12955 (N_12955,N_11157,N_11019);
nor U12956 (N_12956,N_11686,N_11558);
nor U12957 (N_12957,N_11703,N_11097);
and U12958 (N_12958,N_11131,N_11077);
nand U12959 (N_12959,N_11633,N_11003);
or U12960 (N_12960,N_11039,N_11014);
and U12961 (N_12961,N_11165,N_11468);
nor U12962 (N_12962,N_11698,N_11103);
and U12963 (N_12963,N_11052,N_11852);
or U12964 (N_12964,N_11257,N_11378);
nor U12965 (N_12965,N_11989,N_11265);
and U12966 (N_12966,N_11340,N_11381);
nand U12967 (N_12967,N_11905,N_11304);
or U12968 (N_12968,N_11454,N_11143);
nand U12969 (N_12969,N_11350,N_11454);
nand U12970 (N_12970,N_11528,N_11939);
nand U12971 (N_12971,N_11503,N_11017);
nor U12972 (N_12972,N_11093,N_11051);
nand U12973 (N_12973,N_11494,N_11901);
or U12974 (N_12974,N_11469,N_11446);
nand U12975 (N_12975,N_11190,N_11883);
or U12976 (N_12976,N_11387,N_11359);
or U12977 (N_12977,N_11082,N_11803);
nor U12978 (N_12978,N_11679,N_11299);
and U12979 (N_12979,N_11013,N_11470);
nor U12980 (N_12980,N_11599,N_11515);
and U12981 (N_12981,N_11187,N_11327);
nand U12982 (N_12982,N_11709,N_11569);
nor U12983 (N_12983,N_11938,N_11892);
nand U12984 (N_12984,N_11669,N_11186);
and U12985 (N_12985,N_11073,N_11465);
or U12986 (N_12986,N_11713,N_11916);
and U12987 (N_12987,N_11404,N_11608);
nor U12988 (N_12988,N_11594,N_11439);
nor U12989 (N_12989,N_11114,N_11203);
nand U12990 (N_12990,N_11161,N_11745);
nand U12991 (N_12991,N_11486,N_11874);
or U12992 (N_12992,N_11206,N_11712);
and U12993 (N_12993,N_11109,N_11036);
nor U12994 (N_12994,N_11915,N_11636);
nor U12995 (N_12995,N_11049,N_11146);
nor U12996 (N_12996,N_11467,N_11000);
or U12997 (N_12997,N_11181,N_11492);
and U12998 (N_12998,N_11945,N_11186);
nor U12999 (N_12999,N_11645,N_11339);
nand U13000 (N_13000,N_12968,N_12542);
nor U13001 (N_13001,N_12137,N_12430);
nand U13002 (N_13002,N_12153,N_12801);
nor U13003 (N_13003,N_12289,N_12491);
xor U13004 (N_13004,N_12680,N_12477);
nor U13005 (N_13005,N_12252,N_12171);
nor U13006 (N_13006,N_12300,N_12657);
and U13007 (N_13007,N_12602,N_12872);
nor U13008 (N_13008,N_12148,N_12178);
nand U13009 (N_13009,N_12395,N_12995);
or U13010 (N_13010,N_12926,N_12596);
or U13011 (N_13011,N_12907,N_12794);
nand U13012 (N_13012,N_12412,N_12514);
nor U13013 (N_13013,N_12301,N_12941);
nand U13014 (N_13014,N_12690,N_12584);
and U13015 (N_13015,N_12188,N_12822);
or U13016 (N_13016,N_12123,N_12319);
and U13017 (N_13017,N_12746,N_12292);
nand U13018 (N_13018,N_12219,N_12670);
or U13019 (N_13019,N_12362,N_12259);
nor U13020 (N_13020,N_12607,N_12428);
nor U13021 (N_13021,N_12321,N_12250);
nor U13022 (N_13022,N_12504,N_12421);
and U13023 (N_13023,N_12278,N_12061);
or U13024 (N_13024,N_12515,N_12048);
nor U13025 (N_13025,N_12356,N_12106);
nor U13026 (N_13026,N_12672,N_12826);
nor U13027 (N_13027,N_12285,N_12162);
or U13028 (N_13028,N_12627,N_12629);
and U13029 (N_13029,N_12128,N_12913);
nand U13030 (N_13030,N_12409,N_12336);
or U13031 (N_13031,N_12823,N_12540);
or U13032 (N_13032,N_12732,N_12483);
and U13033 (N_13033,N_12223,N_12811);
and U13034 (N_13034,N_12817,N_12979);
and U13035 (N_13035,N_12875,N_12070);
and U13036 (N_13036,N_12551,N_12844);
or U13037 (N_13037,N_12177,N_12677);
and U13038 (N_13038,N_12367,N_12924);
nand U13039 (N_13039,N_12685,N_12029);
nor U13040 (N_13040,N_12282,N_12835);
and U13041 (N_13041,N_12699,N_12803);
or U13042 (N_13042,N_12156,N_12740);
and U13043 (N_13043,N_12813,N_12195);
and U13044 (N_13044,N_12674,N_12098);
nand U13045 (N_13045,N_12706,N_12444);
or U13046 (N_13046,N_12897,N_12807);
or U13047 (N_13047,N_12933,N_12182);
and U13048 (N_13048,N_12091,N_12563);
and U13049 (N_13049,N_12217,N_12088);
nor U13050 (N_13050,N_12829,N_12735);
or U13051 (N_13051,N_12538,N_12325);
nor U13052 (N_13052,N_12304,N_12097);
nor U13053 (N_13053,N_12727,N_12454);
nand U13054 (N_13054,N_12111,N_12914);
nor U13055 (N_13055,N_12413,N_12272);
or U13056 (N_13056,N_12068,N_12274);
or U13057 (N_13057,N_12470,N_12669);
nand U13058 (N_13058,N_12372,N_12013);
nand U13059 (N_13059,N_12196,N_12185);
nor U13060 (N_13060,N_12728,N_12648);
and U13061 (N_13061,N_12764,N_12722);
nor U13062 (N_13062,N_12134,N_12556);
nor U13063 (N_13063,N_12125,N_12855);
nand U13064 (N_13064,N_12131,N_12917);
nand U13065 (N_13065,N_12534,N_12056);
and U13066 (N_13066,N_12838,N_12908);
nor U13067 (N_13067,N_12560,N_12512);
and U13068 (N_13068,N_12054,N_12756);
or U13069 (N_13069,N_12353,N_12998);
nor U13070 (N_13070,N_12885,N_12475);
and U13071 (N_13071,N_12473,N_12346);
and U13072 (N_13072,N_12757,N_12206);
and U13073 (N_13073,N_12574,N_12856);
and U13074 (N_13074,N_12634,N_12696);
nand U13075 (N_13075,N_12624,N_12681);
or U13076 (N_13076,N_12264,N_12120);
nor U13077 (N_13077,N_12022,N_12805);
nand U13078 (N_13078,N_12752,N_12199);
or U13079 (N_13079,N_12451,N_12558);
nor U13080 (N_13080,N_12643,N_12239);
or U13081 (N_13081,N_12482,N_12167);
nor U13082 (N_13082,N_12406,N_12783);
or U13083 (N_13083,N_12378,N_12373);
and U13084 (N_13084,N_12456,N_12880);
nand U13085 (N_13085,N_12291,N_12474);
nand U13086 (N_13086,N_12768,N_12047);
xor U13087 (N_13087,N_12932,N_12407);
nand U13088 (N_13088,N_12956,N_12002);
or U13089 (N_13089,N_12041,N_12747);
and U13090 (N_13090,N_12782,N_12572);
nor U13091 (N_13091,N_12849,N_12647);
and U13092 (N_13092,N_12268,N_12126);
nand U13093 (N_13093,N_12711,N_12507);
and U13094 (N_13094,N_12186,N_12969);
nand U13095 (N_13095,N_12307,N_12775);
nand U13096 (N_13096,N_12149,N_12600);
and U13097 (N_13097,N_12493,N_12820);
nand U13098 (N_13098,N_12737,N_12626);
nor U13099 (N_13099,N_12092,N_12592);
nand U13100 (N_13100,N_12469,N_12462);
nor U13101 (N_13101,N_12175,N_12094);
or U13102 (N_13102,N_12520,N_12074);
or U13103 (N_13103,N_12270,N_12038);
and U13104 (N_13104,N_12508,N_12889);
or U13105 (N_13105,N_12967,N_12492);
nor U13106 (N_13106,N_12539,N_12610);
nand U13107 (N_13107,N_12638,N_12343);
or U13108 (N_13108,N_12121,N_12990);
or U13109 (N_13109,N_12116,N_12400);
or U13110 (N_13110,N_12734,N_12511);
nor U13111 (N_13111,N_12093,N_12103);
or U13112 (N_13112,N_12915,N_12667);
and U13113 (N_13113,N_12637,N_12450);
and U13114 (N_13114,N_12389,N_12609);
or U13115 (N_13115,N_12874,N_12526);
and U13116 (N_13116,N_12050,N_12011);
nor U13117 (N_13117,N_12881,N_12553);
nand U13118 (N_13118,N_12916,N_12973);
nor U13119 (N_13119,N_12843,N_12877);
nand U13120 (N_13120,N_12615,N_12155);
nor U13121 (N_13121,N_12139,N_12345);
nor U13122 (N_13122,N_12660,N_12385);
nor U13123 (N_13123,N_12383,N_12774);
and U13124 (N_13124,N_12950,N_12903);
or U13125 (N_13125,N_12057,N_12927);
and U13126 (N_13126,N_12608,N_12957);
and U13127 (N_13127,N_12159,N_12871);
nand U13128 (N_13128,N_12955,N_12790);
and U13129 (N_13129,N_12277,N_12851);
or U13130 (N_13130,N_12682,N_12815);
or U13131 (N_13131,N_12623,N_12831);
or U13132 (N_13132,N_12890,N_12891);
and U13133 (N_13133,N_12810,N_12145);
and U13134 (N_13134,N_12036,N_12187);
nor U13135 (N_13135,N_12433,N_12459);
and U13136 (N_13136,N_12724,N_12380);
nor U13137 (N_13137,N_12308,N_12117);
nor U13138 (N_13138,N_12401,N_12840);
nand U13139 (N_13139,N_12611,N_12240);
or U13140 (N_13140,N_12269,N_12224);
nand U13141 (N_13141,N_12310,N_12369);
nand U13142 (N_13142,N_12163,N_12288);
nor U13143 (N_13143,N_12925,N_12287);
nor U13144 (N_13144,N_12316,N_12295);
or U13145 (N_13145,N_12644,N_12537);
nand U13146 (N_13146,N_12772,N_12020);
or U13147 (N_13147,N_12220,N_12000);
nand U13148 (N_13148,N_12144,N_12530);
or U13149 (N_13149,N_12987,N_12415);
and U13150 (N_13150,N_12158,N_12639);
or U13151 (N_13151,N_12312,N_12427);
nand U13152 (N_13152,N_12854,N_12435);
nand U13153 (N_13153,N_12693,N_12205);
or U13154 (N_13154,N_12332,N_12049);
nor U13155 (N_13155,N_12652,N_12582);
and U13156 (N_13156,N_12096,N_12464);
nor U13157 (N_13157,N_12500,N_12222);
nor U13158 (N_13158,N_12429,N_12231);
or U13159 (N_13159,N_12816,N_12870);
nand U13160 (N_13160,N_12276,N_12241);
or U13161 (N_13161,N_12620,N_12730);
nor U13162 (N_13162,N_12920,N_12254);
and U13163 (N_13163,N_12005,N_12883);
nand U13164 (N_13164,N_12510,N_12731);
or U13165 (N_13165,N_12351,N_12953);
nand U13166 (N_13166,N_12418,N_12494);
nand U13167 (N_13167,N_12168,N_12804);
or U13168 (N_13168,N_12410,N_12958);
or U13169 (N_13169,N_12065,N_12830);
and U13170 (N_13170,N_12705,N_12069);
and U13171 (N_13171,N_12760,N_12991);
and U13172 (N_13172,N_12478,N_12806);
or U13173 (N_13173,N_12497,N_12296);
nand U13174 (N_13174,N_12115,N_12550);
nand U13175 (N_13175,N_12867,N_12328);
nand U13176 (N_13176,N_12853,N_12232);
nor U13177 (N_13177,N_12850,N_12651);
or U13178 (N_13178,N_12053,N_12960);
or U13179 (N_13179,N_12800,N_12824);
nor U13180 (N_13180,N_12524,N_12702);
nor U13181 (N_13181,N_12320,N_12382);
nand U13182 (N_13182,N_12181,N_12073);
nand U13183 (N_13183,N_12247,N_12084);
and U13184 (N_13184,N_12785,N_12063);
nand U13185 (N_13185,N_12748,N_12173);
nor U13186 (N_13186,N_12703,N_12951);
and U13187 (N_13187,N_12911,N_12329);
nand U13188 (N_13188,N_12857,N_12654);
or U13189 (N_13189,N_12448,N_12212);
nand U13190 (N_13190,N_12588,N_12388);
or U13191 (N_13191,N_12442,N_12165);
or U13192 (N_13192,N_12939,N_12845);
nor U13193 (N_13193,N_12778,N_12355);
and U13194 (N_13194,N_12019,N_12255);
nand U13195 (N_13195,N_12026,N_12081);
or U13196 (N_13196,N_12846,N_12359);
or U13197 (N_13197,N_12993,N_12837);
nand U13198 (N_13198,N_12770,N_12243);
and U13199 (N_13199,N_12513,N_12621);
nor U13200 (N_13200,N_12496,N_12244);
nand U13201 (N_13201,N_12566,N_12438);
or U13202 (N_13202,N_12034,N_12306);
and U13203 (N_13203,N_12318,N_12204);
or U13204 (N_13204,N_12922,N_12899);
or U13205 (N_13205,N_12625,N_12888);
or U13206 (N_13206,N_12402,N_12398);
or U13207 (N_13207,N_12327,N_12150);
nand U13208 (N_13208,N_12417,N_12863);
nor U13209 (N_13209,N_12315,N_12619);
and U13210 (N_13210,N_12436,N_12503);
and U13211 (N_13211,N_12324,N_12750);
nor U13212 (N_13212,N_12980,N_12142);
nand U13213 (N_13213,N_12586,N_12309);
nand U13214 (N_13214,N_12839,N_12909);
and U13215 (N_13215,N_12700,N_12051);
or U13216 (N_13216,N_12635,N_12501);
nand U13217 (N_13217,N_12640,N_12758);
nor U13218 (N_13218,N_12368,N_12465);
or U13219 (N_13219,N_12738,N_12910);
or U13220 (N_13220,N_12802,N_12339);
nor U13221 (N_13221,N_12593,N_12229);
nor U13222 (N_13222,N_12422,N_12555);
and U13223 (N_13223,N_12697,N_12233);
or U13224 (N_13224,N_12719,N_12630);
or U13225 (N_13225,N_12197,N_12604);
and U13226 (N_13226,N_12010,N_12227);
and U13227 (N_13227,N_12860,N_12425);
and U13228 (N_13228,N_12691,N_12921);
nand U13229 (N_13229,N_12532,N_12605);
or U13230 (N_13230,N_12527,N_12426);
or U13231 (N_13231,N_12234,N_12201);
and U13232 (N_13232,N_12789,N_12656);
nor U13233 (N_13233,N_12403,N_12387);
nand U13234 (N_13234,N_12864,N_12808);
nor U13235 (N_13235,N_12873,N_12357);
or U13236 (N_13236,N_12594,N_12058);
or U13237 (N_13237,N_12379,N_12257);
or U13238 (N_13238,N_12313,N_12251);
and U13239 (N_13239,N_12718,N_12330);
or U13240 (N_13240,N_12467,N_12266);
or U13241 (N_13241,N_12107,N_12970);
or U13242 (N_13242,N_12432,N_12761);
and U13243 (N_13243,N_12210,N_12076);
nor U13244 (N_13244,N_12363,N_12848);
or U13245 (N_13245,N_12606,N_12876);
or U13246 (N_13246,N_12636,N_12841);
or U13247 (N_13247,N_12564,N_12420);
or U13248 (N_13248,N_12544,N_12267);
and U13249 (N_13249,N_12027,N_12271);
or U13250 (N_13250,N_12568,N_12008);
and U13251 (N_13251,N_12253,N_12777);
nand U13252 (N_13252,N_12687,N_12906);
nor U13253 (N_13253,N_12533,N_12009);
nand U13254 (N_13254,N_12505,N_12384);
nor U13255 (N_13255,N_12161,N_12381);
nand U13256 (N_13256,N_12791,N_12988);
nand U13257 (N_13257,N_12715,N_12795);
nand U13258 (N_13258,N_12089,N_12834);
nand U13259 (N_13259,N_12443,N_12392);
nand U13260 (N_13260,N_12930,N_12007);
or U13261 (N_13261,N_12982,N_12095);
nand U13262 (N_13262,N_12653,N_12959);
nand U13263 (N_13263,N_12689,N_12112);
or U13264 (N_13264,N_12543,N_12003);
nor U13265 (N_13265,N_12366,N_12974);
nand U13266 (N_13266,N_12631,N_12561);
or U13267 (N_13267,N_12509,N_12323);
nand U13268 (N_13268,N_12157,N_12179);
and U13269 (N_13269,N_12552,N_12242);
and U13270 (N_13270,N_12546,N_12136);
nor U13271 (N_13271,N_12215,N_12683);
nor U13272 (N_13272,N_12799,N_12570);
or U13273 (N_13273,N_12894,N_12765);
and U13274 (N_13274,N_12023,N_12447);
and U13275 (N_13275,N_12248,N_12776);
nor U13276 (N_13276,N_12595,N_12338);
or U13277 (N_13277,N_12754,N_12064);
nor U13278 (N_13278,N_12893,N_12461);
or U13279 (N_13279,N_12071,N_12079);
nand U13280 (N_13280,N_12225,N_12599);
nand U13281 (N_13281,N_12203,N_12869);
and U13282 (N_13282,N_12040,N_12557);
nor U13283 (N_13283,N_12518,N_12997);
and U13284 (N_13284,N_12391,N_12286);
nor U13285 (N_13285,N_12337,N_12457);
and U13286 (N_13286,N_12684,N_12166);
or U13287 (N_13287,N_12714,N_12302);
or U13288 (N_13288,N_12226,N_12878);
or U13289 (N_13289,N_12273,N_12755);
nand U13290 (N_13290,N_12613,N_12085);
nor U13291 (N_13291,N_12364,N_12836);
nand U13292 (N_13292,N_12441,N_12938);
nor U13293 (N_13293,N_12937,N_12127);
and U13294 (N_13294,N_12018,N_12487);
or U13295 (N_13295,N_12349,N_12581);
xor U13296 (N_13296,N_12374,N_12996);
nand U13297 (N_13297,N_12531,N_12169);
or U13298 (N_13298,N_12726,N_12779);
nand U13299 (N_13299,N_12549,N_12039);
nand U13300 (N_13300,N_12375,N_12675);
and U13301 (N_13301,N_12119,N_12460);
nand U13302 (N_13302,N_12386,N_12122);
nor U13303 (N_13303,N_12587,N_12463);
or U13304 (N_13304,N_12942,N_12172);
nor U13305 (N_13305,N_12246,N_12024);
nor U13306 (N_13306,N_12245,N_12861);
nand U13307 (N_13307,N_12954,N_12440);
nor U13308 (N_13308,N_12796,N_12275);
and U13309 (N_13309,N_12192,N_12265);
nor U13310 (N_13310,N_12102,N_12110);
and U13311 (N_13311,N_12439,N_12124);
nor U13312 (N_13312,N_12347,N_12773);
or U13313 (N_13313,N_12214,N_12646);
or U13314 (N_13314,N_12046,N_12965);
or U13315 (N_13315,N_12305,N_12725);
nand U13316 (N_13316,N_12390,N_12101);
nand U13317 (N_13317,N_12576,N_12342);
nor U13318 (N_13318,N_12723,N_12739);
and U13319 (N_13319,N_12590,N_12742);
and U13320 (N_13320,N_12698,N_12879);
nor U13321 (N_13321,N_12695,N_12832);
nor U13322 (N_13322,N_12209,N_12499);
nor U13323 (N_13323,N_12704,N_12299);
nand U13324 (N_13324,N_12075,N_12340);
nor U13325 (N_13325,N_12281,N_12238);
and U13326 (N_13326,N_12862,N_12912);
or U13327 (N_13327,N_12666,N_12376);
xor U13328 (N_13328,N_12283,N_12668);
or U13329 (N_13329,N_12946,N_12350);
nand U13330 (N_13330,N_12180,N_12404);
and U13331 (N_13331,N_12978,N_12710);
nor U13332 (N_13332,N_12377,N_12825);
nor U13333 (N_13333,N_12614,N_12536);
and U13334 (N_13334,N_12781,N_12445);
or U13335 (N_13335,N_12506,N_12972);
and U13336 (N_13336,N_12692,N_12521);
nand U13337 (N_13337,N_12480,N_12080);
nor U13338 (N_13338,N_12154,N_12977);
nand U13339 (N_13339,N_12671,N_12601);
nor U13340 (N_13340,N_12847,N_12767);
or U13341 (N_13341,N_12658,N_12143);
nand U13342 (N_13342,N_12498,N_12709);
nand U13343 (N_13343,N_12567,N_12628);
nor U13344 (N_13344,N_12676,N_12371);
nor U13345 (N_13345,N_12458,N_12033);
nor U13346 (N_13346,N_12529,N_12228);
and U13347 (N_13347,N_12736,N_12519);
nand U13348 (N_13348,N_12293,N_12769);
nor U13349 (N_13349,N_12940,N_12297);
xnor U13350 (N_13350,N_12397,N_12230);
and U13351 (N_13351,N_12753,N_12842);
nand U13352 (N_13352,N_12025,N_12455);
and U13353 (N_13353,N_12017,N_12617);
xor U13354 (N_13354,N_12331,N_12109);
nor U13355 (N_13355,N_12200,N_12612);
nand U13356 (N_13356,N_12784,N_12446);
or U13357 (N_13357,N_12066,N_12100);
or U13358 (N_13358,N_12659,N_12334);
and U13359 (N_13359,N_12986,N_12135);
nand U13360 (N_13360,N_12408,N_12424);
nand U13361 (N_13361,N_12202,N_12211);
nand U13362 (N_13362,N_12035,N_12798);
nor U13363 (N_13363,N_12716,N_12964);
nor U13364 (N_13364,N_12792,N_12189);
and U13365 (N_13365,N_12701,N_12882);
and U13366 (N_13366,N_12661,N_12140);
nand U13367 (N_13367,N_12004,N_12999);
nor U13368 (N_13368,N_12216,N_12597);
xor U13369 (N_13369,N_12006,N_12213);
or U13370 (N_13370,N_12260,N_12087);
nor U13371 (N_13371,N_12522,N_12559);
and U13372 (N_13372,N_12618,N_12062);
or U13373 (N_13373,N_12745,N_12453);
and U13374 (N_13374,N_12868,N_12502);
xor U13375 (N_13375,N_12983,N_12749);
or U13376 (N_13376,N_12193,N_12133);
nand U13377 (N_13377,N_12083,N_12819);
nand U13378 (N_13378,N_12984,N_12904);
or U13379 (N_13379,N_12485,N_12016);
nor U13380 (N_13380,N_12923,N_12471);
nand U13381 (N_13381,N_12012,N_12895);
xor U13382 (N_13382,N_12865,N_12686);
nor U13383 (N_13383,N_12892,N_12554);
nand U13384 (N_13384,N_12944,N_12341);
nand U13385 (N_13385,N_12650,N_12935);
nand U13386 (N_13386,N_12190,N_12573);
and U13387 (N_13387,N_12394,N_12583);
and U13388 (N_13388,N_12472,N_12673);
nand U13389 (N_13389,N_12797,N_12985);
and U13390 (N_13390,N_12766,N_12721);
and U13391 (N_13391,N_12961,N_12788);
nand U13392 (N_13392,N_12918,N_12078);
nor U13393 (N_13393,N_12814,N_12194);
and U13394 (N_13394,N_12416,N_12365);
or U13395 (N_13395,N_12743,N_12712);
nor U13396 (N_13396,N_12393,N_12751);
or U13397 (N_13397,N_12976,N_12633);
and U13398 (N_13398,N_12645,N_12809);
or U13399 (N_13399,N_12476,N_12072);
and U13400 (N_13400,N_12147,N_12021);
or U13401 (N_13401,N_12090,N_12642);
nor U13402 (N_13402,N_12104,N_12771);
or U13403 (N_13403,N_12786,N_12298);
and U13404 (N_13404,N_12949,N_12971);
and U13405 (N_13405,N_12170,N_12077);
nor U13406 (N_13406,N_12067,N_12052);
and U13407 (N_13407,N_12793,N_12317);
and U13408 (N_13408,N_12603,N_12405);
nand U13409 (N_13409,N_12326,N_12060);
nand U13410 (N_13410,N_12947,N_12649);
nor U13411 (N_13411,N_12528,N_12733);
and U13412 (N_13412,N_12523,N_12833);
nor U13413 (N_13413,N_12198,N_12929);
and U13414 (N_13414,N_12237,N_12434);
nand U13415 (N_13415,N_12678,N_12138);
or U13416 (N_13416,N_12481,N_12466);
nand U13417 (N_13417,N_12989,N_12577);
or U13418 (N_13418,N_12720,N_12108);
nand U13419 (N_13419,N_12032,N_12713);
or U13420 (N_13420,N_12992,N_12744);
and U13421 (N_13421,N_12141,N_12207);
nor U13422 (N_13422,N_12896,N_12665);
and U13423 (N_13423,N_12545,N_12105);
nor U13424 (N_13424,N_12707,N_12236);
nand U13425 (N_13425,N_12591,N_12565);
and U13426 (N_13426,N_12905,N_12184);
or U13427 (N_13427,N_12030,N_12484);
and U13428 (N_13428,N_12468,N_12589);
and U13429 (N_13429,N_12452,N_12031);
nor U13430 (N_13430,N_12130,N_12943);
nor U13431 (N_13431,N_12818,N_12360);
nor U13432 (N_13432,N_12152,N_12411);
and U13433 (N_13433,N_12218,N_12151);
or U13434 (N_13434,N_12517,N_12086);
or U13435 (N_13435,N_12044,N_12160);
and U13436 (N_13436,N_12055,N_12164);
and U13437 (N_13437,N_12827,N_12414);
and U13438 (N_13438,N_12859,N_12708);
nand U13439 (N_13439,N_12037,N_12975);
nor U13440 (N_13440,N_12717,N_12221);
nor U13441 (N_13441,N_12541,N_12028);
nor U13442 (N_13442,N_12344,N_12399);
and U13443 (N_13443,N_12902,N_12886);
or U13444 (N_13444,N_12352,N_12001);
or U13445 (N_13445,N_12262,N_12852);
or U13446 (N_13446,N_12578,N_12962);
nor U13447 (N_13447,N_12129,N_12449);
nor U13448 (N_13448,N_12952,N_12045);
or U13449 (N_13449,N_12900,N_12981);
and U13450 (N_13450,N_12729,N_12622);
nor U13451 (N_13451,N_12235,N_12679);
nor U13452 (N_13452,N_12099,N_12114);
nor U13453 (N_13453,N_12354,N_12759);
nor U13454 (N_13454,N_12146,N_12311);
and U13455 (N_13455,N_12208,N_12580);
nor U13456 (N_13456,N_12688,N_12928);
nand U13457 (N_13457,N_12042,N_12258);
nand U13458 (N_13458,N_12575,N_12335);
or U13459 (N_13459,N_12358,N_12994);
nor U13460 (N_13460,N_12919,N_12662);
and U13461 (N_13461,N_12763,N_12132);
and U13462 (N_13462,N_12314,N_12261);
and U13463 (N_13463,N_12113,N_12641);
and U13464 (N_13464,N_12059,N_12437);
or U13465 (N_13465,N_12249,N_12931);
or U13466 (N_13466,N_12348,N_12887);
or U13467 (N_13467,N_12936,N_12585);
and U13468 (N_13468,N_12263,N_12191);
nor U13469 (N_13469,N_12945,N_12280);
nand U13470 (N_13470,N_12015,N_12361);
nand U13471 (N_13471,N_12812,N_12431);
and U13472 (N_13472,N_12082,N_12655);
or U13473 (N_13473,N_12419,N_12616);
nor U13474 (N_13474,N_12694,N_12279);
nand U13475 (N_13475,N_12780,N_12118);
nand U13476 (N_13476,N_12516,N_12934);
nand U13477 (N_13477,N_12664,N_12548);
and U13478 (N_13478,N_12303,N_12571);
nand U13479 (N_13479,N_12256,N_12966);
nor U13480 (N_13480,N_12290,N_12370);
nand U13481 (N_13481,N_12284,N_12489);
nor U13482 (N_13482,N_12525,N_12333);
nor U13483 (N_13483,N_12884,N_12479);
nand U13484 (N_13484,N_12948,N_12963);
and U13485 (N_13485,N_12488,N_12174);
nand U13486 (N_13486,N_12423,N_12821);
and U13487 (N_13487,N_12858,N_12598);
nor U13488 (N_13488,N_12741,N_12787);
or U13489 (N_13489,N_12866,N_12562);
and U13490 (N_13490,N_12043,N_12183);
nor U13491 (N_13491,N_12901,N_12632);
and U13492 (N_13492,N_12396,N_12495);
nor U13493 (N_13493,N_12762,N_12663);
nand U13494 (N_13494,N_12176,N_12322);
and U13495 (N_13495,N_12569,N_12828);
nand U13496 (N_13496,N_12014,N_12547);
or U13497 (N_13497,N_12898,N_12486);
nand U13498 (N_13498,N_12294,N_12579);
xnor U13499 (N_13499,N_12535,N_12490);
and U13500 (N_13500,N_12228,N_12989);
or U13501 (N_13501,N_12653,N_12285);
nor U13502 (N_13502,N_12514,N_12932);
or U13503 (N_13503,N_12232,N_12130);
or U13504 (N_13504,N_12448,N_12278);
or U13505 (N_13505,N_12390,N_12680);
nand U13506 (N_13506,N_12483,N_12160);
or U13507 (N_13507,N_12132,N_12072);
or U13508 (N_13508,N_12659,N_12679);
nor U13509 (N_13509,N_12467,N_12536);
and U13510 (N_13510,N_12934,N_12023);
or U13511 (N_13511,N_12410,N_12768);
nand U13512 (N_13512,N_12174,N_12060);
and U13513 (N_13513,N_12150,N_12348);
or U13514 (N_13514,N_12737,N_12561);
nand U13515 (N_13515,N_12929,N_12178);
nor U13516 (N_13516,N_12844,N_12215);
and U13517 (N_13517,N_12955,N_12841);
nand U13518 (N_13518,N_12106,N_12730);
or U13519 (N_13519,N_12439,N_12187);
or U13520 (N_13520,N_12023,N_12646);
nand U13521 (N_13521,N_12800,N_12481);
nand U13522 (N_13522,N_12183,N_12108);
and U13523 (N_13523,N_12623,N_12275);
and U13524 (N_13524,N_12026,N_12959);
nand U13525 (N_13525,N_12700,N_12926);
nor U13526 (N_13526,N_12449,N_12925);
and U13527 (N_13527,N_12287,N_12445);
nand U13528 (N_13528,N_12386,N_12148);
or U13529 (N_13529,N_12467,N_12406);
or U13530 (N_13530,N_12412,N_12865);
nor U13531 (N_13531,N_12506,N_12015);
nor U13532 (N_13532,N_12570,N_12239);
nor U13533 (N_13533,N_12937,N_12390);
nor U13534 (N_13534,N_12753,N_12000);
nand U13535 (N_13535,N_12593,N_12530);
nor U13536 (N_13536,N_12252,N_12518);
and U13537 (N_13537,N_12413,N_12372);
and U13538 (N_13538,N_12482,N_12777);
nor U13539 (N_13539,N_12016,N_12767);
or U13540 (N_13540,N_12129,N_12057);
and U13541 (N_13541,N_12200,N_12191);
and U13542 (N_13542,N_12172,N_12115);
and U13543 (N_13543,N_12209,N_12411);
or U13544 (N_13544,N_12352,N_12859);
nand U13545 (N_13545,N_12937,N_12452);
nor U13546 (N_13546,N_12995,N_12004);
and U13547 (N_13547,N_12942,N_12036);
nand U13548 (N_13548,N_12445,N_12085);
nand U13549 (N_13549,N_12440,N_12906);
nor U13550 (N_13550,N_12306,N_12008);
nor U13551 (N_13551,N_12793,N_12735);
and U13552 (N_13552,N_12750,N_12094);
and U13553 (N_13553,N_12671,N_12247);
xnor U13554 (N_13554,N_12230,N_12555);
nor U13555 (N_13555,N_12198,N_12833);
nand U13556 (N_13556,N_12653,N_12051);
nor U13557 (N_13557,N_12830,N_12879);
nor U13558 (N_13558,N_12070,N_12668);
nor U13559 (N_13559,N_12394,N_12096);
nor U13560 (N_13560,N_12548,N_12400);
and U13561 (N_13561,N_12207,N_12194);
xor U13562 (N_13562,N_12374,N_12066);
nand U13563 (N_13563,N_12376,N_12530);
or U13564 (N_13564,N_12358,N_12398);
or U13565 (N_13565,N_12032,N_12404);
nand U13566 (N_13566,N_12512,N_12457);
nor U13567 (N_13567,N_12995,N_12134);
nand U13568 (N_13568,N_12320,N_12782);
or U13569 (N_13569,N_12294,N_12553);
nand U13570 (N_13570,N_12177,N_12544);
or U13571 (N_13571,N_12031,N_12592);
nor U13572 (N_13572,N_12152,N_12498);
nor U13573 (N_13573,N_12731,N_12722);
nand U13574 (N_13574,N_12849,N_12481);
and U13575 (N_13575,N_12945,N_12666);
or U13576 (N_13576,N_12455,N_12008);
and U13577 (N_13577,N_12478,N_12200);
or U13578 (N_13578,N_12347,N_12697);
nor U13579 (N_13579,N_12796,N_12506);
xnor U13580 (N_13580,N_12954,N_12247);
and U13581 (N_13581,N_12134,N_12217);
or U13582 (N_13582,N_12471,N_12010);
and U13583 (N_13583,N_12274,N_12854);
or U13584 (N_13584,N_12216,N_12193);
and U13585 (N_13585,N_12090,N_12383);
nand U13586 (N_13586,N_12360,N_12285);
and U13587 (N_13587,N_12580,N_12789);
or U13588 (N_13588,N_12176,N_12787);
nor U13589 (N_13589,N_12816,N_12656);
nor U13590 (N_13590,N_12267,N_12149);
or U13591 (N_13591,N_12213,N_12841);
nor U13592 (N_13592,N_12413,N_12831);
nand U13593 (N_13593,N_12953,N_12196);
nand U13594 (N_13594,N_12642,N_12029);
or U13595 (N_13595,N_12266,N_12858);
nand U13596 (N_13596,N_12494,N_12378);
or U13597 (N_13597,N_12793,N_12491);
or U13598 (N_13598,N_12296,N_12528);
nor U13599 (N_13599,N_12626,N_12658);
and U13600 (N_13600,N_12228,N_12007);
and U13601 (N_13601,N_12369,N_12287);
nand U13602 (N_13602,N_12164,N_12898);
nand U13603 (N_13603,N_12781,N_12322);
nor U13604 (N_13604,N_12645,N_12872);
nand U13605 (N_13605,N_12004,N_12771);
nand U13606 (N_13606,N_12273,N_12113);
nand U13607 (N_13607,N_12499,N_12247);
nor U13608 (N_13608,N_12761,N_12876);
nor U13609 (N_13609,N_12585,N_12974);
nor U13610 (N_13610,N_12344,N_12217);
or U13611 (N_13611,N_12413,N_12481);
and U13612 (N_13612,N_12863,N_12435);
and U13613 (N_13613,N_12120,N_12299);
or U13614 (N_13614,N_12046,N_12159);
and U13615 (N_13615,N_12717,N_12774);
and U13616 (N_13616,N_12503,N_12162);
and U13617 (N_13617,N_12186,N_12032);
and U13618 (N_13618,N_12226,N_12953);
or U13619 (N_13619,N_12579,N_12973);
or U13620 (N_13620,N_12553,N_12693);
and U13621 (N_13621,N_12954,N_12759);
and U13622 (N_13622,N_12360,N_12200);
nand U13623 (N_13623,N_12773,N_12089);
and U13624 (N_13624,N_12373,N_12981);
and U13625 (N_13625,N_12347,N_12618);
or U13626 (N_13626,N_12430,N_12979);
or U13627 (N_13627,N_12743,N_12117);
or U13628 (N_13628,N_12959,N_12491);
and U13629 (N_13629,N_12326,N_12864);
or U13630 (N_13630,N_12548,N_12298);
or U13631 (N_13631,N_12500,N_12267);
and U13632 (N_13632,N_12161,N_12504);
or U13633 (N_13633,N_12212,N_12667);
nor U13634 (N_13634,N_12211,N_12047);
and U13635 (N_13635,N_12419,N_12514);
nand U13636 (N_13636,N_12448,N_12901);
nand U13637 (N_13637,N_12531,N_12940);
nor U13638 (N_13638,N_12292,N_12528);
or U13639 (N_13639,N_12406,N_12558);
nor U13640 (N_13640,N_12572,N_12850);
nor U13641 (N_13641,N_12725,N_12024);
nand U13642 (N_13642,N_12386,N_12762);
and U13643 (N_13643,N_12220,N_12164);
or U13644 (N_13644,N_12524,N_12788);
xnor U13645 (N_13645,N_12182,N_12600);
or U13646 (N_13646,N_12834,N_12665);
or U13647 (N_13647,N_12055,N_12075);
or U13648 (N_13648,N_12596,N_12767);
nand U13649 (N_13649,N_12307,N_12031);
or U13650 (N_13650,N_12478,N_12182);
and U13651 (N_13651,N_12542,N_12241);
or U13652 (N_13652,N_12957,N_12938);
nor U13653 (N_13653,N_12513,N_12088);
nand U13654 (N_13654,N_12429,N_12832);
and U13655 (N_13655,N_12587,N_12734);
nand U13656 (N_13656,N_12309,N_12379);
or U13657 (N_13657,N_12451,N_12414);
or U13658 (N_13658,N_12921,N_12957);
nor U13659 (N_13659,N_12766,N_12565);
or U13660 (N_13660,N_12406,N_12806);
and U13661 (N_13661,N_12098,N_12930);
xnor U13662 (N_13662,N_12418,N_12841);
and U13663 (N_13663,N_12040,N_12831);
or U13664 (N_13664,N_12957,N_12175);
or U13665 (N_13665,N_12980,N_12994);
or U13666 (N_13666,N_12410,N_12950);
nand U13667 (N_13667,N_12445,N_12159);
nor U13668 (N_13668,N_12794,N_12198);
and U13669 (N_13669,N_12427,N_12572);
and U13670 (N_13670,N_12841,N_12840);
nor U13671 (N_13671,N_12052,N_12723);
nand U13672 (N_13672,N_12292,N_12818);
nand U13673 (N_13673,N_12809,N_12588);
or U13674 (N_13674,N_12605,N_12191);
nor U13675 (N_13675,N_12695,N_12795);
nand U13676 (N_13676,N_12962,N_12442);
and U13677 (N_13677,N_12604,N_12688);
nor U13678 (N_13678,N_12597,N_12295);
nand U13679 (N_13679,N_12113,N_12404);
nand U13680 (N_13680,N_12985,N_12480);
or U13681 (N_13681,N_12331,N_12552);
nor U13682 (N_13682,N_12201,N_12345);
nand U13683 (N_13683,N_12404,N_12309);
and U13684 (N_13684,N_12747,N_12712);
nand U13685 (N_13685,N_12239,N_12674);
nor U13686 (N_13686,N_12568,N_12521);
or U13687 (N_13687,N_12417,N_12776);
nand U13688 (N_13688,N_12569,N_12882);
and U13689 (N_13689,N_12727,N_12196);
and U13690 (N_13690,N_12042,N_12950);
nor U13691 (N_13691,N_12367,N_12195);
xor U13692 (N_13692,N_12625,N_12378);
and U13693 (N_13693,N_12313,N_12626);
nand U13694 (N_13694,N_12329,N_12757);
nand U13695 (N_13695,N_12355,N_12859);
and U13696 (N_13696,N_12883,N_12454);
and U13697 (N_13697,N_12764,N_12306);
or U13698 (N_13698,N_12440,N_12320);
nor U13699 (N_13699,N_12042,N_12304);
and U13700 (N_13700,N_12593,N_12472);
and U13701 (N_13701,N_12351,N_12364);
and U13702 (N_13702,N_12898,N_12831);
or U13703 (N_13703,N_12090,N_12235);
nor U13704 (N_13704,N_12372,N_12864);
nor U13705 (N_13705,N_12046,N_12014);
nand U13706 (N_13706,N_12633,N_12900);
or U13707 (N_13707,N_12779,N_12629);
nor U13708 (N_13708,N_12306,N_12507);
nand U13709 (N_13709,N_12704,N_12462);
and U13710 (N_13710,N_12894,N_12131);
nand U13711 (N_13711,N_12326,N_12139);
or U13712 (N_13712,N_12014,N_12302);
and U13713 (N_13713,N_12134,N_12486);
or U13714 (N_13714,N_12527,N_12795);
nor U13715 (N_13715,N_12204,N_12087);
or U13716 (N_13716,N_12000,N_12523);
or U13717 (N_13717,N_12217,N_12337);
and U13718 (N_13718,N_12580,N_12569);
and U13719 (N_13719,N_12610,N_12251);
and U13720 (N_13720,N_12010,N_12484);
nor U13721 (N_13721,N_12457,N_12190);
or U13722 (N_13722,N_12148,N_12701);
nand U13723 (N_13723,N_12284,N_12652);
or U13724 (N_13724,N_12538,N_12467);
nor U13725 (N_13725,N_12487,N_12275);
nor U13726 (N_13726,N_12863,N_12245);
nor U13727 (N_13727,N_12750,N_12108);
and U13728 (N_13728,N_12555,N_12806);
and U13729 (N_13729,N_12382,N_12395);
and U13730 (N_13730,N_12849,N_12522);
nor U13731 (N_13731,N_12608,N_12804);
and U13732 (N_13732,N_12765,N_12101);
and U13733 (N_13733,N_12493,N_12639);
and U13734 (N_13734,N_12418,N_12347);
or U13735 (N_13735,N_12905,N_12172);
nor U13736 (N_13736,N_12728,N_12188);
nand U13737 (N_13737,N_12288,N_12952);
and U13738 (N_13738,N_12032,N_12026);
nor U13739 (N_13739,N_12352,N_12753);
nand U13740 (N_13740,N_12780,N_12172);
and U13741 (N_13741,N_12458,N_12444);
nor U13742 (N_13742,N_12769,N_12954);
or U13743 (N_13743,N_12674,N_12535);
nand U13744 (N_13744,N_12868,N_12377);
nand U13745 (N_13745,N_12057,N_12863);
nand U13746 (N_13746,N_12892,N_12760);
nand U13747 (N_13747,N_12617,N_12252);
nand U13748 (N_13748,N_12288,N_12979);
and U13749 (N_13749,N_12794,N_12642);
nor U13750 (N_13750,N_12821,N_12803);
or U13751 (N_13751,N_12873,N_12131);
nand U13752 (N_13752,N_12219,N_12949);
nand U13753 (N_13753,N_12131,N_12693);
and U13754 (N_13754,N_12886,N_12556);
nor U13755 (N_13755,N_12500,N_12437);
or U13756 (N_13756,N_12321,N_12257);
and U13757 (N_13757,N_12546,N_12857);
or U13758 (N_13758,N_12401,N_12890);
and U13759 (N_13759,N_12622,N_12547);
or U13760 (N_13760,N_12367,N_12681);
or U13761 (N_13761,N_12747,N_12390);
nand U13762 (N_13762,N_12944,N_12882);
nand U13763 (N_13763,N_12412,N_12058);
or U13764 (N_13764,N_12307,N_12733);
nand U13765 (N_13765,N_12441,N_12281);
or U13766 (N_13766,N_12648,N_12857);
or U13767 (N_13767,N_12979,N_12302);
nand U13768 (N_13768,N_12239,N_12100);
and U13769 (N_13769,N_12863,N_12089);
or U13770 (N_13770,N_12747,N_12900);
xor U13771 (N_13771,N_12478,N_12636);
and U13772 (N_13772,N_12325,N_12218);
and U13773 (N_13773,N_12692,N_12986);
xor U13774 (N_13774,N_12405,N_12508);
nor U13775 (N_13775,N_12827,N_12233);
xnor U13776 (N_13776,N_12754,N_12984);
nand U13777 (N_13777,N_12174,N_12796);
nand U13778 (N_13778,N_12683,N_12392);
and U13779 (N_13779,N_12678,N_12050);
or U13780 (N_13780,N_12735,N_12982);
and U13781 (N_13781,N_12296,N_12988);
nor U13782 (N_13782,N_12077,N_12683);
and U13783 (N_13783,N_12260,N_12283);
and U13784 (N_13784,N_12301,N_12926);
or U13785 (N_13785,N_12566,N_12144);
nand U13786 (N_13786,N_12387,N_12721);
or U13787 (N_13787,N_12970,N_12526);
and U13788 (N_13788,N_12886,N_12266);
or U13789 (N_13789,N_12049,N_12947);
nand U13790 (N_13790,N_12076,N_12243);
nand U13791 (N_13791,N_12804,N_12696);
or U13792 (N_13792,N_12593,N_12417);
nand U13793 (N_13793,N_12056,N_12971);
and U13794 (N_13794,N_12100,N_12221);
and U13795 (N_13795,N_12636,N_12298);
nor U13796 (N_13796,N_12957,N_12168);
nor U13797 (N_13797,N_12218,N_12682);
or U13798 (N_13798,N_12537,N_12045);
and U13799 (N_13799,N_12018,N_12908);
nor U13800 (N_13800,N_12311,N_12304);
or U13801 (N_13801,N_12115,N_12835);
xor U13802 (N_13802,N_12197,N_12248);
nor U13803 (N_13803,N_12546,N_12868);
nand U13804 (N_13804,N_12323,N_12661);
nor U13805 (N_13805,N_12874,N_12628);
and U13806 (N_13806,N_12611,N_12873);
nor U13807 (N_13807,N_12372,N_12584);
and U13808 (N_13808,N_12316,N_12135);
nand U13809 (N_13809,N_12580,N_12081);
nor U13810 (N_13810,N_12021,N_12467);
or U13811 (N_13811,N_12681,N_12191);
nor U13812 (N_13812,N_12526,N_12506);
nand U13813 (N_13813,N_12479,N_12271);
or U13814 (N_13814,N_12314,N_12343);
or U13815 (N_13815,N_12638,N_12959);
nor U13816 (N_13816,N_12596,N_12873);
nand U13817 (N_13817,N_12341,N_12640);
or U13818 (N_13818,N_12072,N_12442);
or U13819 (N_13819,N_12124,N_12392);
nand U13820 (N_13820,N_12968,N_12422);
and U13821 (N_13821,N_12904,N_12742);
and U13822 (N_13822,N_12320,N_12218);
nand U13823 (N_13823,N_12029,N_12797);
nor U13824 (N_13824,N_12739,N_12206);
nor U13825 (N_13825,N_12081,N_12356);
nand U13826 (N_13826,N_12271,N_12074);
or U13827 (N_13827,N_12361,N_12236);
or U13828 (N_13828,N_12430,N_12770);
nand U13829 (N_13829,N_12012,N_12958);
and U13830 (N_13830,N_12326,N_12818);
or U13831 (N_13831,N_12322,N_12777);
nor U13832 (N_13832,N_12111,N_12344);
nand U13833 (N_13833,N_12133,N_12610);
nor U13834 (N_13834,N_12353,N_12580);
or U13835 (N_13835,N_12132,N_12022);
or U13836 (N_13836,N_12871,N_12249);
and U13837 (N_13837,N_12035,N_12898);
nand U13838 (N_13838,N_12377,N_12468);
nand U13839 (N_13839,N_12054,N_12568);
nand U13840 (N_13840,N_12701,N_12095);
nand U13841 (N_13841,N_12655,N_12026);
nor U13842 (N_13842,N_12645,N_12185);
and U13843 (N_13843,N_12221,N_12391);
xnor U13844 (N_13844,N_12562,N_12365);
nand U13845 (N_13845,N_12940,N_12116);
and U13846 (N_13846,N_12224,N_12679);
nand U13847 (N_13847,N_12419,N_12255);
or U13848 (N_13848,N_12542,N_12420);
or U13849 (N_13849,N_12376,N_12340);
nor U13850 (N_13850,N_12120,N_12256);
or U13851 (N_13851,N_12459,N_12486);
or U13852 (N_13852,N_12949,N_12580);
nor U13853 (N_13853,N_12193,N_12892);
nand U13854 (N_13854,N_12194,N_12313);
and U13855 (N_13855,N_12503,N_12513);
and U13856 (N_13856,N_12404,N_12354);
and U13857 (N_13857,N_12046,N_12760);
nor U13858 (N_13858,N_12649,N_12826);
and U13859 (N_13859,N_12975,N_12527);
and U13860 (N_13860,N_12888,N_12654);
nor U13861 (N_13861,N_12075,N_12006);
and U13862 (N_13862,N_12480,N_12612);
and U13863 (N_13863,N_12372,N_12570);
nor U13864 (N_13864,N_12137,N_12368);
or U13865 (N_13865,N_12252,N_12411);
or U13866 (N_13866,N_12449,N_12606);
nor U13867 (N_13867,N_12818,N_12507);
or U13868 (N_13868,N_12885,N_12624);
or U13869 (N_13869,N_12746,N_12952);
nand U13870 (N_13870,N_12395,N_12987);
nand U13871 (N_13871,N_12405,N_12263);
or U13872 (N_13872,N_12325,N_12045);
or U13873 (N_13873,N_12542,N_12884);
and U13874 (N_13874,N_12785,N_12651);
nand U13875 (N_13875,N_12599,N_12841);
or U13876 (N_13876,N_12908,N_12258);
nor U13877 (N_13877,N_12421,N_12159);
nand U13878 (N_13878,N_12547,N_12732);
nor U13879 (N_13879,N_12071,N_12414);
and U13880 (N_13880,N_12555,N_12929);
nor U13881 (N_13881,N_12155,N_12421);
nor U13882 (N_13882,N_12987,N_12761);
or U13883 (N_13883,N_12624,N_12275);
and U13884 (N_13884,N_12473,N_12102);
nand U13885 (N_13885,N_12276,N_12845);
nand U13886 (N_13886,N_12181,N_12069);
and U13887 (N_13887,N_12551,N_12222);
or U13888 (N_13888,N_12591,N_12011);
nand U13889 (N_13889,N_12838,N_12859);
or U13890 (N_13890,N_12192,N_12695);
and U13891 (N_13891,N_12143,N_12447);
and U13892 (N_13892,N_12348,N_12394);
and U13893 (N_13893,N_12032,N_12484);
and U13894 (N_13894,N_12440,N_12716);
or U13895 (N_13895,N_12093,N_12022);
nor U13896 (N_13896,N_12057,N_12398);
or U13897 (N_13897,N_12373,N_12744);
or U13898 (N_13898,N_12937,N_12441);
nand U13899 (N_13899,N_12759,N_12984);
and U13900 (N_13900,N_12078,N_12490);
nor U13901 (N_13901,N_12354,N_12313);
xnor U13902 (N_13902,N_12456,N_12086);
and U13903 (N_13903,N_12633,N_12815);
and U13904 (N_13904,N_12564,N_12531);
nor U13905 (N_13905,N_12282,N_12522);
or U13906 (N_13906,N_12920,N_12191);
and U13907 (N_13907,N_12655,N_12156);
and U13908 (N_13908,N_12056,N_12351);
and U13909 (N_13909,N_12885,N_12307);
nand U13910 (N_13910,N_12187,N_12928);
or U13911 (N_13911,N_12491,N_12281);
or U13912 (N_13912,N_12741,N_12192);
and U13913 (N_13913,N_12975,N_12033);
nor U13914 (N_13914,N_12300,N_12316);
and U13915 (N_13915,N_12347,N_12534);
and U13916 (N_13916,N_12293,N_12852);
and U13917 (N_13917,N_12175,N_12681);
and U13918 (N_13918,N_12810,N_12475);
nor U13919 (N_13919,N_12935,N_12786);
and U13920 (N_13920,N_12356,N_12550);
or U13921 (N_13921,N_12329,N_12713);
and U13922 (N_13922,N_12337,N_12184);
and U13923 (N_13923,N_12784,N_12032);
or U13924 (N_13924,N_12026,N_12304);
xor U13925 (N_13925,N_12645,N_12104);
nand U13926 (N_13926,N_12614,N_12074);
nand U13927 (N_13927,N_12860,N_12505);
and U13928 (N_13928,N_12065,N_12959);
nand U13929 (N_13929,N_12498,N_12075);
and U13930 (N_13930,N_12774,N_12323);
and U13931 (N_13931,N_12750,N_12038);
or U13932 (N_13932,N_12077,N_12749);
nor U13933 (N_13933,N_12591,N_12133);
nor U13934 (N_13934,N_12751,N_12273);
nand U13935 (N_13935,N_12583,N_12902);
or U13936 (N_13936,N_12089,N_12306);
nor U13937 (N_13937,N_12679,N_12371);
nand U13938 (N_13938,N_12352,N_12954);
nand U13939 (N_13939,N_12736,N_12491);
nor U13940 (N_13940,N_12068,N_12994);
nand U13941 (N_13941,N_12022,N_12554);
nor U13942 (N_13942,N_12850,N_12658);
and U13943 (N_13943,N_12440,N_12048);
nor U13944 (N_13944,N_12848,N_12342);
and U13945 (N_13945,N_12757,N_12853);
nor U13946 (N_13946,N_12030,N_12156);
nor U13947 (N_13947,N_12312,N_12536);
and U13948 (N_13948,N_12061,N_12863);
and U13949 (N_13949,N_12623,N_12052);
and U13950 (N_13950,N_12994,N_12867);
xor U13951 (N_13951,N_12350,N_12221);
or U13952 (N_13952,N_12628,N_12024);
xnor U13953 (N_13953,N_12378,N_12433);
nand U13954 (N_13954,N_12895,N_12210);
and U13955 (N_13955,N_12410,N_12592);
or U13956 (N_13956,N_12261,N_12681);
nor U13957 (N_13957,N_12781,N_12151);
nor U13958 (N_13958,N_12438,N_12039);
and U13959 (N_13959,N_12399,N_12676);
and U13960 (N_13960,N_12063,N_12165);
nor U13961 (N_13961,N_12819,N_12697);
nor U13962 (N_13962,N_12173,N_12953);
nor U13963 (N_13963,N_12662,N_12676);
nand U13964 (N_13964,N_12006,N_12109);
nor U13965 (N_13965,N_12390,N_12901);
nand U13966 (N_13966,N_12578,N_12544);
or U13967 (N_13967,N_12248,N_12511);
or U13968 (N_13968,N_12556,N_12665);
nand U13969 (N_13969,N_12092,N_12811);
and U13970 (N_13970,N_12623,N_12346);
or U13971 (N_13971,N_12893,N_12504);
or U13972 (N_13972,N_12637,N_12737);
nand U13973 (N_13973,N_12775,N_12623);
nand U13974 (N_13974,N_12560,N_12380);
or U13975 (N_13975,N_12650,N_12491);
or U13976 (N_13976,N_12395,N_12979);
and U13977 (N_13977,N_12893,N_12360);
and U13978 (N_13978,N_12554,N_12859);
nor U13979 (N_13979,N_12335,N_12923);
and U13980 (N_13980,N_12155,N_12937);
and U13981 (N_13981,N_12924,N_12774);
and U13982 (N_13982,N_12629,N_12690);
nor U13983 (N_13983,N_12092,N_12698);
nand U13984 (N_13984,N_12738,N_12850);
nand U13985 (N_13985,N_12815,N_12377);
and U13986 (N_13986,N_12620,N_12145);
or U13987 (N_13987,N_12137,N_12260);
nand U13988 (N_13988,N_12720,N_12128);
or U13989 (N_13989,N_12750,N_12355);
or U13990 (N_13990,N_12228,N_12276);
nor U13991 (N_13991,N_12857,N_12217);
or U13992 (N_13992,N_12966,N_12413);
or U13993 (N_13993,N_12778,N_12310);
or U13994 (N_13994,N_12307,N_12266);
or U13995 (N_13995,N_12667,N_12440);
nand U13996 (N_13996,N_12229,N_12155);
and U13997 (N_13997,N_12312,N_12573);
nor U13998 (N_13998,N_12299,N_12787);
nor U13999 (N_13999,N_12409,N_12478);
nor U14000 (N_14000,N_13716,N_13547);
nand U14001 (N_14001,N_13591,N_13804);
nand U14002 (N_14002,N_13352,N_13977);
nand U14003 (N_14003,N_13443,N_13135);
nand U14004 (N_14004,N_13745,N_13259);
nand U14005 (N_14005,N_13570,N_13142);
nand U14006 (N_14006,N_13153,N_13574);
nand U14007 (N_14007,N_13592,N_13768);
or U14008 (N_14008,N_13278,N_13100);
or U14009 (N_14009,N_13931,N_13654);
or U14010 (N_14010,N_13295,N_13034);
nand U14011 (N_14011,N_13561,N_13718);
and U14012 (N_14012,N_13885,N_13524);
and U14013 (N_14013,N_13713,N_13587);
xnor U14014 (N_14014,N_13971,N_13277);
and U14015 (N_14015,N_13364,N_13498);
or U14016 (N_14016,N_13317,N_13645);
and U14017 (N_14017,N_13377,N_13923);
nor U14018 (N_14018,N_13422,N_13282);
and U14019 (N_14019,N_13534,N_13469);
nand U14020 (N_14020,N_13919,N_13458);
and U14021 (N_14021,N_13476,N_13834);
nand U14022 (N_14022,N_13214,N_13554);
nor U14023 (N_14023,N_13859,N_13240);
nor U14024 (N_14024,N_13179,N_13589);
or U14025 (N_14025,N_13794,N_13399);
xor U14026 (N_14026,N_13462,N_13960);
or U14027 (N_14027,N_13744,N_13509);
nand U14028 (N_14028,N_13480,N_13292);
nor U14029 (N_14029,N_13691,N_13098);
and U14030 (N_14030,N_13661,N_13375);
or U14031 (N_14031,N_13588,N_13037);
and U14032 (N_14032,N_13769,N_13900);
and U14033 (N_14033,N_13218,N_13429);
nand U14034 (N_14034,N_13488,N_13912);
nor U14035 (N_14035,N_13829,N_13950);
and U14036 (N_14036,N_13348,N_13027);
nor U14037 (N_14037,N_13192,N_13263);
nor U14038 (N_14038,N_13898,N_13323);
or U14039 (N_14039,N_13515,N_13230);
nor U14040 (N_14040,N_13467,N_13793);
nor U14041 (N_14041,N_13092,N_13830);
nor U14042 (N_14042,N_13167,N_13594);
nor U14043 (N_14043,N_13123,N_13644);
nor U14044 (N_14044,N_13933,N_13294);
nand U14045 (N_14045,N_13531,N_13017);
nor U14046 (N_14046,N_13300,N_13396);
or U14047 (N_14047,N_13328,N_13679);
and U14048 (N_14048,N_13265,N_13506);
and U14049 (N_14049,N_13023,N_13190);
or U14050 (N_14050,N_13215,N_13684);
and U14051 (N_14051,N_13722,N_13310);
nor U14052 (N_14052,N_13938,N_13775);
nand U14053 (N_14053,N_13852,N_13143);
and U14054 (N_14054,N_13903,N_13372);
nor U14055 (N_14055,N_13992,N_13784);
nand U14056 (N_14056,N_13433,N_13827);
or U14057 (N_14057,N_13464,N_13741);
and U14058 (N_14058,N_13740,N_13557);
nor U14059 (N_14059,N_13417,N_13523);
or U14060 (N_14060,N_13477,N_13795);
or U14061 (N_14061,N_13596,N_13096);
nand U14062 (N_14062,N_13955,N_13978);
and U14063 (N_14063,N_13033,N_13216);
and U14064 (N_14064,N_13086,N_13544);
and U14065 (N_14065,N_13507,N_13370);
nand U14066 (N_14066,N_13389,N_13045);
and U14067 (N_14067,N_13354,N_13281);
nor U14068 (N_14068,N_13669,N_13917);
and U14069 (N_14069,N_13332,N_13351);
nand U14070 (N_14070,N_13670,N_13749);
nor U14071 (N_14071,N_13773,N_13910);
xor U14072 (N_14072,N_13441,N_13787);
nand U14073 (N_14073,N_13656,N_13851);
nand U14074 (N_14074,N_13382,N_13770);
or U14075 (N_14075,N_13831,N_13064);
nor U14076 (N_14076,N_13623,N_13242);
nor U14077 (N_14077,N_13176,N_13502);
xnor U14078 (N_14078,N_13707,N_13867);
nor U14079 (N_14079,N_13863,N_13003);
nor U14080 (N_14080,N_13089,N_13401);
nand U14081 (N_14081,N_13511,N_13520);
and U14082 (N_14082,N_13137,N_13388);
or U14083 (N_14083,N_13193,N_13754);
nand U14084 (N_14084,N_13271,N_13823);
nand U14085 (N_14085,N_13421,N_13896);
nor U14086 (N_14086,N_13457,N_13049);
and U14087 (N_14087,N_13172,N_13493);
and U14088 (N_14088,N_13132,N_13924);
or U14089 (N_14089,N_13657,N_13161);
nand U14090 (N_14090,N_13957,N_13880);
and U14091 (N_14091,N_13942,N_13133);
and U14092 (N_14092,N_13538,N_13334);
and U14093 (N_14093,N_13582,N_13432);
or U14094 (N_14094,N_13427,N_13188);
nor U14095 (N_14095,N_13403,N_13466);
nor U14096 (N_14096,N_13956,N_13168);
and U14097 (N_14097,N_13384,N_13024);
and U14098 (N_14098,N_13288,N_13239);
nand U14099 (N_14099,N_13410,N_13029);
nor U14100 (N_14100,N_13571,N_13129);
nor U14101 (N_14101,N_13616,N_13762);
nor U14102 (N_14102,N_13076,N_13871);
nor U14103 (N_14103,N_13101,N_13597);
or U14104 (N_14104,N_13361,N_13890);
nand U14105 (N_14105,N_13651,N_13455);
nor U14106 (N_14106,N_13012,N_13966);
nand U14107 (N_14107,N_13980,N_13201);
nor U14108 (N_14108,N_13122,N_13365);
nor U14109 (N_14109,N_13822,N_13875);
nor U14110 (N_14110,N_13873,N_13102);
or U14111 (N_14111,N_13811,N_13270);
or U14112 (N_14112,N_13800,N_13131);
nor U14113 (N_14113,N_13854,N_13212);
nor U14114 (N_14114,N_13341,N_13888);
nand U14115 (N_14115,N_13066,N_13330);
and U14116 (N_14116,N_13947,N_13932);
nor U14117 (N_14117,N_13202,N_13110);
and U14118 (N_14118,N_13849,N_13540);
or U14119 (N_14119,N_13513,N_13985);
nor U14120 (N_14120,N_13986,N_13009);
or U14121 (N_14121,N_13695,N_13302);
or U14122 (N_14122,N_13234,N_13580);
and U14123 (N_14123,N_13556,N_13714);
nand U14124 (N_14124,N_13084,N_13519);
or U14125 (N_14125,N_13073,N_13438);
nand U14126 (N_14126,N_13319,N_13094);
or U14127 (N_14127,N_13260,N_13892);
or U14128 (N_14128,N_13810,N_13198);
or U14129 (N_14129,N_13170,N_13573);
or U14130 (N_14130,N_13449,N_13727);
or U14131 (N_14131,N_13191,N_13836);
nand U14132 (N_14132,N_13865,N_13763);
nand U14133 (N_14133,N_13478,N_13991);
or U14134 (N_14134,N_13283,N_13456);
nand U14135 (N_14135,N_13327,N_13549);
or U14136 (N_14136,N_13777,N_13087);
or U14137 (N_14137,N_13247,N_13008);
and U14138 (N_14138,N_13647,N_13376);
nand U14139 (N_14139,N_13968,N_13155);
and U14140 (N_14140,N_13567,N_13864);
or U14141 (N_14141,N_13158,N_13813);
nand U14142 (N_14142,N_13545,N_13610);
nand U14143 (N_14143,N_13901,N_13210);
and U14144 (N_14144,N_13445,N_13759);
and U14145 (N_14145,N_13454,N_13043);
nand U14146 (N_14146,N_13386,N_13815);
and U14147 (N_14147,N_13553,N_13862);
nand U14148 (N_14148,N_13149,N_13847);
nor U14149 (N_14149,N_13621,N_13363);
nor U14150 (N_14150,N_13127,N_13649);
nor U14151 (N_14151,N_13802,N_13126);
or U14152 (N_14152,N_13378,N_13431);
and U14153 (N_14153,N_13374,N_13692);
nor U14154 (N_14154,N_13479,N_13877);
and U14155 (N_14155,N_13020,N_13748);
and U14156 (N_14156,N_13147,N_13079);
nand U14157 (N_14157,N_13371,N_13408);
and U14158 (N_14158,N_13551,N_13252);
nor U14159 (N_14159,N_13850,N_13710);
or U14160 (N_14160,N_13184,N_13514);
and U14161 (N_14161,N_13564,N_13781);
and U14162 (N_14162,N_13952,N_13324);
nor U14163 (N_14163,N_13735,N_13653);
and U14164 (N_14164,N_13720,N_13275);
nand U14165 (N_14165,N_13182,N_13979);
or U14166 (N_14166,N_13208,N_13491);
and U14167 (N_14167,N_13030,N_13090);
nand U14168 (N_14168,N_13696,N_13231);
and U14169 (N_14169,N_13878,N_13313);
or U14170 (N_14170,N_13638,N_13286);
nand U14171 (N_14171,N_13350,N_13533);
nor U14172 (N_14172,N_13088,N_13998);
or U14173 (N_14173,N_13618,N_13044);
and U14174 (N_14174,N_13136,N_13953);
or U14175 (N_14175,N_13093,N_13819);
and U14176 (N_14176,N_13293,N_13765);
and U14177 (N_14177,N_13052,N_13316);
nand U14178 (N_14178,N_13434,N_13289);
and U14179 (N_14179,N_13333,N_13711);
or U14180 (N_14180,N_13171,N_13972);
and U14181 (N_14181,N_13790,N_13887);
or U14182 (N_14182,N_13016,N_13818);
nor U14183 (N_14183,N_13083,N_13672);
nor U14184 (N_14184,N_13632,N_13995);
or U14185 (N_14185,N_13107,N_13255);
and U14186 (N_14186,N_13284,N_13500);
or U14187 (N_14187,N_13848,N_13642);
nor U14188 (N_14188,N_13032,N_13419);
and U14189 (N_14189,N_13204,N_13999);
nor U14190 (N_14190,N_13832,N_13267);
and U14191 (N_14191,N_13505,N_13314);
and U14192 (N_14192,N_13002,N_13673);
and U14193 (N_14193,N_13261,N_13072);
and U14194 (N_14194,N_13633,N_13959);
nor U14195 (N_14195,N_13719,N_13611);
or U14196 (N_14196,N_13468,N_13766);
nand U14197 (N_14197,N_13121,N_13742);
nor U14198 (N_14198,N_13881,N_13050);
nand U14199 (N_14199,N_13211,N_13721);
nand U14200 (N_14200,N_13060,N_13853);
nand U14201 (N_14201,N_13934,N_13413);
or U14202 (N_14202,N_13353,N_13470);
or U14203 (N_14203,N_13563,N_13990);
nor U14204 (N_14204,N_13501,N_13035);
and U14205 (N_14205,N_13307,N_13362);
nor U14206 (N_14206,N_13897,N_13418);
xnor U14207 (N_14207,N_13005,N_13059);
nand U14208 (N_14208,N_13726,N_13447);
and U14209 (N_14209,N_13337,N_13575);
nand U14210 (N_14210,N_13635,N_13648);
nor U14211 (N_14211,N_13228,N_13063);
nor U14212 (N_14212,N_13837,N_13806);
nor U14213 (N_14213,N_13583,N_13843);
nand U14214 (N_14214,N_13304,N_13146);
nor U14215 (N_14215,N_13883,N_13305);
nand U14216 (N_14216,N_13758,N_13785);
nor U14217 (N_14217,N_13015,N_13346);
or U14218 (N_14218,N_13541,N_13199);
nor U14219 (N_14219,N_13976,N_13322);
nand U14220 (N_14220,N_13660,N_13209);
nand U14221 (N_14221,N_13046,N_13522);
nor U14222 (N_14222,N_13537,N_13639);
nor U14223 (N_14223,N_13595,N_13308);
or U14224 (N_14224,N_13816,N_13014);
and U14225 (N_14225,N_13869,N_13593);
or U14226 (N_14226,N_13631,N_13948);
and U14227 (N_14227,N_13886,N_13598);
and U14228 (N_14228,N_13746,N_13951);
and U14229 (N_14229,N_13615,N_13124);
nand U14230 (N_14230,N_13974,N_13075);
nand U14231 (N_14231,N_13628,N_13266);
or U14232 (N_14232,N_13054,N_13680);
nor U14233 (N_14233,N_13803,N_13989);
nor U14234 (N_14234,N_13643,N_13729);
nand U14235 (N_14235,N_13671,N_13569);
or U14236 (N_14236,N_13922,N_13704);
nor U14237 (N_14237,N_13821,N_13926);
and U14238 (N_14238,N_13578,N_13860);
and U14239 (N_14239,N_13961,N_13344);
and U14240 (N_14240,N_13690,N_13516);
and U14241 (N_14241,N_13071,N_13439);
or U14242 (N_14242,N_13559,N_13543);
nand U14243 (N_14243,N_13928,N_13152);
or U14244 (N_14244,N_13258,N_13173);
nor U14245 (N_14245,N_13233,N_13734);
or U14246 (N_14246,N_13475,N_13398);
nand U14247 (N_14247,N_13820,N_13503);
nor U14248 (N_14248,N_13814,N_13700);
nand U14249 (N_14249,N_13941,N_13495);
and U14250 (N_14250,N_13437,N_13566);
or U14251 (N_14251,N_13057,N_13061);
nand U14252 (N_14252,N_13699,N_13982);
or U14253 (N_14253,N_13082,N_13780);
nand U14254 (N_14254,N_13665,N_13508);
nand U14255 (N_14255,N_13577,N_13664);
nand U14256 (N_14256,N_13637,N_13613);
nor U14257 (N_14257,N_13053,N_13915);
or U14258 (N_14258,N_13535,N_13004);
or U14259 (N_14259,N_13962,N_13303);
or U14260 (N_14260,N_13884,N_13459);
nor U14261 (N_14261,N_13117,N_13492);
nand U14262 (N_14262,N_13343,N_13113);
and U14263 (N_14263,N_13156,N_13237);
nand U14264 (N_14264,N_13602,N_13757);
or U14265 (N_14265,N_13141,N_13160);
nand U14266 (N_14266,N_13964,N_13868);
nand U14267 (N_14267,N_13808,N_13080);
and U14268 (N_14268,N_13969,N_13845);
or U14269 (N_14269,N_13169,N_13693);
nand U14270 (N_14270,N_13068,N_13095);
nor U14271 (N_14271,N_13297,N_13130);
nand U14272 (N_14272,N_13272,N_13451);
and U14273 (N_14273,N_13189,N_13743);
and U14274 (N_14274,N_13685,N_13911);
or U14275 (N_14275,N_13461,N_13497);
and U14276 (N_14276,N_13662,N_13311);
and U14277 (N_14277,N_13416,N_13298);
or U14278 (N_14278,N_13213,N_13006);
and U14279 (N_14279,N_13681,N_13021);
or U14280 (N_14280,N_13200,N_13166);
nand U14281 (N_14281,N_13423,N_13779);
nor U14282 (N_14282,N_13390,N_13357);
nor U14283 (N_14283,N_13668,N_13042);
nor U14284 (N_14284,N_13723,N_13750);
nor U14285 (N_14285,N_13655,N_13676);
nand U14286 (N_14286,N_13264,N_13162);
nor U14287 (N_14287,N_13689,N_13724);
nand U14288 (N_14288,N_13636,N_13366);
nand U14289 (N_14289,N_13125,N_13194);
nand U14290 (N_14290,N_13448,N_13791);
nor U14291 (N_14291,N_13512,N_13178);
or U14292 (N_14292,N_13894,N_13504);
and U14293 (N_14293,N_13165,N_13841);
and U14294 (N_14294,N_13530,N_13997);
nand U14295 (N_14295,N_13805,N_13708);
nand U14296 (N_14296,N_13174,N_13617);
and U14297 (N_14297,N_13929,N_13751);
or U14298 (N_14298,N_13356,N_13391);
or U14299 (N_14299,N_13013,N_13335);
or U14300 (N_14300,N_13144,N_13036);
or U14301 (N_14301,N_13097,N_13510);
nor U14302 (N_14302,N_13373,N_13148);
or U14303 (N_14303,N_13181,N_13186);
and U14304 (N_14304,N_13562,N_13930);
nand U14305 (N_14305,N_13529,N_13345);
and U14306 (N_14306,N_13380,N_13250);
nor U14307 (N_14307,N_13450,N_13446);
nand U14308 (N_14308,N_13776,N_13861);
and U14309 (N_14309,N_13331,N_13397);
or U14310 (N_14310,N_13369,N_13177);
nor U14311 (N_14311,N_13175,N_13039);
nand U14312 (N_14312,N_13904,N_13984);
nor U14313 (N_14313,N_13442,N_13667);
or U14314 (N_14314,N_13268,N_13355);
xor U14315 (N_14315,N_13675,N_13663);
and U14316 (N_14316,N_13646,N_13603);
nand U14317 (N_14317,N_13954,N_13725);
and U14318 (N_14318,N_13062,N_13788);
nand U14319 (N_14319,N_13614,N_13484);
and U14320 (N_14320,N_13634,N_13590);
and U14321 (N_14321,N_13460,N_13916);
nor U14322 (N_14322,N_13471,N_13796);
or U14323 (N_14323,N_13607,N_13728);
nand U14324 (N_14324,N_13222,N_13767);
nand U14325 (N_14325,N_13774,N_13279);
nand U14326 (N_14326,N_13440,N_13206);
and U14327 (N_14327,N_13091,N_13140);
nand U14328 (N_14328,N_13424,N_13678);
or U14329 (N_14329,N_13404,N_13855);
nand U14330 (N_14330,N_13605,N_13157);
nor U14331 (N_14331,N_13203,N_13183);
nand U14332 (N_14332,N_13983,N_13251);
nand U14333 (N_14333,N_13846,N_13812);
nand U14334 (N_14334,N_13698,N_13340);
or U14335 (N_14335,N_13921,N_13994);
nand U14336 (N_14336,N_13936,N_13550);
nand U14337 (N_14337,N_13128,N_13078);
or U14338 (N_14338,N_13320,N_13686);
and U14339 (N_14339,N_13817,N_13359);
and U14340 (N_14340,N_13001,N_13975);
nor U14341 (N_14341,N_13532,N_13151);
and U14342 (N_14342,N_13560,N_13889);
and U14343 (N_14343,N_13026,N_13835);
nor U14344 (N_14344,N_13238,N_13402);
nor U14345 (N_14345,N_13879,N_13118);
and U14346 (N_14346,N_13706,N_13326);
nor U14347 (N_14347,N_13565,N_13392);
xnor U14348 (N_14348,N_13712,N_13120);
nor U14349 (N_14349,N_13798,N_13572);
and U14350 (N_14350,N_13866,N_13435);
or U14351 (N_14351,N_13943,N_13274);
nor U14352 (N_14352,N_13601,N_13927);
or U14353 (N_14353,N_13395,N_13772);
or U14354 (N_14354,N_13895,N_13797);
or U14355 (N_14355,N_13620,N_13801);
nand U14356 (N_14356,N_13312,N_13963);
nand U14357 (N_14357,N_13526,N_13760);
or U14358 (N_14358,N_13858,N_13752);
nand U14359 (N_14359,N_13755,N_13058);
and U14360 (N_14360,N_13280,N_13612);
nor U14361 (N_14361,N_13627,N_13925);
nand U14362 (N_14362,N_13379,N_13558);
nor U14363 (N_14363,N_13739,N_13939);
or U14364 (N_14364,N_13619,N_13056);
nor U14365 (N_14365,N_13368,N_13038);
or U14366 (N_14366,N_13257,N_13993);
nor U14367 (N_14367,N_13856,N_13276);
nand U14368 (N_14368,N_13223,N_13109);
or U14369 (N_14369,N_13406,N_13048);
nand U14370 (N_14370,N_13040,N_13996);
or U14371 (N_14371,N_13299,N_13227);
or U14372 (N_14372,N_13273,N_13067);
and U14373 (N_14373,N_13677,N_13254);
and U14374 (N_14374,N_13249,N_13241);
nor U14375 (N_14375,N_13694,N_13367);
and U14376 (N_14376,N_13756,N_13065);
nand U14377 (N_14377,N_13473,N_13906);
nand U14378 (N_14378,N_13907,N_13783);
or U14379 (N_14379,N_13555,N_13463);
nor U14380 (N_14380,N_13290,N_13489);
or U14381 (N_14381,N_13285,N_13518);
nand U14382 (N_14382,N_13321,N_13909);
nor U14383 (N_14383,N_13414,N_13358);
and U14384 (N_14384,N_13217,N_13420);
nand U14385 (N_14385,N_13081,N_13196);
nand U14386 (N_14386,N_13824,N_13010);
and U14387 (N_14387,N_13949,N_13839);
nand U14388 (N_14388,N_13430,N_13246);
or U14389 (N_14389,N_13899,N_13018);
and U14390 (N_14390,N_13486,N_13622);
and U14391 (N_14391,N_13119,N_13426);
nand U14392 (N_14392,N_13652,N_13666);
nor U14393 (N_14393,N_13958,N_13902);
nor U14394 (N_14394,N_13394,N_13220);
nand U14395 (N_14395,N_13225,N_13838);
and U14396 (N_14396,N_13483,N_13347);
and U14397 (N_14397,N_13074,N_13474);
xnor U14398 (N_14398,N_13428,N_13600);
nor U14399 (N_14399,N_13874,N_13683);
nor U14400 (N_14400,N_13164,N_13650);
or U14401 (N_14401,N_13687,N_13070);
nand U14402 (N_14402,N_13625,N_13154);
nand U14403 (N_14403,N_13732,N_13360);
and U14404 (N_14404,N_13658,N_13764);
nor U14405 (N_14405,N_13499,N_13077);
nor U14406 (N_14406,N_13315,N_13920);
nand U14407 (N_14407,N_13047,N_13139);
or U14408 (N_14408,N_13221,N_13905);
nand U14409 (N_14409,N_13940,N_13945);
and U14410 (N_14410,N_13028,N_13778);
nand U14411 (N_14411,N_13262,N_13579);
or U14412 (N_14412,N_13329,N_13306);
and U14413 (N_14413,N_13608,N_13786);
or U14414 (N_14414,N_13581,N_13604);
and U14415 (N_14415,N_13296,N_13891);
and U14416 (N_14416,N_13106,N_13381);
nand U14417 (N_14417,N_13385,N_13715);
and U14418 (N_14418,N_13425,N_13630);
and U14419 (N_14419,N_13055,N_13232);
nand U14420 (N_14420,N_13465,N_13988);
or U14421 (N_14421,N_13548,N_13521);
nor U14422 (N_14422,N_13688,N_13235);
nand U14423 (N_14423,N_13197,N_13185);
or U14424 (N_14424,N_13114,N_13546);
nor U14425 (N_14425,N_13069,N_13496);
nor U14426 (N_14426,N_13000,N_13112);
and U14427 (N_14427,N_13145,N_13527);
or U14428 (N_14428,N_13789,N_13799);
or U14429 (N_14429,N_13609,N_13586);
nor U14430 (N_14430,N_13226,N_13236);
nor U14431 (N_14431,N_13253,N_13411);
nor U14432 (N_14432,N_13412,N_13336);
or U14433 (N_14433,N_13301,N_13937);
nor U14434 (N_14434,N_13485,N_13702);
nor U14435 (N_14435,N_13482,N_13552);
nand U14436 (N_14436,N_13525,N_13807);
nor U14437 (N_14437,N_13674,N_13697);
or U14438 (N_14438,N_13844,N_13967);
and U14439 (N_14439,N_13452,N_13517);
nor U14440 (N_14440,N_13244,N_13935);
nand U14441 (N_14441,N_13104,N_13914);
or U14442 (N_14442,N_13207,N_13453);
and U14443 (N_14443,N_13150,N_13606);
or U14444 (N_14444,N_13245,N_13444);
nor U14445 (N_14445,N_13318,N_13629);
nor U14446 (N_14446,N_13407,N_13753);
or U14447 (N_14447,N_13539,N_13342);
or U14448 (N_14448,N_13624,N_13041);
nand U14449 (N_14449,N_13737,N_13256);
and U14450 (N_14450,N_13876,N_13115);
nand U14451 (N_14451,N_13872,N_13747);
nor U14452 (N_14452,N_13826,N_13782);
and U14453 (N_14453,N_13913,N_13828);
nand U14454 (N_14454,N_13736,N_13882);
nor U14455 (N_14455,N_13659,N_13243);
nand U14456 (N_14456,N_13487,N_13269);
nand U14457 (N_14457,N_13965,N_13325);
and U14458 (N_14458,N_13472,N_13542);
and U14459 (N_14459,N_13857,N_13730);
or U14460 (N_14460,N_13011,N_13717);
nand U14461 (N_14461,N_13025,N_13031);
nand U14462 (N_14462,N_13705,N_13159);
or U14463 (N_14463,N_13981,N_13970);
nor U14464 (N_14464,N_13809,N_13738);
or U14465 (N_14465,N_13436,N_13568);
or U14466 (N_14466,N_13111,N_13022);
nor U14467 (N_14467,N_13219,N_13387);
or U14468 (N_14468,N_13528,N_13287);
nand U14469 (N_14469,N_13309,N_13116);
and U14470 (N_14470,N_13973,N_13833);
or U14471 (N_14471,N_13682,N_13761);
and U14472 (N_14472,N_13584,N_13007);
nor U14473 (N_14473,N_13481,N_13134);
nand U14474 (N_14474,N_13103,N_13893);
nor U14475 (N_14475,N_13944,N_13731);
or U14476 (N_14476,N_13641,N_13599);
and U14477 (N_14477,N_13051,N_13771);
or U14478 (N_14478,N_13908,N_13840);
and U14479 (N_14479,N_13163,N_13393);
or U14480 (N_14480,N_13085,N_13703);
and U14481 (N_14481,N_13405,N_13383);
and U14482 (N_14482,N_13180,N_13105);
or U14483 (N_14483,N_13400,N_13490);
or U14484 (N_14484,N_13195,N_13733);
xor U14485 (N_14485,N_13918,N_13792);
nand U14486 (N_14486,N_13701,N_13205);
or U14487 (N_14487,N_13248,N_13415);
nand U14488 (N_14488,N_13842,N_13494);
nand U14489 (N_14489,N_13576,N_13709);
and U14490 (N_14490,N_13825,N_13339);
or U14491 (N_14491,N_13640,N_13229);
nand U14492 (N_14492,N_13138,N_13987);
nand U14493 (N_14493,N_13291,N_13187);
nor U14494 (N_14494,N_13626,N_13409);
and U14495 (N_14495,N_13585,N_13108);
nor U14496 (N_14496,N_13224,N_13536);
nor U14497 (N_14497,N_13338,N_13019);
nand U14498 (N_14498,N_13099,N_13946);
nor U14499 (N_14499,N_13349,N_13870);
or U14500 (N_14500,N_13756,N_13798);
and U14501 (N_14501,N_13075,N_13693);
nand U14502 (N_14502,N_13814,N_13119);
and U14503 (N_14503,N_13131,N_13363);
and U14504 (N_14504,N_13639,N_13188);
or U14505 (N_14505,N_13783,N_13429);
and U14506 (N_14506,N_13082,N_13148);
nor U14507 (N_14507,N_13477,N_13242);
nand U14508 (N_14508,N_13142,N_13877);
nand U14509 (N_14509,N_13650,N_13054);
and U14510 (N_14510,N_13852,N_13447);
and U14511 (N_14511,N_13122,N_13790);
nand U14512 (N_14512,N_13586,N_13144);
or U14513 (N_14513,N_13341,N_13323);
nand U14514 (N_14514,N_13730,N_13931);
nand U14515 (N_14515,N_13609,N_13430);
nand U14516 (N_14516,N_13641,N_13232);
nand U14517 (N_14517,N_13954,N_13066);
or U14518 (N_14518,N_13629,N_13248);
and U14519 (N_14519,N_13886,N_13907);
nor U14520 (N_14520,N_13449,N_13878);
or U14521 (N_14521,N_13738,N_13737);
and U14522 (N_14522,N_13809,N_13086);
and U14523 (N_14523,N_13928,N_13763);
xnor U14524 (N_14524,N_13499,N_13248);
nor U14525 (N_14525,N_13718,N_13900);
xnor U14526 (N_14526,N_13170,N_13332);
nor U14527 (N_14527,N_13422,N_13667);
and U14528 (N_14528,N_13361,N_13383);
nand U14529 (N_14529,N_13511,N_13392);
nand U14530 (N_14530,N_13400,N_13717);
or U14531 (N_14531,N_13129,N_13646);
and U14532 (N_14532,N_13342,N_13041);
nor U14533 (N_14533,N_13188,N_13175);
nor U14534 (N_14534,N_13995,N_13214);
and U14535 (N_14535,N_13517,N_13658);
or U14536 (N_14536,N_13793,N_13329);
nor U14537 (N_14537,N_13860,N_13863);
nand U14538 (N_14538,N_13739,N_13509);
or U14539 (N_14539,N_13701,N_13790);
or U14540 (N_14540,N_13905,N_13763);
nor U14541 (N_14541,N_13579,N_13283);
nor U14542 (N_14542,N_13561,N_13377);
or U14543 (N_14543,N_13265,N_13485);
nor U14544 (N_14544,N_13702,N_13636);
and U14545 (N_14545,N_13401,N_13397);
nor U14546 (N_14546,N_13388,N_13677);
nor U14547 (N_14547,N_13308,N_13508);
xor U14548 (N_14548,N_13678,N_13146);
and U14549 (N_14549,N_13149,N_13327);
nand U14550 (N_14550,N_13968,N_13702);
and U14551 (N_14551,N_13866,N_13795);
nand U14552 (N_14552,N_13104,N_13892);
nor U14553 (N_14553,N_13307,N_13586);
or U14554 (N_14554,N_13668,N_13152);
nor U14555 (N_14555,N_13494,N_13098);
or U14556 (N_14556,N_13119,N_13661);
nor U14557 (N_14557,N_13823,N_13631);
and U14558 (N_14558,N_13865,N_13970);
nor U14559 (N_14559,N_13366,N_13468);
nor U14560 (N_14560,N_13276,N_13455);
or U14561 (N_14561,N_13540,N_13658);
nand U14562 (N_14562,N_13073,N_13749);
and U14563 (N_14563,N_13636,N_13611);
nand U14564 (N_14564,N_13628,N_13329);
or U14565 (N_14565,N_13014,N_13020);
and U14566 (N_14566,N_13774,N_13960);
nand U14567 (N_14567,N_13234,N_13496);
nor U14568 (N_14568,N_13806,N_13689);
and U14569 (N_14569,N_13294,N_13491);
and U14570 (N_14570,N_13594,N_13516);
nor U14571 (N_14571,N_13020,N_13428);
nand U14572 (N_14572,N_13594,N_13003);
or U14573 (N_14573,N_13492,N_13927);
or U14574 (N_14574,N_13360,N_13292);
or U14575 (N_14575,N_13750,N_13539);
nand U14576 (N_14576,N_13845,N_13832);
nor U14577 (N_14577,N_13519,N_13226);
nor U14578 (N_14578,N_13164,N_13727);
or U14579 (N_14579,N_13934,N_13167);
or U14580 (N_14580,N_13197,N_13632);
nor U14581 (N_14581,N_13177,N_13473);
or U14582 (N_14582,N_13643,N_13041);
nand U14583 (N_14583,N_13807,N_13945);
nor U14584 (N_14584,N_13581,N_13701);
nor U14585 (N_14585,N_13767,N_13980);
nand U14586 (N_14586,N_13094,N_13478);
nor U14587 (N_14587,N_13207,N_13990);
and U14588 (N_14588,N_13221,N_13572);
or U14589 (N_14589,N_13961,N_13628);
nand U14590 (N_14590,N_13162,N_13107);
or U14591 (N_14591,N_13859,N_13806);
or U14592 (N_14592,N_13549,N_13499);
nor U14593 (N_14593,N_13931,N_13268);
nand U14594 (N_14594,N_13776,N_13446);
nand U14595 (N_14595,N_13983,N_13138);
or U14596 (N_14596,N_13734,N_13451);
and U14597 (N_14597,N_13326,N_13989);
or U14598 (N_14598,N_13524,N_13977);
and U14599 (N_14599,N_13024,N_13202);
nor U14600 (N_14600,N_13674,N_13675);
nor U14601 (N_14601,N_13894,N_13213);
nor U14602 (N_14602,N_13236,N_13972);
or U14603 (N_14603,N_13625,N_13450);
nand U14604 (N_14604,N_13936,N_13317);
nor U14605 (N_14605,N_13291,N_13169);
or U14606 (N_14606,N_13332,N_13810);
and U14607 (N_14607,N_13486,N_13847);
or U14608 (N_14608,N_13173,N_13431);
xnor U14609 (N_14609,N_13035,N_13156);
nand U14610 (N_14610,N_13130,N_13634);
or U14611 (N_14611,N_13958,N_13195);
and U14612 (N_14612,N_13630,N_13387);
nand U14613 (N_14613,N_13816,N_13061);
or U14614 (N_14614,N_13388,N_13106);
nand U14615 (N_14615,N_13348,N_13736);
and U14616 (N_14616,N_13570,N_13695);
nor U14617 (N_14617,N_13475,N_13563);
and U14618 (N_14618,N_13916,N_13019);
nand U14619 (N_14619,N_13914,N_13776);
or U14620 (N_14620,N_13767,N_13012);
nor U14621 (N_14621,N_13763,N_13457);
nor U14622 (N_14622,N_13361,N_13844);
nand U14623 (N_14623,N_13233,N_13012);
nand U14624 (N_14624,N_13066,N_13248);
nor U14625 (N_14625,N_13333,N_13608);
and U14626 (N_14626,N_13980,N_13552);
nand U14627 (N_14627,N_13294,N_13719);
nand U14628 (N_14628,N_13991,N_13476);
or U14629 (N_14629,N_13067,N_13465);
nor U14630 (N_14630,N_13563,N_13085);
nor U14631 (N_14631,N_13528,N_13450);
and U14632 (N_14632,N_13157,N_13233);
nor U14633 (N_14633,N_13772,N_13833);
and U14634 (N_14634,N_13116,N_13707);
and U14635 (N_14635,N_13737,N_13357);
or U14636 (N_14636,N_13452,N_13016);
or U14637 (N_14637,N_13996,N_13127);
nand U14638 (N_14638,N_13996,N_13439);
and U14639 (N_14639,N_13461,N_13590);
nand U14640 (N_14640,N_13963,N_13685);
nand U14641 (N_14641,N_13235,N_13587);
and U14642 (N_14642,N_13596,N_13874);
and U14643 (N_14643,N_13862,N_13614);
nor U14644 (N_14644,N_13513,N_13810);
nand U14645 (N_14645,N_13283,N_13711);
nand U14646 (N_14646,N_13155,N_13131);
and U14647 (N_14647,N_13863,N_13637);
nor U14648 (N_14648,N_13234,N_13579);
nand U14649 (N_14649,N_13054,N_13844);
nor U14650 (N_14650,N_13374,N_13572);
nor U14651 (N_14651,N_13494,N_13156);
nor U14652 (N_14652,N_13841,N_13319);
nand U14653 (N_14653,N_13023,N_13288);
or U14654 (N_14654,N_13062,N_13707);
nand U14655 (N_14655,N_13530,N_13844);
nand U14656 (N_14656,N_13895,N_13256);
and U14657 (N_14657,N_13630,N_13756);
nand U14658 (N_14658,N_13029,N_13346);
or U14659 (N_14659,N_13026,N_13077);
or U14660 (N_14660,N_13131,N_13904);
nor U14661 (N_14661,N_13798,N_13668);
or U14662 (N_14662,N_13319,N_13069);
or U14663 (N_14663,N_13247,N_13433);
nor U14664 (N_14664,N_13220,N_13634);
and U14665 (N_14665,N_13577,N_13594);
nor U14666 (N_14666,N_13135,N_13165);
nand U14667 (N_14667,N_13312,N_13406);
nor U14668 (N_14668,N_13062,N_13517);
or U14669 (N_14669,N_13584,N_13392);
nor U14670 (N_14670,N_13965,N_13063);
nor U14671 (N_14671,N_13430,N_13783);
and U14672 (N_14672,N_13513,N_13704);
nor U14673 (N_14673,N_13192,N_13099);
or U14674 (N_14674,N_13020,N_13375);
nand U14675 (N_14675,N_13638,N_13540);
or U14676 (N_14676,N_13239,N_13025);
nor U14677 (N_14677,N_13293,N_13615);
or U14678 (N_14678,N_13252,N_13299);
nand U14679 (N_14679,N_13096,N_13007);
and U14680 (N_14680,N_13194,N_13422);
and U14681 (N_14681,N_13030,N_13457);
and U14682 (N_14682,N_13533,N_13872);
nand U14683 (N_14683,N_13258,N_13353);
nor U14684 (N_14684,N_13592,N_13289);
and U14685 (N_14685,N_13358,N_13319);
nand U14686 (N_14686,N_13499,N_13503);
nor U14687 (N_14687,N_13702,N_13294);
or U14688 (N_14688,N_13683,N_13873);
nor U14689 (N_14689,N_13065,N_13806);
nand U14690 (N_14690,N_13811,N_13347);
and U14691 (N_14691,N_13267,N_13086);
nand U14692 (N_14692,N_13398,N_13743);
and U14693 (N_14693,N_13614,N_13780);
and U14694 (N_14694,N_13026,N_13015);
and U14695 (N_14695,N_13167,N_13076);
nand U14696 (N_14696,N_13413,N_13861);
nand U14697 (N_14697,N_13513,N_13990);
or U14698 (N_14698,N_13698,N_13812);
and U14699 (N_14699,N_13433,N_13811);
or U14700 (N_14700,N_13611,N_13402);
nor U14701 (N_14701,N_13610,N_13970);
or U14702 (N_14702,N_13831,N_13707);
nor U14703 (N_14703,N_13077,N_13466);
or U14704 (N_14704,N_13510,N_13389);
and U14705 (N_14705,N_13193,N_13739);
xor U14706 (N_14706,N_13743,N_13673);
nand U14707 (N_14707,N_13916,N_13644);
nand U14708 (N_14708,N_13232,N_13212);
and U14709 (N_14709,N_13942,N_13691);
or U14710 (N_14710,N_13337,N_13535);
and U14711 (N_14711,N_13070,N_13293);
or U14712 (N_14712,N_13721,N_13899);
or U14713 (N_14713,N_13410,N_13677);
nor U14714 (N_14714,N_13366,N_13361);
and U14715 (N_14715,N_13700,N_13501);
nor U14716 (N_14716,N_13494,N_13663);
or U14717 (N_14717,N_13791,N_13924);
nand U14718 (N_14718,N_13909,N_13834);
or U14719 (N_14719,N_13181,N_13920);
nand U14720 (N_14720,N_13757,N_13241);
or U14721 (N_14721,N_13453,N_13812);
nor U14722 (N_14722,N_13582,N_13829);
and U14723 (N_14723,N_13787,N_13544);
nor U14724 (N_14724,N_13100,N_13317);
and U14725 (N_14725,N_13744,N_13395);
and U14726 (N_14726,N_13657,N_13230);
or U14727 (N_14727,N_13439,N_13010);
and U14728 (N_14728,N_13505,N_13805);
nand U14729 (N_14729,N_13352,N_13035);
nand U14730 (N_14730,N_13038,N_13904);
and U14731 (N_14731,N_13545,N_13052);
or U14732 (N_14732,N_13927,N_13946);
nor U14733 (N_14733,N_13990,N_13536);
nor U14734 (N_14734,N_13600,N_13910);
nor U14735 (N_14735,N_13210,N_13688);
nor U14736 (N_14736,N_13096,N_13960);
and U14737 (N_14737,N_13393,N_13870);
or U14738 (N_14738,N_13048,N_13136);
and U14739 (N_14739,N_13142,N_13579);
or U14740 (N_14740,N_13710,N_13451);
or U14741 (N_14741,N_13970,N_13779);
and U14742 (N_14742,N_13886,N_13983);
nor U14743 (N_14743,N_13973,N_13698);
nor U14744 (N_14744,N_13501,N_13951);
and U14745 (N_14745,N_13490,N_13399);
nor U14746 (N_14746,N_13352,N_13844);
or U14747 (N_14747,N_13884,N_13054);
nor U14748 (N_14748,N_13724,N_13680);
and U14749 (N_14749,N_13121,N_13399);
and U14750 (N_14750,N_13952,N_13969);
or U14751 (N_14751,N_13289,N_13810);
xnor U14752 (N_14752,N_13893,N_13889);
and U14753 (N_14753,N_13433,N_13462);
and U14754 (N_14754,N_13634,N_13062);
or U14755 (N_14755,N_13927,N_13607);
nand U14756 (N_14756,N_13907,N_13268);
nand U14757 (N_14757,N_13931,N_13915);
or U14758 (N_14758,N_13401,N_13568);
xnor U14759 (N_14759,N_13752,N_13012);
nor U14760 (N_14760,N_13396,N_13021);
nor U14761 (N_14761,N_13907,N_13455);
nand U14762 (N_14762,N_13057,N_13797);
and U14763 (N_14763,N_13629,N_13317);
or U14764 (N_14764,N_13062,N_13408);
nor U14765 (N_14765,N_13241,N_13362);
nor U14766 (N_14766,N_13702,N_13517);
or U14767 (N_14767,N_13797,N_13664);
and U14768 (N_14768,N_13506,N_13251);
nor U14769 (N_14769,N_13522,N_13981);
and U14770 (N_14770,N_13312,N_13685);
and U14771 (N_14771,N_13409,N_13466);
nor U14772 (N_14772,N_13307,N_13986);
or U14773 (N_14773,N_13123,N_13968);
nand U14774 (N_14774,N_13959,N_13983);
and U14775 (N_14775,N_13655,N_13420);
nor U14776 (N_14776,N_13762,N_13679);
and U14777 (N_14777,N_13920,N_13983);
and U14778 (N_14778,N_13866,N_13778);
or U14779 (N_14779,N_13200,N_13571);
or U14780 (N_14780,N_13099,N_13820);
xnor U14781 (N_14781,N_13725,N_13829);
and U14782 (N_14782,N_13922,N_13914);
nor U14783 (N_14783,N_13665,N_13175);
nor U14784 (N_14784,N_13598,N_13378);
or U14785 (N_14785,N_13839,N_13871);
and U14786 (N_14786,N_13410,N_13880);
nand U14787 (N_14787,N_13205,N_13707);
and U14788 (N_14788,N_13253,N_13551);
or U14789 (N_14789,N_13251,N_13242);
or U14790 (N_14790,N_13152,N_13415);
nor U14791 (N_14791,N_13532,N_13572);
and U14792 (N_14792,N_13207,N_13843);
nor U14793 (N_14793,N_13016,N_13588);
and U14794 (N_14794,N_13906,N_13739);
nand U14795 (N_14795,N_13583,N_13929);
nor U14796 (N_14796,N_13834,N_13778);
and U14797 (N_14797,N_13720,N_13788);
and U14798 (N_14798,N_13557,N_13633);
and U14799 (N_14799,N_13288,N_13637);
or U14800 (N_14800,N_13821,N_13158);
nor U14801 (N_14801,N_13052,N_13540);
or U14802 (N_14802,N_13777,N_13369);
or U14803 (N_14803,N_13763,N_13687);
nand U14804 (N_14804,N_13263,N_13486);
nand U14805 (N_14805,N_13262,N_13702);
nor U14806 (N_14806,N_13426,N_13091);
or U14807 (N_14807,N_13156,N_13048);
nor U14808 (N_14808,N_13802,N_13948);
and U14809 (N_14809,N_13938,N_13772);
nor U14810 (N_14810,N_13305,N_13836);
nor U14811 (N_14811,N_13626,N_13126);
nor U14812 (N_14812,N_13583,N_13622);
nor U14813 (N_14813,N_13560,N_13214);
and U14814 (N_14814,N_13677,N_13210);
or U14815 (N_14815,N_13017,N_13580);
nand U14816 (N_14816,N_13897,N_13112);
nand U14817 (N_14817,N_13482,N_13248);
or U14818 (N_14818,N_13093,N_13133);
nor U14819 (N_14819,N_13516,N_13193);
nand U14820 (N_14820,N_13033,N_13851);
or U14821 (N_14821,N_13592,N_13606);
nand U14822 (N_14822,N_13364,N_13149);
and U14823 (N_14823,N_13996,N_13133);
nor U14824 (N_14824,N_13242,N_13034);
nor U14825 (N_14825,N_13097,N_13167);
nor U14826 (N_14826,N_13502,N_13026);
nor U14827 (N_14827,N_13203,N_13479);
and U14828 (N_14828,N_13960,N_13011);
and U14829 (N_14829,N_13038,N_13537);
or U14830 (N_14830,N_13376,N_13467);
nor U14831 (N_14831,N_13010,N_13818);
nor U14832 (N_14832,N_13320,N_13109);
nand U14833 (N_14833,N_13699,N_13294);
and U14834 (N_14834,N_13499,N_13315);
and U14835 (N_14835,N_13383,N_13686);
nand U14836 (N_14836,N_13284,N_13384);
nand U14837 (N_14837,N_13952,N_13216);
and U14838 (N_14838,N_13844,N_13560);
nand U14839 (N_14839,N_13986,N_13947);
nor U14840 (N_14840,N_13289,N_13401);
or U14841 (N_14841,N_13956,N_13198);
and U14842 (N_14842,N_13566,N_13429);
nor U14843 (N_14843,N_13832,N_13279);
and U14844 (N_14844,N_13701,N_13244);
nand U14845 (N_14845,N_13745,N_13671);
and U14846 (N_14846,N_13865,N_13375);
and U14847 (N_14847,N_13521,N_13475);
nand U14848 (N_14848,N_13839,N_13533);
nor U14849 (N_14849,N_13190,N_13690);
xor U14850 (N_14850,N_13080,N_13707);
and U14851 (N_14851,N_13197,N_13943);
nor U14852 (N_14852,N_13888,N_13070);
nand U14853 (N_14853,N_13417,N_13839);
nand U14854 (N_14854,N_13912,N_13897);
or U14855 (N_14855,N_13528,N_13391);
nor U14856 (N_14856,N_13715,N_13814);
nand U14857 (N_14857,N_13205,N_13681);
and U14858 (N_14858,N_13672,N_13349);
nor U14859 (N_14859,N_13477,N_13232);
nand U14860 (N_14860,N_13437,N_13638);
nor U14861 (N_14861,N_13240,N_13083);
or U14862 (N_14862,N_13438,N_13970);
nand U14863 (N_14863,N_13865,N_13438);
and U14864 (N_14864,N_13256,N_13141);
nor U14865 (N_14865,N_13844,N_13672);
nor U14866 (N_14866,N_13873,N_13339);
or U14867 (N_14867,N_13228,N_13678);
and U14868 (N_14868,N_13482,N_13339);
and U14869 (N_14869,N_13157,N_13135);
or U14870 (N_14870,N_13262,N_13268);
nand U14871 (N_14871,N_13317,N_13112);
or U14872 (N_14872,N_13642,N_13611);
or U14873 (N_14873,N_13320,N_13638);
nor U14874 (N_14874,N_13403,N_13873);
nand U14875 (N_14875,N_13544,N_13859);
or U14876 (N_14876,N_13583,N_13018);
nand U14877 (N_14877,N_13694,N_13506);
or U14878 (N_14878,N_13609,N_13941);
and U14879 (N_14879,N_13524,N_13855);
nand U14880 (N_14880,N_13269,N_13452);
nor U14881 (N_14881,N_13290,N_13911);
nor U14882 (N_14882,N_13967,N_13666);
nand U14883 (N_14883,N_13704,N_13139);
and U14884 (N_14884,N_13750,N_13286);
and U14885 (N_14885,N_13002,N_13452);
or U14886 (N_14886,N_13398,N_13090);
nor U14887 (N_14887,N_13438,N_13789);
and U14888 (N_14888,N_13750,N_13801);
or U14889 (N_14889,N_13350,N_13234);
or U14890 (N_14890,N_13159,N_13515);
or U14891 (N_14891,N_13320,N_13255);
or U14892 (N_14892,N_13274,N_13095);
nor U14893 (N_14893,N_13996,N_13462);
nand U14894 (N_14894,N_13472,N_13195);
or U14895 (N_14895,N_13517,N_13433);
or U14896 (N_14896,N_13689,N_13558);
and U14897 (N_14897,N_13845,N_13501);
or U14898 (N_14898,N_13685,N_13556);
or U14899 (N_14899,N_13426,N_13526);
or U14900 (N_14900,N_13382,N_13764);
or U14901 (N_14901,N_13123,N_13204);
or U14902 (N_14902,N_13992,N_13277);
nand U14903 (N_14903,N_13215,N_13852);
nand U14904 (N_14904,N_13986,N_13805);
nand U14905 (N_14905,N_13157,N_13625);
or U14906 (N_14906,N_13537,N_13007);
nor U14907 (N_14907,N_13550,N_13698);
xor U14908 (N_14908,N_13414,N_13716);
nor U14909 (N_14909,N_13088,N_13828);
nand U14910 (N_14910,N_13456,N_13475);
and U14911 (N_14911,N_13430,N_13009);
xnor U14912 (N_14912,N_13460,N_13193);
or U14913 (N_14913,N_13144,N_13166);
and U14914 (N_14914,N_13818,N_13357);
or U14915 (N_14915,N_13387,N_13519);
and U14916 (N_14916,N_13964,N_13449);
nand U14917 (N_14917,N_13820,N_13199);
nand U14918 (N_14918,N_13530,N_13635);
nor U14919 (N_14919,N_13863,N_13055);
nor U14920 (N_14920,N_13837,N_13223);
and U14921 (N_14921,N_13645,N_13094);
nor U14922 (N_14922,N_13330,N_13005);
nor U14923 (N_14923,N_13134,N_13007);
and U14924 (N_14924,N_13449,N_13398);
and U14925 (N_14925,N_13004,N_13767);
nand U14926 (N_14926,N_13983,N_13685);
or U14927 (N_14927,N_13645,N_13937);
or U14928 (N_14928,N_13004,N_13622);
nor U14929 (N_14929,N_13065,N_13423);
nand U14930 (N_14930,N_13972,N_13105);
nor U14931 (N_14931,N_13765,N_13504);
and U14932 (N_14932,N_13452,N_13409);
and U14933 (N_14933,N_13392,N_13121);
nor U14934 (N_14934,N_13791,N_13740);
nor U14935 (N_14935,N_13827,N_13234);
and U14936 (N_14936,N_13423,N_13535);
and U14937 (N_14937,N_13543,N_13858);
nand U14938 (N_14938,N_13826,N_13023);
nor U14939 (N_14939,N_13493,N_13599);
nand U14940 (N_14940,N_13262,N_13782);
nor U14941 (N_14941,N_13047,N_13157);
or U14942 (N_14942,N_13207,N_13334);
nor U14943 (N_14943,N_13824,N_13014);
nor U14944 (N_14944,N_13909,N_13644);
or U14945 (N_14945,N_13153,N_13412);
and U14946 (N_14946,N_13363,N_13798);
or U14947 (N_14947,N_13280,N_13910);
or U14948 (N_14948,N_13390,N_13944);
and U14949 (N_14949,N_13610,N_13293);
and U14950 (N_14950,N_13032,N_13589);
nand U14951 (N_14951,N_13882,N_13044);
nor U14952 (N_14952,N_13324,N_13022);
nor U14953 (N_14953,N_13017,N_13538);
and U14954 (N_14954,N_13701,N_13652);
and U14955 (N_14955,N_13442,N_13489);
and U14956 (N_14956,N_13912,N_13811);
or U14957 (N_14957,N_13397,N_13871);
nor U14958 (N_14958,N_13186,N_13148);
or U14959 (N_14959,N_13667,N_13600);
nor U14960 (N_14960,N_13757,N_13754);
nor U14961 (N_14961,N_13844,N_13163);
or U14962 (N_14962,N_13952,N_13135);
nor U14963 (N_14963,N_13527,N_13703);
nand U14964 (N_14964,N_13669,N_13834);
and U14965 (N_14965,N_13446,N_13007);
or U14966 (N_14966,N_13464,N_13891);
nor U14967 (N_14967,N_13004,N_13531);
or U14968 (N_14968,N_13092,N_13908);
and U14969 (N_14969,N_13248,N_13563);
nor U14970 (N_14970,N_13674,N_13271);
or U14971 (N_14971,N_13714,N_13195);
nor U14972 (N_14972,N_13563,N_13479);
or U14973 (N_14973,N_13805,N_13528);
or U14974 (N_14974,N_13915,N_13071);
and U14975 (N_14975,N_13961,N_13194);
and U14976 (N_14976,N_13237,N_13660);
xor U14977 (N_14977,N_13448,N_13649);
or U14978 (N_14978,N_13265,N_13973);
or U14979 (N_14979,N_13221,N_13956);
nor U14980 (N_14980,N_13635,N_13911);
nand U14981 (N_14981,N_13470,N_13037);
or U14982 (N_14982,N_13110,N_13828);
nor U14983 (N_14983,N_13984,N_13396);
and U14984 (N_14984,N_13114,N_13783);
nand U14985 (N_14985,N_13971,N_13125);
nor U14986 (N_14986,N_13842,N_13073);
and U14987 (N_14987,N_13465,N_13289);
nand U14988 (N_14988,N_13190,N_13509);
nand U14989 (N_14989,N_13434,N_13356);
nand U14990 (N_14990,N_13586,N_13932);
nand U14991 (N_14991,N_13016,N_13999);
nor U14992 (N_14992,N_13074,N_13399);
or U14993 (N_14993,N_13684,N_13178);
nand U14994 (N_14994,N_13960,N_13540);
nand U14995 (N_14995,N_13107,N_13930);
nor U14996 (N_14996,N_13378,N_13558);
and U14997 (N_14997,N_13893,N_13531);
or U14998 (N_14998,N_13909,N_13330);
or U14999 (N_14999,N_13153,N_13456);
or UO_0 (O_0,N_14913,N_14246);
nor UO_1 (O_1,N_14344,N_14073);
and UO_2 (O_2,N_14061,N_14728);
and UO_3 (O_3,N_14651,N_14576);
or UO_4 (O_4,N_14461,N_14977);
nor UO_5 (O_5,N_14190,N_14726);
nand UO_6 (O_6,N_14599,N_14792);
and UO_7 (O_7,N_14942,N_14589);
nor UO_8 (O_8,N_14912,N_14544);
or UO_9 (O_9,N_14995,N_14313);
and UO_10 (O_10,N_14415,N_14055);
nand UO_11 (O_11,N_14616,N_14808);
and UO_12 (O_12,N_14564,N_14146);
or UO_13 (O_13,N_14189,N_14103);
or UO_14 (O_14,N_14681,N_14192);
nor UO_15 (O_15,N_14251,N_14637);
nand UO_16 (O_16,N_14868,N_14172);
nand UO_17 (O_17,N_14869,N_14840);
nand UO_18 (O_18,N_14794,N_14899);
nand UO_19 (O_19,N_14843,N_14734);
nand UO_20 (O_20,N_14428,N_14749);
or UO_21 (O_21,N_14937,N_14862);
nand UO_22 (O_22,N_14216,N_14758);
and UO_23 (O_23,N_14662,N_14908);
nor UO_24 (O_24,N_14691,N_14556);
and UO_25 (O_25,N_14279,N_14910);
or UO_26 (O_26,N_14183,N_14391);
nand UO_27 (O_27,N_14459,N_14892);
nor UO_28 (O_28,N_14583,N_14014);
nor UO_29 (O_29,N_14125,N_14443);
nor UO_30 (O_30,N_14557,N_14306);
nor UO_31 (O_31,N_14606,N_14767);
and UO_32 (O_32,N_14880,N_14904);
or UO_33 (O_33,N_14712,N_14200);
or UO_34 (O_34,N_14893,N_14374);
nor UO_35 (O_35,N_14204,N_14261);
nand UO_36 (O_36,N_14573,N_14741);
and UO_37 (O_37,N_14483,N_14960);
nor UO_38 (O_38,N_14439,N_14276);
nand UO_39 (O_39,N_14176,N_14225);
nand UO_40 (O_40,N_14480,N_14962);
or UO_41 (O_41,N_14837,N_14577);
and UO_42 (O_42,N_14881,N_14017);
nor UO_43 (O_43,N_14132,N_14581);
or UO_44 (O_44,N_14285,N_14911);
nor UO_45 (O_45,N_14708,N_14498);
or UO_46 (O_46,N_14610,N_14771);
nand UO_47 (O_47,N_14124,N_14926);
or UO_48 (O_48,N_14860,N_14412);
nand UO_49 (O_49,N_14765,N_14488);
and UO_50 (O_50,N_14803,N_14058);
and UO_51 (O_51,N_14468,N_14473);
nor UO_52 (O_52,N_14453,N_14381);
nor UO_53 (O_53,N_14947,N_14652);
nor UO_54 (O_54,N_14181,N_14250);
xor UO_55 (O_55,N_14955,N_14785);
nor UO_56 (O_56,N_14145,N_14368);
or UO_57 (O_57,N_14602,N_14989);
nand UO_58 (O_58,N_14545,N_14228);
or UO_59 (O_59,N_14232,N_14120);
or UO_60 (O_60,N_14224,N_14328);
nand UO_61 (O_61,N_14507,N_14865);
nor UO_62 (O_62,N_14431,N_14692);
or UO_63 (O_63,N_14160,N_14532);
nor UO_64 (O_64,N_14311,N_14565);
or UO_65 (O_65,N_14922,N_14586);
nor UO_66 (O_66,N_14738,N_14085);
or UO_67 (O_67,N_14781,N_14950);
nand UO_68 (O_68,N_14816,N_14856);
or UO_69 (O_69,N_14082,N_14535);
and UO_70 (O_70,N_14949,N_14541);
and UO_71 (O_71,N_14357,N_14713);
nor UO_72 (O_72,N_14740,N_14477);
or UO_73 (O_73,N_14594,N_14169);
and UO_74 (O_74,N_14819,N_14065);
or UO_75 (O_75,N_14370,N_14917);
or UO_76 (O_76,N_14575,N_14838);
and UO_77 (O_77,N_14288,N_14945);
nand UO_78 (O_78,N_14258,N_14171);
and UO_79 (O_79,N_14001,N_14292);
or UO_80 (O_80,N_14629,N_14976);
and UO_81 (O_81,N_14826,N_14495);
and UO_82 (O_82,N_14824,N_14627);
nor UO_83 (O_83,N_14915,N_14361);
or UO_84 (O_84,N_14158,N_14510);
or UO_85 (O_85,N_14919,N_14939);
and UO_86 (O_86,N_14509,N_14759);
and UO_87 (O_87,N_14798,N_14322);
nand UO_88 (O_88,N_14035,N_14552);
nor UO_89 (O_89,N_14965,N_14283);
or UO_90 (O_90,N_14555,N_14299);
and UO_91 (O_91,N_14486,N_14905);
nand UO_92 (O_92,N_14716,N_14973);
nor UO_93 (O_93,N_14804,N_14400);
nor UO_94 (O_94,N_14147,N_14191);
and UO_95 (O_95,N_14255,N_14677);
nor UO_96 (O_96,N_14502,N_14045);
and UO_97 (O_97,N_14175,N_14214);
nor UO_98 (O_98,N_14077,N_14018);
nor UO_99 (O_99,N_14458,N_14141);
nand UO_100 (O_100,N_14049,N_14828);
nand UO_101 (O_101,N_14793,N_14091);
or UO_102 (O_102,N_14857,N_14520);
nand UO_103 (O_103,N_14426,N_14332);
or UO_104 (O_104,N_14978,N_14605);
nor UO_105 (O_105,N_14956,N_14604);
and UO_106 (O_106,N_14847,N_14536);
and UO_107 (O_107,N_14992,N_14548);
nor UO_108 (O_108,N_14695,N_14517);
and UO_109 (O_109,N_14043,N_14966);
nand UO_110 (O_110,N_14151,N_14900);
and UO_111 (O_111,N_14506,N_14395);
nor UO_112 (O_112,N_14670,N_14199);
nor UO_113 (O_113,N_14696,N_14243);
nor UO_114 (O_114,N_14684,N_14230);
or UO_115 (O_115,N_14280,N_14571);
and UO_116 (O_116,N_14549,N_14036);
and UO_117 (O_117,N_14462,N_14801);
or UO_118 (O_118,N_14063,N_14252);
nor UO_119 (O_119,N_14115,N_14012);
and UO_120 (O_120,N_14388,N_14148);
nor UO_121 (O_121,N_14732,N_14830);
nor UO_122 (O_122,N_14729,N_14613);
nand UO_123 (O_123,N_14807,N_14156);
or UO_124 (O_124,N_14814,N_14831);
or UO_125 (O_125,N_14095,N_14409);
and UO_126 (O_126,N_14496,N_14471);
and UO_127 (O_127,N_14090,N_14825);
and UO_128 (O_128,N_14167,N_14647);
or UO_129 (O_129,N_14273,N_14218);
nand UO_130 (O_130,N_14679,N_14354);
nand UO_131 (O_131,N_14187,N_14603);
and UO_132 (O_132,N_14705,N_14570);
or UO_133 (O_133,N_14072,N_14257);
and UO_134 (O_134,N_14088,N_14957);
nor UO_135 (O_135,N_14429,N_14855);
nor UO_136 (O_136,N_14229,N_14427);
nand UO_137 (O_137,N_14638,N_14419);
nand UO_138 (O_138,N_14274,N_14669);
nand UO_139 (O_139,N_14023,N_14641);
nand UO_140 (O_140,N_14936,N_14051);
and UO_141 (O_141,N_14558,N_14797);
or UO_142 (O_142,N_14524,N_14430);
or UO_143 (O_143,N_14286,N_14263);
and UO_144 (O_144,N_14946,N_14326);
or UO_145 (O_145,N_14040,N_14236);
nand UO_146 (O_146,N_14630,N_14657);
nand UO_147 (O_147,N_14475,N_14454);
nand UO_148 (O_148,N_14970,N_14013);
nor UO_149 (O_149,N_14347,N_14397);
and UO_150 (O_150,N_14991,N_14408);
nor UO_151 (O_151,N_14128,N_14987);
nand UO_152 (O_152,N_14423,N_14940);
nor UO_153 (O_153,N_14437,N_14163);
and UO_154 (O_154,N_14059,N_14247);
nand UO_155 (O_155,N_14711,N_14592);
nand UO_156 (O_156,N_14827,N_14206);
or UO_157 (O_157,N_14634,N_14964);
and UO_158 (O_158,N_14126,N_14746);
or UO_159 (O_159,N_14673,N_14944);
and UO_160 (O_160,N_14866,N_14337);
and UO_161 (O_161,N_14240,N_14667);
or UO_162 (O_162,N_14778,N_14752);
or UO_163 (O_163,N_14829,N_14626);
nand UO_164 (O_164,N_14898,N_14399);
nor UO_165 (O_165,N_14584,N_14319);
nor UO_166 (O_166,N_14254,N_14514);
nand UO_167 (O_167,N_14852,N_14658);
nand UO_168 (O_168,N_14725,N_14390);
nand UO_169 (O_169,N_14440,N_14710);
nor UO_170 (O_170,N_14587,N_14002);
and UO_171 (O_171,N_14513,N_14757);
nor UO_172 (O_172,N_14364,N_14188);
or UO_173 (O_173,N_14007,N_14559);
nand UO_174 (O_174,N_14053,N_14984);
or UO_175 (O_175,N_14024,N_14476);
nor UO_176 (O_176,N_14542,N_14444);
and UO_177 (O_177,N_14918,N_14567);
nand UO_178 (O_178,N_14371,N_14810);
nor UO_179 (O_179,N_14968,N_14066);
or UO_180 (O_180,N_14972,N_14521);
or UO_181 (O_181,N_14052,N_14293);
or UO_182 (O_182,N_14008,N_14467);
nor UO_183 (O_183,N_14452,N_14446);
nor UO_184 (O_184,N_14133,N_14341);
and UO_185 (O_185,N_14231,N_14432);
and UO_186 (O_186,N_14340,N_14135);
and UO_187 (O_187,N_14877,N_14709);
nand UO_188 (O_188,N_14553,N_14974);
nand UO_189 (O_189,N_14718,N_14201);
or UO_190 (O_190,N_14220,N_14403);
and UO_191 (O_191,N_14447,N_14504);
or UO_192 (O_192,N_14768,N_14064);
nor UO_193 (O_193,N_14723,N_14727);
nand UO_194 (O_194,N_14215,N_14821);
nor UO_195 (O_195,N_14068,N_14401);
nand UO_196 (O_196,N_14533,N_14178);
nand UO_197 (O_197,N_14245,N_14435);
and UO_198 (O_198,N_14259,N_14773);
nand UO_199 (O_199,N_14472,N_14766);
nand UO_200 (O_200,N_14796,N_14083);
or UO_201 (O_201,N_14697,N_14282);
or UO_202 (O_202,N_14875,N_14348);
nand UO_203 (O_203,N_14092,N_14835);
or UO_204 (O_204,N_14086,N_14527);
or UO_205 (O_205,N_14318,N_14378);
or UO_206 (O_206,N_14621,N_14355);
and UO_207 (O_207,N_14154,N_14222);
nand UO_208 (O_208,N_14362,N_14591);
and UO_209 (O_209,N_14396,N_14130);
nand UO_210 (O_210,N_14844,N_14537);
nand UO_211 (O_211,N_14479,N_14704);
nor UO_212 (O_212,N_14924,N_14999);
or UO_213 (O_213,N_14101,N_14941);
and UO_214 (O_214,N_14717,N_14640);
nand UO_215 (O_215,N_14518,N_14003);
nor UO_216 (O_216,N_14170,N_14335);
nand UO_217 (O_217,N_14938,N_14887);
nor UO_218 (O_218,N_14470,N_14394);
nor UO_219 (O_219,N_14878,N_14384);
nor UO_220 (O_220,N_14817,N_14097);
or UO_221 (O_221,N_14047,N_14611);
and UO_222 (O_222,N_14031,N_14755);
and UO_223 (O_223,N_14117,N_14398);
nor UO_224 (O_224,N_14790,N_14168);
nor UO_225 (O_225,N_14566,N_14351);
and UO_226 (O_226,N_14237,N_14155);
and UO_227 (O_227,N_14096,N_14449);
and UO_228 (O_228,N_14886,N_14104);
nor UO_229 (O_229,N_14076,N_14223);
nor UO_230 (O_230,N_14295,N_14554);
or UO_231 (O_231,N_14490,N_14687);
nor UO_232 (O_232,N_14004,N_14349);
nand UO_233 (O_233,N_14813,N_14642);
nor UO_234 (O_234,N_14665,N_14563);
and UO_235 (O_235,N_14547,N_14593);
or UO_236 (O_236,N_14360,N_14159);
or UO_237 (O_237,N_14659,N_14182);
nor UO_238 (O_238,N_14574,N_14531);
nor UO_239 (O_239,N_14372,N_14572);
and UO_240 (O_240,N_14241,N_14753);
nand UO_241 (O_241,N_14455,N_14491);
nand UO_242 (O_242,N_14406,N_14497);
nor UO_243 (O_243,N_14540,N_14590);
and UO_244 (O_244,N_14850,N_14105);
nand UO_245 (O_245,N_14110,N_14027);
and UO_246 (O_246,N_14873,N_14721);
nand UO_247 (O_247,N_14656,N_14959);
and UO_248 (O_248,N_14754,N_14745);
or UO_249 (O_249,N_14839,N_14769);
nand UO_250 (O_250,N_14628,N_14208);
nand UO_251 (O_251,N_14811,N_14310);
and UO_252 (O_252,N_14682,N_14981);
nand UO_253 (O_253,N_14969,N_14038);
nand UO_254 (O_254,N_14056,N_14099);
nor UO_255 (O_255,N_14854,N_14832);
and UO_256 (O_256,N_14074,N_14668);
nand UO_257 (O_257,N_14456,N_14882);
nand UO_258 (O_258,N_14815,N_14661);
and UO_259 (O_259,N_14418,N_14935);
nand UO_260 (O_260,N_14762,N_14359);
nor UO_261 (O_261,N_14108,N_14737);
and UO_262 (O_262,N_14185,N_14300);
nor UO_263 (O_263,N_14515,N_14622);
nor UO_264 (O_264,N_14756,N_14791);
and UO_265 (O_265,N_14569,N_14127);
or UO_266 (O_266,N_14744,N_14943);
and UO_267 (O_267,N_14205,N_14909);
or UO_268 (O_268,N_14818,N_14482);
nor UO_269 (O_269,N_14242,N_14113);
nand UO_270 (O_270,N_14290,N_14526);
or UO_271 (O_271,N_14760,N_14660);
or UO_272 (O_272,N_14676,N_14150);
or UO_273 (O_273,N_14820,N_14932);
nor UO_274 (O_274,N_14304,N_14693);
nand UO_275 (O_275,N_14213,N_14783);
nand UO_276 (O_276,N_14275,N_14750);
xor UO_277 (O_277,N_14614,N_14806);
nand UO_278 (O_278,N_14193,N_14071);
and UO_279 (O_279,N_14078,N_14314);
nor UO_280 (O_280,N_14345,N_14469);
and UO_281 (O_281,N_14494,N_14358);
nor UO_282 (O_282,N_14450,N_14138);
and UO_283 (O_283,N_14902,N_14387);
and UO_284 (O_284,N_14339,N_14393);
and UO_285 (O_285,N_14980,N_14998);
nand UO_286 (O_286,N_14184,N_14625);
or UO_287 (O_287,N_14385,N_14897);
or UO_288 (O_288,N_14367,N_14683);
or UO_289 (O_289,N_14648,N_14863);
nand UO_290 (O_290,N_14874,N_14070);
and UO_291 (O_291,N_14107,N_14624);
and UO_292 (O_292,N_14645,N_14451);
nor UO_293 (O_293,N_14081,N_14075);
nor UO_294 (O_294,N_14649,N_14048);
or UO_295 (O_295,N_14841,N_14039);
and UO_296 (O_296,N_14853,N_14129);
and UO_297 (O_297,N_14975,N_14543);
or UO_298 (O_298,N_14149,N_14985);
nor UO_299 (O_299,N_14596,N_14060);
and UO_300 (O_300,N_14165,N_14896);
nor UO_301 (O_301,N_14032,N_14410);
nand UO_302 (O_302,N_14294,N_14884);
and UO_303 (O_303,N_14643,N_14689);
and UO_304 (O_304,N_14226,N_14080);
and UO_305 (O_305,N_14672,N_14353);
nor UO_306 (O_306,N_14463,N_14308);
or UO_307 (O_307,N_14329,N_14162);
nand UO_308 (O_308,N_14719,N_14595);
and UO_309 (O_309,N_14142,N_14883);
nor UO_310 (O_310,N_14383,N_14489);
or UO_311 (O_311,N_14098,N_14352);
or UO_312 (O_312,N_14493,N_14579);
nand UO_313 (O_313,N_14731,N_14281);
nand UO_314 (O_314,N_14993,N_14005);
nand UO_315 (O_315,N_14153,N_14457);
xnor UO_316 (O_316,N_14742,N_14789);
and UO_317 (O_317,N_14179,N_14029);
nor UO_318 (O_318,N_14607,N_14747);
or UO_319 (O_319,N_14788,N_14925);
and UO_320 (O_320,N_14928,N_14033);
or UO_321 (O_321,N_14139,N_14020);
nand UO_322 (O_322,N_14715,N_14538);
nand UO_323 (O_323,N_14441,N_14889);
or UO_324 (O_324,N_14519,N_14685);
nor UO_325 (O_325,N_14414,N_14864);
and UO_326 (O_326,N_14588,N_14653);
and UO_327 (O_327,N_14177,N_14923);
nand UO_328 (O_328,N_14842,N_14774);
and UO_329 (O_329,N_14365,N_14617);
nand UO_330 (O_330,N_14478,N_14407);
or UO_331 (O_331,N_14094,N_14356);
or UO_332 (O_332,N_14872,N_14694);
nor UO_333 (O_333,N_14166,N_14934);
nand UO_334 (O_334,N_14380,N_14334);
nor UO_335 (O_335,N_14623,N_14324);
nor UO_336 (O_336,N_14421,N_14688);
nand UO_337 (O_337,N_14777,N_14775);
nor UO_338 (O_338,N_14265,N_14674);
and UO_339 (O_339,N_14833,N_14028);
nand UO_340 (O_340,N_14582,N_14982);
and UO_341 (O_341,N_14748,N_14903);
or UO_342 (O_342,N_14363,N_14174);
or UO_343 (O_343,N_14289,N_14404);
or UO_344 (O_344,N_14198,N_14784);
nor UO_345 (O_345,N_14500,N_14448);
nand UO_346 (O_346,N_14823,N_14210);
or UO_347 (O_347,N_14000,N_14119);
or UO_348 (O_348,N_14046,N_14870);
nor UO_349 (O_349,N_14834,N_14876);
and UO_350 (O_350,N_14666,N_14221);
and UO_351 (O_351,N_14851,N_14284);
nand UO_352 (O_352,N_14111,N_14631);
and UO_353 (O_353,N_14100,N_14079);
and UO_354 (O_354,N_14822,N_14994);
nor UO_355 (O_355,N_14867,N_14597);
and UO_356 (O_356,N_14618,N_14485);
or UO_357 (O_357,N_14933,N_14433);
nand UO_358 (O_358,N_14173,N_14425);
and UO_359 (O_359,N_14836,N_14022);
and UO_360 (O_360,N_14118,N_14633);
nor UO_361 (O_361,N_14157,N_14186);
nor UO_362 (O_362,N_14010,N_14296);
nand UO_363 (O_363,N_14654,N_14131);
and UO_364 (O_364,N_14009,N_14511);
and UO_365 (O_365,N_14802,N_14015);
nand UO_366 (O_366,N_14202,N_14366);
or UO_367 (O_367,N_14207,N_14327);
or UO_368 (O_368,N_14140,N_14516);
or UO_369 (O_369,N_14735,N_14849);
nand UO_370 (O_370,N_14442,N_14405);
and UO_371 (O_371,N_14266,N_14305);
and UO_372 (O_372,N_14116,N_14782);
or UO_373 (O_373,N_14297,N_14639);
or UO_374 (O_374,N_14260,N_14392);
nand UO_375 (O_375,N_14499,N_14894);
nor UO_376 (O_376,N_14248,N_14707);
nor UO_377 (O_377,N_14346,N_14787);
or UO_378 (O_378,N_14143,N_14612);
nor UO_379 (O_379,N_14699,N_14505);
nor UO_380 (O_380,N_14278,N_14436);
nor UO_381 (O_381,N_14675,N_14523);
or UO_382 (O_382,N_14786,N_14264);
or UO_383 (O_383,N_14585,N_14233);
nor UO_384 (O_384,N_14799,N_14663);
nor UO_385 (O_385,N_14508,N_14312);
nand UO_386 (O_386,N_14763,N_14800);
nand UO_387 (O_387,N_14619,N_14315);
nand UO_388 (O_388,N_14194,N_14011);
or UO_389 (O_389,N_14698,N_14320);
nand UO_390 (O_390,N_14434,N_14714);
nand UO_391 (O_391,N_14733,N_14620);
nor UO_392 (O_392,N_14069,N_14761);
nand UO_393 (O_393,N_14244,N_14958);
or UO_394 (O_394,N_14212,N_14382);
nor UO_395 (O_395,N_14309,N_14891);
or UO_396 (O_396,N_14701,N_14920);
or UO_397 (O_397,N_14019,N_14379);
nand UO_398 (O_398,N_14376,N_14227);
and UO_399 (O_399,N_14287,N_14460);
and UO_400 (O_400,N_14650,N_14034);
and UO_401 (O_401,N_14234,N_14988);
nand UO_402 (O_402,N_14343,N_14256);
and UO_403 (O_403,N_14720,N_14528);
nor UO_404 (O_404,N_14375,N_14809);
nor UO_405 (O_405,N_14269,N_14780);
nand UO_406 (O_406,N_14635,N_14333);
or UO_407 (O_407,N_14861,N_14580);
and UO_408 (O_408,N_14961,N_14986);
xor UO_409 (O_409,N_14772,N_14921);
nor UO_410 (O_410,N_14338,N_14764);
nand UO_411 (O_411,N_14466,N_14044);
and UO_412 (O_412,N_14180,N_14812);
and UO_413 (O_413,N_14914,N_14568);
and UO_414 (O_414,N_14953,N_14253);
and UO_415 (O_415,N_14901,N_14690);
nand UO_416 (O_416,N_14026,N_14235);
and UO_417 (O_417,N_14601,N_14562);
or UO_418 (O_418,N_14386,N_14195);
or UO_419 (O_419,N_14655,N_14238);
and UO_420 (O_420,N_14369,N_14239);
nand UO_421 (O_421,N_14530,N_14330);
or UO_422 (O_422,N_14770,N_14416);
nand UO_423 (O_423,N_14736,N_14931);
nor UO_424 (O_424,N_14951,N_14561);
nand UO_425 (O_425,N_14331,N_14102);
nor UO_426 (O_426,N_14885,N_14703);
or UO_427 (O_427,N_14465,N_14030);
and UO_428 (O_428,N_14967,N_14323);
or UO_429 (O_429,N_14219,N_14929);
nand UO_430 (O_430,N_14271,N_14492);
and UO_431 (O_431,N_14203,N_14211);
nor UO_432 (O_432,N_14021,N_14109);
nor UO_433 (O_433,N_14417,N_14680);
xnor UO_434 (O_434,N_14578,N_14664);
or UO_435 (O_435,N_14445,N_14895);
and UO_436 (O_436,N_14779,N_14996);
nor UO_437 (O_437,N_14871,N_14122);
and UO_438 (O_438,N_14730,N_14845);
or UO_439 (O_439,N_14751,N_14413);
nand UO_440 (O_440,N_14084,N_14859);
or UO_441 (O_441,N_14979,N_14106);
and UO_442 (O_442,N_14301,N_14700);
and UO_443 (O_443,N_14927,N_14302);
or UO_444 (O_444,N_14144,N_14722);
or UO_445 (O_445,N_14411,N_14298);
nand UO_446 (O_446,N_14671,N_14137);
nor UO_447 (O_447,N_14686,N_14529);
nor UO_448 (O_448,N_14481,N_14424);
xnor UO_449 (O_449,N_14609,N_14983);
or UO_450 (O_450,N_14888,N_14350);
nand UO_451 (O_451,N_14632,N_14534);
and UO_452 (O_452,N_14890,N_14501);
nor UO_453 (O_453,N_14041,N_14474);
or UO_454 (O_454,N_14805,N_14307);
and UO_455 (O_455,N_14420,N_14316);
or UO_456 (O_456,N_14724,N_14776);
nor UO_457 (O_457,N_14196,N_14551);
and UO_458 (O_458,N_14487,N_14121);
nor UO_459 (O_459,N_14858,N_14217);
nor UO_460 (O_460,N_14270,N_14321);
or UO_461 (O_461,N_14291,N_14795);
and UO_462 (O_462,N_14123,N_14948);
nand UO_463 (O_463,N_14016,N_14152);
nand UO_464 (O_464,N_14997,N_14743);
nand UO_465 (O_465,N_14646,N_14209);
nand UO_466 (O_466,N_14025,N_14164);
nor UO_467 (O_467,N_14037,N_14336);
or UO_468 (O_468,N_14636,N_14525);
and UO_469 (O_469,N_14267,N_14054);
or UO_470 (O_470,N_14615,N_14389);
and UO_471 (O_471,N_14006,N_14268);
or UO_472 (O_472,N_14560,N_14550);
and UO_473 (O_473,N_14042,N_14971);
nor UO_474 (O_474,N_14057,N_14303);
and UO_475 (O_475,N_14050,N_14678);
or UO_476 (O_476,N_14916,N_14963);
nand UO_477 (O_477,N_14249,N_14503);
nand UO_478 (O_478,N_14484,N_14317);
nor UO_479 (O_479,N_14402,N_14134);
or UO_480 (O_480,N_14087,N_14277);
or UO_481 (O_481,N_14608,N_14067);
nand UO_482 (O_482,N_14422,N_14262);
and UO_483 (O_483,N_14093,N_14952);
nor UO_484 (O_484,N_14272,N_14325);
nor UO_485 (O_485,N_14342,N_14438);
nor UO_486 (O_486,N_14906,N_14114);
nand UO_487 (O_487,N_14600,N_14546);
nand UO_488 (O_488,N_14907,N_14089);
xor UO_489 (O_489,N_14706,N_14377);
or UO_490 (O_490,N_14112,N_14522);
and UO_491 (O_491,N_14954,N_14062);
and UO_492 (O_492,N_14930,N_14990);
or UO_493 (O_493,N_14373,N_14846);
and UO_494 (O_494,N_14197,N_14848);
nor UO_495 (O_495,N_14539,N_14161);
nand UO_496 (O_496,N_14702,N_14644);
and UO_497 (O_497,N_14464,N_14136);
or UO_498 (O_498,N_14512,N_14598);
and UO_499 (O_499,N_14739,N_14879);
or UO_500 (O_500,N_14883,N_14330);
and UO_501 (O_501,N_14624,N_14985);
and UO_502 (O_502,N_14234,N_14745);
nand UO_503 (O_503,N_14501,N_14182);
nand UO_504 (O_504,N_14556,N_14580);
nand UO_505 (O_505,N_14034,N_14882);
or UO_506 (O_506,N_14192,N_14260);
or UO_507 (O_507,N_14821,N_14304);
xnor UO_508 (O_508,N_14249,N_14081);
nor UO_509 (O_509,N_14680,N_14052);
nand UO_510 (O_510,N_14904,N_14445);
nor UO_511 (O_511,N_14415,N_14947);
nor UO_512 (O_512,N_14885,N_14220);
nand UO_513 (O_513,N_14644,N_14793);
or UO_514 (O_514,N_14034,N_14289);
nor UO_515 (O_515,N_14705,N_14477);
nand UO_516 (O_516,N_14942,N_14917);
and UO_517 (O_517,N_14920,N_14459);
nand UO_518 (O_518,N_14541,N_14583);
nand UO_519 (O_519,N_14262,N_14429);
or UO_520 (O_520,N_14083,N_14560);
or UO_521 (O_521,N_14702,N_14983);
nand UO_522 (O_522,N_14429,N_14932);
nand UO_523 (O_523,N_14116,N_14777);
nand UO_524 (O_524,N_14987,N_14415);
nand UO_525 (O_525,N_14851,N_14697);
nor UO_526 (O_526,N_14236,N_14977);
or UO_527 (O_527,N_14832,N_14644);
nor UO_528 (O_528,N_14721,N_14337);
or UO_529 (O_529,N_14759,N_14057);
nand UO_530 (O_530,N_14340,N_14884);
and UO_531 (O_531,N_14536,N_14812);
or UO_532 (O_532,N_14820,N_14314);
nor UO_533 (O_533,N_14499,N_14341);
nand UO_534 (O_534,N_14683,N_14650);
or UO_535 (O_535,N_14811,N_14972);
nand UO_536 (O_536,N_14065,N_14130);
or UO_537 (O_537,N_14159,N_14117);
nand UO_538 (O_538,N_14572,N_14525);
nand UO_539 (O_539,N_14742,N_14819);
or UO_540 (O_540,N_14225,N_14839);
nand UO_541 (O_541,N_14353,N_14478);
and UO_542 (O_542,N_14149,N_14980);
and UO_543 (O_543,N_14725,N_14680);
and UO_544 (O_544,N_14539,N_14214);
nand UO_545 (O_545,N_14750,N_14405);
nand UO_546 (O_546,N_14914,N_14680);
nor UO_547 (O_547,N_14630,N_14440);
nand UO_548 (O_548,N_14183,N_14690);
and UO_549 (O_549,N_14423,N_14072);
or UO_550 (O_550,N_14316,N_14095);
and UO_551 (O_551,N_14086,N_14557);
or UO_552 (O_552,N_14451,N_14734);
nor UO_553 (O_553,N_14561,N_14104);
nand UO_554 (O_554,N_14105,N_14873);
or UO_555 (O_555,N_14828,N_14759);
nor UO_556 (O_556,N_14336,N_14310);
nand UO_557 (O_557,N_14626,N_14780);
nand UO_558 (O_558,N_14437,N_14814);
nor UO_559 (O_559,N_14940,N_14694);
or UO_560 (O_560,N_14520,N_14462);
or UO_561 (O_561,N_14576,N_14352);
nand UO_562 (O_562,N_14341,N_14763);
nand UO_563 (O_563,N_14178,N_14488);
and UO_564 (O_564,N_14136,N_14682);
and UO_565 (O_565,N_14193,N_14543);
nor UO_566 (O_566,N_14111,N_14363);
xor UO_567 (O_567,N_14668,N_14783);
nor UO_568 (O_568,N_14203,N_14209);
or UO_569 (O_569,N_14987,N_14590);
nand UO_570 (O_570,N_14858,N_14663);
and UO_571 (O_571,N_14491,N_14666);
nand UO_572 (O_572,N_14747,N_14440);
nand UO_573 (O_573,N_14725,N_14481);
or UO_574 (O_574,N_14888,N_14847);
and UO_575 (O_575,N_14105,N_14642);
nand UO_576 (O_576,N_14193,N_14446);
and UO_577 (O_577,N_14343,N_14566);
nand UO_578 (O_578,N_14066,N_14597);
nor UO_579 (O_579,N_14825,N_14531);
and UO_580 (O_580,N_14077,N_14140);
and UO_581 (O_581,N_14083,N_14288);
nand UO_582 (O_582,N_14213,N_14202);
or UO_583 (O_583,N_14351,N_14752);
nand UO_584 (O_584,N_14028,N_14394);
and UO_585 (O_585,N_14035,N_14788);
or UO_586 (O_586,N_14516,N_14475);
nand UO_587 (O_587,N_14825,N_14188);
or UO_588 (O_588,N_14751,N_14230);
nor UO_589 (O_589,N_14105,N_14495);
nor UO_590 (O_590,N_14665,N_14902);
or UO_591 (O_591,N_14567,N_14429);
nand UO_592 (O_592,N_14684,N_14681);
and UO_593 (O_593,N_14413,N_14861);
or UO_594 (O_594,N_14217,N_14018);
nor UO_595 (O_595,N_14913,N_14688);
and UO_596 (O_596,N_14983,N_14996);
or UO_597 (O_597,N_14351,N_14180);
nor UO_598 (O_598,N_14942,N_14505);
or UO_599 (O_599,N_14714,N_14885);
nor UO_600 (O_600,N_14970,N_14968);
nand UO_601 (O_601,N_14636,N_14688);
or UO_602 (O_602,N_14191,N_14555);
and UO_603 (O_603,N_14469,N_14539);
nor UO_604 (O_604,N_14712,N_14781);
and UO_605 (O_605,N_14089,N_14026);
and UO_606 (O_606,N_14529,N_14287);
and UO_607 (O_607,N_14645,N_14285);
or UO_608 (O_608,N_14983,N_14857);
and UO_609 (O_609,N_14080,N_14923);
nor UO_610 (O_610,N_14545,N_14308);
or UO_611 (O_611,N_14864,N_14057);
nor UO_612 (O_612,N_14815,N_14262);
nand UO_613 (O_613,N_14872,N_14424);
and UO_614 (O_614,N_14142,N_14618);
nand UO_615 (O_615,N_14665,N_14337);
nand UO_616 (O_616,N_14877,N_14065);
or UO_617 (O_617,N_14883,N_14268);
and UO_618 (O_618,N_14249,N_14353);
nor UO_619 (O_619,N_14996,N_14205);
nand UO_620 (O_620,N_14089,N_14970);
and UO_621 (O_621,N_14271,N_14049);
or UO_622 (O_622,N_14054,N_14729);
nand UO_623 (O_623,N_14006,N_14789);
and UO_624 (O_624,N_14902,N_14184);
or UO_625 (O_625,N_14781,N_14999);
nand UO_626 (O_626,N_14596,N_14804);
nand UO_627 (O_627,N_14687,N_14316);
nand UO_628 (O_628,N_14882,N_14800);
nand UO_629 (O_629,N_14326,N_14007);
and UO_630 (O_630,N_14687,N_14440);
or UO_631 (O_631,N_14369,N_14278);
nand UO_632 (O_632,N_14703,N_14178);
or UO_633 (O_633,N_14322,N_14864);
nor UO_634 (O_634,N_14188,N_14501);
nor UO_635 (O_635,N_14944,N_14591);
nand UO_636 (O_636,N_14536,N_14927);
or UO_637 (O_637,N_14302,N_14442);
nand UO_638 (O_638,N_14115,N_14220);
and UO_639 (O_639,N_14200,N_14118);
nand UO_640 (O_640,N_14938,N_14805);
and UO_641 (O_641,N_14496,N_14114);
nor UO_642 (O_642,N_14640,N_14212);
or UO_643 (O_643,N_14158,N_14460);
and UO_644 (O_644,N_14140,N_14821);
and UO_645 (O_645,N_14270,N_14595);
nand UO_646 (O_646,N_14790,N_14702);
and UO_647 (O_647,N_14809,N_14936);
nor UO_648 (O_648,N_14559,N_14989);
nand UO_649 (O_649,N_14286,N_14193);
nand UO_650 (O_650,N_14242,N_14067);
nand UO_651 (O_651,N_14253,N_14758);
and UO_652 (O_652,N_14557,N_14481);
and UO_653 (O_653,N_14105,N_14970);
and UO_654 (O_654,N_14810,N_14495);
and UO_655 (O_655,N_14611,N_14850);
nand UO_656 (O_656,N_14155,N_14706);
nand UO_657 (O_657,N_14510,N_14340);
nand UO_658 (O_658,N_14175,N_14893);
and UO_659 (O_659,N_14450,N_14216);
and UO_660 (O_660,N_14383,N_14511);
and UO_661 (O_661,N_14568,N_14726);
nand UO_662 (O_662,N_14713,N_14013);
nor UO_663 (O_663,N_14156,N_14459);
or UO_664 (O_664,N_14161,N_14834);
nor UO_665 (O_665,N_14941,N_14408);
and UO_666 (O_666,N_14968,N_14988);
and UO_667 (O_667,N_14013,N_14693);
and UO_668 (O_668,N_14156,N_14087);
or UO_669 (O_669,N_14880,N_14686);
nor UO_670 (O_670,N_14280,N_14821);
nand UO_671 (O_671,N_14164,N_14365);
nor UO_672 (O_672,N_14842,N_14280);
nand UO_673 (O_673,N_14992,N_14189);
nand UO_674 (O_674,N_14510,N_14759);
or UO_675 (O_675,N_14892,N_14422);
nand UO_676 (O_676,N_14711,N_14351);
or UO_677 (O_677,N_14986,N_14870);
and UO_678 (O_678,N_14503,N_14845);
and UO_679 (O_679,N_14603,N_14754);
and UO_680 (O_680,N_14884,N_14692);
nor UO_681 (O_681,N_14639,N_14906);
and UO_682 (O_682,N_14746,N_14065);
nand UO_683 (O_683,N_14728,N_14887);
or UO_684 (O_684,N_14178,N_14456);
nand UO_685 (O_685,N_14397,N_14352);
nand UO_686 (O_686,N_14259,N_14050);
and UO_687 (O_687,N_14735,N_14863);
or UO_688 (O_688,N_14100,N_14195);
or UO_689 (O_689,N_14657,N_14454);
and UO_690 (O_690,N_14894,N_14686);
nand UO_691 (O_691,N_14677,N_14877);
or UO_692 (O_692,N_14168,N_14436);
or UO_693 (O_693,N_14349,N_14924);
xor UO_694 (O_694,N_14329,N_14141);
nand UO_695 (O_695,N_14888,N_14177);
and UO_696 (O_696,N_14516,N_14492);
xnor UO_697 (O_697,N_14596,N_14702);
nand UO_698 (O_698,N_14958,N_14948);
nand UO_699 (O_699,N_14598,N_14385);
or UO_700 (O_700,N_14085,N_14029);
and UO_701 (O_701,N_14099,N_14037);
and UO_702 (O_702,N_14716,N_14540);
and UO_703 (O_703,N_14230,N_14558);
or UO_704 (O_704,N_14746,N_14379);
or UO_705 (O_705,N_14680,N_14718);
and UO_706 (O_706,N_14690,N_14976);
or UO_707 (O_707,N_14051,N_14787);
nand UO_708 (O_708,N_14526,N_14505);
or UO_709 (O_709,N_14128,N_14516);
nand UO_710 (O_710,N_14653,N_14308);
and UO_711 (O_711,N_14255,N_14195);
or UO_712 (O_712,N_14949,N_14103);
nor UO_713 (O_713,N_14748,N_14895);
nor UO_714 (O_714,N_14512,N_14765);
or UO_715 (O_715,N_14897,N_14708);
or UO_716 (O_716,N_14457,N_14709);
nand UO_717 (O_717,N_14057,N_14807);
nor UO_718 (O_718,N_14181,N_14490);
nand UO_719 (O_719,N_14702,N_14158);
or UO_720 (O_720,N_14726,N_14359);
or UO_721 (O_721,N_14203,N_14037);
and UO_722 (O_722,N_14710,N_14717);
or UO_723 (O_723,N_14537,N_14670);
or UO_724 (O_724,N_14705,N_14595);
and UO_725 (O_725,N_14503,N_14546);
nor UO_726 (O_726,N_14354,N_14044);
nand UO_727 (O_727,N_14145,N_14923);
nand UO_728 (O_728,N_14259,N_14646);
nor UO_729 (O_729,N_14641,N_14447);
or UO_730 (O_730,N_14269,N_14863);
nand UO_731 (O_731,N_14869,N_14047);
and UO_732 (O_732,N_14618,N_14934);
nor UO_733 (O_733,N_14473,N_14815);
or UO_734 (O_734,N_14367,N_14247);
or UO_735 (O_735,N_14249,N_14132);
or UO_736 (O_736,N_14604,N_14298);
nor UO_737 (O_737,N_14700,N_14861);
nor UO_738 (O_738,N_14698,N_14147);
nor UO_739 (O_739,N_14094,N_14703);
nor UO_740 (O_740,N_14275,N_14339);
or UO_741 (O_741,N_14804,N_14501);
nor UO_742 (O_742,N_14526,N_14291);
nand UO_743 (O_743,N_14768,N_14579);
and UO_744 (O_744,N_14898,N_14670);
or UO_745 (O_745,N_14198,N_14241);
nand UO_746 (O_746,N_14528,N_14331);
and UO_747 (O_747,N_14265,N_14271);
and UO_748 (O_748,N_14034,N_14422);
and UO_749 (O_749,N_14883,N_14612);
nor UO_750 (O_750,N_14149,N_14364);
nor UO_751 (O_751,N_14972,N_14538);
or UO_752 (O_752,N_14469,N_14494);
or UO_753 (O_753,N_14866,N_14715);
and UO_754 (O_754,N_14024,N_14303);
or UO_755 (O_755,N_14755,N_14364);
nor UO_756 (O_756,N_14036,N_14392);
nand UO_757 (O_757,N_14535,N_14275);
nand UO_758 (O_758,N_14284,N_14485);
or UO_759 (O_759,N_14387,N_14715);
nand UO_760 (O_760,N_14879,N_14733);
or UO_761 (O_761,N_14899,N_14801);
and UO_762 (O_762,N_14385,N_14530);
nor UO_763 (O_763,N_14554,N_14868);
nor UO_764 (O_764,N_14709,N_14708);
and UO_765 (O_765,N_14786,N_14278);
nor UO_766 (O_766,N_14175,N_14518);
and UO_767 (O_767,N_14857,N_14807);
nor UO_768 (O_768,N_14217,N_14276);
or UO_769 (O_769,N_14662,N_14053);
and UO_770 (O_770,N_14065,N_14720);
nand UO_771 (O_771,N_14986,N_14489);
nor UO_772 (O_772,N_14826,N_14916);
nor UO_773 (O_773,N_14037,N_14341);
or UO_774 (O_774,N_14827,N_14290);
nand UO_775 (O_775,N_14183,N_14352);
or UO_776 (O_776,N_14699,N_14979);
nand UO_777 (O_777,N_14596,N_14398);
and UO_778 (O_778,N_14627,N_14322);
and UO_779 (O_779,N_14249,N_14633);
nand UO_780 (O_780,N_14454,N_14557);
nor UO_781 (O_781,N_14766,N_14840);
nand UO_782 (O_782,N_14489,N_14761);
nand UO_783 (O_783,N_14670,N_14839);
and UO_784 (O_784,N_14740,N_14373);
and UO_785 (O_785,N_14473,N_14856);
or UO_786 (O_786,N_14142,N_14162);
or UO_787 (O_787,N_14652,N_14709);
and UO_788 (O_788,N_14172,N_14499);
and UO_789 (O_789,N_14506,N_14069);
or UO_790 (O_790,N_14072,N_14575);
or UO_791 (O_791,N_14342,N_14973);
or UO_792 (O_792,N_14579,N_14892);
and UO_793 (O_793,N_14380,N_14285);
and UO_794 (O_794,N_14899,N_14510);
nand UO_795 (O_795,N_14307,N_14892);
nor UO_796 (O_796,N_14641,N_14327);
and UO_797 (O_797,N_14374,N_14964);
nor UO_798 (O_798,N_14798,N_14774);
nor UO_799 (O_799,N_14416,N_14410);
nor UO_800 (O_800,N_14015,N_14712);
nand UO_801 (O_801,N_14701,N_14992);
or UO_802 (O_802,N_14182,N_14817);
or UO_803 (O_803,N_14962,N_14028);
nand UO_804 (O_804,N_14022,N_14804);
nor UO_805 (O_805,N_14573,N_14114);
nand UO_806 (O_806,N_14946,N_14564);
nor UO_807 (O_807,N_14001,N_14769);
nor UO_808 (O_808,N_14751,N_14626);
nor UO_809 (O_809,N_14196,N_14125);
or UO_810 (O_810,N_14739,N_14380);
and UO_811 (O_811,N_14610,N_14923);
nor UO_812 (O_812,N_14113,N_14934);
nand UO_813 (O_813,N_14562,N_14617);
and UO_814 (O_814,N_14519,N_14006);
nor UO_815 (O_815,N_14039,N_14157);
nor UO_816 (O_816,N_14319,N_14481);
and UO_817 (O_817,N_14987,N_14905);
nor UO_818 (O_818,N_14120,N_14737);
nand UO_819 (O_819,N_14401,N_14658);
or UO_820 (O_820,N_14077,N_14029);
or UO_821 (O_821,N_14644,N_14764);
nand UO_822 (O_822,N_14152,N_14222);
and UO_823 (O_823,N_14314,N_14210);
nor UO_824 (O_824,N_14373,N_14797);
or UO_825 (O_825,N_14773,N_14981);
nand UO_826 (O_826,N_14550,N_14648);
and UO_827 (O_827,N_14439,N_14605);
nor UO_828 (O_828,N_14349,N_14774);
nor UO_829 (O_829,N_14389,N_14872);
nor UO_830 (O_830,N_14734,N_14648);
nand UO_831 (O_831,N_14641,N_14844);
or UO_832 (O_832,N_14812,N_14225);
nand UO_833 (O_833,N_14512,N_14542);
or UO_834 (O_834,N_14289,N_14480);
or UO_835 (O_835,N_14629,N_14475);
nor UO_836 (O_836,N_14578,N_14207);
or UO_837 (O_837,N_14258,N_14115);
nor UO_838 (O_838,N_14636,N_14347);
nor UO_839 (O_839,N_14986,N_14634);
nor UO_840 (O_840,N_14839,N_14247);
and UO_841 (O_841,N_14793,N_14457);
and UO_842 (O_842,N_14578,N_14528);
and UO_843 (O_843,N_14306,N_14982);
nand UO_844 (O_844,N_14354,N_14749);
or UO_845 (O_845,N_14578,N_14977);
and UO_846 (O_846,N_14121,N_14268);
nor UO_847 (O_847,N_14868,N_14089);
nand UO_848 (O_848,N_14138,N_14061);
and UO_849 (O_849,N_14523,N_14279);
and UO_850 (O_850,N_14628,N_14802);
and UO_851 (O_851,N_14747,N_14353);
nor UO_852 (O_852,N_14487,N_14111);
and UO_853 (O_853,N_14062,N_14117);
and UO_854 (O_854,N_14844,N_14542);
or UO_855 (O_855,N_14694,N_14744);
nor UO_856 (O_856,N_14421,N_14126);
and UO_857 (O_857,N_14992,N_14984);
or UO_858 (O_858,N_14282,N_14511);
or UO_859 (O_859,N_14680,N_14664);
nor UO_860 (O_860,N_14135,N_14813);
and UO_861 (O_861,N_14544,N_14987);
or UO_862 (O_862,N_14413,N_14930);
nor UO_863 (O_863,N_14406,N_14336);
nand UO_864 (O_864,N_14202,N_14334);
nand UO_865 (O_865,N_14508,N_14977);
or UO_866 (O_866,N_14968,N_14948);
or UO_867 (O_867,N_14163,N_14869);
and UO_868 (O_868,N_14596,N_14727);
or UO_869 (O_869,N_14537,N_14781);
nor UO_870 (O_870,N_14963,N_14354);
nand UO_871 (O_871,N_14304,N_14542);
or UO_872 (O_872,N_14328,N_14766);
or UO_873 (O_873,N_14406,N_14078);
nand UO_874 (O_874,N_14059,N_14192);
and UO_875 (O_875,N_14878,N_14435);
or UO_876 (O_876,N_14592,N_14923);
and UO_877 (O_877,N_14889,N_14230);
or UO_878 (O_878,N_14679,N_14536);
nand UO_879 (O_879,N_14611,N_14459);
nor UO_880 (O_880,N_14043,N_14119);
nor UO_881 (O_881,N_14624,N_14989);
nor UO_882 (O_882,N_14521,N_14849);
nor UO_883 (O_883,N_14615,N_14937);
nand UO_884 (O_884,N_14589,N_14386);
nand UO_885 (O_885,N_14727,N_14945);
and UO_886 (O_886,N_14938,N_14962);
or UO_887 (O_887,N_14324,N_14619);
or UO_888 (O_888,N_14505,N_14730);
and UO_889 (O_889,N_14847,N_14864);
or UO_890 (O_890,N_14405,N_14606);
or UO_891 (O_891,N_14518,N_14070);
nand UO_892 (O_892,N_14737,N_14474);
and UO_893 (O_893,N_14108,N_14359);
nand UO_894 (O_894,N_14699,N_14106);
or UO_895 (O_895,N_14120,N_14040);
nand UO_896 (O_896,N_14570,N_14777);
or UO_897 (O_897,N_14653,N_14704);
nor UO_898 (O_898,N_14640,N_14227);
nand UO_899 (O_899,N_14452,N_14744);
or UO_900 (O_900,N_14606,N_14747);
and UO_901 (O_901,N_14740,N_14762);
nand UO_902 (O_902,N_14604,N_14227);
nor UO_903 (O_903,N_14484,N_14105);
or UO_904 (O_904,N_14328,N_14104);
nor UO_905 (O_905,N_14742,N_14848);
nand UO_906 (O_906,N_14614,N_14276);
nand UO_907 (O_907,N_14010,N_14503);
xor UO_908 (O_908,N_14854,N_14882);
nor UO_909 (O_909,N_14481,N_14887);
or UO_910 (O_910,N_14572,N_14324);
or UO_911 (O_911,N_14477,N_14303);
nand UO_912 (O_912,N_14205,N_14404);
and UO_913 (O_913,N_14530,N_14045);
nor UO_914 (O_914,N_14707,N_14636);
and UO_915 (O_915,N_14504,N_14643);
nor UO_916 (O_916,N_14720,N_14419);
nand UO_917 (O_917,N_14147,N_14508);
nand UO_918 (O_918,N_14587,N_14657);
and UO_919 (O_919,N_14191,N_14465);
nand UO_920 (O_920,N_14874,N_14400);
and UO_921 (O_921,N_14184,N_14338);
nand UO_922 (O_922,N_14820,N_14299);
or UO_923 (O_923,N_14070,N_14894);
or UO_924 (O_924,N_14203,N_14411);
nand UO_925 (O_925,N_14601,N_14420);
and UO_926 (O_926,N_14299,N_14521);
nand UO_927 (O_927,N_14291,N_14048);
and UO_928 (O_928,N_14562,N_14819);
nor UO_929 (O_929,N_14528,N_14003);
nand UO_930 (O_930,N_14100,N_14584);
nand UO_931 (O_931,N_14774,N_14226);
nand UO_932 (O_932,N_14523,N_14238);
nor UO_933 (O_933,N_14738,N_14594);
or UO_934 (O_934,N_14011,N_14727);
nand UO_935 (O_935,N_14969,N_14546);
nand UO_936 (O_936,N_14077,N_14895);
or UO_937 (O_937,N_14047,N_14174);
and UO_938 (O_938,N_14108,N_14377);
nand UO_939 (O_939,N_14704,N_14473);
nor UO_940 (O_940,N_14792,N_14328);
nor UO_941 (O_941,N_14363,N_14486);
nor UO_942 (O_942,N_14660,N_14977);
nand UO_943 (O_943,N_14506,N_14330);
nor UO_944 (O_944,N_14579,N_14036);
nor UO_945 (O_945,N_14086,N_14971);
nor UO_946 (O_946,N_14987,N_14654);
or UO_947 (O_947,N_14033,N_14951);
or UO_948 (O_948,N_14352,N_14085);
nor UO_949 (O_949,N_14885,N_14468);
nand UO_950 (O_950,N_14892,N_14314);
nand UO_951 (O_951,N_14806,N_14669);
and UO_952 (O_952,N_14251,N_14534);
nor UO_953 (O_953,N_14022,N_14661);
nand UO_954 (O_954,N_14544,N_14591);
nor UO_955 (O_955,N_14560,N_14459);
nand UO_956 (O_956,N_14732,N_14272);
nand UO_957 (O_957,N_14514,N_14259);
and UO_958 (O_958,N_14923,N_14903);
or UO_959 (O_959,N_14693,N_14991);
nand UO_960 (O_960,N_14208,N_14371);
or UO_961 (O_961,N_14786,N_14097);
nand UO_962 (O_962,N_14638,N_14845);
or UO_963 (O_963,N_14813,N_14224);
or UO_964 (O_964,N_14331,N_14256);
nor UO_965 (O_965,N_14659,N_14170);
nand UO_966 (O_966,N_14588,N_14279);
xor UO_967 (O_967,N_14454,N_14625);
nor UO_968 (O_968,N_14635,N_14402);
nand UO_969 (O_969,N_14362,N_14594);
or UO_970 (O_970,N_14822,N_14950);
nand UO_971 (O_971,N_14018,N_14762);
and UO_972 (O_972,N_14596,N_14156);
or UO_973 (O_973,N_14885,N_14321);
and UO_974 (O_974,N_14299,N_14890);
and UO_975 (O_975,N_14881,N_14604);
and UO_976 (O_976,N_14262,N_14222);
nor UO_977 (O_977,N_14934,N_14766);
xnor UO_978 (O_978,N_14295,N_14523);
or UO_979 (O_979,N_14223,N_14344);
nand UO_980 (O_980,N_14962,N_14144);
and UO_981 (O_981,N_14175,N_14966);
nand UO_982 (O_982,N_14720,N_14307);
nor UO_983 (O_983,N_14408,N_14174);
and UO_984 (O_984,N_14430,N_14584);
and UO_985 (O_985,N_14458,N_14662);
nand UO_986 (O_986,N_14084,N_14635);
nand UO_987 (O_987,N_14871,N_14582);
or UO_988 (O_988,N_14378,N_14138);
or UO_989 (O_989,N_14701,N_14634);
and UO_990 (O_990,N_14936,N_14844);
nor UO_991 (O_991,N_14553,N_14753);
and UO_992 (O_992,N_14600,N_14361);
nand UO_993 (O_993,N_14156,N_14812);
or UO_994 (O_994,N_14358,N_14651);
nand UO_995 (O_995,N_14014,N_14960);
nor UO_996 (O_996,N_14903,N_14559);
xor UO_997 (O_997,N_14159,N_14935);
nand UO_998 (O_998,N_14901,N_14156);
or UO_999 (O_999,N_14418,N_14351);
xnor UO_1000 (O_1000,N_14741,N_14756);
nor UO_1001 (O_1001,N_14843,N_14275);
nand UO_1002 (O_1002,N_14693,N_14676);
and UO_1003 (O_1003,N_14338,N_14728);
nor UO_1004 (O_1004,N_14572,N_14236);
or UO_1005 (O_1005,N_14150,N_14854);
or UO_1006 (O_1006,N_14347,N_14125);
nor UO_1007 (O_1007,N_14473,N_14267);
nand UO_1008 (O_1008,N_14716,N_14299);
nor UO_1009 (O_1009,N_14578,N_14038);
nor UO_1010 (O_1010,N_14364,N_14426);
or UO_1011 (O_1011,N_14726,N_14245);
or UO_1012 (O_1012,N_14216,N_14083);
and UO_1013 (O_1013,N_14655,N_14017);
or UO_1014 (O_1014,N_14970,N_14373);
nor UO_1015 (O_1015,N_14125,N_14593);
or UO_1016 (O_1016,N_14271,N_14178);
nor UO_1017 (O_1017,N_14979,N_14568);
and UO_1018 (O_1018,N_14682,N_14909);
and UO_1019 (O_1019,N_14413,N_14333);
nor UO_1020 (O_1020,N_14451,N_14587);
nand UO_1021 (O_1021,N_14538,N_14202);
nor UO_1022 (O_1022,N_14113,N_14416);
and UO_1023 (O_1023,N_14343,N_14600);
and UO_1024 (O_1024,N_14948,N_14060);
and UO_1025 (O_1025,N_14220,N_14204);
and UO_1026 (O_1026,N_14101,N_14386);
and UO_1027 (O_1027,N_14317,N_14489);
nor UO_1028 (O_1028,N_14116,N_14618);
and UO_1029 (O_1029,N_14840,N_14926);
nand UO_1030 (O_1030,N_14698,N_14758);
and UO_1031 (O_1031,N_14835,N_14687);
and UO_1032 (O_1032,N_14997,N_14196);
or UO_1033 (O_1033,N_14479,N_14380);
or UO_1034 (O_1034,N_14696,N_14286);
nor UO_1035 (O_1035,N_14502,N_14874);
nand UO_1036 (O_1036,N_14147,N_14581);
and UO_1037 (O_1037,N_14481,N_14395);
and UO_1038 (O_1038,N_14836,N_14074);
and UO_1039 (O_1039,N_14150,N_14657);
nand UO_1040 (O_1040,N_14051,N_14308);
or UO_1041 (O_1041,N_14592,N_14241);
nor UO_1042 (O_1042,N_14469,N_14051);
or UO_1043 (O_1043,N_14254,N_14537);
nor UO_1044 (O_1044,N_14156,N_14423);
nor UO_1045 (O_1045,N_14884,N_14934);
nand UO_1046 (O_1046,N_14416,N_14790);
nand UO_1047 (O_1047,N_14282,N_14074);
or UO_1048 (O_1048,N_14872,N_14280);
or UO_1049 (O_1049,N_14473,N_14504);
nor UO_1050 (O_1050,N_14293,N_14742);
nand UO_1051 (O_1051,N_14396,N_14194);
or UO_1052 (O_1052,N_14627,N_14113);
and UO_1053 (O_1053,N_14571,N_14195);
or UO_1054 (O_1054,N_14023,N_14105);
or UO_1055 (O_1055,N_14799,N_14851);
or UO_1056 (O_1056,N_14430,N_14229);
and UO_1057 (O_1057,N_14011,N_14942);
nor UO_1058 (O_1058,N_14973,N_14677);
nand UO_1059 (O_1059,N_14219,N_14927);
nand UO_1060 (O_1060,N_14571,N_14286);
and UO_1061 (O_1061,N_14479,N_14115);
and UO_1062 (O_1062,N_14672,N_14845);
nor UO_1063 (O_1063,N_14752,N_14289);
and UO_1064 (O_1064,N_14701,N_14376);
and UO_1065 (O_1065,N_14005,N_14050);
nor UO_1066 (O_1066,N_14126,N_14917);
nand UO_1067 (O_1067,N_14487,N_14742);
and UO_1068 (O_1068,N_14190,N_14140);
nor UO_1069 (O_1069,N_14278,N_14178);
nor UO_1070 (O_1070,N_14924,N_14946);
nand UO_1071 (O_1071,N_14913,N_14796);
or UO_1072 (O_1072,N_14000,N_14481);
nand UO_1073 (O_1073,N_14849,N_14070);
and UO_1074 (O_1074,N_14994,N_14974);
nor UO_1075 (O_1075,N_14658,N_14775);
nor UO_1076 (O_1076,N_14672,N_14149);
nor UO_1077 (O_1077,N_14271,N_14940);
or UO_1078 (O_1078,N_14651,N_14465);
or UO_1079 (O_1079,N_14571,N_14215);
nand UO_1080 (O_1080,N_14154,N_14785);
or UO_1081 (O_1081,N_14405,N_14538);
nand UO_1082 (O_1082,N_14859,N_14173);
nor UO_1083 (O_1083,N_14457,N_14596);
and UO_1084 (O_1084,N_14698,N_14176);
or UO_1085 (O_1085,N_14234,N_14765);
and UO_1086 (O_1086,N_14895,N_14313);
and UO_1087 (O_1087,N_14278,N_14782);
or UO_1088 (O_1088,N_14009,N_14873);
nand UO_1089 (O_1089,N_14656,N_14958);
nor UO_1090 (O_1090,N_14294,N_14185);
nor UO_1091 (O_1091,N_14160,N_14306);
nand UO_1092 (O_1092,N_14933,N_14443);
and UO_1093 (O_1093,N_14277,N_14403);
or UO_1094 (O_1094,N_14095,N_14983);
and UO_1095 (O_1095,N_14596,N_14540);
nand UO_1096 (O_1096,N_14517,N_14780);
nand UO_1097 (O_1097,N_14237,N_14987);
nand UO_1098 (O_1098,N_14535,N_14935);
nor UO_1099 (O_1099,N_14593,N_14319);
or UO_1100 (O_1100,N_14922,N_14594);
and UO_1101 (O_1101,N_14451,N_14327);
and UO_1102 (O_1102,N_14535,N_14665);
or UO_1103 (O_1103,N_14323,N_14560);
nand UO_1104 (O_1104,N_14366,N_14029);
nor UO_1105 (O_1105,N_14374,N_14600);
nor UO_1106 (O_1106,N_14567,N_14917);
nor UO_1107 (O_1107,N_14557,N_14337);
nor UO_1108 (O_1108,N_14173,N_14117);
nand UO_1109 (O_1109,N_14470,N_14347);
or UO_1110 (O_1110,N_14073,N_14695);
nor UO_1111 (O_1111,N_14238,N_14144);
nand UO_1112 (O_1112,N_14472,N_14113);
and UO_1113 (O_1113,N_14231,N_14070);
and UO_1114 (O_1114,N_14754,N_14709);
nand UO_1115 (O_1115,N_14245,N_14838);
nand UO_1116 (O_1116,N_14964,N_14823);
nand UO_1117 (O_1117,N_14131,N_14060);
and UO_1118 (O_1118,N_14730,N_14243);
nand UO_1119 (O_1119,N_14451,N_14777);
or UO_1120 (O_1120,N_14616,N_14114);
or UO_1121 (O_1121,N_14784,N_14916);
nand UO_1122 (O_1122,N_14802,N_14721);
nor UO_1123 (O_1123,N_14915,N_14538);
and UO_1124 (O_1124,N_14620,N_14346);
or UO_1125 (O_1125,N_14286,N_14651);
nor UO_1126 (O_1126,N_14819,N_14575);
nand UO_1127 (O_1127,N_14677,N_14491);
nand UO_1128 (O_1128,N_14857,N_14010);
nand UO_1129 (O_1129,N_14218,N_14612);
nor UO_1130 (O_1130,N_14040,N_14227);
nor UO_1131 (O_1131,N_14333,N_14192);
nand UO_1132 (O_1132,N_14105,N_14405);
nor UO_1133 (O_1133,N_14259,N_14692);
or UO_1134 (O_1134,N_14867,N_14437);
or UO_1135 (O_1135,N_14272,N_14226);
nor UO_1136 (O_1136,N_14402,N_14867);
nand UO_1137 (O_1137,N_14086,N_14477);
or UO_1138 (O_1138,N_14314,N_14357);
nor UO_1139 (O_1139,N_14413,N_14587);
or UO_1140 (O_1140,N_14670,N_14062);
nand UO_1141 (O_1141,N_14032,N_14838);
nand UO_1142 (O_1142,N_14799,N_14426);
nor UO_1143 (O_1143,N_14406,N_14540);
or UO_1144 (O_1144,N_14823,N_14829);
or UO_1145 (O_1145,N_14601,N_14736);
nand UO_1146 (O_1146,N_14172,N_14430);
or UO_1147 (O_1147,N_14773,N_14410);
nand UO_1148 (O_1148,N_14524,N_14747);
nor UO_1149 (O_1149,N_14856,N_14191);
nand UO_1150 (O_1150,N_14713,N_14935);
and UO_1151 (O_1151,N_14383,N_14652);
and UO_1152 (O_1152,N_14872,N_14160);
and UO_1153 (O_1153,N_14436,N_14606);
and UO_1154 (O_1154,N_14877,N_14213);
or UO_1155 (O_1155,N_14220,N_14129);
or UO_1156 (O_1156,N_14225,N_14907);
or UO_1157 (O_1157,N_14067,N_14617);
xor UO_1158 (O_1158,N_14162,N_14712);
nor UO_1159 (O_1159,N_14860,N_14248);
nor UO_1160 (O_1160,N_14130,N_14491);
nor UO_1161 (O_1161,N_14042,N_14791);
and UO_1162 (O_1162,N_14427,N_14255);
nand UO_1163 (O_1163,N_14348,N_14508);
nor UO_1164 (O_1164,N_14107,N_14325);
nor UO_1165 (O_1165,N_14151,N_14769);
nand UO_1166 (O_1166,N_14776,N_14701);
nor UO_1167 (O_1167,N_14583,N_14402);
or UO_1168 (O_1168,N_14672,N_14647);
nand UO_1169 (O_1169,N_14088,N_14618);
or UO_1170 (O_1170,N_14472,N_14804);
or UO_1171 (O_1171,N_14624,N_14913);
or UO_1172 (O_1172,N_14782,N_14484);
nor UO_1173 (O_1173,N_14986,N_14618);
nor UO_1174 (O_1174,N_14780,N_14809);
and UO_1175 (O_1175,N_14694,N_14509);
or UO_1176 (O_1176,N_14787,N_14975);
or UO_1177 (O_1177,N_14015,N_14189);
nand UO_1178 (O_1178,N_14175,N_14329);
nor UO_1179 (O_1179,N_14420,N_14867);
or UO_1180 (O_1180,N_14856,N_14342);
nor UO_1181 (O_1181,N_14571,N_14676);
or UO_1182 (O_1182,N_14568,N_14323);
or UO_1183 (O_1183,N_14832,N_14589);
or UO_1184 (O_1184,N_14068,N_14319);
nand UO_1185 (O_1185,N_14958,N_14403);
and UO_1186 (O_1186,N_14525,N_14028);
and UO_1187 (O_1187,N_14946,N_14888);
xor UO_1188 (O_1188,N_14888,N_14602);
nand UO_1189 (O_1189,N_14038,N_14783);
nand UO_1190 (O_1190,N_14447,N_14648);
and UO_1191 (O_1191,N_14767,N_14432);
nor UO_1192 (O_1192,N_14807,N_14161);
xnor UO_1193 (O_1193,N_14971,N_14981);
or UO_1194 (O_1194,N_14202,N_14185);
and UO_1195 (O_1195,N_14018,N_14389);
and UO_1196 (O_1196,N_14762,N_14995);
nand UO_1197 (O_1197,N_14552,N_14231);
nand UO_1198 (O_1198,N_14633,N_14851);
or UO_1199 (O_1199,N_14286,N_14936);
or UO_1200 (O_1200,N_14431,N_14933);
nor UO_1201 (O_1201,N_14650,N_14042);
nor UO_1202 (O_1202,N_14040,N_14643);
nor UO_1203 (O_1203,N_14836,N_14185);
or UO_1204 (O_1204,N_14666,N_14046);
and UO_1205 (O_1205,N_14689,N_14275);
and UO_1206 (O_1206,N_14374,N_14938);
or UO_1207 (O_1207,N_14102,N_14484);
or UO_1208 (O_1208,N_14633,N_14588);
nand UO_1209 (O_1209,N_14482,N_14399);
and UO_1210 (O_1210,N_14096,N_14176);
or UO_1211 (O_1211,N_14180,N_14251);
nor UO_1212 (O_1212,N_14169,N_14803);
nor UO_1213 (O_1213,N_14633,N_14867);
nand UO_1214 (O_1214,N_14913,N_14798);
nor UO_1215 (O_1215,N_14968,N_14316);
and UO_1216 (O_1216,N_14354,N_14825);
nor UO_1217 (O_1217,N_14016,N_14391);
nor UO_1218 (O_1218,N_14624,N_14586);
nand UO_1219 (O_1219,N_14081,N_14830);
and UO_1220 (O_1220,N_14502,N_14334);
nor UO_1221 (O_1221,N_14780,N_14048);
and UO_1222 (O_1222,N_14092,N_14003);
and UO_1223 (O_1223,N_14348,N_14197);
or UO_1224 (O_1224,N_14613,N_14123);
or UO_1225 (O_1225,N_14568,N_14130);
nor UO_1226 (O_1226,N_14480,N_14141);
and UO_1227 (O_1227,N_14117,N_14570);
nor UO_1228 (O_1228,N_14095,N_14888);
nor UO_1229 (O_1229,N_14347,N_14891);
and UO_1230 (O_1230,N_14696,N_14227);
nand UO_1231 (O_1231,N_14151,N_14060);
and UO_1232 (O_1232,N_14790,N_14917);
nor UO_1233 (O_1233,N_14518,N_14479);
and UO_1234 (O_1234,N_14661,N_14361);
nand UO_1235 (O_1235,N_14689,N_14414);
nand UO_1236 (O_1236,N_14476,N_14474);
nor UO_1237 (O_1237,N_14111,N_14850);
nor UO_1238 (O_1238,N_14770,N_14769);
nor UO_1239 (O_1239,N_14659,N_14829);
or UO_1240 (O_1240,N_14434,N_14642);
nor UO_1241 (O_1241,N_14720,N_14193);
or UO_1242 (O_1242,N_14060,N_14204);
nand UO_1243 (O_1243,N_14201,N_14594);
nor UO_1244 (O_1244,N_14358,N_14132);
or UO_1245 (O_1245,N_14777,N_14990);
and UO_1246 (O_1246,N_14500,N_14841);
or UO_1247 (O_1247,N_14793,N_14428);
nand UO_1248 (O_1248,N_14549,N_14673);
nand UO_1249 (O_1249,N_14042,N_14123);
nand UO_1250 (O_1250,N_14097,N_14913);
nand UO_1251 (O_1251,N_14599,N_14024);
and UO_1252 (O_1252,N_14739,N_14629);
and UO_1253 (O_1253,N_14625,N_14836);
and UO_1254 (O_1254,N_14370,N_14596);
nor UO_1255 (O_1255,N_14578,N_14354);
or UO_1256 (O_1256,N_14033,N_14551);
nor UO_1257 (O_1257,N_14540,N_14826);
xnor UO_1258 (O_1258,N_14208,N_14593);
nand UO_1259 (O_1259,N_14115,N_14308);
and UO_1260 (O_1260,N_14699,N_14809);
or UO_1261 (O_1261,N_14391,N_14081);
nand UO_1262 (O_1262,N_14466,N_14190);
nor UO_1263 (O_1263,N_14140,N_14680);
nand UO_1264 (O_1264,N_14937,N_14471);
nor UO_1265 (O_1265,N_14408,N_14157);
or UO_1266 (O_1266,N_14284,N_14748);
nor UO_1267 (O_1267,N_14311,N_14401);
nor UO_1268 (O_1268,N_14517,N_14224);
or UO_1269 (O_1269,N_14160,N_14492);
and UO_1270 (O_1270,N_14581,N_14946);
nand UO_1271 (O_1271,N_14870,N_14107);
or UO_1272 (O_1272,N_14321,N_14593);
and UO_1273 (O_1273,N_14158,N_14937);
and UO_1274 (O_1274,N_14366,N_14560);
nor UO_1275 (O_1275,N_14993,N_14858);
nand UO_1276 (O_1276,N_14141,N_14762);
or UO_1277 (O_1277,N_14026,N_14665);
nand UO_1278 (O_1278,N_14250,N_14824);
or UO_1279 (O_1279,N_14189,N_14138);
and UO_1280 (O_1280,N_14902,N_14809);
or UO_1281 (O_1281,N_14285,N_14718);
or UO_1282 (O_1282,N_14323,N_14972);
nor UO_1283 (O_1283,N_14993,N_14576);
nor UO_1284 (O_1284,N_14553,N_14729);
nor UO_1285 (O_1285,N_14639,N_14847);
nor UO_1286 (O_1286,N_14566,N_14812);
and UO_1287 (O_1287,N_14150,N_14256);
and UO_1288 (O_1288,N_14945,N_14450);
nor UO_1289 (O_1289,N_14102,N_14229);
nor UO_1290 (O_1290,N_14368,N_14743);
nand UO_1291 (O_1291,N_14309,N_14372);
nand UO_1292 (O_1292,N_14632,N_14796);
or UO_1293 (O_1293,N_14858,N_14534);
nand UO_1294 (O_1294,N_14339,N_14332);
and UO_1295 (O_1295,N_14664,N_14241);
or UO_1296 (O_1296,N_14704,N_14242);
nand UO_1297 (O_1297,N_14224,N_14569);
nand UO_1298 (O_1298,N_14523,N_14102);
nor UO_1299 (O_1299,N_14793,N_14734);
or UO_1300 (O_1300,N_14130,N_14522);
and UO_1301 (O_1301,N_14614,N_14942);
nor UO_1302 (O_1302,N_14242,N_14787);
or UO_1303 (O_1303,N_14588,N_14263);
nand UO_1304 (O_1304,N_14007,N_14300);
and UO_1305 (O_1305,N_14919,N_14470);
and UO_1306 (O_1306,N_14498,N_14145);
nand UO_1307 (O_1307,N_14269,N_14224);
nand UO_1308 (O_1308,N_14082,N_14832);
or UO_1309 (O_1309,N_14973,N_14013);
nor UO_1310 (O_1310,N_14925,N_14182);
or UO_1311 (O_1311,N_14987,N_14397);
nor UO_1312 (O_1312,N_14281,N_14542);
nor UO_1313 (O_1313,N_14326,N_14702);
nand UO_1314 (O_1314,N_14205,N_14434);
or UO_1315 (O_1315,N_14266,N_14186);
nor UO_1316 (O_1316,N_14928,N_14644);
and UO_1317 (O_1317,N_14099,N_14304);
and UO_1318 (O_1318,N_14272,N_14511);
or UO_1319 (O_1319,N_14662,N_14413);
and UO_1320 (O_1320,N_14397,N_14716);
and UO_1321 (O_1321,N_14651,N_14444);
nor UO_1322 (O_1322,N_14882,N_14701);
nand UO_1323 (O_1323,N_14638,N_14383);
or UO_1324 (O_1324,N_14684,N_14670);
and UO_1325 (O_1325,N_14634,N_14535);
or UO_1326 (O_1326,N_14333,N_14535);
nand UO_1327 (O_1327,N_14572,N_14237);
or UO_1328 (O_1328,N_14621,N_14574);
and UO_1329 (O_1329,N_14528,N_14638);
or UO_1330 (O_1330,N_14548,N_14439);
and UO_1331 (O_1331,N_14603,N_14516);
and UO_1332 (O_1332,N_14541,N_14153);
nand UO_1333 (O_1333,N_14474,N_14517);
or UO_1334 (O_1334,N_14790,N_14309);
nor UO_1335 (O_1335,N_14434,N_14132);
or UO_1336 (O_1336,N_14572,N_14808);
and UO_1337 (O_1337,N_14986,N_14568);
nor UO_1338 (O_1338,N_14811,N_14658);
nand UO_1339 (O_1339,N_14705,N_14157);
nand UO_1340 (O_1340,N_14114,N_14931);
or UO_1341 (O_1341,N_14667,N_14372);
and UO_1342 (O_1342,N_14410,N_14362);
nand UO_1343 (O_1343,N_14537,N_14039);
or UO_1344 (O_1344,N_14092,N_14957);
and UO_1345 (O_1345,N_14991,N_14582);
and UO_1346 (O_1346,N_14869,N_14101);
nor UO_1347 (O_1347,N_14617,N_14569);
xor UO_1348 (O_1348,N_14303,N_14315);
and UO_1349 (O_1349,N_14461,N_14784);
nand UO_1350 (O_1350,N_14762,N_14892);
nand UO_1351 (O_1351,N_14658,N_14074);
and UO_1352 (O_1352,N_14717,N_14622);
nand UO_1353 (O_1353,N_14008,N_14188);
nor UO_1354 (O_1354,N_14740,N_14821);
nand UO_1355 (O_1355,N_14691,N_14930);
nor UO_1356 (O_1356,N_14004,N_14877);
nand UO_1357 (O_1357,N_14396,N_14484);
xor UO_1358 (O_1358,N_14866,N_14384);
nand UO_1359 (O_1359,N_14636,N_14469);
nor UO_1360 (O_1360,N_14953,N_14784);
nand UO_1361 (O_1361,N_14152,N_14948);
nand UO_1362 (O_1362,N_14356,N_14222);
and UO_1363 (O_1363,N_14159,N_14188);
or UO_1364 (O_1364,N_14236,N_14049);
or UO_1365 (O_1365,N_14661,N_14880);
or UO_1366 (O_1366,N_14423,N_14928);
or UO_1367 (O_1367,N_14536,N_14280);
or UO_1368 (O_1368,N_14640,N_14630);
nor UO_1369 (O_1369,N_14717,N_14306);
nand UO_1370 (O_1370,N_14840,N_14118);
nand UO_1371 (O_1371,N_14105,N_14202);
and UO_1372 (O_1372,N_14660,N_14161);
nor UO_1373 (O_1373,N_14491,N_14417);
or UO_1374 (O_1374,N_14364,N_14369);
nand UO_1375 (O_1375,N_14464,N_14178);
nor UO_1376 (O_1376,N_14184,N_14080);
and UO_1377 (O_1377,N_14912,N_14414);
and UO_1378 (O_1378,N_14838,N_14448);
nand UO_1379 (O_1379,N_14836,N_14851);
or UO_1380 (O_1380,N_14276,N_14008);
nor UO_1381 (O_1381,N_14976,N_14688);
nor UO_1382 (O_1382,N_14837,N_14795);
nor UO_1383 (O_1383,N_14718,N_14591);
and UO_1384 (O_1384,N_14857,N_14242);
nand UO_1385 (O_1385,N_14137,N_14771);
nor UO_1386 (O_1386,N_14893,N_14445);
nor UO_1387 (O_1387,N_14191,N_14480);
nor UO_1388 (O_1388,N_14515,N_14870);
or UO_1389 (O_1389,N_14812,N_14689);
nor UO_1390 (O_1390,N_14747,N_14541);
and UO_1391 (O_1391,N_14680,N_14265);
or UO_1392 (O_1392,N_14907,N_14497);
nand UO_1393 (O_1393,N_14999,N_14842);
or UO_1394 (O_1394,N_14336,N_14901);
nor UO_1395 (O_1395,N_14711,N_14060);
nand UO_1396 (O_1396,N_14696,N_14124);
nor UO_1397 (O_1397,N_14952,N_14105);
or UO_1398 (O_1398,N_14223,N_14896);
nor UO_1399 (O_1399,N_14142,N_14682);
and UO_1400 (O_1400,N_14120,N_14159);
nor UO_1401 (O_1401,N_14963,N_14274);
nor UO_1402 (O_1402,N_14721,N_14342);
or UO_1403 (O_1403,N_14165,N_14844);
nor UO_1404 (O_1404,N_14757,N_14408);
nand UO_1405 (O_1405,N_14611,N_14628);
or UO_1406 (O_1406,N_14131,N_14198);
nand UO_1407 (O_1407,N_14519,N_14711);
nor UO_1408 (O_1408,N_14406,N_14177);
nand UO_1409 (O_1409,N_14130,N_14420);
and UO_1410 (O_1410,N_14670,N_14523);
and UO_1411 (O_1411,N_14770,N_14937);
nor UO_1412 (O_1412,N_14322,N_14766);
nor UO_1413 (O_1413,N_14758,N_14290);
or UO_1414 (O_1414,N_14797,N_14844);
or UO_1415 (O_1415,N_14815,N_14347);
and UO_1416 (O_1416,N_14272,N_14163);
or UO_1417 (O_1417,N_14907,N_14877);
nor UO_1418 (O_1418,N_14933,N_14341);
nor UO_1419 (O_1419,N_14915,N_14886);
nor UO_1420 (O_1420,N_14033,N_14916);
and UO_1421 (O_1421,N_14828,N_14945);
and UO_1422 (O_1422,N_14673,N_14667);
or UO_1423 (O_1423,N_14501,N_14013);
nand UO_1424 (O_1424,N_14698,N_14169);
and UO_1425 (O_1425,N_14356,N_14038);
and UO_1426 (O_1426,N_14579,N_14298);
nand UO_1427 (O_1427,N_14465,N_14547);
and UO_1428 (O_1428,N_14763,N_14429);
nor UO_1429 (O_1429,N_14068,N_14086);
nor UO_1430 (O_1430,N_14193,N_14249);
nand UO_1431 (O_1431,N_14093,N_14712);
nor UO_1432 (O_1432,N_14680,N_14965);
or UO_1433 (O_1433,N_14350,N_14501);
and UO_1434 (O_1434,N_14385,N_14882);
or UO_1435 (O_1435,N_14456,N_14776);
and UO_1436 (O_1436,N_14812,N_14692);
nand UO_1437 (O_1437,N_14639,N_14193);
and UO_1438 (O_1438,N_14091,N_14042);
and UO_1439 (O_1439,N_14641,N_14301);
or UO_1440 (O_1440,N_14592,N_14011);
nand UO_1441 (O_1441,N_14261,N_14389);
nand UO_1442 (O_1442,N_14368,N_14222);
nand UO_1443 (O_1443,N_14718,N_14087);
nand UO_1444 (O_1444,N_14568,N_14575);
and UO_1445 (O_1445,N_14059,N_14259);
nor UO_1446 (O_1446,N_14138,N_14689);
and UO_1447 (O_1447,N_14393,N_14246);
and UO_1448 (O_1448,N_14570,N_14034);
nand UO_1449 (O_1449,N_14793,N_14393);
and UO_1450 (O_1450,N_14071,N_14130);
and UO_1451 (O_1451,N_14207,N_14522);
and UO_1452 (O_1452,N_14226,N_14429);
and UO_1453 (O_1453,N_14356,N_14111);
nor UO_1454 (O_1454,N_14138,N_14769);
nor UO_1455 (O_1455,N_14735,N_14014);
and UO_1456 (O_1456,N_14644,N_14141);
nand UO_1457 (O_1457,N_14057,N_14342);
xnor UO_1458 (O_1458,N_14996,N_14097);
nand UO_1459 (O_1459,N_14095,N_14365);
nor UO_1460 (O_1460,N_14563,N_14740);
or UO_1461 (O_1461,N_14370,N_14643);
nor UO_1462 (O_1462,N_14334,N_14545);
nand UO_1463 (O_1463,N_14827,N_14524);
nand UO_1464 (O_1464,N_14450,N_14165);
nor UO_1465 (O_1465,N_14874,N_14106);
or UO_1466 (O_1466,N_14958,N_14718);
nand UO_1467 (O_1467,N_14645,N_14496);
nor UO_1468 (O_1468,N_14792,N_14719);
or UO_1469 (O_1469,N_14868,N_14997);
and UO_1470 (O_1470,N_14186,N_14459);
and UO_1471 (O_1471,N_14735,N_14502);
nor UO_1472 (O_1472,N_14852,N_14366);
nand UO_1473 (O_1473,N_14573,N_14223);
nor UO_1474 (O_1474,N_14359,N_14944);
and UO_1475 (O_1475,N_14754,N_14414);
or UO_1476 (O_1476,N_14589,N_14674);
nand UO_1477 (O_1477,N_14563,N_14870);
nand UO_1478 (O_1478,N_14926,N_14412);
and UO_1479 (O_1479,N_14765,N_14537);
and UO_1480 (O_1480,N_14889,N_14165);
nand UO_1481 (O_1481,N_14753,N_14188);
and UO_1482 (O_1482,N_14092,N_14446);
and UO_1483 (O_1483,N_14160,N_14767);
nor UO_1484 (O_1484,N_14738,N_14058);
or UO_1485 (O_1485,N_14389,N_14928);
or UO_1486 (O_1486,N_14346,N_14485);
and UO_1487 (O_1487,N_14837,N_14510);
or UO_1488 (O_1488,N_14566,N_14464);
nor UO_1489 (O_1489,N_14833,N_14213);
nor UO_1490 (O_1490,N_14751,N_14242);
nand UO_1491 (O_1491,N_14739,N_14000);
or UO_1492 (O_1492,N_14311,N_14091);
and UO_1493 (O_1493,N_14727,N_14769);
and UO_1494 (O_1494,N_14441,N_14350);
nor UO_1495 (O_1495,N_14726,N_14036);
nand UO_1496 (O_1496,N_14379,N_14179);
and UO_1497 (O_1497,N_14852,N_14125);
or UO_1498 (O_1498,N_14836,N_14628);
xnor UO_1499 (O_1499,N_14485,N_14788);
or UO_1500 (O_1500,N_14031,N_14837);
nor UO_1501 (O_1501,N_14802,N_14114);
nor UO_1502 (O_1502,N_14576,N_14569);
nor UO_1503 (O_1503,N_14596,N_14294);
and UO_1504 (O_1504,N_14624,N_14353);
nand UO_1505 (O_1505,N_14470,N_14477);
nor UO_1506 (O_1506,N_14961,N_14636);
or UO_1507 (O_1507,N_14428,N_14470);
nand UO_1508 (O_1508,N_14817,N_14885);
nand UO_1509 (O_1509,N_14265,N_14591);
nor UO_1510 (O_1510,N_14316,N_14077);
nor UO_1511 (O_1511,N_14719,N_14610);
nor UO_1512 (O_1512,N_14216,N_14794);
or UO_1513 (O_1513,N_14827,N_14103);
or UO_1514 (O_1514,N_14139,N_14637);
nor UO_1515 (O_1515,N_14859,N_14655);
nand UO_1516 (O_1516,N_14517,N_14894);
or UO_1517 (O_1517,N_14158,N_14728);
or UO_1518 (O_1518,N_14562,N_14446);
or UO_1519 (O_1519,N_14282,N_14661);
nor UO_1520 (O_1520,N_14939,N_14998);
nor UO_1521 (O_1521,N_14459,N_14630);
nor UO_1522 (O_1522,N_14104,N_14631);
nor UO_1523 (O_1523,N_14508,N_14031);
nor UO_1524 (O_1524,N_14448,N_14579);
nand UO_1525 (O_1525,N_14568,N_14170);
and UO_1526 (O_1526,N_14421,N_14697);
or UO_1527 (O_1527,N_14731,N_14916);
and UO_1528 (O_1528,N_14008,N_14493);
and UO_1529 (O_1529,N_14434,N_14833);
and UO_1530 (O_1530,N_14573,N_14885);
or UO_1531 (O_1531,N_14585,N_14848);
or UO_1532 (O_1532,N_14737,N_14886);
nand UO_1533 (O_1533,N_14857,N_14200);
nand UO_1534 (O_1534,N_14645,N_14955);
nand UO_1535 (O_1535,N_14377,N_14966);
and UO_1536 (O_1536,N_14727,N_14565);
and UO_1537 (O_1537,N_14014,N_14385);
xor UO_1538 (O_1538,N_14268,N_14233);
and UO_1539 (O_1539,N_14948,N_14403);
or UO_1540 (O_1540,N_14237,N_14096);
or UO_1541 (O_1541,N_14137,N_14113);
and UO_1542 (O_1542,N_14942,N_14048);
or UO_1543 (O_1543,N_14393,N_14231);
or UO_1544 (O_1544,N_14366,N_14143);
nor UO_1545 (O_1545,N_14763,N_14641);
or UO_1546 (O_1546,N_14611,N_14975);
nor UO_1547 (O_1547,N_14330,N_14437);
or UO_1548 (O_1548,N_14656,N_14980);
nor UO_1549 (O_1549,N_14855,N_14092);
nand UO_1550 (O_1550,N_14992,N_14394);
nor UO_1551 (O_1551,N_14529,N_14192);
or UO_1552 (O_1552,N_14583,N_14619);
nand UO_1553 (O_1553,N_14097,N_14099);
or UO_1554 (O_1554,N_14203,N_14571);
nand UO_1555 (O_1555,N_14862,N_14542);
or UO_1556 (O_1556,N_14435,N_14108);
or UO_1557 (O_1557,N_14334,N_14656);
and UO_1558 (O_1558,N_14490,N_14357);
or UO_1559 (O_1559,N_14419,N_14462);
nand UO_1560 (O_1560,N_14781,N_14037);
and UO_1561 (O_1561,N_14923,N_14242);
nand UO_1562 (O_1562,N_14989,N_14240);
nand UO_1563 (O_1563,N_14536,N_14528);
nand UO_1564 (O_1564,N_14184,N_14573);
nand UO_1565 (O_1565,N_14148,N_14358);
nor UO_1566 (O_1566,N_14454,N_14007);
nand UO_1567 (O_1567,N_14629,N_14759);
or UO_1568 (O_1568,N_14142,N_14652);
nand UO_1569 (O_1569,N_14007,N_14837);
or UO_1570 (O_1570,N_14733,N_14990);
or UO_1571 (O_1571,N_14590,N_14584);
nor UO_1572 (O_1572,N_14913,N_14725);
nand UO_1573 (O_1573,N_14968,N_14229);
or UO_1574 (O_1574,N_14266,N_14988);
and UO_1575 (O_1575,N_14645,N_14551);
or UO_1576 (O_1576,N_14026,N_14449);
nor UO_1577 (O_1577,N_14746,N_14879);
and UO_1578 (O_1578,N_14930,N_14547);
or UO_1579 (O_1579,N_14867,N_14163);
nor UO_1580 (O_1580,N_14541,N_14005);
nand UO_1581 (O_1581,N_14448,N_14027);
and UO_1582 (O_1582,N_14120,N_14980);
nor UO_1583 (O_1583,N_14111,N_14662);
or UO_1584 (O_1584,N_14803,N_14232);
nor UO_1585 (O_1585,N_14188,N_14285);
or UO_1586 (O_1586,N_14135,N_14847);
nor UO_1587 (O_1587,N_14810,N_14127);
nor UO_1588 (O_1588,N_14193,N_14143);
and UO_1589 (O_1589,N_14704,N_14123);
nand UO_1590 (O_1590,N_14482,N_14230);
nand UO_1591 (O_1591,N_14247,N_14729);
and UO_1592 (O_1592,N_14117,N_14027);
nor UO_1593 (O_1593,N_14313,N_14896);
or UO_1594 (O_1594,N_14860,N_14130);
nor UO_1595 (O_1595,N_14843,N_14808);
nor UO_1596 (O_1596,N_14868,N_14463);
nor UO_1597 (O_1597,N_14937,N_14207);
and UO_1598 (O_1598,N_14300,N_14288);
nor UO_1599 (O_1599,N_14045,N_14867);
or UO_1600 (O_1600,N_14002,N_14940);
or UO_1601 (O_1601,N_14059,N_14633);
or UO_1602 (O_1602,N_14173,N_14402);
nor UO_1603 (O_1603,N_14873,N_14313);
and UO_1604 (O_1604,N_14590,N_14223);
nand UO_1605 (O_1605,N_14848,N_14671);
or UO_1606 (O_1606,N_14309,N_14247);
or UO_1607 (O_1607,N_14097,N_14651);
nor UO_1608 (O_1608,N_14646,N_14638);
nand UO_1609 (O_1609,N_14114,N_14946);
nand UO_1610 (O_1610,N_14383,N_14678);
and UO_1611 (O_1611,N_14652,N_14233);
and UO_1612 (O_1612,N_14132,N_14917);
nand UO_1613 (O_1613,N_14040,N_14750);
or UO_1614 (O_1614,N_14696,N_14971);
and UO_1615 (O_1615,N_14173,N_14739);
or UO_1616 (O_1616,N_14375,N_14634);
nand UO_1617 (O_1617,N_14971,N_14853);
and UO_1618 (O_1618,N_14313,N_14284);
nor UO_1619 (O_1619,N_14988,N_14976);
nor UO_1620 (O_1620,N_14029,N_14887);
or UO_1621 (O_1621,N_14685,N_14009);
or UO_1622 (O_1622,N_14893,N_14430);
nand UO_1623 (O_1623,N_14125,N_14779);
xor UO_1624 (O_1624,N_14117,N_14780);
nand UO_1625 (O_1625,N_14386,N_14721);
or UO_1626 (O_1626,N_14004,N_14030);
nand UO_1627 (O_1627,N_14286,N_14386);
nor UO_1628 (O_1628,N_14903,N_14771);
nor UO_1629 (O_1629,N_14421,N_14647);
nor UO_1630 (O_1630,N_14157,N_14292);
or UO_1631 (O_1631,N_14702,N_14749);
or UO_1632 (O_1632,N_14295,N_14335);
nor UO_1633 (O_1633,N_14743,N_14924);
nor UO_1634 (O_1634,N_14123,N_14044);
and UO_1635 (O_1635,N_14570,N_14913);
nor UO_1636 (O_1636,N_14407,N_14243);
or UO_1637 (O_1637,N_14763,N_14478);
nor UO_1638 (O_1638,N_14649,N_14808);
and UO_1639 (O_1639,N_14545,N_14492);
or UO_1640 (O_1640,N_14996,N_14594);
or UO_1641 (O_1641,N_14059,N_14102);
or UO_1642 (O_1642,N_14244,N_14013);
nor UO_1643 (O_1643,N_14348,N_14798);
nor UO_1644 (O_1644,N_14196,N_14758);
nand UO_1645 (O_1645,N_14807,N_14897);
and UO_1646 (O_1646,N_14328,N_14867);
or UO_1647 (O_1647,N_14791,N_14492);
and UO_1648 (O_1648,N_14663,N_14758);
or UO_1649 (O_1649,N_14796,N_14211);
or UO_1650 (O_1650,N_14149,N_14448);
and UO_1651 (O_1651,N_14828,N_14689);
nand UO_1652 (O_1652,N_14038,N_14106);
or UO_1653 (O_1653,N_14259,N_14870);
or UO_1654 (O_1654,N_14305,N_14877);
nand UO_1655 (O_1655,N_14705,N_14933);
nand UO_1656 (O_1656,N_14299,N_14237);
nand UO_1657 (O_1657,N_14143,N_14546);
or UO_1658 (O_1658,N_14968,N_14081);
nand UO_1659 (O_1659,N_14440,N_14653);
nor UO_1660 (O_1660,N_14325,N_14166);
and UO_1661 (O_1661,N_14268,N_14162);
or UO_1662 (O_1662,N_14412,N_14254);
nand UO_1663 (O_1663,N_14543,N_14628);
nor UO_1664 (O_1664,N_14724,N_14914);
nand UO_1665 (O_1665,N_14406,N_14989);
nand UO_1666 (O_1666,N_14373,N_14896);
nand UO_1667 (O_1667,N_14059,N_14991);
nor UO_1668 (O_1668,N_14680,N_14715);
and UO_1669 (O_1669,N_14048,N_14381);
nor UO_1670 (O_1670,N_14827,N_14621);
nor UO_1671 (O_1671,N_14106,N_14601);
nand UO_1672 (O_1672,N_14731,N_14788);
or UO_1673 (O_1673,N_14484,N_14104);
nand UO_1674 (O_1674,N_14617,N_14494);
nor UO_1675 (O_1675,N_14488,N_14228);
nand UO_1676 (O_1676,N_14063,N_14467);
nand UO_1677 (O_1677,N_14497,N_14927);
nand UO_1678 (O_1678,N_14198,N_14629);
or UO_1679 (O_1679,N_14463,N_14094);
or UO_1680 (O_1680,N_14078,N_14468);
or UO_1681 (O_1681,N_14424,N_14110);
and UO_1682 (O_1682,N_14640,N_14791);
or UO_1683 (O_1683,N_14978,N_14355);
nand UO_1684 (O_1684,N_14465,N_14324);
nor UO_1685 (O_1685,N_14932,N_14442);
nor UO_1686 (O_1686,N_14146,N_14270);
or UO_1687 (O_1687,N_14864,N_14702);
or UO_1688 (O_1688,N_14666,N_14090);
or UO_1689 (O_1689,N_14812,N_14003);
and UO_1690 (O_1690,N_14977,N_14822);
nor UO_1691 (O_1691,N_14858,N_14906);
nor UO_1692 (O_1692,N_14729,N_14769);
and UO_1693 (O_1693,N_14691,N_14581);
and UO_1694 (O_1694,N_14197,N_14858);
or UO_1695 (O_1695,N_14264,N_14045);
and UO_1696 (O_1696,N_14913,N_14482);
and UO_1697 (O_1697,N_14397,N_14274);
nand UO_1698 (O_1698,N_14395,N_14104);
nor UO_1699 (O_1699,N_14142,N_14598);
nand UO_1700 (O_1700,N_14367,N_14021);
or UO_1701 (O_1701,N_14161,N_14579);
nand UO_1702 (O_1702,N_14180,N_14995);
and UO_1703 (O_1703,N_14997,N_14042);
or UO_1704 (O_1704,N_14732,N_14827);
nor UO_1705 (O_1705,N_14951,N_14545);
nor UO_1706 (O_1706,N_14669,N_14774);
and UO_1707 (O_1707,N_14832,N_14663);
nor UO_1708 (O_1708,N_14286,N_14975);
or UO_1709 (O_1709,N_14638,N_14992);
and UO_1710 (O_1710,N_14822,N_14109);
or UO_1711 (O_1711,N_14851,N_14447);
and UO_1712 (O_1712,N_14017,N_14337);
or UO_1713 (O_1713,N_14721,N_14174);
nor UO_1714 (O_1714,N_14864,N_14706);
or UO_1715 (O_1715,N_14909,N_14625);
nor UO_1716 (O_1716,N_14116,N_14362);
nor UO_1717 (O_1717,N_14626,N_14679);
nand UO_1718 (O_1718,N_14539,N_14740);
nand UO_1719 (O_1719,N_14224,N_14740);
or UO_1720 (O_1720,N_14445,N_14805);
nand UO_1721 (O_1721,N_14413,N_14793);
or UO_1722 (O_1722,N_14691,N_14407);
or UO_1723 (O_1723,N_14910,N_14114);
nand UO_1724 (O_1724,N_14916,N_14131);
or UO_1725 (O_1725,N_14648,N_14185);
and UO_1726 (O_1726,N_14232,N_14675);
nand UO_1727 (O_1727,N_14498,N_14056);
nand UO_1728 (O_1728,N_14467,N_14261);
and UO_1729 (O_1729,N_14317,N_14590);
and UO_1730 (O_1730,N_14646,N_14941);
nor UO_1731 (O_1731,N_14333,N_14713);
nor UO_1732 (O_1732,N_14463,N_14036);
and UO_1733 (O_1733,N_14259,N_14842);
or UO_1734 (O_1734,N_14761,N_14125);
nand UO_1735 (O_1735,N_14818,N_14069);
nor UO_1736 (O_1736,N_14354,N_14823);
nand UO_1737 (O_1737,N_14287,N_14380);
nor UO_1738 (O_1738,N_14606,N_14656);
nor UO_1739 (O_1739,N_14450,N_14026);
or UO_1740 (O_1740,N_14513,N_14851);
and UO_1741 (O_1741,N_14094,N_14749);
or UO_1742 (O_1742,N_14140,N_14983);
nand UO_1743 (O_1743,N_14766,N_14498);
nand UO_1744 (O_1744,N_14266,N_14194);
or UO_1745 (O_1745,N_14984,N_14320);
nor UO_1746 (O_1746,N_14393,N_14863);
and UO_1747 (O_1747,N_14562,N_14280);
and UO_1748 (O_1748,N_14432,N_14022);
or UO_1749 (O_1749,N_14619,N_14224);
nand UO_1750 (O_1750,N_14277,N_14474);
nand UO_1751 (O_1751,N_14913,N_14522);
and UO_1752 (O_1752,N_14609,N_14668);
nor UO_1753 (O_1753,N_14037,N_14920);
and UO_1754 (O_1754,N_14580,N_14025);
or UO_1755 (O_1755,N_14436,N_14182);
nand UO_1756 (O_1756,N_14020,N_14098);
or UO_1757 (O_1757,N_14136,N_14474);
or UO_1758 (O_1758,N_14697,N_14263);
nor UO_1759 (O_1759,N_14342,N_14557);
nor UO_1760 (O_1760,N_14793,N_14422);
and UO_1761 (O_1761,N_14138,N_14889);
or UO_1762 (O_1762,N_14423,N_14085);
nand UO_1763 (O_1763,N_14201,N_14651);
nor UO_1764 (O_1764,N_14448,N_14979);
nand UO_1765 (O_1765,N_14298,N_14164);
nor UO_1766 (O_1766,N_14498,N_14433);
or UO_1767 (O_1767,N_14398,N_14136);
nor UO_1768 (O_1768,N_14915,N_14508);
or UO_1769 (O_1769,N_14150,N_14146);
nand UO_1770 (O_1770,N_14079,N_14879);
and UO_1771 (O_1771,N_14924,N_14380);
and UO_1772 (O_1772,N_14906,N_14543);
or UO_1773 (O_1773,N_14652,N_14101);
nor UO_1774 (O_1774,N_14493,N_14486);
or UO_1775 (O_1775,N_14420,N_14088);
nor UO_1776 (O_1776,N_14627,N_14505);
nor UO_1777 (O_1777,N_14330,N_14864);
or UO_1778 (O_1778,N_14703,N_14374);
nor UO_1779 (O_1779,N_14555,N_14956);
or UO_1780 (O_1780,N_14451,N_14838);
or UO_1781 (O_1781,N_14026,N_14560);
and UO_1782 (O_1782,N_14822,N_14798);
nand UO_1783 (O_1783,N_14774,N_14971);
nand UO_1784 (O_1784,N_14475,N_14612);
and UO_1785 (O_1785,N_14000,N_14817);
and UO_1786 (O_1786,N_14552,N_14271);
or UO_1787 (O_1787,N_14871,N_14598);
or UO_1788 (O_1788,N_14557,N_14187);
nand UO_1789 (O_1789,N_14999,N_14832);
nand UO_1790 (O_1790,N_14958,N_14983);
nand UO_1791 (O_1791,N_14594,N_14103);
nand UO_1792 (O_1792,N_14375,N_14731);
or UO_1793 (O_1793,N_14034,N_14876);
or UO_1794 (O_1794,N_14478,N_14875);
and UO_1795 (O_1795,N_14698,N_14107);
nand UO_1796 (O_1796,N_14735,N_14756);
or UO_1797 (O_1797,N_14830,N_14238);
nor UO_1798 (O_1798,N_14726,N_14344);
nand UO_1799 (O_1799,N_14338,N_14301);
nor UO_1800 (O_1800,N_14896,N_14889);
or UO_1801 (O_1801,N_14079,N_14980);
and UO_1802 (O_1802,N_14734,N_14263);
nand UO_1803 (O_1803,N_14505,N_14162);
and UO_1804 (O_1804,N_14249,N_14859);
and UO_1805 (O_1805,N_14850,N_14621);
nor UO_1806 (O_1806,N_14016,N_14182);
nand UO_1807 (O_1807,N_14070,N_14590);
and UO_1808 (O_1808,N_14724,N_14310);
nor UO_1809 (O_1809,N_14240,N_14412);
nand UO_1810 (O_1810,N_14985,N_14543);
nor UO_1811 (O_1811,N_14207,N_14647);
and UO_1812 (O_1812,N_14517,N_14424);
nor UO_1813 (O_1813,N_14556,N_14085);
nor UO_1814 (O_1814,N_14731,N_14886);
and UO_1815 (O_1815,N_14433,N_14255);
nor UO_1816 (O_1816,N_14373,N_14915);
nor UO_1817 (O_1817,N_14866,N_14011);
nand UO_1818 (O_1818,N_14155,N_14066);
nor UO_1819 (O_1819,N_14828,N_14948);
or UO_1820 (O_1820,N_14650,N_14541);
or UO_1821 (O_1821,N_14064,N_14676);
and UO_1822 (O_1822,N_14157,N_14889);
nand UO_1823 (O_1823,N_14189,N_14704);
or UO_1824 (O_1824,N_14993,N_14178);
xnor UO_1825 (O_1825,N_14746,N_14427);
or UO_1826 (O_1826,N_14954,N_14364);
or UO_1827 (O_1827,N_14250,N_14887);
or UO_1828 (O_1828,N_14097,N_14504);
nand UO_1829 (O_1829,N_14227,N_14459);
or UO_1830 (O_1830,N_14884,N_14538);
or UO_1831 (O_1831,N_14024,N_14637);
nor UO_1832 (O_1832,N_14780,N_14439);
nor UO_1833 (O_1833,N_14803,N_14676);
and UO_1834 (O_1834,N_14220,N_14852);
nand UO_1835 (O_1835,N_14139,N_14697);
and UO_1836 (O_1836,N_14669,N_14684);
and UO_1837 (O_1837,N_14894,N_14814);
nand UO_1838 (O_1838,N_14351,N_14171);
nor UO_1839 (O_1839,N_14477,N_14957);
nor UO_1840 (O_1840,N_14184,N_14472);
nor UO_1841 (O_1841,N_14131,N_14982);
nor UO_1842 (O_1842,N_14601,N_14440);
nor UO_1843 (O_1843,N_14241,N_14440);
and UO_1844 (O_1844,N_14125,N_14048);
nand UO_1845 (O_1845,N_14122,N_14611);
and UO_1846 (O_1846,N_14023,N_14506);
or UO_1847 (O_1847,N_14051,N_14721);
and UO_1848 (O_1848,N_14635,N_14319);
nand UO_1849 (O_1849,N_14348,N_14051);
xor UO_1850 (O_1850,N_14406,N_14456);
nand UO_1851 (O_1851,N_14613,N_14262);
nor UO_1852 (O_1852,N_14537,N_14565);
nor UO_1853 (O_1853,N_14263,N_14165);
and UO_1854 (O_1854,N_14807,N_14623);
nand UO_1855 (O_1855,N_14309,N_14515);
or UO_1856 (O_1856,N_14732,N_14238);
or UO_1857 (O_1857,N_14164,N_14723);
nand UO_1858 (O_1858,N_14771,N_14675);
nand UO_1859 (O_1859,N_14237,N_14164);
nor UO_1860 (O_1860,N_14908,N_14728);
nand UO_1861 (O_1861,N_14120,N_14042);
or UO_1862 (O_1862,N_14285,N_14511);
nor UO_1863 (O_1863,N_14083,N_14173);
nand UO_1864 (O_1864,N_14349,N_14198);
or UO_1865 (O_1865,N_14018,N_14289);
or UO_1866 (O_1866,N_14372,N_14085);
or UO_1867 (O_1867,N_14584,N_14786);
nand UO_1868 (O_1868,N_14438,N_14003);
and UO_1869 (O_1869,N_14602,N_14348);
nor UO_1870 (O_1870,N_14534,N_14748);
nand UO_1871 (O_1871,N_14341,N_14463);
nand UO_1872 (O_1872,N_14345,N_14850);
or UO_1873 (O_1873,N_14747,N_14391);
nand UO_1874 (O_1874,N_14477,N_14616);
nand UO_1875 (O_1875,N_14798,N_14364);
nor UO_1876 (O_1876,N_14297,N_14910);
or UO_1877 (O_1877,N_14926,N_14332);
nor UO_1878 (O_1878,N_14807,N_14044);
and UO_1879 (O_1879,N_14925,N_14875);
nor UO_1880 (O_1880,N_14848,N_14120);
nor UO_1881 (O_1881,N_14357,N_14498);
and UO_1882 (O_1882,N_14037,N_14285);
or UO_1883 (O_1883,N_14513,N_14658);
nand UO_1884 (O_1884,N_14396,N_14352);
nand UO_1885 (O_1885,N_14091,N_14056);
or UO_1886 (O_1886,N_14154,N_14262);
and UO_1887 (O_1887,N_14705,N_14168);
nand UO_1888 (O_1888,N_14328,N_14368);
and UO_1889 (O_1889,N_14695,N_14197);
and UO_1890 (O_1890,N_14636,N_14894);
or UO_1891 (O_1891,N_14283,N_14044);
nand UO_1892 (O_1892,N_14921,N_14482);
nor UO_1893 (O_1893,N_14809,N_14461);
or UO_1894 (O_1894,N_14823,N_14347);
and UO_1895 (O_1895,N_14404,N_14027);
nand UO_1896 (O_1896,N_14067,N_14603);
and UO_1897 (O_1897,N_14798,N_14421);
and UO_1898 (O_1898,N_14257,N_14328);
or UO_1899 (O_1899,N_14151,N_14221);
or UO_1900 (O_1900,N_14723,N_14315);
nor UO_1901 (O_1901,N_14147,N_14774);
or UO_1902 (O_1902,N_14172,N_14961);
nor UO_1903 (O_1903,N_14576,N_14603);
nand UO_1904 (O_1904,N_14292,N_14988);
and UO_1905 (O_1905,N_14665,N_14114);
nor UO_1906 (O_1906,N_14182,N_14518);
and UO_1907 (O_1907,N_14487,N_14661);
nor UO_1908 (O_1908,N_14666,N_14320);
or UO_1909 (O_1909,N_14795,N_14836);
and UO_1910 (O_1910,N_14831,N_14910);
and UO_1911 (O_1911,N_14117,N_14368);
and UO_1912 (O_1912,N_14334,N_14386);
nor UO_1913 (O_1913,N_14281,N_14244);
nand UO_1914 (O_1914,N_14123,N_14461);
and UO_1915 (O_1915,N_14359,N_14207);
or UO_1916 (O_1916,N_14438,N_14694);
nand UO_1917 (O_1917,N_14672,N_14090);
nor UO_1918 (O_1918,N_14070,N_14808);
and UO_1919 (O_1919,N_14511,N_14602);
and UO_1920 (O_1920,N_14186,N_14602);
and UO_1921 (O_1921,N_14728,N_14740);
nand UO_1922 (O_1922,N_14130,N_14652);
and UO_1923 (O_1923,N_14676,N_14663);
nand UO_1924 (O_1924,N_14719,N_14196);
nand UO_1925 (O_1925,N_14306,N_14984);
or UO_1926 (O_1926,N_14717,N_14905);
nand UO_1927 (O_1927,N_14124,N_14769);
and UO_1928 (O_1928,N_14853,N_14476);
nor UO_1929 (O_1929,N_14992,N_14667);
or UO_1930 (O_1930,N_14506,N_14525);
nor UO_1931 (O_1931,N_14112,N_14697);
or UO_1932 (O_1932,N_14017,N_14838);
and UO_1933 (O_1933,N_14844,N_14026);
nor UO_1934 (O_1934,N_14882,N_14343);
nand UO_1935 (O_1935,N_14208,N_14682);
and UO_1936 (O_1936,N_14773,N_14137);
or UO_1937 (O_1937,N_14576,N_14744);
nand UO_1938 (O_1938,N_14446,N_14148);
nor UO_1939 (O_1939,N_14977,N_14388);
and UO_1940 (O_1940,N_14408,N_14728);
nand UO_1941 (O_1941,N_14617,N_14409);
and UO_1942 (O_1942,N_14821,N_14655);
nand UO_1943 (O_1943,N_14650,N_14957);
nand UO_1944 (O_1944,N_14049,N_14252);
nand UO_1945 (O_1945,N_14960,N_14700);
and UO_1946 (O_1946,N_14497,N_14594);
nand UO_1947 (O_1947,N_14524,N_14242);
or UO_1948 (O_1948,N_14856,N_14173);
nand UO_1949 (O_1949,N_14542,N_14716);
and UO_1950 (O_1950,N_14528,N_14863);
and UO_1951 (O_1951,N_14740,N_14930);
nand UO_1952 (O_1952,N_14702,N_14003);
or UO_1953 (O_1953,N_14196,N_14048);
and UO_1954 (O_1954,N_14079,N_14420);
xnor UO_1955 (O_1955,N_14490,N_14226);
nor UO_1956 (O_1956,N_14619,N_14044);
nand UO_1957 (O_1957,N_14962,N_14678);
and UO_1958 (O_1958,N_14289,N_14356);
nand UO_1959 (O_1959,N_14563,N_14081);
and UO_1960 (O_1960,N_14360,N_14258);
and UO_1961 (O_1961,N_14656,N_14522);
and UO_1962 (O_1962,N_14085,N_14268);
or UO_1963 (O_1963,N_14599,N_14288);
or UO_1964 (O_1964,N_14184,N_14952);
and UO_1965 (O_1965,N_14121,N_14798);
and UO_1966 (O_1966,N_14333,N_14586);
nor UO_1967 (O_1967,N_14615,N_14292);
or UO_1968 (O_1968,N_14534,N_14520);
nand UO_1969 (O_1969,N_14600,N_14158);
nand UO_1970 (O_1970,N_14223,N_14020);
nor UO_1971 (O_1971,N_14962,N_14324);
or UO_1972 (O_1972,N_14509,N_14344);
nand UO_1973 (O_1973,N_14175,N_14915);
or UO_1974 (O_1974,N_14435,N_14338);
or UO_1975 (O_1975,N_14087,N_14378);
nand UO_1976 (O_1976,N_14424,N_14079);
and UO_1977 (O_1977,N_14815,N_14745);
or UO_1978 (O_1978,N_14002,N_14927);
nand UO_1979 (O_1979,N_14133,N_14245);
nor UO_1980 (O_1980,N_14891,N_14027);
and UO_1981 (O_1981,N_14393,N_14963);
and UO_1982 (O_1982,N_14567,N_14176);
and UO_1983 (O_1983,N_14206,N_14468);
or UO_1984 (O_1984,N_14564,N_14500);
nand UO_1985 (O_1985,N_14009,N_14370);
nand UO_1986 (O_1986,N_14432,N_14974);
or UO_1987 (O_1987,N_14365,N_14724);
and UO_1988 (O_1988,N_14217,N_14222);
and UO_1989 (O_1989,N_14797,N_14342);
nor UO_1990 (O_1990,N_14779,N_14784);
and UO_1991 (O_1991,N_14836,N_14968);
nand UO_1992 (O_1992,N_14839,N_14105);
and UO_1993 (O_1993,N_14080,N_14138);
and UO_1994 (O_1994,N_14422,N_14176);
or UO_1995 (O_1995,N_14641,N_14430);
and UO_1996 (O_1996,N_14965,N_14999);
or UO_1997 (O_1997,N_14578,N_14360);
and UO_1998 (O_1998,N_14322,N_14889);
nand UO_1999 (O_1999,N_14122,N_14308);
endmodule