module basic_1000_10000_1500_100_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_153,In_34);
nor U1 (N_1,In_44,In_429);
and U2 (N_2,In_347,In_128);
and U3 (N_3,In_868,In_398);
nor U4 (N_4,In_302,In_395);
or U5 (N_5,In_26,In_134);
or U6 (N_6,In_824,In_122);
nor U7 (N_7,In_378,In_68);
nand U8 (N_8,In_893,In_256);
xnor U9 (N_9,In_486,In_394);
nand U10 (N_10,In_215,In_979);
and U11 (N_11,In_106,In_17);
or U12 (N_12,In_258,In_612);
or U13 (N_13,In_235,In_572);
nor U14 (N_14,In_994,In_896);
or U15 (N_15,In_36,In_875);
or U16 (N_16,In_148,In_200);
or U17 (N_17,In_100,In_748);
and U18 (N_18,In_700,In_178);
nand U19 (N_19,In_877,In_188);
and U20 (N_20,In_871,In_244);
or U21 (N_21,In_112,In_287);
nor U22 (N_22,In_158,In_445);
and U23 (N_23,In_733,In_467);
nand U24 (N_24,In_724,In_262);
nand U25 (N_25,In_130,In_655);
nand U26 (N_26,In_409,In_300);
nand U27 (N_27,In_358,In_731);
nand U28 (N_28,In_276,In_676);
and U29 (N_29,In_630,In_681);
nor U30 (N_30,In_752,In_649);
nor U31 (N_31,In_997,In_760);
and U32 (N_32,In_527,In_853);
nand U33 (N_33,In_746,In_356);
xor U34 (N_34,In_801,In_671);
xor U35 (N_35,In_229,In_74);
or U36 (N_36,In_620,In_545);
nor U37 (N_37,In_856,In_468);
or U38 (N_38,In_702,In_920);
or U39 (N_39,In_46,In_913);
nand U40 (N_40,In_621,In_541);
or U41 (N_41,In_114,In_761);
and U42 (N_42,In_903,In_911);
and U43 (N_43,In_393,In_196);
and U44 (N_44,In_172,In_9);
or U45 (N_45,In_659,In_249);
nand U46 (N_46,In_870,In_758);
and U47 (N_47,In_860,In_452);
nor U48 (N_48,In_810,In_607);
and U49 (N_49,In_532,In_206);
nand U50 (N_50,In_633,In_842);
or U51 (N_51,In_806,In_846);
nand U52 (N_52,In_907,In_594);
and U53 (N_53,In_127,In_462);
nand U54 (N_54,In_73,In_214);
nand U55 (N_55,In_382,In_794);
and U56 (N_56,In_16,In_283);
and U57 (N_57,In_683,In_170);
nor U58 (N_58,In_32,In_892);
and U59 (N_59,In_21,In_253);
or U60 (N_60,In_267,In_368);
nor U61 (N_61,In_147,In_493);
nand U62 (N_62,In_165,In_551);
and U63 (N_63,In_471,In_980);
nand U64 (N_64,In_342,In_270);
nor U65 (N_65,In_446,In_812);
nor U66 (N_66,In_474,In_776);
and U67 (N_67,In_27,In_414);
nand U68 (N_68,In_960,In_243);
nand U69 (N_69,In_54,In_273);
and U70 (N_70,In_970,In_232);
xnor U71 (N_71,In_661,In_764);
nor U72 (N_72,In_438,In_146);
nand U73 (N_73,In_506,In_841);
and U74 (N_74,In_963,In_567);
nor U75 (N_75,In_706,In_247);
or U76 (N_76,In_484,In_201);
nand U77 (N_77,In_837,In_682);
and U78 (N_78,In_540,In_339);
or U79 (N_79,In_408,In_640);
and U80 (N_80,In_882,In_183);
nand U81 (N_81,In_729,In_777);
and U82 (N_82,In_495,In_538);
nand U83 (N_83,In_585,In_522);
nand U84 (N_84,In_605,In_12);
nor U85 (N_85,In_624,In_2);
nand U86 (N_86,In_207,In_922);
and U87 (N_87,In_660,In_935);
or U88 (N_88,In_285,In_718);
nor U89 (N_89,In_677,In_167);
nand U90 (N_90,In_785,In_190);
nor U91 (N_91,In_263,In_505);
or U92 (N_92,In_863,In_861);
or U93 (N_93,In_105,In_432);
or U94 (N_94,In_361,In_182);
nand U95 (N_95,In_370,In_513);
and U96 (N_96,In_738,In_813);
or U97 (N_97,In_116,In_915);
or U98 (N_98,In_646,In_376);
and U99 (N_99,In_547,In_756);
and U100 (N_100,In_530,In_266);
nor U101 (N_101,N_59,In_749);
nor U102 (N_102,In_526,N_33);
nand U103 (N_103,In_701,In_279);
and U104 (N_104,In_595,N_48);
and U105 (N_105,In_515,In_982);
nand U106 (N_106,In_889,N_99);
or U107 (N_107,In_898,In_946);
and U108 (N_108,In_7,In_866);
nand U109 (N_109,In_928,In_163);
and U110 (N_110,N_31,In_216);
and U111 (N_111,In_265,In_783);
or U112 (N_112,In_237,In_419);
or U113 (N_113,N_15,In_867);
nand U114 (N_114,In_511,In_154);
nor U115 (N_115,In_840,In_968);
nor U116 (N_116,In_628,In_383);
nand U117 (N_117,In_140,In_24);
and U118 (N_118,N_69,In_930);
nand U119 (N_119,In_528,In_684);
or U120 (N_120,N_41,In_110);
nand U121 (N_121,In_591,In_502);
nand U122 (N_122,In_145,In_869);
and U123 (N_123,In_821,N_62);
nand U124 (N_124,In_972,In_827);
xnor U125 (N_125,In_331,N_5);
nor U126 (N_126,In_184,In_876);
or U127 (N_127,In_992,In_55);
and U128 (N_128,In_734,In_976);
nand U129 (N_129,In_726,In_135);
nand U130 (N_130,In_407,In_973);
nor U131 (N_131,In_675,In_236);
nor U132 (N_132,In_665,In_619);
or U133 (N_133,In_834,In_63);
nor U134 (N_134,In_259,In_354);
nand U135 (N_135,In_989,In_208);
or U136 (N_136,In_228,In_90);
nor U137 (N_137,In_571,In_195);
nor U138 (N_138,In_353,In_645);
or U139 (N_139,N_54,In_97);
and U140 (N_140,In_780,In_956);
nor U141 (N_141,In_379,In_223);
and U142 (N_142,N_42,In_891);
nand U143 (N_143,In_974,In_103);
nand U144 (N_144,In_473,In_601);
nor U145 (N_145,In_616,In_217);
or U146 (N_146,In_78,In_838);
nand U147 (N_147,In_220,In_131);
nand U148 (N_148,N_97,In_549);
and U149 (N_149,In_653,In_565);
or U150 (N_150,In_156,In_322);
or U151 (N_151,In_152,In_290);
and U152 (N_152,In_350,In_83);
nor U153 (N_153,In_80,In_5);
and U154 (N_154,In_67,In_967);
or U155 (N_155,In_179,In_8);
nor U156 (N_156,In_852,In_168);
nand U157 (N_157,In_656,N_50);
or U158 (N_158,In_521,In_995);
or U159 (N_159,In_346,In_294);
nand U160 (N_160,In_865,In_969);
nor U161 (N_161,In_977,N_7);
nor U162 (N_162,In_472,In_280);
nand U163 (N_163,In_475,N_10);
nand U164 (N_164,In_494,In_643);
nor U165 (N_165,In_47,In_335);
and U166 (N_166,In_464,N_44);
and U167 (N_167,In_599,N_27);
and U168 (N_168,In_574,In_849);
nor U169 (N_169,In_906,In_209);
nor U170 (N_170,In_577,In_711);
nor U171 (N_171,In_49,In_470);
and U172 (N_172,In_453,In_524);
nor U173 (N_173,In_912,In_603);
and U174 (N_174,N_34,In_76);
and U175 (N_175,In_788,In_424);
and U176 (N_176,In_899,In_441);
nor U177 (N_177,N_25,N_11);
nand U178 (N_178,In_772,N_46);
and U179 (N_179,In_321,In_552);
nor U180 (N_180,In_298,In_81);
xnor U181 (N_181,In_299,In_205);
nor U182 (N_182,In_864,In_3);
or U183 (N_183,In_781,N_70);
nor U184 (N_184,In_908,In_962);
or U185 (N_185,In_385,In_98);
and U186 (N_186,In_798,In_480);
or U187 (N_187,In_371,In_485);
nand U188 (N_188,In_874,In_62);
nor U189 (N_189,In_808,N_36);
nor U190 (N_190,In_917,N_29);
and U191 (N_191,In_845,In_844);
nand U192 (N_192,In_560,In_15);
nor U193 (N_193,In_826,In_957);
nor U194 (N_194,In_695,In_28);
nand U195 (N_195,In_86,In_554);
nand U196 (N_196,In_461,In_449);
nor U197 (N_197,In_625,In_598);
xor U198 (N_198,In_314,In_92);
nor U199 (N_199,In_602,In_910);
nand U200 (N_200,N_100,In_850);
or U201 (N_201,In_550,In_650);
and U202 (N_202,In_859,N_135);
nand U203 (N_203,N_45,In_365);
nand U204 (N_204,N_167,In_955);
and U205 (N_205,In_242,N_172);
nor U206 (N_206,N_109,In_292);
nor U207 (N_207,In_58,In_37);
and U208 (N_208,In_180,In_213);
or U209 (N_209,In_117,In_779);
nand U210 (N_210,In_126,In_241);
nor U211 (N_211,In_890,N_52);
or U212 (N_212,In_366,In_425);
and U213 (N_213,In_218,In_454);
and U214 (N_214,In_586,In_138);
nand U215 (N_215,In_512,In_789);
nor U216 (N_216,N_186,In_857);
nand U217 (N_217,In_402,In_987);
nor U218 (N_218,In_582,N_168);
or U219 (N_219,In_820,In_436);
or U220 (N_220,In_93,In_669);
nor U221 (N_221,In_23,In_904);
nor U222 (N_222,N_177,In_288);
nand U223 (N_223,In_631,In_887);
nor U224 (N_224,In_389,In_923);
nand U225 (N_225,In_48,In_177);
or U226 (N_226,N_142,In_744);
nand U227 (N_227,In_119,In_89);
nor U228 (N_228,In_52,In_261);
and U229 (N_229,In_38,In_570);
nor U230 (N_230,In_412,In_1);
and U231 (N_231,In_689,In_947);
nand U232 (N_232,In_670,In_685);
nand U233 (N_233,In_697,N_14);
nand U234 (N_234,In_568,N_180);
nand U235 (N_235,N_107,In_939);
nand U236 (N_236,In_858,In_714);
or U237 (N_237,In_730,N_106);
and U238 (N_238,In_759,In_301);
nand U239 (N_239,In_715,In_442);
nand U240 (N_240,In_699,In_186);
or U241 (N_241,In_828,In_316);
nand U242 (N_242,In_872,In_193);
or U243 (N_243,In_264,N_90);
and U244 (N_244,In_953,In_501);
and U245 (N_245,In_588,In_274);
and U246 (N_246,N_163,In_404);
nor U247 (N_247,In_771,In_897);
and U248 (N_248,In_708,In_648);
and U249 (N_249,In_476,In_144);
and U250 (N_250,In_481,In_377);
and U251 (N_251,In_597,In_459);
or U252 (N_252,N_196,N_83);
nand U253 (N_253,In_765,In_774);
and U254 (N_254,In_735,In_931);
and U255 (N_255,N_193,In_831);
nor U256 (N_256,In_691,N_86);
nor U257 (N_257,N_102,In_988);
nand U258 (N_258,In_364,In_30);
or U259 (N_259,In_750,In_797);
or U260 (N_260,N_8,In_51);
nand U261 (N_261,In_338,In_84);
or U262 (N_262,In_428,In_340);
or U263 (N_263,N_132,N_184);
or U264 (N_264,In_707,In_33);
nor U265 (N_265,In_916,N_188);
or U266 (N_266,In_664,In_465);
nor U267 (N_267,In_349,In_673);
xnor U268 (N_268,In_139,In_975);
nor U269 (N_269,In_647,N_56);
or U270 (N_270,N_28,In_355);
or U271 (N_271,In_203,In_964);
nand U272 (N_272,In_434,In_958);
or U273 (N_273,In_590,N_155);
nand U274 (N_274,In_741,N_190);
nand U275 (N_275,N_47,In_825);
nor U276 (N_276,In_490,In_492);
xnor U277 (N_277,In_72,In_202);
nor U278 (N_278,In_723,In_230);
nor U279 (N_279,N_63,In_142);
or U280 (N_280,In_945,In_634);
xnor U281 (N_281,In_418,In_489);
or U282 (N_282,In_53,In_751);
and U283 (N_283,In_199,In_885);
nor U284 (N_284,In_456,N_182);
and U285 (N_285,In_403,In_770);
nand U286 (N_286,N_195,N_127);
or U287 (N_287,In_141,In_272);
nand U288 (N_288,In_416,N_73);
or U289 (N_289,In_610,In_985);
nand U290 (N_290,N_152,In_909);
and U291 (N_291,N_37,In_657);
and U292 (N_292,N_118,N_141);
nor U293 (N_293,In_900,In_719);
nor U294 (N_294,In_327,N_112);
and U295 (N_295,N_148,In_629);
and U296 (N_296,In_29,In_600);
nand U297 (N_297,N_115,In_96);
nand U298 (N_298,In_477,In_564);
and U299 (N_299,In_488,In_627);
or U300 (N_300,N_61,In_795);
and U301 (N_301,In_224,In_818);
nor U302 (N_302,In_233,In_329);
nor U303 (N_303,N_225,In_936);
or U304 (N_304,In_757,In_658);
nand U305 (N_305,In_31,In_952);
and U306 (N_306,In_85,In_359);
or U307 (N_307,In_546,In_71);
nand U308 (N_308,N_64,In_666);
or U309 (N_309,In_766,In_155);
nand U310 (N_310,In_422,In_822);
or U311 (N_311,In_529,In_192);
nor U312 (N_312,In_637,N_80);
nand U313 (N_313,N_299,In_296);
or U314 (N_314,N_24,In_293);
nor U315 (N_315,In_523,N_176);
and U316 (N_316,In_563,In_622);
nand U317 (N_317,In_252,In_390);
nor U318 (N_318,N_35,N_91);
or U319 (N_319,In_555,In_809);
nand U320 (N_320,In_176,N_20);
nand U321 (N_321,In_251,N_194);
or U322 (N_322,In_914,In_792);
nand U323 (N_323,In_227,N_290);
nor U324 (N_324,In_282,In_159);
nand U325 (N_325,N_26,In_57);
nand U326 (N_326,In_929,In_149);
or U327 (N_327,In_815,N_187);
and U328 (N_328,N_104,N_265);
and U329 (N_329,N_160,In_709);
nand U330 (N_330,In_693,N_147);
and U331 (N_331,In_499,In_884);
and U332 (N_332,In_234,In_615);
or U333 (N_333,In_954,In_517);
or U334 (N_334,In_636,In_663);
nand U335 (N_335,In_632,In_392);
or U336 (N_336,In_687,In_450);
and U337 (N_337,N_292,In_843);
or U338 (N_338,In_642,In_753);
nor U339 (N_339,N_241,N_58);
or U340 (N_340,N_261,N_159);
or U341 (N_341,In_345,In_690);
nand U342 (N_342,N_143,N_0);
or U343 (N_343,In_539,In_310);
and U344 (N_344,In_79,In_173);
nand U345 (N_345,In_773,In_966);
nand U346 (N_346,N_126,In_41);
nand U347 (N_347,In_129,In_886);
or U348 (N_348,N_81,N_215);
nand U349 (N_349,N_236,N_111);
or U350 (N_350,In_397,In_959);
or U351 (N_351,In_983,In_308);
and U352 (N_352,In_786,N_283);
or U353 (N_353,N_79,In_204);
and U354 (N_354,In_938,In_592);
or U355 (N_355,In_520,N_206);
or U356 (N_356,In_623,N_23);
or U357 (N_357,In_851,In_854);
or U358 (N_358,In_796,In_91);
nor U359 (N_359,In_70,In_504);
nor U360 (N_360,N_157,N_150);
or U361 (N_361,In_950,In_304);
nand U362 (N_362,In_118,N_271);
nand U363 (N_363,In_307,In_277);
and U364 (N_364,In_94,In_271);
and U365 (N_365,In_123,N_101);
xor U366 (N_366,In_804,N_138);
nor U367 (N_367,N_60,In_423);
and U368 (N_368,In_755,N_134);
or U369 (N_369,In_18,In_162);
nand U370 (N_370,N_228,In_325);
and U371 (N_371,In_544,In_121);
nor U372 (N_372,In_341,In_313);
or U373 (N_373,In_374,In_732);
nor U374 (N_374,In_557,N_130);
or U375 (N_375,N_113,In_561);
nor U376 (N_376,In_924,In_618);
nand U377 (N_377,In_548,N_203);
nand U378 (N_378,N_255,In_426);
nor U379 (N_379,N_237,N_131);
nor U380 (N_380,In_437,In_401);
xnor U381 (N_381,N_22,In_754);
nand U382 (N_382,In_575,N_139);
nand U383 (N_383,N_239,In_999);
nand U384 (N_384,N_169,In_536);
and U385 (N_385,In_500,N_231);
nor U386 (N_386,In_981,N_178);
nor U387 (N_387,N_129,In_367);
nand U388 (N_388,In_136,In_133);
nand U389 (N_389,In_894,N_192);
nor U390 (N_390,N_173,In_769);
nand U391 (N_391,In_878,In_312);
or U392 (N_392,N_214,In_246);
or U393 (N_393,In_879,In_343);
nand U394 (N_394,In_596,In_143);
and U395 (N_395,N_213,In_921);
and U396 (N_396,N_85,In_888);
nor U397 (N_397,N_119,In_873);
or U398 (N_398,In_406,N_296);
or U399 (N_399,N_71,In_435);
or U400 (N_400,In_311,In_836);
nand U401 (N_401,N_258,In_496);
nor U402 (N_402,In_583,N_137);
and U403 (N_403,N_189,In_881);
nand U404 (N_404,In_614,In_559);
nand U405 (N_405,In_439,In_745);
nand U406 (N_406,N_229,In_805);
nand U407 (N_407,N_222,N_234);
nor U408 (N_408,N_396,In_819);
nor U409 (N_409,In_175,In_45);
nor U410 (N_410,N_13,N_313);
or U411 (N_411,N_276,In_351);
and U412 (N_412,N_165,In_151);
nor U413 (N_413,N_57,N_95);
xnor U414 (N_414,N_337,In_319);
or U415 (N_415,In_169,N_96);
or U416 (N_416,In_286,In_42);
nor U417 (N_417,N_377,In_722);
or U418 (N_418,In_862,In_430);
nand U419 (N_419,In_132,N_343);
xnor U420 (N_420,N_67,In_531);
nand U421 (N_421,In_25,In_638);
nand U422 (N_422,In_231,N_383);
or U423 (N_423,N_375,In_833);
nor U424 (N_424,N_347,In_832);
nor U425 (N_425,In_823,N_397);
nand U426 (N_426,N_392,N_94);
nor U427 (N_427,In_226,N_154);
nand U428 (N_428,N_39,N_220);
nor U429 (N_429,In_166,In_775);
nor U430 (N_430,N_367,In_703);
nand U431 (N_431,N_361,In_417);
and U432 (N_432,In_275,N_318);
xor U433 (N_433,In_509,N_352);
and U434 (N_434,In_626,In_543);
nand U435 (N_435,N_286,N_3);
nand U436 (N_436,N_125,In_839);
or U437 (N_437,In_194,In_728);
or U438 (N_438,N_368,In_56);
nand U439 (N_439,N_72,In_82);
and U440 (N_440,In_662,In_934);
nor U441 (N_441,N_294,N_212);
or U442 (N_442,N_279,N_218);
nand U443 (N_443,In_463,N_242);
or U444 (N_444,In_458,In_932);
and U445 (N_445,In_317,In_508);
or U446 (N_446,N_371,In_360);
xor U447 (N_447,N_278,N_300);
and U448 (N_448,N_317,In_609);
nor U449 (N_449,In_793,In_902);
nor U450 (N_450,N_205,In_533);
nor U451 (N_451,N_207,In_778);
nor U452 (N_452,In_219,In_405);
nor U453 (N_453,In_667,In_381);
or U454 (N_454,N_308,In_400);
or U455 (N_455,N_19,N_145);
and U456 (N_456,N_251,In_587);
nor U457 (N_457,N_274,N_327);
or U458 (N_458,In_427,N_391);
xor U459 (N_459,N_248,N_223);
nand U460 (N_460,N_179,In_455);
or U461 (N_461,In_357,In_883);
nor U462 (N_462,In_60,In_978);
or U463 (N_463,N_211,In_372);
nor U464 (N_464,N_105,N_68);
nand U465 (N_465,In_800,In_767);
nand U466 (N_466,In_210,In_161);
or U467 (N_467,N_314,In_584);
and U468 (N_468,In_942,In_951);
or U469 (N_469,In_120,N_121);
or U470 (N_470,N_144,In_245);
or U471 (N_471,N_307,In_895);
and U472 (N_472,N_362,In_14);
nand U473 (N_473,N_66,In_516);
nand U474 (N_474,In_10,In_413);
or U475 (N_475,N_110,In_535);
or U476 (N_476,In_613,N_297);
nor U477 (N_477,N_330,N_390);
nor U478 (N_478,In_569,N_197);
or U479 (N_479,N_263,In_686);
nand U480 (N_480,In_692,In_940);
and U481 (N_481,N_301,In_807);
nor U482 (N_482,In_925,N_381);
nor U483 (N_483,In_905,N_285);
and U484 (N_484,N_346,N_288);
nand U485 (N_485,N_219,N_341);
nor U486 (N_486,In_802,N_333);
nor U487 (N_487,In_410,N_191);
nor U488 (N_488,N_360,In_104);
and U489 (N_489,N_84,In_380);
or U490 (N_490,N_270,In_606);
nor U491 (N_491,In_716,In_421);
and U492 (N_492,In_652,In_69);
or U493 (N_493,In_212,In_420);
and U494 (N_494,N_287,N_289);
nor U495 (N_495,In_101,In_99);
nor U496 (N_496,N_365,In_944);
and U497 (N_497,In_109,N_124);
nor U498 (N_498,In_580,N_51);
and U499 (N_499,N_356,N_16);
nand U500 (N_500,In_39,N_476);
nand U501 (N_501,N_415,In_113);
nor U502 (N_502,In_717,N_321);
nand U503 (N_503,N_284,N_484);
nor U504 (N_504,N_411,N_114);
nand U505 (N_505,N_473,In_77);
nor U506 (N_506,N_407,In_933);
nor U507 (N_507,In_451,N_266);
nand U508 (N_508,In_19,In_269);
nor U509 (N_509,N_442,N_158);
or U510 (N_510,N_403,In_289);
nand U511 (N_511,N_456,In_617);
nand U512 (N_512,N_434,N_183);
nor U513 (N_513,N_432,In_303);
or U514 (N_514,In_705,N_87);
or U515 (N_515,N_170,N_459);
and U516 (N_516,In_578,N_117);
nor U517 (N_517,In_20,N_463);
or U518 (N_518,In_721,In_710);
nand U519 (N_519,N_149,In_961);
and U520 (N_520,N_238,N_472);
or U521 (N_521,N_488,In_448);
nor U522 (N_522,N_479,N_310);
or U523 (N_523,In_553,In_328);
or U524 (N_524,In_635,N_233);
or U525 (N_525,In_444,N_2);
nand U526 (N_526,N_262,N_406);
nand U527 (N_527,In_816,In_498);
or U528 (N_528,In_352,In_589);
nor U529 (N_529,N_452,N_151);
or U530 (N_530,In_835,In_411);
and U531 (N_531,In_240,N_93);
nand U532 (N_532,In_64,In_225);
nand U533 (N_533,In_306,N_161);
or U534 (N_534,In_787,N_454);
and U535 (N_535,N_230,N_116);
nand U536 (N_536,N_465,In_497);
and U537 (N_537,N_405,N_446);
or U538 (N_538,N_435,In_737);
nor U539 (N_539,N_461,N_338);
nand U540 (N_540,In_696,In_829);
nand U541 (N_541,In_373,In_747);
nor U542 (N_542,In_443,In_698);
nor U543 (N_543,N_146,N_466);
nor U544 (N_544,In_880,In_672);
nor U545 (N_545,In_901,N_489);
nand U546 (N_546,N_18,N_273);
nand U547 (N_547,N_370,In_688);
and U548 (N_548,N_340,N_252);
and U549 (N_549,N_427,N_467);
nor U550 (N_550,N_136,In_257);
xnor U551 (N_551,In_281,N_462);
nand U552 (N_552,In_384,N_49);
nor U553 (N_553,N_12,In_4);
or U554 (N_554,In_817,In_291);
and U555 (N_555,In_248,In_160);
or U556 (N_556,In_491,N_320);
and U557 (N_557,N_491,N_201);
and U558 (N_558,In_197,In_534);
nor U559 (N_559,N_464,N_264);
and U560 (N_560,N_443,N_430);
nor U561 (N_561,N_208,N_319);
nand U562 (N_562,In_124,N_355);
nor U563 (N_563,N_103,In_743);
or U564 (N_564,N_416,In_333);
nor U565 (N_565,In_198,N_447);
or U566 (N_566,In_604,In_157);
nand U567 (N_567,In_674,In_965);
xnor U568 (N_568,N_424,N_247);
nor U569 (N_569,N_385,In_680);
or U570 (N_570,In_0,In_35);
or U571 (N_571,N_277,N_40);
or U572 (N_572,N_282,N_227);
and U573 (N_573,In_191,In_941);
nand U574 (N_574,N_174,In_482);
nand U575 (N_575,In_43,In_334);
nor U576 (N_576,In_137,In_608);
nor U577 (N_577,N_17,N_171);
nor U578 (N_578,N_4,In_150);
or U579 (N_579,N_374,N_302);
nor U580 (N_580,N_349,N_444);
and U581 (N_581,N_487,N_474);
nor U582 (N_582,N_108,N_445);
nor U583 (N_583,N_232,N_245);
nor U584 (N_584,In_510,N_76);
nor U585 (N_585,In_323,N_200);
xnor U586 (N_586,N_417,In_75);
nand U587 (N_587,In_297,N_6);
or U588 (N_588,In_65,N_122);
nand U589 (N_589,In_447,In_479);
and U590 (N_590,N_384,N_326);
nand U591 (N_591,In_254,N_260);
and U592 (N_592,N_376,N_496);
and U593 (N_593,N_140,N_478);
and U594 (N_594,In_431,N_498);
and U595 (N_595,In_998,N_306);
nand U596 (N_596,N_334,In_984);
nor U597 (N_597,N_382,In_396);
and U598 (N_598,N_309,N_450);
nand U599 (N_599,N_354,N_199);
nor U600 (N_600,In_799,N_597);
xor U601 (N_601,N_455,N_589);
or U602 (N_602,N_249,In_562);
nor U603 (N_603,N_325,In_469);
or U604 (N_604,N_552,N_420);
or U605 (N_605,N_418,In_6);
and U606 (N_606,N_181,In_250);
nand U607 (N_607,N_404,N_486);
or U608 (N_608,N_477,N_209);
nor U609 (N_609,N_439,N_304);
nand U610 (N_610,N_74,In_762);
nand U611 (N_611,N_256,N_578);
and U612 (N_612,N_583,N_543);
and U613 (N_613,N_566,N_494);
and U614 (N_614,N_175,N_528);
and U615 (N_615,In_611,N_373);
nand U616 (N_616,In_278,In_971);
and U617 (N_617,N_89,N_128);
and U618 (N_618,N_291,N_562);
and U619 (N_619,N_32,N_386);
and U620 (N_620,In_926,N_400);
and U621 (N_621,In_375,In_558);
xor U622 (N_622,N_221,In_330);
and U623 (N_623,In_295,N_586);
or U624 (N_624,In_22,N_501);
and U625 (N_625,In_440,N_153);
and U626 (N_626,N_522,N_453);
nor U627 (N_627,N_599,N_204);
nor U628 (N_628,N_389,In_487);
or U629 (N_629,In_95,N_588);
or U630 (N_630,N_544,N_398);
or U631 (N_631,N_564,In_433);
and U632 (N_632,N_293,In_742);
nor U633 (N_633,N_495,N_198);
nor U634 (N_634,In_514,N_305);
or U635 (N_635,N_295,N_431);
nor U636 (N_636,N_421,N_584);
or U637 (N_637,N_525,N_529);
nand U638 (N_638,N_545,N_574);
nor U639 (N_639,N_541,In_679);
nand U640 (N_640,In_211,N_590);
or U641 (N_641,In_948,In_525);
and U642 (N_642,N_485,In_694);
or U643 (N_643,N_510,In_221);
or U644 (N_644,N_53,In_320);
or U645 (N_645,N_217,N_441);
nor U646 (N_646,N_323,N_480);
nor U647 (N_647,N_426,N_548);
and U648 (N_648,N_563,In_790);
nand U649 (N_649,N_1,N_598);
nor U650 (N_650,N_359,In_727);
nor U651 (N_651,In_391,N_440);
nor U652 (N_652,N_342,In_644);
nor U653 (N_653,In_337,N_357);
or U654 (N_654,N_438,In_855);
and U655 (N_655,In_651,N_422);
nor U656 (N_656,N_577,In_362);
nor U657 (N_657,N_493,N_504);
or U658 (N_658,N_471,N_585);
or U659 (N_659,N_587,N_55);
or U660 (N_660,N_162,N_393);
nor U661 (N_661,In_399,N_482);
and U662 (N_662,N_268,N_259);
or U663 (N_663,N_312,N_329);
or U664 (N_664,In_164,N_580);
and U665 (N_665,In_566,N_332);
nand U666 (N_666,N_533,N_481);
nand U667 (N_667,N_557,In_326);
nor U668 (N_668,N_576,N_364);
and U669 (N_669,In_415,In_369);
nor U670 (N_670,In_255,In_581);
nor U671 (N_671,N_526,N_569);
and U672 (N_672,In_50,N_521);
nor U673 (N_673,In_704,In_108);
nor U674 (N_674,N_353,N_509);
and U675 (N_675,N_530,In_739);
xnor U676 (N_676,In_102,In_736);
nor U677 (N_677,N_243,In_654);
xor U678 (N_678,N_65,In_107);
or U679 (N_679,N_77,N_78);
or U680 (N_680,In_712,In_811);
nand U681 (N_681,N_513,In_174);
or U682 (N_682,N_520,N_387);
nand U683 (N_683,N_514,N_591);
nand U684 (N_684,N_98,N_515);
nand U685 (N_685,N_517,In_641);
and U686 (N_686,In_324,N_272);
or U687 (N_687,N_246,In_519);
nor U688 (N_688,N_536,N_414);
or U689 (N_689,N_281,In_791);
nand U690 (N_690,N_570,N_550);
or U691 (N_691,N_429,N_592);
and U692 (N_692,In_943,In_763);
and U693 (N_693,N_538,N_298);
nand U694 (N_694,N_345,In_268);
nand U695 (N_695,N_458,N_539);
nand U696 (N_696,N_561,N_502);
nand U697 (N_697,N_470,N_511);
and U698 (N_698,N_448,In_639);
xor U699 (N_699,In_66,N_573);
or U700 (N_700,N_269,N_582);
and U701 (N_701,In_576,N_632);
or U702 (N_702,N_695,In_87);
and U703 (N_703,N_581,N_623);
nor U704 (N_704,N_660,N_685);
or U705 (N_705,In_725,In_187);
nor U706 (N_706,N_625,In_927);
nor U707 (N_707,N_670,N_542);
nand U708 (N_708,N_369,N_559);
nor U709 (N_709,N_649,N_689);
nand U710 (N_710,N_678,In_918);
or U711 (N_711,In_388,N_661);
nand U712 (N_712,N_610,N_614);
nor U713 (N_713,N_555,N_537);
or U714 (N_714,In_720,In_937);
nor U715 (N_715,N_674,N_568);
and U716 (N_716,In_466,In_309);
or U717 (N_717,N_579,N_571);
nand U718 (N_718,N_409,In_336);
nor U719 (N_719,N_656,N_601);
and U720 (N_720,In_483,N_681);
and U721 (N_721,N_433,N_691);
nand U722 (N_722,N_609,N_608);
nor U723 (N_723,N_650,N_624);
nor U724 (N_724,In_238,N_240);
nor U725 (N_725,N_92,In_991);
nand U726 (N_726,In_830,N_469);
or U727 (N_727,N_672,N_512);
and U728 (N_728,N_648,N_667);
and U729 (N_729,In_678,N_602);
and U730 (N_730,N_235,N_394);
nor U731 (N_731,N_30,In_363);
nor U732 (N_732,N_620,In_115);
or U733 (N_733,N_696,N_250);
or U734 (N_734,N_575,N_253);
nand U735 (N_735,In_573,N_535);
and U736 (N_736,N_523,N_638);
or U737 (N_737,In_848,In_740);
and U738 (N_738,N_527,In_814);
xnor U739 (N_739,In_344,In_507);
or U740 (N_740,N_628,N_21);
and U741 (N_741,N_643,In_181);
or U742 (N_742,In_171,N_395);
and U743 (N_743,N_490,In_386);
or U744 (N_744,N_224,In_318);
nor U745 (N_745,N_647,N_499);
nor U746 (N_746,N_492,N_366);
nor U747 (N_747,N_316,N_457);
or U748 (N_748,N_451,N_636);
nand U749 (N_749,N_633,N_344);
or U750 (N_750,N_120,N_88);
nand U751 (N_751,N_551,N_692);
and U752 (N_752,In_593,N_216);
nor U753 (N_753,N_679,N_687);
and U754 (N_754,N_565,N_425);
or U755 (N_755,N_682,N_350);
nor U756 (N_756,N_402,N_519);
or U757 (N_757,N_640,N_38);
nor U758 (N_758,N_690,N_506);
nor U759 (N_759,N_531,N_669);
nor U760 (N_760,In_713,N_596);
nor U761 (N_761,N_500,In_556);
or U762 (N_762,N_412,In_260);
or U763 (N_763,In_668,N_641);
or U764 (N_764,In_518,N_635);
and U765 (N_765,N_572,N_518);
or U766 (N_766,N_558,In_803);
or U767 (N_767,N_505,N_9);
or U768 (N_768,N_677,N_616);
and U769 (N_769,N_388,N_401);
nand U770 (N_770,N_604,N_507);
nand U771 (N_771,N_651,N_372);
or U772 (N_772,N_410,In_13);
and U773 (N_773,N_358,N_43);
nor U774 (N_774,N_413,N_549);
xnor U775 (N_775,In_111,N_303);
nor U776 (N_776,In_782,N_688);
xnor U777 (N_777,N_280,N_605);
nor U778 (N_778,In_996,N_622);
nand U779 (N_779,In_460,N_328);
or U780 (N_780,N_460,N_634);
nand U781 (N_781,N_639,N_693);
nor U782 (N_782,N_399,In_305);
or U783 (N_783,N_567,N_339);
or U784 (N_784,N_419,In_348);
and U785 (N_785,N_475,N_631);
or U786 (N_786,In_185,N_668);
and U787 (N_787,N_408,N_202);
and U788 (N_788,In_189,In_61);
nor U789 (N_789,N_483,N_653);
and U790 (N_790,N_627,N_254);
or U791 (N_791,In_542,N_654);
nor U792 (N_792,N_676,N_348);
nor U793 (N_793,N_185,N_560);
or U794 (N_794,In_284,N_378);
nand U795 (N_795,N_524,N_428);
nor U796 (N_796,N_532,N_331);
nand U797 (N_797,N_593,N_662);
and U798 (N_798,N_267,N_686);
nand U799 (N_799,N_606,In_579);
and U800 (N_800,N_664,In_332);
and U801 (N_801,N_756,N_618);
or U802 (N_802,N_703,N_799);
nor U803 (N_803,N_725,N_646);
nor U804 (N_804,N_757,N_710);
nand U805 (N_805,N_721,N_698);
nand U806 (N_806,N_724,N_335);
or U807 (N_807,N_595,In_387);
or U808 (N_808,N_82,N_706);
nand U809 (N_809,In_919,N_257);
and U810 (N_810,N_226,N_336);
or U811 (N_811,N_755,N_380);
or U812 (N_812,N_720,N_468);
and U813 (N_813,N_671,N_164);
nand U814 (N_814,N_795,N_746);
and U815 (N_815,N_613,N_351);
nand U816 (N_816,N_379,N_423);
and U817 (N_817,N_629,N_556);
nand U818 (N_818,N_699,N_665);
and U819 (N_819,N_315,N_763);
nand U820 (N_820,N_717,N_449);
or U821 (N_821,In_993,In_986);
and U822 (N_822,N_701,N_637);
or U823 (N_823,N_769,N_657);
nor U824 (N_824,N_767,N_733);
nor U825 (N_825,N_700,N_781);
nand U826 (N_826,N_716,N_553);
nor U827 (N_827,N_534,N_792);
nand U828 (N_828,N_621,N_707);
and U829 (N_829,In_478,N_791);
or U830 (N_830,N_630,N_619);
nor U831 (N_831,N_626,N_758);
or U832 (N_832,N_540,N_645);
or U833 (N_833,N_658,N_684);
or U834 (N_834,N_730,N_785);
nand U835 (N_835,N_704,N_702);
nand U836 (N_836,N_777,N_752);
nor U837 (N_837,N_697,N_796);
or U838 (N_838,N_516,In_847);
nand U839 (N_839,N_731,N_786);
nor U840 (N_840,N_783,N_764);
nand U841 (N_841,N_683,N_663);
or U842 (N_842,N_166,In_315);
nand U843 (N_843,N_322,N_600);
nand U844 (N_844,In_239,In_990);
nand U845 (N_845,N_123,N_714);
and U846 (N_846,In_88,N_773);
or U847 (N_847,N_787,N_770);
or U848 (N_848,N_794,N_748);
or U849 (N_849,N_727,N_75);
nand U850 (N_850,N_709,N_719);
or U851 (N_851,N_324,N_789);
nor U852 (N_852,N_713,N_780);
nor U853 (N_853,N_776,In_784);
nor U854 (N_854,In_125,N_722);
nor U855 (N_855,N_508,In_768);
nor U856 (N_856,N_680,N_738);
or U857 (N_857,N_712,N_749);
or U858 (N_858,N_790,N_766);
or U859 (N_859,N_747,N_611);
and U860 (N_860,N_782,N_615);
nand U861 (N_861,In_59,N_761);
or U862 (N_862,N_156,N_675);
and U863 (N_863,N_788,N_723);
nor U864 (N_864,N_133,In_503);
and U865 (N_865,N_751,N_705);
nor U866 (N_866,N_244,N_617);
and U867 (N_867,N_659,N_775);
or U868 (N_868,N_711,N_607);
nand U869 (N_869,N_652,N_784);
or U870 (N_870,N_735,N_797);
and U871 (N_871,N_708,N_753);
or U872 (N_872,N_778,N_772);
and U873 (N_873,N_726,N_715);
nor U874 (N_874,N_793,N_603);
or U875 (N_875,In_537,N_798);
nand U876 (N_876,In_949,N_728);
nand U877 (N_877,N_742,N_363);
or U878 (N_878,N_497,N_760);
nand U879 (N_879,N_655,N_754);
or U880 (N_880,N_762,N_736);
or U881 (N_881,N_673,N_737);
nor U882 (N_882,N_744,N_546);
or U883 (N_883,N_275,N_547);
or U884 (N_884,N_594,N_745);
or U885 (N_885,N_768,In_222);
and U886 (N_886,N_642,N_718);
nor U887 (N_887,N_759,N_771);
nor U888 (N_888,N_774,N_779);
and U889 (N_889,N_612,In_40);
xor U890 (N_890,N_644,N_765);
nand U891 (N_891,N_740,N_554);
nand U892 (N_892,N_750,N_666);
nor U893 (N_893,N_732,N_694);
or U894 (N_894,N_503,N_210);
or U895 (N_895,N_729,N_437);
nand U896 (N_896,In_457,N_436);
or U897 (N_897,N_743,N_739);
nor U898 (N_898,N_311,N_741);
nor U899 (N_899,In_11,N_734);
and U900 (N_900,N_840,N_830);
nor U901 (N_901,N_865,N_863);
nand U902 (N_902,N_835,N_882);
nand U903 (N_903,N_822,N_883);
and U904 (N_904,N_856,N_838);
nand U905 (N_905,N_801,N_869);
and U906 (N_906,N_820,N_843);
nand U907 (N_907,N_897,N_800);
and U908 (N_908,N_825,N_847);
or U909 (N_909,N_808,N_898);
and U910 (N_910,N_829,N_827);
nand U911 (N_911,N_845,N_852);
nand U912 (N_912,N_894,N_862);
xor U913 (N_913,N_864,N_871);
and U914 (N_914,N_804,N_855);
nor U915 (N_915,N_893,N_816);
nand U916 (N_916,N_859,N_889);
nand U917 (N_917,N_876,N_886);
and U918 (N_918,N_826,N_880);
or U919 (N_919,N_848,N_851);
nand U920 (N_920,N_807,N_841);
or U921 (N_921,N_824,N_805);
and U922 (N_922,N_890,N_812);
nor U923 (N_923,N_823,N_818);
xnor U924 (N_924,N_821,N_839);
nor U925 (N_925,N_860,N_850);
nand U926 (N_926,N_809,N_874);
and U927 (N_927,N_803,N_861);
nand U928 (N_928,N_888,N_857);
and U929 (N_929,N_875,N_873);
and U930 (N_930,N_837,N_899);
or U931 (N_931,N_814,N_881);
nor U932 (N_932,N_819,N_833);
or U933 (N_933,N_842,N_896);
and U934 (N_934,N_884,N_891);
and U935 (N_935,N_895,N_877);
xnor U936 (N_936,N_802,N_834);
or U937 (N_937,N_844,N_828);
nor U938 (N_938,N_879,N_892);
nor U939 (N_939,N_846,N_811);
or U940 (N_940,N_866,N_887);
or U941 (N_941,N_815,N_870);
nor U942 (N_942,N_885,N_868);
and U943 (N_943,N_853,N_872);
or U944 (N_944,N_832,N_813);
nand U945 (N_945,N_806,N_867);
or U946 (N_946,N_858,N_810);
nand U947 (N_947,N_878,N_849);
nor U948 (N_948,N_854,N_836);
nand U949 (N_949,N_831,N_817);
nor U950 (N_950,N_862,N_884);
or U951 (N_951,N_815,N_812);
and U952 (N_952,N_821,N_808);
nand U953 (N_953,N_892,N_849);
or U954 (N_954,N_800,N_866);
and U955 (N_955,N_859,N_848);
and U956 (N_956,N_853,N_824);
or U957 (N_957,N_859,N_867);
nor U958 (N_958,N_853,N_834);
or U959 (N_959,N_852,N_826);
and U960 (N_960,N_803,N_830);
or U961 (N_961,N_836,N_845);
and U962 (N_962,N_815,N_833);
and U963 (N_963,N_814,N_850);
nand U964 (N_964,N_872,N_856);
xor U965 (N_965,N_881,N_822);
or U966 (N_966,N_885,N_888);
or U967 (N_967,N_867,N_803);
and U968 (N_968,N_817,N_815);
xnor U969 (N_969,N_802,N_850);
nor U970 (N_970,N_895,N_814);
nor U971 (N_971,N_879,N_816);
nor U972 (N_972,N_858,N_814);
or U973 (N_973,N_827,N_813);
or U974 (N_974,N_806,N_848);
nor U975 (N_975,N_874,N_852);
and U976 (N_976,N_871,N_811);
and U977 (N_977,N_803,N_851);
or U978 (N_978,N_843,N_876);
nand U979 (N_979,N_803,N_838);
and U980 (N_980,N_858,N_801);
or U981 (N_981,N_890,N_888);
nor U982 (N_982,N_859,N_814);
nor U983 (N_983,N_848,N_863);
nor U984 (N_984,N_825,N_899);
nand U985 (N_985,N_839,N_877);
and U986 (N_986,N_821,N_846);
nand U987 (N_987,N_843,N_885);
and U988 (N_988,N_860,N_888);
nor U989 (N_989,N_820,N_857);
or U990 (N_990,N_864,N_803);
nor U991 (N_991,N_835,N_853);
or U992 (N_992,N_870,N_819);
nor U993 (N_993,N_863,N_814);
nor U994 (N_994,N_846,N_832);
nor U995 (N_995,N_881,N_827);
nor U996 (N_996,N_836,N_818);
nor U997 (N_997,N_886,N_817);
nand U998 (N_998,N_889,N_887);
and U999 (N_999,N_828,N_848);
and U1000 (N_1000,N_958,N_985);
and U1001 (N_1001,N_975,N_906);
nor U1002 (N_1002,N_996,N_917);
or U1003 (N_1003,N_999,N_982);
nand U1004 (N_1004,N_910,N_907);
and U1005 (N_1005,N_993,N_913);
nand U1006 (N_1006,N_971,N_938);
or U1007 (N_1007,N_937,N_987);
nand U1008 (N_1008,N_943,N_900);
nor U1009 (N_1009,N_902,N_960);
nand U1010 (N_1010,N_966,N_926);
nor U1011 (N_1011,N_961,N_939);
or U1012 (N_1012,N_945,N_918);
and U1013 (N_1013,N_955,N_935);
and U1014 (N_1014,N_931,N_977);
nor U1015 (N_1015,N_981,N_924);
or U1016 (N_1016,N_928,N_951);
or U1017 (N_1017,N_954,N_933);
nor U1018 (N_1018,N_979,N_923);
nand U1019 (N_1019,N_949,N_984);
nand U1020 (N_1020,N_976,N_932);
and U1021 (N_1021,N_950,N_919);
and U1022 (N_1022,N_957,N_930);
or U1023 (N_1023,N_922,N_973);
nor U1024 (N_1024,N_940,N_988);
or U1025 (N_1025,N_969,N_974);
nand U1026 (N_1026,N_992,N_916);
and U1027 (N_1027,N_952,N_911);
or U1028 (N_1028,N_963,N_994);
and U1029 (N_1029,N_991,N_909);
nor U1030 (N_1030,N_962,N_990);
xor U1031 (N_1031,N_944,N_912);
and U1032 (N_1032,N_948,N_920);
or U1033 (N_1033,N_905,N_998);
and U1034 (N_1034,N_983,N_995);
nor U1035 (N_1035,N_929,N_947);
nand U1036 (N_1036,N_964,N_970);
nor U1037 (N_1037,N_915,N_901);
or U1038 (N_1038,N_978,N_904);
nor U1039 (N_1039,N_967,N_934);
or U1040 (N_1040,N_925,N_903);
nor U1041 (N_1041,N_927,N_953);
or U1042 (N_1042,N_921,N_908);
xnor U1043 (N_1043,N_942,N_956);
nor U1044 (N_1044,N_997,N_968);
nor U1045 (N_1045,N_965,N_941);
nand U1046 (N_1046,N_946,N_914);
nand U1047 (N_1047,N_980,N_986);
and U1048 (N_1048,N_972,N_989);
nand U1049 (N_1049,N_959,N_936);
and U1050 (N_1050,N_967,N_980);
nand U1051 (N_1051,N_991,N_978);
nand U1052 (N_1052,N_977,N_901);
nand U1053 (N_1053,N_944,N_996);
nand U1054 (N_1054,N_940,N_900);
nor U1055 (N_1055,N_997,N_972);
or U1056 (N_1056,N_904,N_971);
nor U1057 (N_1057,N_922,N_942);
nand U1058 (N_1058,N_921,N_944);
and U1059 (N_1059,N_920,N_934);
nor U1060 (N_1060,N_938,N_952);
or U1061 (N_1061,N_908,N_987);
nand U1062 (N_1062,N_981,N_978);
nand U1063 (N_1063,N_975,N_988);
or U1064 (N_1064,N_923,N_913);
or U1065 (N_1065,N_983,N_905);
xor U1066 (N_1066,N_985,N_929);
nand U1067 (N_1067,N_973,N_982);
and U1068 (N_1068,N_945,N_939);
nor U1069 (N_1069,N_958,N_907);
and U1070 (N_1070,N_944,N_986);
or U1071 (N_1071,N_902,N_973);
nor U1072 (N_1072,N_922,N_934);
and U1073 (N_1073,N_950,N_973);
nor U1074 (N_1074,N_909,N_922);
or U1075 (N_1075,N_930,N_973);
nand U1076 (N_1076,N_984,N_968);
nor U1077 (N_1077,N_915,N_992);
nor U1078 (N_1078,N_933,N_917);
or U1079 (N_1079,N_993,N_954);
nand U1080 (N_1080,N_902,N_985);
and U1081 (N_1081,N_990,N_925);
and U1082 (N_1082,N_945,N_979);
nand U1083 (N_1083,N_975,N_920);
and U1084 (N_1084,N_935,N_971);
nor U1085 (N_1085,N_978,N_939);
nor U1086 (N_1086,N_968,N_954);
nor U1087 (N_1087,N_960,N_998);
nor U1088 (N_1088,N_966,N_985);
and U1089 (N_1089,N_966,N_993);
nand U1090 (N_1090,N_943,N_997);
or U1091 (N_1091,N_977,N_955);
nor U1092 (N_1092,N_963,N_980);
or U1093 (N_1093,N_908,N_990);
nand U1094 (N_1094,N_968,N_993);
or U1095 (N_1095,N_977,N_942);
nor U1096 (N_1096,N_942,N_987);
nor U1097 (N_1097,N_975,N_945);
and U1098 (N_1098,N_985,N_984);
nor U1099 (N_1099,N_949,N_912);
nand U1100 (N_1100,N_1024,N_1013);
nor U1101 (N_1101,N_1062,N_1064);
and U1102 (N_1102,N_1090,N_1035);
nor U1103 (N_1103,N_1077,N_1020);
or U1104 (N_1104,N_1083,N_1008);
and U1105 (N_1105,N_1087,N_1068);
and U1106 (N_1106,N_1032,N_1001);
nand U1107 (N_1107,N_1006,N_1086);
or U1108 (N_1108,N_1040,N_1017);
nor U1109 (N_1109,N_1033,N_1003);
and U1110 (N_1110,N_1053,N_1073);
or U1111 (N_1111,N_1039,N_1000);
nand U1112 (N_1112,N_1031,N_1014);
or U1113 (N_1113,N_1036,N_1060);
nor U1114 (N_1114,N_1037,N_1059);
and U1115 (N_1115,N_1061,N_1079);
nand U1116 (N_1116,N_1080,N_1047);
nand U1117 (N_1117,N_1030,N_1051);
nand U1118 (N_1118,N_1048,N_1004);
and U1119 (N_1119,N_1094,N_1071);
and U1120 (N_1120,N_1042,N_1043);
nor U1121 (N_1121,N_1056,N_1029);
xnor U1122 (N_1122,N_1055,N_1066);
or U1123 (N_1123,N_1085,N_1049);
nor U1124 (N_1124,N_1082,N_1088);
and U1125 (N_1125,N_1044,N_1019);
nand U1126 (N_1126,N_1023,N_1016);
or U1127 (N_1127,N_1063,N_1050);
nand U1128 (N_1128,N_1069,N_1093);
or U1129 (N_1129,N_1089,N_1026);
or U1130 (N_1130,N_1010,N_1011);
nor U1131 (N_1131,N_1041,N_1078);
and U1132 (N_1132,N_1072,N_1058);
nand U1133 (N_1133,N_1096,N_1021);
nand U1134 (N_1134,N_1067,N_1046);
nor U1135 (N_1135,N_1091,N_1075);
and U1136 (N_1136,N_1018,N_1074);
nor U1137 (N_1137,N_1081,N_1099);
or U1138 (N_1138,N_1065,N_1038);
and U1139 (N_1139,N_1057,N_1002);
and U1140 (N_1140,N_1098,N_1007);
or U1141 (N_1141,N_1045,N_1025);
or U1142 (N_1142,N_1005,N_1028);
and U1143 (N_1143,N_1097,N_1034);
nand U1144 (N_1144,N_1022,N_1084);
and U1145 (N_1145,N_1015,N_1095);
nor U1146 (N_1146,N_1052,N_1027);
and U1147 (N_1147,N_1054,N_1009);
nand U1148 (N_1148,N_1092,N_1076);
or U1149 (N_1149,N_1070,N_1012);
and U1150 (N_1150,N_1032,N_1020);
nand U1151 (N_1151,N_1066,N_1075);
nand U1152 (N_1152,N_1085,N_1027);
nor U1153 (N_1153,N_1070,N_1085);
or U1154 (N_1154,N_1020,N_1002);
xnor U1155 (N_1155,N_1049,N_1032);
and U1156 (N_1156,N_1027,N_1050);
nor U1157 (N_1157,N_1091,N_1012);
and U1158 (N_1158,N_1056,N_1064);
or U1159 (N_1159,N_1080,N_1049);
nor U1160 (N_1160,N_1037,N_1044);
and U1161 (N_1161,N_1040,N_1061);
xnor U1162 (N_1162,N_1053,N_1033);
and U1163 (N_1163,N_1032,N_1088);
nand U1164 (N_1164,N_1025,N_1089);
and U1165 (N_1165,N_1020,N_1061);
xnor U1166 (N_1166,N_1000,N_1075);
and U1167 (N_1167,N_1099,N_1066);
nor U1168 (N_1168,N_1065,N_1005);
and U1169 (N_1169,N_1059,N_1043);
xor U1170 (N_1170,N_1064,N_1074);
nor U1171 (N_1171,N_1068,N_1078);
nand U1172 (N_1172,N_1090,N_1096);
or U1173 (N_1173,N_1094,N_1051);
or U1174 (N_1174,N_1099,N_1076);
or U1175 (N_1175,N_1091,N_1037);
nand U1176 (N_1176,N_1057,N_1080);
nand U1177 (N_1177,N_1087,N_1082);
and U1178 (N_1178,N_1040,N_1049);
nor U1179 (N_1179,N_1055,N_1040);
nand U1180 (N_1180,N_1010,N_1040);
and U1181 (N_1181,N_1098,N_1016);
nor U1182 (N_1182,N_1054,N_1028);
or U1183 (N_1183,N_1004,N_1039);
and U1184 (N_1184,N_1086,N_1070);
or U1185 (N_1185,N_1039,N_1029);
nand U1186 (N_1186,N_1080,N_1002);
nor U1187 (N_1187,N_1003,N_1099);
and U1188 (N_1188,N_1097,N_1080);
nor U1189 (N_1189,N_1017,N_1025);
nor U1190 (N_1190,N_1003,N_1065);
nand U1191 (N_1191,N_1068,N_1019);
nor U1192 (N_1192,N_1017,N_1097);
nand U1193 (N_1193,N_1090,N_1080);
nor U1194 (N_1194,N_1036,N_1029);
or U1195 (N_1195,N_1065,N_1093);
and U1196 (N_1196,N_1033,N_1084);
nor U1197 (N_1197,N_1019,N_1002);
nand U1198 (N_1198,N_1052,N_1034);
and U1199 (N_1199,N_1002,N_1077);
nand U1200 (N_1200,N_1137,N_1149);
or U1201 (N_1201,N_1152,N_1140);
or U1202 (N_1202,N_1158,N_1181);
and U1203 (N_1203,N_1183,N_1131);
or U1204 (N_1204,N_1128,N_1147);
xor U1205 (N_1205,N_1136,N_1103);
nand U1206 (N_1206,N_1173,N_1150);
xor U1207 (N_1207,N_1100,N_1105);
xnor U1208 (N_1208,N_1113,N_1160);
nand U1209 (N_1209,N_1104,N_1139);
nor U1210 (N_1210,N_1108,N_1117);
nand U1211 (N_1211,N_1166,N_1195);
nor U1212 (N_1212,N_1143,N_1172);
nand U1213 (N_1213,N_1118,N_1159);
or U1214 (N_1214,N_1188,N_1193);
and U1215 (N_1215,N_1138,N_1156);
or U1216 (N_1216,N_1151,N_1164);
nor U1217 (N_1217,N_1178,N_1132);
nor U1218 (N_1218,N_1162,N_1174);
and U1219 (N_1219,N_1194,N_1192);
nand U1220 (N_1220,N_1126,N_1161);
and U1221 (N_1221,N_1106,N_1199);
and U1222 (N_1222,N_1191,N_1107);
nor U1223 (N_1223,N_1180,N_1120);
and U1224 (N_1224,N_1145,N_1125);
nor U1225 (N_1225,N_1185,N_1189);
nor U1226 (N_1226,N_1163,N_1169);
nor U1227 (N_1227,N_1121,N_1119);
or U1228 (N_1228,N_1127,N_1142);
or U1229 (N_1229,N_1116,N_1135);
nand U1230 (N_1230,N_1154,N_1101);
nor U1231 (N_1231,N_1114,N_1130);
nor U1232 (N_1232,N_1153,N_1129);
and U1233 (N_1233,N_1184,N_1133);
nor U1234 (N_1234,N_1171,N_1123);
xor U1235 (N_1235,N_1190,N_1111);
and U1236 (N_1236,N_1168,N_1148);
or U1237 (N_1237,N_1167,N_1196);
nand U1238 (N_1238,N_1175,N_1155);
nor U1239 (N_1239,N_1144,N_1146);
or U1240 (N_1240,N_1179,N_1177);
or U1241 (N_1241,N_1187,N_1186);
and U1242 (N_1242,N_1198,N_1102);
nor U1243 (N_1243,N_1115,N_1182);
or U1244 (N_1244,N_1157,N_1197);
nor U1245 (N_1245,N_1165,N_1176);
nor U1246 (N_1246,N_1170,N_1124);
and U1247 (N_1247,N_1134,N_1109);
or U1248 (N_1248,N_1122,N_1141);
and U1249 (N_1249,N_1112,N_1110);
and U1250 (N_1250,N_1137,N_1168);
nand U1251 (N_1251,N_1114,N_1107);
nand U1252 (N_1252,N_1147,N_1101);
nor U1253 (N_1253,N_1128,N_1117);
nor U1254 (N_1254,N_1104,N_1154);
nand U1255 (N_1255,N_1197,N_1156);
and U1256 (N_1256,N_1167,N_1195);
and U1257 (N_1257,N_1132,N_1189);
nor U1258 (N_1258,N_1169,N_1107);
nand U1259 (N_1259,N_1153,N_1171);
nand U1260 (N_1260,N_1100,N_1137);
nand U1261 (N_1261,N_1111,N_1120);
nand U1262 (N_1262,N_1157,N_1123);
and U1263 (N_1263,N_1146,N_1102);
nand U1264 (N_1264,N_1157,N_1112);
and U1265 (N_1265,N_1101,N_1189);
or U1266 (N_1266,N_1188,N_1110);
nand U1267 (N_1267,N_1120,N_1174);
nor U1268 (N_1268,N_1192,N_1124);
nor U1269 (N_1269,N_1188,N_1173);
and U1270 (N_1270,N_1153,N_1120);
and U1271 (N_1271,N_1127,N_1130);
and U1272 (N_1272,N_1185,N_1193);
nor U1273 (N_1273,N_1134,N_1157);
xor U1274 (N_1274,N_1115,N_1156);
nor U1275 (N_1275,N_1199,N_1155);
nor U1276 (N_1276,N_1175,N_1148);
or U1277 (N_1277,N_1118,N_1106);
nand U1278 (N_1278,N_1119,N_1174);
nor U1279 (N_1279,N_1185,N_1191);
nor U1280 (N_1280,N_1153,N_1148);
and U1281 (N_1281,N_1116,N_1131);
and U1282 (N_1282,N_1170,N_1115);
nand U1283 (N_1283,N_1183,N_1145);
xnor U1284 (N_1284,N_1147,N_1113);
nor U1285 (N_1285,N_1139,N_1132);
nor U1286 (N_1286,N_1199,N_1188);
xnor U1287 (N_1287,N_1188,N_1178);
or U1288 (N_1288,N_1108,N_1190);
or U1289 (N_1289,N_1172,N_1108);
nand U1290 (N_1290,N_1127,N_1185);
nor U1291 (N_1291,N_1174,N_1139);
or U1292 (N_1292,N_1174,N_1118);
nand U1293 (N_1293,N_1126,N_1112);
nor U1294 (N_1294,N_1159,N_1144);
or U1295 (N_1295,N_1155,N_1198);
or U1296 (N_1296,N_1145,N_1138);
xor U1297 (N_1297,N_1144,N_1140);
nor U1298 (N_1298,N_1134,N_1178);
nor U1299 (N_1299,N_1110,N_1134);
or U1300 (N_1300,N_1240,N_1291);
or U1301 (N_1301,N_1255,N_1229);
nand U1302 (N_1302,N_1266,N_1289);
or U1303 (N_1303,N_1269,N_1271);
nor U1304 (N_1304,N_1230,N_1287);
or U1305 (N_1305,N_1254,N_1239);
or U1306 (N_1306,N_1284,N_1231);
nor U1307 (N_1307,N_1264,N_1296);
and U1308 (N_1308,N_1272,N_1223);
or U1309 (N_1309,N_1250,N_1293);
nand U1310 (N_1310,N_1224,N_1292);
nor U1311 (N_1311,N_1218,N_1256);
nor U1312 (N_1312,N_1281,N_1200);
and U1313 (N_1313,N_1245,N_1216);
or U1314 (N_1314,N_1244,N_1290);
and U1315 (N_1315,N_1215,N_1258);
or U1316 (N_1316,N_1273,N_1225);
and U1317 (N_1317,N_1213,N_1247);
nor U1318 (N_1318,N_1210,N_1220);
nor U1319 (N_1319,N_1263,N_1207);
and U1320 (N_1320,N_1288,N_1236);
nor U1321 (N_1321,N_1246,N_1252);
nand U1322 (N_1322,N_1285,N_1276);
nand U1323 (N_1323,N_1203,N_1261);
nand U1324 (N_1324,N_1279,N_1278);
nor U1325 (N_1325,N_1283,N_1275);
or U1326 (N_1326,N_1211,N_1238);
nand U1327 (N_1327,N_1205,N_1274);
or U1328 (N_1328,N_1201,N_1259);
nor U1329 (N_1329,N_1265,N_1257);
nand U1330 (N_1330,N_1249,N_1268);
and U1331 (N_1331,N_1217,N_1282);
and U1332 (N_1332,N_1297,N_1227);
nor U1333 (N_1333,N_1248,N_1270);
and U1334 (N_1334,N_1209,N_1262);
nand U1335 (N_1335,N_1212,N_1234);
and U1336 (N_1336,N_1298,N_1228);
nor U1337 (N_1337,N_1208,N_1222);
nor U1338 (N_1338,N_1260,N_1243);
nand U1339 (N_1339,N_1253,N_1206);
nand U1340 (N_1340,N_1286,N_1232);
nor U1341 (N_1341,N_1235,N_1280);
or U1342 (N_1342,N_1299,N_1267);
nor U1343 (N_1343,N_1277,N_1202);
nand U1344 (N_1344,N_1204,N_1233);
and U1345 (N_1345,N_1214,N_1221);
or U1346 (N_1346,N_1219,N_1295);
xor U1347 (N_1347,N_1237,N_1241);
and U1348 (N_1348,N_1294,N_1226);
or U1349 (N_1349,N_1251,N_1242);
nor U1350 (N_1350,N_1246,N_1245);
nor U1351 (N_1351,N_1210,N_1277);
or U1352 (N_1352,N_1247,N_1265);
and U1353 (N_1353,N_1256,N_1264);
xor U1354 (N_1354,N_1255,N_1288);
and U1355 (N_1355,N_1217,N_1259);
and U1356 (N_1356,N_1279,N_1208);
and U1357 (N_1357,N_1216,N_1293);
or U1358 (N_1358,N_1289,N_1220);
nand U1359 (N_1359,N_1226,N_1293);
or U1360 (N_1360,N_1236,N_1225);
nor U1361 (N_1361,N_1286,N_1243);
nor U1362 (N_1362,N_1275,N_1205);
nand U1363 (N_1363,N_1212,N_1285);
nor U1364 (N_1364,N_1267,N_1226);
nand U1365 (N_1365,N_1257,N_1235);
and U1366 (N_1366,N_1234,N_1268);
or U1367 (N_1367,N_1291,N_1285);
and U1368 (N_1368,N_1277,N_1248);
and U1369 (N_1369,N_1296,N_1247);
and U1370 (N_1370,N_1207,N_1203);
nand U1371 (N_1371,N_1240,N_1234);
nand U1372 (N_1372,N_1231,N_1247);
or U1373 (N_1373,N_1263,N_1298);
nor U1374 (N_1374,N_1258,N_1206);
or U1375 (N_1375,N_1250,N_1244);
or U1376 (N_1376,N_1211,N_1208);
or U1377 (N_1377,N_1264,N_1219);
nand U1378 (N_1378,N_1253,N_1282);
and U1379 (N_1379,N_1257,N_1217);
nand U1380 (N_1380,N_1243,N_1234);
or U1381 (N_1381,N_1218,N_1244);
nor U1382 (N_1382,N_1266,N_1253);
nor U1383 (N_1383,N_1274,N_1235);
nand U1384 (N_1384,N_1272,N_1240);
and U1385 (N_1385,N_1216,N_1233);
nor U1386 (N_1386,N_1206,N_1213);
or U1387 (N_1387,N_1222,N_1261);
nand U1388 (N_1388,N_1295,N_1211);
nand U1389 (N_1389,N_1232,N_1201);
xnor U1390 (N_1390,N_1287,N_1201);
or U1391 (N_1391,N_1203,N_1216);
and U1392 (N_1392,N_1212,N_1247);
or U1393 (N_1393,N_1281,N_1211);
nor U1394 (N_1394,N_1239,N_1284);
or U1395 (N_1395,N_1270,N_1273);
nor U1396 (N_1396,N_1283,N_1277);
nor U1397 (N_1397,N_1296,N_1213);
nor U1398 (N_1398,N_1214,N_1294);
and U1399 (N_1399,N_1253,N_1202);
xor U1400 (N_1400,N_1398,N_1375);
nand U1401 (N_1401,N_1378,N_1381);
or U1402 (N_1402,N_1362,N_1396);
and U1403 (N_1403,N_1370,N_1322);
nand U1404 (N_1404,N_1351,N_1331);
and U1405 (N_1405,N_1350,N_1399);
nor U1406 (N_1406,N_1366,N_1367);
or U1407 (N_1407,N_1315,N_1326);
and U1408 (N_1408,N_1386,N_1348);
or U1409 (N_1409,N_1302,N_1365);
nand U1410 (N_1410,N_1313,N_1377);
nor U1411 (N_1411,N_1358,N_1374);
and U1412 (N_1412,N_1392,N_1333);
nor U1413 (N_1413,N_1300,N_1349);
nor U1414 (N_1414,N_1363,N_1305);
nand U1415 (N_1415,N_1376,N_1371);
and U1416 (N_1416,N_1373,N_1352);
and U1417 (N_1417,N_1321,N_1328);
nor U1418 (N_1418,N_1341,N_1380);
or U1419 (N_1419,N_1337,N_1336);
or U1420 (N_1420,N_1369,N_1382);
nor U1421 (N_1421,N_1359,N_1389);
nand U1422 (N_1422,N_1372,N_1339);
nand U1423 (N_1423,N_1356,N_1368);
and U1424 (N_1424,N_1338,N_1393);
nor U1425 (N_1425,N_1388,N_1320);
or U1426 (N_1426,N_1329,N_1355);
and U1427 (N_1427,N_1311,N_1317);
or U1428 (N_1428,N_1301,N_1361);
and U1429 (N_1429,N_1391,N_1357);
nand U1430 (N_1430,N_1384,N_1335);
nand U1431 (N_1431,N_1307,N_1342);
and U1432 (N_1432,N_1385,N_1397);
and U1433 (N_1433,N_1387,N_1309);
or U1434 (N_1434,N_1324,N_1310);
nor U1435 (N_1435,N_1303,N_1308);
or U1436 (N_1436,N_1360,N_1340);
and U1437 (N_1437,N_1330,N_1379);
nor U1438 (N_1438,N_1353,N_1332);
or U1439 (N_1439,N_1306,N_1314);
nor U1440 (N_1440,N_1304,N_1364);
or U1441 (N_1441,N_1323,N_1345);
nor U1442 (N_1442,N_1344,N_1343);
nand U1443 (N_1443,N_1318,N_1319);
and U1444 (N_1444,N_1325,N_1390);
and U1445 (N_1445,N_1316,N_1346);
nand U1446 (N_1446,N_1327,N_1395);
and U1447 (N_1447,N_1347,N_1312);
nand U1448 (N_1448,N_1334,N_1394);
and U1449 (N_1449,N_1354,N_1383);
and U1450 (N_1450,N_1380,N_1377);
nand U1451 (N_1451,N_1331,N_1348);
nor U1452 (N_1452,N_1335,N_1389);
xor U1453 (N_1453,N_1393,N_1313);
nor U1454 (N_1454,N_1315,N_1308);
or U1455 (N_1455,N_1319,N_1336);
and U1456 (N_1456,N_1398,N_1339);
nor U1457 (N_1457,N_1313,N_1318);
nor U1458 (N_1458,N_1370,N_1323);
nor U1459 (N_1459,N_1360,N_1362);
and U1460 (N_1460,N_1373,N_1310);
nand U1461 (N_1461,N_1328,N_1385);
nand U1462 (N_1462,N_1325,N_1303);
nor U1463 (N_1463,N_1333,N_1316);
or U1464 (N_1464,N_1314,N_1323);
and U1465 (N_1465,N_1394,N_1390);
or U1466 (N_1466,N_1309,N_1375);
nand U1467 (N_1467,N_1374,N_1399);
or U1468 (N_1468,N_1318,N_1310);
or U1469 (N_1469,N_1376,N_1372);
nor U1470 (N_1470,N_1314,N_1334);
nand U1471 (N_1471,N_1340,N_1363);
nor U1472 (N_1472,N_1308,N_1356);
nor U1473 (N_1473,N_1311,N_1357);
nand U1474 (N_1474,N_1351,N_1382);
nand U1475 (N_1475,N_1399,N_1342);
and U1476 (N_1476,N_1376,N_1314);
and U1477 (N_1477,N_1354,N_1399);
nand U1478 (N_1478,N_1370,N_1352);
nand U1479 (N_1479,N_1301,N_1320);
nand U1480 (N_1480,N_1353,N_1301);
nor U1481 (N_1481,N_1335,N_1318);
or U1482 (N_1482,N_1383,N_1365);
nor U1483 (N_1483,N_1336,N_1373);
or U1484 (N_1484,N_1385,N_1350);
nand U1485 (N_1485,N_1350,N_1384);
or U1486 (N_1486,N_1352,N_1366);
nand U1487 (N_1487,N_1364,N_1373);
and U1488 (N_1488,N_1394,N_1363);
nor U1489 (N_1489,N_1347,N_1361);
and U1490 (N_1490,N_1300,N_1398);
nand U1491 (N_1491,N_1387,N_1355);
nor U1492 (N_1492,N_1313,N_1314);
nor U1493 (N_1493,N_1327,N_1306);
and U1494 (N_1494,N_1331,N_1329);
nand U1495 (N_1495,N_1368,N_1326);
or U1496 (N_1496,N_1389,N_1302);
nor U1497 (N_1497,N_1384,N_1302);
xnor U1498 (N_1498,N_1369,N_1357);
and U1499 (N_1499,N_1367,N_1302);
nor U1500 (N_1500,N_1414,N_1478);
nor U1501 (N_1501,N_1405,N_1424);
and U1502 (N_1502,N_1441,N_1467);
nor U1503 (N_1503,N_1495,N_1415);
nor U1504 (N_1504,N_1432,N_1488);
and U1505 (N_1505,N_1491,N_1460);
nor U1506 (N_1506,N_1442,N_1476);
or U1507 (N_1507,N_1492,N_1401);
nand U1508 (N_1508,N_1430,N_1485);
and U1509 (N_1509,N_1434,N_1449);
or U1510 (N_1510,N_1443,N_1472);
nand U1511 (N_1511,N_1407,N_1493);
and U1512 (N_1512,N_1487,N_1484);
or U1513 (N_1513,N_1450,N_1439);
and U1514 (N_1514,N_1466,N_1409);
or U1515 (N_1515,N_1416,N_1490);
nand U1516 (N_1516,N_1497,N_1486);
nor U1517 (N_1517,N_1436,N_1413);
or U1518 (N_1518,N_1422,N_1479);
and U1519 (N_1519,N_1408,N_1453);
nor U1520 (N_1520,N_1406,N_1404);
nand U1521 (N_1521,N_1471,N_1456);
nor U1522 (N_1522,N_1400,N_1428);
xor U1523 (N_1523,N_1482,N_1440);
or U1524 (N_1524,N_1403,N_1447);
or U1525 (N_1525,N_1423,N_1483);
nor U1526 (N_1526,N_1410,N_1480);
nand U1527 (N_1527,N_1455,N_1438);
nor U1528 (N_1528,N_1435,N_1429);
nand U1529 (N_1529,N_1468,N_1445);
nor U1530 (N_1530,N_1402,N_1411);
or U1531 (N_1531,N_1459,N_1464);
or U1532 (N_1532,N_1474,N_1454);
xnor U1533 (N_1533,N_1425,N_1431);
xnor U1534 (N_1534,N_1457,N_1452);
and U1535 (N_1535,N_1470,N_1469);
nand U1536 (N_1536,N_1433,N_1458);
nor U1537 (N_1537,N_1412,N_1451);
and U1538 (N_1538,N_1481,N_1499);
or U1539 (N_1539,N_1421,N_1420);
nor U1540 (N_1540,N_1417,N_1463);
nor U1541 (N_1541,N_1462,N_1494);
nor U1542 (N_1542,N_1489,N_1448);
nand U1543 (N_1543,N_1444,N_1418);
or U1544 (N_1544,N_1446,N_1437);
or U1545 (N_1545,N_1461,N_1465);
and U1546 (N_1546,N_1419,N_1475);
or U1547 (N_1547,N_1427,N_1473);
and U1548 (N_1548,N_1426,N_1477);
or U1549 (N_1549,N_1498,N_1496);
or U1550 (N_1550,N_1483,N_1418);
and U1551 (N_1551,N_1458,N_1465);
nand U1552 (N_1552,N_1490,N_1438);
nor U1553 (N_1553,N_1477,N_1454);
nand U1554 (N_1554,N_1495,N_1467);
nor U1555 (N_1555,N_1409,N_1445);
and U1556 (N_1556,N_1418,N_1470);
or U1557 (N_1557,N_1432,N_1460);
nand U1558 (N_1558,N_1438,N_1403);
or U1559 (N_1559,N_1445,N_1406);
nor U1560 (N_1560,N_1454,N_1402);
or U1561 (N_1561,N_1470,N_1407);
and U1562 (N_1562,N_1465,N_1478);
or U1563 (N_1563,N_1402,N_1400);
xor U1564 (N_1564,N_1429,N_1499);
nor U1565 (N_1565,N_1418,N_1405);
nor U1566 (N_1566,N_1480,N_1488);
and U1567 (N_1567,N_1403,N_1488);
nand U1568 (N_1568,N_1416,N_1415);
nand U1569 (N_1569,N_1403,N_1426);
xnor U1570 (N_1570,N_1433,N_1429);
nand U1571 (N_1571,N_1447,N_1468);
nor U1572 (N_1572,N_1458,N_1415);
nor U1573 (N_1573,N_1485,N_1477);
nor U1574 (N_1574,N_1466,N_1496);
or U1575 (N_1575,N_1447,N_1488);
nand U1576 (N_1576,N_1456,N_1422);
nor U1577 (N_1577,N_1411,N_1408);
nor U1578 (N_1578,N_1432,N_1470);
and U1579 (N_1579,N_1405,N_1448);
nor U1580 (N_1580,N_1430,N_1468);
nor U1581 (N_1581,N_1479,N_1440);
or U1582 (N_1582,N_1460,N_1454);
or U1583 (N_1583,N_1456,N_1423);
nor U1584 (N_1584,N_1495,N_1480);
or U1585 (N_1585,N_1451,N_1470);
or U1586 (N_1586,N_1475,N_1445);
and U1587 (N_1587,N_1447,N_1411);
or U1588 (N_1588,N_1487,N_1407);
and U1589 (N_1589,N_1476,N_1477);
nand U1590 (N_1590,N_1440,N_1443);
or U1591 (N_1591,N_1443,N_1463);
and U1592 (N_1592,N_1421,N_1488);
or U1593 (N_1593,N_1498,N_1435);
or U1594 (N_1594,N_1489,N_1441);
or U1595 (N_1595,N_1408,N_1437);
nand U1596 (N_1596,N_1448,N_1401);
and U1597 (N_1597,N_1475,N_1466);
nand U1598 (N_1598,N_1400,N_1419);
and U1599 (N_1599,N_1459,N_1403);
and U1600 (N_1600,N_1518,N_1582);
nand U1601 (N_1601,N_1566,N_1553);
nor U1602 (N_1602,N_1550,N_1590);
nor U1603 (N_1603,N_1502,N_1538);
or U1604 (N_1604,N_1520,N_1576);
nor U1605 (N_1605,N_1512,N_1571);
nand U1606 (N_1606,N_1595,N_1569);
xnor U1607 (N_1607,N_1504,N_1547);
nand U1608 (N_1608,N_1565,N_1568);
or U1609 (N_1609,N_1555,N_1556);
or U1610 (N_1610,N_1549,N_1545);
and U1611 (N_1611,N_1527,N_1581);
nor U1612 (N_1612,N_1531,N_1597);
or U1613 (N_1613,N_1583,N_1560);
nand U1614 (N_1614,N_1523,N_1505);
and U1615 (N_1615,N_1535,N_1509);
and U1616 (N_1616,N_1567,N_1537);
nand U1617 (N_1617,N_1596,N_1536);
nor U1618 (N_1618,N_1559,N_1511);
nor U1619 (N_1619,N_1570,N_1586);
nand U1620 (N_1620,N_1580,N_1521);
or U1621 (N_1621,N_1574,N_1539);
or U1622 (N_1622,N_1554,N_1564);
or U1623 (N_1623,N_1516,N_1577);
or U1624 (N_1624,N_1525,N_1593);
nand U1625 (N_1625,N_1587,N_1529);
or U1626 (N_1626,N_1585,N_1513);
and U1627 (N_1627,N_1507,N_1552);
and U1628 (N_1628,N_1517,N_1526);
and U1629 (N_1629,N_1515,N_1543);
or U1630 (N_1630,N_1501,N_1551);
nand U1631 (N_1631,N_1589,N_1510);
nand U1632 (N_1632,N_1592,N_1598);
or U1633 (N_1633,N_1563,N_1579);
or U1634 (N_1634,N_1528,N_1540);
or U1635 (N_1635,N_1544,N_1524);
and U1636 (N_1636,N_1519,N_1561);
nor U1637 (N_1637,N_1573,N_1594);
and U1638 (N_1638,N_1530,N_1533);
nor U1639 (N_1639,N_1532,N_1534);
nand U1640 (N_1640,N_1588,N_1558);
nor U1641 (N_1641,N_1503,N_1548);
and U1642 (N_1642,N_1591,N_1546);
and U1643 (N_1643,N_1542,N_1562);
nand U1644 (N_1644,N_1578,N_1514);
nor U1645 (N_1645,N_1522,N_1508);
nor U1646 (N_1646,N_1506,N_1541);
or U1647 (N_1647,N_1599,N_1500);
and U1648 (N_1648,N_1572,N_1575);
nor U1649 (N_1649,N_1557,N_1584);
nand U1650 (N_1650,N_1593,N_1532);
nor U1651 (N_1651,N_1568,N_1517);
nor U1652 (N_1652,N_1557,N_1531);
and U1653 (N_1653,N_1532,N_1515);
nand U1654 (N_1654,N_1513,N_1520);
or U1655 (N_1655,N_1521,N_1539);
xnor U1656 (N_1656,N_1533,N_1512);
and U1657 (N_1657,N_1574,N_1512);
nor U1658 (N_1658,N_1538,N_1504);
nand U1659 (N_1659,N_1568,N_1577);
nand U1660 (N_1660,N_1506,N_1547);
nor U1661 (N_1661,N_1520,N_1566);
nor U1662 (N_1662,N_1514,N_1568);
nand U1663 (N_1663,N_1552,N_1542);
nand U1664 (N_1664,N_1594,N_1599);
nor U1665 (N_1665,N_1597,N_1573);
nor U1666 (N_1666,N_1508,N_1550);
nor U1667 (N_1667,N_1539,N_1579);
and U1668 (N_1668,N_1595,N_1525);
nand U1669 (N_1669,N_1542,N_1587);
nor U1670 (N_1670,N_1521,N_1586);
nor U1671 (N_1671,N_1541,N_1546);
nand U1672 (N_1672,N_1540,N_1510);
and U1673 (N_1673,N_1523,N_1515);
xnor U1674 (N_1674,N_1529,N_1500);
xor U1675 (N_1675,N_1595,N_1553);
or U1676 (N_1676,N_1534,N_1598);
nand U1677 (N_1677,N_1527,N_1573);
or U1678 (N_1678,N_1547,N_1578);
or U1679 (N_1679,N_1566,N_1556);
and U1680 (N_1680,N_1589,N_1593);
nor U1681 (N_1681,N_1514,N_1549);
and U1682 (N_1682,N_1507,N_1575);
or U1683 (N_1683,N_1533,N_1522);
or U1684 (N_1684,N_1563,N_1516);
nand U1685 (N_1685,N_1582,N_1514);
or U1686 (N_1686,N_1590,N_1559);
and U1687 (N_1687,N_1584,N_1565);
and U1688 (N_1688,N_1591,N_1584);
or U1689 (N_1689,N_1525,N_1575);
nor U1690 (N_1690,N_1581,N_1516);
nand U1691 (N_1691,N_1534,N_1572);
and U1692 (N_1692,N_1560,N_1586);
or U1693 (N_1693,N_1526,N_1502);
and U1694 (N_1694,N_1555,N_1525);
or U1695 (N_1695,N_1502,N_1575);
or U1696 (N_1696,N_1527,N_1571);
nor U1697 (N_1697,N_1592,N_1518);
nand U1698 (N_1698,N_1548,N_1529);
nand U1699 (N_1699,N_1566,N_1528);
nand U1700 (N_1700,N_1681,N_1692);
nand U1701 (N_1701,N_1645,N_1695);
nand U1702 (N_1702,N_1667,N_1654);
nor U1703 (N_1703,N_1661,N_1636);
and U1704 (N_1704,N_1683,N_1641);
and U1705 (N_1705,N_1634,N_1638);
or U1706 (N_1706,N_1647,N_1626);
or U1707 (N_1707,N_1656,N_1699);
nand U1708 (N_1708,N_1682,N_1614);
nand U1709 (N_1709,N_1602,N_1663);
nand U1710 (N_1710,N_1622,N_1694);
nand U1711 (N_1711,N_1617,N_1619);
and U1712 (N_1712,N_1616,N_1662);
nand U1713 (N_1713,N_1643,N_1693);
and U1714 (N_1714,N_1675,N_1684);
nand U1715 (N_1715,N_1676,N_1665);
and U1716 (N_1716,N_1608,N_1642);
nand U1717 (N_1717,N_1666,N_1632);
nand U1718 (N_1718,N_1603,N_1659);
or U1719 (N_1719,N_1615,N_1657);
nand U1720 (N_1720,N_1621,N_1673);
nand U1721 (N_1721,N_1697,N_1685);
nor U1722 (N_1722,N_1677,N_1637);
or U1723 (N_1723,N_1670,N_1686);
and U1724 (N_1724,N_1606,N_1628);
nand U1725 (N_1725,N_1668,N_1652);
and U1726 (N_1726,N_1650,N_1610);
or U1727 (N_1727,N_1680,N_1674);
nand U1728 (N_1728,N_1607,N_1627);
or U1729 (N_1729,N_1671,N_1669);
or U1730 (N_1730,N_1644,N_1688);
or U1731 (N_1731,N_1605,N_1629);
or U1732 (N_1732,N_1658,N_1620);
and U1733 (N_1733,N_1651,N_1612);
nand U1734 (N_1734,N_1649,N_1648);
and U1735 (N_1735,N_1633,N_1639);
nor U1736 (N_1736,N_1687,N_1631);
or U1737 (N_1737,N_1664,N_1678);
nand U1738 (N_1738,N_1672,N_1689);
and U1739 (N_1739,N_1609,N_1698);
nand U1740 (N_1740,N_1601,N_1640);
nand U1741 (N_1741,N_1679,N_1624);
nand U1742 (N_1742,N_1604,N_1691);
nor U1743 (N_1743,N_1646,N_1635);
and U1744 (N_1744,N_1613,N_1625);
nand U1745 (N_1745,N_1660,N_1653);
and U1746 (N_1746,N_1611,N_1630);
nor U1747 (N_1747,N_1618,N_1690);
or U1748 (N_1748,N_1696,N_1655);
nor U1749 (N_1749,N_1623,N_1600);
or U1750 (N_1750,N_1656,N_1685);
nor U1751 (N_1751,N_1688,N_1638);
or U1752 (N_1752,N_1691,N_1661);
nor U1753 (N_1753,N_1636,N_1678);
nor U1754 (N_1754,N_1629,N_1627);
and U1755 (N_1755,N_1606,N_1633);
and U1756 (N_1756,N_1658,N_1680);
nand U1757 (N_1757,N_1651,N_1660);
and U1758 (N_1758,N_1688,N_1604);
nand U1759 (N_1759,N_1669,N_1641);
nor U1760 (N_1760,N_1602,N_1621);
and U1761 (N_1761,N_1653,N_1623);
or U1762 (N_1762,N_1617,N_1641);
xor U1763 (N_1763,N_1658,N_1647);
and U1764 (N_1764,N_1651,N_1669);
xnor U1765 (N_1765,N_1689,N_1666);
or U1766 (N_1766,N_1620,N_1645);
nand U1767 (N_1767,N_1699,N_1615);
nand U1768 (N_1768,N_1677,N_1626);
or U1769 (N_1769,N_1631,N_1693);
nor U1770 (N_1770,N_1679,N_1660);
or U1771 (N_1771,N_1646,N_1677);
or U1772 (N_1772,N_1685,N_1624);
nor U1773 (N_1773,N_1623,N_1628);
nor U1774 (N_1774,N_1623,N_1687);
or U1775 (N_1775,N_1614,N_1653);
or U1776 (N_1776,N_1667,N_1635);
and U1777 (N_1777,N_1689,N_1658);
nor U1778 (N_1778,N_1641,N_1692);
or U1779 (N_1779,N_1649,N_1685);
or U1780 (N_1780,N_1670,N_1620);
nor U1781 (N_1781,N_1673,N_1686);
nor U1782 (N_1782,N_1624,N_1664);
and U1783 (N_1783,N_1601,N_1609);
or U1784 (N_1784,N_1615,N_1633);
nand U1785 (N_1785,N_1625,N_1624);
and U1786 (N_1786,N_1654,N_1630);
nand U1787 (N_1787,N_1604,N_1680);
nor U1788 (N_1788,N_1625,N_1660);
nand U1789 (N_1789,N_1669,N_1683);
and U1790 (N_1790,N_1611,N_1636);
or U1791 (N_1791,N_1680,N_1683);
nor U1792 (N_1792,N_1680,N_1644);
nor U1793 (N_1793,N_1667,N_1636);
nor U1794 (N_1794,N_1624,N_1601);
or U1795 (N_1795,N_1600,N_1681);
and U1796 (N_1796,N_1675,N_1607);
nor U1797 (N_1797,N_1673,N_1637);
and U1798 (N_1798,N_1609,N_1696);
nand U1799 (N_1799,N_1641,N_1614);
and U1800 (N_1800,N_1767,N_1703);
and U1801 (N_1801,N_1792,N_1763);
nor U1802 (N_1802,N_1790,N_1742);
nand U1803 (N_1803,N_1772,N_1770);
nor U1804 (N_1804,N_1777,N_1714);
nor U1805 (N_1805,N_1721,N_1724);
nor U1806 (N_1806,N_1756,N_1716);
nand U1807 (N_1807,N_1715,N_1762);
and U1808 (N_1808,N_1737,N_1751);
nand U1809 (N_1809,N_1768,N_1754);
or U1810 (N_1810,N_1723,N_1732);
nor U1811 (N_1811,N_1752,N_1705);
and U1812 (N_1812,N_1774,N_1776);
or U1813 (N_1813,N_1734,N_1782);
and U1814 (N_1814,N_1780,N_1725);
or U1815 (N_1815,N_1797,N_1735);
nand U1816 (N_1816,N_1799,N_1733);
nor U1817 (N_1817,N_1758,N_1798);
and U1818 (N_1818,N_1793,N_1736);
nor U1819 (N_1819,N_1761,N_1729);
nor U1820 (N_1820,N_1726,N_1718);
nand U1821 (N_1821,N_1730,N_1786);
nor U1822 (N_1822,N_1745,N_1738);
and U1823 (N_1823,N_1746,N_1765);
xor U1824 (N_1824,N_1781,N_1712);
nor U1825 (N_1825,N_1787,N_1704);
nor U1826 (N_1826,N_1743,N_1709);
or U1827 (N_1827,N_1708,N_1740);
nand U1828 (N_1828,N_1784,N_1747);
nand U1829 (N_1829,N_1702,N_1741);
and U1830 (N_1830,N_1722,N_1711);
nor U1831 (N_1831,N_1789,N_1731);
nand U1832 (N_1832,N_1706,N_1755);
nand U1833 (N_1833,N_1783,N_1778);
or U1834 (N_1834,N_1707,N_1771);
nand U1835 (N_1835,N_1779,N_1748);
or U1836 (N_1836,N_1749,N_1794);
nand U1837 (N_1837,N_1717,N_1750);
nor U1838 (N_1838,N_1720,N_1710);
nor U1839 (N_1839,N_1700,N_1775);
or U1840 (N_1840,N_1753,N_1760);
or U1841 (N_1841,N_1728,N_1773);
and U1842 (N_1842,N_1788,N_1739);
nand U1843 (N_1843,N_1785,N_1759);
nand U1844 (N_1844,N_1719,N_1796);
nand U1845 (N_1845,N_1757,N_1727);
nand U1846 (N_1846,N_1766,N_1795);
and U1847 (N_1847,N_1744,N_1713);
and U1848 (N_1848,N_1701,N_1769);
nand U1849 (N_1849,N_1791,N_1764);
nand U1850 (N_1850,N_1749,N_1797);
and U1851 (N_1851,N_1744,N_1754);
nand U1852 (N_1852,N_1723,N_1747);
nor U1853 (N_1853,N_1728,N_1725);
or U1854 (N_1854,N_1759,N_1730);
and U1855 (N_1855,N_1775,N_1747);
and U1856 (N_1856,N_1795,N_1720);
or U1857 (N_1857,N_1793,N_1741);
or U1858 (N_1858,N_1768,N_1713);
nor U1859 (N_1859,N_1776,N_1707);
nor U1860 (N_1860,N_1767,N_1774);
nor U1861 (N_1861,N_1779,N_1708);
nand U1862 (N_1862,N_1779,N_1763);
or U1863 (N_1863,N_1783,N_1743);
nor U1864 (N_1864,N_1743,N_1784);
nand U1865 (N_1865,N_1762,N_1727);
nand U1866 (N_1866,N_1757,N_1720);
nand U1867 (N_1867,N_1700,N_1743);
or U1868 (N_1868,N_1736,N_1713);
nor U1869 (N_1869,N_1757,N_1709);
nand U1870 (N_1870,N_1744,N_1720);
or U1871 (N_1871,N_1728,N_1750);
nand U1872 (N_1872,N_1771,N_1767);
and U1873 (N_1873,N_1728,N_1769);
nor U1874 (N_1874,N_1723,N_1771);
or U1875 (N_1875,N_1763,N_1723);
or U1876 (N_1876,N_1717,N_1798);
and U1877 (N_1877,N_1736,N_1782);
nand U1878 (N_1878,N_1770,N_1709);
nand U1879 (N_1879,N_1749,N_1792);
and U1880 (N_1880,N_1753,N_1702);
and U1881 (N_1881,N_1710,N_1731);
nand U1882 (N_1882,N_1779,N_1768);
nand U1883 (N_1883,N_1715,N_1767);
and U1884 (N_1884,N_1710,N_1745);
nand U1885 (N_1885,N_1747,N_1791);
and U1886 (N_1886,N_1719,N_1774);
nand U1887 (N_1887,N_1763,N_1719);
or U1888 (N_1888,N_1779,N_1715);
nand U1889 (N_1889,N_1773,N_1727);
and U1890 (N_1890,N_1709,N_1771);
nand U1891 (N_1891,N_1703,N_1704);
nand U1892 (N_1892,N_1726,N_1727);
or U1893 (N_1893,N_1741,N_1757);
or U1894 (N_1894,N_1744,N_1723);
nand U1895 (N_1895,N_1789,N_1766);
or U1896 (N_1896,N_1787,N_1721);
or U1897 (N_1897,N_1783,N_1775);
nor U1898 (N_1898,N_1779,N_1727);
nor U1899 (N_1899,N_1705,N_1708);
or U1900 (N_1900,N_1894,N_1845);
and U1901 (N_1901,N_1827,N_1899);
or U1902 (N_1902,N_1864,N_1858);
or U1903 (N_1903,N_1849,N_1842);
nand U1904 (N_1904,N_1891,N_1896);
nor U1905 (N_1905,N_1875,N_1847);
or U1906 (N_1906,N_1834,N_1881);
and U1907 (N_1907,N_1812,N_1857);
and U1908 (N_1908,N_1823,N_1862);
or U1909 (N_1909,N_1853,N_1822);
nand U1910 (N_1910,N_1868,N_1839);
nand U1911 (N_1911,N_1872,N_1860);
nor U1912 (N_1912,N_1819,N_1811);
and U1913 (N_1913,N_1826,N_1892);
xor U1914 (N_1914,N_1884,N_1882);
or U1915 (N_1915,N_1841,N_1825);
and U1916 (N_1916,N_1888,N_1846);
nor U1917 (N_1917,N_1824,N_1898);
or U1918 (N_1918,N_1877,N_1856);
nand U1919 (N_1919,N_1805,N_1889);
and U1920 (N_1920,N_1802,N_1800);
nor U1921 (N_1921,N_1818,N_1865);
and U1922 (N_1922,N_1890,N_1821);
nor U1923 (N_1923,N_1828,N_1843);
and U1924 (N_1924,N_1829,N_1832);
and U1925 (N_1925,N_1873,N_1861);
xnor U1926 (N_1926,N_1895,N_1874);
nor U1927 (N_1927,N_1867,N_1880);
and U1928 (N_1928,N_1831,N_1808);
and U1929 (N_1929,N_1803,N_1876);
nor U1930 (N_1930,N_1893,N_1835);
and U1931 (N_1931,N_1859,N_1850);
and U1932 (N_1932,N_1883,N_1852);
nor U1933 (N_1933,N_1886,N_1837);
or U1934 (N_1934,N_1810,N_1830);
nor U1935 (N_1935,N_1897,N_1833);
nand U1936 (N_1936,N_1885,N_1866);
or U1937 (N_1937,N_1870,N_1836);
and U1938 (N_1938,N_1838,N_1871);
and U1939 (N_1939,N_1855,N_1806);
nor U1940 (N_1940,N_1844,N_1807);
nand U1941 (N_1941,N_1854,N_1804);
nand U1942 (N_1942,N_1820,N_1863);
nand U1943 (N_1943,N_1813,N_1815);
nor U1944 (N_1944,N_1801,N_1809);
and U1945 (N_1945,N_1878,N_1816);
and U1946 (N_1946,N_1840,N_1817);
nand U1947 (N_1947,N_1887,N_1879);
and U1948 (N_1948,N_1848,N_1851);
or U1949 (N_1949,N_1814,N_1869);
nand U1950 (N_1950,N_1889,N_1863);
nor U1951 (N_1951,N_1837,N_1821);
or U1952 (N_1952,N_1830,N_1825);
nor U1953 (N_1953,N_1842,N_1808);
nor U1954 (N_1954,N_1834,N_1843);
nand U1955 (N_1955,N_1877,N_1881);
or U1956 (N_1956,N_1821,N_1874);
nand U1957 (N_1957,N_1887,N_1848);
and U1958 (N_1958,N_1833,N_1819);
or U1959 (N_1959,N_1821,N_1886);
and U1960 (N_1960,N_1880,N_1809);
nor U1961 (N_1961,N_1800,N_1806);
nor U1962 (N_1962,N_1877,N_1880);
nor U1963 (N_1963,N_1807,N_1850);
or U1964 (N_1964,N_1810,N_1870);
nor U1965 (N_1965,N_1830,N_1850);
nor U1966 (N_1966,N_1813,N_1869);
or U1967 (N_1967,N_1823,N_1806);
nor U1968 (N_1968,N_1828,N_1878);
or U1969 (N_1969,N_1811,N_1802);
and U1970 (N_1970,N_1841,N_1813);
and U1971 (N_1971,N_1873,N_1804);
nand U1972 (N_1972,N_1854,N_1851);
and U1973 (N_1973,N_1800,N_1845);
nand U1974 (N_1974,N_1882,N_1847);
or U1975 (N_1975,N_1885,N_1897);
xor U1976 (N_1976,N_1885,N_1840);
or U1977 (N_1977,N_1869,N_1895);
or U1978 (N_1978,N_1869,N_1825);
nor U1979 (N_1979,N_1879,N_1876);
and U1980 (N_1980,N_1811,N_1861);
and U1981 (N_1981,N_1827,N_1817);
or U1982 (N_1982,N_1840,N_1852);
and U1983 (N_1983,N_1845,N_1898);
or U1984 (N_1984,N_1829,N_1886);
nor U1985 (N_1985,N_1867,N_1878);
nor U1986 (N_1986,N_1886,N_1882);
and U1987 (N_1987,N_1803,N_1817);
and U1988 (N_1988,N_1876,N_1871);
or U1989 (N_1989,N_1887,N_1834);
nand U1990 (N_1990,N_1860,N_1856);
and U1991 (N_1991,N_1836,N_1894);
nor U1992 (N_1992,N_1845,N_1805);
nand U1993 (N_1993,N_1841,N_1880);
nand U1994 (N_1994,N_1863,N_1802);
nor U1995 (N_1995,N_1894,N_1899);
and U1996 (N_1996,N_1857,N_1868);
or U1997 (N_1997,N_1884,N_1803);
xnor U1998 (N_1998,N_1861,N_1856);
nor U1999 (N_1999,N_1881,N_1835);
and U2000 (N_2000,N_1905,N_1978);
nor U2001 (N_2001,N_1962,N_1999);
or U2002 (N_2002,N_1946,N_1912);
nand U2003 (N_2003,N_1914,N_1901);
and U2004 (N_2004,N_1929,N_1983);
nor U2005 (N_2005,N_1910,N_1959);
xnor U2006 (N_2006,N_1992,N_1967);
nor U2007 (N_2007,N_1957,N_1994);
nor U2008 (N_2008,N_1906,N_1924);
or U2009 (N_2009,N_1956,N_1926);
or U2010 (N_2010,N_1904,N_1961);
and U2011 (N_2011,N_1908,N_1987);
nor U2012 (N_2012,N_1968,N_1921);
or U2013 (N_2013,N_1973,N_1995);
or U2014 (N_2014,N_1951,N_1955);
nor U2015 (N_2015,N_1988,N_1937);
and U2016 (N_2016,N_1981,N_1942);
nor U2017 (N_2017,N_1970,N_1943);
nor U2018 (N_2018,N_1979,N_1931);
nand U2019 (N_2019,N_1960,N_1939);
or U2020 (N_2020,N_1933,N_1984);
and U2021 (N_2021,N_1945,N_1935);
or U2022 (N_2022,N_1928,N_1936);
or U2023 (N_2023,N_1900,N_1907);
nand U2024 (N_2024,N_1954,N_1938);
nor U2025 (N_2025,N_1982,N_1974);
and U2026 (N_2026,N_1997,N_1913);
nand U2027 (N_2027,N_1911,N_1985);
and U2028 (N_2028,N_1948,N_1953);
nand U2029 (N_2029,N_1918,N_1991);
nor U2030 (N_2030,N_1917,N_1927);
and U2031 (N_2031,N_1972,N_1964);
and U2032 (N_2032,N_1941,N_1952);
nand U2033 (N_2033,N_1950,N_1958);
and U2034 (N_2034,N_1977,N_1980);
nand U2035 (N_2035,N_1922,N_1949);
and U2036 (N_2036,N_1903,N_1969);
and U2037 (N_2037,N_1925,N_1919);
or U2038 (N_2038,N_1993,N_1916);
and U2039 (N_2039,N_1971,N_1966);
or U2040 (N_2040,N_1998,N_1976);
nor U2041 (N_2041,N_1934,N_1909);
nor U2042 (N_2042,N_1932,N_1915);
nand U2043 (N_2043,N_1940,N_1989);
and U2044 (N_2044,N_1947,N_1996);
and U2045 (N_2045,N_1902,N_1975);
xor U2046 (N_2046,N_1963,N_1923);
or U2047 (N_2047,N_1944,N_1920);
or U2048 (N_2048,N_1986,N_1930);
and U2049 (N_2049,N_1990,N_1965);
nand U2050 (N_2050,N_1995,N_1961);
nand U2051 (N_2051,N_1951,N_1968);
nor U2052 (N_2052,N_1979,N_1924);
and U2053 (N_2053,N_1904,N_1952);
nor U2054 (N_2054,N_1929,N_1951);
nor U2055 (N_2055,N_1931,N_1935);
xnor U2056 (N_2056,N_1958,N_1972);
and U2057 (N_2057,N_1974,N_1936);
nand U2058 (N_2058,N_1912,N_1915);
or U2059 (N_2059,N_1903,N_1984);
or U2060 (N_2060,N_1980,N_1900);
nor U2061 (N_2061,N_1946,N_1919);
or U2062 (N_2062,N_1947,N_1908);
and U2063 (N_2063,N_1973,N_1971);
or U2064 (N_2064,N_1914,N_1981);
or U2065 (N_2065,N_1925,N_1999);
or U2066 (N_2066,N_1978,N_1913);
xnor U2067 (N_2067,N_1965,N_1992);
or U2068 (N_2068,N_1955,N_1934);
nand U2069 (N_2069,N_1925,N_1997);
xnor U2070 (N_2070,N_1932,N_1970);
nand U2071 (N_2071,N_1954,N_1901);
nor U2072 (N_2072,N_1975,N_1959);
and U2073 (N_2073,N_1971,N_1913);
or U2074 (N_2074,N_1943,N_1992);
or U2075 (N_2075,N_1911,N_1965);
nor U2076 (N_2076,N_1958,N_1991);
or U2077 (N_2077,N_1959,N_1925);
nor U2078 (N_2078,N_1909,N_1925);
nor U2079 (N_2079,N_1947,N_1961);
nand U2080 (N_2080,N_1954,N_1912);
nand U2081 (N_2081,N_1944,N_1916);
nand U2082 (N_2082,N_1921,N_1977);
nand U2083 (N_2083,N_1983,N_1946);
or U2084 (N_2084,N_1914,N_1912);
and U2085 (N_2085,N_1919,N_1928);
nand U2086 (N_2086,N_1991,N_1967);
or U2087 (N_2087,N_1909,N_1976);
and U2088 (N_2088,N_1969,N_1929);
nand U2089 (N_2089,N_1920,N_1965);
or U2090 (N_2090,N_1943,N_1901);
nor U2091 (N_2091,N_1946,N_1935);
nand U2092 (N_2092,N_1950,N_1970);
and U2093 (N_2093,N_1910,N_1978);
or U2094 (N_2094,N_1961,N_1982);
nor U2095 (N_2095,N_1979,N_1954);
and U2096 (N_2096,N_1967,N_1947);
or U2097 (N_2097,N_1938,N_1992);
and U2098 (N_2098,N_1987,N_1933);
and U2099 (N_2099,N_1902,N_1954);
or U2100 (N_2100,N_2004,N_2002);
nor U2101 (N_2101,N_2061,N_2028);
xor U2102 (N_2102,N_2020,N_2090);
and U2103 (N_2103,N_2094,N_2066);
nand U2104 (N_2104,N_2006,N_2069);
and U2105 (N_2105,N_2067,N_2049);
xor U2106 (N_2106,N_2077,N_2011);
xnor U2107 (N_2107,N_2060,N_2050);
nor U2108 (N_2108,N_2082,N_2087);
nor U2109 (N_2109,N_2068,N_2019);
and U2110 (N_2110,N_2072,N_2025);
or U2111 (N_2111,N_2036,N_2086);
or U2112 (N_2112,N_2035,N_2057);
or U2113 (N_2113,N_2051,N_2097);
nand U2114 (N_2114,N_2039,N_2034);
or U2115 (N_2115,N_2024,N_2045);
nor U2116 (N_2116,N_2033,N_2063);
or U2117 (N_2117,N_2021,N_2040);
nor U2118 (N_2118,N_2075,N_2073);
or U2119 (N_2119,N_2014,N_2044);
nor U2120 (N_2120,N_2016,N_2026);
or U2121 (N_2121,N_2078,N_2053);
nand U2122 (N_2122,N_2056,N_2093);
xor U2123 (N_2123,N_2052,N_2047);
nor U2124 (N_2124,N_2048,N_2076);
or U2125 (N_2125,N_2001,N_2084);
nand U2126 (N_2126,N_2059,N_2030);
and U2127 (N_2127,N_2027,N_2032);
and U2128 (N_2128,N_2088,N_2018);
or U2129 (N_2129,N_2010,N_2009);
nor U2130 (N_2130,N_2065,N_2042);
and U2131 (N_2131,N_2043,N_2085);
nor U2132 (N_2132,N_2080,N_2079);
and U2133 (N_2133,N_2064,N_2007);
or U2134 (N_2134,N_2071,N_2031);
and U2135 (N_2135,N_2041,N_2038);
nor U2136 (N_2136,N_2091,N_2005);
and U2137 (N_2137,N_2029,N_2015);
nand U2138 (N_2138,N_2058,N_2092);
and U2139 (N_2139,N_2055,N_2054);
or U2140 (N_2140,N_2023,N_2062);
nand U2141 (N_2141,N_2089,N_2081);
and U2142 (N_2142,N_2098,N_2083);
nand U2143 (N_2143,N_2013,N_2095);
nor U2144 (N_2144,N_2017,N_2074);
nor U2145 (N_2145,N_2099,N_2012);
or U2146 (N_2146,N_2037,N_2096);
or U2147 (N_2147,N_2022,N_2003);
or U2148 (N_2148,N_2008,N_2070);
or U2149 (N_2149,N_2046,N_2000);
and U2150 (N_2150,N_2018,N_2075);
nand U2151 (N_2151,N_2079,N_2077);
nand U2152 (N_2152,N_2082,N_2090);
nand U2153 (N_2153,N_2088,N_2095);
nor U2154 (N_2154,N_2014,N_2092);
xnor U2155 (N_2155,N_2072,N_2008);
nand U2156 (N_2156,N_2091,N_2011);
or U2157 (N_2157,N_2082,N_2069);
or U2158 (N_2158,N_2009,N_2027);
and U2159 (N_2159,N_2007,N_2041);
nor U2160 (N_2160,N_2083,N_2015);
or U2161 (N_2161,N_2018,N_2093);
nor U2162 (N_2162,N_2020,N_2068);
and U2163 (N_2163,N_2099,N_2093);
xor U2164 (N_2164,N_2090,N_2098);
nor U2165 (N_2165,N_2096,N_2006);
nor U2166 (N_2166,N_2054,N_2080);
or U2167 (N_2167,N_2012,N_2066);
or U2168 (N_2168,N_2058,N_2020);
and U2169 (N_2169,N_2086,N_2076);
nor U2170 (N_2170,N_2088,N_2084);
nor U2171 (N_2171,N_2002,N_2074);
or U2172 (N_2172,N_2011,N_2093);
or U2173 (N_2173,N_2053,N_2020);
and U2174 (N_2174,N_2002,N_2077);
nand U2175 (N_2175,N_2072,N_2033);
or U2176 (N_2176,N_2004,N_2057);
or U2177 (N_2177,N_2054,N_2052);
nand U2178 (N_2178,N_2036,N_2009);
and U2179 (N_2179,N_2038,N_2013);
nand U2180 (N_2180,N_2097,N_2079);
or U2181 (N_2181,N_2049,N_2020);
and U2182 (N_2182,N_2067,N_2092);
and U2183 (N_2183,N_2093,N_2061);
or U2184 (N_2184,N_2061,N_2025);
and U2185 (N_2185,N_2040,N_2082);
nor U2186 (N_2186,N_2026,N_2036);
and U2187 (N_2187,N_2074,N_2098);
and U2188 (N_2188,N_2095,N_2005);
or U2189 (N_2189,N_2063,N_2088);
or U2190 (N_2190,N_2070,N_2053);
and U2191 (N_2191,N_2074,N_2058);
and U2192 (N_2192,N_2035,N_2043);
and U2193 (N_2193,N_2031,N_2043);
or U2194 (N_2194,N_2017,N_2057);
and U2195 (N_2195,N_2017,N_2008);
nand U2196 (N_2196,N_2012,N_2037);
and U2197 (N_2197,N_2041,N_2048);
nand U2198 (N_2198,N_2005,N_2040);
nand U2199 (N_2199,N_2058,N_2001);
nand U2200 (N_2200,N_2124,N_2133);
nor U2201 (N_2201,N_2130,N_2178);
or U2202 (N_2202,N_2171,N_2114);
and U2203 (N_2203,N_2148,N_2182);
nor U2204 (N_2204,N_2179,N_2128);
nor U2205 (N_2205,N_2165,N_2192);
and U2206 (N_2206,N_2155,N_2120);
or U2207 (N_2207,N_2140,N_2118);
and U2208 (N_2208,N_2109,N_2123);
and U2209 (N_2209,N_2199,N_2195);
nand U2210 (N_2210,N_2145,N_2159);
xor U2211 (N_2211,N_2173,N_2164);
or U2212 (N_2212,N_2105,N_2136);
or U2213 (N_2213,N_2119,N_2143);
and U2214 (N_2214,N_2186,N_2141);
or U2215 (N_2215,N_2154,N_2193);
nand U2216 (N_2216,N_2142,N_2103);
or U2217 (N_2217,N_2163,N_2139);
and U2218 (N_2218,N_2116,N_2174);
nand U2219 (N_2219,N_2167,N_2168);
and U2220 (N_2220,N_2188,N_2162);
and U2221 (N_2221,N_2187,N_2100);
and U2222 (N_2222,N_2108,N_2161);
and U2223 (N_2223,N_2115,N_2104);
nor U2224 (N_2224,N_2102,N_2197);
and U2225 (N_2225,N_2153,N_2134);
nand U2226 (N_2226,N_2107,N_2122);
nand U2227 (N_2227,N_2156,N_2149);
and U2228 (N_2228,N_2157,N_2177);
and U2229 (N_2229,N_2183,N_2169);
and U2230 (N_2230,N_2121,N_2144);
nor U2231 (N_2231,N_2194,N_2117);
nor U2232 (N_2232,N_2126,N_2166);
nand U2233 (N_2233,N_2176,N_2180);
nand U2234 (N_2234,N_2196,N_2172);
nand U2235 (N_2235,N_2181,N_2131);
and U2236 (N_2236,N_2112,N_2151);
or U2237 (N_2237,N_2190,N_2191);
or U2238 (N_2238,N_2175,N_2138);
nand U2239 (N_2239,N_2152,N_2129);
nand U2240 (N_2240,N_2160,N_2170);
and U2241 (N_2241,N_2106,N_2132);
nor U2242 (N_2242,N_2111,N_2185);
and U2243 (N_2243,N_2135,N_2125);
nand U2244 (N_2244,N_2150,N_2137);
or U2245 (N_2245,N_2146,N_2113);
or U2246 (N_2246,N_2101,N_2158);
nor U2247 (N_2247,N_2184,N_2189);
or U2248 (N_2248,N_2110,N_2147);
nor U2249 (N_2249,N_2198,N_2127);
and U2250 (N_2250,N_2105,N_2161);
nor U2251 (N_2251,N_2182,N_2167);
nor U2252 (N_2252,N_2133,N_2163);
and U2253 (N_2253,N_2171,N_2119);
nor U2254 (N_2254,N_2183,N_2176);
or U2255 (N_2255,N_2139,N_2141);
nand U2256 (N_2256,N_2140,N_2144);
or U2257 (N_2257,N_2106,N_2149);
nor U2258 (N_2258,N_2141,N_2100);
and U2259 (N_2259,N_2137,N_2129);
nand U2260 (N_2260,N_2104,N_2138);
nand U2261 (N_2261,N_2190,N_2113);
or U2262 (N_2262,N_2178,N_2167);
nor U2263 (N_2263,N_2130,N_2106);
or U2264 (N_2264,N_2121,N_2154);
or U2265 (N_2265,N_2146,N_2143);
nand U2266 (N_2266,N_2158,N_2122);
nor U2267 (N_2267,N_2132,N_2181);
nor U2268 (N_2268,N_2154,N_2119);
nand U2269 (N_2269,N_2168,N_2142);
nor U2270 (N_2270,N_2117,N_2101);
and U2271 (N_2271,N_2119,N_2199);
and U2272 (N_2272,N_2194,N_2189);
nor U2273 (N_2273,N_2162,N_2172);
nor U2274 (N_2274,N_2129,N_2126);
nand U2275 (N_2275,N_2193,N_2164);
nand U2276 (N_2276,N_2181,N_2116);
or U2277 (N_2277,N_2196,N_2141);
and U2278 (N_2278,N_2183,N_2108);
nor U2279 (N_2279,N_2151,N_2130);
and U2280 (N_2280,N_2153,N_2168);
nand U2281 (N_2281,N_2107,N_2148);
nand U2282 (N_2282,N_2102,N_2196);
nor U2283 (N_2283,N_2115,N_2191);
nand U2284 (N_2284,N_2178,N_2199);
nand U2285 (N_2285,N_2175,N_2133);
or U2286 (N_2286,N_2145,N_2113);
and U2287 (N_2287,N_2143,N_2100);
nor U2288 (N_2288,N_2132,N_2104);
nand U2289 (N_2289,N_2142,N_2177);
nand U2290 (N_2290,N_2131,N_2122);
or U2291 (N_2291,N_2167,N_2151);
or U2292 (N_2292,N_2122,N_2151);
nand U2293 (N_2293,N_2101,N_2194);
or U2294 (N_2294,N_2136,N_2118);
and U2295 (N_2295,N_2194,N_2145);
nand U2296 (N_2296,N_2141,N_2111);
or U2297 (N_2297,N_2103,N_2198);
or U2298 (N_2298,N_2170,N_2177);
or U2299 (N_2299,N_2187,N_2156);
nand U2300 (N_2300,N_2290,N_2285);
nor U2301 (N_2301,N_2231,N_2269);
nand U2302 (N_2302,N_2281,N_2230);
or U2303 (N_2303,N_2213,N_2255);
nand U2304 (N_2304,N_2256,N_2241);
nor U2305 (N_2305,N_2235,N_2244);
xnor U2306 (N_2306,N_2206,N_2216);
nor U2307 (N_2307,N_2232,N_2280);
nor U2308 (N_2308,N_2267,N_2211);
nand U2309 (N_2309,N_2200,N_2299);
nor U2310 (N_2310,N_2243,N_2298);
nand U2311 (N_2311,N_2275,N_2260);
nand U2312 (N_2312,N_2252,N_2291);
and U2313 (N_2313,N_2242,N_2233);
nor U2314 (N_2314,N_2268,N_2228);
or U2315 (N_2315,N_2248,N_2274);
and U2316 (N_2316,N_2214,N_2217);
nand U2317 (N_2317,N_2223,N_2236);
nand U2318 (N_2318,N_2276,N_2258);
nand U2319 (N_2319,N_2208,N_2239);
nand U2320 (N_2320,N_2238,N_2222);
and U2321 (N_2321,N_2286,N_2212);
nor U2322 (N_2322,N_2283,N_2261);
nor U2323 (N_2323,N_2263,N_2294);
and U2324 (N_2324,N_2254,N_2292);
nand U2325 (N_2325,N_2250,N_2272);
nor U2326 (N_2326,N_2278,N_2224);
and U2327 (N_2327,N_2229,N_2265);
nor U2328 (N_2328,N_2240,N_2259);
nand U2329 (N_2329,N_2273,N_2295);
and U2330 (N_2330,N_2221,N_2271);
nand U2331 (N_2331,N_2234,N_2207);
xnor U2332 (N_2332,N_2202,N_2296);
nand U2333 (N_2333,N_2287,N_2288);
and U2334 (N_2334,N_2253,N_2204);
or U2335 (N_2335,N_2282,N_2249);
nand U2336 (N_2336,N_2277,N_2218);
nor U2337 (N_2337,N_2209,N_2264);
and U2338 (N_2338,N_2245,N_2270);
nor U2339 (N_2339,N_2237,N_2289);
xnor U2340 (N_2340,N_2262,N_2257);
nor U2341 (N_2341,N_2220,N_2266);
or U2342 (N_2342,N_2205,N_2201);
nor U2343 (N_2343,N_2251,N_2284);
and U2344 (N_2344,N_2246,N_2219);
and U2345 (N_2345,N_2279,N_2227);
nand U2346 (N_2346,N_2226,N_2297);
and U2347 (N_2347,N_2293,N_2203);
nand U2348 (N_2348,N_2215,N_2247);
xnor U2349 (N_2349,N_2225,N_2210);
xor U2350 (N_2350,N_2242,N_2264);
or U2351 (N_2351,N_2264,N_2247);
nand U2352 (N_2352,N_2204,N_2264);
nor U2353 (N_2353,N_2237,N_2272);
nand U2354 (N_2354,N_2299,N_2240);
and U2355 (N_2355,N_2296,N_2273);
nand U2356 (N_2356,N_2244,N_2253);
nor U2357 (N_2357,N_2207,N_2284);
nand U2358 (N_2358,N_2266,N_2260);
nand U2359 (N_2359,N_2213,N_2264);
and U2360 (N_2360,N_2242,N_2207);
and U2361 (N_2361,N_2261,N_2213);
nand U2362 (N_2362,N_2293,N_2210);
or U2363 (N_2363,N_2244,N_2221);
and U2364 (N_2364,N_2225,N_2230);
or U2365 (N_2365,N_2249,N_2257);
or U2366 (N_2366,N_2215,N_2238);
or U2367 (N_2367,N_2243,N_2224);
and U2368 (N_2368,N_2295,N_2221);
nor U2369 (N_2369,N_2288,N_2207);
or U2370 (N_2370,N_2260,N_2200);
nand U2371 (N_2371,N_2253,N_2212);
nand U2372 (N_2372,N_2268,N_2288);
and U2373 (N_2373,N_2268,N_2255);
or U2374 (N_2374,N_2253,N_2211);
nand U2375 (N_2375,N_2203,N_2250);
nor U2376 (N_2376,N_2261,N_2228);
and U2377 (N_2377,N_2250,N_2204);
nand U2378 (N_2378,N_2254,N_2245);
or U2379 (N_2379,N_2202,N_2209);
and U2380 (N_2380,N_2268,N_2267);
xor U2381 (N_2381,N_2293,N_2291);
and U2382 (N_2382,N_2286,N_2270);
nand U2383 (N_2383,N_2269,N_2297);
and U2384 (N_2384,N_2216,N_2267);
or U2385 (N_2385,N_2233,N_2201);
nand U2386 (N_2386,N_2256,N_2292);
and U2387 (N_2387,N_2273,N_2204);
xnor U2388 (N_2388,N_2233,N_2290);
nand U2389 (N_2389,N_2296,N_2226);
nand U2390 (N_2390,N_2263,N_2228);
nand U2391 (N_2391,N_2268,N_2250);
nand U2392 (N_2392,N_2227,N_2278);
or U2393 (N_2393,N_2262,N_2247);
and U2394 (N_2394,N_2276,N_2264);
nand U2395 (N_2395,N_2263,N_2271);
and U2396 (N_2396,N_2299,N_2232);
nand U2397 (N_2397,N_2225,N_2267);
or U2398 (N_2398,N_2275,N_2253);
nor U2399 (N_2399,N_2236,N_2294);
or U2400 (N_2400,N_2341,N_2313);
and U2401 (N_2401,N_2325,N_2302);
and U2402 (N_2402,N_2374,N_2335);
or U2403 (N_2403,N_2354,N_2346);
or U2404 (N_2404,N_2307,N_2360);
nand U2405 (N_2405,N_2326,N_2363);
nor U2406 (N_2406,N_2324,N_2333);
and U2407 (N_2407,N_2339,N_2394);
and U2408 (N_2408,N_2305,N_2382);
nand U2409 (N_2409,N_2304,N_2381);
and U2410 (N_2410,N_2301,N_2372);
nor U2411 (N_2411,N_2336,N_2308);
nand U2412 (N_2412,N_2379,N_2389);
or U2413 (N_2413,N_2340,N_2334);
nand U2414 (N_2414,N_2321,N_2384);
nor U2415 (N_2415,N_2392,N_2393);
or U2416 (N_2416,N_2356,N_2391);
or U2417 (N_2417,N_2370,N_2348);
nor U2418 (N_2418,N_2387,N_2371);
nor U2419 (N_2419,N_2310,N_2303);
nand U2420 (N_2420,N_2352,N_2328);
or U2421 (N_2421,N_2375,N_2314);
and U2422 (N_2422,N_2368,N_2369);
or U2423 (N_2423,N_2380,N_2319);
or U2424 (N_2424,N_2331,N_2342);
and U2425 (N_2425,N_2329,N_2337);
or U2426 (N_2426,N_2353,N_2345);
and U2427 (N_2427,N_2359,N_2358);
and U2428 (N_2428,N_2343,N_2349);
and U2429 (N_2429,N_2362,N_2320);
nand U2430 (N_2430,N_2373,N_2351);
and U2431 (N_2431,N_2383,N_2317);
nor U2432 (N_2432,N_2386,N_2364);
nor U2433 (N_2433,N_2312,N_2395);
nand U2434 (N_2434,N_2396,N_2300);
and U2435 (N_2435,N_2332,N_2388);
or U2436 (N_2436,N_2390,N_2378);
nor U2437 (N_2437,N_2357,N_2376);
nand U2438 (N_2438,N_2316,N_2399);
nand U2439 (N_2439,N_2347,N_2397);
nand U2440 (N_2440,N_2355,N_2318);
or U2441 (N_2441,N_2315,N_2366);
or U2442 (N_2442,N_2323,N_2338);
and U2443 (N_2443,N_2385,N_2330);
nor U2444 (N_2444,N_2327,N_2350);
nand U2445 (N_2445,N_2322,N_2309);
and U2446 (N_2446,N_2311,N_2398);
or U2447 (N_2447,N_2344,N_2377);
or U2448 (N_2448,N_2361,N_2306);
nand U2449 (N_2449,N_2365,N_2367);
nor U2450 (N_2450,N_2353,N_2360);
or U2451 (N_2451,N_2386,N_2318);
and U2452 (N_2452,N_2321,N_2315);
or U2453 (N_2453,N_2379,N_2356);
nor U2454 (N_2454,N_2362,N_2303);
nor U2455 (N_2455,N_2376,N_2366);
nand U2456 (N_2456,N_2356,N_2333);
and U2457 (N_2457,N_2329,N_2342);
nand U2458 (N_2458,N_2370,N_2328);
nand U2459 (N_2459,N_2325,N_2363);
nor U2460 (N_2460,N_2352,N_2366);
nand U2461 (N_2461,N_2301,N_2375);
nor U2462 (N_2462,N_2322,N_2339);
nand U2463 (N_2463,N_2373,N_2358);
nor U2464 (N_2464,N_2367,N_2371);
or U2465 (N_2465,N_2356,N_2362);
and U2466 (N_2466,N_2376,N_2359);
nand U2467 (N_2467,N_2342,N_2338);
or U2468 (N_2468,N_2398,N_2326);
nor U2469 (N_2469,N_2331,N_2339);
nand U2470 (N_2470,N_2339,N_2328);
nand U2471 (N_2471,N_2398,N_2374);
and U2472 (N_2472,N_2360,N_2327);
nor U2473 (N_2473,N_2384,N_2322);
nand U2474 (N_2474,N_2387,N_2370);
or U2475 (N_2475,N_2310,N_2379);
and U2476 (N_2476,N_2317,N_2328);
nor U2477 (N_2477,N_2395,N_2300);
or U2478 (N_2478,N_2378,N_2361);
nor U2479 (N_2479,N_2302,N_2337);
nand U2480 (N_2480,N_2356,N_2392);
nor U2481 (N_2481,N_2321,N_2317);
nor U2482 (N_2482,N_2341,N_2365);
or U2483 (N_2483,N_2396,N_2352);
and U2484 (N_2484,N_2311,N_2373);
xnor U2485 (N_2485,N_2389,N_2347);
nand U2486 (N_2486,N_2335,N_2379);
or U2487 (N_2487,N_2362,N_2300);
xnor U2488 (N_2488,N_2312,N_2383);
nand U2489 (N_2489,N_2358,N_2391);
nand U2490 (N_2490,N_2309,N_2352);
nand U2491 (N_2491,N_2370,N_2380);
and U2492 (N_2492,N_2381,N_2331);
nor U2493 (N_2493,N_2337,N_2307);
nor U2494 (N_2494,N_2356,N_2313);
or U2495 (N_2495,N_2310,N_2312);
and U2496 (N_2496,N_2332,N_2324);
nand U2497 (N_2497,N_2310,N_2306);
or U2498 (N_2498,N_2358,N_2375);
or U2499 (N_2499,N_2304,N_2340);
or U2500 (N_2500,N_2486,N_2484);
or U2501 (N_2501,N_2496,N_2433);
or U2502 (N_2502,N_2456,N_2455);
nand U2503 (N_2503,N_2416,N_2479);
or U2504 (N_2504,N_2467,N_2411);
nand U2505 (N_2505,N_2417,N_2448);
nand U2506 (N_2506,N_2418,N_2498);
nand U2507 (N_2507,N_2443,N_2404);
and U2508 (N_2508,N_2485,N_2410);
nor U2509 (N_2509,N_2490,N_2460);
nor U2510 (N_2510,N_2452,N_2489);
nand U2511 (N_2511,N_2428,N_2429);
nand U2512 (N_2512,N_2413,N_2477);
nand U2513 (N_2513,N_2482,N_2466);
nor U2514 (N_2514,N_2431,N_2474);
nand U2515 (N_2515,N_2459,N_2453);
nand U2516 (N_2516,N_2432,N_2434);
or U2517 (N_2517,N_2425,N_2450);
nand U2518 (N_2518,N_2493,N_2463);
xnor U2519 (N_2519,N_2444,N_2461);
nand U2520 (N_2520,N_2472,N_2478);
and U2521 (N_2521,N_2422,N_2408);
nand U2522 (N_2522,N_2407,N_2458);
or U2523 (N_2523,N_2419,N_2415);
and U2524 (N_2524,N_2491,N_2435);
nor U2525 (N_2525,N_2449,N_2481);
xnor U2526 (N_2526,N_2405,N_2470);
nor U2527 (N_2527,N_2451,N_2442);
nor U2528 (N_2528,N_2462,N_2494);
nor U2529 (N_2529,N_2436,N_2468);
or U2530 (N_2530,N_2471,N_2497);
or U2531 (N_2531,N_2447,N_2464);
nand U2532 (N_2532,N_2480,N_2421);
nor U2533 (N_2533,N_2440,N_2401);
xnor U2534 (N_2534,N_2483,N_2475);
or U2535 (N_2535,N_2409,N_2406);
and U2536 (N_2536,N_2437,N_2402);
or U2537 (N_2537,N_2423,N_2426);
nor U2538 (N_2538,N_2439,N_2441);
or U2539 (N_2539,N_2412,N_2420);
nor U2540 (N_2540,N_2427,N_2445);
nand U2541 (N_2541,N_2492,N_2487);
nand U2542 (N_2542,N_2400,N_2499);
or U2543 (N_2543,N_2446,N_2454);
and U2544 (N_2544,N_2488,N_2403);
and U2545 (N_2545,N_2473,N_2438);
and U2546 (N_2546,N_2495,N_2457);
nor U2547 (N_2547,N_2465,N_2414);
or U2548 (N_2548,N_2469,N_2424);
or U2549 (N_2549,N_2476,N_2430);
nor U2550 (N_2550,N_2403,N_2402);
or U2551 (N_2551,N_2426,N_2416);
and U2552 (N_2552,N_2453,N_2475);
nor U2553 (N_2553,N_2457,N_2434);
nand U2554 (N_2554,N_2422,N_2490);
nor U2555 (N_2555,N_2420,N_2406);
nor U2556 (N_2556,N_2441,N_2453);
or U2557 (N_2557,N_2439,N_2435);
and U2558 (N_2558,N_2437,N_2413);
and U2559 (N_2559,N_2459,N_2464);
and U2560 (N_2560,N_2403,N_2445);
nor U2561 (N_2561,N_2417,N_2456);
or U2562 (N_2562,N_2406,N_2482);
nor U2563 (N_2563,N_2428,N_2412);
nand U2564 (N_2564,N_2453,N_2499);
and U2565 (N_2565,N_2406,N_2456);
nand U2566 (N_2566,N_2464,N_2419);
or U2567 (N_2567,N_2443,N_2492);
nand U2568 (N_2568,N_2416,N_2483);
or U2569 (N_2569,N_2455,N_2498);
nand U2570 (N_2570,N_2488,N_2463);
and U2571 (N_2571,N_2431,N_2486);
nand U2572 (N_2572,N_2468,N_2451);
nand U2573 (N_2573,N_2405,N_2421);
and U2574 (N_2574,N_2450,N_2483);
nand U2575 (N_2575,N_2420,N_2466);
or U2576 (N_2576,N_2467,N_2436);
or U2577 (N_2577,N_2493,N_2423);
nand U2578 (N_2578,N_2400,N_2467);
xor U2579 (N_2579,N_2466,N_2472);
nand U2580 (N_2580,N_2479,N_2406);
nand U2581 (N_2581,N_2479,N_2419);
and U2582 (N_2582,N_2473,N_2457);
and U2583 (N_2583,N_2470,N_2461);
or U2584 (N_2584,N_2466,N_2475);
nand U2585 (N_2585,N_2484,N_2464);
or U2586 (N_2586,N_2427,N_2448);
nor U2587 (N_2587,N_2429,N_2455);
nand U2588 (N_2588,N_2425,N_2429);
and U2589 (N_2589,N_2439,N_2429);
nor U2590 (N_2590,N_2452,N_2447);
nor U2591 (N_2591,N_2409,N_2469);
nor U2592 (N_2592,N_2471,N_2421);
or U2593 (N_2593,N_2444,N_2402);
or U2594 (N_2594,N_2475,N_2497);
xor U2595 (N_2595,N_2426,N_2419);
nand U2596 (N_2596,N_2412,N_2415);
nand U2597 (N_2597,N_2469,N_2474);
and U2598 (N_2598,N_2469,N_2433);
nor U2599 (N_2599,N_2495,N_2463);
nor U2600 (N_2600,N_2543,N_2532);
and U2601 (N_2601,N_2565,N_2537);
xor U2602 (N_2602,N_2551,N_2575);
and U2603 (N_2603,N_2553,N_2526);
nand U2604 (N_2604,N_2523,N_2546);
or U2605 (N_2605,N_2509,N_2573);
xor U2606 (N_2606,N_2529,N_2500);
nand U2607 (N_2607,N_2542,N_2520);
nor U2608 (N_2608,N_2541,N_2550);
nand U2609 (N_2609,N_2510,N_2576);
or U2610 (N_2610,N_2507,N_2534);
and U2611 (N_2611,N_2596,N_2564);
nor U2612 (N_2612,N_2547,N_2567);
nor U2613 (N_2613,N_2533,N_2517);
or U2614 (N_2614,N_2593,N_2518);
nand U2615 (N_2615,N_2548,N_2506);
nand U2616 (N_2616,N_2561,N_2535);
and U2617 (N_2617,N_2552,N_2597);
or U2618 (N_2618,N_2577,N_2522);
and U2619 (N_2619,N_2594,N_2559);
nand U2620 (N_2620,N_2581,N_2571);
and U2621 (N_2621,N_2589,N_2568);
nor U2622 (N_2622,N_2572,N_2562);
nand U2623 (N_2623,N_2515,N_2578);
and U2624 (N_2624,N_2554,N_2519);
and U2625 (N_2625,N_2528,N_2527);
nor U2626 (N_2626,N_2514,N_2560);
or U2627 (N_2627,N_2538,N_2563);
nor U2628 (N_2628,N_2516,N_2549);
and U2629 (N_2629,N_2574,N_2504);
and U2630 (N_2630,N_2595,N_2524);
nand U2631 (N_2631,N_2590,N_2598);
and U2632 (N_2632,N_2502,N_2505);
or U2633 (N_2633,N_2513,N_2569);
nand U2634 (N_2634,N_2503,N_2566);
nor U2635 (N_2635,N_2540,N_2591);
nand U2636 (N_2636,N_2599,N_2592);
nand U2637 (N_2637,N_2587,N_2588);
nor U2638 (N_2638,N_2544,N_2580);
nand U2639 (N_2639,N_2558,N_2521);
nand U2640 (N_2640,N_2511,N_2584);
or U2641 (N_2641,N_2531,N_2586);
nand U2642 (N_2642,N_2512,N_2539);
nor U2643 (N_2643,N_2555,N_2530);
and U2644 (N_2644,N_2557,N_2570);
nand U2645 (N_2645,N_2585,N_2536);
or U2646 (N_2646,N_2501,N_2545);
and U2647 (N_2647,N_2579,N_2582);
nor U2648 (N_2648,N_2583,N_2556);
or U2649 (N_2649,N_2525,N_2508);
nand U2650 (N_2650,N_2552,N_2513);
and U2651 (N_2651,N_2551,N_2525);
nand U2652 (N_2652,N_2542,N_2510);
and U2653 (N_2653,N_2530,N_2583);
or U2654 (N_2654,N_2580,N_2599);
or U2655 (N_2655,N_2531,N_2514);
and U2656 (N_2656,N_2597,N_2511);
or U2657 (N_2657,N_2520,N_2556);
and U2658 (N_2658,N_2500,N_2532);
or U2659 (N_2659,N_2564,N_2578);
or U2660 (N_2660,N_2552,N_2594);
and U2661 (N_2661,N_2507,N_2558);
nand U2662 (N_2662,N_2568,N_2594);
and U2663 (N_2663,N_2513,N_2561);
or U2664 (N_2664,N_2570,N_2519);
nand U2665 (N_2665,N_2585,N_2593);
nor U2666 (N_2666,N_2512,N_2506);
and U2667 (N_2667,N_2534,N_2502);
nand U2668 (N_2668,N_2574,N_2533);
and U2669 (N_2669,N_2555,N_2524);
nor U2670 (N_2670,N_2505,N_2548);
nand U2671 (N_2671,N_2514,N_2519);
or U2672 (N_2672,N_2524,N_2588);
nand U2673 (N_2673,N_2567,N_2582);
nor U2674 (N_2674,N_2597,N_2584);
nand U2675 (N_2675,N_2548,N_2553);
nor U2676 (N_2676,N_2588,N_2598);
nor U2677 (N_2677,N_2580,N_2595);
nor U2678 (N_2678,N_2575,N_2519);
and U2679 (N_2679,N_2555,N_2520);
nor U2680 (N_2680,N_2549,N_2529);
nor U2681 (N_2681,N_2508,N_2545);
or U2682 (N_2682,N_2519,N_2506);
or U2683 (N_2683,N_2561,N_2596);
or U2684 (N_2684,N_2533,N_2576);
or U2685 (N_2685,N_2598,N_2553);
nor U2686 (N_2686,N_2536,N_2557);
and U2687 (N_2687,N_2585,N_2524);
and U2688 (N_2688,N_2591,N_2541);
nand U2689 (N_2689,N_2567,N_2541);
and U2690 (N_2690,N_2524,N_2542);
and U2691 (N_2691,N_2542,N_2587);
and U2692 (N_2692,N_2549,N_2548);
or U2693 (N_2693,N_2547,N_2554);
or U2694 (N_2694,N_2577,N_2532);
nand U2695 (N_2695,N_2583,N_2582);
nand U2696 (N_2696,N_2513,N_2598);
xnor U2697 (N_2697,N_2548,N_2577);
nor U2698 (N_2698,N_2542,N_2568);
nor U2699 (N_2699,N_2516,N_2594);
and U2700 (N_2700,N_2648,N_2654);
nor U2701 (N_2701,N_2627,N_2678);
nor U2702 (N_2702,N_2659,N_2624);
nand U2703 (N_2703,N_2690,N_2653);
and U2704 (N_2704,N_2675,N_2639);
or U2705 (N_2705,N_2650,N_2612);
or U2706 (N_2706,N_2658,N_2600);
and U2707 (N_2707,N_2643,N_2683);
xor U2708 (N_2708,N_2603,N_2623);
nand U2709 (N_2709,N_2674,N_2632);
and U2710 (N_2710,N_2604,N_2630);
nand U2711 (N_2711,N_2693,N_2652);
and U2712 (N_2712,N_2685,N_2694);
nand U2713 (N_2713,N_2609,N_2673);
nand U2714 (N_2714,N_2616,N_2640);
and U2715 (N_2715,N_2619,N_2698);
nand U2716 (N_2716,N_2666,N_2672);
or U2717 (N_2717,N_2667,N_2677);
or U2718 (N_2718,N_2638,N_2684);
nor U2719 (N_2719,N_2642,N_2605);
nor U2720 (N_2720,N_2634,N_2607);
nand U2721 (N_2721,N_2651,N_2611);
nand U2722 (N_2722,N_2622,N_2669);
nor U2723 (N_2723,N_2615,N_2621);
or U2724 (N_2724,N_2601,N_2664);
nor U2725 (N_2725,N_2608,N_2657);
nor U2726 (N_2726,N_2617,N_2695);
and U2727 (N_2727,N_2633,N_2671);
or U2728 (N_2728,N_2625,N_2626);
or U2729 (N_2729,N_2655,N_2649);
or U2730 (N_2730,N_2692,N_2699);
nand U2731 (N_2731,N_2637,N_2628);
nor U2732 (N_2732,N_2656,N_2613);
nand U2733 (N_2733,N_2697,N_2662);
nor U2734 (N_2734,N_2660,N_2689);
nand U2735 (N_2735,N_2635,N_2686);
and U2736 (N_2736,N_2647,N_2618);
and U2737 (N_2737,N_2670,N_2661);
nand U2738 (N_2738,N_2606,N_2696);
or U2739 (N_2739,N_2644,N_2668);
and U2740 (N_2740,N_2679,N_2676);
nand U2741 (N_2741,N_2665,N_2663);
nand U2742 (N_2742,N_2691,N_2602);
nand U2743 (N_2743,N_2645,N_2620);
or U2744 (N_2744,N_2610,N_2681);
nor U2745 (N_2745,N_2629,N_2680);
or U2746 (N_2746,N_2687,N_2631);
and U2747 (N_2747,N_2646,N_2641);
nand U2748 (N_2748,N_2682,N_2688);
or U2749 (N_2749,N_2614,N_2636);
and U2750 (N_2750,N_2668,N_2611);
or U2751 (N_2751,N_2629,N_2657);
nor U2752 (N_2752,N_2695,N_2651);
nand U2753 (N_2753,N_2677,N_2679);
or U2754 (N_2754,N_2637,N_2688);
or U2755 (N_2755,N_2642,N_2607);
nand U2756 (N_2756,N_2678,N_2603);
nor U2757 (N_2757,N_2609,N_2649);
and U2758 (N_2758,N_2655,N_2677);
nand U2759 (N_2759,N_2638,N_2639);
or U2760 (N_2760,N_2618,N_2662);
or U2761 (N_2761,N_2605,N_2626);
nand U2762 (N_2762,N_2619,N_2642);
and U2763 (N_2763,N_2621,N_2602);
nor U2764 (N_2764,N_2690,N_2612);
nand U2765 (N_2765,N_2664,N_2671);
nand U2766 (N_2766,N_2604,N_2657);
and U2767 (N_2767,N_2632,N_2615);
and U2768 (N_2768,N_2684,N_2632);
nand U2769 (N_2769,N_2601,N_2617);
nand U2770 (N_2770,N_2658,N_2686);
nand U2771 (N_2771,N_2660,N_2676);
or U2772 (N_2772,N_2695,N_2615);
nor U2773 (N_2773,N_2697,N_2693);
and U2774 (N_2774,N_2670,N_2641);
nand U2775 (N_2775,N_2686,N_2693);
and U2776 (N_2776,N_2638,N_2627);
or U2777 (N_2777,N_2630,N_2672);
nor U2778 (N_2778,N_2665,N_2667);
nor U2779 (N_2779,N_2695,N_2674);
and U2780 (N_2780,N_2607,N_2653);
nand U2781 (N_2781,N_2675,N_2641);
nand U2782 (N_2782,N_2668,N_2664);
nand U2783 (N_2783,N_2688,N_2685);
or U2784 (N_2784,N_2677,N_2698);
nand U2785 (N_2785,N_2689,N_2603);
and U2786 (N_2786,N_2693,N_2671);
nor U2787 (N_2787,N_2642,N_2600);
nor U2788 (N_2788,N_2668,N_2610);
or U2789 (N_2789,N_2644,N_2645);
nor U2790 (N_2790,N_2620,N_2623);
and U2791 (N_2791,N_2602,N_2618);
and U2792 (N_2792,N_2605,N_2609);
nor U2793 (N_2793,N_2671,N_2641);
or U2794 (N_2794,N_2661,N_2646);
nor U2795 (N_2795,N_2624,N_2671);
and U2796 (N_2796,N_2625,N_2664);
and U2797 (N_2797,N_2683,N_2693);
or U2798 (N_2798,N_2689,N_2656);
nor U2799 (N_2799,N_2666,N_2695);
and U2800 (N_2800,N_2718,N_2774);
nor U2801 (N_2801,N_2723,N_2700);
nor U2802 (N_2802,N_2754,N_2726);
nand U2803 (N_2803,N_2734,N_2710);
nand U2804 (N_2804,N_2779,N_2764);
nor U2805 (N_2805,N_2738,N_2746);
or U2806 (N_2806,N_2798,N_2749);
xnor U2807 (N_2807,N_2793,N_2770);
and U2808 (N_2808,N_2791,N_2755);
or U2809 (N_2809,N_2788,N_2728);
nand U2810 (N_2810,N_2796,N_2717);
or U2811 (N_2811,N_2705,N_2730);
nor U2812 (N_2812,N_2794,N_2785);
and U2813 (N_2813,N_2761,N_2767);
or U2814 (N_2814,N_2773,N_2744);
nand U2815 (N_2815,N_2766,N_2762);
or U2816 (N_2816,N_2789,N_2702);
or U2817 (N_2817,N_2772,N_2748);
nand U2818 (N_2818,N_2757,N_2714);
nor U2819 (N_2819,N_2708,N_2765);
or U2820 (N_2820,N_2769,N_2732);
or U2821 (N_2821,N_2733,N_2706);
nand U2822 (N_2822,N_2784,N_2747);
nand U2823 (N_2823,N_2753,N_2790);
nand U2824 (N_2824,N_2752,N_2721);
nor U2825 (N_2825,N_2735,N_2743);
and U2826 (N_2826,N_2778,N_2781);
and U2827 (N_2827,N_2729,N_2756);
or U2828 (N_2828,N_2709,N_2725);
or U2829 (N_2829,N_2750,N_2715);
nand U2830 (N_2830,N_2713,N_2740);
nand U2831 (N_2831,N_2742,N_2768);
and U2832 (N_2832,N_2799,N_2736);
or U2833 (N_2833,N_2795,N_2775);
or U2834 (N_2834,N_2712,N_2759);
or U2835 (N_2835,N_2760,N_2792);
nand U2836 (N_2836,N_2727,N_2701);
xnor U2837 (N_2837,N_2724,N_2780);
and U2838 (N_2838,N_2720,N_2745);
nand U2839 (N_2839,N_2786,N_2758);
nand U2840 (N_2840,N_2797,N_2739);
nand U2841 (N_2841,N_2777,N_2741);
or U2842 (N_2842,N_2737,N_2751);
or U2843 (N_2843,N_2782,N_2704);
or U2844 (N_2844,N_2722,N_2783);
or U2845 (N_2845,N_2776,N_2707);
and U2846 (N_2846,N_2771,N_2719);
nand U2847 (N_2847,N_2731,N_2763);
nor U2848 (N_2848,N_2716,N_2711);
and U2849 (N_2849,N_2703,N_2787);
or U2850 (N_2850,N_2767,N_2738);
or U2851 (N_2851,N_2761,N_2748);
nand U2852 (N_2852,N_2766,N_2720);
nand U2853 (N_2853,N_2756,N_2781);
and U2854 (N_2854,N_2764,N_2724);
nor U2855 (N_2855,N_2745,N_2787);
nand U2856 (N_2856,N_2769,N_2712);
xnor U2857 (N_2857,N_2736,N_2731);
or U2858 (N_2858,N_2776,N_2792);
nand U2859 (N_2859,N_2799,N_2795);
and U2860 (N_2860,N_2757,N_2712);
or U2861 (N_2861,N_2792,N_2766);
and U2862 (N_2862,N_2725,N_2703);
nor U2863 (N_2863,N_2706,N_2787);
nor U2864 (N_2864,N_2732,N_2781);
or U2865 (N_2865,N_2726,N_2723);
or U2866 (N_2866,N_2722,N_2771);
nor U2867 (N_2867,N_2755,N_2760);
nor U2868 (N_2868,N_2794,N_2744);
nand U2869 (N_2869,N_2746,N_2781);
or U2870 (N_2870,N_2724,N_2751);
and U2871 (N_2871,N_2706,N_2776);
and U2872 (N_2872,N_2789,N_2755);
or U2873 (N_2873,N_2745,N_2738);
or U2874 (N_2874,N_2760,N_2756);
nor U2875 (N_2875,N_2754,N_2735);
xnor U2876 (N_2876,N_2794,N_2791);
nand U2877 (N_2877,N_2776,N_2775);
or U2878 (N_2878,N_2759,N_2790);
nand U2879 (N_2879,N_2721,N_2768);
nand U2880 (N_2880,N_2710,N_2792);
and U2881 (N_2881,N_2783,N_2726);
and U2882 (N_2882,N_2787,N_2785);
or U2883 (N_2883,N_2749,N_2764);
xor U2884 (N_2884,N_2739,N_2727);
nor U2885 (N_2885,N_2723,N_2764);
nand U2886 (N_2886,N_2750,N_2777);
xor U2887 (N_2887,N_2792,N_2708);
nand U2888 (N_2888,N_2751,N_2734);
nand U2889 (N_2889,N_2726,N_2719);
nor U2890 (N_2890,N_2750,N_2740);
or U2891 (N_2891,N_2746,N_2745);
nor U2892 (N_2892,N_2741,N_2761);
nor U2893 (N_2893,N_2712,N_2762);
or U2894 (N_2894,N_2770,N_2742);
and U2895 (N_2895,N_2719,N_2731);
or U2896 (N_2896,N_2782,N_2711);
or U2897 (N_2897,N_2788,N_2794);
and U2898 (N_2898,N_2778,N_2772);
nand U2899 (N_2899,N_2790,N_2731);
or U2900 (N_2900,N_2800,N_2890);
nor U2901 (N_2901,N_2851,N_2835);
nand U2902 (N_2902,N_2867,N_2814);
nand U2903 (N_2903,N_2807,N_2804);
nor U2904 (N_2904,N_2857,N_2819);
nor U2905 (N_2905,N_2854,N_2816);
nand U2906 (N_2906,N_2873,N_2843);
or U2907 (N_2907,N_2844,N_2841);
nand U2908 (N_2908,N_2808,N_2853);
and U2909 (N_2909,N_2826,N_2831);
nand U2910 (N_2910,N_2875,N_2809);
nand U2911 (N_2911,N_2837,N_2812);
nand U2912 (N_2912,N_2861,N_2885);
and U2913 (N_2913,N_2888,N_2863);
nor U2914 (N_2914,N_2882,N_2891);
and U2915 (N_2915,N_2876,N_2847);
and U2916 (N_2916,N_2834,N_2805);
and U2917 (N_2917,N_2833,N_2838);
nand U2918 (N_2918,N_2855,N_2846);
and U2919 (N_2919,N_2842,N_2889);
or U2920 (N_2920,N_2828,N_2899);
or U2921 (N_2921,N_2860,N_2818);
nor U2922 (N_2922,N_2822,N_2856);
nand U2923 (N_2923,N_2825,N_2836);
nand U2924 (N_2924,N_2803,N_2892);
nand U2925 (N_2925,N_2852,N_2824);
nor U2926 (N_2926,N_2806,N_2859);
or U2927 (N_2927,N_2832,N_2894);
or U2928 (N_2928,N_2865,N_2895);
nand U2929 (N_2929,N_2858,N_2874);
nand U2930 (N_2930,N_2827,N_2887);
and U2931 (N_2931,N_2813,N_2811);
nand U2932 (N_2932,N_2864,N_2877);
nand U2933 (N_2933,N_2848,N_2810);
xnor U2934 (N_2934,N_2886,N_2872);
nor U2935 (N_2935,N_2840,N_2821);
nor U2936 (N_2936,N_2878,N_2815);
nor U2937 (N_2937,N_2883,N_2850);
nor U2938 (N_2938,N_2823,N_2839);
and U2939 (N_2939,N_2869,N_2820);
and U2940 (N_2940,N_2849,N_2862);
and U2941 (N_2941,N_2897,N_2829);
and U2942 (N_2942,N_2893,N_2870);
or U2943 (N_2943,N_2871,N_2845);
or U2944 (N_2944,N_2898,N_2817);
or U2945 (N_2945,N_2866,N_2884);
nand U2946 (N_2946,N_2801,N_2880);
nand U2947 (N_2947,N_2879,N_2868);
or U2948 (N_2948,N_2881,N_2802);
and U2949 (N_2949,N_2896,N_2830);
and U2950 (N_2950,N_2815,N_2818);
nor U2951 (N_2951,N_2843,N_2864);
nand U2952 (N_2952,N_2850,N_2800);
nor U2953 (N_2953,N_2818,N_2888);
and U2954 (N_2954,N_2871,N_2820);
nor U2955 (N_2955,N_2864,N_2881);
nand U2956 (N_2956,N_2873,N_2886);
nor U2957 (N_2957,N_2855,N_2869);
nand U2958 (N_2958,N_2854,N_2858);
and U2959 (N_2959,N_2804,N_2893);
and U2960 (N_2960,N_2856,N_2847);
nand U2961 (N_2961,N_2805,N_2815);
nor U2962 (N_2962,N_2834,N_2866);
nand U2963 (N_2963,N_2899,N_2848);
or U2964 (N_2964,N_2812,N_2876);
nand U2965 (N_2965,N_2890,N_2826);
and U2966 (N_2966,N_2865,N_2839);
and U2967 (N_2967,N_2808,N_2837);
nor U2968 (N_2968,N_2827,N_2866);
nor U2969 (N_2969,N_2847,N_2854);
or U2970 (N_2970,N_2821,N_2875);
nor U2971 (N_2971,N_2897,N_2818);
or U2972 (N_2972,N_2843,N_2855);
and U2973 (N_2973,N_2821,N_2886);
xnor U2974 (N_2974,N_2885,N_2850);
nand U2975 (N_2975,N_2814,N_2880);
and U2976 (N_2976,N_2879,N_2898);
nand U2977 (N_2977,N_2858,N_2863);
and U2978 (N_2978,N_2848,N_2859);
or U2979 (N_2979,N_2835,N_2862);
or U2980 (N_2980,N_2823,N_2809);
nor U2981 (N_2981,N_2868,N_2800);
or U2982 (N_2982,N_2886,N_2820);
nor U2983 (N_2983,N_2848,N_2847);
nor U2984 (N_2984,N_2838,N_2864);
nor U2985 (N_2985,N_2867,N_2898);
or U2986 (N_2986,N_2887,N_2829);
nand U2987 (N_2987,N_2871,N_2867);
nor U2988 (N_2988,N_2813,N_2845);
nor U2989 (N_2989,N_2814,N_2855);
nor U2990 (N_2990,N_2810,N_2875);
and U2991 (N_2991,N_2872,N_2867);
or U2992 (N_2992,N_2874,N_2827);
and U2993 (N_2993,N_2839,N_2885);
nor U2994 (N_2994,N_2836,N_2813);
and U2995 (N_2995,N_2865,N_2822);
nand U2996 (N_2996,N_2847,N_2842);
nor U2997 (N_2997,N_2882,N_2803);
or U2998 (N_2998,N_2840,N_2893);
nand U2999 (N_2999,N_2838,N_2853);
nand U3000 (N_3000,N_2905,N_2909);
nand U3001 (N_3001,N_2992,N_2942);
nand U3002 (N_3002,N_2951,N_2953);
nand U3003 (N_3003,N_2975,N_2963);
nor U3004 (N_3004,N_2962,N_2924);
nand U3005 (N_3005,N_2900,N_2989);
nor U3006 (N_3006,N_2945,N_2914);
nand U3007 (N_3007,N_2929,N_2908);
or U3008 (N_3008,N_2910,N_2958);
nor U3009 (N_3009,N_2990,N_2932);
or U3010 (N_3010,N_2931,N_2949);
or U3011 (N_3011,N_2980,N_2937);
nor U3012 (N_3012,N_2936,N_2954);
or U3013 (N_3013,N_2997,N_2965);
nor U3014 (N_3014,N_2998,N_2939);
xor U3015 (N_3015,N_2988,N_2981);
nand U3016 (N_3016,N_2933,N_2964);
and U3017 (N_3017,N_2979,N_2977);
nor U3018 (N_3018,N_2946,N_2904);
nor U3019 (N_3019,N_2927,N_2957);
nor U3020 (N_3020,N_2974,N_2906);
nor U3021 (N_3021,N_2920,N_2961);
and U3022 (N_3022,N_2911,N_2968);
and U3023 (N_3023,N_2921,N_2916);
nand U3024 (N_3024,N_2901,N_2996);
nand U3025 (N_3025,N_2983,N_2960);
nand U3026 (N_3026,N_2947,N_2993);
nor U3027 (N_3027,N_2994,N_2918);
nand U3028 (N_3028,N_2925,N_2966);
and U3029 (N_3029,N_2991,N_2978);
and U3030 (N_3030,N_2922,N_2944);
and U3031 (N_3031,N_2986,N_2952);
nor U3032 (N_3032,N_2941,N_2972);
and U3033 (N_3033,N_2955,N_2940);
nand U3034 (N_3034,N_2903,N_2987);
and U3035 (N_3035,N_2928,N_2926);
nand U3036 (N_3036,N_2934,N_2907);
nand U3037 (N_3037,N_2969,N_2985);
nor U3038 (N_3038,N_2935,N_2938);
nor U3039 (N_3039,N_2950,N_2995);
or U3040 (N_3040,N_2923,N_2917);
and U3041 (N_3041,N_2919,N_2915);
nand U3042 (N_3042,N_2943,N_2973);
nand U3043 (N_3043,N_2967,N_2984);
or U3044 (N_3044,N_2902,N_2982);
nor U3045 (N_3045,N_2948,N_2912);
or U3046 (N_3046,N_2971,N_2976);
and U3047 (N_3047,N_2913,N_2970);
and U3048 (N_3048,N_2999,N_2959);
nand U3049 (N_3049,N_2956,N_2930);
nor U3050 (N_3050,N_2931,N_2954);
nand U3051 (N_3051,N_2958,N_2947);
nand U3052 (N_3052,N_2992,N_2991);
nand U3053 (N_3053,N_2944,N_2914);
nor U3054 (N_3054,N_2978,N_2903);
and U3055 (N_3055,N_2940,N_2947);
nor U3056 (N_3056,N_2973,N_2927);
nor U3057 (N_3057,N_2964,N_2941);
or U3058 (N_3058,N_2982,N_2987);
or U3059 (N_3059,N_2994,N_2966);
and U3060 (N_3060,N_2913,N_2944);
or U3061 (N_3061,N_2926,N_2968);
or U3062 (N_3062,N_2927,N_2995);
and U3063 (N_3063,N_2993,N_2966);
nand U3064 (N_3064,N_2931,N_2985);
nor U3065 (N_3065,N_2969,N_2993);
nor U3066 (N_3066,N_2942,N_2983);
nand U3067 (N_3067,N_2916,N_2949);
and U3068 (N_3068,N_2990,N_2986);
and U3069 (N_3069,N_2941,N_2915);
and U3070 (N_3070,N_2972,N_2908);
nand U3071 (N_3071,N_2926,N_2948);
and U3072 (N_3072,N_2972,N_2967);
and U3073 (N_3073,N_2925,N_2955);
nand U3074 (N_3074,N_2947,N_2992);
and U3075 (N_3075,N_2914,N_2941);
nand U3076 (N_3076,N_2930,N_2902);
or U3077 (N_3077,N_2998,N_2938);
or U3078 (N_3078,N_2942,N_2916);
nand U3079 (N_3079,N_2951,N_2906);
nand U3080 (N_3080,N_2950,N_2941);
or U3081 (N_3081,N_2957,N_2993);
and U3082 (N_3082,N_2988,N_2976);
nand U3083 (N_3083,N_2942,N_2910);
nand U3084 (N_3084,N_2919,N_2927);
nand U3085 (N_3085,N_2953,N_2903);
or U3086 (N_3086,N_2983,N_2933);
and U3087 (N_3087,N_2903,N_2940);
nand U3088 (N_3088,N_2931,N_2920);
nor U3089 (N_3089,N_2936,N_2921);
and U3090 (N_3090,N_2907,N_2918);
or U3091 (N_3091,N_2968,N_2963);
and U3092 (N_3092,N_2966,N_2972);
and U3093 (N_3093,N_2981,N_2909);
nor U3094 (N_3094,N_2997,N_2961);
or U3095 (N_3095,N_2917,N_2905);
nand U3096 (N_3096,N_2968,N_2971);
nand U3097 (N_3097,N_2958,N_2988);
nand U3098 (N_3098,N_2913,N_2997);
nand U3099 (N_3099,N_2901,N_2941);
or U3100 (N_3100,N_3080,N_3067);
and U3101 (N_3101,N_3093,N_3009);
or U3102 (N_3102,N_3022,N_3071);
nor U3103 (N_3103,N_3011,N_3076);
or U3104 (N_3104,N_3016,N_3044);
or U3105 (N_3105,N_3063,N_3003);
nor U3106 (N_3106,N_3026,N_3007);
and U3107 (N_3107,N_3052,N_3058);
nor U3108 (N_3108,N_3060,N_3032);
nor U3109 (N_3109,N_3006,N_3087);
or U3110 (N_3110,N_3019,N_3029);
and U3111 (N_3111,N_3061,N_3010);
or U3112 (N_3112,N_3059,N_3089);
nor U3113 (N_3113,N_3085,N_3036);
nor U3114 (N_3114,N_3064,N_3017);
nor U3115 (N_3115,N_3098,N_3086);
or U3116 (N_3116,N_3014,N_3002);
or U3117 (N_3117,N_3088,N_3077);
nor U3118 (N_3118,N_3001,N_3013);
xor U3119 (N_3119,N_3041,N_3096);
nand U3120 (N_3120,N_3099,N_3065);
and U3121 (N_3121,N_3008,N_3043);
and U3122 (N_3122,N_3097,N_3025);
or U3123 (N_3123,N_3005,N_3012);
or U3124 (N_3124,N_3037,N_3049);
and U3125 (N_3125,N_3015,N_3023);
or U3126 (N_3126,N_3082,N_3020);
or U3127 (N_3127,N_3083,N_3040);
nor U3128 (N_3128,N_3074,N_3068);
nand U3129 (N_3129,N_3055,N_3091);
nand U3130 (N_3130,N_3053,N_3039);
or U3131 (N_3131,N_3028,N_3095);
or U3132 (N_3132,N_3024,N_3070);
nor U3133 (N_3133,N_3021,N_3056);
nor U3134 (N_3134,N_3030,N_3066);
nor U3135 (N_3135,N_3033,N_3079);
nand U3136 (N_3136,N_3075,N_3051);
nand U3137 (N_3137,N_3062,N_3034);
or U3138 (N_3138,N_3078,N_3038);
xor U3139 (N_3139,N_3046,N_3031);
and U3140 (N_3140,N_3048,N_3050);
and U3141 (N_3141,N_3072,N_3073);
or U3142 (N_3142,N_3047,N_3094);
nand U3143 (N_3143,N_3018,N_3027);
nand U3144 (N_3144,N_3090,N_3054);
nor U3145 (N_3145,N_3057,N_3000);
and U3146 (N_3146,N_3069,N_3045);
nor U3147 (N_3147,N_3004,N_3081);
nand U3148 (N_3148,N_3092,N_3035);
and U3149 (N_3149,N_3084,N_3042);
and U3150 (N_3150,N_3015,N_3067);
or U3151 (N_3151,N_3053,N_3084);
or U3152 (N_3152,N_3079,N_3057);
or U3153 (N_3153,N_3080,N_3022);
or U3154 (N_3154,N_3020,N_3084);
and U3155 (N_3155,N_3008,N_3075);
nand U3156 (N_3156,N_3014,N_3098);
and U3157 (N_3157,N_3091,N_3014);
and U3158 (N_3158,N_3015,N_3010);
or U3159 (N_3159,N_3052,N_3025);
or U3160 (N_3160,N_3086,N_3095);
nand U3161 (N_3161,N_3003,N_3098);
nor U3162 (N_3162,N_3043,N_3086);
nor U3163 (N_3163,N_3013,N_3058);
and U3164 (N_3164,N_3086,N_3078);
nand U3165 (N_3165,N_3021,N_3053);
and U3166 (N_3166,N_3002,N_3025);
or U3167 (N_3167,N_3074,N_3053);
and U3168 (N_3168,N_3087,N_3096);
nand U3169 (N_3169,N_3084,N_3008);
xnor U3170 (N_3170,N_3025,N_3055);
xor U3171 (N_3171,N_3077,N_3058);
and U3172 (N_3172,N_3030,N_3028);
nor U3173 (N_3173,N_3060,N_3070);
xor U3174 (N_3174,N_3017,N_3052);
nand U3175 (N_3175,N_3015,N_3013);
nand U3176 (N_3176,N_3020,N_3015);
nand U3177 (N_3177,N_3032,N_3047);
nand U3178 (N_3178,N_3082,N_3052);
and U3179 (N_3179,N_3001,N_3096);
and U3180 (N_3180,N_3047,N_3006);
nand U3181 (N_3181,N_3045,N_3099);
and U3182 (N_3182,N_3080,N_3082);
nor U3183 (N_3183,N_3016,N_3049);
and U3184 (N_3184,N_3043,N_3017);
or U3185 (N_3185,N_3096,N_3056);
or U3186 (N_3186,N_3010,N_3081);
nor U3187 (N_3187,N_3019,N_3006);
and U3188 (N_3188,N_3053,N_3059);
nor U3189 (N_3189,N_3082,N_3079);
or U3190 (N_3190,N_3034,N_3042);
and U3191 (N_3191,N_3080,N_3018);
and U3192 (N_3192,N_3098,N_3040);
nor U3193 (N_3193,N_3072,N_3094);
or U3194 (N_3194,N_3031,N_3027);
or U3195 (N_3195,N_3082,N_3003);
and U3196 (N_3196,N_3089,N_3058);
nor U3197 (N_3197,N_3085,N_3019);
or U3198 (N_3198,N_3028,N_3037);
nand U3199 (N_3199,N_3035,N_3067);
and U3200 (N_3200,N_3178,N_3186);
or U3201 (N_3201,N_3156,N_3151);
nand U3202 (N_3202,N_3107,N_3130);
nor U3203 (N_3203,N_3189,N_3140);
or U3204 (N_3204,N_3152,N_3188);
or U3205 (N_3205,N_3101,N_3122);
and U3206 (N_3206,N_3131,N_3191);
and U3207 (N_3207,N_3149,N_3133);
or U3208 (N_3208,N_3163,N_3143);
and U3209 (N_3209,N_3196,N_3134);
nor U3210 (N_3210,N_3177,N_3179);
or U3211 (N_3211,N_3147,N_3146);
and U3212 (N_3212,N_3112,N_3168);
nand U3213 (N_3213,N_3195,N_3117);
or U3214 (N_3214,N_3139,N_3104);
nor U3215 (N_3215,N_3182,N_3118);
nor U3216 (N_3216,N_3170,N_3113);
and U3217 (N_3217,N_3137,N_3169);
nor U3218 (N_3218,N_3172,N_3110);
nand U3219 (N_3219,N_3161,N_3181);
nor U3220 (N_3220,N_3174,N_3100);
nor U3221 (N_3221,N_3160,N_3190);
xor U3222 (N_3222,N_3121,N_3153);
nor U3223 (N_3223,N_3114,N_3184);
nor U3224 (N_3224,N_3197,N_3108);
and U3225 (N_3225,N_3106,N_3119);
nor U3226 (N_3226,N_3175,N_3138);
or U3227 (N_3227,N_3167,N_3194);
nor U3228 (N_3228,N_3105,N_3192);
nand U3229 (N_3229,N_3183,N_3129);
and U3230 (N_3230,N_3115,N_3141);
or U3231 (N_3231,N_3185,N_3159);
and U3232 (N_3232,N_3103,N_3148);
or U3233 (N_3233,N_3155,N_3144);
nor U3234 (N_3234,N_3124,N_3187);
nand U3235 (N_3235,N_3127,N_3171);
xnor U3236 (N_3236,N_3132,N_3198);
and U3237 (N_3237,N_3136,N_3145);
nor U3238 (N_3238,N_3102,N_3166);
and U3239 (N_3239,N_3123,N_3120);
nand U3240 (N_3240,N_3176,N_3126);
nand U3241 (N_3241,N_3180,N_3164);
nor U3242 (N_3242,N_3135,N_3111);
nand U3243 (N_3243,N_3116,N_3193);
nor U3244 (N_3244,N_3109,N_3150);
nand U3245 (N_3245,N_3142,N_3154);
and U3246 (N_3246,N_3165,N_3199);
or U3247 (N_3247,N_3125,N_3158);
nand U3248 (N_3248,N_3162,N_3173);
and U3249 (N_3249,N_3157,N_3128);
and U3250 (N_3250,N_3123,N_3163);
or U3251 (N_3251,N_3114,N_3153);
nand U3252 (N_3252,N_3124,N_3133);
and U3253 (N_3253,N_3176,N_3159);
or U3254 (N_3254,N_3149,N_3103);
and U3255 (N_3255,N_3140,N_3125);
and U3256 (N_3256,N_3155,N_3148);
or U3257 (N_3257,N_3119,N_3156);
and U3258 (N_3258,N_3164,N_3132);
and U3259 (N_3259,N_3143,N_3109);
nor U3260 (N_3260,N_3172,N_3119);
nand U3261 (N_3261,N_3139,N_3190);
or U3262 (N_3262,N_3136,N_3135);
nor U3263 (N_3263,N_3112,N_3103);
nand U3264 (N_3264,N_3125,N_3150);
nor U3265 (N_3265,N_3104,N_3118);
and U3266 (N_3266,N_3131,N_3189);
nand U3267 (N_3267,N_3194,N_3174);
nand U3268 (N_3268,N_3189,N_3129);
or U3269 (N_3269,N_3199,N_3166);
and U3270 (N_3270,N_3110,N_3147);
or U3271 (N_3271,N_3194,N_3147);
or U3272 (N_3272,N_3101,N_3136);
nor U3273 (N_3273,N_3156,N_3106);
and U3274 (N_3274,N_3149,N_3141);
or U3275 (N_3275,N_3150,N_3179);
or U3276 (N_3276,N_3122,N_3108);
nand U3277 (N_3277,N_3144,N_3176);
and U3278 (N_3278,N_3163,N_3148);
nor U3279 (N_3279,N_3167,N_3136);
nand U3280 (N_3280,N_3181,N_3145);
and U3281 (N_3281,N_3196,N_3152);
and U3282 (N_3282,N_3151,N_3124);
or U3283 (N_3283,N_3110,N_3128);
and U3284 (N_3284,N_3197,N_3112);
and U3285 (N_3285,N_3195,N_3155);
nand U3286 (N_3286,N_3196,N_3100);
nor U3287 (N_3287,N_3137,N_3193);
or U3288 (N_3288,N_3171,N_3186);
nand U3289 (N_3289,N_3145,N_3148);
and U3290 (N_3290,N_3197,N_3132);
or U3291 (N_3291,N_3157,N_3171);
and U3292 (N_3292,N_3119,N_3102);
or U3293 (N_3293,N_3141,N_3143);
and U3294 (N_3294,N_3148,N_3142);
and U3295 (N_3295,N_3109,N_3180);
nand U3296 (N_3296,N_3127,N_3169);
and U3297 (N_3297,N_3121,N_3185);
nand U3298 (N_3298,N_3147,N_3111);
nand U3299 (N_3299,N_3100,N_3177);
and U3300 (N_3300,N_3218,N_3217);
nor U3301 (N_3301,N_3256,N_3232);
or U3302 (N_3302,N_3237,N_3276);
and U3303 (N_3303,N_3229,N_3245);
or U3304 (N_3304,N_3213,N_3270);
and U3305 (N_3305,N_3206,N_3277);
nand U3306 (N_3306,N_3240,N_3230);
and U3307 (N_3307,N_3271,N_3211);
nor U3308 (N_3308,N_3269,N_3262);
nand U3309 (N_3309,N_3287,N_3249);
nor U3310 (N_3310,N_3203,N_3288);
nand U3311 (N_3311,N_3285,N_3201);
or U3312 (N_3312,N_3272,N_3281);
and U3313 (N_3313,N_3231,N_3273);
and U3314 (N_3314,N_3208,N_3222);
nand U3315 (N_3315,N_3292,N_3244);
nor U3316 (N_3316,N_3268,N_3242);
or U3317 (N_3317,N_3246,N_3243);
nor U3318 (N_3318,N_3200,N_3226);
nor U3319 (N_3319,N_3223,N_3215);
nand U3320 (N_3320,N_3258,N_3257);
nor U3321 (N_3321,N_3266,N_3250);
or U3322 (N_3322,N_3234,N_3220);
or U3323 (N_3323,N_3233,N_3202);
nor U3324 (N_3324,N_3248,N_3227);
or U3325 (N_3325,N_3207,N_3278);
nand U3326 (N_3326,N_3298,N_3252);
and U3327 (N_3327,N_3283,N_3216);
nor U3328 (N_3328,N_3224,N_3299);
or U3329 (N_3329,N_3267,N_3263);
and U3330 (N_3330,N_3289,N_3235);
and U3331 (N_3331,N_3225,N_3236);
nand U3332 (N_3332,N_3219,N_3247);
nor U3333 (N_3333,N_3259,N_3212);
nor U3334 (N_3334,N_3204,N_3251);
nand U3335 (N_3335,N_3228,N_3239);
nor U3336 (N_3336,N_3253,N_3280);
nor U3337 (N_3337,N_3286,N_3241);
nand U3338 (N_3338,N_3290,N_3291);
or U3339 (N_3339,N_3279,N_3274);
nor U3340 (N_3340,N_3282,N_3210);
nor U3341 (N_3341,N_3209,N_3293);
nand U3342 (N_3342,N_3275,N_3238);
nor U3343 (N_3343,N_3264,N_3260);
nand U3344 (N_3344,N_3221,N_3255);
or U3345 (N_3345,N_3261,N_3297);
nand U3346 (N_3346,N_3296,N_3284);
nand U3347 (N_3347,N_3214,N_3295);
nor U3348 (N_3348,N_3265,N_3294);
and U3349 (N_3349,N_3254,N_3205);
and U3350 (N_3350,N_3295,N_3231);
and U3351 (N_3351,N_3266,N_3296);
xnor U3352 (N_3352,N_3211,N_3265);
xor U3353 (N_3353,N_3206,N_3222);
nand U3354 (N_3354,N_3243,N_3214);
and U3355 (N_3355,N_3257,N_3223);
nor U3356 (N_3356,N_3235,N_3238);
nand U3357 (N_3357,N_3225,N_3297);
and U3358 (N_3358,N_3250,N_3299);
nor U3359 (N_3359,N_3285,N_3289);
and U3360 (N_3360,N_3291,N_3254);
nor U3361 (N_3361,N_3267,N_3251);
or U3362 (N_3362,N_3266,N_3235);
nand U3363 (N_3363,N_3258,N_3270);
or U3364 (N_3364,N_3268,N_3206);
nand U3365 (N_3365,N_3209,N_3240);
nand U3366 (N_3366,N_3222,N_3211);
nor U3367 (N_3367,N_3219,N_3283);
and U3368 (N_3368,N_3259,N_3204);
nand U3369 (N_3369,N_3252,N_3218);
nor U3370 (N_3370,N_3294,N_3280);
nor U3371 (N_3371,N_3231,N_3248);
nand U3372 (N_3372,N_3279,N_3284);
nand U3373 (N_3373,N_3287,N_3207);
nor U3374 (N_3374,N_3232,N_3292);
nand U3375 (N_3375,N_3298,N_3282);
nor U3376 (N_3376,N_3262,N_3254);
and U3377 (N_3377,N_3262,N_3261);
nand U3378 (N_3378,N_3261,N_3274);
or U3379 (N_3379,N_3288,N_3268);
nor U3380 (N_3380,N_3244,N_3200);
and U3381 (N_3381,N_3248,N_3283);
or U3382 (N_3382,N_3260,N_3258);
and U3383 (N_3383,N_3246,N_3211);
or U3384 (N_3384,N_3284,N_3250);
or U3385 (N_3385,N_3237,N_3296);
or U3386 (N_3386,N_3284,N_3272);
or U3387 (N_3387,N_3247,N_3265);
and U3388 (N_3388,N_3232,N_3226);
or U3389 (N_3389,N_3213,N_3272);
nor U3390 (N_3390,N_3242,N_3289);
nor U3391 (N_3391,N_3265,N_3224);
or U3392 (N_3392,N_3239,N_3274);
and U3393 (N_3393,N_3204,N_3207);
nor U3394 (N_3394,N_3270,N_3212);
and U3395 (N_3395,N_3244,N_3285);
or U3396 (N_3396,N_3285,N_3249);
and U3397 (N_3397,N_3268,N_3263);
nand U3398 (N_3398,N_3260,N_3235);
nor U3399 (N_3399,N_3206,N_3273);
nor U3400 (N_3400,N_3387,N_3312);
or U3401 (N_3401,N_3354,N_3328);
nand U3402 (N_3402,N_3331,N_3314);
nand U3403 (N_3403,N_3384,N_3300);
or U3404 (N_3404,N_3315,N_3334);
nand U3405 (N_3405,N_3368,N_3364);
or U3406 (N_3406,N_3391,N_3390);
and U3407 (N_3407,N_3355,N_3339);
and U3408 (N_3408,N_3371,N_3381);
or U3409 (N_3409,N_3394,N_3356);
or U3410 (N_3410,N_3378,N_3335);
or U3411 (N_3411,N_3348,N_3379);
and U3412 (N_3412,N_3377,N_3319);
nand U3413 (N_3413,N_3304,N_3393);
or U3414 (N_3414,N_3359,N_3326);
and U3415 (N_3415,N_3370,N_3389);
nand U3416 (N_3416,N_3374,N_3320);
nor U3417 (N_3417,N_3347,N_3395);
nor U3418 (N_3418,N_3330,N_3317);
and U3419 (N_3419,N_3396,N_3398);
xor U3420 (N_3420,N_3383,N_3349);
nor U3421 (N_3421,N_3376,N_3316);
nand U3422 (N_3422,N_3380,N_3340);
or U3423 (N_3423,N_3323,N_3322);
nor U3424 (N_3424,N_3325,N_3333);
or U3425 (N_3425,N_3329,N_3306);
and U3426 (N_3426,N_3352,N_3307);
or U3427 (N_3427,N_3308,N_3399);
and U3428 (N_3428,N_3382,N_3338);
nor U3429 (N_3429,N_3375,N_3369);
nor U3430 (N_3430,N_3372,N_3373);
nor U3431 (N_3431,N_3385,N_3366);
xnor U3432 (N_3432,N_3361,N_3341);
nand U3433 (N_3433,N_3313,N_3321);
and U3434 (N_3434,N_3342,N_3346);
nor U3435 (N_3435,N_3309,N_3367);
or U3436 (N_3436,N_3311,N_3332);
nand U3437 (N_3437,N_3305,N_3344);
nand U3438 (N_3438,N_3318,N_3345);
xnor U3439 (N_3439,N_3336,N_3388);
nand U3440 (N_3440,N_3351,N_3357);
xor U3441 (N_3441,N_3310,N_3362);
nor U3442 (N_3442,N_3324,N_3358);
or U3443 (N_3443,N_3343,N_3303);
nor U3444 (N_3444,N_3365,N_3397);
and U3445 (N_3445,N_3337,N_3353);
or U3446 (N_3446,N_3327,N_3350);
and U3447 (N_3447,N_3386,N_3363);
nand U3448 (N_3448,N_3301,N_3302);
nand U3449 (N_3449,N_3360,N_3392);
and U3450 (N_3450,N_3350,N_3334);
xnor U3451 (N_3451,N_3395,N_3303);
nor U3452 (N_3452,N_3332,N_3323);
nand U3453 (N_3453,N_3381,N_3346);
and U3454 (N_3454,N_3345,N_3303);
nand U3455 (N_3455,N_3394,N_3321);
or U3456 (N_3456,N_3348,N_3308);
or U3457 (N_3457,N_3399,N_3338);
and U3458 (N_3458,N_3399,N_3343);
and U3459 (N_3459,N_3309,N_3369);
and U3460 (N_3460,N_3325,N_3344);
nand U3461 (N_3461,N_3347,N_3370);
nand U3462 (N_3462,N_3303,N_3370);
or U3463 (N_3463,N_3388,N_3394);
and U3464 (N_3464,N_3335,N_3372);
or U3465 (N_3465,N_3335,N_3312);
and U3466 (N_3466,N_3389,N_3343);
nor U3467 (N_3467,N_3317,N_3350);
or U3468 (N_3468,N_3386,N_3364);
and U3469 (N_3469,N_3306,N_3339);
and U3470 (N_3470,N_3314,N_3368);
nor U3471 (N_3471,N_3377,N_3365);
nand U3472 (N_3472,N_3381,N_3394);
nand U3473 (N_3473,N_3363,N_3308);
nor U3474 (N_3474,N_3397,N_3355);
xnor U3475 (N_3475,N_3309,N_3312);
and U3476 (N_3476,N_3390,N_3318);
nand U3477 (N_3477,N_3394,N_3375);
or U3478 (N_3478,N_3340,N_3360);
and U3479 (N_3479,N_3387,N_3359);
and U3480 (N_3480,N_3330,N_3352);
nor U3481 (N_3481,N_3343,N_3324);
nor U3482 (N_3482,N_3378,N_3353);
nor U3483 (N_3483,N_3307,N_3391);
and U3484 (N_3484,N_3388,N_3314);
nor U3485 (N_3485,N_3306,N_3374);
and U3486 (N_3486,N_3360,N_3398);
nand U3487 (N_3487,N_3305,N_3347);
nand U3488 (N_3488,N_3342,N_3399);
nor U3489 (N_3489,N_3329,N_3366);
nor U3490 (N_3490,N_3340,N_3325);
or U3491 (N_3491,N_3327,N_3333);
or U3492 (N_3492,N_3348,N_3388);
nand U3493 (N_3493,N_3357,N_3336);
nand U3494 (N_3494,N_3391,N_3335);
and U3495 (N_3495,N_3337,N_3382);
and U3496 (N_3496,N_3388,N_3325);
and U3497 (N_3497,N_3391,N_3350);
nand U3498 (N_3498,N_3311,N_3335);
and U3499 (N_3499,N_3336,N_3360);
and U3500 (N_3500,N_3489,N_3407);
or U3501 (N_3501,N_3477,N_3490);
or U3502 (N_3502,N_3445,N_3430);
nand U3503 (N_3503,N_3481,N_3494);
nor U3504 (N_3504,N_3434,N_3436);
or U3505 (N_3505,N_3485,N_3405);
nor U3506 (N_3506,N_3410,N_3422);
xnor U3507 (N_3507,N_3462,N_3483);
nor U3508 (N_3508,N_3460,N_3435);
and U3509 (N_3509,N_3470,N_3418);
nor U3510 (N_3510,N_3471,N_3473);
or U3511 (N_3511,N_3484,N_3466);
nor U3512 (N_3512,N_3474,N_3451);
or U3513 (N_3513,N_3472,N_3414);
and U3514 (N_3514,N_3459,N_3480);
nand U3515 (N_3515,N_3440,N_3403);
nand U3516 (N_3516,N_3411,N_3493);
or U3517 (N_3517,N_3443,N_3495);
nor U3518 (N_3518,N_3448,N_3433);
nand U3519 (N_3519,N_3429,N_3468);
or U3520 (N_3520,N_3450,N_3469);
and U3521 (N_3521,N_3413,N_3424);
and U3522 (N_3522,N_3421,N_3408);
nor U3523 (N_3523,N_3498,N_3499);
or U3524 (N_3524,N_3453,N_3457);
or U3525 (N_3525,N_3416,N_3496);
nor U3526 (N_3526,N_3446,N_3406);
nand U3527 (N_3527,N_3491,N_3417);
nor U3528 (N_3528,N_3400,N_3488);
nor U3529 (N_3529,N_3486,N_3482);
nand U3530 (N_3530,N_3402,N_3415);
nor U3531 (N_3531,N_3441,N_3449);
and U3532 (N_3532,N_3423,N_3420);
nand U3533 (N_3533,N_3438,N_3412);
nand U3534 (N_3534,N_3428,N_3401);
or U3535 (N_3535,N_3465,N_3476);
and U3536 (N_3536,N_3404,N_3455);
nand U3537 (N_3537,N_3458,N_3437);
or U3538 (N_3538,N_3478,N_3425);
or U3539 (N_3539,N_3439,N_3444);
and U3540 (N_3540,N_3456,N_3467);
nor U3541 (N_3541,N_3447,N_3492);
nand U3542 (N_3542,N_3431,N_3479);
or U3543 (N_3543,N_3426,N_3497);
or U3544 (N_3544,N_3475,N_3427);
and U3545 (N_3545,N_3409,N_3442);
nor U3546 (N_3546,N_3452,N_3461);
xor U3547 (N_3547,N_3432,N_3487);
nand U3548 (N_3548,N_3454,N_3463);
or U3549 (N_3549,N_3419,N_3464);
nand U3550 (N_3550,N_3404,N_3410);
nand U3551 (N_3551,N_3484,N_3437);
and U3552 (N_3552,N_3430,N_3437);
nand U3553 (N_3553,N_3487,N_3440);
nand U3554 (N_3554,N_3444,N_3437);
nor U3555 (N_3555,N_3461,N_3418);
nand U3556 (N_3556,N_3414,N_3486);
or U3557 (N_3557,N_3449,N_3484);
nand U3558 (N_3558,N_3456,N_3410);
and U3559 (N_3559,N_3481,N_3473);
or U3560 (N_3560,N_3427,N_3483);
nor U3561 (N_3561,N_3442,N_3477);
nand U3562 (N_3562,N_3448,N_3493);
nand U3563 (N_3563,N_3423,N_3459);
nor U3564 (N_3564,N_3468,N_3403);
nand U3565 (N_3565,N_3491,N_3422);
nor U3566 (N_3566,N_3495,N_3444);
and U3567 (N_3567,N_3494,N_3402);
and U3568 (N_3568,N_3473,N_3479);
and U3569 (N_3569,N_3402,N_3413);
and U3570 (N_3570,N_3403,N_3497);
nor U3571 (N_3571,N_3449,N_3471);
and U3572 (N_3572,N_3463,N_3435);
or U3573 (N_3573,N_3467,N_3431);
nor U3574 (N_3574,N_3409,N_3405);
xnor U3575 (N_3575,N_3451,N_3493);
or U3576 (N_3576,N_3448,N_3444);
and U3577 (N_3577,N_3463,N_3478);
and U3578 (N_3578,N_3403,N_3444);
nand U3579 (N_3579,N_3431,N_3472);
or U3580 (N_3580,N_3483,N_3418);
nand U3581 (N_3581,N_3419,N_3448);
xnor U3582 (N_3582,N_3446,N_3449);
nor U3583 (N_3583,N_3419,N_3414);
or U3584 (N_3584,N_3410,N_3449);
or U3585 (N_3585,N_3440,N_3494);
nand U3586 (N_3586,N_3416,N_3460);
nor U3587 (N_3587,N_3478,N_3461);
and U3588 (N_3588,N_3421,N_3441);
or U3589 (N_3589,N_3439,N_3485);
or U3590 (N_3590,N_3444,N_3478);
nor U3591 (N_3591,N_3491,N_3436);
and U3592 (N_3592,N_3480,N_3422);
nand U3593 (N_3593,N_3456,N_3413);
xor U3594 (N_3594,N_3466,N_3498);
or U3595 (N_3595,N_3442,N_3451);
or U3596 (N_3596,N_3494,N_3472);
or U3597 (N_3597,N_3425,N_3411);
nand U3598 (N_3598,N_3466,N_3402);
or U3599 (N_3599,N_3437,N_3415);
or U3600 (N_3600,N_3530,N_3542);
nor U3601 (N_3601,N_3500,N_3539);
nand U3602 (N_3602,N_3534,N_3514);
nand U3603 (N_3603,N_3505,N_3591);
nand U3604 (N_3604,N_3503,N_3504);
nor U3605 (N_3605,N_3533,N_3592);
nor U3606 (N_3606,N_3548,N_3595);
or U3607 (N_3607,N_3553,N_3519);
nand U3608 (N_3608,N_3521,N_3598);
nand U3609 (N_3609,N_3565,N_3577);
or U3610 (N_3610,N_3515,N_3545);
or U3611 (N_3611,N_3576,N_3568);
nand U3612 (N_3612,N_3543,N_3540);
and U3613 (N_3613,N_3506,N_3527);
nand U3614 (N_3614,N_3554,N_3574);
nand U3615 (N_3615,N_3552,N_3585);
nor U3616 (N_3616,N_3523,N_3575);
and U3617 (N_3617,N_3570,N_3509);
and U3618 (N_3618,N_3562,N_3586);
nor U3619 (N_3619,N_3547,N_3535);
nor U3620 (N_3620,N_3531,N_3549);
nand U3621 (N_3621,N_3511,N_3528);
nand U3622 (N_3622,N_3522,N_3561);
and U3623 (N_3623,N_3520,N_3590);
or U3624 (N_3624,N_3510,N_3507);
nor U3625 (N_3625,N_3513,N_3516);
nand U3626 (N_3626,N_3569,N_3583);
nor U3627 (N_3627,N_3578,N_3594);
or U3628 (N_3628,N_3596,N_3538);
xor U3629 (N_3629,N_3557,N_3597);
xor U3630 (N_3630,N_3571,N_3532);
nand U3631 (N_3631,N_3556,N_3599);
or U3632 (N_3632,N_3544,N_3555);
or U3633 (N_3633,N_3589,N_3508);
or U3634 (N_3634,N_3587,N_3518);
or U3635 (N_3635,N_3579,N_3541);
and U3636 (N_3636,N_3572,N_3537);
or U3637 (N_3637,N_3512,N_3566);
and U3638 (N_3638,N_3588,N_3559);
and U3639 (N_3639,N_3551,N_3502);
nor U3640 (N_3640,N_3529,N_3584);
nor U3641 (N_3641,N_3536,N_3525);
and U3642 (N_3642,N_3558,N_3593);
and U3643 (N_3643,N_3546,N_3582);
nand U3644 (N_3644,N_3580,N_3524);
nand U3645 (N_3645,N_3573,N_3526);
and U3646 (N_3646,N_3550,N_3567);
nor U3647 (N_3647,N_3517,N_3501);
and U3648 (N_3648,N_3564,N_3563);
and U3649 (N_3649,N_3581,N_3560);
nor U3650 (N_3650,N_3551,N_3507);
and U3651 (N_3651,N_3510,N_3563);
or U3652 (N_3652,N_3557,N_3583);
nor U3653 (N_3653,N_3573,N_3553);
nor U3654 (N_3654,N_3589,N_3519);
nor U3655 (N_3655,N_3552,N_3565);
nand U3656 (N_3656,N_3558,N_3585);
nor U3657 (N_3657,N_3510,N_3529);
and U3658 (N_3658,N_3555,N_3534);
or U3659 (N_3659,N_3593,N_3539);
or U3660 (N_3660,N_3519,N_3506);
nor U3661 (N_3661,N_3549,N_3571);
nor U3662 (N_3662,N_3561,N_3521);
or U3663 (N_3663,N_3588,N_3511);
and U3664 (N_3664,N_3500,N_3575);
nor U3665 (N_3665,N_3513,N_3550);
and U3666 (N_3666,N_3539,N_3549);
and U3667 (N_3667,N_3566,N_3519);
and U3668 (N_3668,N_3512,N_3565);
nor U3669 (N_3669,N_3524,N_3528);
nor U3670 (N_3670,N_3568,N_3523);
nor U3671 (N_3671,N_3507,N_3528);
nor U3672 (N_3672,N_3593,N_3541);
and U3673 (N_3673,N_3555,N_3512);
or U3674 (N_3674,N_3583,N_3555);
xor U3675 (N_3675,N_3539,N_3566);
and U3676 (N_3676,N_3568,N_3521);
and U3677 (N_3677,N_3501,N_3586);
or U3678 (N_3678,N_3555,N_3517);
nor U3679 (N_3679,N_3544,N_3567);
and U3680 (N_3680,N_3515,N_3579);
or U3681 (N_3681,N_3558,N_3516);
nand U3682 (N_3682,N_3582,N_3561);
or U3683 (N_3683,N_3560,N_3597);
or U3684 (N_3684,N_3551,N_3559);
and U3685 (N_3685,N_3597,N_3520);
and U3686 (N_3686,N_3518,N_3549);
and U3687 (N_3687,N_3590,N_3595);
nand U3688 (N_3688,N_3515,N_3589);
nor U3689 (N_3689,N_3581,N_3523);
nand U3690 (N_3690,N_3565,N_3545);
or U3691 (N_3691,N_3552,N_3511);
or U3692 (N_3692,N_3554,N_3599);
or U3693 (N_3693,N_3557,N_3511);
nor U3694 (N_3694,N_3590,N_3546);
or U3695 (N_3695,N_3578,N_3589);
and U3696 (N_3696,N_3542,N_3503);
or U3697 (N_3697,N_3550,N_3546);
or U3698 (N_3698,N_3593,N_3591);
or U3699 (N_3699,N_3541,N_3537);
and U3700 (N_3700,N_3683,N_3672);
nor U3701 (N_3701,N_3688,N_3634);
or U3702 (N_3702,N_3679,N_3644);
or U3703 (N_3703,N_3658,N_3605);
xnor U3704 (N_3704,N_3604,N_3684);
or U3705 (N_3705,N_3662,N_3641);
or U3706 (N_3706,N_3686,N_3667);
nand U3707 (N_3707,N_3668,N_3642);
or U3708 (N_3708,N_3613,N_3606);
or U3709 (N_3709,N_3695,N_3612);
and U3710 (N_3710,N_3636,N_3615);
or U3711 (N_3711,N_3653,N_3692);
nand U3712 (N_3712,N_3687,N_3671);
or U3713 (N_3713,N_3623,N_3680);
nand U3714 (N_3714,N_3698,N_3626);
xnor U3715 (N_3715,N_3639,N_3611);
or U3716 (N_3716,N_3652,N_3640);
nand U3717 (N_3717,N_3625,N_3622);
nor U3718 (N_3718,N_3696,N_3670);
nor U3719 (N_3719,N_3651,N_3638);
or U3720 (N_3720,N_3685,N_3621);
and U3721 (N_3721,N_3659,N_3661);
nor U3722 (N_3722,N_3609,N_3690);
or U3723 (N_3723,N_3643,N_3616);
or U3724 (N_3724,N_3673,N_3628);
nand U3725 (N_3725,N_3693,N_3629);
nand U3726 (N_3726,N_3631,N_3655);
and U3727 (N_3727,N_3663,N_3656);
and U3728 (N_3728,N_3601,N_3691);
or U3729 (N_3729,N_3689,N_3650);
nor U3730 (N_3730,N_3678,N_3632);
and U3731 (N_3731,N_3624,N_3618);
nor U3732 (N_3732,N_3660,N_3664);
nor U3733 (N_3733,N_3682,N_3610);
and U3734 (N_3734,N_3602,N_3677);
nand U3735 (N_3735,N_3607,N_3608);
nand U3736 (N_3736,N_3666,N_3633);
nand U3737 (N_3737,N_3697,N_3649);
nand U3738 (N_3738,N_3630,N_3681);
nand U3739 (N_3739,N_3694,N_3645);
nand U3740 (N_3740,N_3617,N_3637);
nand U3741 (N_3741,N_3627,N_3674);
nor U3742 (N_3742,N_3635,N_3648);
nand U3743 (N_3743,N_3676,N_3646);
nor U3744 (N_3744,N_3620,N_3614);
nand U3745 (N_3745,N_3600,N_3619);
or U3746 (N_3746,N_3657,N_3699);
nand U3747 (N_3747,N_3647,N_3675);
nand U3748 (N_3748,N_3654,N_3669);
and U3749 (N_3749,N_3603,N_3665);
or U3750 (N_3750,N_3651,N_3604);
and U3751 (N_3751,N_3674,N_3642);
and U3752 (N_3752,N_3608,N_3648);
and U3753 (N_3753,N_3654,N_3697);
xor U3754 (N_3754,N_3680,N_3673);
nand U3755 (N_3755,N_3644,N_3611);
nor U3756 (N_3756,N_3696,N_3646);
nor U3757 (N_3757,N_3643,N_3624);
and U3758 (N_3758,N_3629,N_3627);
or U3759 (N_3759,N_3631,N_3687);
and U3760 (N_3760,N_3655,N_3614);
or U3761 (N_3761,N_3628,N_3662);
nor U3762 (N_3762,N_3616,N_3653);
xnor U3763 (N_3763,N_3697,N_3688);
nand U3764 (N_3764,N_3688,N_3619);
nor U3765 (N_3765,N_3699,N_3686);
and U3766 (N_3766,N_3684,N_3627);
nor U3767 (N_3767,N_3623,N_3653);
nor U3768 (N_3768,N_3618,N_3649);
and U3769 (N_3769,N_3634,N_3692);
xor U3770 (N_3770,N_3688,N_3649);
or U3771 (N_3771,N_3675,N_3650);
and U3772 (N_3772,N_3680,N_3635);
and U3773 (N_3773,N_3611,N_3605);
or U3774 (N_3774,N_3634,N_3628);
nor U3775 (N_3775,N_3678,N_3670);
nand U3776 (N_3776,N_3621,N_3613);
or U3777 (N_3777,N_3646,N_3655);
or U3778 (N_3778,N_3635,N_3601);
nand U3779 (N_3779,N_3607,N_3674);
and U3780 (N_3780,N_3690,N_3646);
and U3781 (N_3781,N_3686,N_3629);
nand U3782 (N_3782,N_3681,N_3602);
nand U3783 (N_3783,N_3635,N_3627);
nor U3784 (N_3784,N_3681,N_3687);
or U3785 (N_3785,N_3668,N_3614);
or U3786 (N_3786,N_3671,N_3601);
nor U3787 (N_3787,N_3629,N_3665);
or U3788 (N_3788,N_3662,N_3699);
nor U3789 (N_3789,N_3685,N_3679);
nand U3790 (N_3790,N_3678,N_3648);
nand U3791 (N_3791,N_3659,N_3618);
xnor U3792 (N_3792,N_3636,N_3678);
nor U3793 (N_3793,N_3626,N_3604);
nor U3794 (N_3794,N_3637,N_3689);
or U3795 (N_3795,N_3624,N_3665);
nor U3796 (N_3796,N_3634,N_3673);
and U3797 (N_3797,N_3604,N_3679);
and U3798 (N_3798,N_3632,N_3647);
nand U3799 (N_3799,N_3602,N_3626);
or U3800 (N_3800,N_3718,N_3774);
nand U3801 (N_3801,N_3772,N_3784);
and U3802 (N_3802,N_3712,N_3737);
nor U3803 (N_3803,N_3764,N_3738);
and U3804 (N_3804,N_3717,N_3746);
nand U3805 (N_3805,N_3796,N_3765);
nor U3806 (N_3806,N_3742,N_3781);
nor U3807 (N_3807,N_3782,N_3794);
or U3808 (N_3808,N_3729,N_3769);
or U3809 (N_3809,N_3749,N_3778);
or U3810 (N_3810,N_3709,N_3768);
and U3811 (N_3811,N_3779,N_3702);
nor U3812 (N_3812,N_3722,N_3741);
and U3813 (N_3813,N_3786,N_3789);
or U3814 (N_3814,N_3705,N_3734);
and U3815 (N_3815,N_3799,N_3760);
nor U3816 (N_3816,N_3748,N_3770);
nand U3817 (N_3817,N_3750,N_3703);
nor U3818 (N_3818,N_3708,N_3735);
or U3819 (N_3819,N_3771,N_3753);
or U3820 (N_3820,N_3767,N_3798);
and U3821 (N_3821,N_3785,N_3721);
or U3822 (N_3822,N_3783,N_3756);
and U3823 (N_3823,N_3728,N_3706);
xor U3824 (N_3824,N_3777,N_3704);
or U3825 (N_3825,N_3743,N_3795);
or U3826 (N_3826,N_3793,N_3797);
or U3827 (N_3827,N_3720,N_3711);
nor U3828 (N_3828,N_3775,N_3790);
and U3829 (N_3829,N_3700,N_3733);
nand U3830 (N_3830,N_3730,N_3792);
nand U3831 (N_3831,N_3755,N_3736);
or U3832 (N_3832,N_3739,N_3715);
and U3833 (N_3833,N_3744,N_3732);
nand U3834 (N_3834,N_3759,N_3731);
or U3835 (N_3835,N_3776,N_3719);
nor U3836 (N_3836,N_3714,N_3745);
xor U3837 (N_3837,N_3727,N_3701);
or U3838 (N_3838,N_3763,N_3740);
nor U3839 (N_3839,N_3725,N_3791);
and U3840 (N_3840,N_3710,N_3788);
and U3841 (N_3841,N_3747,N_3723);
and U3842 (N_3842,N_3787,N_3751);
or U3843 (N_3843,N_3754,N_3762);
nand U3844 (N_3844,N_3726,N_3761);
or U3845 (N_3845,N_3773,N_3752);
nor U3846 (N_3846,N_3707,N_3780);
or U3847 (N_3847,N_3713,N_3757);
nor U3848 (N_3848,N_3758,N_3724);
nor U3849 (N_3849,N_3716,N_3766);
nand U3850 (N_3850,N_3774,N_3765);
nor U3851 (N_3851,N_3791,N_3718);
or U3852 (N_3852,N_3736,N_3721);
nand U3853 (N_3853,N_3783,N_3707);
or U3854 (N_3854,N_3760,N_3704);
and U3855 (N_3855,N_3748,N_3747);
and U3856 (N_3856,N_3742,N_3703);
nor U3857 (N_3857,N_3705,N_3798);
nor U3858 (N_3858,N_3750,N_3713);
nand U3859 (N_3859,N_3719,N_3702);
nand U3860 (N_3860,N_3718,N_3785);
or U3861 (N_3861,N_3740,N_3733);
nand U3862 (N_3862,N_3794,N_3787);
nand U3863 (N_3863,N_3743,N_3764);
nand U3864 (N_3864,N_3736,N_3703);
nor U3865 (N_3865,N_3790,N_3750);
nand U3866 (N_3866,N_3709,N_3774);
and U3867 (N_3867,N_3741,N_3782);
and U3868 (N_3868,N_3723,N_3775);
or U3869 (N_3869,N_3706,N_3712);
nand U3870 (N_3870,N_3754,N_3789);
and U3871 (N_3871,N_3785,N_3736);
nor U3872 (N_3872,N_3780,N_3738);
nor U3873 (N_3873,N_3765,N_3724);
nor U3874 (N_3874,N_3755,N_3713);
and U3875 (N_3875,N_3705,N_3799);
nor U3876 (N_3876,N_3772,N_3748);
nand U3877 (N_3877,N_3766,N_3793);
nor U3878 (N_3878,N_3713,N_3731);
or U3879 (N_3879,N_3703,N_3752);
and U3880 (N_3880,N_3784,N_3735);
nand U3881 (N_3881,N_3762,N_3749);
or U3882 (N_3882,N_3720,N_3726);
nand U3883 (N_3883,N_3748,N_3700);
nand U3884 (N_3884,N_3770,N_3799);
nor U3885 (N_3885,N_3715,N_3726);
nand U3886 (N_3886,N_3717,N_3784);
or U3887 (N_3887,N_3750,N_3755);
nand U3888 (N_3888,N_3781,N_3747);
nor U3889 (N_3889,N_3793,N_3748);
or U3890 (N_3890,N_3718,N_3759);
nand U3891 (N_3891,N_3748,N_3774);
xor U3892 (N_3892,N_3739,N_3703);
and U3893 (N_3893,N_3784,N_3791);
and U3894 (N_3894,N_3711,N_3734);
nand U3895 (N_3895,N_3778,N_3751);
nor U3896 (N_3896,N_3748,N_3759);
nor U3897 (N_3897,N_3746,N_3750);
and U3898 (N_3898,N_3735,N_3742);
nor U3899 (N_3899,N_3799,N_3797);
xnor U3900 (N_3900,N_3885,N_3826);
nor U3901 (N_3901,N_3896,N_3851);
or U3902 (N_3902,N_3888,N_3898);
nor U3903 (N_3903,N_3852,N_3861);
xnor U3904 (N_3904,N_3822,N_3843);
or U3905 (N_3905,N_3876,N_3835);
and U3906 (N_3906,N_3842,N_3867);
nor U3907 (N_3907,N_3817,N_3877);
and U3908 (N_3908,N_3827,N_3804);
or U3909 (N_3909,N_3809,N_3890);
and U3910 (N_3910,N_3868,N_3862);
nor U3911 (N_3911,N_3849,N_3805);
nand U3912 (N_3912,N_3860,N_3841);
and U3913 (N_3913,N_3857,N_3854);
nand U3914 (N_3914,N_3800,N_3889);
nand U3915 (N_3915,N_3897,N_3875);
or U3916 (N_3916,N_3831,N_3895);
or U3917 (N_3917,N_3893,N_3883);
xnor U3918 (N_3918,N_3886,N_3818);
nor U3919 (N_3919,N_3846,N_3887);
nor U3920 (N_3920,N_3821,N_3836);
or U3921 (N_3921,N_3801,N_3892);
and U3922 (N_3922,N_3833,N_3830);
nand U3923 (N_3923,N_3807,N_3812);
nor U3924 (N_3924,N_3824,N_3864);
and U3925 (N_3925,N_3806,N_3850);
nor U3926 (N_3926,N_3844,N_3874);
and U3927 (N_3927,N_3823,N_3829);
nor U3928 (N_3928,N_3848,N_3853);
or U3929 (N_3929,N_3815,N_3870);
and U3930 (N_3930,N_3882,N_3802);
nor U3931 (N_3931,N_3873,N_3872);
or U3932 (N_3932,N_3819,N_3856);
nor U3933 (N_3933,N_3816,N_3866);
nor U3934 (N_3934,N_3832,N_3839);
and U3935 (N_3935,N_3810,N_3845);
or U3936 (N_3936,N_3847,N_3878);
or U3937 (N_3937,N_3880,N_3840);
nand U3938 (N_3938,N_3814,N_3859);
nor U3939 (N_3939,N_3879,N_3825);
nor U3940 (N_3940,N_3855,N_3811);
nand U3941 (N_3941,N_3863,N_3865);
nand U3942 (N_3942,N_3820,N_3828);
nand U3943 (N_3943,N_3884,N_3891);
nor U3944 (N_3944,N_3899,N_3894);
or U3945 (N_3945,N_3837,N_3808);
and U3946 (N_3946,N_3813,N_3838);
nor U3947 (N_3947,N_3869,N_3803);
nor U3948 (N_3948,N_3834,N_3858);
xnor U3949 (N_3949,N_3871,N_3881);
nor U3950 (N_3950,N_3872,N_3870);
nand U3951 (N_3951,N_3861,N_3813);
nand U3952 (N_3952,N_3827,N_3805);
and U3953 (N_3953,N_3847,N_3827);
or U3954 (N_3954,N_3818,N_3850);
nand U3955 (N_3955,N_3883,N_3843);
xor U3956 (N_3956,N_3858,N_3826);
and U3957 (N_3957,N_3852,N_3804);
and U3958 (N_3958,N_3808,N_3823);
or U3959 (N_3959,N_3805,N_3867);
nor U3960 (N_3960,N_3825,N_3859);
nand U3961 (N_3961,N_3899,N_3853);
nand U3962 (N_3962,N_3837,N_3828);
nor U3963 (N_3963,N_3859,N_3844);
or U3964 (N_3964,N_3846,N_3853);
or U3965 (N_3965,N_3805,N_3893);
or U3966 (N_3966,N_3864,N_3870);
and U3967 (N_3967,N_3842,N_3807);
and U3968 (N_3968,N_3848,N_3889);
nor U3969 (N_3969,N_3891,N_3863);
nor U3970 (N_3970,N_3883,N_3801);
nand U3971 (N_3971,N_3880,N_3820);
and U3972 (N_3972,N_3857,N_3832);
nor U3973 (N_3973,N_3878,N_3833);
nand U3974 (N_3974,N_3818,N_3827);
or U3975 (N_3975,N_3874,N_3806);
nand U3976 (N_3976,N_3874,N_3892);
or U3977 (N_3977,N_3873,N_3868);
and U3978 (N_3978,N_3833,N_3822);
or U3979 (N_3979,N_3857,N_3863);
nand U3980 (N_3980,N_3819,N_3851);
xor U3981 (N_3981,N_3878,N_3816);
nor U3982 (N_3982,N_3821,N_3820);
and U3983 (N_3983,N_3858,N_3890);
nor U3984 (N_3984,N_3825,N_3849);
nor U3985 (N_3985,N_3896,N_3827);
nor U3986 (N_3986,N_3844,N_3892);
and U3987 (N_3987,N_3840,N_3867);
nand U3988 (N_3988,N_3877,N_3816);
and U3989 (N_3989,N_3895,N_3827);
and U3990 (N_3990,N_3844,N_3850);
or U3991 (N_3991,N_3828,N_3867);
and U3992 (N_3992,N_3861,N_3853);
nor U3993 (N_3993,N_3892,N_3878);
or U3994 (N_3994,N_3860,N_3889);
and U3995 (N_3995,N_3856,N_3834);
nand U3996 (N_3996,N_3817,N_3855);
nand U3997 (N_3997,N_3833,N_3819);
nor U3998 (N_3998,N_3804,N_3893);
or U3999 (N_3999,N_3846,N_3873);
or U4000 (N_4000,N_3927,N_3992);
nand U4001 (N_4001,N_3956,N_3983);
and U4002 (N_4002,N_3930,N_3903);
nor U4003 (N_4003,N_3969,N_3904);
nor U4004 (N_4004,N_3978,N_3906);
nand U4005 (N_4005,N_3937,N_3981);
or U4006 (N_4006,N_3924,N_3994);
and U4007 (N_4007,N_3996,N_3967);
nand U4008 (N_4008,N_3988,N_3952);
nand U4009 (N_4009,N_3997,N_3949);
nand U4010 (N_4010,N_3929,N_3914);
and U4011 (N_4011,N_3966,N_3963);
nand U4012 (N_4012,N_3970,N_3923);
nand U4013 (N_4013,N_3954,N_3979);
nor U4014 (N_4014,N_3934,N_3971);
nand U4015 (N_4015,N_3999,N_3936);
and U4016 (N_4016,N_3907,N_3910);
nand U4017 (N_4017,N_3908,N_3912);
and U4018 (N_4018,N_3995,N_3985);
and U4019 (N_4019,N_3987,N_3947);
nor U4020 (N_4020,N_3958,N_3974);
and U4021 (N_4021,N_3977,N_3942);
xnor U4022 (N_4022,N_3959,N_3964);
nor U4023 (N_4023,N_3986,N_3989);
or U4024 (N_4024,N_3955,N_3957);
and U4025 (N_4025,N_3928,N_3975);
nor U4026 (N_4026,N_3915,N_3972);
nor U4027 (N_4027,N_3900,N_3931);
nor U4028 (N_4028,N_3911,N_3933);
and U4029 (N_4029,N_3953,N_3935);
and U4030 (N_4030,N_3913,N_3951);
nor U4031 (N_4031,N_3918,N_3901);
nor U4032 (N_4032,N_3922,N_3944);
nand U4033 (N_4033,N_3991,N_3973);
nand U4034 (N_4034,N_3948,N_3960);
and U4035 (N_4035,N_3902,N_3998);
nor U4036 (N_4036,N_3968,N_3940);
or U4037 (N_4037,N_3905,N_3965);
nor U4038 (N_4038,N_3932,N_3926);
nand U4039 (N_4039,N_3909,N_3982);
nor U4040 (N_4040,N_3945,N_3946);
or U4041 (N_4041,N_3939,N_3990);
and U4042 (N_4042,N_3950,N_3920);
nor U4043 (N_4043,N_3916,N_3921);
nor U4044 (N_4044,N_3976,N_3980);
nand U4045 (N_4045,N_3961,N_3919);
nand U4046 (N_4046,N_3917,N_3938);
xnor U4047 (N_4047,N_3925,N_3993);
nor U4048 (N_4048,N_3943,N_3962);
nor U4049 (N_4049,N_3984,N_3941);
nor U4050 (N_4050,N_3901,N_3977);
and U4051 (N_4051,N_3947,N_3921);
nand U4052 (N_4052,N_3974,N_3907);
and U4053 (N_4053,N_3989,N_3906);
nor U4054 (N_4054,N_3978,N_3912);
or U4055 (N_4055,N_3908,N_3964);
and U4056 (N_4056,N_3936,N_3947);
or U4057 (N_4057,N_3914,N_3927);
or U4058 (N_4058,N_3938,N_3911);
and U4059 (N_4059,N_3962,N_3915);
nor U4060 (N_4060,N_3964,N_3914);
or U4061 (N_4061,N_3977,N_3941);
nand U4062 (N_4062,N_3986,N_3967);
nor U4063 (N_4063,N_3983,N_3949);
and U4064 (N_4064,N_3964,N_3905);
nand U4065 (N_4065,N_3988,N_3946);
nand U4066 (N_4066,N_3967,N_3924);
nor U4067 (N_4067,N_3947,N_3972);
and U4068 (N_4068,N_3915,N_3989);
nand U4069 (N_4069,N_3914,N_3949);
and U4070 (N_4070,N_3947,N_3966);
nor U4071 (N_4071,N_3937,N_3956);
or U4072 (N_4072,N_3956,N_3980);
nand U4073 (N_4073,N_3948,N_3949);
and U4074 (N_4074,N_3979,N_3910);
nand U4075 (N_4075,N_3939,N_3962);
nand U4076 (N_4076,N_3952,N_3900);
or U4077 (N_4077,N_3990,N_3976);
or U4078 (N_4078,N_3982,N_3962);
nand U4079 (N_4079,N_3974,N_3914);
and U4080 (N_4080,N_3929,N_3931);
or U4081 (N_4081,N_3932,N_3943);
nand U4082 (N_4082,N_3994,N_3917);
nor U4083 (N_4083,N_3919,N_3956);
nor U4084 (N_4084,N_3945,N_3919);
and U4085 (N_4085,N_3989,N_3934);
nand U4086 (N_4086,N_3986,N_3973);
nand U4087 (N_4087,N_3916,N_3904);
xnor U4088 (N_4088,N_3991,N_3918);
nor U4089 (N_4089,N_3959,N_3992);
or U4090 (N_4090,N_3943,N_3921);
and U4091 (N_4091,N_3901,N_3927);
nand U4092 (N_4092,N_3912,N_3906);
and U4093 (N_4093,N_3918,N_3911);
and U4094 (N_4094,N_3926,N_3986);
nand U4095 (N_4095,N_3950,N_3959);
nor U4096 (N_4096,N_3950,N_3934);
nand U4097 (N_4097,N_3994,N_3912);
or U4098 (N_4098,N_3968,N_3933);
nand U4099 (N_4099,N_3935,N_3924);
nor U4100 (N_4100,N_4065,N_4039);
or U4101 (N_4101,N_4045,N_4003);
nand U4102 (N_4102,N_4052,N_4024);
or U4103 (N_4103,N_4062,N_4034);
nand U4104 (N_4104,N_4042,N_4068);
or U4105 (N_4105,N_4099,N_4040);
nor U4106 (N_4106,N_4049,N_4009);
and U4107 (N_4107,N_4057,N_4027);
nor U4108 (N_4108,N_4006,N_4063);
nand U4109 (N_4109,N_4002,N_4038);
or U4110 (N_4110,N_4035,N_4077);
nand U4111 (N_4111,N_4096,N_4022);
and U4112 (N_4112,N_4031,N_4095);
and U4113 (N_4113,N_4079,N_4093);
nand U4114 (N_4114,N_4067,N_4004);
and U4115 (N_4115,N_4051,N_4098);
nand U4116 (N_4116,N_4094,N_4029);
nand U4117 (N_4117,N_4012,N_4016);
nand U4118 (N_4118,N_4086,N_4047);
nor U4119 (N_4119,N_4085,N_4054);
and U4120 (N_4120,N_4061,N_4090);
and U4121 (N_4121,N_4007,N_4084);
and U4122 (N_4122,N_4032,N_4064);
and U4123 (N_4123,N_4021,N_4037);
nand U4124 (N_4124,N_4008,N_4078);
nand U4125 (N_4125,N_4015,N_4014);
or U4126 (N_4126,N_4053,N_4066);
or U4127 (N_4127,N_4074,N_4041);
nand U4128 (N_4128,N_4036,N_4073);
nor U4129 (N_4129,N_4019,N_4076);
and U4130 (N_4130,N_4091,N_4013);
and U4131 (N_4131,N_4080,N_4026);
or U4132 (N_4132,N_4033,N_4059);
or U4133 (N_4133,N_4050,N_4081);
nand U4134 (N_4134,N_4082,N_4097);
nor U4135 (N_4135,N_4092,N_4028);
and U4136 (N_4136,N_4071,N_4046);
or U4137 (N_4137,N_4058,N_4020);
nor U4138 (N_4138,N_4069,N_4083);
and U4139 (N_4139,N_4075,N_4011);
and U4140 (N_4140,N_4087,N_4017);
and U4141 (N_4141,N_4010,N_4070);
and U4142 (N_4142,N_4025,N_4018);
xor U4143 (N_4143,N_4060,N_4001);
nand U4144 (N_4144,N_4072,N_4048);
or U4145 (N_4145,N_4043,N_4089);
and U4146 (N_4146,N_4030,N_4000);
and U4147 (N_4147,N_4023,N_4055);
and U4148 (N_4148,N_4005,N_4044);
and U4149 (N_4149,N_4088,N_4056);
nor U4150 (N_4150,N_4006,N_4013);
and U4151 (N_4151,N_4091,N_4041);
and U4152 (N_4152,N_4036,N_4018);
or U4153 (N_4153,N_4054,N_4046);
nand U4154 (N_4154,N_4030,N_4080);
nor U4155 (N_4155,N_4041,N_4062);
and U4156 (N_4156,N_4044,N_4017);
nor U4157 (N_4157,N_4010,N_4056);
nand U4158 (N_4158,N_4063,N_4003);
nor U4159 (N_4159,N_4077,N_4012);
or U4160 (N_4160,N_4041,N_4053);
nand U4161 (N_4161,N_4065,N_4083);
or U4162 (N_4162,N_4030,N_4039);
nand U4163 (N_4163,N_4024,N_4098);
or U4164 (N_4164,N_4085,N_4063);
xnor U4165 (N_4165,N_4042,N_4070);
or U4166 (N_4166,N_4029,N_4034);
xor U4167 (N_4167,N_4040,N_4089);
or U4168 (N_4168,N_4070,N_4023);
or U4169 (N_4169,N_4044,N_4083);
or U4170 (N_4170,N_4075,N_4082);
nand U4171 (N_4171,N_4012,N_4009);
xor U4172 (N_4172,N_4037,N_4038);
nand U4173 (N_4173,N_4001,N_4012);
and U4174 (N_4174,N_4030,N_4071);
nand U4175 (N_4175,N_4029,N_4086);
and U4176 (N_4176,N_4058,N_4046);
nor U4177 (N_4177,N_4033,N_4072);
nand U4178 (N_4178,N_4050,N_4053);
or U4179 (N_4179,N_4006,N_4079);
nor U4180 (N_4180,N_4033,N_4025);
nor U4181 (N_4181,N_4053,N_4089);
or U4182 (N_4182,N_4037,N_4044);
nor U4183 (N_4183,N_4006,N_4098);
nor U4184 (N_4184,N_4090,N_4096);
or U4185 (N_4185,N_4074,N_4089);
and U4186 (N_4186,N_4050,N_4000);
nor U4187 (N_4187,N_4034,N_4059);
and U4188 (N_4188,N_4085,N_4059);
nor U4189 (N_4189,N_4044,N_4031);
and U4190 (N_4190,N_4006,N_4043);
nand U4191 (N_4191,N_4086,N_4096);
and U4192 (N_4192,N_4013,N_4037);
nand U4193 (N_4193,N_4024,N_4036);
nor U4194 (N_4194,N_4093,N_4037);
nand U4195 (N_4195,N_4067,N_4046);
nor U4196 (N_4196,N_4002,N_4032);
nor U4197 (N_4197,N_4062,N_4015);
and U4198 (N_4198,N_4047,N_4056);
nor U4199 (N_4199,N_4092,N_4055);
and U4200 (N_4200,N_4163,N_4198);
nor U4201 (N_4201,N_4146,N_4159);
nand U4202 (N_4202,N_4102,N_4116);
nor U4203 (N_4203,N_4162,N_4100);
nor U4204 (N_4204,N_4123,N_4181);
xnor U4205 (N_4205,N_4176,N_4155);
and U4206 (N_4206,N_4128,N_4186);
or U4207 (N_4207,N_4152,N_4126);
nor U4208 (N_4208,N_4174,N_4105);
nand U4209 (N_4209,N_4192,N_4122);
nand U4210 (N_4210,N_4160,N_4140);
nand U4211 (N_4211,N_4127,N_4117);
xnor U4212 (N_4212,N_4195,N_4125);
nor U4213 (N_4213,N_4131,N_4142);
and U4214 (N_4214,N_4157,N_4144);
nor U4215 (N_4215,N_4164,N_4189);
or U4216 (N_4216,N_4101,N_4183);
and U4217 (N_4217,N_4161,N_4147);
nor U4218 (N_4218,N_4143,N_4166);
or U4219 (N_4219,N_4134,N_4110);
nand U4220 (N_4220,N_4165,N_4172);
or U4221 (N_4221,N_4149,N_4141);
and U4222 (N_4222,N_4133,N_4154);
and U4223 (N_4223,N_4177,N_4194);
and U4224 (N_4224,N_4103,N_4196);
or U4225 (N_4225,N_4187,N_4178);
nor U4226 (N_4226,N_4175,N_4136);
nand U4227 (N_4227,N_4151,N_4184);
nor U4228 (N_4228,N_4106,N_4130);
and U4229 (N_4229,N_4158,N_4115);
and U4230 (N_4230,N_4188,N_4150);
nor U4231 (N_4231,N_4137,N_4107);
and U4232 (N_4232,N_4148,N_4132);
nor U4233 (N_4233,N_4113,N_4171);
or U4234 (N_4234,N_4197,N_4135);
or U4235 (N_4235,N_4129,N_4179);
nor U4236 (N_4236,N_4182,N_4170);
and U4237 (N_4237,N_4120,N_4156);
or U4238 (N_4238,N_4111,N_4112);
or U4239 (N_4239,N_4153,N_4139);
nand U4240 (N_4240,N_4190,N_4191);
nor U4241 (N_4241,N_4169,N_4121);
and U4242 (N_4242,N_4104,N_4180);
nand U4243 (N_4243,N_4167,N_4118);
or U4244 (N_4244,N_4119,N_4124);
nor U4245 (N_4245,N_4173,N_4138);
xor U4246 (N_4246,N_4193,N_4145);
and U4247 (N_4247,N_4109,N_4114);
or U4248 (N_4248,N_4185,N_4199);
nand U4249 (N_4249,N_4168,N_4108);
or U4250 (N_4250,N_4122,N_4184);
or U4251 (N_4251,N_4165,N_4161);
nand U4252 (N_4252,N_4123,N_4125);
nand U4253 (N_4253,N_4115,N_4142);
nand U4254 (N_4254,N_4122,N_4141);
nor U4255 (N_4255,N_4151,N_4122);
or U4256 (N_4256,N_4103,N_4104);
nor U4257 (N_4257,N_4191,N_4182);
nand U4258 (N_4258,N_4106,N_4128);
and U4259 (N_4259,N_4148,N_4103);
nand U4260 (N_4260,N_4157,N_4139);
and U4261 (N_4261,N_4106,N_4102);
and U4262 (N_4262,N_4198,N_4128);
or U4263 (N_4263,N_4106,N_4108);
or U4264 (N_4264,N_4106,N_4156);
xnor U4265 (N_4265,N_4115,N_4182);
and U4266 (N_4266,N_4123,N_4155);
and U4267 (N_4267,N_4176,N_4108);
and U4268 (N_4268,N_4100,N_4105);
nor U4269 (N_4269,N_4193,N_4124);
and U4270 (N_4270,N_4107,N_4128);
nand U4271 (N_4271,N_4194,N_4132);
and U4272 (N_4272,N_4130,N_4180);
or U4273 (N_4273,N_4129,N_4130);
or U4274 (N_4274,N_4115,N_4110);
nor U4275 (N_4275,N_4113,N_4194);
nor U4276 (N_4276,N_4122,N_4167);
and U4277 (N_4277,N_4173,N_4121);
nor U4278 (N_4278,N_4134,N_4152);
nor U4279 (N_4279,N_4183,N_4172);
or U4280 (N_4280,N_4146,N_4155);
or U4281 (N_4281,N_4137,N_4149);
or U4282 (N_4282,N_4166,N_4152);
and U4283 (N_4283,N_4103,N_4129);
nand U4284 (N_4284,N_4116,N_4127);
or U4285 (N_4285,N_4146,N_4176);
and U4286 (N_4286,N_4135,N_4122);
and U4287 (N_4287,N_4168,N_4102);
xor U4288 (N_4288,N_4168,N_4186);
nor U4289 (N_4289,N_4111,N_4161);
or U4290 (N_4290,N_4179,N_4114);
nor U4291 (N_4291,N_4157,N_4183);
or U4292 (N_4292,N_4141,N_4176);
nand U4293 (N_4293,N_4188,N_4105);
nand U4294 (N_4294,N_4178,N_4111);
and U4295 (N_4295,N_4146,N_4186);
nor U4296 (N_4296,N_4172,N_4138);
or U4297 (N_4297,N_4122,N_4104);
or U4298 (N_4298,N_4119,N_4130);
and U4299 (N_4299,N_4166,N_4155);
nand U4300 (N_4300,N_4244,N_4224);
and U4301 (N_4301,N_4206,N_4293);
or U4302 (N_4302,N_4259,N_4213);
nand U4303 (N_4303,N_4273,N_4245);
nand U4304 (N_4304,N_4238,N_4235);
and U4305 (N_4305,N_4265,N_4229);
or U4306 (N_4306,N_4234,N_4222);
and U4307 (N_4307,N_4276,N_4200);
or U4308 (N_4308,N_4226,N_4296);
nand U4309 (N_4309,N_4233,N_4211);
or U4310 (N_4310,N_4258,N_4254);
or U4311 (N_4311,N_4289,N_4207);
or U4312 (N_4312,N_4266,N_4219);
nor U4313 (N_4313,N_4283,N_4294);
nand U4314 (N_4314,N_4242,N_4205);
and U4315 (N_4315,N_4268,N_4220);
and U4316 (N_4316,N_4208,N_4288);
nor U4317 (N_4317,N_4231,N_4267);
and U4318 (N_4318,N_4299,N_4241);
nor U4319 (N_4319,N_4264,N_4221);
or U4320 (N_4320,N_4232,N_4255);
or U4321 (N_4321,N_4285,N_4262);
or U4322 (N_4322,N_4280,N_4260);
nand U4323 (N_4323,N_4249,N_4278);
and U4324 (N_4324,N_4286,N_4217);
or U4325 (N_4325,N_4297,N_4236);
nor U4326 (N_4326,N_4227,N_4257);
or U4327 (N_4327,N_4256,N_4272);
xnor U4328 (N_4328,N_4295,N_4279);
nand U4329 (N_4329,N_4210,N_4298);
xnor U4330 (N_4330,N_4237,N_4204);
and U4331 (N_4331,N_4230,N_4216);
xnor U4332 (N_4332,N_4291,N_4203);
nand U4333 (N_4333,N_4201,N_4270);
and U4334 (N_4334,N_4218,N_4214);
or U4335 (N_4335,N_4277,N_4250);
nand U4336 (N_4336,N_4209,N_4202);
nand U4337 (N_4337,N_4251,N_4252);
or U4338 (N_4338,N_4223,N_4261);
and U4339 (N_4339,N_4240,N_4215);
and U4340 (N_4340,N_4282,N_4246);
nor U4341 (N_4341,N_4243,N_4292);
nor U4342 (N_4342,N_4239,N_4263);
and U4343 (N_4343,N_4287,N_4228);
nor U4344 (N_4344,N_4271,N_4212);
or U4345 (N_4345,N_4274,N_4281);
nor U4346 (N_4346,N_4269,N_4275);
and U4347 (N_4347,N_4248,N_4253);
and U4348 (N_4348,N_4225,N_4284);
and U4349 (N_4349,N_4290,N_4247);
nor U4350 (N_4350,N_4290,N_4241);
nand U4351 (N_4351,N_4289,N_4267);
or U4352 (N_4352,N_4277,N_4229);
or U4353 (N_4353,N_4237,N_4206);
and U4354 (N_4354,N_4258,N_4297);
nor U4355 (N_4355,N_4205,N_4223);
or U4356 (N_4356,N_4234,N_4290);
or U4357 (N_4357,N_4237,N_4238);
nor U4358 (N_4358,N_4208,N_4216);
or U4359 (N_4359,N_4270,N_4298);
nor U4360 (N_4360,N_4233,N_4232);
or U4361 (N_4361,N_4256,N_4252);
nor U4362 (N_4362,N_4263,N_4200);
or U4363 (N_4363,N_4235,N_4221);
xnor U4364 (N_4364,N_4276,N_4271);
and U4365 (N_4365,N_4274,N_4248);
or U4366 (N_4366,N_4204,N_4201);
and U4367 (N_4367,N_4288,N_4297);
and U4368 (N_4368,N_4275,N_4287);
or U4369 (N_4369,N_4223,N_4234);
or U4370 (N_4370,N_4280,N_4297);
or U4371 (N_4371,N_4236,N_4210);
nand U4372 (N_4372,N_4237,N_4281);
and U4373 (N_4373,N_4226,N_4230);
and U4374 (N_4374,N_4293,N_4228);
nor U4375 (N_4375,N_4215,N_4261);
nor U4376 (N_4376,N_4216,N_4204);
nor U4377 (N_4377,N_4216,N_4273);
or U4378 (N_4378,N_4221,N_4278);
nand U4379 (N_4379,N_4255,N_4266);
xor U4380 (N_4380,N_4292,N_4234);
nand U4381 (N_4381,N_4225,N_4238);
and U4382 (N_4382,N_4259,N_4212);
or U4383 (N_4383,N_4255,N_4268);
or U4384 (N_4384,N_4227,N_4236);
or U4385 (N_4385,N_4252,N_4289);
nor U4386 (N_4386,N_4230,N_4273);
and U4387 (N_4387,N_4249,N_4290);
nand U4388 (N_4388,N_4231,N_4259);
and U4389 (N_4389,N_4225,N_4268);
nand U4390 (N_4390,N_4247,N_4236);
and U4391 (N_4391,N_4218,N_4256);
and U4392 (N_4392,N_4291,N_4253);
nor U4393 (N_4393,N_4202,N_4248);
and U4394 (N_4394,N_4279,N_4297);
nor U4395 (N_4395,N_4224,N_4261);
nand U4396 (N_4396,N_4268,N_4233);
or U4397 (N_4397,N_4274,N_4225);
and U4398 (N_4398,N_4277,N_4243);
or U4399 (N_4399,N_4263,N_4255);
nor U4400 (N_4400,N_4352,N_4346);
nand U4401 (N_4401,N_4319,N_4312);
and U4402 (N_4402,N_4313,N_4316);
nand U4403 (N_4403,N_4358,N_4384);
nor U4404 (N_4404,N_4355,N_4343);
nor U4405 (N_4405,N_4324,N_4392);
and U4406 (N_4406,N_4367,N_4325);
nor U4407 (N_4407,N_4365,N_4336);
nand U4408 (N_4408,N_4318,N_4303);
nand U4409 (N_4409,N_4372,N_4305);
nor U4410 (N_4410,N_4301,N_4330);
or U4411 (N_4411,N_4393,N_4310);
and U4412 (N_4412,N_4321,N_4347);
nand U4413 (N_4413,N_4329,N_4380);
and U4414 (N_4414,N_4377,N_4370);
and U4415 (N_4415,N_4385,N_4338);
nand U4416 (N_4416,N_4311,N_4314);
nor U4417 (N_4417,N_4390,N_4383);
and U4418 (N_4418,N_4326,N_4306);
nand U4419 (N_4419,N_4317,N_4364);
or U4420 (N_4420,N_4375,N_4307);
or U4421 (N_4421,N_4361,N_4356);
xor U4422 (N_4422,N_4371,N_4320);
nand U4423 (N_4423,N_4353,N_4332);
or U4424 (N_4424,N_4348,N_4323);
or U4425 (N_4425,N_4335,N_4394);
or U4426 (N_4426,N_4333,N_4381);
and U4427 (N_4427,N_4396,N_4302);
nand U4428 (N_4428,N_4362,N_4351);
nor U4429 (N_4429,N_4345,N_4388);
and U4430 (N_4430,N_4315,N_4376);
and U4431 (N_4431,N_4349,N_4331);
nand U4432 (N_4432,N_4397,N_4340);
and U4433 (N_4433,N_4378,N_4387);
nor U4434 (N_4434,N_4337,N_4344);
nand U4435 (N_4435,N_4360,N_4386);
nor U4436 (N_4436,N_4322,N_4304);
or U4437 (N_4437,N_4339,N_4328);
nor U4438 (N_4438,N_4350,N_4369);
and U4439 (N_4439,N_4357,N_4363);
or U4440 (N_4440,N_4342,N_4374);
nand U4441 (N_4441,N_4368,N_4354);
nor U4442 (N_4442,N_4300,N_4399);
nand U4443 (N_4443,N_4379,N_4391);
nand U4444 (N_4444,N_4359,N_4382);
or U4445 (N_4445,N_4327,N_4334);
nor U4446 (N_4446,N_4398,N_4373);
and U4447 (N_4447,N_4395,N_4308);
nor U4448 (N_4448,N_4341,N_4366);
nand U4449 (N_4449,N_4389,N_4309);
or U4450 (N_4450,N_4304,N_4372);
and U4451 (N_4451,N_4381,N_4319);
and U4452 (N_4452,N_4311,N_4313);
nor U4453 (N_4453,N_4322,N_4398);
nor U4454 (N_4454,N_4315,N_4356);
nand U4455 (N_4455,N_4368,N_4382);
or U4456 (N_4456,N_4317,N_4335);
nand U4457 (N_4457,N_4386,N_4388);
nor U4458 (N_4458,N_4341,N_4349);
or U4459 (N_4459,N_4362,N_4356);
and U4460 (N_4460,N_4346,N_4310);
or U4461 (N_4461,N_4379,N_4396);
or U4462 (N_4462,N_4361,N_4347);
nand U4463 (N_4463,N_4314,N_4326);
nand U4464 (N_4464,N_4316,N_4367);
nor U4465 (N_4465,N_4342,N_4363);
nor U4466 (N_4466,N_4399,N_4311);
and U4467 (N_4467,N_4321,N_4346);
or U4468 (N_4468,N_4332,N_4322);
nor U4469 (N_4469,N_4364,N_4323);
or U4470 (N_4470,N_4370,N_4324);
nand U4471 (N_4471,N_4357,N_4328);
nor U4472 (N_4472,N_4336,N_4388);
or U4473 (N_4473,N_4313,N_4326);
or U4474 (N_4474,N_4333,N_4362);
and U4475 (N_4475,N_4367,N_4318);
nand U4476 (N_4476,N_4336,N_4392);
nand U4477 (N_4477,N_4361,N_4374);
and U4478 (N_4478,N_4352,N_4331);
nand U4479 (N_4479,N_4341,N_4384);
and U4480 (N_4480,N_4361,N_4333);
or U4481 (N_4481,N_4399,N_4359);
nand U4482 (N_4482,N_4339,N_4327);
nor U4483 (N_4483,N_4374,N_4351);
nor U4484 (N_4484,N_4341,N_4336);
and U4485 (N_4485,N_4339,N_4382);
or U4486 (N_4486,N_4370,N_4331);
nor U4487 (N_4487,N_4389,N_4357);
nand U4488 (N_4488,N_4342,N_4371);
and U4489 (N_4489,N_4365,N_4307);
or U4490 (N_4490,N_4385,N_4363);
nor U4491 (N_4491,N_4399,N_4365);
nor U4492 (N_4492,N_4383,N_4301);
or U4493 (N_4493,N_4394,N_4381);
nand U4494 (N_4494,N_4329,N_4320);
and U4495 (N_4495,N_4315,N_4347);
and U4496 (N_4496,N_4384,N_4396);
nand U4497 (N_4497,N_4307,N_4343);
nor U4498 (N_4498,N_4386,N_4311);
nor U4499 (N_4499,N_4391,N_4376);
nand U4500 (N_4500,N_4480,N_4408);
nand U4501 (N_4501,N_4417,N_4431);
or U4502 (N_4502,N_4494,N_4424);
nor U4503 (N_4503,N_4498,N_4497);
and U4504 (N_4504,N_4453,N_4435);
and U4505 (N_4505,N_4461,N_4443);
nand U4506 (N_4506,N_4439,N_4468);
or U4507 (N_4507,N_4401,N_4430);
and U4508 (N_4508,N_4416,N_4407);
nand U4509 (N_4509,N_4444,N_4495);
nor U4510 (N_4510,N_4462,N_4460);
and U4511 (N_4511,N_4485,N_4438);
nand U4512 (N_4512,N_4489,N_4436);
nand U4513 (N_4513,N_4486,N_4474);
and U4514 (N_4514,N_4456,N_4450);
or U4515 (N_4515,N_4484,N_4487);
or U4516 (N_4516,N_4429,N_4412);
or U4517 (N_4517,N_4469,N_4471);
nor U4518 (N_4518,N_4402,N_4413);
nor U4519 (N_4519,N_4477,N_4459);
xor U4520 (N_4520,N_4423,N_4420);
nor U4521 (N_4521,N_4454,N_4448);
or U4522 (N_4522,N_4479,N_4440);
and U4523 (N_4523,N_4437,N_4434);
nor U4524 (N_4524,N_4410,N_4496);
xor U4525 (N_4525,N_4473,N_4419);
nor U4526 (N_4526,N_4427,N_4481);
and U4527 (N_4527,N_4491,N_4432);
or U4528 (N_4528,N_4442,N_4446);
and U4529 (N_4529,N_4403,N_4451);
or U4530 (N_4530,N_4476,N_4478);
nor U4531 (N_4531,N_4488,N_4466);
nor U4532 (N_4532,N_4492,N_4470);
and U4533 (N_4533,N_4499,N_4483);
and U4534 (N_4534,N_4415,N_4421);
nor U4535 (N_4535,N_4452,N_4405);
or U4536 (N_4536,N_4441,N_4465);
nor U4537 (N_4537,N_4422,N_4493);
or U4538 (N_4538,N_4409,N_4411);
nor U4539 (N_4539,N_4404,N_4414);
xnor U4540 (N_4540,N_4418,N_4457);
or U4541 (N_4541,N_4458,N_4490);
nor U4542 (N_4542,N_4428,N_4426);
nand U4543 (N_4543,N_4472,N_4433);
and U4544 (N_4544,N_4475,N_4445);
and U4545 (N_4545,N_4467,N_4425);
nand U4546 (N_4546,N_4463,N_4447);
and U4547 (N_4547,N_4449,N_4482);
nand U4548 (N_4548,N_4406,N_4455);
or U4549 (N_4549,N_4464,N_4400);
and U4550 (N_4550,N_4499,N_4403);
nand U4551 (N_4551,N_4435,N_4456);
and U4552 (N_4552,N_4458,N_4429);
nor U4553 (N_4553,N_4495,N_4485);
nand U4554 (N_4554,N_4420,N_4410);
nand U4555 (N_4555,N_4497,N_4451);
and U4556 (N_4556,N_4439,N_4484);
or U4557 (N_4557,N_4406,N_4445);
and U4558 (N_4558,N_4493,N_4492);
or U4559 (N_4559,N_4408,N_4486);
nor U4560 (N_4560,N_4473,N_4437);
nor U4561 (N_4561,N_4483,N_4417);
nor U4562 (N_4562,N_4457,N_4440);
nand U4563 (N_4563,N_4432,N_4463);
nor U4564 (N_4564,N_4441,N_4484);
nor U4565 (N_4565,N_4421,N_4428);
nor U4566 (N_4566,N_4465,N_4488);
nand U4567 (N_4567,N_4477,N_4452);
or U4568 (N_4568,N_4476,N_4414);
or U4569 (N_4569,N_4406,N_4403);
and U4570 (N_4570,N_4447,N_4423);
and U4571 (N_4571,N_4491,N_4408);
nor U4572 (N_4572,N_4432,N_4408);
nand U4573 (N_4573,N_4479,N_4418);
and U4574 (N_4574,N_4484,N_4433);
nor U4575 (N_4575,N_4427,N_4465);
or U4576 (N_4576,N_4454,N_4469);
nor U4577 (N_4577,N_4475,N_4488);
or U4578 (N_4578,N_4425,N_4411);
nand U4579 (N_4579,N_4498,N_4414);
or U4580 (N_4580,N_4406,N_4439);
and U4581 (N_4581,N_4476,N_4477);
nand U4582 (N_4582,N_4445,N_4450);
or U4583 (N_4583,N_4429,N_4448);
or U4584 (N_4584,N_4498,N_4482);
and U4585 (N_4585,N_4449,N_4474);
or U4586 (N_4586,N_4495,N_4429);
nor U4587 (N_4587,N_4480,N_4405);
nand U4588 (N_4588,N_4427,N_4493);
and U4589 (N_4589,N_4497,N_4419);
and U4590 (N_4590,N_4445,N_4489);
nor U4591 (N_4591,N_4460,N_4441);
nand U4592 (N_4592,N_4417,N_4495);
or U4593 (N_4593,N_4421,N_4491);
or U4594 (N_4594,N_4482,N_4463);
nand U4595 (N_4595,N_4474,N_4405);
nor U4596 (N_4596,N_4489,N_4463);
nor U4597 (N_4597,N_4459,N_4413);
or U4598 (N_4598,N_4444,N_4499);
or U4599 (N_4599,N_4420,N_4491);
and U4600 (N_4600,N_4509,N_4592);
nand U4601 (N_4601,N_4566,N_4501);
or U4602 (N_4602,N_4560,N_4525);
and U4603 (N_4603,N_4517,N_4543);
nor U4604 (N_4604,N_4521,N_4503);
or U4605 (N_4605,N_4565,N_4550);
or U4606 (N_4606,N_4529,N_4570);
and U4607 (N_4607,N_4573,N_4526);
or U4608 (N_4608,N_4545,N_4588);
and U4609 (N_4609,N_4541,N_4534);
xor U4610 (N_4610,N_4564,N_4513);
nand U4611 (N_4611,N_4516,N_4581);
nand U4612 (N_4612,N_4551,N_4585);
and U4613 (N_4613,N_4555,N_4510);
or U4614 (N_4614,N_4532,N_4538);
or U4615 (N_4615,N_4589,N_4522);
nor U4616 (N_4616,N_4531,N_4562);
and U4617 (N_4617,N_4500,N_4552);
nand U4618 (N_4618,N_4559,N_4515);
and U4619 (N_4619,N_4511,N_4549);
nand U4620 (N_4620,N_4548,N_4533);
or U4621 (N_4621,N_4583,N_4558);
and U4622 (N_4622,N_4504,N_4567);
or U4623 (N_4623,N_4553,N_4544);
nor U4624 (N_4624,N_4575,N_4508);
nor U4625 (N_4625,N_4556,N_4547);
nor U4626 (N_4626,N_4536,N_4530);
or U4627 (N_4627,N_4502,N_4586);
nand U4628 (N_4628,N_4540,N_4596);
and U4629 (N_4629,N_4582,N_4594);
nor U4630 (N_4630,N_4563,N_4593);
nor U4631 (N_4631,N_4554,N_4527);
nor U4632 (N_4632,N_4590,N_4579);
nand U4633 (N_4633,N_4505,N_4524);
and U4634 (N_4634,N_4537,N_4557);
or U4635 (N_4635,N_4519,N_4506);
nor U4636 (N_4636,N_4535,N_4597);
nand U4637 (N_4637,N_4584,N_4514);
or U4638 (N_4638,N_4561,N_4539);
nor U4639 (N_4639,N_4518,N_4578);
nor U4640 (N_4640,N_4599,N_4528);
nand U4641 (N_4641,N_4512,N_4568);
nor U4642 (N_4642,N_4542,N_4546);
and U4643 (N_4643,N_4580,N_4595);
and U4644 (N_4644,N_4520,N_4507);
and U4645 (N_4645,N_4591,N_4574);
and U4646 (N_4646,N_4572,N_4523);
nor U4647 (N_4647,N_4587,N_4598);
nor U4648 (N_4648,N_4571,N_4577);
nor U4649 (N_4649,N_4569,N_4576);
nor U4650 (N_4650,N_4514,N_4529);
and U4651 (N_4651,N_4548,N_4531);
nor U4652 (N_4652,N_4515,N_4561);
and U4653 (N_4653,N_4525,N_4545);
and U4654 (N_4654,N_4510,N_4574);
or U4655 (N_4655,N_4553,N_4554);
and U4656 (N_4656,N_4540,N_4543);
nor U4657 (N_4657,N_4552,N_4569);
nand U4658 (N_4658,N_4545,N_4560);
and U4659 (N_4659,N_4585,N_4501);
nand U4660 (N_4660,N_4581,N_4532);
nor U4661 (N_4661,N_4510,N_4506);
or U4662 (N_4662,N_4509,N_4533);
and U4663 (N_4663,N_4554,N_4532);
nand U4664 (N_4664,N_4593,N_4546);
nand U4665 (N_4665,N_4570,N_4548);
nand U4666 (N_4666,N_4555,N_4546);
and U4667 (N_4667,N_4591,N_4505);
nor U4668 (N_4668,N_4552,N_4576);
nor U4669 (N_4669,N_4527,N_4552);
nor U4670 (N_4670,N_4579,N_4507);
nor U4671 (N_4671,N_4504,N_4595);
nand U4672 (N_4672,N_4566,N_4592);
nand U4673 (N_4673,N_4502,N_4555);
or U4674 (N_4674,N_4577,N_4570);
nand U4675 (N_4675,N_4552,N_4504);
nor U4676 (N_4676,N_4500,N_4513);
nand U4677 (N_4677,N_4556,N_4532);
nor U4678 (N_4678,N_4575,N_4513);
and U4679 (N_4679,N_4566,N_4505);
nand U4680 (N_4680,N_4555,N_4519);
nor U4681 (N_4681,N_4522,N_4527);
nand U4682 (N_4682,N_4551,N_4559);
nand U4683 (N_4683,N_4535,N_4501);
or U4684 (N_4684,N_4577,N_4532);
nand U4685 (N_4685,N_4515,N_4575);
nor U4686 (N_4686,N_4597,N_4543);
nor U4687 (N_4687,N_4595,N_4585);
nor U4688 (N_4688,N_4530,N_4587);
nor U4689 (N_4689,N_4558,N_4568);
nand U4690 (N_4690,N_4583,N_4595);
nor U4691 (N_4691,N_4537,N_4577);
nand U4692 (N_4692,N_4582,N_4523);
nor U4693 (N_4693,N_4562,N_4597);
nand U4694 (N_4694,N_4501,N_4561);
nor U4695 (N_4695,N_4597,N_4560);
nand U4696 (N_4696,N_4588,N_4569);
nor U4697 (N_4697,N_4573,N_4522);
nand U4698 (N_4698,N_4586,N_4504);
nor U4699 (N_4699,N_4541,N_4515);
nor U4700 (N_4700,N_4613,N_4661);
nor U4701 (N_4701,N_4696,N_4663);
and U4702 (N_4702,N_4607,N_4614);
and U4703 (N_4703,N_4612,N_4640);
or U4704 (N_4704,N_4645,N_4606);
nand U4705 (N_4705,N_4652,N_4671);
and U4706 (N_4706,N_4632,N_4610);
nor U4707 (N_4707,N_4649,N_4697);
and U4708 (N_4708,N_4694,N_4679);
xnor U4709 (N_4709,N_4600,N_4617);
nor U4710 (N_4710,N_4686,N_4668);
and U4711 (N_4711,N_4665,N_4626);
or U4712 (N_4712,N_4627,N_4689);
or U4713 (N_4713,N_4654,N_4620);
nand U4714 (N_4714,N_4664,N_4644);
or U4715 (N_4715,N_4621,N_4630);
and U4716 (N_4716,N_4646,N_4682);
nor U4717 (N_4717,N_4636,N_4660);
and U4718 (N_4718,N_4615,N_4639);
nand U4719 (N_4719,N_4603,N_4670);
nand U4720 (N_4720,N_4651,N_4692);
or U4721 (N_4721,N_4690,N_4631);
and U4722 (N_4722,N_4623,N_4688);
nor U4723 (N_4723,N_4658,N_4666);
nand U4724 (N_4724,N_4662,N_4619);
and U4725 (N_4725,N_4655,N_4698);
or U4726 (N_4726,N_4678,N_4681);
and U4727 (N_4727,N_4624,N_4602);
or U4728 (N_4728,N_4673,N_4611);
or U4729 (N_4729,N_4667,N_4643);
nand U4730 (N_4730,N_4672,N_4683);
and U4731 (N_4731,N_4635,N_4691);
nor U4732 (N_4732,N_4601,N_4608);
and U4733 (N_4733,N_4625,N_4669);
nor U4734 (N_4734,N_4677,N_4629);
nand U4735 (N_4735,N_4650,N_4638);
or U4736 (N_4736,N_4637,N_4687);
and U4737 (N_4737,N_4693,N_4699);
nor U4738 (N_4738,N_4628,N_4674);
or U4739 (N_4739,N_4648,N_4684);
nor U4740 (N_4740,N_4622,N_4676);
and U4741 (N_4741,N_4653,N_4609);
and U4742 (N_4742,N_4656,N_4680);
nor U4743 (N_4743,N_4641,N_4618);
nor U4744 (N_4744,N_4604,N_4659);
xor U4745 (N_4745,N_4605,N_4657);
nor U4746 (N_4746,N_4695,N_4647);
and U4747 (N_4747,N_4675,N_4634);
nand U4748 (N_4748,N_4685,N_4616);
nand U4749 (N_4749,N_4642,N_4633);
and U4750 (N_4750,N_4676,N_4695);
nor U4751 (N_4751,N_4634,N_4604);
nor U4752 (N_4752,N_4610,N_4626);
nor U4753 (N_4753,N_4697,N_4620);
nor U4754 (N_4754,N_4647,N_4666);
or U4755 (N_4755,N_4671,N_4611);
xor U4756 (N_4756,N_4629,N_4630);
and U4757 (N_4757,N_4624,N_4632);
or U4758 (N_4758,N_4664,N_4662);
and U4759 (N_4759,N_4692,N_4697);
or U4760 (N_4760,N_4660,N_4629);
nor U4761 (N_4761,N_4609,N_4642);
and U4762 (N_4762,N_4664,N_4689);
nor U4763 (N_4763,N_4642,N_4641);
nor U4764 (N_4764,N_4602,N_4671);
or U4765 (N_4765,N_4622,N_4697);
and U4766 (N_4766,N_4620,N_4695);
nor U4767 (N_4767,N_4622,N_4635);
or U4768 (N_4768,N_4617,N_4699);
and U4769 (N_4769,N_4605,N_4612);
and U4770 (N_4770,N_4644,N_4687);
and U4771 (N_4771,N_4606,N_4635);
or U4772 (N_4772,N_4695,N_4662);
and U4773 (N_4773,N_4644,N_4699);
and U4774 (N_4774,N_4639,N_4643);
or U4775 (N_4775,N_4638,N_4675);
or U4776 (N_4776,N_4673,N_4632);
nand U4777 (N_4777,N_4611,N_4685);
or U4778 (N_4778,N_4603,N_4698);
and U4779 (N_4779,N_4680,N_4604);
and U4780 (N_4780,N_4602,N_4647);
and U4781 (N_4781,N_4680,N_4686);
nor U4782 (N_4782,N_4642,N_4651);
nor U4783 (N_4783,N_4697,N_4611);
nand U4784 (N_4784,N_4637,N_4646);
xor U4785 (N_4785,N_4696,N_4669);
or U4786 (N_4786,N_4625,N_4667);
nand U4787 (N_4787,N_4665,N_4645);
nand U4788 (N_4788,N_4664,N_4622);
or U4789 (N_4789,N_4604,N_4623);
nor U4790 (N_4790,N_4627,N_4603);
nand U4791 (N_4791,N_4646,N_4677);
and U4792 (N_4792,N_4620,N_4606);
and U4793 (N_4793,N_4630,N_4622);
nor U4794 (N_4794,N_4656,N_4654);
or U4795 (N_4795,N_4695,N_4684);
and U4796 (N_4796,N_4612,N_4677);
or U4797 (N_4797,N_4657,N_4666);
or U4798 (N_4798,N_4627,N_4628);
and U4799 (N_4799,N_4679,N_4685);
and U4800 (N_4800,N_4750,N_4708);
and U4801 (N_4801,N_4794,N_4784);
nor U4802 (N_4802,N_4762,N_4776);
and U4803 (N_4803,N_4753,N_4755);
nand U4804 (N_4804,N_4702,N_4733);
and U4805 (N_4805,N_4731,N_4769);
nor U4806 (N_4806,N_4775,N_4780);
nand U4807 (N_4807,N_4779,N_4742);
nor U4808 (N_4808,N_4746,N_4735);
or U4809 (N_4809,N_4715,N_4730);
and U4810 (N_4810,N_4754,N_4752);
nand U4811 (N_4811,N_4707,N_4738);
and U4812 (N_4812,N_4777,N_4714);
xnor U4813 (N_4813,N_4744,N_4797);
and U4814 (N_4814,N_4796,N_4717);
nor U4815 (N_4815,N_4791,N_4761);
nand U4816 (N_4816,N_4725,N_4700);
and U4817 (N_4817,N_4736,N_4795);
nand U4818 (N_4818,N_4745,N_4758);
or U4819 (N_4819,N_4721,N_4792);
or U4820 (N_4820,N_4728,N_4701);
and U4821 (N_4821,N_4766,N_4704);
nand U4822 (N_4822,N_4782,N_4787);
nand U4823 (N_4823,N_4747,N_4741);
and U4824 (N_4824,N_4798,N_4773);
or U4825 (N_4825,N_4749,N_4719);
or U4826 (N_4826,N_4759,N_4726);
or U4827 (N_4827,N_4722,N_4768);
nand U4828 (N_4828,N_4778,N_4743);
or U4829 (N_4829,N_4757,N_4770);
nand U4830 (N_4830,N_4799,N_4789);
nor U4831 (N_4831,N_4712,N_4774);
or U4832 (N_4832,N_4703,N_4711);
or U4833 (N_4833,N_4720,N_4786);
nand U4834 (N_4834,N_4748,N_4713);
and U4835 (N_4835,N_4790,N_4751);
nor U4836 (N_4836,N_4732,N_4760);
nand U4837 (N_4837,N_4737,N_4756);
or U4838 (N_4838,N_4729,N_4709);
and U4839 (N_4839,N_4727,N_4710);
and U4840 (N_4840,N_4788,N_4705);
and U4841 (N_4841,N_4740,N_4783);
nand U4842 (N_4842,N_4764,N_4723);
nor U4843 (N_4843,N_4781,N_4734);
nor U4844 (N_4844,N_4771,N_4716);
nor U4845 (N_4845,N_4706,N_4765);
and U4846 (N_4846,N_4763,N_4767);
or U4847 (N_4847,N_4785,N_4772);
nor U4848 (N_4848,N_4724,N_4739);
or U4849 (N_4849,N_4793,N_4718);
and U4850 (N_4850,N_4708,N_4714);
xnor U4851 (N_4851,N_4768,N_4739);
nor U4852 (N_4852,N_4781,N_4749);
and U4853 (N_4853,N_4767,N_4778);
or U4854 (N_4854,N_4715,N_4709);
nand U4855 (N_4855,N_4756,N_4745);
and U4856 (N_4856,N_4740,N_4743);
nand U4857 (N_4857,N_4717,N_4780);
nand U4858 (N_4858,N_4728,N_4761);
nor U4859 (N_4859,N_4736,N_4789);
or U4860 (N_4860,N_4787,N_4705);
or U4861 (N_4861,N_4769,N_4788);
or U4862 (N_4862,N_4778,N_4798);
and U4863 (N_4863,N_4738,N_4769);
or U4864 (N_4864,N_4787,N_4763);
or U4865 (N_4865,N_4715,N_4727);
or U4866 (N_4866,N_4791,N_4759);
and U4867 (N_4867,N_4776,N_4793);
nor U4868 (N_4868,N_4772,N_4711);
nor U4869 (N_4869,N_4711,N_4783);
or U4870 (N_4870,N_4741,N_4723);
nor U4871 (N_4871,N_4764,N_4727);
and U4872 (N_4872,N_4700,N_4752);
nor U4873 (N_4873,N_4732,N_4754);
nand U4874 (N_4874,N_4707,N_4743);
or U4875 (N_4875,N_4758,N_4734);
nor U4876 (N_4876,N_4719,N_4708);
nor U4877 (N_4877,N_4758,N_4718);
nand U4878 (N_4878,N_4790,N_4786);
or U4879 (N_4879,N_4743,N_4796);
nor U4880 (N_4880,N_4756,N_4769);
and U4881 (N_4881,N_4791,N_4796);
or U4882 (N_4882,N_4751,N_4705);
nand U4883 (N_4883,N_4784,N_4753);
nand U4884 (N_4884,N_4793,N_4745);
and U4885 (N_4885,N_4744,N_4751);
nor U4886 (N_4886,N_4741,N_4707);
and U4887 (N_4887,N_4774,N_4744);
and U4888 (N_4888,N_4718,N_4732);
nand U4889 (N_4889,N_4725,N_4722);
nor U4890 (N_4890,N_4711,N_4786);
nand U4891 (N_4891,N_4727,N_4713);
xnor U4892 (N_4892,N_4756,N_4743);
nand U4893 (N_4893,N_4762,N_4733);
and U4894 (N_4894,N_4781,N_4759);
nor U4895 (N_4895,N_4734,N_4723);
nand U4896 (N_4896,N_4740,N_4757);
nor U4897 (N_4897,N_4701,N_4781);
or U4898 (N_4898,N_4776,N_4748);
nor U4899 (N_4899,N_4785,N_4732);
and U4900 (N_4900,N_4882,N_4801);
nand U4901 (N_4901,N_4848,N_4847);
nor U4902 (N_4902,N_4863,N_4898);
nor U4903 (N_4903,N_4852,N_4876);
and U4904 (N_4904,N_4851,N_4850);
nor U4905 (N_4905,N_4893,N_4812);
nor U4906 (N_4906,N_4872,N_4888);
and U4907 (N_4907,N_4892,N_4861);
and U4908 (N_4908,N_4871,N_4811);
and U4909 (N_4909,N_4835,N_4891);
or U4910 (N_4910,N_4829,N_4849);
or U4911 (N_4911,N_4844,N_4856);
or U4912 (N_4912,N_4808,N_4804);
nand U4913 (N_4913,N_4837,N_4867);
nand U4914 (N_4914,N_4862,N_4884);
or U4915 (N_4915,N_4827,N_4890);
or U4916 (N_4916,N_4825,N_4886);
nor U4917 (N_4917,N_4896,N_4815);
nor U4918 (N_4918,N_4805,N_4806);
nor U4919 (N_4919,N_4819,N_4834);
and U4920 (N_4920,N_4887,N_4866);
and U4921 (N_4921,N_4869,N_4878);
and U4922 (N_4922,N_4889,N_4836);
or U4923 (N_4923,N_4874,N_4858);
or U4924 (N_4924,N_4838,N_4857);
or U4925 (N_4925,N_4859,N_4883);
and U4926 (N_4926,N_4899,N_4807);
or U4927 (N_4927,N_4875,N_4897);
nand U4928 (N_4928,N_4845,N_4841);
or U4929 (N_4929,N_4870,N_4809);
and U4930 (N_4930,N_4813,N_4877);
nand U4931 (N_4931,N_4879,N_4823);
or U4932 (N_4932,N_4803,N_4868);
and U4933 (N_4933,N_4830,N_4839);
nor U4934 (N_4934,N_4826,N_4853);
or U4935 (N_4935,N_4816,N_4833);
nor U4936 (N_4936,N_4873,N_4810);
nor U4937 (N_4937,N_4818,N_4843);
or U4938 (N_4938,N_4817,N_4860);
nor U4939 (N_4939,N_4895,N_4842);
or U4940 (N_4940,N_4881,N_4802);
nand U4941 (N_4941,N_4822,N_4854);
and U4942 (N_4942,N_4840,N_4800);
nand U4943 (N_4943,N_4865,N_4821);
nand U4944 (N_4944,N_4828,N_4824);
nor U4945 (N_4945,N_4880,N_4894);
and U4946 (N_4946,N_4832,N_4846);
nand U4947 (N_4947,N_4885,N_4831);
nand U4948 (N_4948,N_4814,N_4864);
and U4949 (N_4949,N_4855,N_4820);
nor U4950 (N_4950,N_4876,N_4840);
nand U4951 (N_4951,N_4868,N_4867);
nor U4952 (N_4952,N_4810,N_4850);
and U4953 (N_4953,N_4851,N_4840);
nand U4954 (N_4954,N_4816,N_4898);
nand U4955 (N_4955,N_4835,N_4827);
nand U4956 (N_4956,N_4816,N_4887);
or U4957 (N_4957,N_4825,N_4882);
or U4958 (N_4958,N_4800,N_4848);
nand U4959 (N_4959,N_4818,N_4809);
nand U4960 (N_4960,N_4818,N_4835);
or U4961 (N_4961,N_4888,N_4826);
and U4962 (N_4962,N_4870,N_4800);
nand U4963 (N_4963,N_4825,N_4829);
or U4964 (N_4964,N_4800,N_4866);
or U4965 (N_4965,N_4848,N_4819);
or U4966 (N_4966,N_4895,N_4886);
and U4967 (N_4967,N_4856,N_4896);
nor U4968 (N_4968,N_4860,N_4845);
or U4969 (N_4969,N_4887,N_4885);
and U4970 (N_4970,N_4820,N_4890);
nand U4971 (N_4971,N_4815,N_4887);
or U4972 (N_4972,N_4895,N_4814);
nand U4973 (N_4973,N_4893,N_4800);
nand U4974 (N_4974,N_4855,N_4877);
or U4975 (N_4975,N_4852,N_4865);
or U4976 (N_4976,N_4850,N_4831);
nor U4977 (N_4977,N_4836,N_4820);
nand U4978 (N_4978,N_4881,N_4896);
nand U4979 (N_4979,N_4865,N_4875);
and U4980 (N_4980,N_4815,N_4808);
nor U4981 (N_4981,N_4872,N_4853);
or U4982 (N_4982,N_4862,N_4824);
and U4983 (N_4983,N_4803,N_4828);
nand U4984 (N_4984,N_4834,N_4868);
and U4985 (N_4985,N_4833,N_4835);
nor U4986 (N_4986,N_4845,N_4808);
and U4987 (N_4987,N_4894,N_4891);
nor U4988 (N_4988,N_4897,N_4818);
and U4989 (N_4989,N_4899,N_4850);
nor U4990 (N_4990,N_4896,N_4878);
nor U4991 (N_4991,N_4895,N_4812);
and U4992 (N_4992,N_4870,N_4802);
nor U4993 (N_4993,N_4868,N_4802);
or U4994 (N_4994,N_4870,N_4880);
and U4995 (N_4995,N_4849,N_4807);
and U4996 (N_4996,N_4870,N_4883);
and U4997 (N_4997,N_4802,N_4838);
nor U4998 (N_4998,N_4841,N_4879);
nand U4999 (N_4999,N_4879,N_4815);
xor U5000 (N_5000,N_4994,N_4966);
or U5001 (N_5001,N_4998,N_4995);
nand U5002 (N_5002,N_4937,N_4972);
and U5003 (N_5003,N_4952,N_4971);
xor U5004 (N_5004,N_4960,N_4936);
or U5005 (N_5005,N_4997,N_4919);
nand U5006 (N_5006,N_4955,N_4976);
or U5007 (N_5007,N_4922,N_4949);
or U5008 (N_5008,N_4991,N_4904);
and U5009 (N_5009,N_4905,N_4988);
and U5010 (N_5010,N_4987,N_4929);
or U5011 (N_5011,N_4915,N_4957);
or U5012 (N_5012,N_4969,N_4975);
nand U5013 (N_5013,N_4942,N_4916);
or U5014 (N_5014,N_4990,N_4903);
or U5015 (N_5015,N_4909,N_4931);
and U5016 (N_5016,N_4950,N_4918);
and U5017 (N_5017,N_4963,N_4978);
or U5018 (N_5018,N_4947,N_4927);
nor U5019 (N_5019,N_4934,N_4928);
xor U5020 (N_5020,N_4953,N_4911);
or U5021 (N_5021,N_4958,N_4962);
or U5022 (N_5022,N_4984,N_4940);
and U5023 (N_5023,N_4970,N_4943);
or U5024 (N_5024,N_4906,N_4954);
nand U5025 (N_5025,N_4992,N_4935);
xor U5026 (N_5026,N_4946,N_4967);
and U5027 (N_5027,N_4923,N_4996);
and U5028 (N_5028,N_4917,N_4956);
or U5029 (N_5029,N_4932,N_4982);
nor U5030 (N_5030,N_4985,N_4980);
nand U5031 (N_5031,N_4951,N_4921);
and U5032 (N_5032,N_4907,N_4910);
nor U5033 (N_5033,N_4941,N_4933);
nor U5034 (N_5034,N_4979,N_4913);
and U5035 (N_5035,N_4930,N_4914);
nor U5036 (N_5036,N_4961,N_4901);
and U5037 (N_5037,N_4908,N_4945);
or U5038 (N_5038,N_4974,N_4900);
nand U5039 (N_5039,N_4965,N_4999);
nor U5040 (N_5040,N_4977,N_4981);
nand U5041 (N_5041,N_4948,N_4986);
or U5042 (N_5042,N_4989,N_4964);
nor U5043 (N_5043,N_4902,N_4993);
nand U5044 (N_5044,N_4968,N_4959);
and U5045 (N_5045,N_4939,N_4926);
nand U5046 (N_5046,N_4944,N_4920);
or U5047 (N_5047,N_4924,N_4925);
or U5048 (N_5048,N_4973,N_4983);
nand U5049 (N_5049,N_4912,N_4938);
nor U5050 (N_5050,N_4928,N_4937);
and U5051 (N_5051,N_4959,N_4962);
nand U5052 (N_5052,N_4966,N_4906);
or U5053 (N_5053,N_4954,N_4947);
nand U5054 (N_5054,N_4969,N_4964);
nor U5055 (N_5055,N_4916,N_4953);
or U5056 (N_5056,N_4965,N_4968);
or U5057 (N_5057,N_4909,N_4976);
nand U5058 (N_5058,N_4932,N_4934);
nor U5059 (N_5059,N_4979,N_4922);
nand U5060 (N_5060,N_4936,N_4940);
nor U5061 (N_5061,N_4974,N_4924);
or U5062 (N_5062,N_4933,N_4970);
or U5063 (N_5063,N_4936,N_4922);
or U5064 (N_5064,N_4921,N_4963);
nor U5065 (N_5065,N_4937,N_4989);
nor U5066 (N_5066,N_4974,N_4946);
or U5067 (N_5067,N_4959,N_4966);
or U5068 (N_5068,N_4977,N_4980);
nand U5069 (N_5069,N_4944,N_4998);
and U5070 (N_5070,N_4986,N_4971);
and U5071 (N_5071,N_4911,N_4926);
or U5072 (N_5072,N_4971,N_4999);
and U5073 (N_5073,N_4939,N_4982);
and U5074 (N_5074,N_4979,N_4905);
and U5075 (N_5075,N_4973,N_4900);
nor U5076 (N_5076,N_4923,N_4969);
nand U5077 (N_5077,N_4947,N_4919);
and U5078 (N_5078,N_4915,N_4934);
and U5079 (N_5079,N_4914,N_4978);
nand U5080 (N_5080,N_4981,N_4903);
or U5081 (N_5081,N_4985,N_4992);
or U5082 (N_5082,N_4915,N_4941);
or U5083 (N_5083,N_4979,N_4940);
and U5084 (N_5084,N_4911,N_4959);
nor U5085 (N_5085,N_4937,N_4921);
or U5086 (N_5086,N_4951,N_4926);
nand U5087 (N_5087,N_4914,N_4993);
nor U5088 (N_5088,N_4936,N_4979);
nand U5089 (N_5089,N_4980,N_4953);
nor U5090 (N_5090,N_4932,N_4917);
and U5091 (N_5091,N_4953,N_4928);
nand U5092 (N_5092,N_4988,N_4928);
nand U5093 (N_5093,N_4982,N_4981);
or U5094 (N_5094,N_4945,N_4966);
nor U5095 (N_5095,N_4942,N_4985);
nand U5096 (N_5096,N_4992,N_4903);
and U5097 (N_5097,N_4996,N_4967);
nand U5098 (N_5098,N_4921,N_4938);
or U5099 (N_5099,N_4995,N_4910);
nand U5100 (N_5100,N_5079,N_5015);
nor U5101 (N_5101,N_5021,N_5084);
or U5102 (N_5102,N_5075,N_5011);
nand U5103 (N_5103,N_5053,N_5002);
xor U5104 (N_5104,N_5070,N_5001);
nor U5105 (N_5105,N_5033,N_5018);
nand U5106 (N_5106,N_5067,N_5058);
nand U5107 (N_5107,N_5099,N_5046);
nor U5108 (N_5108,N_5041,N_5069);
nand U5109 (N_5109,N_5036,N_5062);
nand U5110 (N_5110,N_5071,N_5095);
or U5111 (N_5111,N_5048,N_5056);
nand U5112 (N_5112,N_5030,N_5078);
and U5113 (N_5113,N_5020,N_5073);
nor U5114 (N_5114,N_5022,N_5064);
or U5115 (N_5115,N_5019,N_5038);
nor U5116 (N_5116,N_5098,N_5066);
nand U5117 (N_5117,N_5094,N_5081);
nor U5118 (N_5118,N_5010,N_5080);
or U5119 (N_5119,N_5052,N_5047);
and U5120 (N_5120,N_5037,N_5072);
or U5121 (N_5121,N_5082,N_5083);
and U5122 (N_5122,N_5027,N_5032);
nor U5123 (N_5123,N_5004,N_5013);
nor U5124 (N_5124,N_5074,N_5025);
nor U5125 (N_5125,N_5063,N_5049);
or U5126 (N_5126,N_5003,N_5097);
or U5127 (N_5127,N_5028,N_5024);
nand U5128 (N_5128,N_5068,N_5088);
nor U5129 (N_5129,N_5008,N_5050);
nor U5130 (N_5130,N_5085,N_5065);
nor U5131 (N_5131,N_5059,N_5000);
nand U5132 (N_5132,N_5086,N_5043);
or U5133 (N_5133,N_5016,N_5093);
nand U5134 (N_5134,N_5034,N_5017);
and U5135 (N_5135,N_5055,N_5089);
nand U5136 (N_5136,N_5006,N_5023);
and U5137 (N_5137,N_5007,N_5012);
and U5138 (N_5138,N_5040,N_5045);
xnor U5139 (N_5139,N_5061,N_5092);
nor U5140 (N_5140,N_5031,N_5051);
nand U5141 (N_5141,N_5026,N_5042);
nor U5142 (N_5142,N_5087,N_5076);
nand U5143 (N_5143,N_5057,N_5014);
nor U5144 (N_5144,N_5009,N_5005);
or U5145 (N_5145,N_5096,N_5044);
or U5146 (N_5146,N_5077,N_5029);
and U5147 (N_5147,N_5060,N_5035);
and U5148 (N_5148,N_5054,N_5090);
and U5149 (N_5149,N_5039,N_5091);
or U5150 (N_5150,N_5017,N_5071);
and U5151 (N_5151,N_5094,N_5059);
nand U5152 (N_5152,N_5027,N_5000);
and U5153 (N_5153,N_5041,N_5014);
and U5154 (N_5154,N_5068,N_5053);
nor U5155 (N_5155,N_5050,N_5047);
and U5156 (N_5156,N_5021,N_5044);
and U5157 (N_5157,N_5000,N_5039);
and U5158 (N_5158,N_5026,N_5054);
nand U5159 (N_5159,N_5021,N_5015);
or U5160 (N_5160,N_5080,N_5044);
nand U5161 (N_5161,N_5063,N_5092);
and U5162 (N_5162,N_5044,N_5055);
nand U5163 (N_5163,N_5092,N_5089);
or U5164 (N_5164,N_5048,N_5093);
nor U5165 (N_5165,N_5021,N_5010);
and U5166 (N_5166,N_5071,N_5081);
and U5167 (N_5167,N_5046,N_5094);
or U5168 (N_5168,N_5013,N_5003);
and U5169 (N_5169,N_5014,N_5065);
or U5170 (N_5170,N_5078,N_5011);
nand U5171 (N_5171,N_5077,N_5059);
nand U5172 (N_5172,N_5066,N_5071);
nor U5173 (N_5173,N_5086,N_5013);
or U5174 (N_5174,N_5061,N_5027);
and U5175 (N_5175,N_5072,N_5029);
or U5176 (N_5176,N_5039,N_5083);
nor U5177 (N_5177,N_5002,N_5003);
nand U5178 (N_5178,N_5080,N_5045);
nand U5179 (N_5179,N_5045,N_5029);
nand U5180 (N_5180,N_5024,N_5020);
nand U5181 (N_5181,N_5016,N_5084);
nand U5182 (N_5182,N_5021,N_5048);
and U5183 (N_5183,N_5019,N_5078);
xnor U5184 (N_5184,N_5072,N_5075);
nand U5185 (N_5185,N_5046,N_5001);
nor U5186 (N_5186,N_5064,N_5074);
nor U5187 (N_5187,N_5099,N_5067);
or U5188 (N_5188,N_5088,N_5035);
and U5189 (N_5189,N_5040,N_5006);
nand U5190 (N_5190,N_5011,N_5082);
nor U5191 (N_5191,N_5081,N_5037);
and U5192 (N_5192,N_5033,N_5009);
and U5193 (N_5193,N_5007,N_5018);
nand U5194 (N_5194,N_5071,N_5048);
nor U5195 (N_5195,N_5013,N_5079);
nor U5196 (N_5196,N_5040,N_5048);
and U5197 (N_5197,N_5068,N_5033);
nand U5198 (N_5198,N_5095,N_5000);
nand U5199 (N_5199,N_5052,N_5017);
or U5200 (N_5200,N_5112,N_5174);
nor U5201 (N_5201,N_5133,N_5182);
or U5202 (N_5202,N_5170,N_5142);
nand U5203 (N_5203,N_5162,N_5199);
and U5204 (N_5204,N_5197,N_5181);
and U5205 (N_5205,N_5189,N_5149);
and U5206 (N_5206,N_5163,N_5137);
or U5207 (N_5207,N_5136,N_5126);
nand U5208 (N_5208,N_5131,N_5140);
and U5209 (N_5209,N_5100,N_5184);
and U5210 (N_5210,N_5129,N_5195);
and U5211 (N_5211,N_5151,N_5108);
nor U5212 (N_5212,N_5138,N_5168);
or U5213 (N_5213,N_5115,N_5121);
and U5214 (N_5214,N_5193,N_5190);
nand U5215 (N_5215,N_5175,N_5183);
or U5216 (N_5216,N_5132,N_5110);
nand U5217 (N_5217,N_5166,N_5143);
or U5218 (N_5218,N_5188,N_5116);
and U5219 (N_5219,N_5134,N_5164);
or U5220 (N_5220,N_5160,N_5111);
or U5221 (N_5221,N_5153,N_5147);
or U5222 (N_5222,N_5145,N_5104);
nand U5223 (N_5223,N_5186,N_5155);
or U5224 (N_5224,N_5173,N_5130);
nand U5225 (N_5225,N_5109,N_5122);
and U5226 (N_5226,N_5107,N_5141);
or U5227 (N_5227,N_5165,N_5178);
nand U5228 (N_5228,N_5152,N_5180);
nor U5229 (N_5229,N_5196,N_5171);
and U5230 (N_5230,N_5156,N_5124);
and U5231 (N_5231,N_5185,N_5118);
nor U5232 (N_5232,N_5125,N_5198);
nand U5233 (N_5233,N_5176,N_5154);
nand U5234 (N_5234,N_5120,N_5161);
and U5235 (N_5235,N_5150,N_5127);
nand U5236 (N_5236,N_5105,N_5102);
nor U5237 (N_5237,N_5179,N_5144);
or U5238 (N_5238,N_5172,N_5169);
and U5239 (N_5239,N_5106,N_5123);
or U5240 (N_5240,N_5158,N_5191);
nor U5241 (N_5241,N_5119,N_5167);
nand U5242 (N_5242,N_5148,N_5187);
nor U5243 (N_5243,N_5135,N_5192);
and U5244 (N_5244,N_5194,N_5157);
and U5245 (N_5245,N_5128,N_5114);
nand U5246 (N_5246,N_5103,N_5113);
nor U5247 (N_5247,N_5139,N_5159);
nand U5248 (N_5248,N_5146,N_5101);
or U5249 (N_5249,N_5117,N_5177);
nor U5250 (N_5250,N_5138,N_5118);
and U5251 (N_5251,N_5181,N_5139);
or U5252 (N_5252,N_5104,N_5162);
or U5253 (N_5253,N_5188,N_5112);
nand U5254 (N_5254,N_5193,N_5136);
or U5255 (N_5255,N_5171,N_5111);
nor U5256 (N_5256,N_5188,N_5149);
and U5257 (N_5257,N_5140,N_5114);
nor U5258 (N_5258,N_5136,N_5125);
nand U5259 (N_5259,N_5159,N_5138);
or U5260 (N_5260,N_5139,N_5125);
or U5261 (N_5261,N_5109,N_5169);
or U5262 (N_5262,N_5131,N_5162);
or U5263 (N_5263,N_5108,N_5127);
or U5264 (N_5264,N_5151,N_5114);
or U5265 (N_5265,N_5183,N_5139);
nor U5266 (N_5266,N_5193,N_5191);
nand U5267 (N_5267,N_5107,N_5193);
nor U5268 (N_5268,N_5108,N_5156);
or U5269 (N_5269,N_5160,N_5143);
and U5270 (N_5270,N_5127,N_5101);
nand U5271 (N_5271,N_5138,N_5115);
nor U5272 (N_5272,N_5154,N_5187);
nand U5273 (N_5273,N_5186,N_5176);
nand U5274 (N_5274,N_5157,N_5120);
nor U5275 (N_5275,N_5120,N_5166);
or U5276 (N_5276,N_5125,N_5176);
or U5277 (N_5277,N_5142,N_5163);
nand U5278 (N_5278,N_5143,N_5150);
or U5279 (N_5279,N_5136,N_5103);
nand U5280 (N_5280,N_5180,N_5155);
or U5281 (N_5281,N_5197,N_5110);
and U5282 (N_5282,N_5132,N_5120);
nand U5283 (N_5283,N_5130,N_5144);
and U5284 (N_5284,N_5120,N_5183);
nor U5285 (N_5285,N_5159,N_5147);
or U5286 (N_5286,N_5139,N_5161);
or U5287 (N_5287,N_5105,N_5197);
and U5288 (N_5288,N_5180,N_5163);
and U5289 (N_5289,N_5148,N_5118);
nand U5290 (N_5290,N_5152,N_5113);
nor U5291 (N_5291,N_5168,N_5118);
and U5292 (N_5292,N_5129,N_5111);
and U5293 (N_5293,N_5129,N_5182);
or U5294 (N_5294,N_5180,N_5143);
and U5295 (N_5295,N_5165,N_5176);
or U5296 (N_5296,N_5132,N_5199);
or U5297 (N_5297,N_5107,N_5197);
nand U5298 (N_5298,N_5143,N_5136);
nand U5299 (N_5299,N_5129,N_5192);
and U5300 (N_5300,N_5203,N_5210);
and U5301 (N_5301,N_5293,N_5264);
nand U5302 (N_5302,N_5220,N_5225);
nor U5303 (N_5303,N_5214,N_5211);
nand U5304 (N_5304,N_5237,N_5280);
and U5305 (N_5305,N_5229,N_5209);
nand U5306 (N_5306,N_5275,N_5265);
xnor U5307 (N_5307,N_5285,N_5202);
or U5308 (N_5308,N_5289,N_5241);
nand U5309 (N_5309,N_5267,N_5256);
nand U5310 (N_5310,N_5271,N_5299);
or U5311 (N_5311,N_5288,N_5244);
or U5312 (N_5312,N_5218,N_5292);
nor U5313 (N_5313,N_5223,N_5282);
and U5314 (N_5314,N_5249,N_5227);
and U5315 (N_5315,N_5246,N_5258);
and U5316 (N_5316,N_5272,N_5200);
nor U5317 (N_5317,N_5286,N_5296);
nand U5318 (N_5318,N_5262,N_5221);
nor U5319 (N_5319,N_5260,N_5277);
and U5320 (N_5320,N_5233,N_5253);
or U5321 (N_5321,N_5206,N_5224);
nand U5322 (N_5322,N_5216,N_5269);
nand U5323 (N_5323,N_5204,N_5243);
nor U5324 (N_5324,N_5242,N_5232);
nor U5325 (N_5325,N_5266,N_5294);
or U5326 (N_5326,N_5248,N_5230);
or U5327 (N_5327,N_5250,N_5291);
nand U5328 (N_5328,N_5222,N_5297);
nand U5329 (N_5329,N_5207,N_5234);
nor U5330 (N_5330,N_5284,N_5231);
nand U5331 (N_5331,N_5236,N_5226);
and U5332 (N_5332,N_5217,N_5261);
nand U5333 (N_5333,N_5213,N_5273);
nand U5334 (N_5334,N_5283,N_5205);
and U5335 (N_5335,N_5254,N_5295);
nor U5336 (N_5336,N_5263,N_5235);
nor U5337 (N_5337,N_5257,N_5268);
nand U5338 (N_5338,N_5208,N_5287);
and U5339 (N_5339,N_5298,N_5219);
and U5340 (N_5340,N_5290,N_5276);
nor U5341 (N_5341,N_5247,N_5278);
nor U5342 (N_5342,N_5228,N_5255);
nand U5343 (N_5343,N_5212,N_5238);
nor U5344 (N_5344,N_5281,N_5201);
and U5345 (N_5345,N_5279,N_5245);
and U5346 (N_5346,N_5274,N_5215);
or U5347 (N_5347,N_5251,N_5259);
and U5348 (N_5348,N_5239,N_5240);
nand U5349 (N_5349,N_5270,N_5252);
nor U5350 (N_5350,N_5208,N_5291);
nor U5351 (N_5351,N_5249,N_5224);
nor U5352 (N_5352,N_5208,N_5216);
and U5353 (N_5353,N_5218,N_5250);
nand U5354 (N_5354,N_5267,N_5290);
nor U5355 (N_5355,N_5248,N_5269);
or U5356 (N_5356,N_5270,N_5293);
and U5357 (N_5357,N_5226,N_5203);
and U5358 (N_5358,N_5209,N_5265);
or U5359 (N_5359,N_5220,N_5223);
and U5360 (N_5360,N_5200,N_5225);
nand U5361 (N_5361,N_5248,N_5229);
nor U5362 (N_5362,N_5208,N_5293);
nor U5363 (N_5363,N_5239,N_5224);
or U5364 (N_5364,N_5201,N_5283);
nor U5365 (N_5365,N_5261,N_5202);
nand U5366 (N_5366,N_5260,N_5249);
or U5367 (N_5367,N_5219,N_5266);
nor U5368 (N_5368,N_5254,N_5237);
nor U5369 (N_5369,N_5294,N_5249);
nor U5370 (N_5370,N_5265,N_5241);
nor U5371 (N_5371,N_5231,N_5216);
and U5372 (N_5372,N_5260,N_5263);
and U5373 (N_5373,N_5215,N_5224);
and U5374 (N_5374,N_5257,N_5276);
nor U5375 (N_5375,N_5238,N_5223);
nand U5376 (N_5376,N_5271,N_5243);
nand U5377 (N_5377,N_5207,N_5227);
nor U5378 (N_5378,N_5210,N_5207);
xor U5379 (N_5379,N_5213,N_5235);
xor U5380 (N_5380,N_5238,N_5283);
nand U5381 (N_5381,N_5226,N_5211);
and U5382 (N_5382,N_5227,N_5261);
or U5383 (N_5383,N_5275,N_5247);
nand U5384 (N_5384,N_5255,N_5251);
or U5385 (N_5385,N_5224,N_5252);
nand U5386 (N_5386,N_5267,N_5275);
and U5387 (N_5387,N_5214,N_5243);
nor U5388 (N_5388,N_5278,N_5254);
or U5389 (N_5389,N_5244,N_5270);
or U5390 (N_5390,N_5265,N_5247);
nand U5391 (N_5391,N_5215,N_5262);
nand U5392 (N_5392,N_5274,N_5291);
and U5393 (N_5393,N_5265,N_5266);
or U5394 (N_5394,N_5278,N_5230);
and U5395 (N_5395,N_5279,N_5284);
nand U5396 (N_5396,N_5233,N_5282);
nand U5397 (N_5397,N_5280,N_5221);
nand U5398 (N_5398,N_5218,N_5230);
nor U5399 (N_5399,N_5209,N_5261);
nor U5400 (N_5400,N_5327,N_5305);
or U5401 (N_5401,N_5317,N_5386);
nor U5402 (N_5402,N_5364,N_5374);
or U5403 (N_5403,N_5306,N_5344);
or U5404 (N_5404,N_5313,N_5300);
and U5405 (N_5405,N_5359,N_5394);
or U5406 (N_5406,N_5360,N_5341);
nor U5407 (N_5407,N_5362,N_5399);
nand U5408 (N_5408,N_5388,N_5348);
or U5409 (N_5409,N_5321,N_5363);
or U5410 (N_5410,N_5358,N_5366);
nand U5411 (N_5411,N_5379,N_5377);
and U5412 (N_5412,N_5320,N_5372);
nor U5413 (N_5413,N_5310,N_5376);
or U5414 (N_5414,N_5307,N_5346);
nor U5415 (N_5415,N_5302,N_5345);
or U5416 (N_5416,N_5334,N_5304);
and U5417 (N_5417,N_5356,N_5390);
nor U5418 (N_5418,N_5350,N_5322);
or U5419 (N_5419,N_5333,N_5336);
nor U5420 (N_5420,N_5319,N_5315);
or U5421 (N_5421,N_5397,N_5371);
or U5422 (N_5422,N_5340,N_5368);
or U5423 (N_5423,N_5329,N_5342);
nand U5424 (N_5424,N_5331,N_5332);
and U5425 (N_5425,N_5398,N_5393);
and U5426 (N_5426,N_5349,N_5301);
nand U5427 (N_5427,N_5354,N_5369);
nand U5428 (N_5428,N_5343,N_5396);
or U5429 (N_5429,N_5365,N_5353);
nor U5430 (N_5430,N_5378,N_5395);
or U5431 (N_5431,N_5326,N_5357);
nand U5432 (N_5432,N_5323,N_5339);
or U5433 (N_5433,N_5309,N_5337);
nand U5434 (N_5434,N_5380,N_5361);
and U5435 (N_5435,N_5391,N_5325);
and U5436 (N_5436,N_5392,N_5385);
or U5437 (N_5437,N_5318,N_5389);
or U5438 (N_5438,N_5347,N_5308);
and U5439 (N_5439,N_5381,N_5352);
and U5440 (N_5440,N_5367,N_5355);
or U5441 (N_5441,N_5330,N_5324);
nand U5442 (N_5442,N_5338,N_5384);
nor U5443 (N_5443,N_5335,N_5316);
nand U5444 (N_5444,N_5314,N_5383);
or U5445 (N_5445,N_5370,N_5311);
nand U5446 (N_5446,N_5387,N_5328);
and U5447 (N_5447,N_5303,N_5382);
and U5448 (N_5448,N_5312,N_5375);
and U5449 (N_5449,N_5373,N_5351);
nor U5450 (N_5450,N_5317,N_5362);
and U5451 (N_5451,N_5308,N_5336);
and U5452 (N_5452,N_5349,N_5383);
or U5453 (N_5453,N_5326,N_5328);
and U5454 (N_5454,N_5324,N_5316);
nor U5455 (N_5455,N_5332,N_5329);
nand U5456 (N_5456,N_5376,N_5355);
or U5457 (N_5457,N_5338,N_5357);
nor U5458 (N_5458,N_5330,N_5372);
nor U5459 (N_5459,N_5337,N_5354);
nand U5460 (N_5460,N_5310,N_5322);
nor U5461 (N_5461,N_5394,N_5333);
nor U5462 (N_5462,N_5386,N_5348);
or U5463 (N_5463,N_5306,N_5307);
and U5464 (N_5464,N_5329,N_5395);
and U5465 (N_5465,N_5335,N_5367);
nand U5466 (N_5466,N_5354,N_5322);
and U5467 (N_5467,N_5329,N_5372);
nor U5468 (N_5468,N_5356,N_5368);
nor U5469 (N_5469,N_5365,N_5377);
or U5470 (N_5470,N_5316,N_5370);
xnor U5471 (N_5471,N_5361,N_5392);
nor U5472 (N_5472,N_5306,N_5348);
or U5473 (N_5473,N_5333,N_5356);
and U5474 (N_5474,N_5328,N_5359);
xnor U5475 (N_5475,N_5355,N_5396);
or U5476 (N_5476,N_5345,N_5383);
nand U5477 (N_5477,N_5347,N_5310);
and U5478 (N_5478,N_5399,N_5306);
nor U5479 (N_5479,N_5363,N_5344);
and U5480 (N_5480,N_5326,N_5307);
and U5481 (N_5481,N_5342,N_5379);
or U5482 (N_5482,N_5342,N_5358);
nand U5483 (N_5483,N_5353,N_5325);
nand U5484 (N_5484,N_5374,N_5304);
nand U5485 (N_5485,N_5312,N_5367);
and U5486 (N_5486,N_5328,N_5345);
or U5487 (N_5487,N_5370,N_5372);
nand U5488 (N_5488,N_5300,N_5392);
nor U5489 (N_5489,N_5361,N_5300);
nand U5490 (N_5490,N_5357,N_5355);
and U5491 (N_5491,N_5395,N_5341);
nand U5492 (N_5492,N_5393,N_5375);
nand U5493 (N_5493,N_5379,N_5365);
nand U5494 (N_5494,N_5366,N_5305);
nor U5495 (N_5495,N_5360,N_5375);
nand U5496 (N_5496,N_5323,N_5311);
nand U5497 (N_5497,N_5317,N_5361);
or U5498 (N_5498,N_5322,N_5363);
nand U5499 (N_5499,N_5304,N_5380);
or U5500 (N_5500,N_5414,N_5407);
and U5501 (N_5501,N_5454,N_5467);
and U5502 (N_5502,N_5469,N_5489);
and U5503 (N_5503,N_5411,N_5416);
nand U5504 (N_5504,N_5403,N_5449);
nor U5505 (N_5505,N_5412,N_5406);
nor U5506 (N_5506,N_5493,N_5466);
and U5507 (N_5507,N_5415,N_5464);
or U5508 (N_5508,N_5462,N_5495);
or U5509 (N_5509,N_5477,N_5409);
or U5510 (N_5510,N_5441,N_5463);
and U5511 (N_5511,N_5440,N_5482);
nand U5512 (N_5512,N_5405,N_5430);
or U5513 (N_5513,N_5436,N_5460);
and U5514 (N_5514,N_5451,N_5424);
and U5515 (N_5515,N_5434,N_5459);
xor U5516 (N_5516,N_5481,N_5444);
and U5517 (N_5517,N_5452,N_5450);
and U5518 (N_5518,N_5400,N_5458);
and U5519 (N_5519,N_5401,N_5479);
or U5520 (N_5520,N_5408,N_5465);
and U5521 (N_5521,N_5437,N_5473);
or U5522 (N_5522,N_5417,N_5443);
and U5523 (N_5523,N_5427,N_5420);
and U5524 (N_5524,N_5484,N_5442);
nand U5525 (N_5525,N_5488,N_5419);
nor U5526 (N_5526,N_5499,N_5446);
or U5527 (N_5527,N_5480,N_5438);
nand U5528 (N_5528,N_5455,N_5496);
and U5529 (N_5529,N_5428,N_5468);
nand U5530 (N_5530,N_5431,N_5483);
nand U5531 (N_5531,N_5435,N_5471);
or U5532 (N_5532,N_5413,N_5492);
and U5533 (N_5533,N_5497,N_5475);
and U5534 (N_5534,N_5486,N_5447);
or U5535 (N_5535,N_5418,N_5433);
and U5536 (N_5536,N_5426,N_5494);
or U5537 (N_5537,N_5478,N_5485);
and U5538 (N_5538,N_5498,N_5410);
xor U5539 (N_5539,N_5453,N_5421);
or U5540 (N_5540,N_5491,N_5425);
nor U5541 (N_5541,N_5487,N_5457);
or U5542 (N_5542,N_5432,N_5404);
nor U5543 (N_5543,N_5402,N_5439);
nand U5544 (N_5544,N_5429,N_5423);
nand U5545 (N_5545,N_5422,N_5456);
or U5546 (N_5546,N_5474,N_5461);
or U5547 (N_5547,N_5476,N_5445);
or U5548 (N_5548,N_5470,N_5490);
nand U5549 (N_5549,N_5448,N_5472);
nor U5550 (N_5550,N_5422,N_5401);
nand U5551 (N_5551,N_5437,N_5429);
and U5552 (N_5552,N_5444,N_5477);
nand U5553 (N_5553,N_5434,N_5415);
nand U5554 (N_5554,N_5413,N_5474);
nor U5555 (N_5555,N_5434,N_5435);
or U5556 (N_5556,N_5447,N_5467);
or U5557 (N_5557,N_5442,N_5434);
xor U5558 (N_5558,N_5418,N_5406);
and U5559 (N_5559,N_5406,N_5448);
and U5560 (N_5560,N_5465,N_5416);
and U5561 (N_5561,N_5471,N_5460);
or U5562 (N_5562,N_5476,N_5426);
nor U5563 (N_5563,N_5453,N_5423);
and U5564 (N_5564,N_5452,N_5476);
nor U5565 (N_5565,N_5406,N_5414);
nor U5566 (N_5566,N_5449,N_5418);
and U5567 (N_5567,N_5495,N_5415);
or U5568 (N_5568,N_5464,N_5421);
nand U5569 (N_5569,N_5440,N_5409);
nor U5570 (N_5570,N_5486,N_5408);
and U5571 (N_5571,N_5412,N_5445);
nor U5572 (N_5572,N_5420,N_5475);
and U5573 (N_5573,N_5467,N_5435);
and U5574 (N_5574,N_5468,N_5465);
and U5575 (N_5575,N_5434,N_5484);
nand U5576 (N_5576,N_5472,N_5439);
or U5577 (N_5577,N_5426,N_5453);
or U5578 (N_5578,N_5489,N_5405);
or U5579 (N_5579,N_5421,N_5411);
nor U5580 (N_5580,N_5401,N_5499);
xor U5581 (N_5581,N_5428,N_5451);
nand U5582 (N_5582,N_5482,N_5445);
nor U5583 (N_5583,N_5456,N_5480);
and U5584 (N_5584,N_5456,N_5479);
nand U5585 (N_5585,N_5408,N_5409);
or U5586 (N_5586,N_5488,N_5484);
nor U5587 (N_5587,N_5402,N_5435);
or U5588 (N_5588,N_5497,N_5431);
nand U5589 (N_5589,N_5442,N_5449);
and U5590 (N_5590,N_5414,N_5467);
and U5591 (N_5591,N_5401,N_5402);
nand U5592 (N_5592,N_5414,N_5497);
or U5593 (N_5593,N_5464,N_5497);
nand U5594 (N_5594,N_5460,N_5489);
or U5595 (N_5595,N_5489,N_5491);
nand U5596 (N_5596,N_5437,N_5406);
or U5597 (N_5597,N_5466,N_5471);
nand U5598 (N_5598,N_5469,N_5488);
nand U5599 (N_5599,N_5490,N_5473);
nor U5600 (N_5600,N_5568,N_5515);
or U5601 (N_5601,N_5540,N_5584);
and U5602 (N_5602,N_5545,N_5516);
nor U5603 (N_5603,N_5585,N_5575);
nand U5604 (N_5604,N_5533,N_5505);
nor U5605 (N_5605,N_5581,N_5569);
nand U5606 (N_5606,N_5573,N_5594);
or U5607 (N_5607,N_5541,N_5513);
nand U5608 (N_5608,N_5521,N_5552);
and U5609 (N_5609,N_5599,N_5514);
nor U5610 (N_5610,N_5534,N_5562);
and U5611 (N_5611,N_5537,N_5577);
nand U5612 (N_5612,N_5549,N_5565);
nor U5613 (N_5613,N_5557,N_5598);
nor U5614 (N_5614,N_5548,N_5566);
and U5615 (N_5615,N_5501,N_5524);
or U5616 (N_5616,N_5578,N_5597);
nand U5617 (N_5617,N_5588,N_5555);
or U5618 (N_5618,N_5520,N_5589);
nand U5619 (N_5619,N_5509,N_5593);
and U5620 (N_5620,N_5587,N_5596);
and U5621 (N_5621,N_5556,N_5504);
or U5622 (N_5622,N_5517,N_5511);
and U5623 (N_5623,N_5530,N_5576);
and U5624 (N_5624,N_5583,N_5563);
or U5625 (N_5625,N_5547,N_5527);
or U5626 (N_5626,N_5544,N_5553);
nor U5627 (N_5627,N_5539,N_5532);
nand U5628 (N_5628,N_5567,N_5510);
or U5629 (N_5629,N_5500,N_5523);
or U5630 (N_5630,N_5572,N_5580);
nand U5631 (N_5631,N_5582,N_5543);
nand U5632 (N_5632,N_5551,N_5519);
or U5633 (N_5633,N_5591,N_5528);
nor U5634 (N_5634,N_5564,N_5571);
or U5635 (N_5635,N_5502,N_5518);
or U5636 (N_5636,N_5579,N_5559);
nand U5637 (N_5637,N_5550,N_5561);
or U5638 (N_5638,N_5560,N_5506);
and U5639 (N_5639,N_5529,N_5512);
nor U5640 (N_5640,N_5592,N_5574);
nor U5641 (N_5641,N_5558,N_5503);
and U5642 (N_5642,N_5590,N_5536);
nor U5643 (N_5643,N_5542,N_5595);
and U5644 (N_5644,N_5535,N_5526);
and U5645 (N_5645,N_5525,N_5508);
or U5646 (N_5646,N_5538,N_5586);
nand U5647 (N_5647,N_5570,N_5522);
or U5648 (N_5648,N_5531,N_5507);
nand U5649 (N_5649,N_5546,N_5554);
nor U5650 (N_5650,N_5575,N_5573);
and U5651 (N_5651,N_5503,N_5570);
nor U5652 (N_5652,N_5575,N_5507);
nand U5653 (N_5653,N_5502,N_5550);
nor U5654 (N_5654,N_5584,N_5556);
nand U5655 (N_5655,N_5555,N_5583);
nor U5656 (N_5656,N_5544,N_5521);
nor U5657 (N_5657,N_5514,N_5548);
or U5658 (N_5658,N_5515,N_5511);
nor U5659 (N_5659,N_5580,N_5557);
xnor U5660 (N_5660,N_5536,N_5519);
or U5661 (N_5661,N_5507,N_5544);
xnor U5662 (N_5662,N_5522,N_5554);
or U5663 (N_5663,N_5585,N_5545);
nand U5664 (N_5664,N_5563,N_5524);
nand U5665 (N_5665,N_5533,N_5546);
and U5666 (N_5666,N_5594,N_5507);
nand U5667 (N_5667,N_5575,N_5545);
and U5668 (N_5668,N_5543,N_5556);
nor U5669 (N_5669,N_5511,N_5532);
and U5670 (N_5670,N_5596,N_5583);
nand U5671 (N_5671,N_5564,N_5522);
or U5672 (N_5672,N_5599,N_5550);
and U5673 (N_5673,N_5599,N_5501);
nor U5674 (N_5674,N_5521,N_5564);
nand U5675 (N_5675,N_5508,N_5554);
nand U5676 (N_5676,N_5557,N_5593);
or U5677 (N_5677,N_5589,N_5525);
or U5678 (N_5678,N_5519,N_5529);
nand U5679 (N_5679,N_5592,N_5590);
nor U5680 (N_5680,N_5519,N_5580);
nand U5681 (N_5681,N_5519,N_5533);
nand U5682 (N_5682,N_5568,N_5550);
or U5683 (N_5683,N_5543,N_5540);
or U5684 (N_5684,N_5544,N_5543);
nor U5685 (N_5685,N_5512,N_5552);
or U5686 (N_5686,N_5587,N_5508);
and U5687 (N_5687,N_5512,N_5541);
or U5688 (N_5688,N_5584,N_5538);
nand U5689 (N_5689,N_5548,N_5500);
and U5690 (N_5690,N_5597,N_5514);
and U5691 (N_5691,N_5511,N_5582);
xor U5692 (N_5692,N_5544,N_5569);
or U5693 (N_5693,N_5581,N_5513);
nor U5694 (N_5694,N_5599,N_5502);
or U5695 (N_5695,N_5599,N_5574);
nor U5696 (N_5696,N_5522,N_5581);
nor U5697 (N_5697,N_5585,N_5547);
and U5698 (N_5698,N_5522,N_5556);
nor U5699 (N_5699,N_5569,N_5596);
nand U5700 (N_5700,N_5675,N_5695);
nor U5701 (N_5701,N_5678,N_5669);
or U5702 (N_5702,N_5673,N_5618);
nand U5703 (N_5703,N_5622,N_5603);
nand U5704 (N_5704,N_5689,N_5682);
nand U5705 (N_5705,N_5607,N_5666);
and U5706 (N_5706,N_5627,N_5686);
nor U5707 (N_5707,N_5625,N_5645);
and U5708 (N_5708,N_5640,N_5667);
and U5709 (N_5709,N_5609,N_5613);
nor U5710 (N_5710,N_5680,N_5661);
nor U5711 (N_5711,N_5693,N_5639);
or U5712 (N_5712,N_5605,N_5624);
nor U5713 (N_5713,N_5628,N_5674);
xnor U5714 (N_5714,N_5629,N_5617);
or U5715 (N_5715,N_5650,N_5692);
or U5716 (N_5716,N_5641,N_5698);
or U5717 (N_5717,N_5600,N_5604);
nand U5718 (N_5718,N_5638,N_5615);
and U5719 (N_5719,N_5649,N_5691);
nand U5720 (N_5720,N_5697,N_5687);
nor U5721 (N_5721,N_5608,N_5671);
or U5722 (N_5722,N_5620,N_5637);
and U5723 (N_5723,N_5663,N_5616);
xnor U5724 (N_5724,N_5677,N_5614);
nor U5725 (N_5725,N_5633,N_5657);
nor U5726 (N_5726,N_5665,N_5631);
nand U5727 (N_5727,N_5648,N_5668);
nand U5728 (N_5728,N_5643,N_5626);
nor U5729 (N_5729,N_5684,N_5654);
nand U5730 (N_5730,N_5644,N_5690);
nand U5731 (N_5731,N_5659,N_5623);
or U5732 (N_5732,N_5602,N_5681);
and U5733 (N_5733,N_5610,N_5647);
and U5734 (N_5734,N_5655,N_5619);
nor U5735 (N_5735,N_5672,N_5676);
xor U5736 (N_5736,N_5652,N_5636);
and U5737 (N_5737,N_5653,N_5646);
nand U5738 (N_5738,N_5679,N_5685);
or U5739 (N_5739,N_5612,N_5664);
nand U5740 (N_5740,N_5660,N_5601);
and U5741 (N_5741,N_5632,N_5630);
nor U5742 (N_5742,N_5662,N_5606);
and U5743 (N_5743,N_5658,N_5635);
and U5744 (N_5744,N_5651,N_5621);
and U5745 (N_5745,N_5683,N_5611);
and U5746 (N_5746,N_5696,N_5642);
nand U5747 (N_5747,N_5670,N_5699);
and U5748 (N_5748,N_5656,N_5688);
and U5749 (N_5749,N_5634,N_5694);
or U5750 (N_5750,N_5612,N_5651);
or U5751 (N_5751,N_5663,N_5660);
and U5752 (N_5752,N_5671,N_5601);
nand U5753 (N_5753,N_5671,N_5678);
nor U5754 (N_5754,N_5671,N_5630);
nand U5755 (N_5755,N_5666,N_5665);
or U5756 (N_5756,N_5628,N_5690);
and U5757 (N_5757,N_5615,N_5604);
and U5758 (N_5758,N_5602,N_5645);
nor U5759 (N_5759,N_5682,N_5639);
nand U5760 (N_5760,N_5653,N_5685);
nand U5761 (N_5761,N_5660,N_5644);
nor U5762 (N_5762,N_5610,N_5652);
and U5763 (N_5763,N_5671,N_5621);
and U5764 (N_5764,N_5629,N_5680);
or U5765 (N_5765,N_5657,N_5660);
nand U5766 (N_5766,N_5662,N_5685);
nor U5767 (N_5767,N_5695,N_5638);
nor U5768 (N_5768,N_5664,N_5616);
nand U5769 (N_5769,N_5623,N_5656);
nand U5770 (N_5770,N_5625,N_5642);
and U5771 (N_5771,N_5626,N_5693);
nor U5772 (N_5772,N_5652,N_5678);
nand U5773 (N_5773,N_5625,N_5675);
or U5774 (N_5774,N_5689,N_5643);
nor U5775 (N_5775,N_5666,N_5619);
nor U5776 (N_5776,N_5612,N_5678);
nor U5777 (N_5777,N_5633,N_5683);
and U5778 (N_5778,N_5605,N_5687);
nand U5779 (N_5779,N_5685,N_5675);
or U5780 (N_5780,N_5692,N_5640);
nand U5781 (N_5781,N_5651,N_5630);
nor U5782 (N_5782,N_5666,N_5638);
nand U5783 (N_5783,N_5661,N_5642);
nand U5784 (N_5784,N_5605,N_5656);
nand U5785 (N_5785,N_5610,N_5675);
nand U5786 (N_5786,N_5668,N_5678);
nand U5787 (N_5787,N_5688,N_5694);
or U5788 (N_5788,N_5629,N_5677);
or U5789 (N_5789,N_5681,N_5642);
nand U5790 (N_5790,N_5698,N_5633);
and U5791 (N_5791,N_5606,N_5681);
or U5792 (N_5792,N_5684,N_5641);
and U5793 (N_5793,N_5657,N_5644);
and U5794 (N_5794,N_5621,N_5665);
or U5795 (N_5795,N_5627,N_5650);
or U5796 (N_5796,N_5626,N_5653);
and U5797 (N_5797,N_5600,N_5602);
and U5798 (N_5798,N_5603,N_5655);
or U5799 (N_5799,N_5635,N_5657);
and U5800 (N_5800,N_5793,N_5743);
or U5801 (N_5801,N_5734,N_5783);
nand U5802 (N_5802,N_5731,N_5710);
nor U5803 (N_5803,N_5779,N_5745);
or U5804 (N_5804,N_5754,N_5713);
nor U5805 (N_5805,N_5705,N_5776);
or U5806 (N_5806,N_5719,N_5789);
and U5807 (N_5807,N_5746,N_5727);
or U5808 (N_5808,N_5768,N_5750);
nand U5809 (N_5809,N_5715,N_5781);
or U5810 (N_5810,N_5758,N_5704);
or U5811 (N_5811,N_5794,N_5712);
or U5812 (N_5812,N_5786,N_5770);
nand U5813 (N_5813,N_5764,N_5780);
nor U5814 (N_5814,N_5733,N_5724);
and U5815 (N_5815,N_5778,N_5707);
or U5816 (N_5816,N_5765,N_5767);
and U5817 (N_5817,N_5756,N_5744);
and U5818 (N_5818,N_5708,N_5752);
and U5819 (N_5819,N_5714,N_5742);
nand U5820 (N_5820,N_5725,N_5762);
and U5821 (N_5821,N_5700,N_5728);
nor U5822 (N_5822,N_5763,N_5777);
nor U5823 (N_5823,N_5735,N_5753);
nand U5824 (N_5824,N_5773,N_5792);
nor U5825 (N_5825,N_5751,N_5720);
nor U5826 (N_5826,N_5772,N_5711);
and U5827 (N_5827,N_5723,N_5749);
nand U5828 (N_5828,N_5701,N_5760);
nor U5829 (N_5829,N_5782,N_5702);
nor U5830 (N_5830,N_5788,N_5717);
or U5831 (N_5831,N_5739,N_5785);
or U5832 (N_5832,N_5732,N_5797);
nor U5833 (N_5833,N_5774,N_5755);
nor U5834 (N_5834,N_5759,N_5798);
and U5835 (N_5835,N_5790,N_5761);
and U5836 (N_5836,N_5738,N_5799);
nand U5837 (N_5837,N_5737,N_5716);
nor U5838 (N_5838,N_5722,N_5740);
or U5839 (N_5839,N_5729,N_5757);
nand U5840 (N_5840,N_5766,N_5726);
or U5841 (N_5841,N_5709,N_5721);
nor U5842 (N_5842,N_5748,N_5784);
nand U5843 (N_5843,N_5771,N_5706);
nor U5844 (N_5844,N_5741,N_5769);
or U5845 (N_5845,N_5795,N_5736);
nor U5846 (N_5846,N_5718,N_5796);
nand U5847 (N_5847,N_5791,N_5787);
and U5848 (N_5848,N_5730,N_5775);
nand U5849 (N_5849,N_5703,N_5747);
nand U5850 (N_5850,N_5740,N_5762);
nor U5851 (N_5851,N_5773,N_5729);
or U5852 (N_5852,N_5711,N_5773);
and U5853 (N_5853,N_5727,N_5735);
and U5854 (N_5854,N_5750,N_5714);
nor U5855 (N_5855,N_5765,N_5798);
and U5856 (N_5856,N_5765,N_5749);
or U5857 (N_5857,N_5754,N_5719);
nor U5858 (N_5858,N_5735,N_5785);
nor U5859 (N_5859,N_5753,N_5773);
nand U5860 (N_5860,N_5736,N_5724);
nor U5861 (N_5861,N_5753,N_5762);
nand U5862 (N_5862,N_5771,N_5713);
nand U5863 (N_5863,N_5746,N_5709);
nor U5864 (N_5864,N_5764,N_5783);
or U5865 (N_5865,N_5781,N_5768);
and U5866 (N_5866,N_5748,N_5715);
nand U5867 (N_5867,N_5720,N_5708);
and U5868 (N_5868,N_5745,N_5771);
nor U5869 (N_5869,N_5785,N_5737);
xnor U5870 (N_5870,N_5770,N_5785);
xnor U5871 (N_5871,N_5770,N_5789);
or U5872 (N_5872,N_5777,N_5709);
and U5873 (N_5873,N_5785,N_5715);
xnor U5874 (N_5874,N_5713,N_5728);
and U5875 (N_5875,N_5744,N_5791);
and U5876 (N_5876,N_5753,N_5784);
nor U5877 (N_5877,N_5727,N_5716);
or U5878 (N_5878,N_5792,N_5749);
or U5879 (N_5879,N_5734,N_5793);
or U5880 (N_5880,N_5745,N_5706);
and U5881 (N_5881,N_5754,N_5736);
or U5882 (N_5882,N_5709,N_5756);
nor U5883 (N_5883,N_5798,N_5763);
nor U5884 (N_5884,N_5722,N_5761);
nand U5885 (N_5885,N_5765,N_5776);
or U5886 (N_5886,N_5751,N_5773);
or U5887 (N_5887,N_5796,N_5783);
nand U5888 (N_5888,N_5780,N_5723);
or U5889 (N_5889,N_5766,N_5714);
nand U5890 (N_5890,N_5701,N_5771);
nand U5891 (N_5891,N_5797,N_5705);
or U5892 (N_5892,N_5726,N_5777);
nand U5893 (N_5893,N_5713,N_5776);
and U5894 (N_5894,N_5799,N_5789);
nor U5895 (N_5895,N_5760,N_5738);
nor U5896 (N_5896,N_5717,N_5702);
nor U5897 (N_5897,N_5723,N_5782);
or U5898 (N_5898,N_5713,N_5785);
or U5899 (N_5899,N_5723,N_5768);
and U5900 (N_5900,N_5862,N_5819);
nor U5901 (N_5901,N_5857,N_5812);
and U5902 (N_5902,N_5849,N_5885);
nor U5903 (N_5903,N_5889,N_5838);
nand U5904 (N_5904,N_5817,N_5846);
or U5905 (N_5905,N_5873,N_5887);
xnor U5906 (N_5906,N_5897,N_5813);
and U5907 (N_5907,N_5800,N_5847);
nor U5908 (N_5908,N_5852,N_5875);
or U5909 (N_5909,N_5872,N_5884);
or U5910 (N_5910,N_5881,N_5871);
nand U5911 (N_5911,N_5818,N_5833);
and U5912 (N_5912,N_5854,N_5830);
or U5913 (N_5913,N_5880,N_5858);
nand U5914 (N_5914,N_5868,N_5877);
nand U5915 (N_5915,N_5883,N_5837);
nand U5916 (N_5916,N_5899,N_5896);
nor U5917 (N_5917,N_5848,N_5856);
nand U5918 (N_5918,N_5845,N_5882);
nand U5919 (N_5919,N_5886,N_5863);
or U5920 (N_5920,N_5893,N_5844);
and U5921 (N_5921,N_5892,N_5827);
and U5922 (N_5922,N_5866,N_5842);
nand U5923 (N_5923,N_5804,N_5824);
nand U5924 (N_5924,N_5864,N_5831);
nor U5925 (N_5925,N_5822,N_5851);
nand U5926 (N_5926,N_5869,N_5891);
nor U5927 (N_5927,N_5865,N_5834);
or U5928 (N_5928,N_5820,N_5876);
or U5929 (N_5929,N_5853,N_5879);
and U5930 (N_5930,N_5836,N_5810);
nor U5931 (N_5931,N_5826,N_5839);
nand U5932 (N_5932,N_5894,N_5803);
nand U5933 (N_5933,N_5835,N_5855);
nand U5934 (N_5934,N_5861,N_5860);
nand U5935 (N_5935,N_5841,N_5816);
nand U5936 (N_5936,N_5821,N_5825);
nor U5937 (N_5937,N_5843,N_5808);
nor U5938 (N_5938,N_5850,N_5809);
and U5939 (N_5939,N_5811,N_5805);
nand U5940 (N_5940,N_5898,N_5888);
xor U5941 (N_5941,N_5867,N_5815);
nand U5942 (N_5942,N_5832,N_5840);
nand U5943 (N_5943,N_5801,N_5814);
nor U5944 (N_5944,N_5859,N_5806);
xor U5945 (N_5945,N_5828,N_5874);
nor U5946 (N_5946,N_5895,N_5870);
nor U5947 (N_5947,N_5890,N_5829);
or U5948 (N_5948,N_5878,N_5807);
and U5949 (N_5949,N_5823,N_5802);
or U5950 (N_5950,N_5813,N_5800);
and U5951 (N_5951,N_5882,N_5879);
or U5952 (N_5952,N_5847,N_5825);
nor U5953 (N_5953,N_5813,N_5885);
nor U5954 (N_5954,N_5899,N_5834);
or U5955 (N_5955,N_5851,N_5888);
or U5956 (N_5956,N_5822,N_5833);
nand U5957 (N_5957,N_5875,N_5836);
and U5958 (N_5958,N_5884,N_5804);
nand U5959 (N_5959,N_5892,N_5818);
nor U5960 (N_5960,N_5875,N_5863);
nor U5961 (N_5961,N_5893,N_5882);
nor U5962 (N_5962,N_5870,N_5852);
nand U5963 (N_5963,N_5806,N_5827);
nand U5964 (N_5964,N_5803,N_5845);
nand U5965 (N_5965,N_5811,N_5897);
nand U5966 (N_5966,N_5886,N_5843);
nand U5967 (N_5967,N_5874,N_5806);
or U5968 (N_5968,N_5838,N_5893);
xor U5969 (N_5969,N_5851,N_5877);
and U5970 (N_5970,N_5879,N_5805);
nand U5971 (N_5971,N_5831,N_5812);
nand U5972 (N_5972,N_5804,N_5814);
and U5973 (N_5973,N_5870,N_5889);
nor U5974 (N_5974,N_5842,N_5863);
or U5975 (N_5975,N_5872,N_5894);
nand U5976 (N_5976,N_5852,N_5897);
nand U5977 (N_5977,N_5843,N_5892);
nand U5978 (N_5978,N_5857,N_5883);
nand U5979 (N_5979,N_5838,N_5801);
and U5980 (N_5980,N_5889,N_5862);
nand U5981 (N_5981,N_5851,N_5874);
nor U5982 (N_5982,N_5843,N_5874);
and U5983 (N_5983,N_5887,N_5806);
nand U5984 (N_5984,N_5820,N_5809);
or U5985 (N_5985,N_5851,N_5854);
and U5986 (N_5986,N_5818,N_5840);
and U5987 (N_5987,N_5807,N_5869);
nor U5988 (N_5988,N_5841,N_5824);
or U5989 (N_5989,N_5885,N_5882);
and U5990 (N_5990,N_5837,N_5861);
nor U5991 (N_5991,N_5850,N_5807);
nor U5992 (N_5992,N_5874,N_5890);
or U5993 (N_5993,N_5814,N_5840);
nand U5994 (N_5994,N_5821,N_5810);
nor U5995 (N_5995,N_5889,N_5886);
nor U5996 (N_5996,N_5840,N_5878);
and U5997 (N_5997,N_5808,N_5899);
and U5998 (N_5998,N_5856,N_5855);
and U5999 (N_5999,N_5845,N_5841);
nand U6000 (N_6000,N_5936,N_5925);
or U6001 (N_6001,N_5955,N_5972);
nor U6002 (N_6002,N_5983,N_5937);
or U6003 (N_6003,N_5918,N_5967);
nor U6004 (N_6004,N_5964,N_5924);
nand U6005 (N_6005,N_5959,N_5958);
nand U6006 (N_6006,N_5986,N_5970);
and U6007 (N_6007,N_5912,N_5901);
or U6008 (N_6008,N_5923,N_5952);
nand U6009 (N_6009,N_5926,N_5900);
and U6010 (N_6010,N_5914,N_5990);
nor U6011 (N_6011,N_5911,N_5902);
nand U6012 (N_6012,N_5919,N_5963);
nand U6013 (N_6013,N_5962,N_5980);
and U6014 (N_6014,N_5993,N_5987);
nor U6015 (N_6015,N_5968,N_5985);
nor U6016 (N_6016,N_5973,N_5945);
and U6017 (N_6017,N_5981,N_5954);
or U6018 (N_6018,N_5915,N_5978);
nor U6019 (N_6019,N_5944,N_5951);
nand U6020 (N_6020,N_5976,N_5984);
and U6021 (N_6021,N_5982,N_5991);
or U6022 (N_6022,N_5920,N_5975);
nand U6023 (N_6023,N_5907,N_5953);
nand U6024 (N_6024,N_5916,N_5960);
nand U6025 (N_6025,N_5996,N_5988);
and U6026 (N_6026,N_5943,N_5940);
nor U6027 (N_6027,N_5957,N_5909);
and U6028 (N_6028,N_5956,N_5950);
nor U6029 (N_6029,N_5929,N_5949);
and U6030 (N_6030,N_5998,N_5966);
or U6031 (N_6031,N_5999,N_5965);
and U6032 (N_6032,N_5946,N_5930);
or U6033 (N_6033,N_5942,N_5947);
and U6034 (N_6034,N_5994,N_5908);
and U6035 (N_6035,N_5969,N_5932);
nor U6036 (N_6036,N_5974,N_5910);
or U6037 (N_6037,N_5921,N_5905);
nand U6038 (N_6038,N_5904,N_5939);
and U6039 (N_6039,N_5979,N_5917);
and U6040 (N_6040,N_5971,N_5938);
or U6041 (N_6041,N_5903,N_5927);
nand U6042 (N_6042,N_5977,N_5933);
or U6043 (N_6043,N_5913,N_5906);
and U6044 (N_6044,N_5997,N_5961);
or U6045 (N_6045,N_5995,N_5948);
nor U6046 (N_6046,N_5989,N_5941);
and U6047 (N_6047,N_5922,N_5931);
or U6048 (N_6048,N_5992,N_5935);
and U6049 (N_6049,N_5928,N_5934);
and U6050 (N_6050,N_5923,N_5966);
nor U6051 (N_6051,N_5923,N_5930);
or U6052 (N_6052,N_5980,N_5948);
or U6053 (N_6053,N_5996,N_5925);
or U6054 (N_6054,N_5928,N_5905);
nand U6055 (N_6055,N_5967,N_5936);
nand U6056 (N_6056,N_5903,N_5965);
or U6057 (N_6057,N_5954,N_5948);
nand U6058 (N_6058,N_5973,N_5920);
and U6059 (N_6059,N_5999,N_5944);
xnor U6060 (N_6060,N_5966,N_5917);
nand U6061 (N_6061,N_5958,N_5912);
or U6062 (N_6062,N_5957,N_5972);
nor U6063 (N_6063,N_5962,N_5939);
nand U6064 (N_6064,N_5947,N_5962);
and U6065 (N_6065,N_5939,N_5907);
nor U6066 (N_6066,N_5963,N_5910);
and U6067 (N_6067,N_5966,N_5926);
nand U6068 (N_6068,N_5963,N_5944);
nand U6069 (N_6069,N_5919,N_5937);
nand U6070 (N_6070,N_5947,N_5948);
nand U6071 (N_6071,N_5978,N_5922);
nand U6072 (N_6072,N_5913,N_5951);
and U6073 (N_6073,N_5924,N_5920);
and U6074 (N_6074,N_5921,N_5990);
or U6075 (N_6075,N_5935,N_5989);
and U6076 (N_6076,N_5910,N_5914);
or U6077 (N_6077,N_5996,N_5923);
or U6078 (N_6078,N_5927,N_5910);
or U6079 (N_6079,N_5906,N_5932);
xnor U6080 (N_6080,N_5959,N_5916);
nor U6081 (N_6081,N_5929,N_5964);
nand U6082 (N_6082,N_5989,N_5942);
nand U6083 (N_6083,N_5996,N_5930);
nand U6084 (N_6084,N_5909,N_5938);
nand U6085 (N_6085,N_5932,N_5965);
nand U6086 (N_6086,N_5994,N_5950);
and U6087 (N_6087,N_5955,N_5993);
nand U6088 (N_6088,N_5935,N_5942);
and U6089 (N_6089,N_5950,N_5980);
or U6090 (N_6090,N_5911,N_5965);
nor U6091 (N_6091,N_5972,N_5945);
nand U6092 (N_6092,N_5943,N_5955);
nor U6093 (N_6093,N_5946,N_5900);
nand U6094 (N_6094,N_5999,N_5945);
nor U6095 (N_6095,N_5911,N_5993);
and U6096 (N_6096,N_5978,N_5960);
and U6097 (N_6097,N_5963,N_5988);
nor U6098 (N_6098,N_5909,N_5904);
nand U6099 (N_6099,N_5991,N_5912);
and U6100 (N_6100,N_6048,N_6028);
or U6101 (N_6101,N_6073,N_6095);
nor U6102 (N_6102,N_6035,N_6092);
nand U6103 (N_6103,N_6021,N_6096);
xnor U6104 (N_6104,N_6003,N_6041);
nand U6105 (N_6105,N_6065,N_6029);
or U6106 (N_6106,N_6060,N_6059);
nor U6107 (N_6107,N_6085,N_6025);
or U6108 (N_6108,N_6033,N_6009);
xnor U6109 (N_6109,N_6089,N_6049);
and U6110 (N_6110,N_6005,N_6000);
nand U6111 (N_6111,N_6084,N_6062);
or U6112 (N_6112,N_6001,N_6020);
nand U6113 (N_6113,N_6040,N_6070);
nor U6114 (N_6114,N_6076,N_6013);
or U6115 (N_6115,N_6077,N_6088);
and U6116 (N_6116,N_6052,N_6030);
or U6117 (N_6117,N_6051,N_6066);
nand U6118 (N_6118,N_6055,N_6008);
and U6119 (N_6119,N_6090,N_6044);
or U6120 (N_6120,N_6093,N_6026);
nor U6121 (N_6121,N_6063,N_6061);
and U6122 (N_6122,N_6004,N_6080);
or U6123 (N_6123,N_6094,N_6036);
nand U6124 (N_6124,N_6012,N_6016);
nand U6125 (N_6125,N_6069,N_6067);
nand U6126 (N_6126,N_6038,N_6010);
and U6127 (N_6127,N_6002,N_6082);
nor U6128 (N_6128,N_6017,N_6014);
nor U6129 (N_6129,N_6091,N_6064);
or U6130 (N_6130,N_6053,N_6006);
nand U6131 (N_6131,N_6074,N_6045);
nor U6132 (N_6132,N_6034,N_6022);
and U6133 (N_6133,N_6032,N_6018);
nand U6134 (N_6134,N_6075,N_6072);
nor U6135 (N_6135,N_6098,N_6087);
and U6136 (N_6136,N_6042,N_6056);
or U6137 (N_6137,N_6058,N_6043);
nor U6138 (N_6138,N_6079,N_6054);
nand U6139 (N_6139,N_6047,N_6011);
nor U6140 (N_6140,N_6057,N_6099);
or U6141 (N_6141,N_6086,N_6037);
and U6142 (N_6142,N_6071,N_6046);
and U6143 (N_6143,N_6083,N_6023);
nand U6144 (N_6144,N_6015,N_6068);
nand U6145 (N_6145,N_6019,N_6050);
and U6146 (N_6146,N_6097,N_6078);
nand U6147 (N_6147,N_6081,N_6031);
nor U6148 (N_6148,N_6027,N_6039);
or U6149 (N_6149,N_6007,N_6024);
nor U6150 (N_6150,N_6071,N_6048);
and U6151 (N_6151,N_6037,N_6031);
and U6152 (N_6152,N_6048,N_6064);
or U6153 (N_6153,N_6074,N_6091);
or U6154 (N_6154,N_6096,N_6079);
nor U6155 (N_6155,N_6002,N_6080);
xor U6156 (N_6156,N_6097,N_6030);
nor U6157 (N_6157,N_6049,N_6011);
nor U6158 (N_6158,N_6008,N_6086);
or U6159 (N_6159,N_6091,N_6006);
nand U6160 (N_6160,N_6095,N_6063);
and U6161 (N_6161,N_6098,N_6020);
nor U6162 (N_6162,N_6092,N_6025);
nor U6163 (N_6163,N_6026,N_6056);
nor U6164 (N_6164,N_6068,N_6048);
or U6165 (N_6165,N_6008,N_6025);
nand U6166 (N_6166,N_6033,N_6090);
nand U6167 (N_6167,N_6092,N_6023);
or U6168 (N_6168,N_6084,N_6037);
nand U6169 (N_6169,N_6068,N_6003);
xor U6170 (N_6170,N_6025,N_6022);
or U6171 (N_6171,N_6037,N_6016);
nor U6172 (N_6172,N_6056,N_6002);
or U6173 (N_6173,N_6049,N_6096);
nand U6174 (N_6174,N_6080,N_6006);
or U6175 (N_6175,N_6042,N_6004);
or U6176 (N_6176,N_6057,N_6073);
or U6177 (N_6177,N_6015,N_6061);
or U6178 (N_6178,N_6009,N_6062);
nand U6179 (N_6179,N_6038,N_6023);
nor U6180 (N_6180,N_6024,N_6076);
nor U6181 (N_6181,N_6003,N_6053);
and U6182 (N_6182,N_6044,N_6095);
nor U6183 (N_6183,N_6086,N_6080);
nand U6184 (N_6184,N_6014,N_6013);
or U6185 (N_6185,N_6040,N_6060);
nor U6186 (N_6186,N_6012,N_6024);
nor U6187 (N_6187,N_6060,N_6090);
and U6188 (N_6188,N_6034,N_6070);
nor U6189 (N_6189,N_6047,N_6063);
nand U6190 (N_6190,N_6050,N_6015);
or U6191 (N_6191,N_6010,N_6033);
or U6192 (N_6192,N_6095,N_6075);
and U6193 (N_6193,N_6031,N_6033);
nor U6194 (N_6194,N_6045,N_6084);
nand U6195 (N_6195,N_6008,N_6015);
or U6196 (N_6196,N_6098,N_6005);
nor U6197 (N_6197,N_6035,N_6075);
or U6198 (N_6198,N_6048,N_6092);
nor U6199 (N_6199,N_6084,N_6080);
nor U6200 (N_6200,N_6101,N_6170);
nor U6201 (N_6201,N_6108,N_6104);
or U6202 (N_6202,N_6158,N_6121);
nand U6203 (N_6203,N_6188,N_6164);
nor U6204 (N_6204,N_6177,N_6172);
nor U6205 (N_6205,N_6133,N_6176);
and U6206 (N_6206,N_6186,N_6192);
nand U6207 (N_6207,N_6138,N_6167);
or U6208 (N_6208,N_6152,N_6189);
and U6209 (N_6209,N_6130,N_6115);
nand U6210 (N_6210,N_6142,N_6131);
nand U6211 (N_6211,N_6109,N_6113);
nor U6212 (N_6212,N_6129,N_6155);
and U6213 (N_6213,N_6154,N_6124);
or U6214 (N_6214,N_6126,N_6150);
nor U6215 (N_6215,N_6106,N_6196);
or U6216 (N_6216,N_6144,N_6145);
and U6217 (N_6217,N_6122,N_6114);
or U6218 (N_6218,N_6123,N_6194);
or U6219 (N_6219,N_6163,N_6136);
or U6220 (N_6220,N_6139,N_6102);
nor U6221 (N_6221,N_6127,N_6169);
nand U6222 (N_6222,N_6107,N_6171);
and U6223 (N_6223,N_6153,N_6181);
nor U6224 (N_6224,N_6168,N_6162);
nand U6225 (N_6225,N_6190,N_6149);
or U6226 (N_6226,N_6103,N_6185);
and U6227 (N_6227,N_6166,N_6198);
or U6228 (N_6228,N_6141,N_6147);
nor U6229 (N_6229,N_6135,N_6184);
nor U6230 (N_6230,N_6128,N_6148);
and U6231 (N_6231,N_6193,N_6116);
nand U6232 (N_6232,N_6146,N_6183);
nor U6233 (N_6233,N_6100,N_6105);
or U6234 (N_6234,N_6125,N_6143);
nor U6235 (N_6235,N_6157,N_6197);
nand U6236 (N_6236,N_6161,N_6175);
or U6237 (N_6237,N_6165,N_6187);
and U6238 (N_6238,N_6119,N_6111);
xnor U6239 (N_6239,N_6182,N_6151);
or U6240 (N_6240,N_6110,N_6137);
xnor U6241 (N_6241,N_6160,N_6199);
or U6242 (N_6242,N_6191,N_6134);
or U6243 (N_6243,N_6180,N_6156);
and U6244 (N_6244,N_6132,N_6179);
or U6245 (N_6245,N_6173,N_6178);
or U6246 (N_6246,N_6118,N_6174);
and U6247 (N_6247,N_6112,N_6195);
and U6248 (N_6248,N_6140,N_6120);
or U6249 (N_6249,N_6159,N_6117);
nand U6250 (N_6250,N_6147,N_6109);
or U6251 (N_6251,N_6148,N_6157);
and U6252 (N_6252,N_6133,N_6149);
nand U6253 (N_6253,N_6129,N_6148);
nor U6254 (N_6254,N_6158,N_6178);
and U6255 (N_6255,N_6142,N_6105);
and U6256 (N_6256,N_6173,N_6180);
nor U6257 (N_6257,N_6184,N_6144);
nand U6258 (N_6258,N_6185,N_6161);
and U6259 (N_6259,N_6154,N_6127);
or U6260 (N_6260,N_6192,N_6185);
or U6261 (N_6261,N_6181,N_6168);
nor U6262 (N_6262,N_6191,N_6107);
nor U6263 (N_6263,N_6125,N_6151);
nor U6264 (N_6264,N_6116,N_6181);
nand U6265 (N_6265,N_6183,N_6191);
and U6266 (N_6266,N_6199,N_6166);
or U6267 (N_6267,N_6143,N_6194);
nor U6268 (N_6268,N_6102,N_6107);
and U6269 (N_6269,N_6116,N_6111);
or U6270 (N_6270,N_6111,N_6120);
nor U6271 (N_6271,N_6108,N_6105);
nand U6272 (N_6272,N_6129,N_6140);
or U6273 (N_6273,N_6173,N_6168);
and U6274 (N_6274,N_6145,N_6151);
or U6275 (N_6275,N_6189,N_6178);
nand U6276 (N_6276,N_6140,N_6112);
nand U6277 (N_6277,N_6169,N_6174);
and U6278 (N_6278,N_6138,N_6105);
nand U6279 (N_6279,N_6138,N_6196);
nor U6280 (N_6280,N_6144,N_6139);
nand U6281 (N_6281,N_6121,N_6189);
and U6282 (N_6282,N_6126,N_6168);
or U6283 (N_6283,N_6189,N_6150);
nor U6284 (N_6284,N_6173,N_6129);
xnor U6285 (N_6285,N_6166,N_6189);
nand U6286 (N_6286,N_6189,N_6162);
nor U6287 (N_6287,N_6122,N_6165);
nand U6288 (N_6288,N_6161,N_6103);
nor U6289 (N_6289,N_6148,N_6190);
nor U6290 (N_6290,N_6177,N_6121);
nand U6291 (N_6291,N_6106,N_6110);
nand U6292 (N_6292,N_6121,N_6188);
nand U6293 (N_6293,N_6148,N_6108);
nor U6294 (N_6294,N_6148,N_6184);
or U6295 (N_6295,N_6140,N_6111);
and U6296 (N_6296,N_6189,N_6185);
nor U6297 (N_6297,N_6138,N_6128);
xnor U6298 (N_6298,N_6127,N_6142);
nand U6299 (N_6299,N_6183,N_6192);
and U6300 (N_6300,N_6261,N_6268);
nand U6301 (N_6301,N_6280,N_6200);
nand U6302 (N_6302,N_6256,N_6253);
nand U6303 (N_6303,N_6238,N_6271);
and U6304 (N_6304,N_6288,N_6279);
nor U6305 (N_6305,N_6212,N_6298);
nand U6306 (N_6306,N_6277,N_6259);
nand U6307 (N_6307,N_6244,N_6224);
or U6308 (N_6308,N_6248,N_6230);
or U6309 (N_6309,N_6269,N_6245);
nor U6310 (N_6310,N_6206,N_6275);
nor U6311 (N_6311,N_6228,N_6235);
nand U6312 (N_6312,N_6281,N_6222);
or U6313 (N_6313,N_6272,N_6299);
nor U6314 (N_6314,N_6229,N_6239);
nand U6315 (N_6315,N_6243,N_6263);
nand U6316 (N_6316,N_6234,N_6241);
and U6317 (N_6317,N_6295,N_6209);
and U6318 (N_6318,N_6210,N_6262);
or U6319 (N_6319,N_6293,N_6273);
or U6320 (N_6320,N_6242,N_6231);
or U6321 (N_6321,N_6266,N_6225);
nand U6322 (N_6322,N_6289,N_6208);
and U6323 (N_6323,N_6216,N_6237);
or U6324 (N_6324,N_6260,N_6278);
or U6325 (N_6325,N_6246,N_6292);
nor U6326 (N_6326,N_6258,N_6251);
nand U6327 (N_6327,N_6217,N_6264);
or U6328 (N_6328,N_6285,N_6287);
and U6329 (N_6329,N_6205,N_6233);
xor U6330 (N_6330,N_6296,N_6203);
nand U6331 (N_6331,N_6211,N_6236);
nand U6332 (N_6332,N_6255,N_6218);
nand U6333 (N_6333,N_6214,N_6223);
nand U6334 (N_6334,N_6204,N_6254);
or U6335 (N_6335,N_6290,N_6219);
or U6336 (N_6336,N_6274,N_6252);
nand U6337 (N_6337,N_6226,N_6232);
and U6338 (N_6338,N_6284,N_6247);
nor U6339 (N_6339,N_6276,N_6283);
or U6340 (N_6340,N_6286,N_6240);
nand U6341 (N_6341,N_6270,N_6227);
nand U6342 (N_6342,N_6249,N_6221);
or U6343 (N_6343,N_6207,N_6267);
or U6344 (N_6344,N_6297,N_6215);
or U6345 (N_6345,N_6257,N_6291);
or U6346 (N_6346,N_6265,N_6294);
nor U6347 (N_6347,N_6213,N_6282);
nand U6348 (N_6348,N_6202,N_6250);
or U6349 (N_6349,N_6220,N_6201);
nor U6350 (N_6350,N_6207,N_6293);
nor U6351 (N_6351,N_6212,N_6250);
and U6352 (N_6352,N_6269,N_6288);
or U6353 (N_6353,N_6272,N_6211);
or U6354 (N_6354,N_6218,N_6240);
and U6355 (N_6355,N_6295,N_6224);
nor U6356 (N_6356,N_6284,N_6216);
or U6357 (N_6357,N_6272,N_6245);
nand U6358 (N_6358,N_6254,N_6248);
or U6359 (N_6359,N_6271,N_6248);
nand U6360 (N_6360,N_6296,N_6274);
nor U6361 (N_6361,N_6294,N_6295);
and U6362 (N_6362,N_6237,N_6209);
and U6363 (N_6363,N_6216,N_6264);
and U6364 (N_6364,N_6262,N_6217);
or U6365 (N_6365,N_6281,N_6267);
nor U6366 (N_6366,N_6241,N_6207);
nand U6367 (N_6367,N_6215,N_6200);
and U6368 (N_6368,N_6240,N_6219);
or U6369 (N_6369,N_6236,N_6269);
or U6370 (N_6370,N_6274,N_6268);
or U6371 (N_6371,N_6228,N_6203);
or U6372 (N_6372,N_6256,N_6270);
nor U6373 (N_6373,N_6238,N_6214);
nor U6374 (N_6374,N_6266,N_6222);
and U6375 (N_6375,N_6209,N_6229);
xnor U6376 (N_6376,N_6284,N_6291);
and U6377 (N_6377,N_6222,N_6295);
nor U6378 (N_6378,N_6262,N_6254);
and U6379 (N_6379,N_6230,N_6219);
nor U6380 (N_6380,N_6283,N_6247);
or U6381 (N_6381,N_6225,N_6226);
or U6382 (N_6382,N_6224,N_6290);
xor U6383 (N_6383,N_6223,N_6278);
nor U6384 (N_6384,N_6201,N_6208);
nand U6385 (N_6385,N_6277,N_6241);
nand U6386 (N_6386,N_6286,N_6243);
or U6387 (N_6387,N_6262,N_6293);
nor U6388 (N_6388,N_6202,N_6254);
nor U6389 (N_6389,N_6231,N_6204);
nor U6390 (N_6390,N_6286,N_6237);
nand U6391 (N_6391,N_6294,N_6232);
or U6392 (N_6392,N_6267,N_6223);
or U6393 (N_6393,N_6293,N_6256);
or U6394 (N_6394,N_6202,N_6200);
or U6395 (N_6395,N_6265,N_6235);
or U6396 (N_6396,N_6275,N_6295);
or U6397 (N_6397,N_6268,N_6220);
xnor U6398 (N_6398,N_6203,N_6255);
xor U6399 (N_6399,N_6267,N_6205);
and U6400 (N_6400,N_6382,N_6387);
or U6401 (N_6401,N_6325,N_6306);
and U6402 (N_6402,N_6304,N_6357);
nor U6403 (N_6403,N_6336,N_6318);
xor U6404 (N_6404,N_6345,N_6307);
and U6405 (N_6405,N_6353,N_6392);
or U6406 (N_6406,N_6363,N_6328);
nand U6407 (N_6407,N_6395,N_6380);
nor U6408 (N_6408,N_6398,N_6364);
or U6409 (N_6409,N_6319,N_6366);
and U6410 (N_6410,N_6374,N_6361);
and U6411 (N_6411,N_6394,N_6321);
nand U6412 (N_6412,N_6376,N_6393);
or U6413 (N_6413,N_6350,N_6302);
or U6414 (N_6414,N_6343,N_6338);
nor U6415 (N_6415,N_6397,N_6370);
or U6416 (N_6416,N_6388,N_6355);
nor U6417 (N_6417,N_6391,N_6308);
nor U6418 (N_6418,N_6326,N_6359);
nand U6419 (N_6419,N_6327,N_6332);
and U6420 (N_6420,N_6312,N_6351);
nand U6421 (N_6421,N_6316,N_6372);
or U6422 (N_6422,N_6375,N_6389);
nand U6423 (N_6423,N_6313,N_6309);
nand U6424 (N_6424,N_6323,N_6303);
nand U6425 (N_6425,N_6314,N_6378);
nand U6426 (N_6426,N_6354,N_6385);
and U6427 (N_6427,N_6386,N_6333);
and U6428 (N_6428,N_6301,N_6311);
nand U6429 (N_6429,N_6377,N_6330);
or U6430 (N_6430,N_6356,N_6310);
or U6431 (N_6431,N_6334,N_6305);
nand U6432 (N_6432,N_6371,N_6344);
or U6433 (N_6433,N_6365,N_6390);
xnor U6434 (N_6434,N_6337,N_6324);
nand U6435 (N_6435,N_6369,N_6331);
or U6436 (N_6436,N_6381,N_6346);
and U6437 (N_6437,N_6317,N_6335);
nand U6438 (N_6438,N_6348,N_6320);
nand U6439 (N_6439,N_6396,N_6373);
and U6440 (N_6440,N_6384,N_6358);
nor U6441 (N_6441,N_6399,N_6340);
or U6442 (N_6442,N_6347,N_6329);
nor U6443 (N_6443,N_6341,N_6379);
nor U6444 (N_6444,N_6368,N_6383);
and U6445 (N_6445,N_6339,N_6360);
or U6446 (N_6446,N_6367,N_6362);
nor U6447 (N_6447,N_6352,N_6322);
and U6448 (N_6448,N_6315,N_6342);
nand U6449 (N_6449,N_6349,N_6300);
and U6450 (N_6450,N_6314,N_6301);
nand U6451 (N_6451,N_6346,N_6314);
or U6452 (N_6452,N_6334,N_6390);
nand U6453 (N_6453,N_6324,N_6322);
nor U6454 (N_6454,N_6324,N_6361);
nand U6455 (N_6455,N_6319,N_6386);
or U6456 (N_6456,N_6346,N_6338);
nor U6457 (N_6457,N_6359,N_6354);
or U6458 (N_6458,N_6351,N_6372);
and U6459 (N_6459,N_6353,N_6386);
nor U6460 (N_6460,N_6333,N_6325);
or U6461 (N_6461,N_6395,N_6304);
or U6462 (N_6462,N_6380,N_6366);
or U6463 (N_6463,N_6369,N_6338);
nand U6464 (N_6464,N_6326,N_6369);
nor U6465 (N_6465,N_6335,N_6338);
or U6466 (N_6466,N_6378,N_6368);
xnor U6467 (N_6467,N_6329,N_6309);
nand U6468 (N_6468,N_6333,N_6319);
nand U6469 (N_6469,N_6345,N_6348);
and U6470 (N_6470,N_6351,N_6384);
and U6471 (N_6471,N_6325,N_6330);
nand U6472 (N_6472,N_6340,N_6342);
nand U6473 (N_6473,N_6341,N_6396);
or U6474 (N_6474,N_6343,N_6305);
or U6475 (N_6475,N_6310,N_6311);
or U6476 (N_6476,N_6325,N_6338);
nor U6477 (N_6477,N_6350,N_6347);
and U6478 (N_6478,N_6386,N_6335);
nand U6479 (N_6479,N_6301,N_6322);
nand U6480 (N_6480,N_6356,N_6322);
or U6481 (N_6481,N_6390,N_6353);
or U6482 (N_6482,N_6335,N_6336);
and U6483 (N_6483,N_6325,N_6337);
or U6484 (N_6484,N_6388,N_6392);
nor U6485 (N_6485,N_6311,N_6380);
nor U6486 (N_6486,N_6331,N_6314);
nand U6487 (N_6487,N_6312,N_6396);
or U6488 (N_6488,N_6343,N_6330);
nand U6489 (N_6489,N_6350,N_6314);
nand U6490 (N_6490,N_6384,N_6397);
or U6491 (N_6491,N_6378,N_6322);
or U6492 (N_6492,N_6350,N_6329);
or U6493 (N_6493,N_6374,N_6378);
nand U6494 (N_6494,N_6350,N_6322);
nor U6495 (N_6495,N_6360,N_6394);
and U6496 (N_6496,N_6351,N_6340);
or U6497 (N_6497,N_6366,N_6383);
and U6498 (N_6498,N_6390,N_6300);
and U6499 (N_6499,N_6349,N_6342);
and U6500 (N_6500,N_6423,N_6497);
or U6501 (N_6501,N_6417,N_6462);
nand U6502 (N_6502,N_6456,N_6430);
nor U6503 (N_6503,N_6411,N_6450);
nand U6504 (N_6504,N_6463,N_6453);
and U6505 (N_6505,N_6457,N_6405);
nor U6506 (N_6506,N_6482,N_6498);
nand U6507 (N_6507,N_6445,N_6495);
nand U6508 (N_6508,N_6477,N_6487);
or U6509 (N_6509,N_6490,N_6481);
and U6510 (N_6510,N_6427,N_6451);
or U6511 (N_6511,N_6439,N_6435);
and U6512 (N_6512,N_6479,N_6449);
nand U6513 (N_6513,N_6419,N_6438);
nor U6514 (N_6514,N_6493,N_6415);
or U6515 (N_6515,N_6454,N_6408);
or U6516 (N_6516,N_6468,N_6425);
nand U6517 (N_6517,N_6474,N_6418);
or U6518 (N_6518,N_6409,N_6424);
or U6519 (N_6519,N_6492,N_6486);
nand U6520 (N_6520,N_6480,N_6432);
or U6521 (N_6521,N_6437,N_6401);
nor U6522 (N_6522,N_6422,N_6494);
and U6523 (N_6523,N_6429,N_6471);
nor U6524 (N_6524,N_6473,N_6460);
nand U6525 (N_6525,N_6403,N_6484);
nand U6526 (N_6526,N_6499,N_6414);
and U6527 (N_6527,N_6413,N_6440);
and U6528 (N_6528,N_6443,N_6489);
nand U6529 (N_6529,N_6466,N_6470);
nor U6530 (N_6530,N_6433,N_6442);
or U6531 (N_6531,N_6452,N_6496);
nand U6532 (N_6532,N_6467,N_6441);
or U6533 (N_6533,N_6459,N_6476);
nor U6534 (N_6534,N_6434,N_6446);
xor U6535 (N_6535,N_6448,N_6436);
nand U6536 (N_6536,N_6421,N_6464);
or U6537 (N_6537,N_6491,N_6412);
and U6538 (N_6538,N_6485,N_6400);
nor U6539 (N_6539,N_6428,N_6406);
nor U6540 (N_6540,N_6410,N_6488);
or U6541 (N_6541,N_6404,N_6444);
and U6542 (N_6542,N_6472,N_6455);
or U6543 (N_6543,N_6431,N_6407);
or U6544 (N_6544,N_6426,N_6458);
nor U6545 (N_6545,N_6483,N_6465);
nand U6546 (N_6546,N_6402,N_6420);
and U6547 (N_6547,N_6478,N_6469);
nand U6548 (N_6548,N_6416,N_6461);
nor U6549 (N_6549,N_6447,N_6475);
or U6550 (N_6550,N_6474,N_6432);
and U6551 (N_6551,N_6455,N_6475);
nand U6552 (N_6552,N_6402,N_6436);
nor U6553 (N_6553,N_6474,N_6491);
nor U6554 (N_6554,N_6452,N_6476);
nor U6555 (N_6555,N_6452,N_6483);
and U6556 (N_6556,N_6411,N_6415);
nor U6557 (N_6557,N_6472,N_6400);
nand U6558 (N_6558,N_6446,N_6487);
or U6559 (N_6559,N_6470,N_6479);
or U6560 (N_6560,N_6491,N_6430);
nand U6561 (N_6561,N_6405,N_6450);
nand U6562 (N_6562,N_6474,N_6446);
nand U6563 (N_6563,N_6486,N_6476);
nand U6564 (N_6564,N_6420,N_6409);
nand U6565 (N_6565,N_6458,N_6407);
or U6566 (N_6566,N_6476,N_6496);
nor U6567 (N_6567,N_6459,N_6483);
or U6568 (N_6568,N_6493,N_6459);
nor U6569 (N_6569,N_6488,N_6492);
and U6570 (N_6570,N_6460,N_6426);
and U6571 (N_6571,N_6460,N_6462);
and U6572 (N_6572,N_6443,N_6401);
or U6573 (N_6573,N_6460,N_6449);
or U6574 (N_6574,N_6472,N_6435);
nor U6575 (N_6575,N_6455,N_6498);
or U6576 (N_6576,N_6492,N_6405);
or U6577 (N_6577,N_6444,N_6458);
and U6578 (N_6578,N_6437,N_6446);
nor U6579 (N_6579,N_6403,N_6407);
nor U6580 (N_6580,N_6474,N_6451);
nand U6581 (N_6581,N_6428,N_6485);
or U6582 (N_6582,N_6419,N_6463);
or U6583 (N_6583,N_6400,N_6448);
nor U6584 (N_6584,N_6459,N_6479);
and U6585 (N_6585,N_6468,N_6478);
and U6586 (N_6586,N_6468,N_6482);
or U6587 (N_6587,N_6432,N_6459);
nor U6588 (N_6588,N_6401,N_6404);
nand U6589 (N_6589,N_6427,N_6480);
xnor U6590 (N_6590,N_6478,N_6499);
or U6591 (N_6591,N_6488,N_6411);
and U6592 (N_6592,N_6457,N_6468);
nand U6593 (N_6593,N_6449,N_6482);
or U6594 (N_6594,N_6449,N_6408);
and U6595 (N_6595,N_6452,N_6412);
nor U6596 (N_6596,N_6426,N_6449);
or U6597 (N_6597,N_6431,N_6414);
and U6598 (N_6598,N_6461,N_6417);
nor U6599 (N_6599,N_6433,N_6477);
nand U6600 (N_6600,N_6573,N_6539);
xor U6601 (N_6601,N_6588,N_6546);
nand U6602 (N_6602,N_6520,N_6565);
and U6603 (N_6603,N_6512,N_6574);
and U6604 (N_6604,N_6524,N_6569);
and U6605 (N_6605,N_6580,N_6567);
nor U6606 (N_6606,N_6547,N_6576);
and U6607 (N_6607,N_6592,N_6502);
nand U6608 (N_6608,N_6522,N_6550);
nor U6609 (N_6609,N_6509,N_6599);
nor U6610 (N_6610,N_6513,N_6518);
or U6611 (N_6611,N_6538,N_6535);
or U6612 (N_6612,N_6545,N_6598);
or U6613 (N_6613,N_6560,N_6594);
and U6614 (N_6614,N_6585,N_6591);
nand U6615 (N_6615,N_6596,N_6577);
nor U6616 (N_6616,N_6561,N_6571);
nand U6617 (N_6617,N_6534,N_6552);
or U6618 (N_6618,N_6541,N_6515);
nor U6619 (N_6619,N_6553,N_6528);
nor U6620 (N_6620,N_6523,N_6559);
nor U6621 (N_6621,N_6554,N_6564);
nand U6622 (N_6622,N_6548,N_6506);
nor U6623 (N_6623,N_6556,N_6500);
or U6624 (N_6624,N_6507,N_6589);
or U6625 (N_6625,N_6551,N_6570);
or U6626 (N_6626,N_6508,N_6575);
and U6627 (N_6627,N_6579,N_6537);
or U6628 (N_6628,N_6530,N_6503);
nand U6629 (N_6629,N_6540,N_6555);
nor U6630 (N_6630,N_6514,N_6525);
nand U6631 (N_6631,N_6531,N_6529);
nand U6632 (N_6632,N_6501,N_6511);
nand U6633 (N_6633,N_6521,N_6584);
or U6634 (N_6634,N_6563,N_6505);
or U6635 (N_6635,N_6593,N_6543);
nor U6636 (N_6636,N_6583,N_6510);
and U6637 (N_6637,N_6566,N_6572);
nor U6638 (N_6638,N_6544,N_6542);
nand U6639 (N_6639,N_6519,N_6590);
nor U6640 (N_6640,N_6504,N_6558);
or U6641 (N_6641,N_6586,N_6595);
or U6642 (N_6642,N_6597,N_6532);
and U6643 (N_6643,N_6533,N_6568);
and U6644 (N_6644,N_6587,N_6516);
and U6645 (N_6645,N_6578,N_6517);
and U6646 (N_6646,N_6527,N_6557);
or U6647 (N_6647,N_6581,N_6526);
and U6648 (N_6648,N_6562,N_6582);
and U6649 (N_6649,N_6549,N_6536);
and U6650 (N_6650,N_6504,N_6516);
or U6651 (N_6651,N_6510,N_6512);
or U6652 (N_6652,N_6590,N_6514);
nor U6653 (N_6653,N_6590,N_6525);
or U6654 (N_6654,N_6529,N_6574);
nand U6655 (N_6655,N_6549,N_6566);
and U6656 (N_6656,N_6558,N_6586);
or U6657 (N_6657,N_6556,N_6548);
nand U6658 (N_6658,N_6599,N_6520);
or U6659 (N_6659,N_6543,N_6595);
or U6660 (N_6660,N_6535,N_6592);
nor U6661 (N_6661,N_6507,N_6581);
or U6662 (N_6662,N_6546,N_6585);
or U6663 (N_6663,N_6520,N_6547);
nor U6664 (N_6664,N_6542,N_6533);
nor U6665 (N_6665,N_6555,N_6566);
nor U6666 (N_6666,N_6500,N_6552);
or U6667 (N_6667,N_6563,N_6534);
nand U6668 (N_6668,N_6535,N_6567);
nor U6669 (N_6669,N_6560,N_6543);
nand U6670 (N_6670,N_6533,N_6555);
nand U6671 (N_6671,N_6561,N_6518);
and U6672 (N_6672,N_6570,N_6528);
nor U6673 (N_6673,N_6543,N_6592);
or U6674 (N_6674,N_6596,N_6502);
and U6675 (N_6675,N_6597,N_6535);
and U6676 (N_6676,N_6581,N_6579);
nor U6677 (N_6677,N_6540,N_6550);
and U6678 (N_6678,N_6570,N_6592);
nand U6679 (N_6679,N_6594,N_6518);
nor U6680 (N_6680,N_6540,N_6552);
and U6681 (N_6681,N_6594,N_6595);
or U6682 (N_6682,N_6528,N_6506);
or U6683 (N_6683,N_6508,N_6536);
or U6684 (N_6684,N_6546,N_6587);
or U6685 (N_6685,N_6525,N_6531);
and U6686 (N_6686,N_6549,N_6553);
nand U6687 (N_6687,N_6508,N_6589);
nand U6688 (N_6688,N_6535,N_6590);
and U6689 (N_6689,N_6528,N_6571);
nand U6690 (N_6690,N_6514,N_6564);
nand U6691 (N_6691,N_6523,N_6596);
and U6692 (N_6692,N_6567,N_6573);
nor U6693 (N_6693,N_6588,N_6590);
or U6694 (N_6694,N_6581,N_6552);
nor U6695 (N_6695,N_6599,N_6514);
nand U6696 (N_6696,N_6509,N_6569);
or U6697 (N_6697,N_6530,N_6521);
and U6698 (N_6698,N_6518,N_6562);
and U6699 (N_6699,N_6536,N_6548);
or U6700 (N_6700,N_6606,N_6622);
nor U6701 (N_6701,N_6632,N_6669);
or U6702 (N_6702,N_6620,N_6618);
and U6703 (N_6703,N_6611,N_6633);
or U6704 (N_6704,N_6684,N_6619);
nand U6705 (N_6705,N_6671,N_6615);
nand U6706 (N_6706,N_6681,N_6677);
or U6707 (N_6707,N_6610,N_6693);
and U6708 (N_6708,N_6697,N_6602);
nor U6709 (N_6709,N_6699,N_6656);
nand U6710 (N_6710,N_6692,N_6666);
and U6711 (N_6711,N_6609,N_6655);
nand U6712 (N_6712,N_6635,N_6649);
or U6713 (N_6713,N_6694,N_6690);
and U6714 (N_6714,N_6667,N_6680);
or U6715 (N_6715,N_6647,N_6689);
nor U6716 (N_6716,N_6621,N_6634);
or U6717 (N_6717,N_6696,N_6644);
or U6718 (N_6718,N_6657,N_6641);
and U6719 (N_6719,N_6637,N_6676);
nor U6720 (N_6720,N_6668,N_6600);
nand U6721 (N_6721,N_6646,N_6613);
nand U6722 (N_6722,N_6652,N_6695);
and U6723 (N_6723,N_6643,N_6679);
or U6724 (N_6724,N_6665,N_6654);
and U6725 (N_6725,N_6614,N_6626);
nor U6726 (N_6726,N_6678,N_6686);
or U6727 (N_6727,N_6603,N_6658);
nor U6728 (N_6728,N_6608,N_6687);
and U6729 (N_6729,N_6640,N_6659);
and U6730 (N_6730,N_6682,N_6648);
or U6731 (N_6731,N_6660,N_6661);
nand U6732 (N_6732,N_6625,N_6638);
nor U6733 (N_6733,N_6645,N_6673);
or U6734 (N_6734,N_6691,N_6601);
or U6735 (N_6735,N_6616,N_6624);
nor U6736 (N_6736,N_6612,N_6674);
nor U6737 (N_6737,N_6698,N_6683);
or U6738 (N_6738,N_6685,N_6636);
nor U6739 (N_6739,N_6623,N_6670);
nand U6740 (N_6740,N_6653,N_6607);
nor U6741 (N_6741,N_6605,N_6650);
nor U6742 (N_6742,N_6688,N_6663);
nand U6743 (N_6743,N_6672,N_6662);
nor U6744 (N_6744,N_6639,N_6604);
nor U6745 (N_6745,N_6627,N_6629);
and U6746 (N_6746,N_6617,N_6630);
nand U6747 (N_6747,N_6651,N_6631);
and U6748 (N_6748,N_6628,N_6664);
xor U6749 (N_6749,N_6675,N_6642);
nand U6750 (N_6750,N_6648,N_6693);
and U6751 (N_6751,N_6689,N_6602);
xor U6752 (N_6752,N_6634,N_6614);
nand U6753 (N_6753,N_6657,N_6647);
xnor U6754 (N_6754,N_6682,N_6664);
nand U6755 (N_6755,N_6654,N_6639);
or U6756 (N_6756,N_6624,N_6684);
nand U6757 (N_6757,N_6644,N_6634);
nand U6758 (N_6758,N_6617,N_6646);
nor U6759 (N_6759,N_6683,N_6618);
nor U6760 (N_6760,N_6692,N_6634);
or U6761 (N_6761,N_6695,N_6677);
and U6762 (N_6762,N_6665,N_6648);
nand U6763 (N_6763,N_6678,N_6628);
nor U6764 (N_6764,N_6629,N_6662);
and U6765 (N_6765,N_6657,N_6630);
nor U6766 (N_6766,N_6667,N_6603);
nand U6767 (N_6767,N_6647,N_6625);
nand U6768 (N_6768,N_6609,N_6660);
nand U6769 (N_6769,N_6677,N_6664);
nor U6770 (N_6770,N_6612,N_6648);
and U6771 (N_6771,N_6681,N_6645);
nand U6772 (N_6772,N_6656,N_6602);
or U6773 (N_6773,N_6681,N_6678);
and U6774 (N_6774,N_6618,N_6653);
and U6775 (N_6775,N_6654,N_6675);
and U6776 (N_6776,N_6625,N_6667);
and U6777 (N_6777,N_6643,N_6695);
and U6778 (N_6778,N_6635,N_6662);
nor U6779 (N_6779,N_6663,N_6613);
or U6780 (N_6780,N_6609,N_6677);
nand U6781 (N_6781,N_6647,N_6613);
or U6782 (N_6782,N_6663,N_6655);
and U6783 (N_6783,N_6686,N_6651);
or U6784 (N_6784,N_6611,N_6613);
and U6785 (N_6785,N_6617,N_6610);
nor U6786 (N_6786,N_6667,N_6614);
or U6787 (N_6787,N_6661,N_6675);
nand U6788 (N_6788,N_6695,N_6692);
nand U6789 (N_6789,N_6611,N_6691);
or U6790 (N_6790,N_6693,N_6644);
and U6791 (N_6791,N_6655,N_6622);
nor U6792 (N_6792,N_6613,N_6688);
nand U6793 (N_6793,N_6660,N_6664);
nor U6794 (N_6794,N_6639,N_6627);
nor U6795 (N_6795,N_6600,N_6651);
and U6796 (N_6796,N_6680,N_6638);
nor U6797 (N_6797,N_6620,N_6657);
nand U6798 (N_6798,N_6609,N_6614);
and U6799 (N_6799,N_6660,N_6688);
nand U6800 (N_6800,N_6706,N_6747);
and U6801 (N_6801,N_6739,N_6743);
nand U6802 (N_6802,N_6756,N_6730);
and U6803 (N_6803,N_6733,N_6765);
or U6804 (N_6804,N_6758,N_6787);
nor U6805 (N_6805,N_6795,N_6770);
nand U6806 (N_6806,N_6735,N_6729);
or U6807 (N_6807,N_6768,N_6785);
and U6808 (N_6808,N_6726,N_6736);
and U6809 (N_6809,N_6746,N_6789);
and U6810 (N_6810,N_6759,N_6777);
nand U6811 (N_6811,N_6760,N_6797);
nand U6812 (N_6812,N_6796,N_6761);
and U6813 (N_6813,N_6757,N_6709);
nor U6814 (N_6814,N_6798,N_6719);
and U6815 (N_6815,N_6715,N_6755);
or U6816 (N_6816,N_6741,N_6779);
nor U6817 (N_6817,N_6763,N_6792);
nand U6818 (N_6818,N_6794,N_6714);
and U6819 (N_6819,N_6717,N_6725);
and U6820 (N_6820,N_6751,N_6703);
nor U6821 (N_6821,N_6700,N_6716);
nor U6822 (N_6822,N_6780,N_6712);
nand U6823 (N_6823,N_6788,N_6718);
nand U6824 (N_6824,N_6721,N_6754);
nor U6825 (N_6825,N_6781,N_6786);
nand U6826 (N_6826,N_6737,N_6723);
or U6827 (N_6827,N_6720,N_6771);
or U6828 (N_6828,N_6707,N_6748);
nand U6829 (N_6829,N_6711,N_6702);
or U6830 (N_6830,N_6774,N_6775);
and U6831 (N_6831,N_6752,N_6764);
nor U6832 (N_6832,N_6753,N_6778);
nor U6833 (N_6833,N_6713,N_6791);
or U6834 (N_6834,N_6724,N_6773);
and U6835 (N_6835,N_6710,N_6704);
nor U6836 (N_6836,N_6783,N_6745);
nand U6837 (N_6837,N_6705,N_6769);
xnor U6838 (N_6838,N_6734,N_6708);
or U6839 (N_6839,N_6742,N_6793);
nor U6840 (N_6840,N_6731,N_6727);
nor U6841 (N_6841,N_6790,N_6732);
or U6842 (N_6842,N_6738,N_6766);
and U6843 (N_6843,N_6799,N_6776);
nand U6844 (N_6844,N_6740,N_6744);
nand U6845 (N_6845,N_6784,N_6750);
nand U6846 (N_6846,N_6772,N_6767);
and U6847 (N_6847,N_6762,N_6728);
nor U6848 (N_6848,N_6749,N_6701);
nand U6849 (N_6849,N_6722,N_6782);
nor U6850 (N_6850,N_6786,N_6794);
and U6851 (N_6851,N_6773,N_6720);
or U6852 (N_6852,N_6720,N_6785);
nand U6853 (N_6853,N_6738,N_6745);
or U6854 (N_6854,N_6779,N_6726);
nor U6855 (N_6855,N_6734,N_6712);
and U6856 (N_6856,N_6706,N_6704);
and U6857 (N_6857,N_6782,N_6778);
and U6858 (N_6858,N_6764,N_6744);
nand U6859 (N_6859,N_6704,N_6749);
and U6860 (N_6860,N_6709,N_6793);
and U6861 (N_6861,N_6701,N_6798);
or U6862 (N_6862,N_6795,N_6704);
nand U6863 (N_6863,N_6761,N_6739);
nand U6864 (N_6864,N_6703,N_6702);
or U6865 (N_6865,N_6738,N_6760);
or U6866 (N_6866,N_6789,N_6776);
nor U6867 (N_6867,N_6700,N_6784);
nand U6868 (N_6868,N_6727,N_6708);
and U6869 (N_6869,N_6731,N_6710);
nor U6870 (N_6870,N_6785,N_6767);
nor U6871 (N_6871,N_6797,N_6728);
and U6872 (N_6872,N_6724,N_6736);
or U6873 (N_6873,N_6725,N_6753);
nand U6874 (N_6874,N_6752,N_6788);
nand U6875 (N_6875,N_6735,N_6765);
and U6876 (N_6876,N_6716,N_6711);
nor U6877 (N_6877,N_6769,N_6764);
or U6878 (N_6878,N_6724,N_6772);
nor U6879 (N_6879,N_6748,N_6783);
and U6880 (N_6880,N_6710,N_6779);
or U6881 (N_6881,N_6733,N_6751);
and U6882 (N_6882,N_6755,N_6784);
and U6883 (N_6883,N_6779,N_6708);
xor U6884 (N_6884,N_6716,N_6709);
or U6885 (N_6885,N_6765,N_6718);
and U6886 (N_6886,N_6708,N_6725);
or U6887 (N_6887,N_6773,N_6766);
and U6888 (N_6888,N_6754,N_6797);
and U6889 (N_6889,N_6750,N_6778);
nand U6890 (N_6890,N_6782,N_6721);
nand U6891 (N_6891,N_6712,N_6788);
and U6892 (N_6892,N_6705,N_6791);
nand U6893 (N_6893,N_6739,N_6783);
or U6894 (N_6894,N_6730,N_6771);
and U6895 (N_6895,N_6736,N_6798);
nand U6896 (N_6896,N_6761,N_6707);
nand U6897 (N_6897,N_6741,N_6740);
nand U6898 (N_6898,N_6743,N_6789);
and U6899 (N_6899,N_6706,N_6770);
nor U6900 (N_6900,N_6834,N_6815);
nor U6901 (N_6901,N_6849,N_6885);
nand U6902 (N_6902,N_6839,N_6826);
nor U6903 (N_6903,N_6837,N_6846);
and U6904 (N_6904,N_6825,N_6824);
xnor U6905 (N_6905,N_6855,N_6812);
and U6906 (N_6906,N_6866,N_6879);
nor U6907 (N_6907,N_6847,N_6831);
nand U6908 (N_6908,N_6808,N_6854);
nor U6909 (N_6909,N_6873,N_6801);
or U6910 (N_6910,N_6872,N_6841);
nor U6911 (N_6911,N_6888,N_6845);
and U6912 (N_6912,N_6836,N_6862);
nor U6913 (N_6913,N_6897,N_6894);
and U6914 (N_6914,N_6829,N_6870);
or U6915 (N_6915,N_6875,N_6867);
and U6916 (N_6916,N_6817,N_6865);
nand U6917 (N_6917,N_6840,N_6800);
and U6918 (N_6918,N_6884,N_6810);
or U6919 (N_6919,N_6818,N_6887);
nor U6920 (N_6920,N_6858,N_6807);
nor U6921 (N_6921,N_6880,N_6821);
or U6922 (N_6922,N_6878,N_6848);
nand U6923 (N_6923,N_6883,N_6833);
and U6924 (N_6924,N_6899,N_6898);
nand U6925 (N_6925,N_6819,N_6835);
or U6926 (N_6926,N_6871,N_6868);
and U6927 (N_6927,N_6893,N_6843);
and U6928 (N_6928,N_6860,N_6828);
nor U6929 (N_6929,N_6822,N_6838);
xnor U6930 (N_6930,N_6851,N_6803);
and U6931 (N_6931,N_6813,N_6856);
and U6932 (N_6932,N_6877,N_6891);
and U6933 (N_6933,N_6830,N_6844);
and U6934 (N_6934,N_6852,N_6814);
nor U6935 (N_6935,N_6895,N_6853);
and U6936 (N_6936,N_6864,N_6802);
or U6937 (N_6937,N_6882,N_6850);
and U6938 (N_6938,N_6881,N_6863);
and U6939 (N_6939,N_6886,N_6874);
nand U6940 (N_6940,N_6832,N_6809);
nor U6941 (N_6941,N_6869,N_6890);
nor U6942 (N_6942,N_6892,N_6842);
and U6943 (N_6943,N_6820,N_6816);
or U6944 (N_6944,N_6827,N_6804);
and U6945 (N_6945,N_6861,N_6859);
nor U6946 (N_6946,N_6889,N_6805);
nor U6947 (N_6947,N_6811,N_6896);
nor U6948 (N_6948,N_6806,N_6876);
nor U6949 (N_6949,N_6857,N_6823);
and U6950 (N_6950,N_6875,N_6873);
nor U6951 (N_6951,N_6822,N_6846);
and U6952 (N_6952,N_6854,N_6845);
or U6953 (N_6953,N_6813,N_6865);
nor U6954 (N_6954,N_6854,N_6894);
nor U6955 (N_6955,N_6829,N_6831);
xor U6956 (N_6956,N_6863,N_6805);
nor U6957 (N_6957,N_6824,N_6802);
xor U6958 (N_6958,N_6814,N_6859);
nor U6959 (N_6959,N_6884,N_6839);
and U6960 (N_6960,N_6806,N_6809);
nand U6961 (N_6961,N_6890,N_6812);
nor U6962 (N_6962,N_6854,N_6891);
or U6963 (N_6963,N_6851,N_6853);
or U6964 (N_6964,N_6879,N_6849);
nand U6965 (N_6965,N_6870,N_6833);
or U6966 (N_6966,N_6875,N_6803);
nand U6967 (N_6967,N_6866,N_6833);
or U6968 (N_6968,N_6860,N_6813);
or U6969 (N_6969,N_6816,N_6828);
and U6970 (N_6970,N_6817,N_6866);
nor U6971 (N_6971,N_6874,N_6860);
or U6972 (N_6972,N_6837,N_6800);
or U6973 (N_6973,N_6853,N_6863);
nand U6974 (N_6974,N_6833,N_6811);
or U6975 (N_6975,N_6888,N_6847);
and U6976 (N_6976,N_6846,N_6897);
nand U6977 (N_6977,N_6870,N_6860);
and U6978 (N_6978,N_6803,N_6823);
or U6979 (N_6979,N_6891,N_6827);
or U6980 (N_6980,N_6862,N_6856);
nor U6981 (N_6981,N_6899,N_6852);
xnor U6982 (N_6982,N_6855,N_6807);
and U6983 (N_6983,N_6818,N_6800);
or U6984 (N_6984,N_6893,N_6830);
and U6985 (N_6985,N_6828,N_6802);
nor U6986 (N_6986,N_6869,N_6852);
and U6987 (N_6987,N_6845,N_6876);
or U6988 (N_6988,N_6884,N_6890);
nor U6989 (N_6989,N_6804,N_6837);
and U6990 (N_6990,N_6852,N_6812);
and U6991 (N_6991,N_6870,N_6880);
nor U6992 (N_6992,N_6851,N_6826);
and U6993 (N_6993,N_6825,N_6822);
or U6994 (N_6994,N_6826,N_6899);
or U6995 (N_6995,N_6817,N_6808);
nor U6996 (N_6996,N_6804,N_6840);
and U6997 (N_6997,N_6842,N_6899);
nand U6998 (N_6998,N_6846,N_6812);
or U6999 (N_6999,N_6877,N_6869);
nand U7000 (N_7000,N_6913,N_6955);
or U7001 (N_7001,N_6958,N_6973);
nand U7002 (N_7002,N_6921,N_6911);
or U7003 (N_7003,N_6927,N_6938);
nor U7004 (N_7004,N_6985,N_6965);
or U7005 (N_7005,N_6923,N_6989);
nor U7006 (N_7006,N_6967,N_6962);
or U7007 (N_7007,N_6988,N_6916);
or U7008 (N_7008,N_6954,N_6909);
or U7009 (N_7009,N_6978,N_6946);
nor U7010 (N_7010,N_6972,N_6977);
or U7011 (N_7011,N_6960,N_6937);
or U7012 (N_7012,N_6957,N_6915);
or U7013 (N_7013,N_6944,N_6932);
or U7014 (N_7014,N_6918,N_6941);
nor U7015 (N_7015,N_6997,N_6969);
or U7016 (N_7016,N_6994,N_6914);
nor U7017 (N_7017,N_6908,N_6948);
nand U7018 (N_7018,N_6925,N_6974);
xor U7019 (N_7019,N_6961,N_6971);
nor U7020 (N_7020,N_6963,N_6933);
or U7021 (N_7021,N_6984,N_6990);
or U7022 (N_7022,N_6917,N_6929);
nand U7023 (N_7023,N_6949,N_6953);
nor U7024 (N_7024,N_6922,N_6993);
or U7025 (N_7025,N_6980,N_6934);
nor U7026 (N_7026,N_6970,N_6919);
or U7027 (N_7027,N_6903,N_6998);
nand U7028 (N_7028,N_6995,N_6968);
or U7029 (N_7029,N_6956,N_6935);
nor U7030 (N_7030,N_6983,N_6930);
and U7031 (N_7031,N_6959,N_6991);
nand U7032 (N_7032,N_6951,N_6931);
nor U7033 (N_7033,N_6924,N_6900);
or U7034 (N_7034,N_6926,N_6947);
and U7035 (N_7035,N_6966,N_6907);
and U7036 (N_7036,N_6901,N_6992);
nor U7037 (N_7037,N_6981,N_6996);
nand U7038 (N_7038,N_6976,N_6975);
or U7039 (N_7039,N_6979,N_6939);
nor U7040 (N_7040,N_6945,N_6910);
nand U7041 (N_7041,N_6902,N_6904);
nand U7042 (N_7042,N_6999,N_6952);
nor U7043 (N_7043,N_6986,N_6928);
or U7044 (N_7044,N_6920,N_6905);
and U7045 (N_7045,N_6964,N_6940);
nor U7046 (N_7046,N_6982,N_6906);
nand U7047 (N_7047,N_6943,N_6950);
or U7048 (N_7048,N_6942,N_6987);
xor U7049 (N_7049,N_6936,N_6912);
nor U7050 (N_7050,N_6916,N_6974);
nor U7051 (N_7051,N_6998,N_6973);
and U7052 (N_7052,N_6963,N_6954);
nand U7053 (N_7053,N_6917,N_6984);
nor U7054 (N_7054,N_6982,N_6943);
and U7055 (N_7055,N_6932,N_6934);
or U7056 (N_7056,N_6909,N_6918);
and U7057 (N_7057,N_6914,N_6926);
nand U7058 (N_7058,N_6971,N_6939);
or U7059 (N_7059,N_6972,N_6989);
nor U7060 (N_7060,N_6943,N_6910);
nand U7061 (N_7061,N_6926,N_6945);
or U7062 (N_7062,N_6955,N_6963);
nor U7063 (N_7063,N_6993,N_6914);
and U7064 (N_7064,N_6951,N_6914);
nand U7065 (N_7065,N_6935,N_6984);
and U7066 (N_7066,N_6951,N_6935);
and U7067 (N_7067,N_6961,N_6999);
and U7068 (N_7068,N_6950,N_6901);
or U7069 (N_7069,N_6966,N_6999);
nor U7070 (N_7070,N_6969,N_6985);
or U7071 (N_7071,N_6993,N_6986);
or U7072 (N_7072,N_6920,N_6980);
and U7073 (N_7073,N_6976,N_6922);
or U7074 (N_7074,N_6989,N_6953);
or U7075 (N_7075,N_6976,N_6925);
nand U7076 (N_7076,N_6970,N_6942);
nor U7077 (N_7077,N_6903,N_6947);
and U7078 (N_7078,N_6972,N_6913);
nor U7079 (N_7079,N_6981,N_6921);
or U7080 (N_7080,N_6937,N_6959);
or U7081 (N_7081,N_6908,N_6991);
and U7082 (N_7082,N_6936,N_6979);
nand U7083 (N_7083,N_6985,N_6936);
or U7084 (N_7084,N_6956,N_6961);
and U7085 (N_7085,N_6959,N_6990);
and U7086 (N_7086,N_6940,N_6983);
and U7087 (N_7087,N_6938,N_6976);
xor U7088 (N_7088,N_6936,N_6904);
nor U7089 (N_7089,N_6967,N_6945);
nand U7090 (N_7090,N_6920,N_6918);
and U7091 (N_7091,N_6985,N_6955);
nor U7092 (N_7092,N_6943,N_6973);
or U7093 (N_7093,N_6934,N_6949);
or U7094 (N_7094,N_6955,N_6950);
nor U7095 (N_7095,N_6954,N_6939);
or U7096 (N_7096,N_6997,N_6925);
and U7097 (N_7097,N_6909,N_6990);
and U7098 (N_7098,N_6919,N_6954);
nor U7099 (N_7099,N_6907,N_6967);
and U7100 (N_7100,N_7040,N_7041);
nand U7101 (N_7101,N_7047,N_7097);
nand U7102 (N_7102,N_7034,N_7074);
nor U7103 (N_7103,N_7059,N_7013);
and U7104 (N_7104,N_7070,N_7081);
nor U7105 (N_7105,N_7020,N_7021);
nor U7106 (N_7106,N_7098,N_7027);
nor U7107 (N_7107,N_7011,N_7045);
nand U7108 (N_7108,N_7075,N_7035);
or U7109 (N_7109,N_7048,N_7089);
nor U7110 (N_7110,N_7024,N_7022);
nand U7111 (N_7111,N_7030,N_7001);
or U7112 (N_7112,N_7004,N_7054);
or U7113 (N_7113,N_7007,N_7071);
nand U7114 (N_7114,N_7053,N_7032);
and U7115 (N_7115,N_7087,N_7086);
nand U7116 (N_7116,N_7037,N_7039);
nand U7117 (N_7117,N_7058,N_7065);
or U7118 (N_7118,N_7029,N_7019);
and U7119 (N_7119,N_7015,N_7050);
or U7120 (N_7120,N_7008,N_7006);
nor U7121 (N_7121,N_7023,N_7061);
nand U7122 (N_7122,N_7031,N_7056);
nand U7123 (N_7123,N_7016,N_7080);
or U7124 (N_7124,N_7049,N_7018);
or U7125 (N_7125,N_7009,N_7068);
nand U7126 (N_7126,N_7063,N_7025);
and U7127 (N_7127,N_7078,N_7084);
nand U7128 (N_7128,N_7099,N_7060);
nand U7129 (N_7129,N_7091,N_7062);
nor U7130 (N_7130,N_7073,N_7083);
nor U7131 (N_7131,N_7092,N_7014);
nand U7132 (N_7132,N_7088,N_7072);
nor U7133 (N_7133,N_7093,N_7090);
nand U7134 (N_7134,N_7026,N_7038);
and U7135 (N_7135,N_7005,N_7042);
and U7136 (N_7136,N_7067,N_7028);
or U7137 (N_7137,N_7003,N_7052);
nand U7138 (N_7138,N_7000,N_7002);
and U7139 (N_7139,N_7085,N_7051);
and U7140 (N_7140,N_7036,N_7017);
and U7141 (N_7141,N_7076,N_7010);
or U7142 (N_7142,N_7066,N_7064);
nor U7143 (N_7143,N_7033,N_7046);
and U7144 (N_7144,N_7077,N_7096);
nor U7145 (N_7145,N_7057,N_7095);
nor U7146 (N_7146,N_7044,N_7069);
or U7147 (N_7147,N_7012,N_7079);
nor U7148 (N_7148,N_7082,N_7094);
nor U7149 (N_7149,N_7055,N_7043);
or U7150 (N_7150,N_7012,N_7002);
and U7151 (N_7151,N_7013,N_7098);
xnor U7152 (N_7152,N_7039,N_7001);
or U7153 (N_7153,N_7078,N_7089);
nand U7154 (N_7154,N_7040,N_7059);
nand U7155 (N_7155,N_7089,N_7057);
or U7156 (N_7156,N_7098,N_7062);
and U7157 (N_7157,N_7019,N_7041);
nor U7158 (N_7158,N_7060,N_7086);
or U7159 (N_7159,N_7017,N_7078);
and U7160 (N_7160,N_7020,N_7000);
nor U7161 (N_7161,N_7016,N_7052);
and U7162 (N_7162,N_7056,N_7083);
and U7163 (N_7163,N_7003,N_7014);
or U7164 (N_7164,N_7091,N_7053);
nor U7165 (N_7165,N_7020,N_7052);
nand U7166 (N_7166,N_7088,N_7044);
and U7167 (N_7167,N_7068,N_7051);
nand U7168 (N_7168,N_7015,N_7013);
and U7169 (N_7169,N_7040,N_7037);
or U7170 (N_7170,N_7002,N_7073);
or U7171 (N_7171,N_7010,N_7061);
and U7172 (N_7172,N_7053,N_7051);
xor U7173 (N_7173,N_7022,N_7026);
or U7174 (N_7174,N_7026,N_7000);
or U7175 (N_7175,N_7093,N_7075);
and U7176 (N_7176,N_7056,N_7092);
and U7177 (N_7177,N_7079,N_7020);
and U7178 (N_7178,N_7018,N_7091);
nand U7179 (N_7179,N_7081,N_7033);
xnor U7180 (N_7180,N_7002,N_7013);
nand U7181 (N_7181,N_7029,N_7038);
or U7182 (N_7182,N_7075,N_7041);
nor U7183 (N_7183,N_7040,N_7090);
and U7184 (N_7184,N_7062,N_7083);
and U7185 (N_7185,N_7097,N_7046);
nand U7186 (N_7186,N_7017,N_7088);
nand U7187 (N_7187,N_7004,N_7041);
and U7188 (N_7188,N_7061,N_7021);
and U7189 (N_7189,N_7059,N_7034);
or U7190 (N_7190,N_7034,N_7088);
nor U7191 (N_7191,N_7083,N_7055);
nand U7192 (N_7192,N_7011,N_7004);
and U7193 (N_7193,N_7043,N_7002);
nor U7194 (N_7194,N_7025,N_7013);
or U7195 (N_7195,N_7074,N_7076);
nor U7196 (N_7196,N_7018,N_7023);
and U7197 (N_7197,N_7090,N_7015);
xnor U7198 (N_7198,N_7071,N_7020);
nand U7199 (N_7199,N_7075,N_7022);
nor U7200 (N_7200,N_7162,N_7140);
or U7201 (N_7201,N_7100,N_7119);
nor U7202 (N_7202,N_7144,N_7173);
and U7203 (N_7203,N_7123,N_7125);
nor U7204 (N_7204,N_7155,N_7107);
and U7205 (N_7205,N_7104,N_7158);
and U7206 (N_7206,N_7116,N_7182);
nor U7207 (N_7207,N_7141,N_7166);
nor U7208 (N_7208,N_7169,N_7190);
xor U7209 (N_7209,N_7136,N_7132);
nor U7210 (N_7210,N_7124,N_7193);
nand U7211 (N_7211,N_7168,N_7131);
nand U7212 (N_7212,N_7179,N_7154);
or U7213 (N_7213,N_7114,N_7167);
xnor U7214 (N_7214,N_7194,N_7165);
or U7215 (N_7215,N_7161,N_7121);
and U7216 (N_7216,N_7110,N_7152);
nor U7217 (N_7217,N_7184,N_7151);
or U7218 (N_7218,N_7103,N_7127);
or U7219 (N_7219,N_7159,N_7102);
or U7220 (N_7220,N_7164,N_7139);
and U7221 (N_7221,N_7138,N_7192);
nor U7222 (N_7222,N_7191,N_7195);
nand U7223 (N_7223,N_7185,N_7108);
nand U7224 (N_7224,N_7115,N_7178);
or U7225 (N_7225,N_7174,N_7186);
nand U7226 (N_7226,N_7199,N_7171);
nor U7227 (N_7227,N_7122,N_7111);
or U7228 (N_7228,N_7137,N_7160);
or U7229 (N_7229,N_7106,N_7143);
or U7230 (N_7230,N_7112,N_7109);
xor U7231 (N_7231,N_7170,N_7187);
nor U7232 (N_7232,N_7145,N_7130);
and U7233 (N_7233,N_7113,N_7118);
nor U7234 (N_7234,N_7133,N_7120);
xor U7235 (N_7235,N_7135,N_7126);
nor U7236 (N_7236,N_7189,N_7176);
and U7237 (N_7237,N_7198,N_7181);
nor U7238 (N_7238,N_7156,N_7180);
nand U7239 (N_7239,N_7134,N_7197);
nand U7240 (N_7240,N_7101,N_7188);
and U7241 (N_7241,N_7183,N_7142);
nand U7242 (N_7242,N_7148,N_7149);
and U7243 (N_7243,N_7147,N_7172);
or U7244 (N_7244,N_7117,N_7177);
nand U7245 (N_7245,N_7157,N_7196);
xor U7246 (N_7246,N_7163,N_7146);
and U7247 (N_7247,N_7175,N_7153);
or U7248 (N_7248,N_7129,N_7105);
and U7249 (N_7249,N_7128,N_7150);
nand U7250 (N_7250,N_7176,N_7198);
nor U7251 (N_7251,N_7106,N_7132);
or U7252 (N_7252,N_7154,N_7120);
nor U7253 (N_7253,N_7125,N_7116);
nand U7254 (N_7254,N_7146,N_7168);
nor U7255 (N_7255,N_7154,N_7193);
and U7256 (N_7256,N_7197,N_7164);
nand U7257 (N_7257,N_7152,N_7108);
and U7258 (N_7258,N_7136,N_7142);
and U7259 (N_7259,N_7180,N_7148);
nand U7260 (N_7260,N_7114,N_7141);
nand U7261 (N_7261,N_7187,N_7139);
and U7262 (N_7262,N_7154,N_7157);
and U7263 (N_7263,N_7141,N_7128);
or U7264 (N_7264,N_7116,N_7112);
or U7265 (N_7265,N_7179,N_7161);
and U7266 (N_7266,N_7124,N_7139);
or U7267 (N_7267,N_7191,N_7126);
nor U7268 (N_7268,N_7178,N_7141);
nor U7269 (N_7269,N_7167,N_7178);
and U7270 (N_7270,N_7155,N_7194);
xor U7271 (N_7271,N_7102,N_7189);
xor U7272 (N_7272,N_7115,N_7150);
nand U7273 (N_7273,N_7123,N_7155);
nor U7274 (N_7274,N_7116,N_7162);
nor U7275 (N_7275,N_7121,N_7195);
and U7276 (N_7276,N_7100,N_7177);
nand U7277 (N_7277,N_7173,N_7197);
nand U7278 (N_7278,N_7143,N_7146);
and U7279 (N_7279,N_7199,N_7132);
nor U7280 (N_7280,N_7132,N_7144);
and U7281 (N_7281,N_7176,N_7155);
nor U7282 (N_7282,N_7152,N_7196);
or U7283 (N_7283,N_7188,N_7144);
and U7284 (N_7284,N_7131,N_7164);
or U7285 (N_7285,N_7114,N_7128);
or U7286 (N_7286,N_7170,N_7186);
and U7287 (N_7287,N_7171,N_7145);
and U7288 (N_7288,N_7165,N_7180);
or U7289 (N_7289,N_7142,N_7115);
nor U7290 (N_7290,N_7129,N_7178);
or U7291 (N_7291,N_7171,N_7134);
nand U7292 (N_7292,N_7190,N_7111);
nor U7293 (N_7293,N_7111,N_7159);
xnor U7294 (N_7294,N_7152,N_7160);
or U7295 (N_7295,N_7107,N_7189);
nor U7296 (N_7296,N_7108,N_7198);
nor U7297 (N_7297,N_7137,N_7143);
nand U7298 (N_7298,N_7139,N_7199);
nor U7299 (N_7299,N_7106,N_7117);
nand U7300 (N_7300,N_7240,N_7286);
and U7301 (N_7301,N_7229,N_7233);
and U7302 (N_7302,N_7221,N_7218);
nor U7303 (N_7303,N_7255,N_7282);
nand U7304 (N_7304,N_7242,N_7291);
and U7305 (N_7305,N_7281,N_7214);
or U7306 (N_7306,N_7292,N_7200);
or U7307 (N_7307,N_7283,N_7275);
nor U7308 (N_7308,N_7208,N_7236);
nand U7309 (N_7309,N_7257,N_7266);
and U7310 (N_7310,N_7213,N_7243);
and U7311 (N_7311,N_7270,N_7256);
nor U7312 (N_7312,N_7272,N_7210);
or U7313 (N_7313,N_7224,N_7238);
xnor U7314 (N_7314,N_7290,N_7299);
or U7315 (N_7315,N_7293,N_7220);
and U7316 (N_7316,N_7264,N_7217);
or U7317 (N_7317,N_7279,N_7274);
or U7318 (N_7318,N_7215,N_7297);
and U7319 (N_7319,N_7262,N_7204);
nand U7320 (N_7320,N_7244,N_7294);
nor U7321 (N_7321,N_7280,N_7260);
nor U7322 (N_7322,N_7237,N_7268);
or U7323 (N_7323,N_7246,N_7223);
and U7324 (N_7324,N_7209,N_7230);
and U7325 (N_7325,N_7235,N_7206);
nand U7326 (N_7326,N_7285,N_7228);
xor U7327 (N_7327,N_7271,N_7267);
xnor U7328 (N_7328,N_7239,N_7247);
nor U7329 (N_7329,N_7278,N_7254);
and U7330 (N_7330,N_7205,N_7245);
and U7331 (N_7331,N_7219,N_7207);
or U7332 (N_7332,N_7277,N_7227);
nor U7333 (N_7333,N_7250,N_7203);
and U7334 (N_7334,N_7216,N_7248);
xor U7335 (N_7335,N_7212,N_7253);
nand U7336 (N_7336,N_7269,N_7211);
or U7337 (N_7337,N_7265,N_7241);
nor U7338 (N_7338,N_7234,N_7273);
nor U7339 (N_7339,N_7276,N_7261);
and U7340 (N_7340,N_7252,N_7263);
or U7341 (N_7341,N_7202,N_7296);
nand U7342 (N_7342,N_7298,N_7288);
nand U7343 (N_7343,N_7226,N_7232);
and U7344 (N_7344,N_7258,N_7231);
and U7345 (N_7345,N_7259,N_7222);
nand U7346 (N_7346,N_7249,N_7289);
nor U7347 (N_7347,N_7201,N_7284);
nor U7348 (N_7348,N_7287,N_7251);
nand U7349 (N_7349,N_7225,N_7295);
or U7350 (N_7350,N_7294,N_7270);
nor U7351 (N_7351,N_7207,N_7237);
or U7352 (N_7352,N_7222,N_7216);
or U7353 (N_7353,N_7213,N_7261);
or U7354 (N_7354,N_7280,N_7293);
nor U7355 (N_7355,N_7203,N_7246);
and U7356 (N_7356,N_7214,N_7232);
nor U7357 (N_7357,N_7256,N_7216);
nand U7358 (N_7358,N_7228,N_7274);
nor U7359 (N_7359,N_7293,N_7215);
xor U7360 (N_7360,N_7267,N_7241);
and U7361 (N_7361,N_7260,N_7240);
and U7362 (N_7362,N_7226,N_7223);
or U7363 (N_7363,N_7293,N_7236);
nand U7364 (N_7364,N_7234,N_7257);
nand U7365 (N_7365,N_7257,N_7291);
nand U7366 (N_7366,N_7225,N_7293);
and U7367 (N_7367,N_7223,N_7231);
or U7368 (N_7368,N_7230,N_7222);
xor U7369 (N_7369,N_7272,N_7234);
nand U7370 (N_7370,N_7260,N_7237);
nor U7371 (N_7371,N_7205,N_7253);
nor U7372 (N_7372,N_7215,N_7233);
nand U7373 (N_7373,N_7250,N_7287);
nand U7374 (N_7374,N_7270,N_7289);
or U7375 (N_7375,N_7276,N_7246);
and U7376 (N_7376,N_7243,N_7286);
and U7377 (N_7377,N_7237,N_7288);
nand U7378 (N_7378,N_7230,N_7276);
and U7379 (N_7379,N_7282,N_7277);
or U7380 (N_7380,N_7257,N_7242);
or U7381 (N_7381,N_7250,N_7226);
or U7382 (N_7382,N_7206,N_7273);
nor U7383 (N_7383,N_7295,N_7252);
nor U7384 (N_7384,N_7201,N_7279);
or U7385 (N_7385,N_7218,N_7207);
nor U7386 (N_7386,N_7241,N_7287);
or U7387 (N_7387,N_7265,N_7205);
or U7388 (N_7388,N_7217,N_7294);
nand U7389 (N_7389,N_7237,N_7241);
xnor U7390 (N_7390,N_7261,N_7210);
and U7391 (N_7391,N_7213,N_7257);
nand U7392 (N_7392,N_7283,N_7208);
or U7393 (N_7393,N_7239,N_7283);
nor U7394 (N_7394,N_7244,N_7259);
nor U7395 (N_7395,N_7288,N_7201);
nor U7396 (N_7396,N_7209,N_7276);
and U7397 (N_7397,N_7245,N_7295);
or U7398 (N_7398,N_7264,N_7241);
xnor U7399 (N_7399,N_7257,N_7295);
nor U7400 (N_7400,N_7396,N_7338);
and U7401 (N_7401,N_7374,N_7321);
nor U7402 (N_7402,N_7317,N_7389);
nand U7403 (N_7403,N_7346,N_7367);
nand U7404 (N_7404,N_7364,N_7327);
or U7405 (N_7405,N_7379,N_7319);
or U7406 (N_7406,N_7391,N_7304);
or U7407 (N_7407,N_7365,N_7324);
and U7408 (N_7408,N_7395,N_7308);
nand U7409 (N_7409,N_7376,N_7325);
nand U7410 (N_7410,N_7310,N_7353);
and U7411 (N_7411,N_7323,N_7378);
nor U7412 (N_7412,N_7345,N_7300);
nand U7413 (N_7413,N_7326,N_7383);
and U7414 (N_7414,N_7301,N_7390);
or U7415 (N_7415,N_7316,N_7388);
and U7416 (N_7416,N_7348,N_7320);
nor U7417 (N_7417,N_7344,N_7352);
nor U7418 (N_7418,N_7386,N_7372);
and U7419 (N_7419,N_7394,N_7380);
nand U7420 (N_7420,N_7358,N_7303);
nor U7421 (N_7421,N_7315,N_7349);
or U7422 (N_7422,N_7328,N_7375);
nand U7423 (N_7423,N_7351,N_7318);
or U7424 (N_7424,N_7363,N_7336);
nand U7425 (N_7425,N_7399,N_7360);
nor U7426 (N_7426,N_7361,N_7312);
and U7427 (N_7427,N_7357,N_7354);
or U7428 (N_7428,N_7392,N_7382);
nand U7429 (N_7429,N_7333,N_7398);
nor U7430 (N_7430,N_7332,N_7387);
xor U7431 (N_7431,N_7342,N_7355);
and U7432 (N_7432,N_7368,N_7340);
nor U7433 (N_7433,N_7322,N_7331);
nand U7434 (N_7434,N_7359,N_7377);
or U7435 (N_7435,N_7371,N_7311);
nor U7436 (N_7436,N_7347,N_7329);
nand U7437 (N_7437,N_7337,N_7381);
nor U7438 (N_7438,N_7307,N_7373);
nor U7439 (N_7439,N_7339,N_7384);
nand U7440 (N_7440,N_7350,N_7335);
nor U7441 (N_7441,N_7313,N_7314);
or U7442 (N_7442,N_7397,N_7334);
nand U7443 (N_7443,N_7343,N_7362);
nor U7444 (N_7444,N_7306,N_7369);
nor U7445 (N_7445,N_7366,N_7341);
and U7446 (N_7446,N_7385,N_7370);
or U7447 (N_7447,N_7330,N_7356);
and U7448 (N_7448,N_7305,N_7393);
nor U7449 (N_7449,N_7309,N_7302);
nor U7450 (N_7450,N_7374,N_7361);
and U7451 (N_7451,N_7346,N_7344);
or U7452 (N_7452,N_7328,N_7373);
nand U7453 (N_7453,N_7361,N_7397);
nor U7454 (N_7454,N_7376,N_7383);
and U7455 (N_7455,N_7319,N_7364);
nand U7456 (N_7456,N_7354,N_7343);
and U7457 (N_7457,N_7372,N_7332);
and U7458 (N_7458,N_7386,N_7332);
or U7459 (N_7459,N_7353,N_7337);
or U7460 (N_7460,N_7338,N_7360);
nor U7461 (N_7461,N_7314,N_7302);
and U7462 (N_7462,N_7398,N_7379);
or U7463 (N_7463,N_7377,N_7334);
or U7464 (N_7464,N_7333,N_7304);
and U7465 (N_7465,N_7385,N_7382);
or U7466 (N_7466,N_7313,N_7343);
nor U7467 (N_7467,N_7309,N_7356);
or U7468 (N_7468,N_7367,N_7320);
nor U7469 (N_7469,N_7354,N_7326);
and U7470 (N_7470,N_7330,N_7379);
nand U7471 (N_7471,N_7375,N_7315);
or U7472 (N_7472,N_7399,N_7347);
nand U7473 (N_7473,N_7362,N_7348);
nor U7474 (N_7474,N_7312,N_7338);
and U7475 (N_7475,N_7378,N_7310);
or U7476 (N_7476,N_7356,N_7316);
nand U7477 (N_7477,N_7378,N_7392);
nand U7478 (N_7478,N_7328,N_7325);
xnor U7479 (N_7479,N_7300,N_7308);
or U7480 (N_7480,N_7346,N_7395);
or U7481 (N_7481,N_7324,N_7342);
nor U7482 (N_7482,N_7399,N_7325);
nor U7483 (N_7483,N_7333,N_7328);
or U7484 (N_7484,N_7330,N_7393);
nand U7485 (N_7485,N_7338,N_7358);
nor U7486 (N_7486,N_7326,N_7391);
nand U7487 (N_7487,N_7320,N_7324);
or U7488 (N_7488,N_7369,N_7365);
nor U7489 (N_7489,N_7376,N_7397);
nor U7490 (N_7490,N_7335,N_7317);
and U7491 (N_7491,N_7393,N_7335);
and U7492 (N_7492,N_7380,N_7316);
or U7493 (N_7493,N_7368,N_7303);
nand U7494 (N_7494,N_7338,N_7307);
and U7495 (N_7495,N_7313,N_7342);
or U7496 (N_7496,N_7364,N_7392);
nor U7497 (N_7497,N_7336,N_7317);
or U7498 (N_7498,N_7391,N_7318);
nand U7499 (N_7499,N_7374,N_7343);
nand U7500 (N_7500,N_7479,N_7470);
or U7501 (N_7501,N_7402,N_7421);
or U7502 (N_7502,N_7484,N_7443);
and U7503 (N_7503,N_7465,N_7423);
nor U7504 (N_7504,N_7488,N_7461);
and U7505 (N_7505,N_7434,N_7477);
nand U7506 (N_7506,N_7401,N_7440);
nor U7507 (N_7507,N_7493,N_7472);
and U7508 (N_7508,N_7432,N_7403);
or U7509 (N_7509,N_7438,N_7408);
or U7510 (N_7510,N_7492,N_7439);
xnor U7511 (N_7511,N_7415,N_7485);
or U7512 (N_7512,N_7483,N_7495);
or U7513 (N_7513,N_7499,N_7441);
and U7514 (N_7514,N_7427,N_7453);
or U7515 (N_7515,N_7422,N_7425);
nand U7516 (N_7516,N_7406,N_7436);
and U7517 (N_7517,N_7450,N_7400);
or U7518 (N_7518,N_7429,N_7491);
or U7519 (N_7519,N_7431,N_7433);
and U7520 (N_7520,N_7418,N_7444);
nor U7521 (N_7521,N_7469,N_7486);
nand U7522 (N_7522,N_7458,N_7466);
or U7523 (N_7523,N_7471,N_7409);
or U7524 (N_7524,N_7480,N_7455);
nor U7525 (N_7525,N_7481,N_7426);
nand U7526 (N_7526,N_7462,N_7478);
nor U7527 (N_7527,N_7489,N_7487);
and U7528 (N_7528,N_7405,N_7474);
nand U7529 (N_7529,N_7467,N_7437);
and U7530 (N_7530,N_7473,N_7490);
or U7531 (N_7531,N_7417,N_7413);
nand U7532 (N_7532,N_7464,N_7445);
nor U7533 (N_7533,N_7446,N_7496);
and U7534 (N_7534,N_7463,N_7416);
nand U7535 (N_7535,N_7414,N_7442);
or U7536 (N_7536,N_7424,N_7460);
and U7537 (N_7537,N_7457,N_7449);
or U7538 (N_7538,N_7420,N_7451);
nand U7539 (N_7539,N_7419,N_7410);
nor U7540 (N_7540,N_7407,N_7428);
and U7541 (N_7541,N_7494,N_7412);
nor U7542 (N_7542,N_7456,N_7475);
and U7543 (N_7543,N_7430,N_7468);
nand U7544 (N_7544,N_7498,N_7411);
nor U7545 (N_7545,N_7452,N_7476);
and U7546 (N_7546,N_7482,N_7454);
or U7547 (N_7547,N_7448,N_7497);
nor U7548 (N_7548,N_7435,N_7459);
or U7549 (N_7549,N_7404,N_7447);
nand U7550 (N_7550,N_7423,N_7439);
or U7551 (N_7551,N_7428,N_7409);
and U7552 (N_7552,N_7484,N_7418);
or U7553 (N_7553,N_7496,N_7423);
nor U7554 (N_7554,N_7409,N_7452);
nor U7555 (N_7555,N_7477,N_7459);
nand U7556 (N_7556,N_7433,N_7442);
nor U7557 (N_7557,N_7458,N_7426);
or U7558 (N_7558,N_7496,N_7411);
or U7559 (N_7559,N_7456,N_7448);
nand U7560 (N_7560,N_7489,N_7450);
nor U7561 (N_7561,N_7454,N_7491);
nand U7562 (N_7562,N_7480,N_7410);
nor U7563 (N_7563,N_7403,N_7482);
and U7564 (N_7564,N_7433,N_7413);
or U7565 (N_7565,N_7464,N_7425);
nand U7566 (N_7566,N_7477,N_7458);
and U7567 (N_7567,N_7438,N_7490);
and U7568 (N_7568,N_7419,N_7496);
and U7569 (N_7569,N_7448,N_7428);
or U7570 (N_7570,N_7402,N_7446);
or U7571 (N_7571,N_7473,N_7440);
nand U7572 (N_7572,N_7416,N_7456);
or U7573 (N_7573,N_7401,N_7416);
and U7574 (N_7574,N_7443,N_7482);
nor U7575 (N_7575,N_7459,N_7420);
nand U7576 (N_7576,N_7499,N_7487);
and U7577 (N_7577,N_7435,N_7461);
nor U7578 (N_7578,N_7466,N_7474);
or U7579 (N_7579,N_7437,N_7454);
or U7580 (N_7580,N_7431,N_7430);
and U7581 (N_7581,N_7435,N_7412);
nor U7582 (N_7582,N_7416,N_7440);
or U7583 (N_7583,N_7465,N_7462);
xnor U7584 (N_7584,N_7443,N_7416);
nor U7585 (N_7585,N_7430,N_7405);
nand U7586 (N_7586,N_7433,N_7437);
nand U7587 (N_7587,N_7408,N_7470);
nor U7588 (N_7588,N_7470,N_7452);
or U7589 (N_7589,N_7487,N_7431);
and U7590 (N_7590,N_7467,N_7498);
and U7591 (N_7591,N_7421,N_7419);
nand U7592 (N_7592,N_7487,N_7437);
and U7593 (N_7593,N_7420,N_7455);
nand U7594 (N_7594,N_7415,N_7477);
nor U7595 (N_7595,N_7412,N_7472);
nand U7596 (N_7596,N_7444,N_7479);
nor U7597 (N_7597,N_7488,N_7428);
nor U7598 (N_7598,N_7483,N_7476);
and U7599 (N_7599,N_7400,N_7477);
and U7600 (N_7600,N_7568,N_7545);
or U7601 (N_7601,N_7505,N_7593);
and U7602 (N_7602,N_7595,N_7575);
or U7603 (N_7603,N_7586,N_7565);
and U7604 (N_7604,N_7596,N_7589);
and U7605 (N_7605,N_7539,N_7522);
nand U7606 (N_7606,N_7562,N_7580);
or U7607 (N_7607,N_7532,N_7518);
nand U7608 (N_7608,N_7517,N_7546);
and U7609 (N_7609,N_7525,N_7579);
nor U7610 (N_7610,N_7547,N_7503);
nand U7611 (N_7611,N_7566,N_7561);
or U7612 (N_7612,N_7585,N_7536);
nand U7613 (N_7613,N_7571,N_7512);
xor U7614 (N_7614,N_7557,N_7513);
and U7615 (N_7615,N_7543,N_7581);
nor U7616 (N_7616,N_7515,N_7569);
nand U7617 (N_7617,N_7552,N_7540);
nor U7618 (N_7618,N_7519,N_7576);
nor U7619 (N_7619,N_7526,N_7502);
nand U7620 (N_7620,N_7553,N_7507);
xor U7621 (N_7621,N_7599,N_7572);
nor U7622 (N_7622,N_7570,N_7506);
or U7623 (N_7623,N_7584,N_7583);
or U7624 (N_7624,N_7542,N_7544);
and U7625 (N_7625,N_7582,N_7531);
nor U7626 (N_7626,N_7578,N_7510);
and U7627 (N_7627,N_7520,N_7509);
nand U7628 (N_7628,N_7591,N_7527);
nand U7629 (N_7629,N_7516,N_7551);
or U7630 (N_7630,N_7533,N_7554);
or U7631 (N_7631,N_7559,N_7592);
nand U7632 (N_7632,N_7538,N_7594);
and U7633 (N_7633,N_7588,N_7534);
nand U7634 (N_7634,N_7555,N_7529);
nor U7635 (N_7635,N_7577,N_7528);
and U7636 (N_7636,N_7587,N_7560);
nor U7637 (N_7637,N_7537,N_7564);
nor U7638 (N_7638,N_7597,N_7567);
or U7639 (N_7639,N_7573,N_7511);
nor U7640 (N_7640,N_7558,N_7541);
nand U7641 (N_7641,N_7549,N_7550);
and U7642 (N_7642,N_7504,N_7548);
nor U7643 (N_7643,N_7524,N_7521);
nor U7644 (N_7644,N_7501,N_7514);
or U7645 (N_7645,N_7563,N_7500);
nand U7646 (N_7646,N_7523,N_7598);
nand U7647 (N_7647,N_7556,N_7508);
or U7648 (N_7648,N_7535,N_7574);
nor U7649 (N_7649,N_7530,N_7590);
nor U7650 (N_7650,N_7583,N_7550);
nand U7651 (N_7651,N_7592,N_7574);
nand U7652 (N_7652,N_7552,N_7520);
and U7653 (N_7653,N_7575,N_7551);
nor U7654 (N_7654,N_7563,N_7588);
or U7655 (N_7655,N_7563,N_7508);
or U7656 (N_7656,N_7503,N_7555);
nor U7657 (N_7657,N_7555,N_7596);
and U7658 (N_7658,N_7534,N_7579);
nor U7659 (N_7659,N_7507,N_7581);
xor U7660 (N_7660,N_7574,N_7533);
or U7661 (N_7661,N_7597,N_7570);
nand U7662 (N_7662,N_7544,N_7553);
nor U7663 (N_7663,N_7504,N_7552);
and U7664 (N_7664,N_7595,N_7529);
and U7665 (N_7665,N_7525,N_7534);
nor U7666 (N_7666,N_7541,N_7500);
and U7667 (N_7667,N_7530,N_7580);
nand U7668 (N_7668,N_7564,N_7576);
or U7669 (N_7669,N_7516,N_7575);
nor U7670 (N_7670,N_7515,N_7576);
and U7671 (N_7671,N_7525,N_7582);
or U7672 (N_7672,N_7523,N_7507);
or U7673 (N_7673,N_7580,N_7510);
xor U7674 (N_7674,N_7546,N_7568);
xor U7675 (N_7675,N_7560,N_7590);
and U7676 (N_7676,N_7515,N_7519);
nand U7677 (N_7677,N_7555,N_7523);
nand U7678 (N_7678,N_7511,N_7563);
nor U7679 (N_7679,N_7587,N_7504);
nand U7680 (N_7680,N_7517,N_7524);
nand U7681 (N_7681,N_7535,N_7517);
and U7682 (N_7682,N_7540,N_7597);
nor U7683 (N_7683,N_7548,N_7529);
or U7684 (N_7684,N_7555,N_7592);
nor U7685 (N_7685,N_7563,N_7570);
nand U7686 (N_7686,N_7551,N_7541);
or U7687 (N_7687,N_7549,N_7521);
and U7688 (N_7688,N_7508,N_7526);
and U7689 (N_7689,N_7500,N_7596);
and U7690 (N_7690,N_7539,N_7556);
and U7691 (N_7691,N_7582,N_7528);
and U7692 (N_7692,N_7554,N_7546);
nor U7693 (N_7693,N_7524,N_7587);
and U7694 (N_7694,N_7561,N_7548);
nand U7695 (N_7695,N_7501,N_7554);
or U7696 (N_7696,N_7558,N_7527);
nand U7697 (N_7697,N_7546,N_7561);
and U7698 (N_7698,N_7580,N_7520);
or U7699 (N_7699,N_7509,N_7573);
and U7700 (N_7700,N_7644,N_7666);
or U7701 (N_7701,N_7659,N_7636);
or U7702 (N_7702,N_7650,N_7699);
nor U7703 (N_7703,N_7693,N_7660);
or U7704 (N_7704,N_7678,N_7611);
nor U7705 (N_7705,N_7661,N_7604);
and U7706 (N_7706,N_7608,N_7691);
nor U7707 (N_7707,N_7663,N_7600);
nand U7708 (N_7708,N_7641,N_7623);
or U7709 (N_7709,N_7645,N_7655);
or U7710 (N_7710,N_7673,N_7610);
and U7711 (N_7711,N_7648,N_7629);
or U7712 (N_7712,N_7690,N_7643);
and U7713 (N_7713,N_7689,N_7697);
or U7714 (N_7714,N_7632,N_7620);
and U7715 (N_7715,N_7627,N_7621);
and U7716 (N_7716,N_7686,N_7683);
nand U7717 (N_7717,N_7625,N_7667);
or U7718 (N_7718,N_7649,N_7635);
nand U7719 (N_7719,N_7642,N_7616);
nand U7720 (N_7720,N_7630,N_7646);
and U7721 (N_7721,N_7612,N_7607);
nor U7722 (N_7722,N_7652,N_7609);
nor U7723 (N_7723,N_7613,N_7688);
or U7724 (N_7724,N_7692,N_7617);
and U7725 (N_7725,N_7681,N_7638);
xor U7726 (N_7726,N_7624,N_7694);
or U7727 (N_7727,N_7679,N_7658);
nand U7728 (N_7728,N_7605,N_7614);
nor U7729 (N_7729,N_7626,N_7672);
nor U7730 (N_7730,N_7631,N_7619);
or U7731 (N_7731,N_7671,N_7695);
nor U7732 (N_7732,N_7675,N_7639);
nor U7733 (N_7733,N_7628,N_7677);
nor U7734 (N_7734,N_7676,N_7601);
or U7735 (N_7735,N_7682,N_7640);
nand U7736 (N_7736,N_7687,N_7662);
nor U7737 (N_7737,N_7606,N_7647);
nand U7738 (N_7738,N_7668,N_7654);
or U7739 (N_7739,N_7696,N_7633);
xnor U7740 (N_7740,N_7618,N_7669);
nand U7741 (N_7741,N_7653,N_7684);
nand U7742 (N_7742,N_7680,N_7664);
nor U7743 (N_7743,N_7685,N_7657);
xor U7744 (N_7744,N_7656,N_7674);
nor U7745 (N_7745,N_7665,N_7634);
nor U7746 (N_7746,N_7602,N_7670);
or U7747 (N_7747,N_7615,N_7651);
nor U7748 (N_7748,N_7698,N_7637);
nand U7749 (N_7749,N_7603,N_7622);
or U7750 (N_7750,N_7652,N_7675);
or U7751 (N_7751,N_7604,N_7673);
nor U7752 (N_7752,N_7638,N_7694);
nor U7753 (N_7753,N_7665,N_7691);
or U7754 (N_7754,N_7649,N_7657);
nor U7755 (N_7755,N_7652,N_7650);
nor U7756 (N_7756,N_7680,N_7604);
nand U7757 (N_7757,N_7623,N_7619);
nand U7758 (N_7758,N_7624,N_7648);
nor U7759 (N_7759,N_7699,N_7649);
or U7760 (N_7760,N_7675,N_7610);
nor U7761 (N_7761,N_7646,N_7685);
nor U7762 (N_7762,N_7628,N_7634);
nand U7763 (N_7763,N_7615,N_7654);
and U7764 (N_7764,N_7657,N_7637);
and U7765 (N_7765,N_7661,N_7693);
nand U7766 (N_7766,N_7666,N_7674);
or U7767 (N_7767,N_7615,N_7618);
and U7768 (N_7768,N_7666,N_7662);
and U7769 (N_7769,N_7655,N_7610);
nor U7770 (N_7770,N_7634,N_7699);
nand U7771 (N_7771,N_7683,N_7630);
and U7772 (N_7772,N_7651,N_7658);
or U7773 (N_7773,N_7656,N_7669);
and U7774 (N_7774,N_7658,N_7630);
nor U7775 (N_7775,N_7634,N_7663);
nand U7776 (N_7776,N_7634,N_7636);
nor U7777 (N_7777,N_7643,N_7620);
and U7778 (N_7778,N_7607,N_7686);
nor U7779 (N_7779,N_7665,N_7698);
nor U7780 (N_7780,N_7608,N_7624);
or U7781 (N_7781,N_7657,N_7688);
or U7782 (N_7782,N_7630,N_7653);
and U7783 (N_7783,N_7650,N_7690);
nand U7784 (N_7784,N_7684,N_7643);
nor U7785 (N_7785,N_7629,N_7686);
or U7786 (N_7786,N_7637,N_7672);
or U7787 (N_7787,N_7609,N_7691);
and U7788 (N_7788,N_7631,N_7651);
or U7789 (N_7789,N_7648,N_7673);
nor U7790 (N_7790,N_7699,N_7683);
nor U7791 (N_7791,N_7647,N_7679);
nand U7792 (N_7792,N_7621,N_7697);
xor U7793 (N_7793,N_7694,N_7605);
and U7794 (N_7794,N_7672,N_7650);
nor U7795 (N_7795,N_7697,N_7686);
nand U7796 (N_7796,N_7614,N_7679);
and U7797 (N_7797,N_7625,N_7604);
or U7798 (N_7798,N_7630,N_7609);
nor U7799 (N_7799,N_7661,N_7639);
nor U7800 (N_7800,N_7769,N_7794);
and U7801 (N_7801,N_7745,N_7766);
nand U7802 (N_7802,N_7702,N_7761);
or U7803 (N_7803,N_7726,N_7759);
or U7804 (N_7804,N_7728,N_7729);
and U7805 (N_7805,N_7723,N_7760);
or U7806 (N_7806,N_7724,N_7756);
and U7807 (N_7807,N_7700,N_7793);
or U7808 (N_7808,N_7734,N_7709);
and U7809 (N_7809,N_7784,N_7764);
nor U7810 (N_7810,N_7713,N_7785);
nor U7811 (N_7811,N_7742,N_7767);
nand U7812 (N_7812,N_7791,N_7787);
nand U7813 (N_7813,N_7733,N_7750);
nand U7814 (N_7814,N_7735,N_7779);
nor U7815 (N_7815,N_7722,N_7738);
xor U7816 (N_7816,N_7708,N_7762);
or U7817 (N_7817,N_7725,N_7707);
and U7818 (N_7818,N_7703,N_7792);
and U7819 (N_7819,N_7798,N_7739);
or U7820 (N_7820,N_7719,N_7711);
nor U7821 (N_7821,N_7797,N_7776);
nand U7822 (N_7822,N_7753,N_7746);
or U7823 (N_7823,N_7768,N_7757);
or U7824 (N_7824,N_7718,N_7775);
xnor U7825 (N_7825,N_7789,N_7790);
nand U7826 (N_7826,N_7727,N_7772);
or U7827 (N_7827,N_7773,N_7783);
nand U7828 (N_7828,N_7736,N_7770);
or U7829 (N_7829,N_7737,N_7705);
nand U7830 (N_7830,N_7799,N_7740);
xor U7831 (N_7831,N_7765,N_7782);
nand U7832 (N_7832,N_7715,N_7781);
and U7833 (N_7833,N_7780,N_7754);
and U7834 (N_7834,N_7795,N_7796);
nor U7835 (N_7835,N_7706,N_7758);
nand U7836 (N_7836,N_7747,N_7788);
and U7837 (N_7837,N_7771,N_7763);
and U7838 (N_7838,N_7717,N_7755);
nor U7839 (N_7839,N_7752,N_7774);
nor U7840 (N_7840,N_7749,N_7741);
nand U7841 (N_7841,N_7704,N_7786);
and U7842 (N_7842,N_7744,N_7732);
nor U7843 (N_7843,N_7731,N_7743);
nor U7844 (N_7844,N_7730,N_7721);
xor U7845 (N_7845,N_7777,N_7778);
or U7846 (N_7846,N_7751,N_7716);
and U7847 (N_7847,N_7714,N_7710);
nor U7848 (N_7848,N_7701,N_7712);
or U7849 (N_7849,N_7720,N_7748);
nor U7850 (N_7850,N_7772,N_7717);
or U7851 (N_7851,N_7724,N_7716);
nor U7852 (N_7852,N_7763,N_7724);
or U7853 (N_7853,N_7735,N_7790);
or U7854 (N_7854,N_7716,N_7752);
nand U7855 (N_7855,N_7737,N_7754);
nand U7856 (N_7856,N_7723,N_7767);
nand U7857 (N_7857,N_7742,N_7785);
nor U7858 (N_7858,N_7733,N_7764);
or U7859 (N_7859,N_7747,N_7797);
or U7860 (N_7860,N_7732,N_7710);
or U7861 (N_7861,N_7785,N_7788);
nor U7862 (N_7862,N_7782,N_7701);
nor U7863 (N_7863,N_7717,N_7783);
nand U7864 (N_7864,N_7799,N_7754);
and U7865 (N_7865,N_7728,N_7772);
nand U7866 (N_7866,N_7705,N_7717);
and U7867 (N_7867,N_7766,N_7765);
or U7868 (N_7868,N_7707,N_7793);
nor U7869 (N_7869,N_7742,N_7714);
nor U7870 (N_7870,N_7763,N_7762);
nor U7871 (N_7871,N_7787,N_7735);
and U7872 (N_7872,N_7703,N_7765);
nand U7873 (N_7873,N_7743,N_7784);
nand U7874 (N_7874,N_7710,N_7716);
nand U7875 (N_7875,N_7788,N_7797);
and U7876 (N_7876,N_7700,N_7711);
nor U7877 (N_7877,N_7784,N_7728);
nor U7878 (N_7878,N_7761,N_7797);
nor U7879 (N_7879,N_7709,N_7764);
or U7880 (N_7880,N_7717,N_7792);
or U7881 (N_7881,N_7786,N_7797);
and U7882 (N_7882,N_7777,N_7768);
or U7883 (N_7883,N_7727,N_7721);
nor U7884 (N_7884,N_7786,N_7726);
or U7885 (N_7885,N_7766,N_7722);
nor U7886 (N_7886,N_7713,N_7789);
and U7887 (N_7887,N_7703,N_7771);
or U7888 (N_7888,N_7750,N_7701);
nor U7889 (N_7889,N_7711,N_7796);
nor U7890 (N_7890,N_7776,N_7751);
nor U7891 (N_7891,N_7751,N_7790);
xnor U7892 (N_7892,N_7760,N_7759);
or U7893 (N_7893,N_7792,N_7787);
or U7894 (N_7894,N_7712,N_7736);
or U7895 (N_7895,N_7708,N_7715);
or U7896 (N_7896,N_7754,N_7795);
and U7897 (N_7897,N_7700,N_7778);
nand U7898 (N_7898,N_7707,N_7732);
and U7899 (N_7899,N_7704,N_7749);
or U7900 (N_7900,N_7867,N_7897);
nand U7901 (N_7901,N_7806,N_7813);
nor U7902 (N_7902,N_7820,N_7875);
or U7903 (N_7903,N_7825,N_7849);
and U7904 (N_7904,N_7848,N_7882);
and U7905 (N_7905,N_7835,N_7870);
nor U7906 (N_7906,N_7893,N_7840);
nand U7907 (N_7907,N_7803,N_7886);
nor U7908 (N_7908,N_7843,N_7890);
or U7909 (N_7909,N_7853,N_7811);
and U7910 (N_7910,N_7857,N_7823);
nor U7911 (N_7911,N_7880,N_7898);
and U7912 (N_7912,N_7829,N_7885);
nand U7913 (N_7913,N_7850,N_7845);
nand U7914 (N_7914,N_7846,N_7865);
and U7915 (N_7915,N_7896,N_7805);
and U7916 (N_7916,N_7810,N_7858);
or U7917 (N_7917,N_7891,N_7837);
xnor U7918 (N_7918,N_7879,N_7872);
xor U7919 (N_7919,N_7808,N_7873);
nand U7920 (N_7920,N_7877,N_7856);
nor U7921 (N_7921,N_7809,N_7859);
or U7922 (N_7922,N_7801,N_7855);
nor U7923 (N_7923,N_7826,N_7844);
nand U7924 (N_7924,N_7861,N_7815);
nor U7925 (N_7925,N_7804,N_7830);
nor U7926 (N_7926,N_7812,N_7868);
nor U7927 (N_7927,N_7822,N_7802);
or U7928 (N_7928,N_7838,N_7828);
or U7929 (N_7929,N_7866,N_7827);
or U7930 (N_7930,N_7841,N_7854);
or U7931 (N_7931,N_7869,N_7833);
and U7932 (N_7932,N_7895,N_7874);
and U7933 (N_7933,N_7836,N_7842);
nor U7934 (N_7934,N_7894,N_7824);
and U7935 (N_7935,N_7871,N_7887);
nor U7936 (N_7936,N_7817,N_7819);
nor U7937 (N_7937,N_7888,N_7800);
or U7938 (N_7938,N_7832,N_7847);
and U7939 (N_7939,N_7899,N_7839);
nand U7940 (N_7940,N_7816,N_7862);
or U7941 (N_7941,N_7878,N_7814);
nand U7942 (N_7942,N_7889,N_7884);
nor U7943 (N_7943,N_7851,N_7834);
and U7944 (N_7944,N_7860,N_7864);
or U7945 (N_7945,N_7852,N_7883);
and U7946 (N_7946,N_7831,N_7821);
or U7947 (N_7947,N_7818,N_7892);
nor U7948 (N_7948,N_7881,N_7863);
or U7949 (N_7949,N_7807,N_7876);
or U7950 (N_7950,N_7891,N_7884);
nand U7951 (N_7951,N_7877,N_7805);
and U7952 (N_7952,N_7810,N_7827);
xor U7953 (N_7953,N_7825,N_7858);
nand U7954 (N_7954,N_7896,N_7892);
or U7955 (N_7955,N_7850,N_7861);
or U7956 (N_7956,N_7880,N_7828);
nand U7957 (N_7957,N_7823,N_7856);
nor U7958 (N_7958,N_7880,N_7832);
xnor U7959 (N_7959,N_7818,N_7882);
and U7960 (N_7960,N_7848,N_7803);
nand U7961 (N_7961,N_7803,N_7869);
nand U7962 (N_7962,N_7844,N_7847);
or U7963 (N_7963,N_7800,N_7810);
nor U7964 (N_7964,N_7816,N_7896);
and U7965 (N_7965,N_7865,N_7811);
nor U7966 (N_7966,N_7816,N_7863);
or U7967 (N_7967,N_7886,N_7891);
and U7968 (N_7968,N_7831,N_7826);
or U7969 (N_7969,N_7838,N_7826);
nor U7970 (N_7970,N_7894,N_7806);
or U7971 (N_7971,N_7877,N_7898);
or U7972 (N_7972,N_7899,N_7830);
nand U7973 (N_7973,N_7896,N_7854);
and U7974 (N_7974,N_7823,N_7884);
nand U7975 (N_7975,N_7825,N_7887);
and U7976 (N_7976,N_7838,N_7842);
nor U7977 (N_7977,N_7824,N_7893);
or U7978 (N_7978,N_7825,N_7843);
or U7979 (N_7979,N_7838,N_7867);
nand U7980 (N_7980,N_7855,N_7833);
nor U7981 (N_7981,N_7897,N_7851);
or U7982 (N_7982,N_7877,N_7839);
nor U7983 (N_7983,N_7802,N_7846);
nor U7984 (N_7984,N_7824,N_7825);
nor U7985 (N_7985,N_7866,N_7841);
xor U7986 (N_7986,N_7882,N_7832);
nand U7987 (N_7987,N_7811,N_7884);
or U7988 (N_7988,N_7839,N_7832);
nand U7989 (N_7989,N_7862,N_7883);
nand U7990 (N_7990,N_7845,N_7822);
and U7991 (N_7991,N_7877,N_7867);
nor U7992 (N_7992,N_7827,N_7811);
nor U7993 (N_7993,N_7848,N_7812);
nor U7994 (N_7994,N_7889,N_7842);
nor U7995 (N_7995,N_7811,N_7871);
or U7996 (N_7996,N_7892,N_7878);
nand U7997 (N_7997,N_7822,N_7878);
and U7998 (N_7998,N_7858,N_7872);
nor U7999 (N_7999,N_7880,N_7809);
and U8000 (N_8000,N_7946,N_7936);
nand U8001 (N_8001,N_7930,N_7955);
and U8002 (N_8002,N_7918,N_7904);
nand U8003 (N_8003,N_7971,N_7957);
nor U8004 (N_8004,N_7973,N_7937);
nor U8005 (N_8005,N_7966,N_7920);
or U8006 (N_8006,N_7921,N_7939);
nor U8007 (N_8007,N_7919,N_7963);
and U8008 (N_8008,N_7941,N_7956);
or U8009 (N_8009,N_7984,N_7903);
nand U8010 (N_8010,N_7913,N_7901);
nor U8011 (N_8011,N_7922,N_7931);
and U8012 (N_8012,N_7934,N_7987);
nor U8013 (N_8013,N_7951,N_7905);
nor U8014 (N_8014,N_7983,N_7916);
xnor U8015 (N_8015,N_7938,N_7978);
nor U8016 (N_8016,N_7962,N_7967);
nor U8017 (N_8017,N_7960,N_7965);
nor U8018 (N_8018,N_7968,N_7950);
nor U8019 (N_8019,N_7908,N_7900);
nor U8020 (N_8020,N_7902,N_7952);
nand U8021 (N_8021,N_7997,N_7932);
nor U8022 (N_8022,N_7995,N_7912);
and U8023 (N_8023,N_7990,N_7907);
nor U8024 (N_8024,N_7928,N_7993);
nand U8025 (N_8025,N_7974,N_7989);
or U8026 (N_8026,N_7906,N_7954);
nor U8027 (N_8027,N_7992,N_7927);
nand U8028 (N_8028,N_7925,N_7953);
nor U8029 (N_8029,N_7948,N_7999);
and U8030 (N_8030,N_7911,N_7979);
nor U8031 (N_8031,N_7985,N_7942);
and U8032 (N_8032,N_7970,N_7976);
and U8033 (N_8033,N_7945,N_7910);
and U8034 (N_8034,N_7975,N_7929);
xnor U8035 (N_8035,N_7909,N_7981);
nor U8036 (N_8036,N_7940,N_7972);
nand U8037 (N_8037,N_7998,N_7947);
or U8038 (N_8038,N_7924,N_7926);
and U8039 (N_8039,N_7944,N_7977);
and U8040 (N_8040,N_7923,N_7986);
nand U8041 (N_8041,N_7958,N_7980);
or U8042 (N_8042,N_7935,N_7988);
nand U8043 (N_8043,N_7914,N_7959);
nand U8044 (N_8044,N_7994,N_7949);
or U8045 (N_8045,N_7964,N_7915);
nand U8046 (N_8046,N_7991,N_7982);
and U8047 (N_8047,N_7933,N_7917);
nor U8048 (N_8048,N_7996,N_7961);
nor U8049 (N_8049,N_7943,N_7969);
or U8050 (N_8050,N_7922,N_7978);
or U8051 (N_8051,N_7994,N_7967);
and U8052 (N_8052,N_7959,N_7909);
or U8053 (N_8053,N_7900,N_7910);
and U8054 (N_8054,N_7995,N_7904);
nand U8055 (N_8055,N_7963,N_7965);
or U8056 (N_8056,N_7907,N_7947);
nand U8057 (N_8057,N_7924,N_7949);
or U8058 (N_8058,N_7925,N_7903);
xnor U8059 (N_8059,N_7981,N_7957);
and U8060 (N_8060,N_7969,N_7904);
and U8061 (N_8061,N_7940,N_7957);
and U8062 (N_8062,N_7996,N_7997);
nor U8063 (N_8063,N_7973,N_7904);
nor U8064 (N_8064,N_7918,N_7925);
or U8065 (N_8065,N_7977,N_7954);
and U8066 (N_8066,N_7928,N_7916);
and U8067 (N_8067,N_7933,N_7991);
or U8068 (N_8068,N_7983,N_7951);
xor U8069 (N_8069,N_7996,N_7990);
xnor U8070 (N_8070,N_7981,N_7949);
or U8071 (N_8071,N_7995,N_7911);
nand U8072 (N_8072,N_7975,N_7912);
nand U8073 (N_8073,N_7903,N_7999);
and U8074 (N_8074,N_7989,N_7982);
xnor U8075 (N_8075,N_7906,N_7966);
nand U8076 (N_8076,N_7929,N_7950);
or U8077 (N_8077,N_7904,N_7934);
nand U8078 (N_8078,N_7964,N_7981);
and U8079 (N_8079,N_7933,N_7964);
nor U8080 (N_8080,N_7912,N_7900);
or U8081 (N_8081,N_7936,N_7969);
nor U8082 (N_8082,N_7938,N_7962);
nor U8083 (N_8083,N_7972,N_7964);
nor U8084 (N_8084,N_7996,N_7982);
nand U8085 (N_8085,N_7993,N_7978);
or U8086 (N_8086,N_7902,N_7914);
or U8087 (N_8087,N_7965,N_7955);
nor U8088 (N_8088,N_7919,N_7959);
nor U8089 (N_8089,N_7975,N_7963);
nor U8090 (N_8090,N_7922,N_7912);
nor U8091 (N_8091,N_7962,N_7915);
nor U8092 (N_8092,N_7957,N_7901);
or U8093 (N_8093,N_7928,N_7962);
nand U8094 (N_8094,N_7984,N_7999);
nand U8095 (N_8095,N_7980,N_7941);
nand U8096 (N_8096,N_7969,N_7968);
nand U8097 (N_8097,N_7999,N_7902);
nor U8098 (N_8098,N_7927,N_7973);
nand U8099 (N_8099,N_7913,N_7904);
or U8100 (N_8100,N_8006,N_8050);
and U8101 (N_8101,N_8054,N_8053);
xor U8102 (N_8102,N_8091,N_8014);
nand U8103 (N_8103,N_8048,N_8060);
and U8104 (N_8104,N_8075,N_8007);
nand U8105 (N_8105,N_8079,N_8099);
nand U8106 (N_8106,N_8022,N_8017);
and U8107 (N_8107,N_8094,N_8031);
or U8108 (N_8108,N_8095,N_8015);
and U8109 (N_8109,N_8071,N_8039);
nand U8110 (N_8110,N_8051,N_8086);
and U8111 (N_8111,N_8081,N_8063);
and U8112 (N_8112,N_8011,N_8044);
xor U8113 (N_8113,N_8073,N_8027);
or U8114 (N_8114,N_8058,N_8056);
or U8115 (N_8115,N_8018,N_8012);
or U8116 (N_8116,N_8078,N_8000);
or U8117 (N_8117,N_8047,N_8055);
nand U8118 (N_8118,N_8089,N_8023);
nor U8119 (N_8119,N_8008,N_8046);
nor U8120 (N_8120,N_8025,N_8062);
nand U8121 (N_8121,N_8059,N_8001);
nor U8122 (N_8122,N_8090,N_8085);
nand U8123 (N_8123,N_8020,N_8038);
nor U8124 (N_8124,N_8013,N_8002);
nor U8125 (N_8125,N_8074,N_8024);
and U8126 (N_8126,N_8035,N_8087);
nor U8127 (N_8127,N_8066,N_8049);
and U8128 (N_8128,N_8040,N_8029);
nor U8129 (N_8129,N_8057,N_8033);
and U8130 (N_8130,N_8093,N_8065);
nor U8131 (N_8131,N_8036,N_8009);
nand U8132 (N_8132,N_8021,N_8084);
xor U8133 (N_8133,N_8043,N_8032);
or U8134 (N_8134,N_8097,N_8037);
nand U8135 (N_8135,N_8028,N_8082);
or U8136 (N_8136,N_8083,N_8070);
nor U8137 (N_8137,N_8030,N_8077);
nand U8138 (N_8138,N_8096,N_8019);
nor U8139 (N_8139,N_8061,N_8016);
or U8140 (N_8140,N_8010,N_8067);
or U8141 (N_8141,N_8005,N_8041);
nor U8142 (N_8142,N_8080,N_8088);
nor U8143 (N_8143,N_8003,N_8098);
nand U8144 (N_8144,N_8042,N_8076);
and U8145 (N_8145,N_8069,N_8045);
or U8146 (N_8146,N_8052,N_8064);
or U8147 (N_8147,N_8092,N_8072);
xnor U8148 (N_8148,N_8068,N_8034);
nor U8149 (N_8149,N_8004,N_8026);
nor U8150 (N_8150,N_8066,N_8090);
or U8151 (N_8151,N_8067,N_8094);
or U8152 (N_8152,N_8032,N_8080);
nor U8153 (N_8153,N_8084,N_8088);
and U8154 (N_8154,N_8087,N_8056);
and U8155 (N_8155,N_8064,N_8025);
or U8156 (N_8156,N_8051,N_8061);
nand U8157 (N_8157,N_8044,N_8081);
nor U8158 (N_8158,N_8045,N_8080);
and U8159 (N_8159,N_8029,N_8064);
or U8160 (N_8160,N_8037,N_8009);
and U8161 (N_8161,N_8052,N_8083);
or U8162 (N_8162,N_8071,N_8064);
or U8163 (N_8163,N_8001,N_8051);
nand U8164 (N_8164,N_8099,N_8028);
or U8165 (N_8165,N_8007,N_8082);
nand U8166 (N_8166,N_8037,N_8010);
and U8167 (N_8167,N_8048,N_8029);
nand U8168 (N_8168,N_8049,N_8086);
and U8169 (N_8169,N_8085,N_8091);
nor U8170 (N_8170,N_8054,N_8057);
and U8171 (N_8171,N_8020,N_8006);
or U8172 (N_8172,N_8085,N_8017);
nor U8173 (N_8173,N_8066,N_8016);
nand U8174 (N_8174,N_8042,N_8008);
nand U8175 (N_8175,N_8001,N_8079);
and U8176 (N_8176,N_8057,N_8000);
nand U8177 (N_8177,N_8086,N_8034);
nand U8178 (N_8178,N_8036,N_8022);
nor U8179 (N_8179,N_8094,N_8017);
and U8180 (N_8180,N_8050,N_8098);
nand U8181 (N_8181,N_8098,N_8088);
nor U8182 (N_8182,N_8022,N_8065);
and U8183 (N_8183,N_8086,N_8000);
nor U8184 (N_8184,N_8024,N_8087);
nand U8185 (N_8185,N_8016,N_8000);
nand U8186 (N_8186,N_8093,N_8083);
nand U8187 (N_8187,N_8006,N_8035);
nand U8188 (N_8188,N_8085,N_8093);
xnor U8189 (N_8189,N_8015,N_8051);
and U8190 (N_8190,N_8009,N_8043);
or U8191 (N_8191,N_8054,N_8070);
nor U8192 (N_8192,N_8068,N_8083);
nand U8193 (N_8193,N_8013,N_8083);
xor U8194 (N_8194,N_8099,N_8073);
nand U8195 (N_8195,N_8031,N_8058);
xnor U8196 (N_8196,N_8042,N_8051);
and U8197 (N_8197,N_8092,N_8074);
nor U8198 (N_8198,N_8049,N_8025);
or U8199 (N_8199,N_8039,N_8078);
nor U8200 (N_8200,N_8102,N_8182);
nand U8201 (N_8201,N_8197,N_8198);
nor U8202 (N_8202,N_8115,N_8137);
nand U8203 (N_8203,N_8172,N_8188);
and U8204 (N_8204,N_8150,N_8189);
nor U8205 (N_8205,N_8116,N_8144);
nand U8206 (N_8206,N_8108,N_8173);
or U8207 (N_8207,N_8103,N_8161);
and U8208 (N_8208,N_8190,N_8129);
or U8209 (N_8209,N_8152,N_8126);
nand U8210 (N_8210,N_8151,N_8119);
nor U8211 (N_8211,N_8113,N_8123);
and U8212 (N_8212,N_8196,N_8183);
or U8213 (N_8213,N_8146,N_8185);
nand U8214 (N_8214,N_8174,N_8194);
or U8215 (N_8215,N_8132,N_8180);
nor U8216 (N_8216,N_8159,N_8178);
nor U8217 (N_8217,N_8112,N_8100);
nand U8218 (N_8218,N_8193,N_8140);
and U8219 (N_8219,N_8158,N_8156);
and U8220 (N_8220,N_8135,N_8128);
nand U8221 (N_8221,N_8195,N_8121);
nor U8222 (N_8222,N_8153,N_8114);
and U8223 (N_8223,N_8184,N_8162);
and U8224 (N_8224,N_8145,N_8105);
or U8225 (N_8225,N_8175,N_8167);
nor U8226 (N_8226,N_8170,N_8139);
nand U8227 (N_8227,N_8155,N_8147);
nor U8228 (N_8228,N_8192,N_8109);
nor U8229 (N_8229,N_8107,N_8133);
nand U8230 (N_8230,N_8124,N_8160);
and U8231 (N_8231,N_8166,N_8149);
or U8232 (N_8232,N_8143,N_8177);
nand U8233 (N_8233,N_8179,N_8110);
nand U8234 (N_8234,N_8169,N_8157);
and U8235 (N_8235,N_8142,N_8136);
and U8236 (N_8236,N_8176,N_8187);
nor U8237 (N_8237,N_8181,N_8127);
nor U8238 (N_8238,N_8141,N_8134);
and U8239 (N_8239,N_8101,N_8154);
or U8240 (N_8240,N_8163,N_8104);
nor U8241 (N_8241,N_8106,N_8131);
or U8242 (N_8242,N_8125,N_8171);
nand U8243 (N_8243,N_8168,N_8148);
and U8244 (N_8244,N_8130,N_8164);
nor U8245 (N_8245,N_8117,N_8186);
and U8246 (N_8246,N_8165,N_8111);
nor U8247 (N_8247,N_8199,N_8191);
nand U8248 (N_8248,N_8138,N_8118);
and U8249 (N_8249,N_8120,N_8122);
and U8250 (N_8250,N_8198,N_8166);
nand U8251 (N_8251,N_8180,N_8116);
nor U8252 (N_8252,N_8197,N_8156);
nand U8253 (N_8253,N_8135,N_8151);
nand U8254 (N_8254,N_8158,N_8184);
nand U8255 (N_8255,N_8150,N_8113);
and U8256 (N_8256,N_8172,N_8192);
nand U8257 (N_8257,N_8131,N_8195);
nor U8258 (N_8258,N_8144,N_8131);
or U8259 (N_8259,N_8133,N_8189);
nor U8260 (N_8260,N_8130,N_8122);
or U8261 (N_8261,N_8108,N_8169);
or U8262 (N_8262,N_8171,N_8138);
and U8263 (N_8263,N_8122,N_8151);
nand U8264 (N_8264,N_8132,N_8183);
and U8265 (N_8265,N_8137,N_8116);
or U8266 (N_8266,N_8123,N_8159);
nand U8267 (N_8267,N_8112,N_8147);
xnor U8268 (N_8268,N_8141,N_8180);
nand U8269 (N_8269,N_8106,N_8100);
and U8270 (N_8270,N_8161,N_8160);
and U8271 (N_8271,N_8160,N_8119);
and U8272 (N_8272,N_8161,N_8114);
or U8273 (N_8273,N_8118,N_8148);
nand U8274 (N_8274,N_8147,N_8143);
and U8275 (N_8275,N_8123,N_8126);
and U8276 (N_8276,N_8115,N_8187);
xnor U8277 (N_8277,N_8168,N_8170);
nor U8278 (N_8278,N_8183,N_8124);
or U8279 (N_8279,N_8174,N_8169);
and U8280 (N_8280,N_8139,N_8145);
and U8281 (N_8281,N_8154,N_8169);
nor U8282 (N_8282,N_8134,N_8145);
and U8283 (N_8283,N_8182,N_8125);
nand U8284 (N_8284,N_8142,N_8197);
nand U8285 (N_8285,N_8192,N_8151);
and U8286 (N_8286,N_8136,N_8156);
xor U8287 (N_8287,N_8104,N_8171);
or U8288 (N_8288,N_8164,N_8199);
nor U8289 (N_8289,N_8148,N_8117);
or U8290 (N_8290,N_8181,N_8152);
and U8291 (N_8291,N_8188,N_8154);
nor U8292 (N_8292,N_8106,N_8158);
nor U8293 (N_8293,N_8134,N_8173);
or U8294 (N_8294,N_8156,N_8184);
nor U8295 (N_8295,N_8110,N_8151);
nand U8296 (N_8296,N_8192,N_8148);
or U8297 (N_8297,N_8177,N_8184);
or U8298 (N_8298,N_8168,N_8179);
nand U8299 (N_8299,N_8160,N_8120);
or U8300 (N_8300,N_8233,N_8220);
nor U8301 (N_8301,N_8250,N_8201);
nor U8302 (N_8302,N_8251,N_8262);
and U8303 (N_8303,N_8298,N_8240);
nand U8304 (N_8304,N_8291,N_8252);
or U8305 (N_8305,N_8232,N_8259);
nand U8306 (N_8306,N_8289,N_8255);
and U8307 (N_8307,N_8280,N_8212);
and U8308 (N_8308,N_8202,N_8238);
and U8309 (N_8309,N_8268,N_8285);
nor U8310 (N_8310,N_8237,N_8260);
nand U8311 (N_8311,N_8234,N_8226);
nand U8312 (N_8312,N_8235,N_8282);
nor U8313 (N_8313,N_8200,N_8261);
and U8314 (N_8314,N_8204,N_8276);
and U8315 (N_8315,N_8203,N_8244);
and U8316 (N_8316,N_8242,N_8297);
xor U8317 (N_8317,N_8211,N_8265);
nand U8318 (N_8318,N_8236,N_8224);
nor U8319 (N_8319,N_8214,N_8273);
nor U8320 (N_8320,N_8213,N_8288);
or U8321 (N_8321,N_8248,N_8281);
nor U8322 (N_8322,N_8221,N_8243);
or U8323 (N_8323,N_8253,N_8293);
nor U8324 (N_8324,N_8267,N_8287);
or U8325 (N_8325,N_8241,N_8256);
nor U8326 (N_8326,N_8205,N_8222);
and U8327 (N_8327,N_8299,N_8208);
nor U8328 (N_8328,N_8275,N_8294);
nand U8329 (N_8329,N_8278,N_8270);
nand U8330 (N_8330,N_8239,N_8295);
nand U8331 (N_8331,N_8210,N_8264);
nor U8332 (N_8332,N_8272,N_8247);
and U8333 (N_8333,N_8216,N_8209);
or U8334 (N_8334,N_8249,N_8271);
or U8335 (N_8335,N_8228,N_8269);
nor U8336 (N_8336,N_8274,N_8296);
nand U8337 (N_8337,N_8215,N_8206);
or U8338 (N_8338,N_8219,N_8277);
nor U8339 (N_8339,N_8217,N_8246);
and U8340 (N_8340,N_8257,N_8283);
or U8341 (N_8341,N_8225,N_8279);
nor U8342 (N_8342,N_8229,N_8266);
and U8343 (N_8343,N_8207,N_8223);
nand U8344 (N_8344,N_8245,N_8292);
nand U8345 (N_8345,N_8218,N_8254);
nor U8346 (N_8346,N_8284,N_8231);
nand U8347 (N_8347,N_8230,N_8263);
or U8348 (N_8348,N_8286,N_8227);
or U8349 (N_8349,N_8290,N_8258);
and U8350 (N_8350,N_8239,N_8283);
or U8351 (N_8351,N_8284,N_8288);
nor U8352 (N_8352,N_8257,N_8238);
and U8353 (N_8353,N_8201,N_8205);
nand U8354 (N_8354,N_8269,N_8299);
and U8355 (N_8355,N_8249,N_8289);
and U8356 (N_8356,N_8213,N_8286);
nor U8357 (N_8357,N_8282,N_8251);
and U8358 (N_8358,N_8221,N_8209);
and U8359 (N_8359,N_8254,N_8200);
and U8360 (N_8360,N_8295,N_8222);
and U8361 (N_8361,N_8267,N_8262);
nor U8362 (N_8362,N_8269,N_8215);
nor U8363 (N_8363,N_8271,N_8222);
nand U8364 (N_8364,N_8218,N_8251);
or U8365 (N_8365,N_8283,N_8282);
and U8366 (N_8366,N_8215,N_8267);
nand U8367 (N_8367,N_8268,N_8235);
and U8368 (N_8368,N_8264,N_8275);
or U8369 (N_8369,N_8230,N_8214);
nor U8370 (N_8370,N_8212,N_8259);
and U8371 (N_8371,N_8229,N_8255);
nand U8372 (N_8372,N_8221,N_8286);
or U8373 (N_8373,N_8275,N_8299);
or U8374 (N_8374,N_8204,N_8278);
nand U8375 (N_8375,N_8215,N_8285);
or U8376 (N_8376,N_8271,N_8245);
xor U8377 (N_8377,N_8241,N_8265);
or U8378 (N_8378,N_8213,N_8269);
nor U8379 (N_8379,N_8217,N_8277);
nand U8380 (N_8380,N_8287,N_8296);
nand U8381 (N_8381,N_8200,N_8292);
nand U8382 (N_8382,N_8234,N_8241);
and U8383 (N_8383,N_8247,N_8261);
nor U8384 (N_8384,N_8209,N_8257);
nor U8385 (N_8385,N_8249,N_8226);
nand U8386 (N_8386,N_8236,N_8245);
and U8387 (N_8387,N_8221,N_8288);
and U8388 (N_8388,N_8293,N_8249);
and U8389 (N_8389,N_8202,N_8212);
nand U8390 (N_8390,N_8293,N_8212);
or U8391 (N_8391,N_8277,N_8284);
or U8392 (N_8392,N_8270,N_8219);
and U8393 (N_8393,N_8200,N_8251);
nor U8394 (N_8394,N_8256,N_8217);
or U8395 (N_8395,N_8267,N_8224);
and U8396 (N_8396,N_8206,N_8266);
or U8397 (N_8397,N_8228,N_8223);
nand U8398 (N_8398,N_8218,N_8210);
nand U8399 (N_8399,N_8221,N_8235);
and U8400 (N_8400,N_8371,N_8373);
or U8401 (N_8401,N_8332,N_8361);
or U8402 (N_8402,N_8313,N_8328);
or U8403 (N_8403,N_8321,N_8379);
or U8404 (N_8404,N_8308,N_8309);
or U8405 (N_8405,N_8383,N_8364);
nand U8406 (N_8406,N_8329,N_8344);
nand U8407 (N_8407,N_8347,N_8395);
nor U8408 (N_8408,N_8314,N_8399);
and U8409 (N_8409,N_8331,N_8349);
and U8410 (N_8410,N_8348,N_8394);
nand U8411 (N_8411,N_8334,N_8336);
and U8412 (N_8412,N_8388,N_8306);
nor U8413 (N_8413,N_8350,N_8335);
or U8414 (N_8414,N_8391,N_8300);
nor U8415 (N_8415,N_8343,N_8324);
nand U8416 (N_8416,N_8323,N_8318);
nand U8417 (N_8417,N_8340,N_8359);
and U8418 (N_8418,N_8365,N_8390);
nand U8419 (N_8419,N_8385,N_8301);
and U8420 (N_8420,N_8376,N_8375);
nand U8421 (N_8421,N_8333,N_8315);
nor U8422 (N_8422,N_8320,N_8302);
or U8423 (N_8423,N_8304,N_8369);
nor U8424 (N_8424,N_8377,N_8393);
nor U8425 (N_8425,N_8342,N_8338);
nand U8426 (N_8426,N_8389,N_8322);
nand U8427 (N_8427,N_8345,N_8356);
nor U8428 (N_8428,N_8354,N_8398);
and U8429 (N_8429,N_8353,N_8382);
and U8430 (N_8430,N_8346,N_8310);
or U8431 (N_8431,N_8330,N_8358);
or U8432 (N_8432,N_8351,N_8378);
or U8433 (N_8433,N_8363,N_8339);
and U8434 (N_8434,N_8360,N_8386);
and U8435 (N_8435,N_8312,N_8355);
and U8436 (N_8436,N_8311,N_8368);
or U8437 (N_8437,N_8325,N_8387);
nand U8438 (N_8438,N_8327,N_8397);
or U8439 (N_8439,N_8357,N_8366);
nor U8440 (N_8440,N_8319,N_8305);
nor U8441 (N_8441,N_8307,N_8392);
nand U8442 (N_8442,N_8380,N_8384);
nand U8443 (N_8443,N_8374,N_8337);
nand U8444 (N_8444,N_8367,N_8303);
xor U8445 (N_8445,N_8341,N_8326);
nor U8446 (N_8446,N_8352,N_8316);
nand U8447 (N_8447,N_8381,N_8317);
or U8448 (N_8448,N_8396,N_8372);
nand U8449 (N_8449,N_8370,N_8362);
or U8450 (N_8450,N_8366,N_8313);
or U8451 (N_8451,N_8318,N_8374);
or U8452 (N_8452,N_8354,N_8325);
and U8453 (N_8453,N_8383,N_8363);
or U8454 (N_8454,N_8370,N_8332);
or U8455 (N_8455,N_8360,N_8374);
nand U8456 (N_8456,N_8303,N_8375);
or U8457 (N_8457,N_8342,N_8328);
nand U8458 (N_8458,N_8315,N_8363);
or U8459 (N_8459,N_8311,N_8317);
or U8460 (N_8460,N_8363,N_8302);
and U8461 (N_8461,N_8315,N_8323);
nor U8462 (N_8462,N_8378,N_8350);
and U8463 (N_8463,N_8352,N_8375);
nor U8464 (N_8464,N_8387,N_8328);
and U8465 (N_8465,N_8300,N_8369);
nand U8466 (N_8466,N_8353,N_8396);
and U8467 (N_8467,N_8347,N_8362);
nand U8468 (N_8468,N_8384,N_8344);
nor U8469 (N_8469,N_8322,N_8343);
nor U8470 (N_8470,N_8301,N_8395);
or U8471 (N_8471,N_8366,N_8354);
or U8472 (N_8472,N_8351,N_8360);
or U8473 (N_8473,N_8354,N_8397);
or U8474 (N_8474,N_8335,N_8353);
and U8475 (N_8475,N_8311,N_8361);
and U8476 (N_8476,N_8382,N_8343);
nor U8477 (N_8477,N_8315,N_8314);
and U8478 (N_8478,N_8384,N_8345);
or U8479 (N_8479,N_8359,N_8392);
or U8480 (N_8480,N_8378,N_8314);
nor U8481 (N_8481,N_8389,N_8383);
xnor U8482 (N_8482,N_8322,N_8307);
nor U8483 (N_8483,N_8339,N_8357);
or U8484 (N_8484,N_8376,N_8393);
nor U8485 (N_8485,N_8312,N_8327);
nor U8486 (N_8486,N_8346,N_8308);
and U8487 (N_8487,N_8332,N_8302);
or U8488 (N_8488,N_8334,N_8308);
or U8489 (N_8489,N_8350,N_8381);
or U8490 (N_8490,N_8341,N_8380);
nand U8491 (N_8491,N_8318,N_8370);
nand U8492 (N_8492,N_8388,N_8356);
or U8493 (N_8493,N_8368,N_8378);
and U8494 (N_8494,N_8373,N_8382);
nor U8495 (N_8495,N_8329,N_8366);
or U8496 (N_8496,N_8307,N_8359);
nand U8497 (N_8497,N_8360,N_8362);
or U8498 (N_8498,N_8347,N_8386);
nor U8499 (N_8499,N_8340,N_8380);
nand U8500 (N_8500,N_8460,N_8477);
xor U8501 (N_8501,N_8406,N_8426);
nor U8502 (N_8502,N_8470,N_8433);
and U8503 (N_8503,N_8497,N_8411);
or U8504 (N_8504,N_8483,N_8427);
nand U8505 (N_8505,N_8403,N_8445);
nor U8506 (N_8506,N_8441,N_8456);
or U8507 (N_8507,N_8462,N_8416);
nor U8508 (N_8508,N_8401,N_8437);
or U8509 (N_8509,N_8418,N_8404);
nand U8510 (N_8510,N_8481,N_8461);
nand U8511 (N_8511,N_8423,N_8405);
or U8512 (N_8512,N_8431,N_8436);
nand U8513 (N_8513,N_8402,N_8415);
nand U8514 (N_8514,N_8451,N_8409);
or U8515 (N_8515,N_8408,N_8417);
and U8516 (N_8516,N_8459,N_8484);
and U8517 (N_8517,N_8474,N_8468);
nand U8518 (N_8518,N_8465,N_8458);
or U8519 (N_8519,N_8488,N_8414);
and U8520 (N_8520,N_8450,N_8442);
and U8521 (N_8521,N_8466,N_8457);
and U8522 (N_8522,N_8498,N_8439);
nor U8523 (N_8523,N_8444,N_8464);
or U8524 (N_8524,N_8440,N_8479);
nand U8525 (N_8525,N_8422,N_8434);
nand U8526 (N_8526,N_8428,N_8487);
nor U8527 (N_8527,N_8478,N_8432);
nand U8528 (N_8528,N_8475,N_8429);
nand U8529 (N_8529,N_8467,N_8495);
or U8530 (N_8530,N_8496,N_8463);
or U8531 (N_8531,N_8419,N_8447);
nor U8532 (N_8532,N_8452,N_8494);
nor U8533 (N_8533,N_8471,N_8443);
and U8534 (N_8534,N_8499,N_8430);
nand U8535 (N_8535,N_8472,N_8424);
nand U8536 (N_8536,N_8453,N_8473);
nand U8537 (N_8537,N_8493,N_8448);
or U8538 (N_8538,N_8438,N_8425);
nor U8539 (N_8539,N_8455,N_8485);
or U8540 (N_8540,N_8413,N_8476);
or U8541 (N_8541,N_8420,N_8400);
or U8542 (N_8542,N_8491,N_8482);
nor U8543 (N_8543,N_8490,N_8421);
or U8544 (N_8544,N_8410,N_8486);
nand U8545 (N_8545,N_8454,N_8449);
xnor U8546 (N_8546,N_8435,N_8492);
nor U8547 (N_8547,N_8407,N_8480);
and U8548 (N_8548,N_8446,N_8469);
and U8549 (N_8549,N_8489,N_8412);
or U8550 (N_8550,N_8433,N_8406);
nor U8551 (N_8551,N_8469,N_8484);
nand U8552 (N_8552,N_8490,N_8433);
xor U8553 (N_8553,N_8418,N_8434);
and U8554 (N_8554,N_8486,N_8432);
and U8555 (N_8555,N_8445,N_8480);
nand U8556 (N_8556,N_8463,N_8440);
and U8557 (N_8557,N_8487,N_8485);
and U8558 (N_8558,N_8478,N_8433);
nor U8559 (N_8559,N_8407,N_8451);
and U8560 (N_8560,N_8462,N_8465);
nor U8561 (N_8561,N_8400,N_8475);
nor U8562 (N_8562,N_8407,N_8453);
nand U8563 (N_8563,N_8486,N_8425);
and U8564 (N_8564,N_8441,N_8481);
nor U8565 (N_8565,N_8492,N_8494);
nand U8566 (N_8566,N_8494,N_8476);
nor U8567 (N_8567,N_8411,N_8436);
nor U8568 (N_8568,N_8447,N_8401);
and U8569 (N_8569,N_8435,N_8451);
or U8570 (N_8570,N_8404,N_8417);
and U8571 (N_8571,N_8415,N_8447);
and U8572 (N_8572,N_8483,N_8448);
nor U8573 (N_8573,N_8409,N_8464);
and U8574 (N_8574,N_8486,N_8478);
nand U8575 (N_8575,N_8414,N_8450);
nor U8576 (N_8576,N_8494,N_8442);
nand U8577 (N_8577,N_8488,N_8420);
and U8578 (N_8578,N_8497,N_8458);
nand U8579 (N_8579,N_8497,N_8481);
or U8580 (N_8580,N_8441,N_8465);
nand U8581 (N_8581,N_8404,N_8492);
and U8582 (N_8582,N_8457,N_8414);
nor U8583 (N_8583,N_8423,N_8467);
nor U8584 (N_8584,N_8421,N_8422);
or U8585 (N_8585,N_8478,N_8460);
and U8586 (N_8586,N_8435,N_8476);
and U8587 (N_8587,N_8491,N_8455);
and U8588 (N_8588,N_8445,N_8460);
nor U8589 (N_8589,N_8472,N_8459);
and U8590 (N_8590,N_8459,N_8461);
and U8591 (N_8591,N_8437,N_8469);
nand U8592 (N_8592,N_8460,N_8459);
nor U8593 (N_8593,N_8438,N_8461);
or U8594 (N_8594,N_8461,N_8419);
nand U8595 (N_8595,N_8493,N_8473);
nor U8596 (N_8596,N_8411,N_8402);
nand U8597 (N_8597,N_8412,N_8446);
or U8598 (N_8598,N_8430,N_8492);
and U8599 (N_8599,N_8420,N_8499);
or U8600 (N_8600,N_8523,N_8552);
nand U8601 (N_8601,N_8588,N_8576);
nor U8602 (N_8602,N_8575,N_8502);
or U8603 (N_8603,N_8560,N_8574);
and U8604 (N_8604,N_8536,N_8571);
or U8605 (N_8605,N_8572,N_8532);
nand U8606 (N_8606,N_8547,N_8587);
nor U8607 (N_8607,N_8581,N_8548);
xor U8608 (N_8608,N_8521,N_8512);
nor U8609 (N_8609,N_8522,N_8545);
nor U8610 (N_8610,N_8517,N_8584);
nand U8611 (N_8611,N_8557,N_8566);
or U8612 (N_8612,N_8562,N_8596);
nand U8613 (N_8613,N_8540,N_8589);
nor U8614 (N_8614,N_8582,N_8568);
nand U8615 (N_8615,N_8509,N_8591);
and U8616 (N_8616,N_8515,N_8529);
and U8617 (N_8617,N_8577,N_8599);
nand U8618 (N_8618,N_8555,N_8506);
nand U8619 (N_8619,N_8503,N_8593);
nand U8620 (N_8620,N_8508,N_8530);
nor U8621 (N_8621,N_8553,N_8550);
and U8622 (N_8622,N_8501,N_8546);
nor U8623 (N_8623,N_8544,N_8510);
or U8624 (N_8624,N_8592,N_8537);
and U8625 (N_8625,N_8585,N_8514);
and U8626 (N_8626,N_8569,N_8518);
nor U8627 (N_8627,N_8541,N_8583);
or U8628 (N_8628,N_8570,N_8563);
or U8629 (N_8629,N_8543,N_8561);
nand U8630 (N_8630,N_8519,N_8535);
nor U8631 (N_8631,N_8520,N_8567);
or U8632 (N_8632,N_8526,N_8542);
nand U8633 (N_8633,N_8500,N_8579);
or U8634 (N_8634,N_8565,N_8549);
nor U8635 (N_8635,N_8533,N_8580);
or U8636 (N_8636,N_8558,N_8554);
and U8637 (N_8637,N_8597,N_8516);
and U8638 (N_8638,N_8595,N_8539);
or U8639 (N_8639,N_8513,N_8511);
nand U8640 (N_8640,N_8505,N_8504);
or U8641 (N_8641,N_8525,N_8556);
nor U8642 (N_8642,N_8551,N_8598);
nand U8643 (N_8643,N_8531,N_8586);
nor U8644 (N_8644,N_8538,N_8534);
nor U8645 (N_8645,N_8594,N_8524);
nor U8646 (N_8646,N_8564,N_8528);
or U8647 (N_8647,N_8578,N_8559);
and U8648 (N_8648,N_8527,N_8507);
nor U8649 (N_8649,N_8573,N_8590);
and U8650 (N_8650,N_8536,N_8590);
nor U8651 (N_8651,N_8582,N_8588);
nor U8652 (N_8652,N_8568,N_8503);
nand U8653 (N_8653,N_8545,N_8579);
or U8654 (N_8654,N_8550,N_8568);
nand U8655 (N_8655,N_8553,N_8554);
nor U8656 (N_8656,N_8572,N_8561);
nor U8657 (N_8657,N_8592,N_8539);
or U8658 (N_8658,N_8525,N_8506);
xor U8659 (N_8659,N_8532,N_8501);
and U8660 (N_8660,N_8569,N_8515);
and U8661 (N_8661,N_8531,N_8542);
nor U8662 (N_8662,N_8515,N_8554);
or U8663 (N_8663,N_8541,N_8517);
or U8664 (N_8664,N_8575,N_8577);
and U8665 (N_8665,N_8590,N_8543);
nand U8666 (N_8666,N_8531,N_8507);
or U8667 (N_8667,N_8526,N_8556);
nand U8668 (N_8668,N_8533,N_8520);
nor U8669 (N_8669,N_8561,N_8575);
or U8670 (N_8670,N_8539,N_8544);
nand U8671 (N_8671,N_8536,N_8588);
and U8672 (N_8672,N_8567,N_8582);
and U8673 (N_8673,N_8521,N_8532);
and U8674 (N_8674,N_8536,N_8598);
or U8675 (N_8675,N_8515,N_8510);
nand U8676 (N_8676,N_8563,N_8568);
and U8677 (N_8677,N_8520,N_8549);
and U8678 (N_8678,N_8500,N_8529);
nor U8679 (N_8679,N_8521,N_8515);
or U8680 (N_8680,N_8533,N_8585);
and U8681 (N_8681,N_8517,N_8570);
nand U8682 (N_8682,N_8589,N_8590);
and U8683 (N_8683,N_8579,N_8563);
and U8684 (N_8684,N_8527,N_8502);
nand U8685 (N_8685,N_8556,N_8594);
nor U8686 (N_8686,N_8536,N_8526);
or U8687 (N_8687,N_8574,N_8569);
nand U8688 (N_8688,N_8583,N_8569);
or U8689 (N_8689,N_8502,N_8548);
nand U8690 (N_8690,N_8502,N_8513);
nand U8691 (N_8691,N_8590,N_8563);
nand U8692 (N_8692,N_8543,N_8587);
nand U8693 (N_8693,N_8511,N_8554);
nand U8694 (N_8694,N_8598,N_8518);
and U8695 (N_8695,N_8589,N_8581);
nand U8696 (N_8696,N_8513,N_8553);
or U8697 (N_8697,N_8518,N_8590);
or U8698 (N_8698,N_8502,N_8572);
and U8699 (N_8699,N_8586,N_8574);
and U8700 (N_8700,N_8640,N_8679);
nand U8701 (N_8701,N_8685,N_8676);
nand U8702 (N_8702,N_8664,N_8668);
xnor U8703 (N_8703,N_8633,N_8603);
and U8704 (N_8704,N_8608,N_8637);
and U8705 (N_8705,N_8632,N_8652);
and U8706 (N_8706,N_8627,N_8604);
nand U8707 (N_8707,N_8600,N_8617);
and U8708 (N_8708,N_8648,N_8689);
and U8709 (N_8709,N_8602,N_8663);
and U8710 (N_8710,N_8658,N_8670);
nor U8711 (N_8711,N_8634,N_8677);
and U8712 (N_8712,N_8691,N_8612);
or U8713 (N_8713,N_8662,N_8614);
or U8714 (N_8714,N_8696,N_8626);
and U8715 (N_8715,N_8650,N_8654);
or U8716 (N_8716,N_8674,N_8623);
nor U8717 (N_8717,N_8636,N_8688);
or U8718 (N_8718,N_8684,N_8651);
and U8719 (N_8719,N_8615,N_8660);
nand U8720 (N_8720,N_8628,N_8669);
and U8721 (N_8721,N_8610,N_8697);
or U8722 (N_8722,N_8649,N_8659);
nand U8723 (N_8723,N_8695,N_8661);
or U8724 (N_8724,N_8672,N_8682);
nor U8725 (N_8725,N_8618,N_8643);
and U8726 (N_8726,N_8631,N_8646);
nor U8727 (N_8727,N_8690,N_8607);
xor U8728 (N_8728,N_8645,N_8680);
and U8729 (N_8729,N_8655,N_8621);
or U8730 (N_8730,N_8667,N_8629);
and U8731 (N_8731,N_8619,N_8683);
or U8732 (N_8732,N_8635,N_8698);
xor U8733 (N_8733,N_8675,N_8678);
or U8734 (N_8734,N_8606,N_8605);
nand U8735 (N_8735,N_8641,N_8622);
nor U8736 (N_8736,N_8666,N_8671);
or U8737 (N_8737,N_8657,N_8620);
and U8738 (N_8738,N_8609,N_8694);
and U8739 (N_8739,N_8686,N_8625);
or U8740 (N_8740,N_8647,N_8644);
nand U8741 (N_8741,N_8616,N_8611);
nor U8742 (N_8742,N_8681,N_8665);
or U8743 (N_8743,N_8624,N_8613);
or U8744 (N_8744,N_8601,N_8653);
or U8745 (N_8745,N_8639,N_8693);
or U8746 (N_8746,N_8699,N_8687);
and U8747 (N_8747,N_8692,N_8642);
or U8748 (N_8748,N_8630,N_8656);
or U8749 (N_8749,N_8673,N_8638);
nand U8750 (N_8750,N_8657,N_8668);
xor U8751 (N_8751,N_8613,N_8659);
nor U8752 (N_8752,N_8637,N_8653);
and U8753 (N_8753,N_8635,N_8670);
nor U8754 (N_8754,N_8642,N_8675);
or U8755 (N_8755,N_8601,N_8660);
and U8756 (N_8756,N_8653,N_8639);
nand U8757 (N_8757,N_8601,N_8627);
xor U8758 (N_8758,N_8670,N_8639);
and U8759 (N_8759,N_8667,N_8653);
nor U8760 (N_8760,N_8690,N_8638);
nand U8761 (N_8761,N_8620,N_8675);
and U8762 (N_8762,N_8620,N_8690);
or U8763 (N_8763,N_8674,N_8626);
or U8764 (N_8764,N_8626,N_8671);
nand U8765 (N_8765,N_8661,N_8624);
or U8766 (N_8766,N_8695,N_8685);
nor U8767 (N_8767,N_8683,N_8663);
nand U8768 (N_8768,N_8697,N_8602);
nand U8769 (N_8769,N_8646,N_8618);
nor U8770 (N_8770,N_8689,N_8639);
nor U8771 (N_8771,N_8674,N_8617);
or U8772 (N_8772,N_8629,N_8631);
nand U8773 (N_8773,N_8692,N_8639);
or U8774 (N_8774,N_8650,N_8692);
or U8775 (N_8775,N_8695,N_8626);
xnor U8776 (N_8776,N_8646,N_8609);
or U8777 (N_8777,N_8612,N_8610);
nor U8778 (N_8778,N_8682,N_8650);
nor U8779 (N_8779,N_8679,N_8608);
or U8780 (N_8780,N_8618,N_8641);
nand U8781 (N_8781,N_8684,N_8638);
nand U8782 (N_8782,N_8661,N_8606);
nand U8783 (N_8783,N_8675,N_8600);
nor U8784 (N_8784,N_8611,N_8687);
nand U8785 (N_8785,N_8629,N_8647);
xnor U8786 (N_8786,N_8680,N_8687);
nor U8787 (N_8787,N_8601,N_8699);
and U8788 (N_8788,N_8653,N_8675);
and U8789 (N_8789,N_8605,N_8633);
and U8790 (N_8790,N_8665,N_8669);
nor U8791 (N_8791,N_8645,N_8690);
nand U8792 (N_8792,N_8695,N_8694);
and U8793 (N_8793,N_8643,N_8612);
nand U8794 (N_8794,N_8676,N_8681);
nand U8795 (N_8795,N_8635,N_8677);
and U8796 (N_8796,N_8697,N_8672);
or U8797 (N_8797,N_8609,N_8606);
and U8798 (N_8798,N_8661,N_8603);
nand U8799 (N_8799,N_8603,N_8606);
nor U8800 (N_8800,N_8735,N_8737);
and U8801 (N_8801,N_8717,N_8744);
or U8802 (N_8802,N_8753,N_8731);
nor U8803 (N_8803,N_8768,N_8723);
and U8804 (N_8804,N_8728,N_8725);
and U8805 (N_8805,N_8764,N_8772);
or U8806 (N_8806,N_8799,N_8700);
nand U8807 (N_8807,N_8787,N_8721);
xnor U8808 (N_8808,N_8775,N_8751);
nand U8809 (N_8809,N_8734,N_8797);
and U8810 (N_8810,N_8784,N_8759);
and U8811 (N_8811,N_8779,N_8783);
or U8812 (N_8812,N_8796,N_8757);
or U8813 (N_8813,N_8713,N_8777);
nand U8814 (N_8814,N_8712,N_8786);
or U8815 (N_8815,N_8782,N_8724);
or U8816 (N_8816,N_8733,N_8761);
nor U8817 (N_8817,N_8792,N_8708);
or U8818 (N_8818,N_8766,N_8705);
nor U8819 (N_8819,N_8707,N_8739);
nor U8820 (N_8820,N_8736,N_8719);
nand U8821 (N_8821,N_8789,N_8722);
nand U8822 (N_8822,N_8765,N_8755);
nor U8823 (N_8823,N_8740,N_8747);
nand U8824 (N_8824,N_8701,N_8704);
nand U8825 (N_8825,N_8770,N_8750);
or U8826 (N_8826,N_8726,N_8711);
and U8827 (N_8827,N_8718,N_8746);
or U8828 (N_8828,N_8710,N_8732);
nand U8829 (N_8829,N_8715,N_8794);
nand U8830 (N_8830,N_8769,N_8702);
or U8831 (N_8831,N_8742,N_8720);
and U8832 (N_8832,N_8785,N_8743);
and U8833 (N_8833,N_8780,N_8729);
and U8834 (N_8834,N_8788,N_8763);
nand U8835 (N_8835,N_8762,N_8774);
nor U8836 (N_8836,N_8760,N_8773);
nor U8837 (N_8837,N_8714,N_8738);
xnor U8838 (N_8838,N_8752,N_8709);
and U8839 (N_8839,N_8749,N_8754);
and U8840 (N_8840,N_8706,N_8793);
or U8841 (N_8841,N_8727,N_8741);
or U8842 (N_8842,N_8758,N_8776);
nor U8843 (N_8843,N_8730,N_8790);
and U8844 (N_8844,N_8767,N_8703);
or U8845 (N_8845,N_8798,N_8795);
nor U8846 (N_8846,N_8781,N_8771);
nor U8847 (N_8847,N_8756,N_8745);
or U8848 (N_8848,N_8748,N_8791);
nand U8849 (N_8849,N_8778,N_8716);
nand U8850 (N_8850,N_8715,N_8757);
nand U8851 (N_8851,N_8781,N_8718);
or U8852 (N_8852,N_8717,N_8701);
xnor U8853 (N_8853,N_8799,N_8781);
and U8854 (N_8854,N_8703,N_8768);
nor U8855 (N_8855,N_8764,N_8760);
nor U8856 (N_8856,N_8797,N_8744);
or U8857 (N_8857,N_8728,N_8796);
nor U8858 (N_8858,N_8771,N_8734);
or U8859 (N_8859,N_8796,N_8798);
nor U8860 (N_8860,N_8743,N_8798);
or U8861 (N_8861,N_8746,N_8761);
and U8862 (N_8862,N_8725,N_8741);
and U8863 (N_8863,N_8759,N_8704);
nor U8864 (N_8864,N_8779,N_8760);
nor U8865 (N_8865,N_8773,N_8755);
or U8866 (N_8866,N_8799,N_8738);
nor U8867 (N_8867,N_8783,N_8766);
nand U8868 (N_8868,N_8777,N_8766);
nand U8869 (N_8869,N_8784,N_8738);
and U8870 (N_8870,N_8745,N_8717);
nor U8871 (N_8871,N_8770,N_8735);
nor U8872 (N_8872,N_8756,N_8701);
xor U8873 (N_8873,N_8755,N_8718);
or U8874 (N_8874,N_8714,N_8772);
nand U8875 (N_8875,N_8782,N_8728);
nand U8876 (N_8876,N_8787,N_8742);
nand U8877 (N_8877,N_8797,N_8789);
nand U8878 (N_8878,N_8709,N_8723);
and U8879 (N_8879,N_8731,N_8792);
nand U8880 (N_8880,N_8701,N_8793);
or U8881 (N_8881,N_8739,N_8753);
and U8882 (N_8882,N_8737,N_8720);
and U8883 (N_8883,N_8729,N_8720);
and U8884 (N_8884,N_8740,N_8720);
nor U8885 (N_8885,N_8770,N_8768);
nor U8886 (N_8886,N_8701,N_8768);
nor U8887 (N_8887,N_8730,N_8714);
nor U8888 (N_8888,N_8715,N_8746);
nor U8889 (N_8889,N_8720,N_8735);
nor U8890 (N_8890,N_8709,N_8737);
and U8891 (N_8891,N_8723,N_8741);
nor U8892 (N_8892,N_8793,N_8764);
nand U8893 (N_8893,N_8779,N_8764);
xnor U8894 (N_8894,N_8712,N_8771);
nand U8895 (N_8895,N_8777,N_8765);
or U8896 (N_8896,N_8702,N_8779);
nor U8897 (N_8897,N_8768,N_8710);
nor U8898 (N_8898,N_8772,N_8718);
or U8899 (N_8899,N_8703,N_8799);
and U8900 (N_8900,N_8828,N_8882);
nor U8901 (N_8901,N_8879,N_8880);
or U8902 (N_8902,N_8830,N_8859);
and U8903 (N_8903,N_8874,N_8819);
and U8904 (N_8904,N_8869,N_8888);
or U8905 (N_8905,N_8802,N_8818);
nor U8906 (N_8906,N_8862,N_8816);
nand U8907 (N_8907,N_8840,N_8868);
nor U8908 (N_8908,N_8865,N_8856);
nand U8909 (N_8909,N_8817,N_8853);
or U8910 (N_8910,N_8836,N_8872);
nand U8911 (N_8911,N_8863,N_8895);
xor U8912 (N_8912,N_8878,N_8838);
and U8913 (N_8913,N_8841,N_8864);
nand U8914 (N_8914,N_8822,N_8839);
nand U8915 (N_8915,N_8899,N_8871);
nor U8916 (N_8916,N_8894,N_8881);
nand U8917 (N_8917,N_8820,N_8805);
nor U8918 (N_8918,N_8844,N_8875);
nand U8919 (N_8919,N_8889,N_8834);
nand U8920 (N_8920,N_8807,N_8854);
and U8921 (N_8921,N_8826,N_8809);
nor U8922 (N_8922,N_8815,N_8877);
and U8923 (N_8923,N_8835,N_8849);
nand U8924 (N_8924,N_8855,N_8885);
nand U8925 (N_8925,N_8803,N_8887);
nor U8926 (N_8926,N_8804,N_8861);
or U8927 (N_8927,N_8829,N_8896);
nor U8928 (N_8928,N_8870,N_8848);
nor U8929 (N_8929,N_8883,N_8821);
nand U8930 (N_8930,N_8800,N_8801);
nand U8931 (N_8931,N_8831,N_8846);
and U8932 (N_8932,N_8814,N_8825);
and U8933 (N_8933,N_8852,N_8811);
and U8934 (N_8934,N_8860,N_8813);
nand U8935 (N_8935,N_8806,N_8886);
or U8936 (N_8936,N_8867,N_8808);
and U8937 (N_8937,N_8876,N_8873);
and U8938 (N_8938,N_8851,N_8810);
nand U8939 (N_8939,N_8884,N_8845);
or U8940 (N_8940,N_8890,N_8843);
nand U8941 (N_8941,N_8832,N_8833);
or U8942 (N_8942,N_8891,N_8897);
and U8943 (N_8943,N_8824,N_8823);
and U8944 (N_8944,N_8866,N_8898);
and U8945 (N_8945,N_8827,N_8847);
and U8946 (N_8946,N_8842,N_8857);
or U8947 (N_8947,N_8892,N_8850);
nand U8948 (N_8948,N_8812,N_8893);
nor U8949 (N_8949,N_8858,N_8837);
and U8950 (N_8950,N_8828,N_8888);
or U8951 (N_8951,N_8840,N_8852);
and U8952 (N_8952,N_8864,N_8808);
nor U8953 (N_8953,N_8868,N_8816);
nand U8954 (N_8954,N_8896,N_8841);
nand U8955 (N_8955,N_8862,N_8873);
xnor U8956 (N_8956,N_8854,N_8882);
and U8957 (N_8957,N_8830,N_8802);
and U8958 (N_8958,N_8879,N_8899);
and U8959 (N_8959,N_8834,N_8809);
nor U8960 (N_8960,N_8832,N_8841);
nand U8961 (N_8961,N_8824,N_8812);
and U8962 (N_8962,N_8836,N_8893);
or U8963 (N_8963,N_8855,N_8899);
and U8964 (N_8964,N_8830,N_8890);
nor U8965 (N_8965,N_8801,N_8830);
nor U8966 (N_8966,N_8872,N_8843);
or U8967 (N_8967,N_8862,N_8896);
nand U8968 (N_8968,N_8816,N_8824);
nand U8969 (N_8969,N_8876,N_8886);
and U8970 (N_8970,N_8879,N_8835);
nand U8971 (N_8971,N_8885,N_8888);
or U8972 (N_8972,N_8860,N_8847);
and U8973 (N_8973,N_8836,N_8855);
nand U8974 (N_8974,N_8875,N_8896);
nand U8975 (N_8975,N_8855,N_8829);
nor U8976 (N_8976,N_8841,N_8820);
nand U8977 (N_8977,N_8811,N_8863);
and U8978 (N_8978,N_8849,N_8879);
nor U8979 (N_8979,N_8855,N_8861);
xnor U8980 (N_8980,N_8894,N_8890);
nor U8981 (N_8981,N_8889,N_8887);
nand U8982 (N_8982,N_8882,N_8802);
and U8983 (N_8983,N_8896,N_8860);
nand U8984 (N_8984,N_8870,N_8850);
nand U8985 (N_8985,N_8860,N_8880);
and U8986 (N_8986,N_8803,N_8857);
or U8987 (N_8987,N_8818,N_8816);
and U8988 (N_8988,N_8873,N_8825);
nand U8989 (N_8989,N_8821,N_8846);
and U8990 (N_8990,N_8876,N_8835);
or U8991 (N_8991,N_8890,N_8827);
or U8992 (N_8992,N_8831,N_8841);
or U8993 (N_8993,N_8897,N_8824);
or U8994 (N_8994,N_8806,N_8854);
nor U8995 (N_8995,N_8874,N_8811);
nand U8996 (N_8996,N_8858,N_8844);
nand U8997 (N_8997,N_8808,N_8844);
nand U8998 (N_8998,N_8807,N_8818);
nor U8999 (N_8999,N_8878,N_8830);
or U9000 (N_9000,N_8925,N_8951);
nand U9001 (N_9001,N_8940,N_8942);
nand U9002 (N_9002,N_8937,N_8914);
nor U9003 (N_9003,N_8955,N_8911);
nand U9004 (N_9004,N_8933,N_8997);
or U9005 (N_9005,N_8908,N_8974);
or U9006 (N_9006,N_8975,N_8988);
nor U9007 (N_9007,N_8993,N_8959);
nand U9008 (N_9008,N_8901,N_8947);
and U9009 (N_9009,N_8922,N_8961);
or U9010 (N_9010,N_8968,N_8987);
and U9011 (N_9011,N_8977,N_8913);
and U9012 (N_9012,N_8982,N_8966);
and U9013 (N_9013,N_8915,N_8992);
or U9014 (N_9014,N_8972,N_8960);
and U9015 (N_9015,N_8946,N_8917);
or U9016 (N_9016,N_8973,N_8967);
nor U9017 (N_9017,N_8998,N_8926);
nor U9018 (N_9018,N_8996,N_8905);
and U9019 (N_9019,N_8934,N_8989);
or U9020 (N_9020,N_8970,N_8938);
nor U9021 (N_9021,N_8980,N_8907);
or U9022 (N_9022,N_8924,N_8990);
nor U9023 (N_9023,N_8948,N_8981);
xnor U9024 (N_9024,N_8929,N_8927);
nor U9025 (N_9025,N_8920,N_8935);
and U9026 (N_9026,N_8958,N_8965);
or U9027 (N_9027,N_8909,N_8949);
nor U9028 (N_9028,N_8941,N_8903);
or U9029 (N_9029,N_8932,N_8912);
or U9030 (N_9030,N_8931,N_8956);
nand U9031 (N_9031,N_8976,N_8950);
or U9032 (N_9032,N_8936,N_8939);
or U9033 (N_9033,N_8945,N_8904);
and U9034 (N_9034,N_8930,N_8962);
or U9035 (N_9035,N_8985,N_8923);
nor U9036 (N_9036,N_8902,N_8971);
and U9037 (N_9037,N_8994,N_8963);
or U9038 (N_9038,N_8969,N_8954);
nand U9039 (N_9039,N_8999,N_8957);
or U9040 (N_9040,N_8983,N_8952);
or U9041 (N_9041,N_8921,N_8919);
and U9042 (N_9042,N_8991,N_8986);
nand U9043 (N_9043,N_8978,N_8928);
or U9044 (N_9044,N_8943,N_8918);
or U9045 (N_9045,N_8953,N_8984);
nand U9046 (N_9046,N_8906,N_8900);
nor U9047 (N_9047,N_8979,N_8964);
nor U9048 (N_9048,N_8995,N_8910);
and U9049 (N_9049,N_8944,N_8916);
nand U9050 (N_9050,N_8905,N_8910);
xnor U9051 (N_9051,N_8969,N_8980);
nor U9052 (N_9052,N_8995,N_8928);
or U9053 (N_9053,N_8945,N_8996);
nor U9054 (N_9054,N_8990,N_8975);
and U9055 (N_9055,N_8941,N_8926);
and U9056 (N_9056,N_8956,N_8905);
and U9057 (N_9057,N_8908,N_8903);
or U9058 (N_9058,N_8986,N_8914);
or U9059 (N_9059,N_8970,N_8962);
and U9060 (N_9060,N_8987,N_8939);
or U9061 (N_9061,N_8908,N_8997);
nor U9062 (N_9062,N_8952,N_8951);
and U9063 (N_9063,N_8950,N_8991);
or U9064 (N_9064,N_8970,N_8994);
nand U9065 (N_9065,N_8961,N_8920);
or U9066 (N_9066,N_8988,N_8954);
and U9067 (N_9067,N_8940,N_8903);
nor U9068 (N_9068,N_8953,N_8975);
nand U9069 (N_9069,N_8995,N_8961);
or U9070 (N_9070,N_8952,N_8928);
nand U9071 (N_9071,N_8932,N_8945);
nand U9072 (N_9072,N_8991,N_8948);
xor U9073 (N_9073,N_8977,N_8931);
and U9074 (N_9074,N_8997,N_8919);
and U9075 (N_9075,N_8916,N_8993);
nand U9076 (N_9076,N_8921,N_8973);
nand U9077 (N_9077,N_8914,N_8946);
or U9078 (N_9078,N_8955,N_8960);
nand U9079 (N_9079,N_8987,N_8936);
or U9080 (N_9080,N_8936,N_8901);
and U9081 (N_9081,N_8940,N_8931);
nor U9082 (N_9082,N_8914,N_8976);
and U9083 (N_9083,N_8962,N_8901);
nor U9084 (N_9084,N_8913,N_8975);
and U9085 (N_9085,N_8915,N_8973);
and U9086 (N_9086,N_8956,N_8989);
nor U9087 (N_9087,N_8908,N_8906);
or U9088 (N_9088,N_8988,N_8964);
or U9089 (N_9089,N_8979,N_8982);
xnor U9090 (N_9090,N_8952,N_8961);
and U9091 (N_9091,N_8908,N_8942);
nor U9092 (N_9092,N_8988,N_8967);
nor U9093 (N_9093,N_8941,N_8938);
nand U9094 (N_9094,N_8950,N_8969);
nor U9095 (N_9095,N_8949,N_8986);
and U9096 (N_9096,N_8974,N_8920);
nand U9097 (N_9097,N_8998,N_8942);
and U9098 (N_9098,N_8984,N_8960);
nand U9099 (N_9099,N_8972,N_8942);
nand U9100 (N_9100,N_9025,N_9006);
xor U9101 (N_9101,N_9050,N_9013);
or U9102 (N_9102,N_9067,N_9018);
nor U9103 (N_9103,N_9068,N_9074);
nand U9104 (N_9104,N_9017,N_9058);
nand U9105 (N_9105,N_9080,N_9044);
and U9106 (N_9106,N_9086,N_9037);
and U9107 (N_9107,N_9046,N_9053);
and U9108 (N_9108,N_9007,N_9008);
and U9109 (N_9109,N_9054,N_9031);
nand U9110 (N_9110,N_9004,N_9011);
nand U9111 (N_9111,N_9002,N_9066);
and U9112 (N_9112,N_9087,N_9069);
nand U9113 (N_9113,N_9033,N_9009);
nand U9114 (N_9114,N_9014,N_9073);
nand U9115 (N_9115,N_9052,N_9095);
and U9116 (N_9116,N_9015,N_9029);
nor U9117 (N_9117,N_9084,N_9085);
nand U9118 (N_9118,N_9049,N_9083);
nand U9119 (N_9119,N_9026,N_9056);
nor U9120 (N_9120,N_9065,N_9071);
nand U9121 (N_9121,N_9091,N_9036);
nor U9122 (N_9122,N_9059,N_9077);
xor U9123 (N_9123,N_9028,N_9062);
nor U9124 (N_9124,N_9010,N_9020);
and U9125 (N_9125,N_9097,N_9098);
nand U9126 (N_9126,N_9055,N_9070);
and U9127 (N_9127,N_9061,N_9089);
nor U9128 (N_9128,N_9032,N_9005);
nand U9129 (N_9129,N_9027,N_9003);
and U9130 (N_9130,N_9042,N_9021);
nor U9131 (N_9131,N_9040,N_9000);
nand U9132 (N_9132,N_9099,N_9043);
or U9133 (N_9133,N_9019,N_9024);
or U9134 (N_9134,N_9081,N_9057);
nand U9135 (N_9135,N_9038,N_9034);
nor U9136 (N_9136,N_9076,N_9001);
or U9137 (N_9137,N_9048,N_9092);
nand U9138 (N_9138,N_9012,N_9072);
or U9139 (N_9139,N_9041,N_9039);
or U9140 (N_9140,N_9045,N_9051);
nor U9141 (N_9141,N_9022,N_9075);
nand U9142 (N_9142,N_9096,N_9088);
or U9143 (N_9143,N_9093,N_9078);
and U9144 (N_9144,N_9016,N_9030);
and U9145 (N_9145,N_9079,N_9023);
and U9146 (N_9146,N_9094,N_9060);
nor U9147 (N_9147,N_9035,N_9047);
and U9148 (N_9148,N_9082,N_9090);
or U9149 (N_9149,N_9063,N_9064);
or U9150 (N_9150,N_9059,N_9010);
nor U9151 (N_9151,N_9014,N_9029);
or U9152 (N_9152,N_9002,N_9029);
and U9153 (N_9153,N_9006,N_9023);
or U9154 (N_9154,N_9073,N_9031);
nor U9155 (N_9155,N_9022,N_9024);
nand U9156 (N_9156,N_9059,N_9072);
or U9157 (N_9157,N_9006,N_9029);
nand U9158 (N_9158,N_9043,N_9090);
or U9159 (N_9159,N_9076,N_9074);
and U9160 (N_9160,N_9082,N_9092);
and U9161 (N_9161,N_9041,N_9079);
and U9162 (N_9162,N_9019,N_9022);
or U9163 (N_9163,N_9021,N_9093);
or U9164 (N_9164,N_9080,N_9038);
or U9165 (N_9165,N_9032,N_9001);
nor U9166 (N_9166,N_9068,N_9009);
or U9167 (N_9167,N_9064,N_9087);
or U9168 (N_9168,N_9079,N_9007);
nor U9169 (N_9169,N_9056,N_9024);
nand U9170 (N_9170,N_9040,N_9022);
nor U9171 (N_9171,N_9004,N_9002);
and U9172 (N_9172,N_9017,N_9016);
or U9173 (N_9173,N_9032,N_9041);
and U9174 (N_9174,N_9062,N_9083);
or U9175 (N_9175,N_9067,N_9005);
or U9176 (N_9176,N_9028,N_9035);
or U9177 (N_9177,N_9098,N_9045);
or U9178 (N_9178,N_9096,N_9018);
xor U9179 (N_9179,N_9002,N_9012);
nand U9180 (N_9180,N_9069,N_9056);
nor U9181 (N_9181,N_9088,N_9023);
or U9182 (N_9182,N_9013,N_9045);
or U9183 (N_9183,N_9010,N_9007);
or U9184 (N_9184,N_9082,N_9004);
nor U9185 (N_9185,N_9004,N_9060);
nor U9186 (N_9186,N_9015,N_9074);
or U9187 (N_9187,N_9077,N_9042);
and U9188 (N_9188,N_9004,N_9024);
and U9189 (N_9189,N_9057,N_9075);
and U9190 (N_9190,N_9009,N_9039);
nand U9191 (N_9191,N_9099,N_9049);
and U9192 (N_9192,N_9066,N_9044);
and U9193 (N_9193,N_9091,N_9031);
nand U9194 (N_9194,N_9018,N_9027);
or U9195 (N_9195,N_9002,N_9070);
and U9196 (N_9196,N_9001,N_9080);
nor U9197 (N_9197,N_9044,N_9091);
or U9198 (N_9198,N_9071,N_9037);
and U9199 (N_9199,N_9049,N_9036);
and U9200 (N_9200,N_9139,N_9113);
xnor U9201 (N_9201,N_9178,N_9103);
or U9202 (N_9202,N_9161,N_9123);
nor U9203 (N_9203,N_9153,N_9106);
nor U9204 (N_9204,N_9150,N_9131);
or U9205 (N_9205,N_9147,N_9171);
or U9206 (N_9206,N_9143,N_9107);
or U9207 (N_9207,N_9117,N_9145);
nor U9208 (N_9208,N_9124,N_9149);
or U9209 (N_9209,N_9180,N_9184);
nand U9210 (N_9210,N_9134,N_9186);
or U9211 (N_9211,N_9173,N_9125);
or U9212 (N_9212,N_9111,N_9104);
or U9213 (N_9213,N_9194,N_9154);
nor U9214 (N_9214,N_9105,N_9141);
nand U9215 (N_9215,N_9199,N_9108);
nor U9216 (N_9216,N_9151,N_9142);
nand U9217 (N_9217,N_9114,N_9115);
nor U9218 (N_9218,N_9198,N_9160);
nand U9219 (N_9219,N_9156,N_9167);
or U9220 (N_9220,N_9176,N_9177);
or U9221 (N_9221,N_9155,N_9126);
and U9222 (N_9222,N_9133,N_9182);
nor U9223 (N_9223,N_9165,N_9192);
or U9224 (N_9224,N_9118,N_9157);
nand U9225 (N_9225,N_9140,N_9196);
or U9226 (N_9226,N_9120,N_9185);
nor U9227 (N_9227,N_9130,N_9175);
nand U9228 (N_9228,N_9148,N_9144);
nor U9229 (N_9229,N_9179,N_9100);
nand U9230 (N_9230,N_9132,N_9166);
and U9231 (N_9231,N_9119,N_9135);
nand U9232 (N_9232,N_9189,N_9188);
nor U9233 (N_9233,N_9138,N_9169);
and U9234 (N_9234,N_9116,N_9170);
or U9235 (N_9235,N_9110,N_9197);
or U9236 (N_9236,N_9136,N_9195);
and U9237 (N_9237,N_9129,N_9174);
nand U9238 (N_9238,N_9137,N_9172);
nor U9239 (N_9239,N_9158,N_9162);
and U9240 (N_9240,N_9122,N_9181);
or U9241 (N_9241,N_9127,N_9102);
nand U9242 (N_9242,N_9146,N_9101);
or U9243 (N_9243,N_9163,N_9183);
and U9244 (N_9244,N_9159,N_9112);
or U9245 (N_9245,N_9193,N_9191);
nand U9246 (N_9246,N_9128,N_9164);
nor U9247 (N_9247,N_9168,N_9152);
or U9248 (N_9248,N_9190,N_9121);
nand U9249 (N_9249,N_9109,N_9187);
and U9250 (N_9250,N_9149,N_9173);
or U9251 (N_9251,N_9185,N_9152);
or U9252 (N_9252,N_9136,N_9143);
nand U9253 (N_9253,N_9135,N_9160);
or U9254 (N_9254,N_9154,N_9184);
nand U9255 (N_9255,N_9152,N_9188);
nor U9256 (N_9256,N_9165,N_9164);
or U9257 (N_9257,N_9166,N_9179);
or U9258 (N_9258,N_9180,N_9139);
nand U9259 (N_9259,N_9153,N_9166);
or U9260 (N_9260,N_9187,N_9110);
nand U9261 (N_9261,N_9109,N_9183);
or U9262 (N_9262,N_9157,N_9186);
and U9263 (N_9263,N_9159,N_9199);
and U9264 (N_9264,N_9115,N_9183);
nand U9265 (N_9265,N_9166,N_9109);
and U9266 (N_9266,N_9129,N_9135);
and U9267 (N_9267,N_9150,N_9186);
nor U9268 (N_9268,N_9185,N_9197);
nor U9269 (N_9269,N_9136,N_9151);
nor U9270 (N_9270,N_9159,N_9169);
and U9271 (N_9271,N_9170,N_9106);
nor U9272 (N_9272,N_9120,N_9145);
nand U9273 (N_9273,N_9135,N_9112);
nand U9274 (N_9274,N_9171,N_9102);
or U9275 (N_9275,N_9132,N_9111);
nand U9276 (N_9276,N_9168,N_9102);
nand U9277 (N_9277,N_9104,N_9199);
nor U9278 (N_9278,N_9150,N_9101);
and U9279 (N_9279,N_9107,N_9155);
and U9280 (N_9280,N_9166,N_9175);
or U9281 (N_9281,N_9148,N_9189);
and U9282 (N_9282,N_9194,N_9116);
or U9283 (N_9283,N_9134,N_9100);
or U9284 (N_9284,N_9168,N_9194);
or U9285 (N_9285,N_9184,N_9134);
or U9286 (N_9286,N_9125,N_9195);
nand U9287 (N_9287,N_9149,N_9172);
nor U9288 (N_9288,N_9134,N_9109);
nor U9289 (N_9289,N_9107,N_9137);
and U9290 (N_9290,N_9159,N_9173);
nand U9291 (N_9291,N_9146,N_9165);
or U9292 (N_9292,N_9152,N_9108);
nand U9293 (N_9293,N_9161,N_9167);
nor U9294 (N_9294,N_9144,N_9188);
nand U9295 (N_9295,N_9189,N_9142);
and U9296 (N_9296,N_9114,N_9112);
nor U9297 (N_9297,N_9162,N_9119);
and U9298 (N_9298,N_9108,N_9180);
nand U9299 (N_9299,N_9120,N_9155);
nand U9300 (N_9300,N_9292,N_9296);
nand U9301 (N_9301,N_9285,N_9235);
or U9302 (N_9302,N_9260,N_9211);
and U9303 (N_9303,N_9277,N_9244);
xor U9304 (N_9304,N_9262,N_9201);
nand U9305 (N_9305,N_9212,N_9224);
nand U9306 (N_9306,N_9246,N_9264);
or U9307 (N_9307,N_9297,N_9286);
and U9308 (N_9308,N_9233,N_9293);
nand U9309 (N_9309,N_9220,N_9214);
xnor U9310 (N_9310,N_9250,N_9278);
and U9311 (N_9311,N_9206,N_9268);
nand U9312 (N_9312,N_9275,N_9240);
nand U9313 (N_9313,N_9245,N_9215);
nor U9314 (N_9314,N_9259,N_9282);
nor U9315 (N_9315,N_9248,N_9256);
xor U9316 (N_9316,N_9251,N_9267);
nand U9317 (N_9317,N_9257,N_9208);
and U9318 (N_9318,N_9234,N_9271);
nand U9319 (N_9319,N_9290,N_9230);
nor U9320 (N_9320,N_9247,N_9219);
or U9321 (N_9321,N_9222,N_9284);
or U9322 (N_9322,N_9265,N_9291);
nand U9323 (N_9323,N_9203,N_9202);
and U9324 (N_9324,N_9226,N_9232);
nor U9325 (N_9325,N_9273,N_9241);
nor U9326 (N_9326,N_9204,N_9255);
nand U9327 (N_9327,N_9279,N_9263);
and U9328 (N_9328,N_9283,N_9205);
and U9329 (N_9329,N_9288,N_9200);
nand U9330 (N_9330,N_9258,N_9287);
and U9331 (N_9331,N_9217,N_9261);
or U9332 (N_9332,N_9229,N_9274);
nand U9333 (N_9333,N_9276,N_9231);
nor U9334 (N_9334,N_9242,N_9266);
and U9335 (N_9335,N_9269,N_9254);
xor U9336 (N_9336,N_9281,N_9227);
or U9337 (N_9337,N_9294,N_9272);
and U9338 (N_9338,N_9209,N_9249);
nand U9339 (N_9339,N_9213,N_9270);
nand U9340 (N_9340,N_9239,N_9280);
nand U9341 (N_9341,N_9207,N_9253);
or U9342 (N_9342,N_9243,N_9228);
nor U9343 (N_9343,N_9289,N_9237);
or U9344 (N_9344,N_9299,N_9223);
nand U9345 (N_9345,N_9221,N_9216);
or U9346 (N_9346,N_9218,N_9225);
nand U9347 (N_9347,N_9252,N_9295);
or U9348 (N_9348,N_9238,N_9298);
or U9349 (N_9349,N_9236,N_9210);
or U9350 (N_9350,N_9210,N_9291);
nand U9351 (N_9351,N_9242,N_9209);
or U9352 (N_9352,N_9222,N_9288);
nand U9353 (N_9353,N_9213,N_9217);
or U9354 (N_9354,N_9271,N_9250);
or U9355 (N_9355,N_9206,N_9207);
nor U9356 (N_9356,N_9224,N_9293);
nor U9357 (N_9357,N_9261,N_9228);
nor U9358 (N_9358,N_9207,N_9238);
nand U9359 (N_9359,N_9227,N_9284);
nand U9360 (N_9360,N_9253,N_9250);
and U9361 (N_9361,N_9294,N_9219);
and U9362 (N_9362,N_9293,N_9244);
nand U9363 (N_9363,N_9262,N_9204);
and U9364 (N_9364,N_9224,N_9226);
or U9365 (N_9365,N_9210,N_9211);
nor U9366 (N_9366,N_9234,N_9279);
or U9367 (N_9367,N_9257,N_9243);
nor U9368 (N_9368,N_9298,N_9204);
and U9369 (N_9369,N_9229,N_9217);
nor U9370 (N_9370,N_9247,N_9207);
or U9371 (N_9371,N_9282,N_9208);
nor U9372 (N_9372,N_9229,N_9281);
nor U9373 (N_9373,N_9226,N_9293);
nor U9374 (N_9374,N_9249,N_9232);
nor U9375 (N_9375,N_9221,N_9272);
nand U9376 (N_9376,N_9256,N_9271);
nand U9377 (N_9377,N_9201,N_9220);
nand U9378 (N_9378,N_9292,N_9224);
nand U9379 (N_9379,N_9213,N_9249);
or U9380 (N_9380,N_9233,N_9251);
and U9381 (N_9381,N_9270,N_9207);
nand U9382 (N_9382,N_9240,N_9226);
xnor U9383 (N_9383,N_9211,N_9204);
nor U9384 (N_9384,N_9202,N_9251);
or U9385 (N_9385,N_9211,N_9275);
xnor U9386 (N_9386,N_9277,N_9278);
nand U9387 (N_9387,N_9231,N_9212);
and U9388 (N_9388,N_9295,N_9203);
and U9389 (N_9389,N_9261,N_9294);
or U9390 (N_9390,N_9242,N_9243);
nand U9391 (N_9391,N_9257,N_9256);
and U9392 (N_9392,N_9267,N_9233);
nand U9393 (N_9393,N_9224,N_9247);
nand U9394 (N_9394,N_9227,N_9219);
and U9395 (N_9395,N_9202,N_9264);
and U9396 (N_9396,N_9234,N_9287);
nand U9397 (N_9397,N_9263,N_9238);
and U9398 (N_9398,N_9215,N_9219);
nand U9399 (N_9399,N_9252,N_9260);
or U9400 (N_9400,N_9301,N_9391);
and U9401 (N_9401,N_9374,N_9398);
nand U9402 (N_9402,N_9370,N_9372);
and U9403 (N_9403,N_9305,N_9304);
or U9404 (N_9404,N_9332,N_9365);
xor U9405 (N_9405,N_9348,N_9360);
nor U9406 (N_9406,N_9339,N_9335);
or U9407 (N_9407,N_9363,N_9327);
and U9408 (N_9408,N_9355,N_9345);
or U9409 (N_9409,N_9313,N_9342);
nor U9410 (N_9410,N_9340,N_9308);
and U9411 (N_9411,N_9315,N_9382);
nor U9412 (N_9412,N_9323,N_9344);
nand U9413 (N_9413,N_9383,N_9367);
nand U9414 (N_9414,N_9399,N_9351);
nand U9415 (N_9415,N_9333,N_9395);
and U9416 (N_9416,N_9371,N_9373);
nand U9417 (N_9417,N_9390,N_9359);
xnor U9418 (N_9418,N_9389,N_9311);
and U9419 (N_9419,N_9386,N_9364);
xor U9420 (N_9420,N_9381,N_9366);
nor U9421 (N_9421,N_9331,N_9312);
and U9422 (N_9422,N_9356,N_9352);
and U9423 (N_9423,N_9357,N_9337);
and U9424 (N_9424,N_9361,N_9393);
and U9425 (N_9425,N_9316,N_9336);
nor U9426 (N_9426,N_9314,N_9347);
nor U9427 (N_9427,N_9397,N_9343);
xnor U9428 (N_9428,N_9369,N_9309);
or U9429 (N_9429,N_9338,N_9346);
and U9430 (N_9430,N_9396,N_9328);
nand U9431 (N_9431,N_9350,N_9319);
nand U9432 (N_9432,N_9324,N_9392);
and U9433 (N_9433,N_9354,N_9303);
nor U9434 (N_9434,N_9325,N_9362);
and U9435 (N_9435,N_9377,N_9320);
or U9436 (N_9436,N_9378,N_9322);
and U9437 (N_9437,N_9379,N_9358);
nand U9438 (N_9438,N_9376,N_9353);
nand U9439 (N_9439,N_9317,N_9388);
and U9440 (N_9440,N_9310,N_9329);
and U9441 (N_9441,N_9321,N_9318);
or U9442 (N_9442,N_9334,N_9387);
and U9443 (N_9443,N_9349,N_9341);
or U9444 (N_9444,N_9385,N_9300);
and U9445 (N_9445,N_9375,N_9302);
nand U9446 (N_9446,N_9307,N_9326);
nor U9447 (N_9447,N_9380,N_9330);
and U9448 (N_9448,N_9394,N_9306);
and U9449 (N_9449,N_9368,N_9384);
or U9450 (N_9450,N_9302,N_9356);
nand U9451 (N_9451,N_9371,N_9310);
or U9452 (N_9452,N_9317,N_9302);
nor U9453 (N_9453,N_9361,N_9382);
or U9454 (N_9454,N_9394,N_9368);
or U9455 (N_9455,N_9325,N_9351);
and U9456 (N_9456,N_9399,N_9332);
nor U9457 (N_9457,N_9330,N_9348);
nor U9458 (N_9458,N_9375,N_9325);
xnor U9459 (N_9459,N_9386,N_9343);
or U9460 (N_9460,N_9344,N_9353);
and U9461 (N_9461,N_9392,N_9389);
and U9462 (N_9462,N_9361,N_9306);
and U9463 (N_9463,N_9378,N_9388);
and U9464 (N_9464,N_9388,N_9373);
nor U9465 (N_9465,N_9384,N_9389);
nand U9466 (N_9466,N_9301,N_9313);
nor U9467 (N_9467,N_9306,N_9337);
nand U9468 (N_9468,N_9357,N_9308);
or U9469 (N_9469,N_9318,N_9320);
and U9470 (N_9470,N_9314,N_9359);
nor U9471 (N_9471,N_9325,N_9339);
nor U9472 (N_9472,N_9342,N_9363);
or U9473 (N_9473,N_9322,N_9319);
and U9474 (N_9474,N_9347,N_9373);
or U9475 (N_9475,N_9369,N_9342);
nand U9476 (N_9476,N_9380,N_9335);
or U9477 (N_9477,N_9302,N_9348);
nand U9478 (N_9478,N_9309,N_9316);
nand U9479 (N_9479,N_9323,N_9360);
and U9480 (N_9480,N_9357,N_9303);
and U9481 (N_9481,N_9321,N_9368);
nor U9482 (N_9482,N_9343,N_9340);
nor U9483 (N_9483,N_9357,N_9382);
nand U9484 (N_9484,N_9393,N_9310);
and U9485 (N_9485,N_9338,N_9312);
nor U9486 (N_9486,N_9303,N_9341);
nand U9487 (N_9487,N_9362,N_9363);
nand U9488 (N_9488,N_9354,N_9338);
or U9489 (N_9489,N_9394,N_9338);
and U9490 (N_9490,N_9338,N_9322);
and U9491 (N_9491,N_9392,N_9359);
nand U9492 (N_9492,N_9398,N_9331);
and U9493 (N_9493,N_9326,N_9355);
nand U9494 (N_9494,N_9315,N_9333);
xnor U9495 (N_9495,N_9350,N_9393);
nand U9496 (N_9496,N_9392,N_9323);
nor U9497 (N_9497,N_9371,N_9389);
and U9498 (N_9498,N_9340,N_9306);
and U9499 (N_9499,N_9341,N_9340);
or U9500 (N_9500,N_9479,N_9480);
and U9501 (N_9501,N_9467,N_9497);
and U9502 (N_9502,N_9452,N_9473);
nand U9503 (N_9503,N_9432,N_9447);
nand U9504 (N_9504,N_9406,N_9465);
or U9505 (N_9505,N_9462,N_9449);
nand U9506 (N_9506,N_9491,N_9430);
or U9507 (N_9507,N_9468,N_9429);
nor U9508 (N_9508,N_9410,N_9419);
and U9509 (N_9509,N_9422,N_9400);
nor U9510 (N_9510,N_9427,N_9418);
or U9511 (N_9511,N_9482,N_9408);
and U9512 (N_9512,N_9414,N_9490);
or U9513 (N_9513,N_9412,N_9436);
and U9514 (N_9514,N_9454,N_9461);
and U9515 (N_9515,N_9416,N_9433);
nand U9516 (N_9516,N_9420,N_9435);
nand U9517 (N_9517,N_9474,N_9496);
nor U9518 (N_9518,N_9469,N_9428);
nor U9519 (N_9519,N_9456,N_9481);
nor U9520 (N_9520,N_9458,N_9489);
or U9521 (N_9521,N_9440,N_9403);
and U9522 (N_9522,N_9459,N_9424);
nor U9523 (N_9523,N_9402,N_9487);
and U9524 (N_9524,N_9426,N_9455);
nand U9525 (N_9525,N_9405,N_9475);
nand U9526 (N_9526,N_9446,N_9464);
nor U9527 (N_9527,N_9448,N_9450);
nor U9528 (N_9528,N_9498,N_9477);
nand U9529 (N_9529,N_9444,N_9486);
and U9530 (N_9530,N_9421,N_9443);
nor U9531 (N_9531,N_9434,N_9409);
nor U9532 (N_9532,N_9451,N_9488);
nor U9533 (N_9533,N_9413,N_9417);
or U9534 (N_9534,N_9439,N_9470);
nand U9535 (N_9535,N_9401,N_9495);
and U9536 (N_9536,N_9407,N_9476);
or U9537 (N_9537,N_9411,N_9438);
nand U9538 (N_9538,N_9478,N_9453);
nor U9539 (N_9539,N_9493,N_9442);
or U9540 (N_9540,N_9472,N_9483);
nor U9541 (N_9541,N_9445,N_9404);
or U9542 (N_9542,N_9466,N_9499);
nor U9543 (N_9543,N_9441,N_9431);
and U9544 (N_9544,N_9492,N_9457);
nand U9545 (N_9545,N_9485,N_9460);
or U9546 (N_9546,N_9484,N_9415);
nor U9547 (N_9547,N_9423,N_9471);
nor U9548 (N_9548,N_9437,N_9494);
nor U9549 (N_9549,N_9425,N_9463);
nor U9550 (N_9550,N_9448,N_9455);
and U9551 (N_9551,N_9451,N_9489);
or U9552 (N_9552,N_9491,N_9469);
nor U9553 (N_9553,N_9450,N_9440);
or U9554 (N_9554,N_9459,N_9467);
or U9555 (N_9555,N_9408,N_9478);
and U9556 (N_9556,N_9472,N_9435);
nand U9557 (N_9557,N_9494,N_9402);
and U9558 (N_9558,N_9489,N_9410);
nor U9559 (N_9559,N_9408,N_9428);
and U9560 (N_9560,N_9412,N_9472);
nor U9561 (N_9561,N_9433,N_9484);
or U9562 (N_9562,N_9433,N_9401);
nor U9563 (N_9563,N_9405,N_9487);
or U9564 (N_9564,N_9470,N_9401);
nor U9565 (N_9565,N_9463,N_9429);
nand U9566 (N_9566,N_9453,N_9456);
or U9567 (N_9567,N_9414,N_9450);
and U9568 (N_9568,N_9405,N_9469);
nand U9569 (N_9569,N_9430,N_9489);
nand U9570 (N_9570,N_9404,N_9468);
nand U9571 (N_9571,N_9459,N_9447);
and U9572 (N_9572,N_9419,N_9422);
nand U9573 (N_9573,N_9412,N_9402);
or U9574 (N_9574,N_9413,N_9453);
nor U9575 (N_9575,N_9477,N_9442);
nand U9576 (N_9576,N_9409,N_9406);
or U9577 (N_9577,N_9474,N_9468);
or U9578 (N_9578,N_9438,N_9403);
xnor U9579 (N_9579,N_9417,N_9420);
and U9580 (N_9580,N_9496,N_9484);
nor U9581 (N_9581,N_9453,N_9438);
and U9582 (N_9582,N_9438,N_9463);
nand U9583 (N_9583,N_9413,N_9494);
or U9584 (N_9584,N_9498,N_9415);
nand U9585 (N_9585,N_9423,N_9487);
nor U9586 (N_9586,N_9421,N_9428);
or U9587 (N_9587,N_9441,N_9421);
nor U9588 (N_9588,N_9469,N_9476);
nor U9589 (N_9589,N_9425,N_9462);
or U9590 (N_9590,N_9472,N_9467);
nor U9591 (N_9591,N_9473,N_9469);
and U9592 (N_9592,N_9419,N_9478);
nor U9593 (N_9593,N_9438,N_9457);
and U9594 (N_9594,N_9496,N_9410);
or U9595 (N_9595,N_9478,N_9456);
or U9596 (N_9596,N_9424,N_9457);
nand U9597 (N_9597,N_9430,N_9483);
nor U9598 (N_9598,N_9425,N_9435);
nor U9599 (N_9599,N_9495,N_9494);
nand U9600 (N_9600,N_9564,N_9569);
and U9601 (N_9601,N_9509,N_9532);
nand U9602 (N_9602,N_9575,N_9523);
and U9603 (N_9603,N_9522,N_9505);
nor U9604 (N_9604,N_9521,N_9546);
or U9605 (N_9605,N_9571,N_9535);
and U9606 (N_9606,N_9560,N_9584);
and U9607 (N_9607,N_9594,N_9570);
nand U9608 (N_9608,N_9565,N_9596);
nor U9609 (N_9609,N_9562,N_9538);
nand U9610 (N_9610,N_9589,N_9588);
nor U9611 (N_9611,N_9508,N_9536);
or U9612 (N_9612,N_9529,N_9520);
or U9613 (N_9613,N_9501,N_9574);
and U9614 (N_9614,N_9548,N_9507);
and U9615 (N_9615,N_9513,N_9540);
nor U9616 (N_9616,N_9518,N_9578);
nand U9617 (N_9617,N_9597,N_9544);
or U9618 (N_9618,N_9515,N_9561);
nor U9619 (N_9619,N_9517,N_9556);
nor U9620 (N_9620,N_9512,N_9581);
or U9621 (N_9621,N_9504,N_9549);
and U9622 (N_9622,N_9567,N_9554);
and U9623 (N_9623,N_9591,N_9526);
nor U9624 (N_9624,N_9582,N_9559);
and U9625 (N_9625,N_9587,N_9573);
or U9626 (N_9626,N_9595,N_9593);
or U9627 (N_9627,N_9527,N_9541);
nor U9628 (N_9628,N_9503,N_9531);
nor U9629 (N_9629,N_9547,N_9555);
nor U9630 (N_9630,N_9583,N_9528);
nand U9631 (N_9631,N_9580,N_9553);
nor U9632 (N_9632,N_9534,N_9577);
nor U9633 (N_9633,N_9542,N_9524);
nor U9634 (N_9634,N_9510,N_9599);
nand U9635 (N_9635,N_9519,N_9506);
nor U9636 (N_9636,N_9558,N_9551);
xnor U9637 (N_9637,N_9550,N_9500);
and U9638 (N_9638,N_9516,N_9543);
nand U9639 (N_9639,N_9579,N_9514);
and U9640 (N_9640,N_9590,N_9539);
nor U9641 (N_9641,N_9530,N_9545);
or U9642 (N_9642,N_9502,N_9566);
or U9643 (N_9643,N_9511,N_9576);
and U9644 (N_9644,N_9537,N_9598);
nor U9645 (N_9645,N_9563,N_9552);
xnor U9646 (N_9646,N_9572,N_9568);
nand U9647 (N_9647,N_9592,N_9533);
xor U9648 (N_9648,N_9586,N_9585);
and U9649 (N_9649,N_9525,N_9557);
nor U9650 (N_9650,N_9563,N_9546);
or U9651 (N_9651,N_9520,N_9550);
or U9652 (N_9652,N_9502,N_9506);
nor U9653 (N_9653,N_9555,N_9584);
nor U9654 (N_9654,N_9504,N_9535);
nor U9655 (N_9655,N_9506,N_9535);
nor U9656 (N_9656,N_9505,N_9562);
nor U9657 (N_9657,N_9594,N_9549);
or U9658 (N_9658,N_9549,N_9526);
nand U9659 (N_9659,N_9543,N_9560);
nand U9660 (N_9660,N_9512,N_9583);
nand U9661 (N_9661,N_9532,N_9557);
and U9662 (N_9662,N_9529,N_9509);
xor U9663 (N_9663,N_9597,N_9537);
nand U9664 (N_9664,N_9519,N_9538);
nor U9665 (N_9665,N_9566,N_9565);
or U9666 (N_9666,N_9525,N_9523);
nand U9667 (N_9667,N_9504,N_9508);
nand U9668 (N_9668,N_9510,N_9502);
and U9669 (N_9669,N_9548,N_9525);
and U9670 (N_9670,N_9582,N_9566);
nor U9671 (N_9671,N_9562,N_9571);
nand U9672 (N_9672,N_9594,N_9519);
nor U9673 (N_9673,N_9541,N_9540);
nor U9674 (N_9674,N_9505,N_9521);
or U9675 (N_9675,N_9518,N_9564);
nor U9676 (N_9676,N_9566,N_9501);
nor U9677 (N_9677,N_9504,N_9536);
nor U9678 (N_9678,N_9500,N_9529);
nand U9679 (N_9679,N_9578,N_9531);
and U9680 (N_9680,N_9581,N_9505);
or U9681 (N_9681,N_9553,N_9598);
or U9682 (N_9682,N_9589,N_9532);
nor U9683 (N_9683,N_9565,N_9591);
nand U9684 (N_9684,N_9536,N_9519);
nand U9685 (N_9685,N_9561,N_9566);
or U9686 (N_9686,N_9542,N_9529);
nand U9687 (N_9687,N_9596,N_9551);
and U9688 (N_9688,N_9578,N_9561);
nor U9689 (N_9689,N_9578,N_9508);
and U9690 (N_9690,N_9597,N_9575);
nor U9691 (N_9691,N_9516,N_9529);
or U9692 (N_9692,N_9511,N_9521);
nor U9693 (N_9693,N_9524,N_9515);
nand U9694 (N_9694,N_9534,N_9539);
and U9695 (N_9695,N_9527,N_9539);
and U9696 (N_9696,N_9596,N_9532);
nand U9697 (N_9697,N_9589,N_9542);
or U9698 (N_9698,N_9547,N_9511);
or U9699 (N_9699,N_9558,N_9555);
and U9700 (N_9700,N_9639,N_9630);
and U9701 (N_9701,N_9651,N_9680);
nand U9702 (N_9702,N_9600,N_9677);
and U9703 (N_9703,N_9683,N_9668);
nand U9704 (N_9704,N_9674,N_9637);
or U9705 (N_9705,N_9678,N_9687);
or U9706 (N_9706,N_9669,N_9656);
and U9707 (N_9707,N_9634,N_9629);
and U9708 (N_9708,N_9620,N_9684);
nor U9709 (N_9709,N_9698,N_9675);
and U9710 (N_9710,N_9641,N_9626);
or U9711 (N_9711,N_9670,N_9621);
xor U9712 (N_9712,N_9688,N_9661);
and U9713 (N_9713,N_9603,N_9608);
or U9714 (N_9714,N_9609,N_9618);
and U9715 (N_9715,N_9645,N_9633);
or U9716 (N_9716,N_9636,N_9648);
and U9717 (N_9717,N_9655,N_9664);
xor U9718 (N_9718,N_9671,N_9663);
xor U9719 (N_9719,N_9610,N_9686);
or U9720 (N_9720,N_9602,N_9622);
nand U9721 (N_9721,N_9647,N_9659);
nand U9722 (N_9722,N_9667,N_9654);
nor U9723 (N_9723,N_9628,N_9601);
xnor U9724 (N_9724,N_9644,N_9662);
nor U9725 (N_9725,N_9623,N_9643);
and U9726 (N_9726,N_9638,N_9657);
and U9727 (N_9727,N_9691,N_9606);
nand U9728 (N_9728,N_9632,N_9665);
nor U9729 (N_9729,N_9614,N_9619);
and U9730 (N_9730,N_9685,N_9660);
xnor U9731 (N_9731,N_9682,N_9693);
nand U9732 (N_9732,N_9690,N_9604);
nor U9733 (N_9733,N_9649,N_9697);
and U9734 (N_9734,N_9615,N_9653);
and U9735 (N_9735,N_9650,N_9611);
nand U9736 (N_9736,N_9627,N_9689);
nor U9737 (N_9737,N_9658,N_9613);
and U9738 (N_9738,N_9676,N_9624);
and U9739 (N_9739,N_9679,N_9616);
or U9740 (N_9740,N_9673,N_9607);
or U9741 (N_9741,N_9625,N_9681);
nand U9742 (N_9742,N_9699,N_9696);
nor U9743 (N_9743,N_9642,N_9694);
and U9744 (N_9744,N_9646,N_9640);
and U9745 (N_9745,N_9635,N_9695);
and U9746 (N_9746,N_9605,N_9652);
nand U9747 (N_9747,N_9631,N_9672);
nor U9748 (N_9748,N_9666,N_9612);
nor U9749 (N_9749,N_9617,N_9692);
or U9750 (N_9750,N_9613,N_9639);
and U9751 (N_9751,N_9604,N_9687);
or U9752 (N_9752,N_9621,N_9665);
or U9753 (N_9753,N_9660,N_9616);
nand U9754 (N_9754,N_9647,N_9679);
nand U9755 (N_9755,N_9634,N_9696);
nand U9756 (N_9756,N_9610,N_9676);
nand U9757 (N_9757,N_9612,N_9693);
or U9758 (N_9758,N_9660,N_9654);
or U9759 (N_9759,N_9667,N_9670);
nand U9760 (N_9760,N_9686,N_9690);
nor U9761 (N_9761,N_9640,N_9630);
nand U9762 (N_9762,N_9631,N_9619);
nand U9763 (N_9763,N_9627,N_9648);
or U9764 (N_9764,N_9602,N_9699);
nand U9765 (N_9765,N_9677,N_9699);
or U9766 (N_9766,N_9653,N_9677);
nor U9767 (N_9767,N_9677,N_9611);
nor U9768 (N_9768,N_9606,N_9695);
or U9769 (N_9769,N_9616,N_9607);
nand U9770 (N_9770,N_9672,N_9693);
nand U9771 (N_9771,N_9644,N_9674);
nand U9772 (N_9772,N_9643,N_9658);
and U9773 (N_9773,N_9646,N_9675);
nand U9774 (N_9774,N_9679,N_9698);
nand U9775 (N_9775,N_9665,N_9638);
or U9776 (N_9776,N_9636,N_9620);
nand U9777 (N_9777,N_9617,N_9642);
and U9778 (N_9778,N_9603,N_9605);
nand U9779 (N_9779,N_9616,N_9647);
and U9780 (N_9780,N_9611,N_9667);
nand U9781 (N_9781,N_9669,N_9651);
nand U9782 (N_9782,N_9639,N_9647);
nor U9783 (N_9783,N_9676,N_9654);
or U9784 (N_9784,N_9694,N_9603);
nor U9785 (N_9785,N_9641,N_9672);
nor U9786 (N_9786,N_9673,N_9679);
nor U9787 (N_9787,N_9600,N_9669);
nor U9788 (N_9788,N_9620,N_9608);
nor U9789 (N_9789,N_9663,N_9669);
or U9790 (N_9790,N_9624,N_9609);
nand U9791 (N_9791,N_9613,N_9637);
or U9792 (N_9792,N_9669,N_9649);
nor U9793 (N_9793,N_9659,N_9676);
nor U9794 (N_9794,N_9668,N_9684);
or U9795 (N_9795,N_9665,N_9684);
and U9796 (N_9796,N_9645,N_9616);
nor U9797 (N_9797,N_9639,N_9635);
and U9798 (N_9798,N_9663,N_9615);
or U9799 (N_9799,N_9692,N_9684);
or U9800 (N_9800,N_9722,N_9782);
and U9801 (N_9801,N_9794,N_9770);
and U9802 (N_9802,N_9743,N_9741);
or U9803 (N_9803,N_9729,N_9777);
nand U9804 (N_9804,N_9793,N_9749);
or U9805 (N_9805,N_9748,N_9764);
nand U9806 (N_9806,N_9763,N_9751);
nand U9807 (N_9807,N_9740,N_9715);
nor U9808 (N_9808,N_9765,N_9775);
and U9809 (N_9809,N_9732,N_9727);
nor U9810 (N_9810,N_9772,N_9720);
nor U9811 (N_9811,N_9768,N_9735);
and U9812 (N_9812,N_9713,N_9788);
nand U9813 (N_9813,N_9787,N_9718);
or U9814 (N_9814,N_9711,N_9795);
nor U9815 (N_9815,N_9716,N_9717);
and U9816 (N_9816,N_9706,N_9708);
and U9817 (N_9817,N_9734,N_9744);
or U9818 (N_9818,N_9726,N_9756);
nor U9819 (N_9819,N_9730,N_9789);
and U9820 (N_9820,N_9725,N_9738);
nor U9821 (N_9821,N_9773,N_9737);
nand U9822 (N_9822,N_9753,N_9701);
and U9823 (N_9823,N_9707,N_9742);
xor U9824 (N_9824,N_9728,N_9745);
nor U9825 (N_9825,N_9778,N_9719);
nand U9826 (N_9826,N_9783,N_9731);
or U9827 (N_9827,N_9771,N_9724);
and U9828 (N_9828,N_9797,N_9761);
nor U9829 (N_9829,N_9784,N_9774);
and U9830 (N_9830,N_9733,N_9798);
or U9831 (N_9831,N_9747,N_9752);
nand U9832 (N_9832,N_9700,N_9757);
nor U9833 (N_9833,N_9760,N_9766);
nor U9834 (N_9834,N_9791,N_9785);
or U9835 (N_9835,N_9712,N_9736);
and U9836 (N_9836,N_9780,N_9709);
or U9837 (N_9837,N_9704,N_9796);
or U9838 (N_9838,N_9779,N_9762);
and U9839 (N_9839,N_9714,N_9710);
or U9840 (N_9840,N_9767,N_9723);
nand U9841 (N_9841,N_9759,N_9792);
nor U9842 (N_9842,N_9703,N_9746);
nor U9843 (N_9843,N_9799,N_9750);
nand U9844 (N_9844,N_9776,N_9754);
nand U9845 (N_9845,N_9769,N_9702);
or U9846 (N_9846,N_9705,N_9739);
nor U9847 (N_9847,N_9781,N_9721);
xnor U9848 (N_9848,N_9758,N_9755);
nor U9849 (N_9849,N_9786,N_9790);
and U9850 (N_9850,N_9708,N_9738);
nor U9851 (N_9851,N_9744,N_9750);
nand U9852 (N_9852,N_9773,N_9789);
and U9853 (N_9853,N_9781,N_9785);
or U9854 (N_9854,N_9766,N_9733);
nand U9855 (N_9855,N_9775,N_9753);
or U9856 (N_9856,N_9744,N_9714);
nor U9857 (N_9857,N_9775,N_9790);
or U9858 (N_9858,N_9705,N_9745);
or U9859 (N_9859,N_9749,N_9739);
and U9860 (N_9860,N_9735,N_9779);
nor U9861 (N_9861,N_9722,N_9769);
nor U9862 (N_9862,N_9704,N_9755);
and U9863 (N_9863,N_9783,N_9748);
nand U9864 (N_9864,N_9774,N_9738);
nand U9865 (N_9865,N_9775,N_9702);
nand U9866 (N_9866,N_9709,N_9787);
or U9867 (N_9867,N_9764,N_9762);
and U9868 (N_9868,N_9739,N_9707);
nand U9869 (N_9869,N_9747,N_9702);
nor U9870 (N_9870,N_9799,N_9795);
and U9871 (N_9871,N_9718,N_9702);
or U9872 (N_9872,N_9726,N_9797);
or U9873 (N_9873,N_9789,N_9772);
nor U9874 (N_9874,N_9702,N_9720);
nand U9875 (N_9875,N_9783,N_9706);
nand U9876 (N_9876,N_9748,N_9746);
nand U9877 (N_9877,N_9739,N_9717);
or U9878 (N_9878,N_9727,N_9763);
and U9879 (N_9879,N_9760,N_9762);
or U9880 (N_9880,N_9785,N_9727);
nor U9881 (N_9881,N_9774,N_9719);
and U9882 (N_9882,N_9729,N_9750);
nor U9883 (N_9883,N_9743,N_9769);
nand U9884 (N_9884,N_9760,N_9730);
nand U9885 (N_9885,N_9705,N_9784);
xnor U9886 (N_9886,N_9739,N_9796);
nor U9887 (N_9887,N_9737,N_9785);
nor U9888 (N_9888,N_9717,N_9784);
nor U9889 (N_9889,N_9759,N_9788);
nand U9890 (N_9890,N_9770,N_9718);
nand U9891 (N_9891,N_9793,N_9724);
nand U9892 (N_9892,N_9701,N_9788);
nand U9893 (N_9893,N_9754,N_9731);
and U9894 (N_9894,N_9745,N_9765);
nor U9895 (N_9895,N_9732,N_9759);
nand U9896 (N_9896,N_9798,N_9741);
and U9897 (N_9897,N_9785,N_9782);
nor U9898 (N_9898,N_9748,N_9739);
nand U9899 (N_9899,N_9769,N_9724);
nand U9900 (N_9900,N_9812,N_9814);
nand U9901 (N_9901,N_9840,N_9862);
or U9902 (N_9902,N_9893,N_9844);
xor U9903 (N_9903,N_9889,N_9810);
nand U9904 (N_9904,N_9819,N_9859);
and U9905 (N_9905,N_9850,N_9895);
nor U9906 (N_9906,N_9891,N_9864);
nor U9907 (N_9907,N_9865,N_9899);
nand U9908 (N_9908,N_9834,N_9830);
nor U9909 (N_9909,N_9890,N_9871);
nor U9910 (N_9910,N_9820,N_9885);
nand U9911 (N_9911,N_9887,N_9855);
and U9912 (N_9912,N_9881,N_9858);
nand U9913 (N_9913,N_9886,N_9898);
nand U9914 (N_9914,N_9868,N_9822);
and U9915 (N_9915,N_9831,N_9808);
nor U9916 (N_9916,N_9807,N_9870);
xnor U9917 (N_9917,N_9860,N_9854);
nand U9918 (N_9918,N_9805,N_9828);
nor U9919 (N_9919,N_9836,N_9832);
and U9920 (N_9920,N_9880,N_9888);
nor U9921 (N_9921,N_9827,N_9835);
xor U9922 (N_9922,N_9802,N_9843);
and U9923 (N_9923,N_9826,N_9824);
or U9924 (N_9924,N_9892,N_9853);
or U9925 (N_9925,N_9866,N_9845);
nand U9926 (N_9926,N_9849,N_9823);
and U9927 (N_9927,N_9878,N_9882);
nor U9928 (N_9928,N_9809,N_9896);
or U9929 (N_9929,N_9872,N_9837);
and U9930 (N_9930,N_9833,N_9873);
or U9931 (N_9931,N_9884,N_9848);
or U9932 (N_9932,N_9816,N_9879);
and U9933 (N_9933,N_9801,N_9829);
and U9934 (N_9934,N_9897,N_9851);
nand U9935 (N_9935,N_9818,N_9800);
or U9936 (N_9936,N_9883,N_9869);
and U9937 (N_9937,N_9846,N_9857);
and U9938 (N_9938,N_9856,N_9852);
or U9939 (N_9939,N_9867,N_9863);
or U9940 (N_9940,N_9804,N_9838);
and U9941 (N_9941,N_9806,N_9861);
or U9942 (N_9942,N_9821,N_9842);
and U9943 (N_9943,N_9811,N_9874);
or U9944 (N_9944,N_9815,N_9875);
nor U9945 (N_9945,N_9841,N_9817);
and U9946 (N_9946,N_9839,N_9894);
nor U9947 (N_9947,N_9803,N_9877);
or U9948 (N_9948,N_9813,N_9825);
and U9949 (N_9949,N_9847,N_9876);
or U9950 (N_9950,N_9825,N_9864);
nand U9951 (N_9951,N_9816,N_9890);
and U9952 (N_9952,N_9889,N_9898);
nand U9953 (N_9953,N_9817,N_9839);
xnor U9954 (N_9954,N_9839,N_9886);
and U9955 (N_9955,N_9857,N_9852);
nand U9956 (N_9956,N_9815,N_9882);
and U9957 (N_9957,N_9899,N_9885);
or U9958 (N_9958,N_9842,N_9824);
nand U9959 (N_9959,N_9835,N_9857);
or U9960 (N_9960,N_9854,N_9846);
and U9961 (N_9961,N_9841,N_9835);
or U9962 (N_9962,N_9817,N_9879);
nand U9963 (N_9963,N_9829,N_9807);
nand U9964 (N_9964,N_9826,N_9846);
or U9965 (N_9965,N_9807,N_9884);
and U9966 (N_9966,N_9888,N_9860);
nand U9967 (N_9967,N_9830,N_9815);
nand U9968 (N_9968,N_9804,N_9854);
or U9969 (N_9969,N_9800,N_9882);
nor U9970 (N_9970,N_9815,N_9872);
or U9971 (N_9971,N_9860,N_9834);
or U9972 (N_9972,N_9850,N_9800);
nand U9973 (N_9973,N_9827,N_9842);
nor U9974 (N_9974,N_9800,N_9883);
or U9975 (N_9975,N_9825,N_9820);
nand U9976 (N_9976,N_9884,N_9881);
or U9977 (N_9977,N_9841,N_9885);
nor U9978 (N_9978,N_9897,N_9824);
or U9979 (N_9979,N_9846,N_9895);
and U9980 (N_9980,N_9812,N_9876);
and U9981 (N_9981,N_9872,N_9821);
nor U9982 (N_9982,N_9827,N_9893);
or U9983 (N_9983,N_9817,N_9897);
xor U9984 (N_9984,N_9848,N_9849);
and U9985 (N_9985,N_9841,N_9881);
and U9986 (N_9986,N_9844,N_9831);
nand U9987 (N_9987,N_9890,N_9898);
and U9988 (N_9988,N_9872,N_9874);
nor U9989 (N_9989,N_9833,N_9851);
nor U9990 (N_9990,N_9875,N_9872);
or U9991 (N_9991,N_9805,N_9852);
nand U9992 (N_9992,N_9829,N_9835);
nand U9993 (N_9993,N_9886,N_9861);
or U9994 (N_9994,N_9813,N_9868);
and U9995 (N_9995,N_9889,N_9802);
nand U9996 (N_9996,N_9865,N_9884);
and U9997 (N_9997,N_9889,N_9819);
nor U9998 (N_9998,N_9808,N_9869);
nand U9999 (N_9999,N_9898,N_9874);
xnor UO_0 (O_0,N_9906,N_9913);
nor UO_1 (O_1,N_9998,N_9951);
and UO_2 (O_2,N_9964,N_9975);
nand UO_3 (O_3,N_9977,N_9979);
and UO_4 (O_4,N_9920,N_9991);
or UO_5 (O_5,N_9994,N_9970);
or UO_6 (O_6,N_9936,N_9927);
and UO_7 (O_7,N_9972,N_9909);
nor UO_8 (O_8,N_9945,N_9955);
nand UO_9 (O_9,N_9956,N_9938);
nand UO_10 (O_10,N_9971,N_9931);
nand UO_11 (O_11,N_9905,N_9999);
nand UO_12 (O_12,N_9980,N_9940);
and UO_13 (O_13,N_9922,N_9966);
nor UO_14 (O_14,N_9982,N_9904);
or UO_15 (O_15,N_9919,N_9932);
and UO_16 (O_16,N_9993,N_9948);
and UO_17 (O_17,N_9928,N_9923);
nand UO_18 (O_18,N_9984,N_9992);
nor UO_19 (O_19,N_9987,N_9926);
nor UO_20 (O_20,N_9974,N_9934);
xnor UO_21 (O_21,N_9953,N_9969);
xor UO_22 (O_22,N_9910,N_9986);
xnor UO_23 (O_23,N_9960,N_9958);
nor UO_24 (O_24,N_9973,N_9989);
and UO_25 (O_25,N_9917,N_9942);
or UO_26 (O_26,N_9968,N_9985);
or UO_27 (O_27,N_9959,N_9925);
nand UO_28 (O_28,N_9978,N_9911);
nor UO_29 (O_29,N_9939,N_9907);
nand UO_30 (O_30,N_9933,N_9963);
nor UO_31 (O_31,N_9983,N_9947);
and UO_32 (O_32,N_9962,N_9912);
or UO_33 (O_33,N_9952,N_9943);
and UO_34 (O_34,N_9954,N_9957);
and UO_35 (O_35,N_9997,N_9967);
or UO_36 (O_36,N_9990,N_9981);
nand UO_37 (O_37,N_9915,N_9949);
and UO_38 (O_38,N_9908,N_9921);
and UO_39 (O_39,N_9901,N_9930);
nand UO_40 (O_40,N_9996,N_9937);
xnor UO_41 (O_41,N_9988,N_9961);
nand UO_42 (O_42,N_9902,N_9916);
nand UO_43 (O_43,N_9903,N_9935);
and UO_44 (O_44,N_9929,N_9946);
and UO_45 (O_45,N_9941,N_9944);
nor UO_46 (O_46,N_9918,N_9995);
or UO_47 (O_47,N_9965,N_9914);
nand UO_48 (O_48,N_9976,N_9950);
and UO_49 (O_49,N_9900,N_9924);
and UO_50 (O_50,N_9993,N_9979);
nand UO_51 (O_51,N_9940,N_9986);
or UO_52 (O_52,N_9972,N_9963);
and UO_53 (O_53,N_9994,N_9954);
or UO_54 (O_54,N_9956,N_9996);
nand UO_55 (O_55,N_9900,N_9979);
or UO_56 (O_56,N_9915,N_9925);
and UO_57 (O_57,N_9958,N_9931);
nand UO_58 (O_58,N_9962,N_9922);
or UO_59 (O_59,N_9901,N_9941);
and UO_60 (O_60,N_9900,N_9943);
and UO_61 (O_61,N_9959,N_9939);
nor UO_62 (O_62,N_9964,N_9909);
nor UO_63 (O_63,N_9901,N_9970);
nor UO_64 (O_64,N_9981,N_9919);
nand UO_65 (O_65,N_9912,N_9964);
nor UO_66 (O_66,N_9921,N_9958);
nand UO_67 (O_67,N_9989,N_9937);
and UO_68 (O_68,N_9981,N_9956);
and UO_69 (O_69,N_9991,N_9931);
nand UO_70 (O_70,N_9923,N_9936);
nand UO_71 (O_71,N_9964,N_9916);
nand UO_72 (O_72,N_9957,N_9964);
xor UO_73 (O_73,N_9971,N_9973);
nor UO_74 (O_74,N_9944,N_9912);
and UO_75 (O_75,N_9983,N_9964);
or UO_76 (O_76,N_9929,N_9994);
nand UO_77 (O_77,N_9901,N_9966);
nor UO_78 (O_78,N_9904,N_9990);
nand UO_79 (O_79,N_9933,N_9905);
nor UO_80 (O_80,N_9924,N_9956);
or UO_81 (O_81,N_9905,N_9953);
or UO_82 (O_82,N_9982,N_9944);
or UO_83 (O_83,N_9979,N_9963);
or UO_84 (O_84,N_9905,N_9943);
nand UO_85 (O_85,N_9945,N_9905);
nor UO_86 (O_86,N_9983,N_9925);
or UO_87 (O_87,N_9908,N_9987);
and UO_88 (O_88,N_9992,N_9901);
nor UO_89 (O_89,N_9909,N_9908);
and UO_90 (O_90,N_9929,N_9967);
or UO_91 (O_91,N_9980,N_9911);
nor UO_92 (O_92,N_9958,N_9927);
nand UO_93 (O_93,N_9964,N_9955);
or UO_94 (O_94,N_9967,N_9998);
and UO_95 (O_95,N_9959,N_9921);
nor UO_96 (O_96,N_9914,N_9934);
or UO_97 (O_97,N_9907,N_9941);
nand UO_98 (O_98,N_9993,N_9995);
xor UO_99 (O_99,N_9933,N_9934);
nand UO_100 (O_100,N_9981,N_9909);
xor UO_101 (O_101,N_9902,N_9987);
and UO_102 (O_102,N_9910,N_9966);
nor UO_103 (O_103,N_9922,N_9959);
nor UO_104 (O_104,N_9955,N_9986);
and UO_105 (O_105,N_9944,N_9988);
nand UO_106 (O_106,N_9997,N_9901);
nand UO_107 (O_107,N_9975,N_9966);
or UO_108 (O_108,N_9978,N_9989);
nand UO_109 (O_109,N_9948,N_9901);
or UO_110 (O_110,N_9904,N_9966);
and UO_111 (O_111,N_9974,N_9953);
nand UO_112 (O_112,N_9975,N_9933);
xor UO_113 (O_113,N_9951,N_9979);
and UO_114 (O_114,N_9907,N_9934);
nor UO_115 (O_115,N_9998,N_9989);
or UO_116 (O_116,N_9924,N_9951);
or UO_117 (O_117,N_9973,N_9947);
or UO_118 (O_118,N_9996,N_9979);
xor UO_119 (O_119,N_9934,N_9962);
nor UO_120 (O_120,N_9922,N_9957);
and UO_121 (O_121,N_9993,N_9957);
nor UO_122 (O_122,N_9921,N_9987);
and UO_123 (O_123,N_9940,N_9976);
xor UO_124 (O_124,N_9987,N_9910);
or UO_125 (O_125,N_9946,N_9955);
nand UO_126 (O_126,N_9976,N_9975);
nor UO_127 (O_127,N_9913,N_9910);
nand UO_128 (O_128,N_9973,N_9946);
and UO_129 (O_129,N_9944,N_9978);
xor UO_130 (O_130,N_9983,N_9987);
nand UO_131 (O_131,N_9925,N_9969);
and UO_132 (O_132,N_9924,N_9938);
and UO_133 (O_133,N_9947,N_9956);
or UO_134 (O_134,N_9961,N_9964);
nor UO_135 (O_135,N_9956,N_9923);
or UO_136 (O_136,N_9910,N_9900);
xor UO_137 (O_137,N_9922,N_9982);
and UO_138 (O_138,N_9919,N_9989);
nand UO_139 (O_139,N_9915,N_9978);
or UO_140 (O_140,N_9956,N_9945);
or UO_141 (O_141,N_9960,N_9910);
nand UO_142 (O_142,N_9915,N_9993);
or UO_143 (O_143,N_9904,N_9955);
nor UO_144 (O_144,N_9981,N_9918);
and UO_145 (O_145,N_9981,N_9942);
and UO_146 (O_146,N_9972,N_9956);
nand UO_147 (O_147,N_9983,N_9970);
nand UO_148 (O_148,N_9984,N_9927);
nand UO_149 (O_149,N_9928,N_9986);
nor UO_150 (O_150,N_9908,N_9997);
nand UO_151 (O_151,N_9930,N_9909);
nor UO_152 (O_152,N_9919,N_9920);
and UO_153 (O_153,N_9926,N_9951);
nor UO_154 (O_154,N_9979,N_9950);
or UO_155 (O_155,N_9990,N_9915);
or UO_156 (O_156,N_9967,N_9953);
nor UO_157 (O_157,N_9995,N_9923);
nand UO_158 (O_158,N_9903,N_9900);
and UO_159 (O_159,N_9930,N_9988);
nand UO_160 (O_160,N_9966,N_9970);
and UO_161 (O_161,N_9968,N_9996);
nand UO_162 (O_162,N_9994,N_9923);
and UO_163 (O_163,N_9937,N_9981);
and UO_164 (O_164,N_9948,N_9932);
and UO_165 (O_165,N_9949,N_9937);
nand UO_166 (O_166,N_9955,N_9906);
nand UO_167 (O_167,N_9944,N_9989);
or UO_168 (O_168,N_9956,N_9943);
or UO_169 (O_169,N_9938,N_9917);
xor UO_170 (O_170,N_9902,N_9946);
nand UO_171 (O_171,N_9976,N_9967);
nor UO_172 (O_172,N_9924,N_9992);
nand UO_173 (O_173,N_9975,N_9921);
nand UO_174 (O_174,N_9943,N_9979);
nand UO_175 (O_175,N_9981,N_9984);
or UO_176 (O_176,N_9959,N_9919);
nand UO_177 (O_177,N_9903,N_9941);
or UO_178 (O_178,N_9971,N_9946);
nand UO_179 (O_179,N_9993,N_9972);
nand UO_180 (O_180,N_9963,N_9920);
nor UO_181 (O_181,N_9923,N_9947);
and UO_182 (O_182,N_9973,N_9979);
nor UO_183 (O_183,N_9982,N_9985);
nand UO_184 (O_184,N_9923,N_9946);
nand UO_185 (O_185,N_9942,N_9928);
nand UO_186 (O_186,N_9912,N_9981);
and UO_187 (O_187,N_9967,N_9961);
and UO_188 (O_188,N_9980,N_9921);
nand UO_189 (O_189,N_9990,N_9906);
nand UO_190 (O_190,N_9927,N_9957);
nor UO_191 (O_191,N_9920,N_9949);
nor UO_192 (O_192,N_9906,N_9976);
or UO_193 (O_193,N_9934,N_9956);
and UO_194 (O_194,N_9902,N_9974);
nand UO_195 (O_195,N_9931,N_9954);
nor UO_196 (O_196,N_9976,N_9935);
nand UO_197 (O_197,N_9960,N_9941);
nand UO_198 (O_198,N_9985,N_9967);
or UO_199 (O_199,N_9923,N_9911);
nor UO_200 (O_200,N_9912,N_9907);
xnor UO_201 (O_201,N_9916,N_9937);
nand UO_202 (O_202,N_9935,N_9985);
and UO_203 (O_203,N_9965,N_9909);
nor UO_204 (O_204,N_9901,N_9944);
and UO_205 (O_205,N_9957,N_9997);
nand UO_206 (O_206,N_9959,N_9984);
and UO_207 (O_207,N_9936,N_9991);
nor UO_208 (O_208,N_9936,N_9922);
or UO_209 (O_209,N_9954,N_9916);
nand UO_210 (O_210,N_9927,N_9926);
or UO_211 (O_211,N_9980,N_9907);
nor UO_212 (O_212,N_9999,N_9966);
and UO_213 (O_213,N_9991,N_9987);
or UO_214 (O_214,N_9963,N_9903);
and UO_215 (O_215,N_9998,N_9960);
nand UO_216 (O_216,N_9929,N_9973);
nor UO_217 (O_217,N_9946,N_9937);
nor UO_218 (O_218,N_9902,N_9997);
nand UO_219 (O_219,N_9949,N_9964);
nor UO_220 (O_220,N_9957,N_9902);
or UO_221 (O_221,N_9960,N_9918);
or UO_222 (O_222,N_9944,N_9910);
nand UO_223 (O_223,N_9900,N_9963);
xnor UO_224 (O_224,N_9920,N_9952);
or UO_225 (O_225,N_9948,N_9923);
nor UO_226 (O_226,N_9986,N_9977);
and UO_227 (O_227,N_9918,N_9958);
nor UO_228 (O_228,N_9942,N_9950);
and UO_229 (O_229,N_9936,N_9904);
and UO_230 (O_230,N_9911,N_9966);
nor UO_231 (O_231,N_9928,N_9945);
or UO_232 (O_232,N_9924,N_9998);
or UO_233 (O_233,N_9970,N_9941);
nand UO_234 (O_234,N_9990,N_9901);
and UO_235 (O_235,N_9919,N_9914);
nor UO_236 (O_236,N_9935,N_9981);
and UO_237 (O_237,N_9982,N_9936);
nor UO_238 (O_238,N_9905,N_9964);
nor UO_239 (O_239,N_9903,N_9989);
nand UO_240 (O_240,N_9996,N_9930);
and UO_241 (O_241,N_9961,N_9957);
and UO_242 (O_242,N_9938,N_9922);
nor UO_243 (O_243,N_9962,N_9937);
or UO_244 (O_244,N_9963,N_9904);
or UO_245 (O_245,N_9931,N_9939);
nor UO_246 (O_246,N_9994,N_9992);
and UO_247 (O_247,N_9911,N_9913);
nand UO_248 (O_248,N_9994,N_9930);
nand UO_249 (O_249,N_9937,N_9923);
nor UO_250 (O_250,N_9911,N_9960);
or UO_251 (O_251,N_9967,N_9919);
or UO_252 (O_252,N_9902,N_9900);
and UO_253 (O_253,N_9901,N_9961);
or UO_254 (O_254,N_9948,N_9945);
and UO_255 (O_255,N_9911,N_9904);
and UO_256 (O_256,N_9972,N_9908);
nor UO_257 (O_257,N_9955,N_9925);
nor UO_258 (O_258,N_9971,N_9993);
nand UO_259 (O_259,N_9917,N_9981);
and UO_260 (O_260,N_9970,N_9932);
nor UO_261 (O_261,N_9902,N_9949);
nor UO_262 (O_262,N_9995,N_9957);
nand UO_263 (O_263,N_9962,N_9960);
nand UO_264 (O_264,N_9916,N_9959);
nor UO_265 (O_265,N_9924,N_9989);
or UO_266 (O_266,N_9937,N_9992);
nor UO_267 (O_267,N_9962,N_9977);
or UO_268 (O_268,N_9976,N_9905);
and UO_269 (O_269,N_9992,N_9956);
nor UO_270 (O_270,N_9950,N_9964);
nor UO_271 (O_271,N_9963,N_9948);
nor UO_272 (O_272,N_9991,N_9988);
nand UO_273 (O_273,N_9958,N_9914);
nor UO_274 (O_274,N_9964,N_9995);
or UO_275 (O_275,N_9966,N_9945);
nor UO_276 (O_276,N_9912,N_9990);
nor UO_277 (O_277,N_9995,N_9971);
and UO_278 (O_278,N_9982,N_9935);
or UO_279 (O_279,N_9994,N_9913);
nand UO_280 (O_280,N_9985,N_9920);
or UO_281 (O_281,N_9937,N_9997);
or UO_282 (O_282,N_9966,N_9987);
and UO_283 (O_283,N_9946,N_9991);
and UO_284 (O_284,N_9934,N_9951);
or UO_285 (O_285,N_9961,N_9904);
nor UO_286 (O_286,N_9902,N_9982);
nand UO_287 (O_287,N_9956,N_9993);
and UO_288 (O_288,N_9905,N_9932);
nand UO_289 (O_289,N_9938,N_9942);
or UO_290 (O_290,N_9922,N_9950);
or UO_291 (O_291,N_9917,N_9963);
nand UO_292 (O_292,N_9922,N_9964);
nand UO_293 (O_293,N_9938,N_9950);
nor UO_294 (O_294,N_9975,N_9912);
or UO_295 (O_295,N_9946,N_9961);
nand UO_296 (O_296,N_9975,N_9984);
nor UO_297 (O_297,N_9905,N_9981);
nand UO_298 (O_298,N_9978,N_9955);
or UO_299 (O_299,N_9946,N_9922);
nor UO_300 (O_300,N_9931,N_9966);
and UO_301 (O_301,N_9915,N_9917);
or UO_302 (O_302,N_9966,N_9926);
or UO_303 (O_303,N_9962,N_9964);
xnor UO_304 (O_304,N_9903,N_9940);
nor UO_305 (O_305,N_9993,N_9953);
or UO_306 (O_306,N_9984,N_9951);
or UO_307 (O_307,N_9949,N_9996);
nor UO_308 (O_308,N_9945,N_9954);
and UO_309 (O_309,N_9978,N_9974);
or UO_310 (O_310,N_9962,N_9904);
or UO_311 (O_311,N_9909,N_9984);
nand UO_312 (O_312,N_9913,N_9947);
or UO_313 (O_313,N_9946,N_9921);
or UO_314 (O_314,N_9912,N_9978);
nand UO_315 (O_315,N_9921,N_9979);
nand UO_316 (O_316,N_9970,N_9931);
and UO_317 (O_317,N_9950,N_9934);
nand UO_318 (O_318,N_9971,N_9947);
nor UO_319 (O_319,N_9983,N_9923);
nand UO_320 (O_320,N_9938,N_9927);
and UO_321 (O_321,N_9903,N_9932);
and UO_322 (O_322,N_9973,N_9952);
or UO_323 (O_323,N_9953,N_9958);
and UO_324 (O_324,N_9928,N_9900);
or UO_325 (O_325,N_9996,N_9999);
nor UO_326 (O_326,N_9943,N_9989);
and UO_327 (O_327,N_9937,N_9979);
nand UO_328 (O_328,N_9979,N_9924);
nand UO_329 (O_329,N_9905,N_9961);
and UO_330 (O_330,N_9960,N_9940);
xnor UO_331 (O_331,N_9949,N_9922);
and UO_332 (O_332,N_9979,N_9920);
xnor UO_333 (O_333,N_9952,N_9927);
nand UO_334 (O_334,N_9981,N_9991);
or UO_335 (O_335,N_9953,N_9981);
or UO_336 (O_336,N_9940,N_9994);
nand UO_337 (O_337,N_9974,N_9983);
or UO_338 (O_338,N_9949,N_9982);
and UO_339 (O_339,N_9902,N_9937);
and UO_340 (O_340,N_9905,N_9918);
nand UO_341 (O_341,N_9901,N_9951);
nor UO_342 (O_342,N_9930,N_9958);
nor UO_343 (O_343,N_9993,N_9967);
or UO_344 (O_344,N_9934,N_9986);
and UO_345 (O_345,N_9912,N_9954);
and UO_346 (O_346,N_9925,N_9939);
nor UO_347 (O_347,N_9930,N_9922);
nand UO_348 (O_348,N_9976,N_9907);
nor UO_349 (O_349,N_9924,N_9945);
nand UO_350 (O_350,N_9978,N_9984);
and UO_351 (O_351,N_9916,N_9957);
or UO_352 (O_352,N_9995,N_9937);
and UO_353 (O_353,N_9991,N_9998);
nand UO_354 (O_354,N_9903,N_9986);
or UO_355 (O_355,N_9937,N_9986);
nor UO_356 (O_356,N_9992,N_9997);
nor UO_357 (O_357,N_9996,N_9953);
or UO_358 (O_358,N_9907,N_9942);
nor UO_359 (O_359,N_9986,N_9978);
nand UO_360 (O_360,N_9945,N_9983);
or UO_361 (O_361,N_9988,N_9950);
xor UO_362 (O_362,N_9979,N_9955);
nor UO_363 (O_363,N_9929,N_9984);
and UO_364 (O_364,N_9920,N_9923);
and UO_365 (O_365,N_9935,N_9970);
nand UO_366 (O_366,N_9924,N_9974);
nor UO_367 (O_367,N_9924,N_9949);
and UO_368 (O_368,N_9950,N_9907);
and UO_369 (O_369,N_9989,N_9947);
nor UO_370 (O_370,N_9991,N_9903);
and UO_371 (O_371,N_9990,N_9948);
nor UO_372 (O_372,N_9903,N_9974);
nand UO_373 (O_373,N_9932,N_9992);
or UO_374 (O_374,N_9946,N_9914);
nor UO_375 (O_375,N_9915,N_9907);
and UO_376 (O_376,N_9942,N_9960);
nand UO_377 (O_377,N_9913,N_9950);
and UO_378 (O_378,N_9956,N_9919);
nor UO_379 (O_379,N_9950,N_9930);
or UO_380 (O_380,N_9998,N_9999);
and UO_381 (O_381,N_9998,N_9927);
nand UO_382 (O_382,N_9970,N_9938);
and UO_383 (O_383,N_9995,N_9932);
and UO_384 (O_384,N_9980,N_9953);
or UO_385 (O_385,N_9981,N_9914);
or UO_386 (O_386,N_9908,N_9911);
or UO_387 (O_387,N_9953,N_9948);
nor UO_388 (O_388,N_9914,N_9990);
or UO_389 (O_389,N_9951,N_9961);
nand UO_390 (O_390,N_9976,N_9937);
and UO_391 (O_391,N_9923,N_9940);
nor UO_392 (O_392,N_9902,N_9989);
nor UO_393 (O_393,N_9905,N_9938);
or UO_394 (O_394,N_9917,N_9908);
or UO_395 (O_395,N_9927,N_9920);
nor UO_396 (O_396,N_9983,N_9961);
nand UO_397 (O_397,N_9969,N_9998);
and UO_398 (O_398,N_9974,N_9946);
nor UO_399 (O_399,N_9984,N_9933);
and UO_400 (O_400,N_9996,N_9958);
and UO_401 (O_401,N_9903,N_9947);
or UO_402 (O_402,N_9960,N_9931);
or UO_403 (O_403,N_9991,N_9922);
or UO_404 (O_404,N_9900,N_9965);
nand UO_405 (O_405,N_9911,N_9996);
and UO_406 (O_406,N_9997,N_9988);
nor UO_407 (O_407,N_9918,N_9980);
nand UO_408 (O_408,N_9980,N_9912);
and UO_409 (O_409,N_9925,N_9935);
or UO_410 (O_410,N_9958,N_9962);
nand UO_411 (O_411,N_9907,N_9960);
nor UO_412 (O_412,N_9946,N_9959);
nor UO_413 (O_413,N_9983,N_9959);
and UO_414 (O_414,N_9945,N_9980);
nor UO_415 (O_415,N_9987,N_9955);
nand UO_416 (O_416,N_9941,N_9925);
and UO_417 (O_417,N_9971,N_9916);
nor UO_418 (O_418,N_9974,N_9999);
nor UO_419 (O_419,N_9959,N_9908);
or UO_420 (O_420,N_9976,N_9984);
nand UO_421 (O_421,N_9930,N_9959);
nand UO_422 (O_422,N_9914,N_9966);
and UO_423 (O_423,N_9984,N_9922);
nor UO_424 (O_424,N_9965,N_9995);
and UO_425 (O_425,N_9928,N_9933);
and UO_426 (O_426,N_9937,N_9984);
nand UO_427 (O_427,N_9944,N_9979);
and UO_428 (O_428,N_9968,N_9902);
and UO_429 (O_429,N_9948,N_9900);
nand UO_430 (O_430,N_9933,N_9917);
nor UO_431 (O_431,N_9901,N_9958);
nor UO_432 (O_432,N_9981,N_9916);
and UO_433 (O_433,N_9980,N_9989);
nand UO_434 (O_434,N_9922,N_9989);
or UO_435 (O_435,N_9906,N_9939);
nand UO_436 (O_436,N_9924,N_9952);
nand UO_437 (O_437,N_9999,N_9951);
or UO_438 (O_438,N_9930,N_9910);
nand UO_439 (O_439,N_9976,N_9961);
nor UO_440 (O_440,N_9912,N_9948);
and UO_441 (O_441,N_9928,N_9921);
nand UO_442 (O_442,N_9920,N_9934);
or UO_443 (O_443,N_9997,N_9906);
nand UO_444 (O_444,N_9912,N_9972);
xnor UO_445 (O_445,N_9996,N_9940);
and UO_446 (O_446,N_9997,N_9965);
nor UO_447 (O_447,N_9975,N_9954);
or UO_448 (O_448,N_9942,N_9965);
or UO_449 (O_449,N_9950,N_9955);
nor UO_450 (O_450,N_9914,N_9933);
and UO_451 (O_451,N_9960,N_9970);
or UO_452 (O_452,N_9958,N_9969);
nor UO_453 (O_453,N_9908,N_9902);
nor UO_454 (O_454,N_9969,N_9957);
nand UO_455 (O_455,N_9968,N_9931);
nand UO_456 (O_456,N_9999,N_9927);
and UO_457 (O_457,N_9976,N_9903);
and UO_458 (O_458,N_9957,N_9996);
or UO_459 (O_459,N_9981,N_9908);
or UO_460 (O_460,N_9984,N_9974);
nand UO_461 (O_461,N_9905,N_9935);
or UO_462 (O_462,N_9987,N_9969);
nor UO_463 (O_463,N_9985,N_9926);
and UO_464 (O_464,N_9974,N_9930);
or UO_465 (O_465,N_9919,N_9901);
or UO_466 (O_466,N_9917,N_9983);
nand UO_467 (O_467,N_9921,N_9910);
and UO_468 (O_468,N_9919,N_9934);
nor UO_469 (O_469,N_9964,N_9989);
nor UO_470 (O_470,N_9983,N_9916);
or UO_471 (O_471,N_9906,N_9965);
nand UO_472 (O_472,N_9996,N_9988);
nor UO_473 (O_473,N_9913,N_9940);
nor UO_474 (O_474,N_9905,N_9967);
and UO_475 (O_475,N_9999,N_9959);
and UO_476 (O_476,N_9932,N_9943);
nor UO_477 (O_477,N_9976,N_9927);
and UO_478 (O_478,N_9996,N_9997);
or UO_479 (O_479,N_9931,N_9919);
nor UO_480 (O_480,N_9903,N_9981);
or UO_481 (O_481,N_9919,N_9976);
and UO_482 (O_482,N_9950,N_9940);
nor UO_483 (O_483,N_9959,N_9932);
nor UO_484 (O_484,N_9918,N_9931);
or UO_485 (O_485,N_9958,N_9906);
and UO_486 (O_486,N_9960,N_9947);
or UO_487 (O_487,N_9961,N_9955);
or UO_488 (O_488,N_9969,N_9936);
nand UO_489 (O_489,N_9969,N_9963);
or UO_490 (O_490,N_9974,N_9919);
nor UO_491 (O_491,N_9978,N_9909);
nor UO_492 (O_492,N_9975,N_9948);
and UO_493 (O_493,N_9934,N_9985);
or UO_494 (O_494,N_9931,N_9990);
or UO_495 (O_495,N_9948,N_9943);
nor UO_496 (O_496,N_9930,N_9934);
and UO_497 (O_497,N_9976,N_9988);
xnor UO_498 (O_498,N_9926,N_9961);
nor UO_499 (O_499,N_9932,N_9963);
and UO_500 (O_500,N_9947,N_9955);
nor UO_501 (O_501,N_9925,N_9950);
xnor UO_502 (O_502,N_9907,N_9988);
nand UO_503 (O_503,N_9990,N_9910);
or UO_504 (O_504,N_9950,N_9987);
nor UO_505 (O_505,N_9901,N_9923);
nand UO_506 (O_506,N_9910,N_9999);
nor UO_507 (O_507,N_9964,N_9960);
nand UO_508 (O_508,N_9999,N_9923);
nand UO_509 (O_509,N_9951,N_9990);
nand UO_510 (O_510,N_9930,N_9931);
or UO_511 (O_511,N_9935,N_9934);
and UO_512 (O_512,N_9970,N_9944);
xnor UO_513 (O_513,N_9962,N_9952);
nor UO_514 (O_514,N_9986,N_9925);
nand UO_515 (O_515,N_9930,N_9954);
or UO_516 (O_516,N_9978,N_9901);
nand UO_517 (O_517,N_9928,N_9920);
nand UO_518 (O_518,N_9942,N_9905);
nor UO_519 (O_519,N_9936,N_9998);
and UO_520 (O_520,N_9923,N_9914);
or UO_521 (O_521,N_9987,N_9937);
or UO_522 (O_522,N_9925,N_9988);
and UO_523 (O_523,N_9981,N_9979);
or UO_524 (O_524,N_9931,N_9952);
or UO_525 (O_525,N_9920,N_9930);
nor UO_526 (O_526,N_9963,N_9983);
nor UO_527 (O_527,N_9957,N_9947);
and UO_528 (O_528,N_9967,N_9930);
or UO_529 (O_529,N_9943,N_9907);
or UO_530 (O_530,N_9988,N_9955);
and UO_531 (O_531,N_9906,N_9957);
nand UO_532 (O_532,N_9901,N_9960);
and UO_533 (O_533,N_9996,N_9912);
and UO_534 (O_534,N_9977,N_9938);
and UO_535 (O_535,N_9997,N_9905);
or UO_536 (O_536,N_9931,N_9948);
nor UO_537 (O_537,N_9972,N_9930);
or UO_538 (O_538,N_9963,N_9968);
or UO_539 (O_539,N_9949,N_9910);
nand UO_540 (O_540,N_9997,N_9933);
or UO_541 (O_541,N_9973,N_9999);
or UO_542 (O_542,N_9966,N_9906);
and UO_543 (O_543,N_9901,N_9953);
and UO_544 (O_544,N_9953,N_9982);
nor UO_545 (O_545,N_9977,N_9931);
nor UO_546 (O_546,N_9941,N_9906);
nand UO_547 (O_547,N_9942,N_9994);
and UO_548 (O_548,N_9984,N_9967);
nand UO_549 (O_549,N_9923,N_9998);
and UO_550 (O_550,N_9911,N_9971);
and UO_551 (O_551,N_9947,N_9952);
and UO_552 (O_552,N_9912,N_9963);
and UO_553 (O_553,N_9993,N_9966);
xnor UO_554 (O_554,N_9998,N_9920);
nor UO_555 (O_555,N_9990,N_9963);
or UO_556 (O_556,N_9995,N_9901);
nor UO_557 (O_557,N_9938,N_9963);
nand UO_558 (O_558,N_9907,N_9933);
nor UO_559 (O_559,N_9906,N_9944);
nor UO_560 (O_560,N_9992,N_9928);
nor UO_561 (O_561,N_9952,N_9907);
nand UO_562 (O_562,N_9961,N_9953);
nor UO_563 (O_563,N_9909,N_9997);
nand UO_564 (O_564,N_9985,N_9987);
nand UO_565 (O_565,N_9914,N_9996);
or UO_566 (O_566,N_9920,N_9909);
nor UO_567 (O_567,N_9967,N_9951);
and UO_568 (O_568,N_9986,N_9996);
or UO_569 (O_569,N_9961,N_9921);
and UO_570 (O_570,N_9935,N_9900);
and UO_571 (O_571,N_9948,N_9906);
and UO_572 (O_572,N_9906,N_9978);
and UO_573 (O_573,N_9960,N_9936);
nand UO_574 (O_574,N_9933,N_9906);
nor UO_575 (O_575,N_9958,N_9981);
nand UO_576 (O_576,N_9992,N_9925);
nand UO_577 (O_577,N_9979,N_9910);
or UO_578 (O_578,N_9935,N_9941);
and UO_579 (O_579,N_9932,N_9906);
and UO_580 (O_580,N_9968,N_9906);
nand UO_581 (O_581,N_9996,N_9907);
nand UO_582 (O_582,N_9965,N_9939);
and UO_583 (O_583,N_9942,N_9919);
and UO_584 (O_584,N_9944,N_9926);
nor UO_585 (O_585,N_9974,N_9969);
nand UO_586 (O_586,N_9948,N_9921);
and UO_587 (O_587,N_9988,N_9951);
or UO_588 (O_588,N_9972,N_9934);
nor UO_589 (O_589,N_9902,N_9972);
nor UO_590 (O_590,N_9982,N_9942);
or UO_591 (O_591,N_9984,N_9982);
and UO_592 (O_592,N_9902,N_9951);
or UO_593 (O_593,N_9931,N_9981);
or UO_594 (O_594,N_9937,N_9959);
nor UO_595 (O_595,N_9974,N_9912);
or UO_596 (O_596,N_9950,N_9978);
or UO_597 (O_597,N_9915,N_9941);
or UO_598 (O_598,N_9998,N_9975);
and UO_599 (O_599,N_9941,N_9930);
nand UO_600 (O_600,N_9986,N_9948);
xor UO_601 (O_601,N_9929,N_9958);
nand UO_602 (O_602,N_9919,N_9994);
nand UO_603 (O_603,N_9947,N_9999);
and UO_604 (O_604,N_9971,N_9987);
xnor UO_605 (O_605,N_9996,N_9966);
or UO_606 (O_606,N_9967,N_9920);
or UO_607 (O_607,N_9996,N_9918);
or UO_608 (O_608,N_9918,N_9920);
nand UO_609 (O_609,N_9977,N_9967);
or UO_610 (O_610,N_9926,N_9928);
xnor UO_611 (O_611,N_9986,N_9988);
and UO_612 (O_612,N_9966,N_9973);
xor UO_613 (O_613,N_9933,N_9970);
and UO_614 (O_614,N_9937,N_9940);
or UO_615 (O_615,N_9955,N_9954);
or UO_616 (O_616,N_9999,N_9906);
nand UO_617 (O_617,N_9916,N_9988);
nand UO_618 (O_618,N_9994,N_9959);
and UO_619 (O_619,N_9948,N_9903);
and UO_620 (O_620,N_9945,N_9979);
or UO_621 (O_621,N_9941,N_9951);
nor UO_622 (O_622,N_9957,N_9951);
nand UO_623 (O_623,N_9985,N_9998);
and UO_624 (O_624,N_9915,N_9934);
nand UO_625 (O_625,N_9903,N_9925);
and UO_626 (O_626,N_9973,N_9982);
nand UO_627 (O_627,N_9956,N_9954);
or UO_628 (O_628,N_9942,N_9906);
or UO_629 (O_629,N_9924,N_9966);
nand UO_630 (O_630,N_9960,N_9966);
nand UO_631 (O_631,N_9944,N_9936);
nand UO_632 (O_632,N_9909,N_9962);
or UO_633 (O_633,N_9915,N_9942);
and UO_634 (O_634,N_9911,N_9912);
or UO_635 (O_635,N_9974,N_9936);
nand UO_636 (O_636,N_9956,N_9939);
and UO_637 (O_637,N_9990,N_9902);
nand UO_638 (O_638,N_9917,N_9988);
or UO_639 (O_639,N_9942,N_9976);
nor UO_640 (O_640,N_9991,N_9935);
and UO_641 (O_641,N_9975,N_9987);
nor UO_642 (O_642,N_9989,N_9954);
xor UO_643 (O_643,N_9995,N_9936);
or UO_644 (O_644,N_9952,N_9988);
nand UO_645 (O_645,N_9916,N_9950);
nand UO_646 (O_646,N_9904,N_9948);
and UO_647 (O_647,N_9906,N_9961);
or UO_648 (O_648,N_9957,N_9970);
or UO_649 (O_649,N_9906,N_9903);
nor UO_650 (O_650,N_9999,N_9942);
or UO_651 (O_651,N_9946,N_9989);
and UO_652 (O_652,N_9983,N_9938);
or UO_653 (O_653,N_9982,N_9909);
nor UO_654 (O_654,N_9948,N_9939);
xor UO_655 (O_655,N_9923,N_9971);
or UO_656 (O_656,N_9971,N_9985);
and UO_657 (O_657,N_9942,N_9921);
and UO_658 (O_658,N_9914,N_9955);
nor UO_659 (O_659,N_9961,N_9900);
nand UO_660 (O_660,N_9904,N_9905);
and UO_661 (O_661,N_9953,N_9926);
nor UO_662 (O_662,N_9992,N_9926);
nand UO_663 (O_663,N_9967,N_9983);
nand UO_664 (O_664,N_9968,N_9908);
nand UO_665 (O_665,N_9941,N_9965);
or UO_666 (O_666,N_9915,N_9965);
nand UO_667 (O_667,N_9988,N_9903);
and UO_668 (O_668,N_9936,N_9989);
nand UO_669 (O_669,N_9943,N_9975);
and UO_670 (O_670,N_9904,N_9981);
or UO_671 (O_671,N_9924,N_9968);
and UO_672 (O_672,N_9964,N_9937);
nor UO_673 (O_673,N_9963,N_9964);
nor UO_674 (O_674,N_9916,N_9926);
or UO_675 (O_675,N_9935,N_9998);
and UO_676 (O_676,N_9979,N_9938);
or UO_677 (O_677,N_9907,N_9997);
and UO_678 (O_678,N_9984,N_9915);
nor UO_679 (O_679,N_9939,N_9915);
and UO_680 (O_680,N_9969,N_9900);
nor UO_681 (O_681,N_9926,N_9990);
or UO_682 (O_682,N_9900,N_9999);
nor UO_683 (O_683,N_9924,N_9959);
nand UO_684 (O_684,N_9974,N_9949);
nand UO_685 (O_685,N_9949,N_9932);
or UO_686 (O_686,N_9952,N_9972);
nor UO_687 (O_687,N_9951,N_9962);
nor UO_688 (O_688,N_9951,N_9963);
and UO_689 (O_689,N_9948,N_9997);
nor UO_690 (O_690,N_9976,N_9999);
nor UO_691 (O_691,N_9912,N_9929);
or UO_692 (O_692,N_9913,N_9930);
nand UO_693 (O_693,N_9954,N_9919);
nor UO_694 (O_694,N_9919,N_9917);
or UO_695 (O_695,N_9968,N_9909);
nor UO_696 (O_696,N_9999,N_9912);
nand UO_697 (O_697,N_9920,N_9987);
and UO_698 (O_698,N_9965,N_9908);
and UO_699 (O_699,N_9914,N_9969);
and UO_700 (O_700,N_9912,N_9983);
and UO_701 (O_701,N_9993,N_9980);
nand UO_702 (O_702,N_9901,N_9947);
and UO_703 (O_703,N_9941,N_9964);
and UO_704 (O_704,N_9948,N_9956);
or UO_705 (O_705,N_9907,N_9948);
or UO_706 (O_706,N_9994,N_9918);
nand UO_707 (O_707,N_9922,N_9993);
nand UO_708 (O_708,N_9929,N_9945);
nand UO_709 (O_709,N_9936,N_9949);
or UO_710 (O_710,N_9909,N_9922);
nor UO_711 (O_711,N_9931,N_9924);
nor UO_712 (O_712,N_9927,N_9974);
nor UO_713 (O_713,N_9992,N_9948);
nand UO_714 (O_714,N_9982,N_9906);
nor UO_715 (O_715,N_9964,N_9954);
and UO_716 (O_716,N_9963,N_9940);
and UO_717 (O_717,N_9914,N_9900);
nand UO_718 (O_718,N_9927,N_9932);
and UO_719 (O_719,N_9996,N_9977);
or UO_720 (O_720,N_9902,N_9958);
and UO_721 (O_721,N_9970,N_9956);
xor UO_722 (O_722,N_9966,N_9907);
nand UO_723 (O_723,N_9958,N_9932);
nand UO_724 (O_724,N_9928,N_9946);
or UO_725 (O_725,N_9950,N_9975);
and UO_726 (O_726,N_9917,N_9927);
or UO_727 (O_727,N_9975,N_9938);
nor UO_728 (O_728,N_9993,N_9982);
nand UO_729 (O_729,N_9937,N_9915);
or UO_730 (O_730,N_9946,N_9942);
and UO_731 (O_731,N_9987,N_9900);
nand UO_732 (O_732,N_9913,N_9927);
nor UO_733 (O_733,N_9972,N_9983);
nor UO_734 (O_734,N_9906,N_9953);
nor UO_735 (O_735,N_9923,N_9989);
nor UO_736 (O_736,N_9908,N_9920);
and UO_737 (O_737,N_9916,N_9943);
nor UO_738 (O_738,N_9972,N_9981);
and UO_739 (O_739,N_9991,N_9961);
or UO_740 (O_740,N_9963,N_9982);
and UO_741 (O_741,N_9937,N_9921);
nand UO_742 (O_742,N_9990,N_9920);
and UO_743 (O_743,N_9943,N_9959);
and UO_744 (O_744,N_9994,N_9960);
and UO_745 (O_745,N_9918,N_9936);
or UO_746 (O_746,N_9936,N_9900);
nor UO_747 (O_747,N_9971,N_9935);
nor UO_748 (O_748,N_9955,N_9966);
and UO_749 (O_749,N_9972,N_9999);
and UO_750 (O_750,N_9917,N_9907);
nand UO_751 (O_751,N_9946,N_9977);
nand UO_752 (O_752,N_9904,N_9992);
nor UO_753 (O_753,N_9999,N_9908);
nor UO_754 (O_754,N_9998,N_9914);
and UO_755 (O_755,N_9918,N_9902);
nand UO_756 (O_756,N_9990,N_9986);
or UO_757 (O_757,N_9927,N_9928);
nor UO_758 (O_758,N_9978,N_9932);
nor UO_759 (O_759,N_9975,N_9924);
or UO_760 (O_760,N_9971,N_9994);
nand UO_761 (O_761,N_9950,N_9928);
nor UO_762 (O_762,N_9923,N_9964);
xor UO_763 (O_763,N_9917,N_9973);
or UO_764 (O_764,N_9947,N_9987);
nor UO_765 (O_765,N_9949,N_9923);
nor UO_766 (O_766,N_9933,N_9998);
and UO_767 (O_767,N_9949,N_9921);
and UO_768 (O_768,N_9960,N_9993);
nand UO_769 (O_769,N_9988,N_9928);
nand UO_770 (O_770,N_9994,N_9908);
nand UO_771 (O_771,N_9947,N_9980);
nor UO_772 (O_772,N_9975,N_9914);
nor UO_773 (O_773,N_9917,N_9964);
nor UO_774 (O_774,N_9989,N_9987);
and UO_775 (O_775,N_9923,N_9912);
or UO_776 (O_776,N_9999,N_9933);
and UO_777 (O_777,N_9924,N_9929);
nor UO_778 (O_778,N_9914,N_9936);
and UO_779 (O_779,N_9993,N_9936);
and UO_780 (O_780,N_9930,N_9955);
nand UO_781 (O_781,N_9965,N_9977);
and UO_782 (O_782,N_9990,N_9938);
or UO_783 (O_783,N_9942,N_9939);
and UO_784 (O_784,N_9976,N_9979);
or UO_785 (O_785,N_9911,N_9934);
and UO_786 (O_786,N_9975,N_9901);
or UO_787 (O_787,N_9958,N_9944);
nor UO_788 (O_788,N_9900,N_9956);
or UO_789 (O_789,N_9950,N_9996);
and UO_790 (O_790,N_9942,N_9961);
and UO_791 (O_791,N_9949,N_9961);
or UO_792 (O_792,N_9976,N_9948);
nor UO_793 (O_793,N_9977,N_9952);
nor UO_794 (O_794,N_9944,N_9950);
or UO_795 (O_795,N_9977,N_9936);
and UO_796 (O_796,N_9958,N_9966);
nand UO_797 (O_797,N_9923,N_9970);
and UO_798 (O_798,N_9907,N_9909);
and UO_799 (O_799,N_9986,N_9921);
and UO_800 (O_800,N_9926,N_9931);
or UO_801 (O_801,N_9983,N_9958);
nand UO_802 (O_802,N_9995,N_9975);
nor UO_803 (O_803,N_9973,N_9925);
and UO_804 (O_804,N_9978,N_9951);
or UO_805 (O_805,N_9979,N_9970);
and UO_806 (O_806,N_9952,N_9984);
and UO_807 (O_807,N_9906,N_9967);
or UO_808 (O_808,N_9932,N_9922);
nor UO_809 (O_809,N_9949,N_9957);
nor UO_810 (O_810,N_9922,N_9912);
xor UO_811 (O_811,N_9971,N_9953);
or UO_812 (O_812,N_9992,N_9920);
nand UO_813 (O_813,N_9920,N_9915);
nor UO_814 (O_814,N_9993,N_9983);
or UO_815 (O_815,N_9954,N_9952);
or UO_816 (O_816,N_9997,N_9985);
or UO_817 (O_817,N_9916,N_9979);
or UO_818 (O_818,N_9940,N_9992);
nand UO_819 (O_819,N_9952,N_9902);
or UO_820 (O_820,N_9928,N_9918);
or UO_821 (O_821,N_9918,N_9969);
and UO_822 (O_822,N_9929,N_9910);
nor UO_823 (O_823,N_9977,N_9995);
and UO_824 (O_824,N_9992,N_9902);
and UO_825 (O_825,N_9932,N_9920);
and UO_826 (O_826,N_9999,N_9925);
or UO_827 (O_827,N_9965,N_9969);
and UO_828 (O_828,N_9993,N_9933);
nand UO_829 (O_829,N_9985,N_9910);
or UO_830 (O_830,N_9914,N_9983);
nand UO_831 (O_831,N_9919,N_9986);
nand UO_832 (O_832,N_9915,N_9959);
and UO_833 (O_833,N_9969,N_9972);
or UO_834 (O_834,N_9900,N_9912);
nor UO_835 (O_835,N_9903,N_9936);
nor UO_836 (O_836,N_9945,N_9982);
nand UO_837 (O_837,N_9933,N_9964);
nor UO_838 (O_838,N_9924,N_9913);
nand UO_839 (O_839,N_9930,N_9936);
or UO_840 (O_840,N_9957,N_9928);
nand UO_841 (O_841,N_9999,N_9970);
nand UO_842 (O_842,N_9940,N_9945);
or UO_843 (O_843,N_9908,N_9935);
nor UO_844 (O_844,N_9900,N_9971);
and UO_845 (O_845,N_9970,N_9922);
nor UO_846 (O_846,N_9956,N_9958);
xnor UO_847 (O_847,N_9987,N_9934);
or UO_848 (O_848,N_9983,N_9941);
and UO_849 (O_849,N_9926,N_9920);
nand UO_850 (O_850,N_9949,N_9919);
nor UO_851 (O_851,N_9997,N_9976);
or UO_852 (O_852,N_9913,N_9980);
and UO_853 (O_853,N_9905,N_9954);
nand UO_854 (O_854,N_9904,N_9913);
nor UO_855 (O_855,N_9990,N_9937);
nor UO_856 (O_856,N_9977,N_9982);
nor UO_857 (O_857,N_9979,N_9936);
xnor UO_858 (O_858,N_9998,N_9921);
nor UO_859 (O_859,N_9959,N_9958);
or UO_860 (O_860,N_9955,N_9938);
nand UO_861 (O_861,N_9973,N_9941);
nor UO_862 (O_862,N_9938,N_9936);
and UO_863 (O_863,N_9994,N_9979);
nand UO_864 (O_864,N_9956,N_9950);
and UO_865 (O_865,N_9995,N_9939);
and UO_866 (O_866,N_9983,N_9979);
nand UO_867 (O_867,N_9927,N_9903);
and UO_868 (O_868,N_9981,N_9992);
or UO_869 (O_869,N_9999,N_9919);
or UO_870 (O_870,N_9957,N_9903);
nor UO_871 (O_871,N_9999,N_9983);
or UO_872 (O_872,N_9930,N_9933);
or UO_873 (O_873,N_9905,N_9915);
nand UO_874 (O_874,N_9953,N_9923);
nor UO_875 (O_875,N_9908,N_9988);
nand UO_876 (O_876,N_9932,N_9950);
nor UO_877 (O_877,N_9916,N_9942);
nor UO_878 (O_878,N_9924,N_9958);
or UO_879 (O_879,N_9961,N_9915);
or UO_880 (O_880,N_9966,N_9948);
nand UO_881 (O_881,N_9969,N_9909);
or UO_882 (O_882,N_9966,N_9961);
or UO_883 (O_883,N_9982,N_9981);
nand UO_884 (O_884,N_9991,N_9943);
nor UO_885 (O_885,N_9948,N_9959);
nor UO_886 (O_886,N_9949,N_9911);
nand UO_887 (O_887,N_9911,N_9988);
xor UO_888 (O_888,N_9980,N_9962);
nor UO_889 (O_889,N_9983,N_9946);
xor UO_890 (O_890,N_9951,N_9904);
nor UO_891 (O_891,N_9909,N_9990);
nor UO_892 (O_892,N_9974,N_9975);
nor UO_893 (O_893,N_9904,N_9974);
and UO_894 (O_894,N_9937,N_9973);
or UO_895 (O_895,N_9928,N_9982);
nand UO_896 (O_896,N_9963,N_9941);
nor UO_897 (O_897,N_9980,N_9984);
nor UO_898 (O_898,N_9956,N_9999);
nand UO_899 (O_899,N_9967,N_9970);
nand UO_900 (O_900,N_9960,N_9930);
nand UO_901 (O_901,N_9921,N_9925);
and UO_902 (O_902,N_9901,N_9906);
and UO_903 (O_903,N_9990,N_9985);
nand UO_904 (O_904,N_9986,N_9920);
nand UO_905 (O_905,N_9909,N_9936);
nand UO_906 (O_906,N_9935,N_9919);
or UO_907 (O_907,N_9978,N_9993);
or UO_908 (O_908,N_9914,N_9929);
or UO_909 (O_909,N_9915,N_9930);
and UO_910 (O_910,N_9976,N_9952);
or UO_911 (O_911,N_9938,N_9915);
or UO_912 (O_912,N_9916,N_9985);
nor UO_913 (O_913,N_9944,N_9977);
and UO_914 (O_914,N_9949,N_9994);
nor UO_915 (O_915,N_9933,N_9958);
and UO_916 (O_916,N_9996,N_9973);
nor UO_917 (O_917,N_9993,N_9977);
or UO_918 (O_918,N_9908,N_9962);
and UO_919 (O_919,N_9929,N_9920);
nor UO_920 (O_920,N_9941,N_9926);
nor UO_921 (O_921,N_9931,N_9917);
and UO_922 (O_922,N_9951,N_9972);
or UO_923 (O_923,N_9920,N_9901);
and UO_924 (O_924,N_9958,N_9965);
or UO_925 (O_925,N_9936,N_9965);
nor UO_926 (O_926,N_9943,N_9927);
or UO_927 (O_927,N_9969,N_9959);
or UO_928 (O_928,N_9964,N_9935);
nand UO_929 (O_929,N_9911,N_9981);
and UO_930 (O_930,N_9916,N_9949);
or UO_931 (O_931,N_9985,N_9970);
nand UO_932 (O_932,N_9977,N_9959);
or UO_933 (O_933,N_9966,N_9994);
or UO_934 (O_934,N_9918,N_9950);
or UO_935 (O_935,N_9918,N_9971);
nand UO_936 (O_936,N_9914,N_9915);
and UO_937 (O_937,N_9919,N_9958);
or UO_938 (O_938,N_9937,N_9963);
xnor UO_939 (O_939,N_9974,N_9943);
nor UO_940 (O_940,N_9992,N_9978);
nor UO_941 (O_941,N_9958,N_9997);
and UO_942 (O_942,N_9962,N_9979);
nand UO_943 (O_943,N_9979,N_9987);
or UO_944 (O_944,N_9931,N_9943);
nand UO_945 (O_945,N_9935,N_9977);
nor UO_946 (O_946,N_9984,N_9968);
or UO_947 (O_947,N_9966,N_9923);
or UO_948 (O_948,N_9937,N_9974);
and UO_949 (O_949,N_9960,N_9967);
nor UO_950 (O_950,N_9972,N_9913);
nor UO_951 (O_951,N_9919,N_9977);
and UO_952 (O_952,N_9954,N_9939);
nor UO_953 (O_953,N_9946,N_9958);
or UO_954 (O_954,N_9922,N_9923);
and UO_955 (O_955,N_9991,N_9983);
xnor UO_956 (O_956,N_9969,N_9943);
nor UO_957 (O_957,N_9971,N_9952);
or UO_958 (O_958,N_9965,N_9949);
nand UO_959 (O_959,N_9963,N_9974);
or UO_960 (O_960,N_9989,N_9900);
and UO_961 (O_961,N_9956,N_9951);
and UO_962 (O_962,N_9978,N_9969);
or UO_963 (O_963,N_9906,N_9981);
and UO_964 (O_964,N_9952,N_9978);
nand UO_965 (O_965,N_9906,N_9980);
nand UO_966 (O_966,N_9993,N_9949);
nor UO_967 (O_967,N_9997,N_9940);
nor UO_968 (O_968,N_9978,N_9914);
or UO_969 (O_969,N_9971,N_9976);
nor UO_970 (O_970,N_9910,N_9952);
or UO_971 (O_971,N_9964,N_9952);
nor UO_972 (O_972,N_9931,N_9940);
nor UO_973 (O_973,N_9945,N_9994);
nor UO_974 (O_974,N_9942,N_9926);
nor UO_975 (O_975,N_9978,N_9975);
and UO_976 (O_976,N_9929,N_9904);
or UO_977 (O_977,N_9970,N_9993);
nand UO_978 (O_978,N_9993,N_9958);
and UO_979 (O_979,N_9999,N_9944);
or UO_980 (O_980,N_9985,N_9979);
or UO_981 (O_981,N_9915,N_9928);
or UO_982 (O_982,N_9935,N_9957);
nand UO_983 (O_983,N_9990,N_9998);
nand UO_984 (O_984,N_9950,N_9936);
or UO_985 (O_985,N_9925,N_9963);
or UO_986 (O_986,N_9910,N_9974);
nand UO_987 (O_987,N_9980,N_9909);
and UO_988 (O_988,N_9982,N_9908);
or UO_989 (O_989,N_9968,N_9966);
and UO_990 (O_990,N_9986,N_9997);
or UO_991 (O_991,N_9957,N_9980);
nor UO_992 (O_992,N_9916,N_9990);
xor UO_993 (O_993,N_9989,N_9920);
nor UO_994 (O_994,N_9939,N_9978);
nor UO_995 (O_995,N_9993,N_9943);
nand UO_996 (O_996,N_9999,N_9975);
nor UO_997 (O_997,N_9944,N_9925);
nand UO_998 (O_998,N_9946,N_9999);
nor UO_999 (O_999,N_9951,N_9936);
xnor UO_1000 (O_1000,N_9973,N_9904);
and UO_1001 (O_1001,N_9987,N_9923);
and UO_1002 (O_1002,N_9938,N_9954);
or UO_1003 (O_1003,N_9953,N_9991);
nor UO_1004 (O_1004,N_9933,N_9915);
nor UO_1005 (O_1005,N_9988,N_9946);
nor UO_1006 (O_1006,N_9913,N_9935);
and UO_1007 (O_1007,N_9924,N_9962);
nand UO_1008 (O_1008,N_9960,N_9983);
and UO_1009 (O_1009,N_9922,N_9990);
and UO_1010 (O_1010,N_9944,N_9915);
or UO_1011 (O_1011,N_9991,N_9979);
xnor UO_1012 (O_1012,N_9901,N_9979);
nor UO_1013 (O_1013,N_9947,N_9939);
nand UO_1014 (O_1014,N_9964,N_9976);
nor UO_1015 (O_1015,N_9970,N_9954);
xor UO_1016 (O_1016,N_9910,N_9911);
or UO_1017 (O_1017,N_9957,N_9967);
or UO_1018 (O_1018,N_9913,N_9929);
nor UO_1019 (O_1019,N_9965,N_9954);
and UO_1020 (O_1020,N_9946,N_9982);
nor UO_1021 (O_1021,N_9949,N_9901);
or UO_1022 (O_1022,N_9994,N_9921);
nor UO_1023 (O_1023,N_9945,N_9975);
and UO_1024 (O_1024,N_9933,N_9972);
or UO_1025 (O_1025,N_9997,N_9950);
or UO_1026 (O_1026,N_9918,N_9915);
or UO_1027 (O_1027,N_9953,N_9932);
and UO_1028 (O_1028,N_9902,N_9905);
nor UO_1029 (O_1029,N_9980,N_9931);
nor UO_1030 (O_1030,N_9931,N_9949);
nand UO_1031 (O_1031,N_9927,N_9960);
nor UO_1032 (O_1032,N_9968,N_9911);
nand UO_1033 (O_1033,N_9931,N_9944);
or UO_1034 (O_1034,N_9960,N_9913);
and UO_1035 (O_1035,N_9917,N_9989);
nand UO_1036 (O_1036,N_9961,N_9902);
nor UO_1037 (O_1037,N_9956,N_9937);
and UO_1038 (O_1038,N_9931,N_9923);
nand UO_1039 (O_1039,N_9934,N_9989);
nor UO_1040 (O_1040,N_9961,N_9963);
xnor UO_1041 (O_1041,N_9957,N_9929);
or UO_1042 (O_1042,N_9957,N_9919);
nand UO_1043 (O_1043,N_9939,N_9920);
or UO_1044 (O_1044,N_9986,N_9935);
nand UO_1045 (O_1045,N_9940,N_9956);
nor UO_1046 (O_1046,N_9929,N_9956);
xnor UO_1047 (O_1047,N_9984,N_9964);
nand UO_1048 (O_1048,N_9926,N_9910);
nand UO_1049 (O_1049,N_9958,N_9989);
nor UO_1050 (O_1050,N_9933,N_9968);
and UO_1051 (O_1051,N_9939,N_9982);
and UO_1052 (O_1052,N_9994,N_9925);
nand UO_1053 (O_1053,N_9943,N_9970);
nor UO_1054 (O_1054,N_9973,N_9927);
nor UO_1055 (O_1055,N_9990,N_9903);
or UO_1056 (O_1056,N_9971,N_9910);
xnor UO_1057 (O_1057,N_9911,N_9921);
and UO_1058 (O_1058,N_9981,N_9989);
nand UO_1059 (O_1059,N_9960,N_9919);
nand UO_1060 (O_1060,N_9917,N_9993);
xnor UO_1061 (O_1061,N_9937,N_9955);
or UO_1062 (O_1062,N_9940,N_9964);
nand UO_1063 (O_1063,N_9904,N_9940);
nand UO_1064 (O_1064,N_9965,N_9910);
and UO_1065 (O_1065,N_9957,N_9905);
nand UO_1066 (O_1066,N_9971,N_9950);
nor UO_1067 (O_1067,N_9920,N_9968);
nand UO_1068 (O_1068,N_9906,N_9904);
and UO_1069 (O_1069,N_9964,N_9985);
and UO_1070 (O_1070,N_9980,N_9968);
and UO_1071 (O_1071,N_9954,N_9902);
nand UO_1072 (O_1072,N_9930,N_9987);
nor UO_1073 (O_1073,N_9984,N_9983);
xor UO_1074 (O_1074,N_9916,N_9932);
nor UO_1075 (O_1075,N_9979,N_9935);
nand UO_1076 (O_1076,N_9945,N_9926);
nor UO_1077 (O_1077,N_9973,N_9939);
or UO_1078 (O_1078,N_9908,N_9950);
nor UO_1079 (O_1079,N_9967,N_9978);
or UO_1080 (O_1080,N_9990,N_9992);
nor UO_1081 (O_1081,N_9972,N_9971);
nor UO_1082 (O_1082,N_9971,N_9945);
or UO_1083 (O_1083,N_9929,N_9934);
nor UO_1084 (O_1084,N_9960,N_9912);
or UO_1085 (O_1085,N_9920,N_9937);
and UO_1086 (O_1086,N_9982,N_9997);
or UO_1087 (O_1087,N_9919,N_9937);
nor UO_1088 (O_1088,N_9999,N_9931);
nor UO_1089 (O_1089,N_9913,N_9973);
xor UO_1090 (O_1090,N_9911,N_9955);
or UO_1091 (O_1091,N_9958,N_9982);
and UO_1092 (O_1092,N_9964,N_9903);
nor UO_1093 (O_1093,N_9931,N_9941);
nor UO_1094 (O_1094,N_9926,N_9922);
nand UO_1095 (O_1095,N_9951,N_9968);
or UO_1096 (O_1096,N_9957,N_9972);
nor UO_1097 (O_1097,N_9918,N_9979);
and UO_1098 (O_1098,N_9956,N_9971);
nand UO_1099 (O_1099,N_9947,N_9916);
or UO_1100 (O_1100,N_9948,N_9941);
nor UO_1101 (O_1101,N_9918,N_9937);
nand UO_1102 (O_1102,N_9988,N_9924);
and UO_1103 (O_1103,N_9932,N_9979);
nor UO_1104 (O_1104,N_9984,N_9997);
nand UO_1105 (O_1105,N_9988,N_9977);
and UO_1106 (O_1106,N_9941,N_9916);
and UO_1107 (O_1107,N_9927,N_9911);
nand UO_1108 (O_1108,N_9913,N_9990);
or UO_1109 (O_1109,N_9920,N_9917);
nor UO_1110 (O_1110,N_9956,N_9968);
and UO_1111 (O_1111,N_9992,N_9908);
nand UO_1112 (O_1112,N_9918,N_9983);
or UO_1113 (O_1113,N_9982,N_9966);
nand UO_1114 (O_1114,N_9969,N_9994);
nand UO_1115 (O_1115,N_9978,N_9917);
nand UO_1116 (O_1116,N_9993,N_9923);
nor UO_1117 (O_1117,N_9933,N_9957);
or UO_1118 (O_1118,N_9989,N_9945);
or UO_1119 (O_1119,N_9914,N_9971);
or UO_1120 (O_1120,N_9920,N_9912);
nand UO_1121 (O_1121,N_9930,N_9980);
nand UO_1122 (O_1122,N_9958,N_9951);
or UO_1123 (O_1123,N_9972,N_9931);
or UO_1124 (O_1124,N_9961,N_9937);
nor UO_1125 (O_1125,N_9936,N_9970);
or UO_1126 (O_1126,N_9906,N_9971);
and UO_1127 (O_1127,N_9939,N_9958);
and UO_1128 (O_1128,N_9969,N_9960);
and UO_1129 (O_1129,N_9921,N_9993);
or UO_1130 (O_1130,N_9955,N_9949);
or UO_1131 (O_1131,N_9940,N_9942);
nor UO_1132 (O_1132,N_9917,N_9979);
nand UO_1133 (O_1133,N_9957,N_9991);
or UO_1134 (O_1134,N_9960,N_9934);
xnor UO_1135 (O_1135,N_9991,N_9945);
nor UO_1136 (O_1136,N_9934,N_9938);
nor UO_1137 (O_1137,N_9951,N_9975);
and UO_1138 (O_1138,N_9908,N_9907);
nor UO_1139 (O_1139,N_9917,N_9903);
and UO_1140 (O_1140,N_9963,N_9905);
nor UO_1141 (O_1141,N_9910,N_9963);
nand UO_1142 (O_1142,N_9940,N_9978);
and UO_1143 (O_1143,N_9931,N_9929);
nand UO_1144 (O_1144,N_9926,N_9993);
or UO_1145 (O_1145,N_9921,N_9901);
and UO_1146 (O_1146,N_9955,N_9952);
nand UO_1147 (O_1147,N_9944,N_9961);
nand UO_1148 (O_1148,N_9911,N_9938);
or UO_1149 (O_1149,N_9914,N_9964);
nand UO_1150 (O_1150,N_9957,N_9977);
and UO_1151 (O_1151,N_9980,N_9971);
nor UO_1152 (O_1152,N_9925,N_9995);
nand UO_1153 (O_1153,N_9967,N_9955);
nor UO_1154 (O_1154,N_9977,N_9912);
and UO_1155 (O_1155,N_9950,N_9904);
or UO_1156 (O_1156,N_9985,N_9986);
and UO_1157 (O_1157,N_9975,N_9944);
nand UO_1158 (O_1158,N_9993,N_9937);
nand UO_1159 (O_1159,N_9959,N_9980);
nor UO_1160 (O_1160,N_9937,N_9994);
and UO_1161 (O_1161,N_9917,N_9940);
nor UO_1162 (O_1162,N_9909,N_9915);
and UO_1163 (O_1163,N_9931,N_9938);
or UO_1164 (O_1164,N_9913,N_9982);
or UO_1165 (O_1165,N_9974,N_9987);
xor UO_1166 (O_1166,N_9970,N_9919);
or UO_1167 (O_1167,N_9901,N_9973);
or UO_1168 (O_1168,N_9986,N_9987);
and UO_1169 (O_1169,N_9960,N_9980);
nor UO_1170 (O_1170,N_9913,N_9916);
or UO_1171 (O_1171,N_9955,N_9977);
nand UO_1172 (O_1172,N_9928,N_9937);
nor UO_1173 (O_1173,N_9994,N_9946);
nand UO_1174 (O_1174,N_9941,N_9924);
or UO_1175 (O_1175,N_9958,N_9948);
nand UO_1176 (O_1176,N_9998,N_9909);
nand UO_1177 (O_1177,N_9976,N_9995);
and UO_1178 (O_1178,N_9944,N_9969);
nand UO_1179 (O_1179,N_9914,N_9907);
or UO_1180 (O_1180,N_9963,N_9952);
nor UO_1181 (O_1181,N_9929,N_9995);
nor UO_1182 (O_1182,N_9939,N_9985);
nor UO_1183 (O_1183,N_9982,N_9914);
nor UO_1184 (O_1184,N_9954,N_9999);
nor UO_1185 (O_1185,N_9924,N_9957);
or UO_1186 (O_1186,N_9965,N_9925);
or UO_1187 (O_1187,N_9978,N_9937);
and UO_1188 (O_1188,N_9985,N_9959);
and UO_1189 (O_1189,N_9953,N_9918);
and UO_1190 (O_1190,N_9916,N_9918);
nor UO_1191 (O_1191,N_9942,N_9945);
nand UO_1192 (O_1192,N_9937,N_9972);
nand UO_1193 (O_1193,N_9950,N_9992);
and UO_1194 (O_1194,N_9928,N_9974);
and UO_1195 (O_1195,N_9976,N_9966);
nand UO_1196 (O_1196,N_9955,N_9956);
nor UO_1197 (O_1197,N_9936,N_9962);
nand UO_1198 (O_1198,N_9932,N_9944);
nor UO_1199 (O_1199,N_9917,N_9906);
nor UO_1200 (O_1200,N_9974,N_9970);
nand UO_1201 (O_1201,N_9948,N_9909);
nor UO_1202 (O_1202,N_9990,N_9907);
or UO_1203 (O_1203,N_9902,N_9978);
nor UO_1204 (O_1204,N_9933,N_9942);
or UO_1205 (O_1205,N_9955,N_9932);
and UO_1206 (O_1206,N_9957,N_9986);
nand UO_1207 (O_1207,N_9953,N_9913);
and UO_1208 (O_1208,N_9980,N_9986);
nor UO_1209 (O_1209,N_9986,N_9964);
nor UO_1210 (O_1210,N_9910,N_9928);
nor UO_1211 (O_1211,N_9966,N_9936);
or UO_1212 (O_1212,N_9936,N_9932);
nor UO_1213 (O_1213,N_9900,N_9954);
or UO_1214 (O_1214,N_9961,N_9924);
nand UO_1215 (O_1215,N_9943,N_9912);
nor UO_1216 (O_1216,N_9968,N_9967);
nor UO_1217 (O_1217,N_9904,N_9978);
and UO_1218 (O_1218,N_9965,N_9996);
or UO_1219 (O_1219,N_9991,N_9999);
nor UO_1220 (O_1220,N_9916,N_9991);
nand UO_1221 (O_1221,N_9968,N_9921);
and UO_1222 (O_1222,N_9909,N_9944);
and UO_1223 (O_1223,N_9984,N_9925);
or UO_1224 (O_1224,N_9902,N_9928);
nor UO_1225 (O_1225,N_9966,N_9991);
nor UO_1226 (O_1226,N_9928,N_9964);
nor UO_1227 (O_1227,N_9940,N_9954);
and UO_1228 (O_1228,N_9940,N_9901);
nand UO_1229 (O_1229,N_9904,N_9999);
nor UO_1230 (O_1230,N_9915,N_9916);
or UO_1231 (O_1231,N_9976,N_9992);
and UO_1232 (O_1232,N_9973,N_9955);
and UO_1233 (O_1233,N_9931,N_9953);
nor UO_1234 (O_1234,N_9962,N_9933);
nand UO_1235 (O_1235,N_9908,N_9951);
or UO_1236 (O_1236,N_9954,N_9918);
or UO_1237 (O_1237,N_9960,N_9961);
nor UO_1238 (O_1238,N_9943,N_9985);
nand UO_1239 (O_1239,N_9930,N_9905);
nor UO_1240 (O_1240,N_9936,N_9981);
and UO_1241 (O_1241,N_9961,N_9920);
and UO_1242 (O_1242,N_9946,N_9936);
or UO_1243 (O_1243,N_9961,N_9984);
and UO_1244 (O_1244,N_9976,N_9924);
or UO_1245 (O_1245,N_9950,N_9903);
and UO_1246 (O_1246,N_9952,N_9936);
or UO_1247 (O_1247,N_9981,N_9934);
and UO_1248 (O_1248,N_9944,N_9923);
nor UO_1249 (O_1249,N_9915,N_9957);
and UO_1250 (O_1250,N_9947,N_9969);
or UO_1251 (O_1251,N_9944,N_9904);
nor UO_1252 (O_1252,N_9990,N_9954);
nand UO_1253 (O_1253,N_9972,N_9992);
nor UO_1254 (O_1254,N_9987,N_9968);
or UO_1255 (O_1255,N_9944,N_9902);
and UO_1256 (O_1256,N_9957,N_9901);
or UO_1257 (O_1257,N_9998,N_9937);
or UO_1258 (O_1258,N_9964,N_9990);
or UO_1259 (O_1259,N_9987,N_9931);
nand UO_1260 (O_1260,N_9900,N_9952);
nand UO_1261 (O_1261,N_9969,N_9903);
nand UO_1262 (O_1262,N_9923,N_9915);
or UO_1263 (O_1263,N_9986,N_9902);
or UO_1264 (O_1264,N_9978,N_9953);
and UO_1265 (O_1265,N_9997,N_9920);
nor UO_1266 (O_1266,N_9908,N_9914);
nor UO_1267 (O_1267,N_9982,N_9901);
or UO_1268 (O_1268,N_9972,N_9987);
and UO_1269 (O_1269,N_9939,N_9935);
nand UO_1270 (O_1270,N_9938,N_9981);
or UO_1271 (O_1271,N_9905,N_9962);
and UO_1272 (O_1272,N_9930,N_9937);
xor UO_1273 (O_1273,N_9995,N_9953);
or UO_1274 (O_1274,N_9916,N_9930);
nor UO_1275 (O_1275,N_9939,N_9929);
or UO_1276 (O_1276,N_9932,N_9928);
or UO_1277 (O_1277,N_9947,N_9979);
nand UO_1278 (O_1278,N_9907,N_9967);
nor UO_1279 (O_1279,N_9912,N_9991);
nand UO_1280 (O_1280,N_9938,N_9978);
xnor UO_1281 (O_1281,N_9974,N_9973);
nor UO_1282 (O_1282,N_9985,N_9901);
nor UO_1283 (O_1283,N_9933,N_9985);
nand UO_1284 (O_1284,N_9914,N_9953);
and UO_1285 (O_1285,N_9990,N_9941);
nand UO_1286 (O_1286,N_9984,N_9948);
and UO_1287 (O_1287,N_9946,N_9948);
and UO_1288 (O_1288,N_9935,N_9980);
nor UO_1289 (O_1289,N_9973,N_9902);
and UO_1290 (O_1290,N_9947,N_9968);
or UO_1291 (O_1291,N_9957,N_9950);
or UO_1292 (O_1292,N_9994,N_9989);
nor UO_1293 (O_1293,N_9926,N_9911);
or UO_1294 (O_1294,N_9934,N_9942);
nor UO_1295 (O_1295,N_9913,N_9993);
or UO_1296 (O_1296,N_9907,N_9954);
nand UO_1297 (O_1297,N_9939,N_9977);
or UO_1298 (O_1298,N_9938,N_9996);
nor UO_1299 (O_1299,N_9984,N_9923);
nor UO_1300 (O_1300,N_9993,N_9911);
nor UO_1301 (O_1301,N_9904,N_9958);
or UO_1302 (O_1302,N_9988,N_9958);
nor UO_1303 (O_1303,N_9956,N_9994);
nor UO_1304 (O_1304,N_9943,N_9921);
and UO_1305 (O_1305,N_9909,N_9903);
and UO_1306 (O_1306,N_9915,N_9999);
nand UO_1307 (O_1307,N_9971,N_9915);
nor UO_1308 (O_1308,N_9938,N_9918);
and UO_1309 (O_1309,N_9933,N_9947);
nor UO_1310 (O_1310,N_9904,N_9912);
nand UO_1311 (O_1311,N_9948,N_9952);
and UO_1312 (O_1312,N_9913,N_9968);
nor UO_1313 (O_1313,N_9927,N_9919);
or UO_1314 (O_1314,N_9989,N_9940);
or UO_1315 (O_1315,N_9903,N_9977);
and UO_1316 (O_1316,N_9945,N_9967);
nand UO_1317 (O_1317,N_9911,N_9987);
or UO_1318 (O_1318,N_9925,N_9976);
or UO_1319 (O_1319,N_9966,N_9913);
nand UO_1320 (O_1320,N_9995,N_9992);
nand UO_1321 (O_1321,N_9921,N_9917);
nand UO_1322 (O_1322,N_9992,N_9930);
or UO_1323 (O_1323,N_9932,N_9985);
nor UO_1324 (O_1324,N_9933,N_9916);
and UO_1325 (O_1325,N_9904,N_9934);
nor UO_1326 (O_1326,N_9920,N_9946);
nand UO_1327 (O_1327,N_9983,N_9990);
and UO_1328 (O_1328,N_9931,N_9993);
nand UO_1329 (O_1329,N_9957,N_9981);
nor UO_1330 (O_1330,N_9971,N_9933);
nand UO_1331 (O_1331,N_9977,N_9907);
or UO_1332 (O_1332,N_9932,N_9973);
or UO_1333 (O_1333,N_9911,N_9920);
and UO_1334 (O_1334,N_9997,N_9922);
nor UO_1335 (O_1335,N_9916,N_9962);
nand UO_1336 (O_1336,N_9964,N_9936);
nor UO_1337 (O_1337,N_9980,N_9926);
nand UO_1338 (O_1338,N_9996,N_9939);
nor UO_1339 (O_1339,N_9981,N_9941);
nand UO_1340 (O_1340,N_9970,N_9981);
and UO_1341 (O_1341,N_9903,N_9926);
or UO_1342 (O_1342,N_9951,N_9996);
nand UO_1343 (O_1343,N_9927,N_9963);
nand UO_1344 (O_1344,N_9989,N_9952);
nand UO_1345 (O_1345,N_9907,N_9964);
and UO_1346 (O_1346,N_9901,N_9968);
or UO_1347 (O_1347,N_9955,N_9934);
and UO_1348 (O_1348,N_9996,N_9983);
nor UO_1349 (O_1349,N_9953,N_9968);
xnor UO_1350 (O_1350,N_9927,N_9906);
or UO_1351 (O_1351,N_9991,N_9950);
or UO_1352 (O_1352,N_9938,N_9961);
or UO_1353 (O_1353,N_9916,N_9978);
or UO_1354 (O_1354,N_9999,N_9949);
nor UO_1355 (O_1355,N_9947,N_9938);
or UO_1356 (O_1356,N_9967,N_9934);
or UO_1357 (O_1357,N_9900,N_9957);
nand UO_1358 (O_1358,N_9962,N_9939);
and UO_1359 (O_1359,N_9905,N_9974);
xnor UO_1360 (O_1360,N_9906,N_9926);
nor UO_1361 (O_1361,N_9991,N_9937);
nor UO_1362 (O_1362,N_9949,N_9929);
nand UO_1363 (O_1363,N_9990,N_9976);
and UO_1364 (O_1364,N_9903,N_9968);
nand UO_1365 (O_1365,N_9929,N_9948);
nor UO_1366 (O_1366,N_9943,N_9954);
or UO_1367 (O_1367,N_9968,N_9916);
nand UO_1368 (O_1368,N_9958,N_9920);
and UO_1369 (O_1369,N_9981,N_9915);
nor UO_1370 (O_1370,N_9931,N_9912);
and UO_1371 (O_1371,N_9983,N_9986);
nand UO_1372 (O_1372,N_9968,N_9990);
and UO_1373 (O_1373,N_9970,N_9940);
nand UO_1374 (O_1374,N_9949,N_9908);
nand UO_1375 (O_1375,N_9940,N_9993);
nor UO_1376 (O_1376,N_9943,N_9994);
and UO_1377 (O_1377,N_9909,N_9901);
nand UO_1378 (O_1378,N_9961,N_9908);
nand UO_1379 (O_1379,N_9959,N_9986);
or UO_1380 (O_1380,N_9938,N_9957);
xor UO_1381 (O_1381,N_9957,N_9910);
nand UO_1382 (O_1382,N_9931,N_9901);
and UO_1383 (O_1383,N_9906,N_9920);
nor UO_1384 (O_1384,N_9971,N_9968);
nor UO_1385 (O_1385,N_9913,N_9922);
nand UO_1386 (O_1386,N_9937,N_9980);
or UO_1387 (O_1387,N_9937,N_9969);
or UO_1388 (O_1388,N_9976,N_9929);
nor UO_1389 (O_1389,N_9943,N_9971);
and UO_1390 (O_1390,N_9956,N_9984);
nand UO_1391 (O_1391,N_9909,N_9957);
and UO_1392 (O_1392,N_9936,N_9984);
nor UO_1393 (O_1393,N_9931,N_9915);
and UO_1394 (O_1394,N_9968,N_9930);
nor UO_1395 (O_1395,N_9907,N_9984);
and UO_1396 (O_1396,N_9971,N_9917);
or UO_1397 (O_1397,N_9961,N_9917);
or UO_1398 (O_1398,N_9944,N_9949);
nand UO_1399 (O_1399,N_9976,N_9986);
nor UO_1400 (O_1400,N_9915,N_9936);
nand UO_1401 (O_1401,N_9922,N_9915);
nand UO_1402 (O_1402,N_9985,N_9928);
and UO_1403 (O_1403,N_9900,N_9932);
or UO_1404 (O_1404,N_9962,N_9999);
nor UO_1405 (O_1405,N_9975,N_9909);
and UO_1406 (O_1406,N_9995,N_9930);
or UO_1407 (O_1407,N_9999,N_9930);
nand UO_1408 (O_1408,N_9915,N_9986);
xor UO_1409 (O_1409,N_9955,N_9901);
and UO_1410 (O_1410,N_9930,N_9939);
and UO_1411 (O_1411,N_9933,N_9904);
or UO_1412 (O_1412,N_9987,N_9940);
nor UO_1413 (O_1413,N_9947,N_9977);
or UO_1414 (O_1414,N_9933,N_9918);
and UO_1415 (O_1415,N_9993,N_9938);
nor UO_1416 (O_1416,N_9928,N_9943);
nand UO_1417 (O_1417,N_9973,N_9943);
or UO_1418 (O_1418,N_9957,N_9940);
nand UO_1419 (O_1419,N_9900,N_9980);
and UO_1420 (O_1420,N_9942,N_9929);
and UO_1421 (O_1421,N_9958,N_9934);
nand UO_1422 (O_1422,N_9974,N_9982);
and UO_1423 (O_1423,N_9905,N_9992);
nor UO_1424 (O_1424,N_9991,N_9970);
nand UO_1425 (O_1425,N_9999,N_9938);
or UO_1426 (O_1426,N_9948,N_9934);
and UO_1427 (O_1427,N_9910,N_9956);
nand UO_1428 (O_1428,N_9938,N_9991);
nor UO_1429 (O_1429,N_9900,N_9946);
nor UO_1430 (O_1430,N_9997,N_9935);
or UO_1431 (O_1431,N_9920,N_9907);
or UO_1432 (O_1432,N_9998,N_9917);
or UO_1433 (O_1433,N_9929,N_9955);
and UO_1434 (O_1434,N_9973,N_9988);
and UO_1435 (O_1435,N_9947,N_9964);
nor UO_1436 (O_1436,N_9949,N_9947);
nor UO_1437 (O_1437,N_9954,N_9972);
nor UO_1438 (O_1438,N_9987,N_9980);
and UO_1439 (O_1439,N_9977,N_9909);
and UO_1440 (O_1440,N_9976,N_9914);
nor UO_1441 (O_1441,N_9965,N_9992);
nor UO_1442 (O_1442,N_9907,N_9971);
and UO_1443 (O_1443,N_9915,N_9977);
and UO_1444 (O_1444,N_9957,N_9955);
and UO_1445 (O_1445,N_9914,N_9973);
nor UO_1446 (O_1446,N_9936,N_9935);
and UO_1447 (O_1447,N_9995,N_9974);
or UO_1448 (O_1448,N_9949,N_9900);
nor UO_1449 (O_1449,N_9990,N_9947);
nand UO_1450 (O_1450,N_9910,N_9976);
and UO_1451 (O_1451,N_9959,N_9900);
nor UO_1452 (O_1452,N_9926,N_9958);
nand UO_1453 (O_1453,N_9987,N_9914);
and UO_1454 (O_1454,N_9991,N_9952);
nand UO_1455 (O_1455,N_9944,N_9966);
or UO_1456 (O_1456,N_9969,N_9975);
or UO_1457 (O_1457,N_9944,N_9911);
nor UO_1458 (O_1458,N_9978,N_9959);
and UO_1459 (O_1459,N_9903,N_9995);
nor UO_1460 (O_1460,N_9965,N_9982);
nand UO_1461 (O_1461,N_9911,N_9964);
and UO_1462 (O_1462,N_9939,N_9905);
or UO_1463 (O_1463,N_9913,N_9912);
and UO_1464 (O_1464,N_9949,N_9945);
and UO_1465 (O_1465,N_9983,N_9948);
nand UO_1466 (O_1466,N_9938,N_9926);
nand UO_1467 (O_1467,N_9938,N_9904);
or UO_1468 (O_1468,N_9963,N_9975);
nand UO_1469 (O_1469,N_9960,N_9974);
and UO_1470 (O_1470,N_9989,N_9942);
nand UO_1471 (O_1471,N_9937,N_9988);
nand UO_1472 (O_1472,N_9926,N_9998);
nand UO_1473 (O_1473,N_9931,N_9979);
or UO_1474 (O_1474,N_9943,N_9960);
xor UO_1475 (O_1475,N_9975,N_9973);
or UO_1476 (O_1476,N_9925,N_9971);
or UO_1477 (O_1477,N_9987,N_9956);
or UO_1478 (O_1478,N_9990,N_9993);
or UO_1479 (O_1479,N_9980,N_9973);
or UO_1480 (O_1480,N_9995,N_9983);
or UO_1481 (O_1481,N_9953,N_9908);
and UO_1482 (O_1482,N_9965,N_9947);
or UO_1483 (O_1483,N_9909,N_9916);
or UO_1484 (O_1484,N_9932,N_9951);
nand UO_1485 (O_1485,N_9949,N_9950);
and UO_1486 (O_1486,N_9921,N_9915);
nand UO_1487 (O_1487,N_9978,N_9933);
nor UO_1488 (O_1488,N_9950,N_9980);
or UO_1489 (O_1489,N_9993,N_9991);
nand UO_1490 (O_1490,N_9936,N_9912);
and UO_1491 (O_1491,N_9940,N_9921);
and UO_1492 (O_1492,N_9926,N_9930);
or UO_1493 (O_1493,N_9913,N_9939);
or UO_1494 (O_1494,N_9994,N_9991);
nor UO_1495 (O_1495,N_9989,N_9938);
or UO_1496 (O_1496,N_9902,N_9950);
or UO_1497 (O_1497,N_9984,N_9966);
nor UO_1498 (O_1498,N_9983,N_9940);
and UO_1499 (O_1499,N_9918,N_9972);
endmodule