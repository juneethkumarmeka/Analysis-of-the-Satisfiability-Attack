module basic_1500_15000_2000_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_597,In_422);
xnor U1 (N_1,In_339,In_48);
nand U2 (N_2,In_466,In_935);
and U3 (N_3,In_461,In_471);
and U4 (N_4,In_1383,In_641);
nand U5 (N_5,In_396,In_1247);
xnor U6 (N_6,In_241,In_221);
xnor U7 (N_7,In_76,In_41);
nand U8 (N_8,In_1060,In_982);
and U9 (N_9,In_1348,In_253);
nor U10 (N_10,In_1279,In_995);
xor U11 (N_11,In_1386,In_197);
and U12 (N_12,In_605,In_963);
nor U13 (N_13,In_341,In_64);
xnor U14 (N_14,In_565,In_366);
xnor U15 (N_15,In_1108,In_1462);
nand U16 (N_16,In_187,In_5);
and U17 (N_17,In_582,In_139);
xnor U18 (N_18,In_259,In_214);
and U19 (N_19,In_711,In_53);
nor U20 (N_20,In_643,In_1358);
and U21 (N_21,In_440,In_9);
xor U22 (N_22,In_1481,In_1143);
nor U23 (N_23,In_491,In_1306);
or U24 (N_24,In_1374,In_1157);
or U25 (N_25,In_68,In_1120);
xnor U26 (N_26,In_26,In_473);
nand U27 (N_27,In_1221,In_634);
xnor U28 (N_28,In_1008,In_560);
and U29 (N_29,In_854,In_934);
nor U30 (N_30,In_195,In_651);
xnor U31 (N_31,In_1458,In_783);
nor U32 (N_32,In_1249,In_355);
and U33 (N_33,In_744,In_117);
nor U34 (N_34,In_137,In_799);
nor U35 (N_35,In_1052,In_67);
nand U36 (N_36,In_1361,In_198);
or U37 (N_37,In_989,In_1127);
and U38 (N_38,In_445,In_147);
or U39 (N_39,In_219,In_1225);
xor U40 (N_40,In_365,In_488);
and U41 (N_41,In_468,In_811);
nor U42 (N_42,In_1230,In_718);
or U43 (N_43,In_533,In_408);
and U44 (N_44,In_880,In_1350);
and U45 (N_45,In_1441,In_826);
and U46 (N_46,In_324,In_1362);
or U47 (N_47,In_820,In_248);
and U48 (N_48,In_1357,In_988);
and U49 (N_49,In_1433,In_169);
or U50 (N_50,In_953,In_1250);
and U51 (N_51,In_792,In_1319);
or U52 (N_52,In_1465,In_872);
nor U53 (N_53,In_98,In_1236);
nand U54 (N_54,In_706,In_805);
nand U55 (N_55,In_454,In_512);
nor U56 (N_56,In_272,In_886);
xnor U57 (N_57,In_516,In_812);
nor U58 (N_58,In_648,In_133);
or U59 (N_59,In_1446,In_238);
nand U60 (N_60,In_91,In_126);
and U61 (N_61,In_979,In_367);
nor U62 (N_62,In_288,In_642);
xor U63 (N_63,In_1258,In_1103);
nand U64 (N_64,In_665,In_1497);
nand U65 (N_65,In_1005,In_112);
and U66 (N_66,In_520,In_65);
and U67 (N_67,In_1283,In_196);
or U68 (N_68,In_142,In_1064);
nand U69 (N_69,In_255,In_120);
xnor U70 (N_70,In_443,In_758);
nand U71 (N_71,In_246,In_791);
nand U72 (N_72,In_121,In_69);
or U73 (N_73,In_376,In_1025);
nand U74 (N_74,In_870,In_1244);
and U75 (N_75,In_1340,In_1309);
nor U76 (N_76,In_920,In_261);
nor U77 (N_77,In_316,In_318);
and U78 (N_78,In_1296,In_1047);
and U79 (N_79,In_1254,In_1292);
or U80 (N_80,In_1149,In_1171);
nand U81 (N_81,In_178,In_431);
xnor U82 (N_82,In_130,In_20);
nand U83 (N_83,In_1499,In_1493);
or U84 (N_84,In_680,In_668);
or U85 (N_85,In_245,In_291);
xnor U86 (N_86,In_229,In_300);
nor U87 (N_87,In_1488,In_110);
nand U88 (N_88,In_536,In_916);
or U89 (N_89,In_1097,In_691);
nand U90 (N_90,In_606,In_774);
nand U91 (N_91,In_150,In_715);
nor U92 (N_92,In_961,In_556);
xor U93 (N_93,In_859,In_284);
nand U94 (N_94,In_1475,In_1241);
nand U95 (N_95,In_185,In_144);
and U96 (N_96,In_476,In_729);
nor U97 (N_97,In_1017,In_759);
or U98 (N_98,In_1086,In_1396);
or U99 (N_99,In_435,In_302);
or U100 (N_100,In_1045,In_1427);
nor U101 (N_101,In_309,In_604);
and U102 (N_102,In_1422,In_100);
or U103 (N_103,In_1484,In_702);
xor U104 (N_104,In_1341,In_1478);
nand U105 (N_105,In_1233,In_497);
nor U106 (N_106,In_1214,In_1451);
and U107 (N_107,In_732,In_1243);
nor U108 (N_108,In_1414,In_1425);
xnor U109 (N_109,In_60,In_118);
or U110 (N_110,In_456,In_849);
nor U111 (N_111,In_1156,In_1454);
nor U112 (N_112,In_297,In_1286);
and U113 (N_113,In_1401,In_1032);
nor U114 (N_114,In_1030,In_393);
nand U115 (N_115,In_1138,In_1257);
and U116 (N_116,In_972,In_1429);
or U117 (N_117,In_1022,In_696);
nor U118 (N_118,In_1150,In_433);
nand U119 (N_119,In_384,In_787);
nand U120 (N_120,In_1310,In_1016);
or U121 (N_121,In_692,In_447);
nor U122 (N_122,In_1308,In_678);
xor U123 (N_123,In_1046,In_924);
and U124 (N_124,In_751,In_1187);
xnor U125 (N_125,In_994,In_1106);
or U126 (N_126,In_448,In_205);
xor U127 (N_127,In_596,In_901);
nor U128 (N_128,In_776,In_176);
nand U129 (N_129,In_136,In_727);
and U130 (N_130,In_855,In_188);
nor U131 (N_131,In_1265,In_1373);
xor U132 (N_132,In_1402,In_830);
nor U133 (N_133,In_814,In_925);
or U134 (N_134,In_1082,In_171);
or U135 (N_135,In_406,In_1067);
or U136 (N_136,In_521,In_168);
xor U137 (N_137,In_518,In_839);
and U138 (N_138,In_1169,In_987);
nand U139 (N_139,In_1463,In_223);
nand U140 (N_140,In_186,In_162);
and U141 (N_141,In_194,In_1194);
nor U142 (N_142,In_501,In_54);
and U143 (N_143,In_270,In_623);
nand U144 (N_144,In_1347,In_107);
nand U145 (N_145,In_1491,In_1232);
and U146 (N_146,In_145,In_1062);
or U147 (N_147,In_489,In_1075);
and U148 (N_148,In_667,In_1173);
and U149 (N_149,In_37,In_247);
nor U150 (N_150,In_170,In_1161);
nand U151 (N_151,In_424,In_103);
and U152 (N_152,In_1264,In_612);
nor U153 (N_153,In_1113,In_917);
xnor U154 (N_154,In_469,In_1080);
nand U155 (N_155,In_189,In_1158);
xnor U156 (N_156,In_1412,In_371);
xnor U157 (N_157,In_1364,In_1333);
or U158 (N_158,In_389,In_1365);
or U159 (N_159,In_412,In_1227);
nor U160 (N_160,In_1163,In_1431);
nand U161 (N_161,In_981,In_784);
and U162 (N_162,In_958,In_598);
or U163 (N_163,In_1144,In_174);
nor U164 (N_164,In_421,In_350);
nor U165 (N_165,In_699,In_904);
nor U166 (N_166,In_588,In_708);
and U167 (N_167,In_1185,In_1384);
nand U168 (N_168,In_985,In_1343);
nand U169 (N_169,In_1039,In_1311);
or U170 (N_170,In_617,In_1159);
nor U171 (N_171,In_243,In_277);
nand U172 (N_172,In_747,In_704);
and U173 (N_173,In_330,In_1302);
or U174 (N_174,In_879,In_964);
nor U175 (N_175,In_77,In_1167);
nand U176 (N_176,In_281,In_16);
xnor U177 (N_177,In_1141,In_449);
or U178 (N_178,In_959,In_1092);
nand U179 (N_179,In_1215,In_111);
nand U180 (N_180,In_608,In_673);
nor U181 (N_181,In_1034,In_1212);
and U182 (N_182,In_362,In_452);
nor U183 (N_183,In_167,In_1222);
nor U184 (N_184,In_211,In_620);
nand U185 (N_185,In_13,In_1000);
and U186 (N_186,In_311,In_1485);
nand U187 (N_187,In_1395,In_881);
nor U188 (N_188,In_1153,In_102);
or U189 (N_189,In_768,In_506);
and U190 (N_190,In_477,In_374);
nor U191 (N_191,In_141,In_731);
nand U192 (N_192,In_965,In_1420);
xnor U193 (N_193,In_1048,In_1002);
or U194 (N_194,In_43,In_538);
or U195 (N_195,In_1188,In_234);
and U196 (N_196,In_282,In_816);
nor U197 (N_197,In_603,In_535);
or U198 (N_198,In_383,In_1);
and U199 (N_199,In_321,In_1419);
xor U200 (N_200,In_662,In_1281);
xnor U201 (N_201,In_1346,In_1124);
xor U202 (N_202,In_1487,In_153);
or U203 (N_203,In_356,In_573);
or U204 (N_204,In_562,In_626);
nor U205 (N_205,In_1455,In_998);
xnor U206 (N_206,In_1162,In_1133);
nand U207 (N_207,In_1177,In_1139);
xor U208 (N_208,In_1331,In_481);
nand U209 (N_209,In_55,In_1399);
and U210 (N_210,In_1111,In_1090);
xnor U211 (N_211,In_584,In_1423);
and U212 (N_212,In_6,In_619);
and U213 (N_213,In_306,In_114);
and U214 (N_214,In_1136,In_465);
and U215 (N_215,In_403,In_1043);
nand U216 (N_216,In_908,In_610);
and U217 (N_217,In_22,In_423);
nor U218 (N_218,In_1245,In_1303);
nand U219 (N_219,In_1466,In_498);
or U220 (N_220,In_803,In_1077);
nor U221 (N_221,In_400,In_286);
nand U222 (N_222,In_1010,In_1007);
xnor U223 (N_223,In_530,In_322);
nand U224 (N_224,In_2,In_652);
xor U225 (N_225,In_191,In_1326);
nand U226 (N_226,In_1262,In_1224);
nand U227 (N_227,In_1129,In_804);
xor U228 (N_228,In_707,In_1059);
nor U229 (N_229,In_546,In_19);
nand U230 (N_230,In_1226,In_761);
or U231 (N_231,In_609,In_1029);
xnor U232 (N_232,In_50,In_1206);
or U233 (N_233,In_1342,In_158);
nand U234 (N_234,In_474,In_1256);
or U235 (N_235,In_765,In_1457);
nand U236 (N_236,In_1426,In_441);
or U237 (N_237,In_1179,In_84);
and U238 (N_238,In_332,In_864);
nand U239 (N_239,In_511,In_900);
and U240 (N_240,In_515,In_716);
and U241 (N_241,In_559,In_88);
xnor U242 (N_242,In_889,In_618);
or U243 (N_243,In_1444,In_601);
and U244 (N_244,In_1440,In_1359);
xor U245 (N_245,In_1411,In_738);
nand U246 (N_246,In_1261,In_1290);
nand U247 (N_247,In_1211,In_347);
or U248 (N_248,In_1018,In_1449);
xor U249 (N_249,In_821,In_779);
nor U250 (N_250,In_1014,In_1316);
and U251 (N_251,In_192,In_554);
and U252 (N_252,In_1155,In_653);
and U253 (N_253,In_996,In_762);
and U254 (N_254,In_17,In_694);
and U255 (N_255,In_392,In_777);
nor U256 (N_256,In_1207,In_359);
or U257 (N_257,In_36,In_841);
xor U258 (N_258,In_1471,In_1028);
nand U259 (N_259,In_1335,In_18);
nor U260 (N_260,In_125,In_225);
nand U261 (N_261,In_978,In_929);
nor U262 (N_262,In_342,In_268);
nor U263 (N_263,In_258,In_381);
xor U264 (N_264,In_1154,In_482);
xor U265 (N_265,In_717,In_660);
nand U266 (N_266,In_845,In_1324);
xor U267 (N_267,In_254,In_1439);
and U268 (N_268,In_1006,In_952);
nand U269 (N_269,In_713,In_1489);
and U270 (N_270,In_640,In_970);
and U271 (N_271,In_838,In_574);
xnor U272 (N_272,In_1021,In_486);
and U273 (N_273,In_1069,In_1368);
and U274 (N_274,In_470,In_459);
and U275 (N_275,In_467,In_567);
and U276 (N_276,In_1375,In_577);
or U277 (N_277,In_1267,In_892);
xor U278 (N_278,In_1255,In_1087);
nor U279 (N_279,In_1389,In_1229);
xnor U280 (N_280,In_1218,In_655);
or U281 (N_281,In_262,In_1360);
nor U282 (N_282,In_884,In_157);
nor U283 (N_283,In_1300,In_428);
or U284 (N_284,In_303,In_1416);
nand U285 (N_285,In_1436,In_911);
nand U286 (N_286,In_541,In_861);
nand U287 (N_287,In_129,In_1418);
or U288 (N_288,In_1410,In_944);
nand U289 (N_289,In_1118,In_782);
or U290 (N_290,In_1321,In_453);
nand U291 (N_291,In_96,In_264);
nor U292 (N_292,In_375,In_720);
nor U293 (N_293,In_148,In_1352);
nand U294 (N_294,In_793,In_921);
xnor U295 (N_295,In_1040,In_1195);
nor U296 (N_296,In_317,In_83);
or U297 (N_297,In_677,In_539);
or U298 (N_298,In_462,In_1011);
or U299 (N_299,In_217,In_1100);
and U300 (N_300,In_583,In_1209);
and U301 (N_301,In_730,In_1234);
xor U302 (N_302,In_278,In_585);
nand U303 (N_303,In_740,In_1417);
nand U304 (N_304,In_1474,In_368);
nand U305 (N_305,In_95,In_496);
xnor U306 (N_306,In_1054,In_1354);
xor U307 (N_307,In_106,In_822);
nor U308 (N_308,In_1088,In_999);
or U309 (N_309,In_1482,In_1024);
or U310 (N_310,In_420,In_1178);
xnor U311 (N_311,In_670,In_47);
nor U312 (N_312,In_134,In_542);
or U313 (N_313,In_75,In_992);
nor U314 (N_314,In_1210,In_79);
and U315 (N_315,In_646,In_955);
xor U316 (N_316,In_639,In_1235);
nand U317 (N_317,In_1404,In_66);
nand U318 (N_318,In_946,In_1351);
nand U319 (N_319,In_401,In_856);
xnor U320 (N_320,In_745,In_877);
nor U321 (N_321,In_1381,In_907);
nand U322 (N_322,In_686,In_1313);
xnor U323 (N_323,In_1282,In_296);
xor U324 (N_324,In_885,In_684);
and U325 (N_325,In_918,In_301);
nor U326 (N_326,In_780,In_714);
or U327 (N_327,In_1130,In_1370);
or U328 (N_328,In_685,In_625);
nor U329 (N_329,In_89,In_775);
nor U330 (N_330,In_746,In_226);
xor U331 (N_331,In_343,In_832);
or U332 (N_332,In_1304,In_388);
xor U333 (N_333,In_320,In_292);
nand U334 (N_334,In_32,In_1307);
and U335 (N_335,In_231,In_1469);
and U336 (N_336,In_109,In_200);
xor U337 (N_337,In_1074,In_42);
xor U338 (N_338,In_1033,In_1152);
xnor U339 (N_339,In_1200,In_1242);
or U340 (N_340,In_1083,In_1322);
nand U341 (N_341,In_1170,In_1252);
nor U342 (N_342,In_70,In_1231);
xor U343 (N_343,In_755,In_517);
and U344 (N_344,In_349,In_558);
or U345 (N_345,In_1098,In_502);
xnor U346 (N_346,In_1430,In_980);
nor U347 (N_347,In_1470,In_1066);
or U348 (N_348,In_1228,In_0);
nor U349 (N_349,In_644,In_834);
and U350 (N_350,In_455,In_1263);
and U351 (N_351,In_119,In_1091);
or U352 (N_352,In_661,In_1398);
xnor U353 (N_353,In_969,In_569);
and U354 (N_354,In_926,In_1330);
nand U355 (N_355,In_1084,In_394);
and U356 (N_356,In_1174,In_913);
or U357 (N_357,In_806,In_1192);
nand U358 (N_358,In_578,In_1145);
or U359 (N_359,In_664,In_887);
or U360 (N_360,In_363,In_257);
nand U361 (N_361,In_681,In_507);
nand U362 (N_362,In_968,In_915);
nor U363 (N_363,In_687,In_1085);
and U364 (N_364,In_1004,In_809);
nor U365 (N_365,In_1142,In_1438);
and U366 (N_366,In_439,In_798);
and U367 (N_367,In_712,In_275);
and U368 (N_368,In_202,In_271);
and U369 (N_369,In_116,In_1219);
xor U370 (N_370,In_847,In_947);
xnor U371 (N_371,In_1134,In_397);
nand U372 (N_372,In_1334,In_337);
and U373 (N_373,In_293,In_1121);
and U374 (N_374,In_416,In_15);
nand U375 (N_375,In_624,In_1151);
and U376 (N_376,In_310,In_549);
nor U377 (N_377,In_682,In_1371);
nand U378 (N_378,In_790,In_236);
nor U379 (N_379,In_338,In_446);
nand U380 (N_380,In_207,In_671);
nand U381 (N_381,In_1239,In_635);
nor U382 (N_382,In_1201,In_7);
and U383 (N_383,In_483,In_23);
xnor U384 (N_384,In_1394,In_1477);
and U385 (N_385,In_58,In_1405);
nand U386 (N_386,In_127,In_571);
xnor U387 (N_387,In_524,In_239);
xor U388 (N_388,In_224,In_951);
or U389 (N_389,In_352,In_260);
nand U390 (N_390,In_748,In_846);
xnor U391 (N_391,In_544,In_1176);
nand U392 (N_392,In_1293,In_1023);
or U393 (N_393,In_974,In_163);
xor U394 (N_394,In_563,In_1435);
nand U395 (N_395,In_490,In_801);
and U396 (N_396,In_657,In_829);
nand U397 (N_397,In_897,In_1146);
nand U398 (N_398,In_629,In_519);
or U399 (N_399,In_1336,In_1403);
xnor U400 (N_400,In_1367,In_132);
nor U401 (N_401,In_950,In_99);
nand U402 (N_402,In_1442,In_611);
and U403 (N_403,In_631,In_1205);
and U404 (N_404,In_1388,In_74);
xnor U405 (N_405,In_430,In_882);
xor U406 (N_406,In_244,In_616);
xnor U407 (N_407,In_1392,In_1058);
nand U408 (N_408,In_1285,In_46);
and U409 (N_409,In_331,In_1012);
nand U410 (N_410,In_410,In_531);
xor U411 (N_411,In_1056,In_51);
nor U412 (N_412,In_326,In_910);
or U413 (N_413,In_1314,In_115);
nand U414 (N_414,In_723,In_698);
xnor U415 (N_415,In_123,In_532);
xnor U416 (N_416,In_44,In_636);
nor U417 (N_417,In_1128,In_576);
nand U418 (N_418,In_1203,In_510);
nor U419 (N_419,In_160,In_92);
xnor U420 (N_420,In_927,In_1180);
nand U421 (N_421,In_39,In_590);
and U422 (N_422,In_1223,In_369);
or U423 (N_423,In_402,In_334);
or U424 (N_424,In_525,In_1496);
or U425 (N_425,In_426,In_672);
and U426 (N_426,In_31,In_312);
nand U427 (N_427,In_1432,In_30);
and U428 (N_428,In_1345,In_984);
or U429 (N_429,In_945,In_1093);
or U430 (N_430,In_155,In_561);
nor U431 (N_431,In_14,In_570);
nor U432 (N_432,In_1437,In_464);
xor U433 (N_433,In_690,In_177);
nand U434 (N_434,In_1494,In_1363);
and U435 (N_435,In_1278,In_213);
and U436 (N_436,In_266,In_1182);
xnor U437 (N_437,In_848,In_249);
nand U438 (N_438,In_658,In_97);
nand U439 (N_439,In_1044,In_432);
xnor U440 (N_440,In_728,In_807);
nor U441 (N_441,In_954,In_28);
xnor U442 (N_442,In_1165,In_346);
nor U443 (N_443,In_1125,In_372);
xor U444 (N_444,In_404,In_895);
or U445 (N_445,In_939,In_869);
nand U446 (N_446,In_263,In_1081);
nor U447 (N_447,In_695,In_796);
nand U448 (N_448,In_943,In_852);
xor U449 (N_449,In_437,In_1198);
or U450 (N_450,In_860,In_743);
nor U451 (N_451,In_418,In_844);
nand U452 (N_452,In_553,In_1015);
nor U453 (N_453,In_242,In_1037);
nor U454 (N_454,In_851,In_298);
nor U455 (N_455,In_11,In_164);
xor U456 (N_456,In_735,In_705);
or U457 (N_457,In_1073,In_269);
xnor U458 (N_458,In_1001,In_1240);
nor U459 (N_459,In_547,In_866);
nor U460 (N_460,In_166,In_587);
nand U461 (N_461,In_592,In_767);
xnor U462 (N_462,In_1372,In_1329);
xor U463 (N_463,In_206,In_1041);
nor U464 (N_464,In_1137,In_764);
nand U465 (N_465,In_1377,In_333);
and U466 (N_466,In_267,In_57);
nand U467 (N_467,In_122,In_523);
and U468 (N_468,In_201,In_813);
nand U469 (N_469,In_997,In_1332);
xor U470 (N_470,In_290,In_1275);
and U471 (N_471,In_545,In_526);
xnor U472 (N_472,In_938,In_283);
and U473 (N_473,In_415,In_613);
or U474 (N_474,In_81,In_819);
nand U475 (N_475,In_450,In_893);
nand U476 (N_476,In_701,In_429);
and U477 (N_477,In_902,In_1495);
nor U478 (N_478,In_78,In_875);
or U479 (N_479,In_1038,In_500);
or U480 (N_480,In_865,In_627);
xor U481 (N_481,In_632,In_210);
and U482 (N_482,In_1102,In_1390);
or U483 (N_483,In_199,In_1190);
xor U484 (N_484,In_390,In_3);
xor U485 (N_485,In_600,In_86);
xor U486 (N_486,In_82,In_579);
xor U487 (N_487,In_1049,In_760);
and U488 (N_488,In_1301,In_750);
nor U489 (N_489,In_548,In_1328);
nor U490 (N_490,In_1382,In_8);
and U491 (N_491,In_551,In_1294);
nor U492 (N_492,In_357,In_949);
nand U493 (N_493,In_29,In_252);
and U494 (N_494,In_940,In_514);
or U495 (N_495,In_581,In_1096);
nand U496 (N_496,In_360,In_1216);
nor U497 (N_497,In_328,In_1110);
or U498 (N_498,In_912,In_863);
and U499 (N_499,In_1453,In_344);
xor U500 (N_500,In_937,In_825);
nor U501 (N_501,In_928,In_1183);
nor U502 (N_502,In_227,In_179);
and U503 (N_503,In_1027,In_1238);
nor U504 (N_504,In_1270,In_1107);
or U505 (N_505,In_222,In_572);
nand U506 (N_506,In_124,In_599);
nor U507 (N_507,In_1445,In_930);
nand U508 (N_508,In_1327,In_308);
nor U509 (N_509,In_184,In_1400);
or U510 (N_510,In_1325,In_1095);
nand U511 (N_511,In_1406,In_1135);
xnor U512 (N_512,In_753,In_1237);
nor U513 (N_513,In_494,In_1184);
xor U514 (N_514,In_1276,In_1160);
xor U515 (N_515,In_128,In_679);
xor U516 (N_516,In_734,In_580);
nand U517 (N_517,In_1467,In_1447);
or U518 (N_518,In_786,In_12);
and U519 (N_519,In_138,In_444);
nand U520 (N_520,In_721,In_663);
nor U521 (N_521,In_151,In_1298);
and U522 (N_522,In_1288,In_967);
or U523 (N_523,In_1315,In_237);
nor U524 (N_524,In_1117,In_1119);
nor U525 (N_525,In_522,In_817);
nand U526 (N_526,In_71,In_203);
nand U527 (N_527,In_319,In_492);
nor U528 (N_528,In_1186,In_645);
and U529 (N_529,In_1376,In_1369);
nor U530 (N_530,In_1013,In_1112);
and U531 (N_531,In_305,In_990);
nor U532 (N_532,In_105,In_1397);
nor U533 (N_533,In_85,In_216);
nand U534 (N_534,In_1248,In_1339);
or U535 (N_535,In_1166,In_40);
or U536 (N_536,In_649,In_183);
or U537 (N_537,In_479,In_1366);
xor U538 (N_538,In_135,In_919);
and U539 (N_539,In_1280,In_472);
and U540 (N_540,In_72,In_621);
xnor U541 (N_541,In_399,In_914);
xnor U542 (N_542,In_669,In_983);
or U543 (N_543,In_922,In_1337);
or U544 (N_544,In_1213,In_769);
nand U545 (N_545,In_348,In_458);
nand U546 (N_546,In_905,In_867);
and U547 (N_547,In_94,In_909);
and U548 (N_548,In_250,In_299);
xnor U549 (N_549,In_1197,In_380);
and U550 (N_550,In_1385,In_1476);
nand U551 (N_551,In_552,In_828);
and U552 (N_552,In_1109,In_1353);
xnor U553 (N_553,In_529,In_874);
nand U554 (N_554,In_193,In_256);
nand U555 (N_555,In_1126,In_1055);
nand U556 (N_556,In_1448,In_827);
and U557 (N_557,In_434,In_478);
xnor U558 (N_558,In_175,In_931);
nor U559 (N_559,In_749,In_1253);
nor U560 (N_560,In_149,In_414);
and U561 (N_561,In_700,In_485);
and U562 (N_562,In_528,In_10);
nand U563 (N_563,In_1140,In_1019);
nand U564 (N_564,In_903,In_52);
nor U565 (N_565,In_45,In_1204);
and U566 (N_566,In_836,In_21);
or U567 (N_567,In_1480,In_59);
and U568 (N_568,In_1456,In_1393);
nor U569 (N_569,In_1259,In_891);
nand U570 (N_570,In_973,In_736);
and U571 (N_571,In_628,In_493);
and U572 (N_572,In_1271,In_789);
nor U573 (N_573,In_1260,In_614);
or U574 (N_574,In_487,In_56);
nand U575 (N_575,In_1421,In_1409);
nand U576 (N_576,In_287,In_304);
xor U577 (N_577,In_173,In_1492);
xor U578 (N_578,In_742,In_991);
nor U579 (N_579,In_858,In_1434);
nand U580 (N_580,In_325,In_329);
nor U581 (N_581,In_1408,In_285);
or U582 (N_582,In_725,In_87);
and U583 (N_583,In_868,In_899);
nor U584 (N_584,In_1168,In_741);
or U585 (N_585,In_505,In_4);
and U586 (N_586,In_733,In_824);
and U587 (N_587,In_1486,In_273);
nand U588 (N_588,In_1317,In_407);
nor U589 (N_589,In_557,In_888);
xnor U590 (N_590,In_754,In_960);
nor U591 (N_591,In_818,In_763);
and U592 (N_592,In_209,In_93);
xor U593 (N_593,In_417,In_391);
and U594 (N_594,In_878,In_35);
or U595 (N_595,In_1202,In_1172);
nor U596 (N_596,In_1191,In_638);
nand U597 (N_597,In_413,In_1181);
xnor U598 (N_598,In_361,In_977);
xor U599 (N_599,In_1057,In_49);
or U600 (N_600,In_156,In_1312);
xnor U601 (N_601,In_586,In_794);
or U602 (N_602,In_315,In_364);
nand U603 (N_603,In_1070,In_499);
nor U604 (N_604,In_513,In_1305);
and U605 (N_605,In_1003,In_451);
nor U606 (N_606,In_1026,In_25);
and U607 (N_607,In_757,In_674);
and U608 (N_608,In_1356,In_161);
and U609 (N_609,In_387,In_370);
nor U610 (N_610,In_1413,In_140);
nor U611 (N_611,In_33,In_104);
nand U612 (N_612,In_143,In_208);
nor U613 (N_613,In_154,In_382);
or U614 (N_614,In_923,In_802);
nand U615 (N_615,In_379,In_377);
nand U616 (N_616,In_737,In_411);
nand U617 (N_617,In_647,In_1175);
nand U618 (N_618,In_575,In_795);
xnor U619 (N_619,In_1428,In_726);
nor U620 (N_620,In_182,In_962);
and U621 (N_621,In_480,In_1147);
nor U622 (N_622,In_228,In_113);
xnor U623 (N_623,In_395,In_336);
nand U624 (N_624,In_1072,In_833);
nor U625 (N_625,In_1415,In_986);
nor U626 (N_626,In_823,In_527);
nand U627 (N_627,In_1391,In_220);
xnor U628 (N_628,In_1076,In_594);
nor U629 (N_629,In_265,In_1246);
and U630 (N_630,In_276,In_1031);
nor U631 (N_631,In_463,In_883);
or U632 (N_632,In_373,In_108);
and U633 (N_633,In_537,In_1284);
or U634 (N_634,In_906,In_815);
nand U635 (N_635,In_484,In_898);
and U636 (N_636,In_351,In_405);
and U637 (N_637,In_327,In_637);
nand U638 (N_638,In_703,In_948);
and U639 (N_639,In_1189,In_1105);
xor U640 (N_640,In_280,In_976);
or U641 (N_641,In_666,In_1068);
nor U642 (N_642,In_1114,In_442);
or U643 (N_643,In_1461,In_1268);
xnor U644 (N_644,In_1490,In_890);
and U645 (N_645,In_1387,In_1115);
and U646 (N_646,In_181,In_1407);
and U647 (N_647,In_314,In_800);
nor U648 (N_648,In_218,In_1220);
xnor U649 (N_649,In_756,In_1061);
xnor U650 (N_650,In_475,In_1208);
or U651 (N_651,In_34,In_340);
and U652 (N_652,In_1460,In_38);
and U653 (N_653,In_165,In_693);
or U654 (N_654,In_504,In_771);
xor U655 (N_655,In_1450,In_543);
or U656 (N_656,In_1078,In_1318);
nand U657 (N_657,In_436,In_1020);
or U658 (N_658,In_73,In_1101);
nand U659 (N_659,In_564,In_1123);
and U660 (N_660,In_862,In_146);
or U661 (N_661,In_425,In_295);
and U662 (N_662,In_1131,In_1132);
nand U663 (N_663,In_409,In_1344);
nand U664 (N_664,In_622,In_1036);
nor U665 (N_665,In_152,In_781);
nand U666 (N_666,In_654,In_233);
and U667 (N_667,In_1269,In_850);
or U668 (N_668,In_689,In_788);
or U669 (N_669,In_555,In_1063);
and U670 (N_670,In_80,In_589);
or U671 (N_671,In_419,In_971);
and U672 (N_672,In_495,In_710);
or U673 (N_673,In_1035,In_1483);
nand U674 (N_674,In_101,In_797);
nand U675 (N_675,In_837,In_27);
or U676 (N_676,In_633,In_932);
and U677 (N_677,In_894,In_1065);
nor U678 (N_678,In_773,In_190);
and U679 (N_679,In_785,In_131);
and U680 (N_680,In_896,In_251);
or U681 (N_681,In_550,In_770);
or U682 (N_682,In_1079,In_1196);
nor U683 (N_683,In_534,In_1473);
and U684 (N_684,In_1009,In_1053);
or U685 (N_685,In_1050,In_602);
nor U686 (N_686,In_1289,In_61);
nand U687 (N_687,In_810,In_358);
xnor U688 (N_688,In_724,In_843);
or U689 (N_689,In_956,In_709);
nor U690 (N_690,In_1472,In_159);
nor U691 (N_691,In_204,In_1272);
or U692 (N_692,In_540,In_993);
and U693 (N_693,In_1273,In_378);
or U694 (N_694,In_739,In_427);
or U695 (N_695,In_1299,In_62);
and U696 (N_696,In_853,In_871);
nand U697 (N_697,In_1498,In_1193);
nor U698 (N_698,In_335,In_180);
nand U699 (N_699,In_386,In_1295);
or U700 (N_700,In_1349,In_240);
nor U701 (N_701,In_460,In_212);
xnor U702 (N_702,In_1042,In_508);
nand U703 (N_703,In_1452,In_941);
or U704 (N_704,In_840,In_697);
or U705 (N_705,In_615,In_1116);
nor U706 (N_706,In_215,In_772);
and U707 (N_707,In_966,In_1355);
nand U708 (N_708,In_1379,In_933);
xor U709 (N_709,In_398,In_1323);
or U710 (N_710,In_857,In_842);
or U711 (N_711,In_438,In_1051);
xor U712 (N_712,In_323,In_503);
xnor U713 (N_713,In_1266,In_1164);
and U714 (N_714,In_778,In_274);
nor U715 (N_715,In_957,In_63);
xor U716 (N_716,In_566,In_1148);
and U717 (N_717,In_1071,In_1251);
nor U718 (N_718,In_385,In_656);
xor U719 (N_719,In_1199,In_1443);
xnor U720 (N_720,In_591,In_595);
nor U721 (N_721,In_676,In_975);
and U722 (N_722,In_688,In_1338);
nor U723 (N_723,In_593,In_650);
and U724 (N_724,In_1464,In_90);
nor U725 (N_725,In_942,In_831);
nand U726 (N_726,In_1297,In_509);
and U727 (N_727,In_354,In_230);
and U728 (N_728,In_353,In_279);
nand U729 (N_729,In_1320,In_873);
or U730 (N_730,In_936,In_1291);
nor U731 (N_731,In_1217,In_675);
xnor U732 (N_732,In_232,In_307);
nand U733 (N_733,In_568,In_835);
or U734 (N_734,In_1089,In_1094);
nand U735 (N_735,In_766,In_1277);
nand U736 (N_736,In_289,In_1274);
and U737 (N_737,In_876,In_1468);
or U738 (N_738,In_457,In_1378);
nor U739 (N_739,In_808,In_294);
xnor U740 (N_740,In_607,In_235);
xnor U741 (N_741,In_752,In_1122);
or U742 (N_742,In_722,In_1459);
xnor U743 (N_743,In_172,In_1104);
and U744 (N_744,In_659,In_1380);
nor U745 (N_745,In_683,In_1424);
xnor U746 (N_746,In_1479,In_1099);
xnor U747 (N_747,In_24,In_345);
or U748 (N_748,In_313,In_630);
nor U749 (N_749,In_1287,In_719);
and U750 (N_750,N_330,N_70);
and U751 (N_751,N_476,N_123);
nor U752 (N_752,N_299,N_646);
and U753 (N_753,N_453,N_213);
nor U754 (N_754,N_87,N_712);
and U755 (N_755,N_252,N_422);
xnor U756 (N_756,N_388,N_734);
and U757 (N_757,N_429,N_568);
nand U758 (N_758,N_524,N_490);
nand U759 (N_759,N_120,N_426);
or U760 (N_760,N_84,N_259);
xor U761 (N_761,N_468,N_88);
or U762 (N_762,N_415,N_203);
xor U763 (N_763,N_147,N_258);
nor U764 (N_764,N_565,N_585);
or U765 (N_765,N_127,N_362);
and U766 (N_766,N_232,N_484);
xnor U767 (N_767,N_738,N_178);
nor U768 (N_768,N_79,N_139);
xor U769 (N_769,N_518,N_511);
xor U770 (N_770,N_412,N_242);
nand U771 (N_771,N_647,N_354);
nand U772 (N_772,N_221,N_684);
or U773 (N_773,N_576,N_327);
nor U774 (N_774,N_472,N_6);
xor U775 (N_775,N_621,N_133);
nand U776 (N_776,N_705,N_627);
nor U777 (N_777,N_690,N_204);
xor U778 (N_778,N_340,N_248);
nor U779 (N_779,N_143,N_142);
or U780 (N_780,N_477,N_391);
or U781 (N_781,N_77,N_282);
and U782 (N_782,N_372,N_152);
or U783 (N_783,N_706,N_250);
and U784 (N_784,N_377,N_651);
nand U785 (N_785,N_102,N_369);
and U786 (N_786,N_664,N_487);
nor U787 (N_787,N_385,N_708);
or U788 (N_788,N_243,N_82);
nor U789 (N_789,N_14,N_549);
xnor U790 (N_790,N_50,N_447);
or U791 (N_791,N_305,N_557);
xnor U792 (N_792,N_680,N_236);
nor U793 (N_793,N_360,N_473);
nand U794 (N_794,N_608,N_177);
or U795 (N_795,N_295,N_498);
nand U796 (N_796,N_520,N_556);
or U797 (N_797,N_215,N_669);
nor U798 (N_798,N_464,N_471);
or U799 (N_799,N_676,N_54);
or U800 (N_800,N_408,N_643);
nand U801 (N_801,N_34,N_430);
nand U802 (N_802,N_626,N_170);
xnor U803 (N_803,N_732,N_470);
nand U804 (N_804,N_210,N_719);
or U805 (N_805,N_431,N_502);
nor U806 (N_806,N_261,N_654);
and U807 (N_807,N_224,N_235);
or U808 (N_808,N_673,N_93);
nor U809 (N_809,N_548,N_713);
and U810 (N_810,N_95,N_314);
and U811 (N_811,N_16,N_118);
and U812 (N_812,N_322,N_659);
or U813 (N_813,N_191,N_403);
nand U814 (N_814,N_695,N_615);
nand U815 (N_815,N_343,N_688);
nand U816 (N_816,N_485,N_272);
or U817 (N_817,N_0,N_237);
and U818 (N_818,N_53,N_559);
nor U819 (N_819,N_728,N_440);
xor U820 (N_820,N_287,N_749);
xor U821 (N_821,N_163,N_641);
xnor U822 (N_822,N_709,N_103);
nor U823 (N_823,N_479,N_513);
xor U824 (N_824,N_386,N_32);
nand U825 (N_825,N_397,N_745);
nor U826 (N_826,N_625,N_463);
nor U827 (N_827,N_655,N_365);
nor U828 (N_828,N_200,N_219);
xnor U829 (N_829,N_742,N_355);
xnor U830 (N_830,N_11,N_162);
xor U831 (N_831,N_636,N_467);
nor U832 (N_832,N_353,N_459);
nand U833 (N_833,N_73,N_122);
or U834 (N_834,N_727,N_185);
xnor U835 (N_835,N_414,N_211);
xor U836 (N_836,N_80,N_668);
and U837 (N_837,N_125,N_547);
and U838 (N_838,N_543,N_492);
nor U839 (N_839,N_566,N_230);
or U840 (N_840,N_715,N_29);
or U841 (N_841,N_370,N_40);
xnor U842 (N_842,N_509,N_279);
and U843 (N_843,N_746,N_285);
nor U844 (N_844,N_721,N_181);
nand U845 (N_845,N_5,N_26);
xnor U846 (N_846,N_681,N_229);
or U847 (N_847,N_602,N_493);
nor U848 (N_848,N_387,N_106);
nand U849 (N_849,N_197,N_631);
nor U850 (N_850,N_268,N_686);
nor U851 (N_851,N_17,N_300);
nor U852 (N_852,N_214,N_244);
or U853 (N_853,N_281,N_182);
or U854 (N_854,N_171,N_13);
xor U855 (N_855,N_270,N_363);
nor U856 (N_856,N_164,N_112);
or U857 (N_857,N_373,N_278);
nand U858 (N_858,N_76,N_640);
xor U859 (N_859,N_263,N_128);
nand U860 (N_860,N_642,N_666);
xor U861 (N_861,N_491,N_501);
and U862 (N_862,N_682,N_591);
nand U863 (N_863,N_685,N_420);
nand U864 (N_864,N_292,N_510);
or U865 (N_865,N_207,N_672);
nand U866 (N_866,N_569,N_358);
xor U867 (N_867,N_717,N_156);
or U868 (N_868,N_338,N_670);
or U869 (N_869,N_246,N_231);
nor U870 (N_870,N_97,N_739);
nand U871 (N_871,N_298,N_561);
nand U872 (N_872,N_108,N_716);
xor U873 (N_873,N_435,N_452);
or U874 (N_874,N_645,N_582);
nor U875 (N_875,N_500,N_544);
nor U876 (N_876,N_44,N_606);
nor U877 (N_877,N_89,N_316);
xor U878 (N_878,N_633,N_38);
or U879 (N_879,N_318,N_276);
or U880 (N_880,N_448,N_564);
xnor U881 (N_881,N_21,N_31);
nand U882 (N_882,N_528,N_743);
xor U883 (N_883,N_290,N_283);
and U884 (N_884,N_22,N_126);
nand U885 (N_885,N_346,N_161);
nand U886 (N_886,N_86,N_425);
nor U887 (N_887,N_489,N_653);
nor U888 (N_888,N_644,N_687);
xor U889 (N_889,N_710,N_540);
xor U890 (N_890,N_262,N_271);
nor U891 (N_891,N_45,N_184);
nor U892 (N_892,N_56,N_445);
nand U893 (N_893,N_587,N_329);
and U894 (N_894,N_136,N_41);
and U895 (N_895,N_454,N_109);
nor U896 (N_896,N_151,N_517);
nor U897 (N_897,N_351,N_427);
nand U898 (N_898,N_522,N_619);
xor U899 (N_899,N_506,N_368);
xor U900 (N_900,N_598,N_629);
nor U901 (N_901,N_9,N_658);
nor U902 (N_902,N_35,N_707);
nor U903 (N_903,N_726,N_260);
and U904 (N_904,N_172,N_736);
nor U905 (N_905,N_567,N_63);
or U906 (N_906,N_432,N_652);
xor U907 (N_907,N_534,N_24);
and U908 (N_908,N_66,N_7);
and U909 (N_909,N_132,N_442);
nor U910 (N_910,N_189,N_20);
nand U911 (N_911,N_226,N_451);
nand U912 (N_912,N_321,N_4);
or U913 (N_913,N_579,N_700);
or U914 (N_914,N_55,N_465);
or U915 (N_915,N_731,N_98);
and U916 (N_916,N_563,N_313);
nand U917 (N_917,N_42,N_698);
and U918 (N_918,N_328,N_304);
and U919 (N_919,N_59,N_434);
and U920 (N_920,N_124,N_206);
or U921 (N_921,N_497,N_538);
and U922 (N_922,N_597,N_293);
nor U923 (N_923,N_662,N_704);
nand U924 (N_924,N_390,N_15);
xnor U925 (N_925,N_198,N_428);
nand U926 (N_926,N_90,N_671);
nor U927 (N_927,N_33,N_192);
and U928 (N_928,N_637,N_458);
or U929 (N_929,N_352,N_649);
nor U930 (N_930,N_165,N_3);
or U931 (N_931,N_196,N_416);
and U932 (N_932,N_628,N_105);
xnor U933 (N_933,N_382,N_334);
xnor U934 (N_934,N_179,N_30);
or U935 (N_935,N_62,N_675);
nor U936 (N_936,N_296,N_12);
nand U937 (N_937,N_542,N_495);
and U938 (N_938,N_635,N_166);
nor U939 (N_939,N_515,N_616);
nor U940 (N_940,N_137,N_389);
and U941 (N_941,N_150,N_43);
nor U942 (N_942,N_180,N_741);
nor U943 (N_943,N_154,N_60);
or U944 (N_944,N_104,N_595);
or U945 (N_945,N_724,N_475);
nor U946 (N_946,N_696,N_74);
nand U947 (N_947,N_275,N_323);
nand U948 (N_948,N_404,N_536);
or U949 (N_949,N_371,N_570);
nand U950 (N_950,N_380,N_545);
nor U951 (N_951,N_332,N_552);
xor U952 (N_952,N_512,N_100);
xnor U953 (N_953,N_581,N_302);
nor U954 (N_954,N_663,N_496);
nor U955 (N_955,N_148,N_280);
and U956 (N_956,N_737,N_326);
xor U957 (N_957,N_450,N_578);
xor U958 (N_958,N_421,N_361);
or U959 (N_959,N_722,N_194);
nor U960 (N_960,N_508,N_665);
or U961 (N_961,N_315,N_610);
nor U962 (N_962,N_378,N_212);
and U963 (N_963,N_96,N_69);
nor U964 (N_964,N_324,N_601);
nor U965 (N_965,N_618,N_488);
nand U966 (N_966,N_306,N_584);
xnor U967 (N_967,N_466,N_594);
nand U968 (N_968,N_2,N_160);
or U969 (N_969,N_8,N_679);
xor U970 (N_970,N_350,N_411);
and U971 (N_971,N_560,N_381);
or U972 (N_972,N_516,N_577);
nor U973 (N_973,N_336,N_384);
nand U974 (N_974,N_257,N_460);
nor U975 (N_975,N_632,N_209);
nand U976 (N_976,N_222,N_599);
nand U977 (N_977,N_474,N_228);
xnor U978 (N_978,N_61,N_309);
or U979 (N_979,N_553,N_67);
nand U980 (N_980,N_469,N_396);
nand U981 (N_981,N_253,N_532);
and U982 (N_982,N_729,N_574);
and U983 (N_983,N_319,N_437);
xor U984 (N_984,N_269,N_521);
nand U985 (N_985,N_342,N_85);
or U986 (N_986,N_402,N_638);
nand U987 (N_987,N_691,N_72);
or U988 (N_988,N_273,N_550);
xor U989 (N_989,N_526,N_92);
or U990 (N_990,N_503,N_392);
or U991 (N_991,N_418,N_740);
and U992 (N_992,N_27,N_220);
nor U993 (N_993,N_505,N_701);
nand U994 (N_994,N_345,N_410);
and U995 (N_995,N_134,N_419);
and U996 (N_996,N_121,N_444);
xnor U997 (N_997,N_173,N_57);
nor U998 (N_998,N_504,N_167);
xnor U999 (N_999,N_75,N_223);
and U1000 (N_1000,N_277,N_49);
or U1001 (N_1001,N_590,N_247);
or U1002 (N_1002,N_650,N_284);
or U1003 (N_1003,N_580,N_720);
nor U1004 (N_1004,N_308,N_541);
nand U1005 (N_1005,N_39,N_58);
or U1006 (N_1006,N_449,N_183);
nor U1007 (N_1007,N_158,N_399);
xnor U1008 (N_1008,N_661,N_462);
and U1009 (N_1009,N_48,N_455);
or U1010 (N_1010,N_47,N_593);
nor U1011 (N_1011,N_169,N_81);
xor U1012 (N_1012,N_604,N_303);
nor U1013 (N_1013,N_99,N_115);
nor U1014 (N_1014,N_718,N_91);
and U1015 (N_1015,N_135,N_395);
nor U1016 (N_1016,N_530,N_195);
nand U1017 (N_1017,N_613,N_310);
or U1018 (N_1018,N_537,N_379);
xor U1019 (N_1019,N_249,N_630);
or U1020 (N_1020,N_357,N_611);
xnor U1021 (N_1021,N_562,N_110);
nand U1022 (N_1022,N_307,N_406);
nand U1023 (N_1023,N_400,N_187);
and U1024 (N_1024,N_483,N_347);
nand U1025 (N_1025,N_320,N_417);
nor U1026 (N_1026,N_130,N_605);
or U1027 (N_1027,N_401,N_693);
xnor U1028 (N_1028,N_592,N_193);
nand U1029 (N_1029,N_744,N_694);
xnor U1030 (N_1030,N_393,N_617);
and U1031 (N_1031,N_571,N_441);
or U1032 (N_1032,N_703,N_551);
nor U1033 (N_1033,N_71,N_176);
xnor U1034 (N_1034,N_714,N_486);
and U1035 (N_1035,N_364,N_678);
nor U1036 (N_1036,N_344,N_37);
nor U1037 (N_1037,N_119,N_639);
nor U1038 (N_1038,N_349,N_311);
nand U1039 (N_1039,N_107,N_286);
nor U1040 (N_1040,N_254,N_341);
nor U1041 (N_1041,N_239,N_433);
xnor U1042 (N_1042,N_461,N_114);
xnor U1043 (N_1043,N_117,N_554);
nor U1044 (N_1044,N_589,N_730);
and U1045 (N_1045,N_603,N_234);
nand U1046 (N_1046,N_238,N_201);
nand U1047 (N_1047,N_374,N_146);
xnor U1048 (N_1048,N_558,N_46);
and U1049 (N_1049,N_656,N_101);
nand U1050 (N_1050,N_409,N_439);
or U1051 (N_1051,N_199,N_359);
nand U1052 (N_1052,N_190,N_331);
xnor U1053 (N_1053,N_51,N_335);
nor U1054 (N_1054,N_407,N_648);
and U1055 (N_1055,N_65,N_241);
and U1056 (N_1056,N_494,N_573);
nand U1057 (N_1057,N_113,N_634);
or U1058 (N_1058,N_523,N_240);
xor U1059 (N_1059,N_186,N_267);
nor U1060 (N_1060,N_131,N_376);
xor U1061 (N_1061,N_294,N_348);
nand U1062 (N_1062,N_586,N_140);
and U1063 (N_1063,N_18,N_266);
xnor U1064 (N_1064,N_622,N_202);
or U1065 (N_1065,N_623,N_697);
and U1066 (N_1066,N_83,N_527);
or U1067 (N_1067,N_413,N_614);
and U1068 (N_1068,N_383,N_149);
nand U1069 (N_1069,N_216,N_394);
nor U1070 (N_1070,N_657,N_436);
nand U1071 (N_1071,N_144,N_531);
and U1072 (N_1072,N_233,N_25);
and U1073 (N_1073,N_10,N_291);
or U1074 (N_1074,N_289,N_747);
xor U1075 (N_1075,N_667,N_94);
nand U1076 (N_1076,N_68,N_36);
xor U1077 (N_1077,N_529,N_174);
nor U1078 (N_1078,N_367,N_265);
and U1079 (N_1079,N_225,N_583);
and U1080 (N_1080,N_138,N_535);
xor U1081 (N_1081,N_255,N_337);
or U1082 (N_1082,N_446,N_735);
xor U1083 (N_1083,N_168,N_533);
or U1084 (N_1084,N_443,N_481);
nor U1085 (N_1085,N_600,N_297);
or U1086 (N_1086,N_546,N_227);
xnor U1087 (N_1087,N_609,N_375);
or U1088 (N_1088,N_175,N_702);
nand U1089 (N_1089,N_699,N_325);
and U1090 (N_1090,N_514,N_689);
or U1091 (N_1091,N_301,N_208);
xor U1092 (N_1092,N_217,N_456);
nand U1093 (N_1093,N_28,N_218);
or U1094 (N_1094,N_116,N_507);
or U1095 (N_1095,N_288,N_23);
or U1096 (N_1096,N_607,N_424);
xnor U1097 (N_1097,N_78,N_499);
nor U1098 (N_1098,N_145,N_478);
or U1099 (N_1099,N_572,N_725);
nor U1100 (N_1100,N_438,N_157);
nor U1101 (N_1101,N_312,N_64);
nand U1102 (N_1102,N_539,N_205);
nor U1103 (N_1103,N_711,N_339);
and U1104 (N_1104,N_1,N_256);
nor U1105 (N_1105,N_457,N_153);
nor U1106 (N_1106,N_333,N_683);
or U1107 (N_1107,N_480,N_555);
or U1108 (N_1108,N_612,N_356);
and U1109 (N_1109,N_188,N_251);
and U1110 (N_1110,N_129,N_141);
nand U1111 (N_1111,N_677,N_748);
or U1112 (N_1112,N_405,N_525);
and U1113 (N_1113,N_723,N_692);
or U1114 (N_1114,N_624,N_366);
nor U1115 (N_1115,N_19,N_274);
xor U1116 (N_1116,N_674,N_575);
nor U1117 (N_1117,N_733,N_111);
xor U1118 (N_1118,N_52,N_660);
nand U1119 (N_1119,N_482,N_398);
xnor U1120 (N_1120,N_245,N_620);
or U1121 (N_1121,N_596,N_264);
xnor U1122 (N_1122,N_159,N_423);
or U1123 (N_1123,N_519,N_588);
and U1124 (N_1124,N_155,N_317);
or U1125 (N_1125,N_561,N_109);
or U1126 (N_1126,N_199,N_132);
and U1127 (N_1127,N_373,N_325);
nand U1128 (N_1128,N_564,N_203);
xor U1129 (N_1129,N_350,N_554);
xnor U1130 (N_1130,N_94,N_57);
or U1131 (N_1131,N_267,N_333);
xor U1132 (N_1132,N_735,N_699);
xnor U1133 (N_1133,N_236,N_18);
xor U1134 (N_1134,N_156,N_136);
xnor U1135 (N_1135,N_495,N_66);
nand U1136 (N_1136,N_525,N_194);
xor U1137 (N_1137,N_127,N_629);
nand U1138 (N_1138,N_507,N_748);
or U1139 (N_1139,N_258,N_583);
nand U1140 (N_1140,N_357,N_460);
or U1141 (N_1141,N_115,N_430);
xor U1142 (N_1142,N_630,N_200);
or U1143 (N_1143,N_574,N_619);
or U1144 (N_1144,N_522,N_66);
xor U1145 (N_1145,N_25,N_16);
and U1146 (N_1146,N_227,N_573);
nand U1147 (N_1147,N_264,N_179);
xor U1148 (N_1148,N_707,N_10);
and U1149 (N_1149,N_409,N_652);
nor U1150 (N_1150,N_326,N_498);
xnor U1151 (N_1151,N_588,N_412);
nor U1152 (N_1152,N_612,N_506);
or U1153 (N_1153,N_561,N_107);
nand U1154 (N_1154,N_638,N_27);
nand U1155 (N_1155,N_92,N_463);
nor U1156 (N_1156,N_394,N_736);
nor U1157 (N_1157,N_685,N_72);
or U1158 (N_1158,N_554,N_279);
xor U1159 (N_1159,N_98,N_106);
xnor U1160 (N_1160,N_545,N_108);
nand U1161 (N_1161,N_540,N_41);
xor U1162 (N_1162,N_91,N_206);
xnor U1163 (N_1163,N_603,N_382);
nor U1164 (N_1164,N_713,N_668);
and U1165 (N_1165,N_559,N_279);
nand U1166 (N_1166,N_543,N_72);
nand U1167 (N_1167,N_475,N_556);
nand U1168 (N_1168,N_366,N_28);
nor U1169 (N_1169,N_405,N_498);
and U1170 (N_1170,N_332,N_237);
and U1171 (N_1171,N_644,N_224);
and U1172 (N_1172,N_463,N_718);
nor U1173 (N_1173,N_90,N_559);
xor U1174 (N_1174,N_509,N_694);
nor U1175 (N_1175,N_218,N_208);
nand U1176 (N_1176,N_174,N_368);
nor U1177 (N_1177,N_572,N_117);
nand U1178 (N_1178,N_483,N_467);
and U1179 (N_1179,N_300,N_740);
nand U1180 (N_1180,N_673,N_508);
or U1181 (N_1181,N_741,N_386);
nor U1182 (N_1182,N_435,N_535);
or U1183 (N_1183,N_724,N_492);
or U1184 (N_1184,N_274,N_191);
or U1185 (N_1185,N_678,N_578);
or U1186 (N_1186,N_377,N_383);
or U1187 (N_1187,N_238,N_112);
nor U1188 (N_1188,N_318,N_735);
xor U1189 (N_1189,N_580,N_147);
nand U1190 (N_1190,N_565,N_206);
xnor U1191 (N_1191,N_692,N_18);
nand U1192 (N_1192,N_244,N_260);
nand U1193 (N_1193,N_33,N_357);
xnor U1194 (N_1194,N_37,N_11);
or U1195 (N_1195,N_160,N_303);
nand U1196 (N_1196,N_640,N_151);
nor U1197 (N_1197,N_376,N_77);
nor U1198 (N_1198,N_254,N_553);
xnor U1199 (N_1199,N_669,N_564);
nor U1200 (N_1200,N_502,N_746);
or U1201 (N_1201,N_38,N_255);
nand U1202 (N_1202,N_21,N_290);
and U1203 (N_1203,N_365,N_0);
xor U1204 (N_1204,N_706,N_559);
nor U1205 (N_1205,N_14,N_563);
and U1206 (N_1206,N_453,N_367);
nand U1207 (N_1207,N_596,N_446);
xor U1208 (N_1208,N_352,N_695);
nor U1209 (N_1209,N_315,N_18);
xor U1210 (N_1210,N_420,N_478);
xnor U1211 (N_1211,N_160,N_191);
xor U1212 (N_1212,N_128,N_717);
nand U1213 (N_1213,N_437,N_200);
nand U1214 (N_1214,N_174,N_592);
xnor U1215 (N_1215,N_693,N_606);
or U1216 (N_1216,N_335,N_571);
nand U1217 (N_1217,N_0,N_270);
or U1218 (N_1218,N_13,N_125);
nand U1219 (N_1219,N_661,N_79);
nand U1220 (N_1220,N_622,N_608);
and U1221 (N_1221,N_495,N_133);
nor U1222 (N_1222,N_209,N_420);
and U1223 (N_1223,N_170,N_722);
nor U1224 (N_1224,N_295,N_478);
and U1225 (N_1225,N_664,N_577);
and U1226 (N_1226,N_473,N_652);
and U1227 (N_1227,N_425,N_721);
xor U1228 (N_1228,N_566,N_658);
or U1229 (N_1229,N_67,N_429);
and U1230 (N_1230,N_77,N_151);
xor U1231 (N_1231,N_523,N_148);
or U1232 (N_1232,N_313,N_525);
and U1233 (N_1233,N_245,N_449);
xnor U1234 (N_1234,N_365,N_704);
and U1235 (N_1235,N_349,N_479);
nand U1236 (N_1236,N_356,N_493);
and U1237 (N_1237,N_430,N_745);
nor U1238 (N_1238,N_326,N_193);
xnor U1239 (N_1239,N_225,N_695);
nor U1240 (N_1240,N_716,N_158);
or U1241 (N_1241,N_519,N_340);
xor U1242 (N_1242,N_324,N_351);
nand U1243 (N_1243,N_505,N_680);
nor U1244 (N_1244,N_604,N_509);
nor U1245 (N_1245,N_206,N_695);
nor U1246 (N_1246,N_274,N_413);
and U1247 (N_1247,N_58,N_597);
nand U1248 (N_1248,N_725,N_418);
xor U1249 (N_1249,N_508,N_605);
and U1250 (N_1250,N_216,N_203);
nand U1251 (N_1251,N_209,N_227);
xnor U1252 (N_1252,N_67,N_724);
and U1253 (N_1253,N_333,N_295);
nand U1254 (N_1254,N_111,N_458);
nor U1255 (N_1255,N_148,N_98);
and U1256 (N_1256,N_280,N_185);
and U1257 (N_1257,N_587,N_482);
and U1258 (N_1258,N_690,N_298);
and U1259 (N_1259,N_602,N_363);
nand U1260 (N_1260,N_165,N_299);
xnor U1261 (N_1261,N_178,N_518);
xnor U1262 (N_1262,N_378,N_510);
or U1263 (N_1263,N_615,N_515);
nand U1264 (N_1264,N_519,N_197);
xor U1265 (N_1265,N_455,N_40);
nor U1266 (N_1266,N_185,N_204);
xnor U1267 (N_1267,N_55,N_299);
nor U1268 (N_1268,N_392,N_466);
and U1269 (N_1269,N_189,N_250);
xor U1270 (N_1270,N_717,N_541);
or U1271 (N_1271,N_603,N_650);
nand U1272 (N_1272,N_191,N_701);
or U1273 (N_1273,N_127,N_352);
and U1274 (N_1274,N_443,N_665);
nor U1275 (N_1275,N_129,N_679);
or U1276 (N_1276,N_152,N_724);
nor U1277 (N_1277,N_417,N_351);
and U1278 (N_1278,N_361,N_211);
nand U1279 (N_1279,N_693,N_613);
xor U1280 (N_1280,N_83,N_713);
and U1281 (N_1281,N_302,N_255);
and U1282 (N_1282,N_211,N_18);
nand U1283 (N_1283,N_223,N_200);
nand U1284 (N_1284,N_147,N_214);
nand U1285 (N_1285,N_375,N_64);
or U1286 (N_1286,N_369,N_109);
xnor U1287 (N_1287,N_282,N_96);
nor U1288 (N_1288,N_355,N_401);
nand U1289 (N_1289,N_186,N_535);
nor U1290 (N_1290,N_125,N_688);
nor U1291 (N_1291,N_67,N_592);
nor U1292 (N_1292,N_642,N_709);
and U1293 (N_1293,N_531,N_522);
nor U1294 (N_1294,N_337,N_498);
nor U1295 (N_1295,N_326,N_725);
nand U1296 (N_1296,N_673,N_510);
or U1297 (N_1297,N_524,N_734);
or U1298 (N_1298,N_239,N_503);
or U1299 (N_1299,N_470,N_232);
xor U1300 (N_1300,N_30,N_611);
nor U1301 (N_1301,N_655,N_193);
xor U1302 (N_1302,N_728,N_685);
xnor U1303 (N_1303,N_334,N_541);
xor U1304 (N_1304,N_228,N_245);
or U1305 (N_1305,N_517,N_525);
nor U1306 (N_1306,N_458,N_266);
nor U1307 (N_1307,N_24,N_443);
or U1308 (N_1308,N_713,N_15);
and U1309 (N_1309,N_487,N_306);
nand U1310 (N_1310,N_144,N_634);
and U1311 (N_1311,N_154,N_624);
and U1312 (N_1312,N_523,N_238);
nand U1313 (N_1313,N_295,N_599);
or U1314 (N_1314,N_234,N_540);
or U1315 (N_1315,N_542,N_72);
or U1316 (N_1316,N_215,N_679);
or U1317 (N_1317,N_504,N_319);
xor U1318 (N_1318,N_461,N_85);
or U1319 (N_1319,N_335,N_708);
nand U1320 (N_1320,N_648,N_469);
nor U1321 (N_1321,N_34,N_549);
nor U1322 (N_1322,N_275,N_736);
xor U1323 (N_1323,N_596,N_120);
and U1324 (N_1324,N_95,N_220);
nand U1325 (N_1325,N_392,N_144);
nand U1326 (N_1326,N_192,N_366);
xnor U1327 (N_1327,N_143,N_696);
nor U1328 (N_1328,N_101,N_718);
or U1329 (N_1329,N_9,N_93);
xnor U1330 (N_1330,N_16,N_243);
nand U1331 (N_1331,N_252,N_350);
nor U1332 (N_1332,N_129,N_588);
xnor U1333 (N_1333,N_239,N_241);
or U1334 (N_1334,N_231,N_127);
and U1335 (N_1335,N_95,N_355);
or U1336 (N_1336,N_642,N_66);
nand U1337 (N_1337,N_72,N_301);
nand U1338 (N_1338,N_380,N_178);
nor U1339 (N_1339,N_200,N_220);
and U1340 (N_1340,N_461,N_744);
or U1341 (N_1341,N_407,N_568);
nor U1342 (N_1342,N_236,N_176);
xor U1343 (N_1343,N_452,N_138);
nor U1344 (N_1344,N_56,N_628);
or U1345 (N_1345,N_222,N_200);
and U1346 (N_1346,N_705,N_171);
xor U1347 (N_1347,N_269,N_499);
or U1348 (N_1348,N_377,N_421);
or U1349 (N_1349,N_205,N_255);
xor U1350 (N_1350,N_50,N_407);
xor U1351 (N_1351,N_159,N_121);
or U1352 (N_1352,N_644,N_414);
xor U1353 (N_1353,N_193,N_170);
and U1354 (N_1354,N_205,N_613);
xnor U1355 (N_1355,N_454,N_232);
and U1356 (N_1356,N_283,N_147);
and U1357 (N_1357,N_410,N_655);
nand U1358 (N_1358,N_439,N_490);
xor U1359 (N_1359,N_619,N_370);
or U1360 (N_1360,N_621,N_667);
or U1361 (N_1361,N_177,N_203);
or U1362 (N_1362,N_405,N_582);
xor U1363 (N_1363,N_681,N_84);
xnor U1364 (N_1364,N_572,N_310);
nor U1365 (N_1365,N_290,N_418);
xor U1366 (N_1366,N_9,N_362);
nor U1367 (N_1367,N_474,N_451);
or U1368 (N_1368,N_441,N_90);
nor U1369 (N_1369,N_273,N_606);
nor U1370 (N_1370,N_18,N_685);
or U1371 (N_1371,N_108,N_150);
nand U1372 (N_1372,N_702,N_202);
nor U1373 (N_1373,N_195,N_383);
xor U1374 (N_1374,N_718,N_210);
xor U1375 (N_1375,N_323,N_518);
and U1376 (N_1376,N_475,N_123);
nand U1377 (N_1377,N_535,N_264);
nand U1378 (N_1378,N_283,N_379);
nand U1379 (N_1379,N_199,N_451);
or U1380 (N_1380,N_8,N_144);
nand U1381 (N_1381,N_57,N_270);
or U1382 (N_1382,N_668,N_83);
nand U1383 (N_1383,N_405,N_14);
xor U1384 (N_1384,N_324,N_90);
and U1385 (N_1385,N_552,N_51);
xor U1386 (N_1386,N_491,N_558);
xor U1387 (N_1387,N_584,N_107);
and U1388 (N_1388,N_534,N_274);
nor U1389 (N_1389,N_616,N_619);
nand U1390 (N_1390,N_308,N_621);
nand U1391 (N_1391,N_514,N_34);
nor U1392 (N_1392,N_64,N_671);
xor U1393 (N_1393,N_135,N_184);
xnor U1394 (N_1394,N_721,N_491);
or U1395 (N_1395,N_502,N_234);
xnor U1396 (N_1396,N_342,N_263);
or U1397 (N_1397,N_435,N_245);
nand U1398 (N_1398,N_244,N_380);
xnor U1399 (N_1399,N_659,N_78);
and U1400 (N_1400,N_73,N_375);
and U1401 (N_1401,N_111,N_52);
or U1402 (N_1402,N_202,N_64);
or U1403 (N_1403,N_214,N_241);
or U1404 (N_1404,N_273,N_636);
xor U1405 (N_1405,N_747,N_566);
nor U1406 (N_1406,N_332,N_235);
xnor U1407 (N_1407,N_426,N_547);
and U1408 (N_1408,N_470,N_509);
and U1409 (N_1409,N_658,N_175);
nor U1410 (N_1410,N_205,N_399);
xnor U1411 (N_1411,N_211,N_587);
nand U1412 (N_1412,N_572,N_614);
and U1413 (N_1413,N_565,N_697);
nor U1414 (N_1414,N_713,N_584);
or U1415 (N_1415,N_695,N_209);
nor U1416 (N_1416,N_206,N_448);
or U1417 (N_1417,N_707,N_598);
nand U1418 (N_1418,N_418,N_362);
or U1419 (N_1419,N_14,N_415);
nand U1420 (N_1420,N_158,N_415);
xor U1421 (N_1421,N_386,N_725);
nor U1422 (N_1422,N_613,N_687);
nor U1423 (N_1423,N_83,N_745);
xor U1424 (N_1424,N_218,N_284);
and U1425 (N_1425,N_721,N_300);
or U1426 (N_1426,N_29,N_443);
or U1427 (N_1427,N_568,N_525);
nand U1428 (N_1428,N_303,N_612);
nand U1429 (N_1429,N_305,N_418);
nor U1430 (N_1430,N_210,N_29);
xor U1431 (N_1431,N_8,N_496);
or U1432 (N_1432,N_274,N_151);
and U1433 (N_1433,N_318,N_288);
or U1434 (N_1434,N_474,N_157);
nand U1435 (N_1435,N_420,N_268);
nor U1436 (N_1436,N_543,N_315);
xor U1437 (N_1437,N_698,N_224);
and U1438 (N_1438,N_475,N_8);
and U1439 (N_1439,N_631,N_36);
nor U1440 (N_1440,N_37,N_607);
or U1441 (N_1441,N_476,N_513);
nor U1442 (N_1442,N_5,N_13);
nor U1443 (N_1443,N_20,N_248);
nor U1444 (N_1444,N_72,N_716);
nand U1445 (N_1445,N_209,N_593);
nand U1446 (N_1446,N_501,N_197);
nand U1447 (N_1447,N_78,N_283);
or U1448 (N_1448,N_30,N_95);
nor U1449 (N_1449,N_680,N_89);
xnor U1450 (N_1450,N_414,N_395);
nor U1451 (N_1451,N_517,N_203);
nand U1452 (N_1452,N_114,N_719);
xor U1453 (N_1453,N_69,N_343);
xor U1454 (N_1454,N_577,N_728);
xnor U1455 (N_1455,N_366,N_293);
xor U1456 (N_1456,N_536,N_410);
nor U1457 (N_1457,N_62,N_101);
and U1458 (N_1458,N_361,N_171);
nand U1459 (N_1459,N_361,N_29);
and U1460 (N_1460,N_205,N_516);
or U1461 (N_1461,N_458,N_57);
nand U1462 (N_1462,N_579,N_267);
nor U1463 (N_1463,N_532,N_536);
nand U1464 (N_1464,N_258,N_592);
or U1465 (N_1465,N_393,N_414);
nor U1466 (N_1466,N_654,N_376);
nand U1467 (N_1467,N_358,N_698);
nor U1468 (N_1468,N_650,N_137);
xnor U1469 (N_1469,N_485,N_472);
or U1470 (N_1470,N_175,N_279);
xor U1471 (N_1471,N_500,N_303);
or U1472 (N_1472,N_99,N_20);
or U1473 (N_1473,N_179,N_207);
and U1474 (N_1474,N_412,N_657);
xnor U1475 (N_1475,N_606,N_290);
nor U1476 (N_1476,N_311,N_262);
nor U1477 (N_1477,N_477,N_300);
nand U1478 (N_1478,N_175,N_682);
nand U1479 (N_1479,N_215,N_449);
nor U1480 (N_1480,N_590,N_329);
and U1481 (N_1481,N_323,N_628);
nor U1482 (N_1482,N_44,N_107);
nand U1483 (N_1483,N_93,N_315);
or U1484 (N_1484,N_70,N_656);
and U1485 (N_1485,N_394,N_48);
nand U1486 (N_1486,N_60,N_705);
or U1487 (N_1487,N_240,N_326);
nor U1488 (N_1488,N_723,N_713);
nor U1489 (N_1489,N_506,N_512);
and U1490 (N_1490,N_559,N_521);
or U1491 (N_1491,N_261,N_553);
or U1492 (N_1492,N_230,N_433);
or U1493 (N_1493,N_154,N_1);
nor U1494 (N_1494,N_698,N_133);
xnor U1495 (N_1495,N_701,N_714);
or U1496 (N_1496,N_116,N_494);
xnor U1497 (N_1497,N_718,N_287);
nand U1498 (N_1498,N_96,N_313);
nor U1499 (N_1499,N_51,N_237);
or U1500 (N_1500,N_1373,N_867);
and U1501 (N_1501,N_984,N_831);
nor U1502 (N_1502,N_1401,N_1491);
and U1503 (N_1503,N_1386,N_952);
and U1504 (N_1504,N_1423,N_1467);
nor U1505 (N_1505,N_1322,N_1025);
nor U1506 (N_1506,N_1324,N_1437);
nand U1507 (N_1507,N_1361,N_1457);
and U1508 (N_1508,N_1033,N_752);
or U1509 (N_1509,N_971,N_1047);
nor U1510 (N_1510,N_1140,N_1421);
xor U1511 (N_1511,N_1416,N_945);
nand U1512 (N_1512,N_1405,N_1382);
nand U1513 (N_1513,N_1155,N_1282);
xnor U1514 (N_1514,N_1428,N_1489);
nor U1515 (N_1515,N_1399,N_1352);
nor U1516 (N_1516,N_947,N_1188);
or U1517 (N_1517,N_1366,N_1003);
nor U1518 (N_1518,N_1359,N_1240);
xnor U1519 (N_1519,N_1223,N_1376);
nand U1520 (N_1520,N_1000,N_1079);
and U1521 (N_1521,N_1023,N_1292);
xnor U1522 (N_1522,N_1090,N_803);
nor U1523 (N_1523,N_785,N_1124);
and U1524 (N_1524,N_1462,N_974);
xor U1525 (N_1525,N_1314,N_859);
and U1526 (N_1526,N_929,N_1184);
nand U1527 (N_1527,N_1161,N_758);
xor U1528 (N_1528,N_1144,N_772);
and U1529 (N_1529,N_1302,N_1492);
nand U1530 (N_1530,N_1368,N_1127);
and U1531 (N_1531,N_1160,N_812);
or U1532 (N_1532,N_987,N_1348);
nand U1533 (N_1533,N_1358,N_1378);
or U1534 (N_1534,N_896,N_1259);
nor U1535 (N_1535,N_855,N_754);
nor U1536 (N_1536,N_1443,N_1414);
nand U1537 (N_1537,N_1007,N_1305);
xor U1538 (N_1538,N_1430,N_1083);
and U1539 (N_1539,N_1107,N_1189);
and U1540 (N_1540,N_1284,N_1122);
and U1541 (N_1541,N_900,N_1479);
nor U1542 (N_1542,N_1211,N_1114);
xor U1543 (N_1543,N_798,N_783);
and U1544 (N_1544,N_775,N_1315);
or U1545 (N_1545,N_1167,N_765);
nor U1546 (N_1546,N_759,N_1431);
xnor U1547 (N_1547,N_1283,N_1029);
and U1548 (N_1548,N_790,N_903);
xnor U1549 (N_1549,N_1463,N_1228);
nor U1550 (N_1550,N_1334,N_1235);
nor U1551 (N_1551,N_1118,N_1388);
xor U1552 (N_1552,N_982,N_1233);
or U1553 (N_1553,N_981,N_941);
or U1554 (N_1554,N_1438,N_1449);
xnor U1555 (N_1555,N_916,N_934);
or U1556 (N_1556,N_1295,N_1032);
nand U1557 (N_1557,N_930,N_1065);
and U1558 (N_1558,N_1207,N_1060);
nor U1559 (N_1559,N_1180,N_1193);
nand U1560 (N_1560,N_1277,N_902);
or U1561 (N_1561,N_1187,N_1267);
nand U1562 (N_1562,N_977,N_1218);
and U1563 (N_1563,N_1464,N_1304);
nor U1564 (N_1564,N_1174,N_849);
or U1565 (N_1565,N_1012,N_860);
or U1566 (N_1566,N_826,N_865);
nor U1567 (N_1567,N_1054,N_1084);
and U1568 (N_1568,N_893,N_968);
nand U1569 (N_1569,N_1372,N_1126);
nor U1570 (N_1570,N_1097,N_781);
and U1571 (N_1571,N_1196,N_764);
nand U1572 (N_1572,N_1362,N_773);
xor U1573 (N_1573,N_1450,N_850);
xnor U1574 (N_1574,N_1141,N_802);
and U1575 (N_1575,N_906,N_1460);
nand U1576 (N_1576,N_852,N_1156);
nor U1577 (N_1577,N_1119,N_887);
or U1578 (N_1578,N_1128,N_1459);
nand U1579 (N_1579,N_1063,N_1338);
and U1580 (N_1580,N_960,N_787);
xnor U1581 (N_1581,N_797,N_1471);
nand U1582 (N_1582,N_1293,N_1070);
and U1583 (N_1583,N_1015,N_811);
and U1584 (N_1584,N_1075,N_875);
or U1585 (N_1585,N_1204,N_805);
nor U1586 (N_1586,N_872,N_1006);
nand U1587 (N_1587,N_1487,N_1321);
xnor U1588 (N_1588,N_793,N_1016);
or U1589 (N_1589,N_1266,N_1076);
or U1590 (N_1590,N_1275,N_961);
nor U1591 (N_1591,N_1274,N_1036);
and U1592 (N_1592,N_993,N_931);
nor U1593 (N_1593,N_1152,N_1225);
and U1594 (N_1594,N_1357,N_975);
or U1595 (N_1595,N_925,N_1364);
and U1596 (N_1596,N_776,N_1417);
xor U1597 (N_1597,N_1498,N_1476);
nor U1598 (N_1598,N_1175,N_1085);
nand U1599 (N_1599,N_813,N_1485);
nor U1600 (N_1600,N_923,N_878);
xnor U1601 (N_1601,N_766,N_1415);
and U1602 (N_1602,N_1289,N_1468);
nor U1603 (N_1603,N_1093,N_1387);
or U1604 (N_1604,N_1385,N_840);
nor U1605 (N_1605,N_1280,N_1086);
nand U1606 (N_1606,N_1217,N_1342);
nand U1607 (N_1607,N_1116,N_1213);
nor U1608 (N_1608,N_914,N_1360);
nor U1609 (N_1609,N_908,N_963);
or U1610 (N_1610,N_1080,N_1209);
nor U1611 (N_1611,N_970,N_922);
nor U1612 (N_1612,N_949,N_1406);
xnor U1613 (N_1613,N_1202,N_1030);
and U1614 (N_1614,N_1397,N_842);
xnor U1615 (N_1615,N_763,N_774);
and U1616 (N_1616,N_1291,N_864);
xnor U1617 (N_1617,N_901,N_964);
nor U1618 (N_1618,N_1044,N_1465);
and U1619 (N_1619,N_1215,N_834);
nor U1620 (N_1620,N_841,N_1276);
nand U1621 (N_1621,N_1154,N_1129);
nand U1622 (N_1622,N_814,N_898);
nand U1623 (N_1623,N_1216,N_1336);
or U1624 (N_1624,N_1299,N_913);
xnor U1625 (N_1625,N_1453,N_1339);
nand U1626 (N_1626,N_1017,N_816);
nand U1627 (N_1627,N_1192,N_1432);
or U1628 (N_1628,N_1271,N_830);
nand U1629 (N_1629,N_991,N_801);
xor U1630 (N_1630,N_924,N_1045);
or U1631 (N_1631,N_1197,N_1311);
or U1632 (N_1632,N_1312,N_762);
nand U1633 (N_1633,N_1263,N_1384);
nand U1634 (N_1634,N_1191,N_1363);
nand U1635 (N_1635,N_1481,N_897);
nand U1636 (N_1636,N_1260,N_869);
or U1637 (N_1637,N_936,N_1350);
nand U1638 (N_1638,N_1490,N_1182);
and U1639 (N_1639,N_1049,N_835);
and U1640 (N_1640,N_1057,N_881);
xnor U1641 (N_1641,N_1108,N_780);
xnor U1642 (N_1642,N_989,N_1112);
nor U1643 (N_1643,N_967,N_1345);
or U1644 (N_1644,N_1496,N_804);
nand U1645 (N_1645,N_1374,N_933);
xor U1646 (N_1646,N_1001,N_1037);
nor U1647 (N_1647,N_810,N_895);
xnor U1648 (N_1648,N_825,N_771);
and U1649 (N_1649,N_1461,N_1330);
nand U1650 (N_1650,N_1138,N_1246);
xnor U1651 (N_1651,N_862,N_1480);
xnor U1652 (N_1652,N_1400,N_1328);
and U1653 (N_1653,N_938,N_1447);
nand U1654 (N_1654,N_796,N_1046);
or U1655 (N_1655,N_1026,N_1418);
nor U1656 (N_1656,N_777,N_1199);
nor U1657 (N_1657,N_1190,N_1035);
xor U1658 (N_1658,N_817,N_1021);
nand U1659 (N_1659,N_823,N_980);
or U1660 (N_1660,N_1488,N_1041);
nor U1661 (N_1661,N_1176,N_1102);
or U1662 (N_1662,N_1148,N_1226);
nand U1663 (N_1663,N_1043,N_828);
or U1664 (N_1664,N_1059,N_1261);
xor U1665 (N_1665,N_1482,N_1310);
nand U1666 (N_1666,N_1194,N_1168);
xnor U1667 (N_1667,N_1137,N_808);
nand U1668 (N_1668,N_1031,N_1436);
nor U1669 (N_1669,N_1227,N_1142);
or U1670 (N_1670,N_1343,N_1278);
and U1671 (N_1671,N_1092,N_789);
and U1672 (N_1672,N_1494,N_1071);
nor U1673 (N_1673,N_876,N_845);
and U1674 (N_1674,N_1326,N_1200);
or U1675 (N_1675,N_959,N_1153);
nor U1676 (N_1676,N_1214,N_1183);
and U1677 (N_1677,N_1420,N_809);
and U1678 (N_1678,N_1206,N_919);
xnor U1679 (N_1679,N_1281,N_1178);
or U1680 (N_1680,N_969,N_1301);
xnor U1681 (N_1681,N_1028,N_1120);
nand U1682 (N_1682,N_1377,N_951);
or U1683 (N_1683,N_909,N_996);
nor U1684 (N_1684,N_1493,N_770);
nand U1685 (N_1685,N_939,N_1087);
xnor U1686 (N_1686,N_1484,N_1323);
nand U1687 (N_1687,N_853,N_1195);
or U1688 (N_1688,N_944,N_1354);
and U1689 (N_1689,N_1444,N_753);
or U1690 (N_1690,N_1270,N_1151);
nand U1691 (N_1691,N_833,N_1058);
nor U1692 (N_1692,N_1410,N_932);
nor U1693 (N_1693,N_985,N_1300);
or U1694 (N_1694,N_829,N_761);
or U1695 (N_1695,N_1327,N_1099);
or U1696 (N_1696,N_844,N_1356);
or U1697 (N_1697,N_904,N_954);
xor U1698 (N_1698,N_1051,N_1146);
or U1699 (N_1699,N_751,N_1298);
and U1700 (N_1700,N_994,N_1210);
nor U1701 (N_1701,N_778,N_1150);
or U1702 (N_1702,N_858,N_784);
and U1703 (N_1703,N_1177,N_915);
nor U1704 (N_1704,N_948,N_1470);
or U1705 (N_1705,N_1091,N_958);
xor U1706 (N_1706,N_1157,N_1332);
or U1707 (N_1707,N_1239,N_1222);
xor U1708 (N_1708,N_1212,N_1448);
nand U1709 (N_1709,N_1318,N_1011);
and U1710 (N_1710,N_1136,N_1344);
or U1711 (N_1711,N_1412,N_1313);
or U1712 (N_1712,N_1367,N_1268);
or U1713 (N_1713,N_827,N_978);
and U1714 (N_1714,N_979,N_1307);
or U1715 (N_1715,N_1411,N_1486);
or U1716 (N_1716,N_1383,N_1117);
nor U1717 (N_1717,N_1433,N_1139);
and U1718 (N_1718,N_894,N_1251);
xor U1719 (N_1719,N_1455,N_1098);
xnor U1720 (N_1720,N_846,N_1048);
xnor U1721 (N_1721,N_1115,N_750);
and U1722 (N_1722,N_799,N_1395);
and U1723 (N_1723,N_873,N_822);
nand U1724 (N_1724,N_1186,N_966);
xor U1725 (N_1725,N_1288,N_1434);
and U1726 (N_1726,N_863,N_1052);
xnor U1727 (N_1727,N_868,N_1252);
nor U1728 (N_1728,N_866,N_917);
or U1729 (N_1729,N_946,N_1133);
or U1730 (N_1730,N_1454,N_943);
or U1731 (N_1731,N_1095,N_836);
and U1732 (N_1732,N_1101,N_1103);
or U1733 (N_1733,N_1181,N_1230);
or U1734 (N_1734,N_1243,N_911);
and U1735 (N_1735,N_1381,N_1064);
xnor U1736 (N_1736,N_767,N_1004);
and U1737 (N_1737,N_819,N_1069);
xor U1738 (N_1738,N_1403,N_1340);
nor U1739 (N_1739,N_1205,N_1452);
nand U1740 (N_1740,N_1309,N_888);
and U1741 (N_1741,N_1053,N_905);
nand U1742 (N_1742,N_1072,N_884);
nand U1743 (N_1743,N_1391,N_1375);
nor U1744 (N_1744,N_1237,N_882);
nand U1745 (N_1745,N_1143,N_1077);
and U1746 (N_1746,N_1149,N_768);
xor U1747 (N_1747,N_965,N_1249);
xnor U1748 (N_1748,N_1169,N_1242);
nand U1749 (N_1749,N_973,N_1123);
xor U1750 (N_1750,N_1074,N_1179);
nor U1751 (N_1751,N_1427,N_992);
or U1752 (N_1752,N_1408,N_1113);
nor U1753 (N_1753,N_1220,N_1171);
or U1754 (N_1754,N_1273,N_1134);
nand U1755 (N_1755,N_1472,N_920);
nor U1756 (N_1756,N_891,N_1499);
xnor U1757 (N_1757,N_857,N_856);
and U1758 (N_1758,N_1287,N_1020);
and U1759 (N_1759,N_1125,N_1066);
or U1760 (N_1760,N_1008,N_794);
and U1761 (N_1761,N_1018,N_1475);
or U1762 (N_1762,N_818,N_1407);
nor U1763 (N_1763,N_1005,N_1166);
nor U1764 (N_1764,N_1351,N_1474);
nor U1765 (N_1765,N_1050,N_1042);
or U1766 (N_1766,N_1390,N_847);
or U1767 (N_1767,N_986,N_815);
nor U1768 (N_1768,N_1346,N_1265);
xor U1769 (N_1769,N_1104,N_1389);
or U1770 (N_1770,N_1068,N_1078);
and U1771 (N_1771,N_861,N_1320);
and U1772 (N_1772,N_1040,N_1473);
or U1773 (N_1773,N_1337,N_927);
nor U1774 (N_1774,N_972,N_1162);
and U1775 (N_1775,N_1130,N_1147);
xor U1776 (N_1776,N_779,N_1442);
xor U1777 (N_1777,N_1105,N_760);
xor U1778 (N_1778,N_1371,N_883);
or U1779 (N_1779,N_1317,N_1100);
nand U1780 (N_1780,N_1290,N_1425);
and U1781 (N_1781,N_880,N_1445);
nor U1782 (N_1782,N_1446,N_1306);
nor U1783 (N_1783,N_1329,N_1229);
xor U1784 (N_1784,N_955,N_1109);
xnor U1785 (N_1785,N_782,N_871);
or U1786 (N_1786,N_889,N_892);
or U1787 (N_1787,N_1316,N_1440);
nand U1788 (N_1788,N_1254,N_890);
and U1789 (N_1789,N_824,N_1231);
or U1790 (N_1790,N_1341,N_937);
and U1791 (N_1791,N_843,N_1296);
xnor U1792 (N_1792,N_839,N_1398);
and U1793 (N_1793,N_1279,N_1034);
or U1794 (N_1794,N_1014,N_1495);
nand U1795 (N_1795,N_1335,N_1219);
xnor U1796 (N_1796,N_1250,N_997);
and U1797 (N_1797,N_1294,N_899);
or U1798 (N_1798,N_1185,N_998);
or U1799 (N_1799,N_1081,N_1253);
and U1800 (N_1800,N_1286,N_1247);
or U1801 (N_1801,N_928,N_1419);
nand U1802 (N_1802,N_1232,N_1198);
and U1803 (N_1803,N_1145,N_1402);
or U1804 (N_1804,N_792,N_807);
or U1805 (N_1805,N_1404,N_1435);
or U1806 (N_1806,N_1055,N_886);
nor U1807 (N_1807,N_1257,N_942);
or U1808 (N_1808,N_821,N_854);
nor U1809 (N_1809,N_1458,N_1027);
xor U1810 (N_1810,N_1413,N_1002);
xor U1811 (N_1811,N_1308,N_1221);
nor U1812 (N_1812,N_988,N_1456);
xor U1813 (N_1813,N_1347,N_976);
nand U1814 (N_1814,N_1319,N_1038);
nor U1815 (N_1815,N_837,N_1477);
and U1816 (N_1816,N_806,N_1164);
and U1817 (N_1817,N_877,N_1325);
or U1818 (N_1818,N_874,N_1245);
nand U1819 (N_1819,N_1241,N_910);
xnor U1820 (N_1820,N_1441,N_1067);
nor U1821 (N_1821,N_795,N_1089);
nand U1822 (N_1822,N_1061,N_950);
nor U1823 (N_1823,N_1234,N_957);
and U1824 (N_1824,N_832,N_755);
and U1825 (N_1825,N_1082,N_1497);
and U1826 (N_1826,N_956,N_1135);
xor U1827 (N_1827,N_1062,N_1173);
and U1828 (N_1828,N_1285,N_788);
nand U1829 (N_1829,N_1172,N_1096);
nand U1830 (N_1830,N_1262,N_1370);
xor U1831 (N_1831,N_1158,N_1170);
or U1832 (N_1832,N_1422,N_1478);
or U1833 (N_1833,N_1369,N_1396);
xnor U1834 (N_1834,N_1256,N_1426);
nor U1835 (N_1835,N_1303,N_1073);
nor U1836 (N_1836,N_1469,N_1258);
and U1837 (N_1837,N_1236,N_1244);
xnor U1838 (N_1838,N_1269,N_1165);
xnor U1839 (N_1839,N_1451,N_907);
xnor U1840 (N_1840,N_879,N_786);
or U1841 (N_1841,N_953,N_1365);
and U1842 (N_1842,N_848,N_935);
nor U1843 (N_1843,N_1238,N_1392);
xnor U1844 (N_1844,N_1224,N_1110);
nand U1845 (N_1845,N_940,N_1394);
xor U1846 (N_1846,N_1379,N_851);
nand U1847 (N_1847,N_1039,N_1333);
nand U1848 (N_1848,N_1131,N_820);
nor U1849 (N_1849,N_1163,N_1264);
and U1850 (N_1850,N_1393,N_1056);
and U1851 (N_1851,N_1022,N_1409);
or U1852 (N_1852,N_1439,N_1208);
xnor U1853 (N_1853,N_1349,N_1331);
nand U1854 (N_1854,N_1019,N_1010);
nor U1855 (N_1855,N_1121,N_962);
or U1856 (N_1856,N_1380,N_1429);
nor U1857 (N_1857,N_1297,N_995);
nand U1858 (N_1858,N_999,N_918);
nand U1859 (N_1859,N_870,N_1111);
nand U1860 (N_1860,N_1424,N_1088);
and U1861 (N_1861,N_1203,N_921);
nand U1862 (N_1862,N_1483,N_1009);
and U1863 (N_1863,N_1013,N_1201);
or U1864 (N_1864,N_1132,N_1353);
or U1865 (N_1865,N_990,N_1024);
and U1866 (N_1866,N_885,N_757);
or U1867 (N_1867,N_769,N_926);
and U1868 (N_1868,N_1466,N_1355);
xnor U1869 (N_1869,N_1272,N_791);
xnor U1870 (N_1870,N_983,N_1255);
and U1871 (N_1871,N_912,N_1159);
nor U1872 (N_1872,N_838,N_1094);
xor U1873 (N_1873,N_1248,N_1106);
nor U1874 (N_1874,N_756,N_800);
nand U1875 (N_1875,N_862,N_1292);
nor U1876 (N_1876,N_1437,N_945);
nand U1877 (N_1877,N_1128,N_915);
or U1878 (N_1878,N_1208,N_1050);
nand U1879 (N_1879,N_863,N_1218);
xnor U1880 (N_1880,N_879,N_1000);
nand U1881 (N_1881,N_1398,N_983);
and U1882 (N_1882,N_1356,N_1311);
xnor U1883 (N_1883,N_868,N_1119);
and U1884 (N_1884,N_1199,N_874);
and U1885 (N_1885,N_1137,N_1012);
xnor U1886 (N_1886,N_968,N_834);
or U1887 (N_1887,N_840,N_1314);
xor U1888 (N_1888,N_1095,N_1303);
or U1889 (N_1889,N_1015,N_1271);
or U1890 (N_1890,N_1305,N_808);
nand U1891 (N_1891,N_1298,N_1402);
xnor U1892 (N_1892,N_877,N_1162);
xor U1893 (N_1893,N_1482,N_1059);
or U1894 (N_1894,N_1089,N_846);
xnor U1895 (N_1895,N_1072,N_788);
or U1896 (N_1896,N_1084,N_1175);
xor U1897 (N_1897,N_1130,N_1382);
and U1898 (N_1898,N_827,N_795);
xor U1899 (N_1899,N_953,N_1453);
or U1900 (N_1900,N_1285,N_1158);
nor U1901 (N_1901,N_1368,N_830);
xnor U1902 (N_1902,N_937,N_892);
or U1903 (N_1903,N_1011,N_1320);
or U1904 (N_1904,N_1461,N_1344);
or U1905 (N_1905,N_1296,N_1237);
nor U1906 (N_1906,N_1325,N_777);
or U1907 (N_1907,N_1312,N_1264);
nand U1908 (N_1908,N_934,N_1376);
and U1909 (N_1909,N_878,N_1450);
nor U1910 (N_1910,N_1191,N_1070);
and U1911 (N_1911,N_1133,N_865);
xnor U1912 (N_1912,N_1326,N_1402);
nor U1913 (N_1913,N_1333,N_1107);
or U1914 (N_1914,N_779,N_797);
or U1915 (N_1915,N_839,N_1007);
nor U1916 (N_1916,N_1295,N_1180);
and U1917 (N_1917,N_1218,N_956);
nand U1918 (N_1918,N_1039,N_1015);
and U1919 (N_1919,N_1057,N_1149);
xor U1920 (N_1920,N_751,N_1080);
nor U1921 (N_1921,N_1361,N_1077);
and U1922 (N_1922,N_914,N_907);
or U1923 (N_1923,N_1144,N_953);
or U1924 (N_1924,N_872,N_764);
and U1925 (N_1925,N_1038,N_1294);
and U1926 (N_1926,N_771,N_1089);
or U1927 (N_1927,N_901,N_1452);
or U1928 (N_1928,N_1301,N_829);
and U1929 (N_1929,N_1115,N_1096);
and U1930 (N_1930,N_1113,N_840);
or U1931 (N_1931,N_822,N_1166);
nand U1932 (N_1932,N_807,N_1270);
and U1933 (N_1933,N_1058,N_1280);
or U1934 (N_1934,N_1465,N_911);
or U1935 (N_1935,N_796,N_1203);
nor U1936 (N_1936,N_1204,N_841);
nand U1937 (N_1937,N_936,N_1174);
xor U1938 (N_1938,N_1067,N_839);
or U1939 (N_1939,N_1280,N_918);
nor U1940 (N_1940,N_889,N_1151);
or U1941 (N_1941,N_1265,N_1042);
nor U1942 (N_1942,N_1185,N_1308);
nand U1943 (N_1943,N_1458,N_1024);
nand U1944 (N_1944,N_761,N_752);
nor U1945 (N_1945,N_1192,N_1050);
and U1946 (N_1946,N_1305,N_995);
nand U1947 (N_1947,N_962,N_1162);
nor U1948 (N_1948,N_1409,N_1207);
nor U1949 (N_1949,N_1380,N_809);
or U1950 (N_1950,N_1355,N_1184);
and U1951 (N_1951,N_1199,N_1175);
xor U1952 (N_1952,N_1118,N_1220);
nor U1953 (N_1953,N_1294,N_1198);
and U1954 (N_1954,N_995,N_1431);
nand U1955 (N_1955,N_1281,N_1466);
nor U1956 (N_1956,N_1339,N_1327);
xnor U1957 (N_1957,N_990,N_1416);
nand U1958 (N_1958,N_1325,N_1405);
and U1959 (N_1959,N_773,N_806);
nand U1960 (N_1960,N_1474,N_1160);
nor U1961 (N_1961,N_1279,N_822);
nand U1962 (N_1962,N_890,N_837);
and U1963 (N_1963,N_884,N_825);
or U1964 (N_1964,N_994,N_1247);
nand U1965 (N_1965,N_1231,N_968);
or U1966 (N_1966,N_1361,N_810);
nand U1967 (N_1967,N_1243,N_1236);
nor U1968 (N_1968,N_769,N_1169);
and U1969 (N_1969,N_941,N_949);
or U1970 (N_1970,N_1332,N_1167);
nor U1971 (N_1971,N_992,N_1152);
nor U1972 (N_1972,N_1453,N_776);
and U1973 (N_1973,N_1145,N_934);
xnor U1974 (N_1974,N_1242,N_998);
xor U1975 (N_1975,N_1193,N_954);
nand U1976 (N_1976,N_1461,N_1360);
nand U1977 (N_1977,N_1037,N_1209);
or U1978 (N_1978,N_871,N_1085);
nand U1979 (N_1979,N_1294,N_892);
or U1980 (N_1980,N_1010,N_1195);
and U1981 (N_1981,N_1374,N_1113);
nor U1982 (N_1982,N_1224,N_1228);
nor U1983 (N_1983,N_1281,N_1236);
nor U1984 (N_1984,N_1209,N_905);
and U1985 (N_1985,N_1352,N_780);
nand U1986 (N_1986,N_1477,N_1041);
and U1987 (N_1987,N_904,N_1193);
nand U1988 (N_1988,N_1108,N_1314);
xnor U1989 (N_1989,N_818,N_1482);
nand U1990 (N_1990,N_762,N_989);
and U1991 (N_1991,N_1132,N_1176);
nor U1992 (N_1992,N_1371,N_850);
xor U1993 (N_1993,N_842,N_1396);
nor U1994 (N_1994,N_769,N_1366);
xnor U1995 (N_1995,N_1392,N_1431);
nor U1996 (N_1996,N_1276,N_1032);
nor U1997 (N_1997,N_795,N_1345);
xor U1998 (N_1998,N_1287,N_1325);
xor U1999 (N_1999,N_1128,N_1009);
nand U2000 (N_2000,N_785,N_1390);
or U2001 (N_2001,N_782,N_1376);
nand U2002 (N_2002,N_1407,N_1149);
and U2003 (N_2003,N_991,N_954);
xnor U2004 (N_2004,N_1468,N_1011);
and U2005 (N_2005,N_1400,N_1037);
xnor U2006 (N_2006,N_754,N_939);
xor U2007 (N_2007,N_1424,N_1226);
and U2008 (N_2008,N_993,N_1403);
nand U2009 (N_2009,N_1262,N_922);
nand U2010 (N_2010,N_1434,N_1257);
or U2011 (N_2011,N_1196,N_781);
nor U2012 (N_2012,N_1198,N_779);
or U2013 (N_2013,N_1308,N_947);
or U2014 (N_2014,N_1494,N_1126);
or U2015 (N_2015,N_1340,N_1166);
nor U2016 (N_2016,N_885,N_1453);
nand U2017 (N_2017,N_1389,N_896);
and U2018 (N_2018,N_1409,N_931);
or U2019 (N_2019,N_1144,N_992);
and U2020 (N_2020,N_1418,N_1158);
and U2021 (N_2021,N_794,N_1312);
xnor U2022 (N_2022,N_1004,N_1357);
xnor U2023 (N_2023,N_1297,N_1336);
nand U2024 (N_2024,N_840,N_1429);
or U2025 (N_2025,N_1358,N_1383);
and U2026 (N_2026,N_1082,N_844);
or U2027 (N_2027,N_1494,N_845);
nand U2028 (N_2028,N_990,N_1159);
and U2029 (N_2029,N_1118,N_878);
or U2030 (N_2030,N_1042,N_1481);
nand U2031 (N_2031,N_838,N_877);
and U2032 (N_2032,N_1349,N_1103);
nor U2033 (N_2033,N_844,N_1374);
nor U2034 (N_2034,N_1342,N_774);
xor U2035 (N_2035,N_1238,N_1194);
nor U2036 (N_2036,N_1132,N_1139);
nand U2037 (N_2037,N_1316,N_777);
and U2038 (N_2038,N_857,N_999);
nor U2039 (N_2039,N_907,N_1204);
xor U2040 (N_2040,N_952,N_1429);
nor U2041 (N_2041,N_797,N_1482);
and U2042 (N_2042,N_851,N_960);
and U2043 (N_2043,N_1033,N_1253);
xor U2044 (N_2044,N_1385,N_1145);
nor U2045 (N_2045,N_1390,N_840);
nand U2046 (N_2046,N_1372,N_1142);
nor U2047 (N_2047,N_1399,N_963);
or U2048 (N_2048,N_1489,N_1278);
nor U2049 (N_2049,N_1303,N_1211);
nor U2050 (N_2050,N_1268,N_1459);
and U2051 (N_2051,N_1296,N_1322);
xnor U2052 (N_2052,N_835,N_1309);
nand U2053 (N_2053,N_1088,N_1355);
or U2054 (N_2054,N_1178,N_997);
xor U2055 (N_2055,N_1417,N_887);
nand U2056 (N_2056,N_752,N_1072);
xnor U2057 (N_2057,N_919,N_818);
nand U2058 (N_2058,N_1322,N_1439);
nor U2059 (N_2059,N_884,N_1441);
nand U2060 (N_2060,N_1036,N_1222);
or U2061 (N_2061,N_1017,N_1391);
and U2062 (N_2062,N_1178,N_839);
nor U2063 (N_2063,N_1157,N_1290);
xor U2064 (N_2064,N_923,N_1057);
or U2065 (N_2065,N_1046,N_1191);
or U2066 (N_2066,N_1340,N_906);
nor U2067 (N_2067,N_1172,N_1260);
nand U2068 (N_2068,N_1454,N_1146);
nand U2069 (N_2069,N_1377,N_1252);
xor U2070 (N_2070,N_1118,N_1098);
xnor U2071 (N_2071,N_1415,N_1059);
xor U2072 (N_2072,N_789,N_818);
nor U2073 (N_2073,N_889,N_1027);
or U2074 (N_2074,N_1085,N_1046);
nor U2075 (N_2075,N_1104,N_1374);
or U2076 (N_2076,N_1152,N_1194);
or U2077 (N_2077,N_1027,N_864);
nor U2078 (N_2078,N_1141,N_763);
xnor U2079 (N_2079,N_1363,N_1233);
nor U2080 (N_2080,N_1136,N_841);
xor U2081 (N_2081,N_1321,N_1422);
nand U2082 (N_2082,N_786,N_1352);
or U2083 (N_2083,N_855,N_1357);
nor U2084 (N_2084,N_1191,N_1239);
xnor U2085 (N_2085,N_1305,N_1318);
and U2086 (N_2086,N_995,N_1344);
nor U2087 (N_2087,N_1105,N_1051);
nor U2088 (N_2088,N_1152,N_982);
nor U2089 (N_2089,N_999,N_1075);
nor U2090 (N_2090,N_970,N_793);
xor U2091 (N_2091,N_773,N_1133);
xor U2092 (N_2092,N_1421,N_963);
and U2093 (N_2093,N_1086,N_909);
or U2094 (N_2094,N_1019,N_1051);
and U2095 (N_2095,N_1250,N_881);
or U2096 (N_2096,N_1052,N_1029);
and U2097 (N_2097,N_847,N_1381);
nand U2098 (N_2098,N_1468,N_1273);
and U2099 (N_2099,N_1400,N_924);
nand U2100 (N_2100,N_1063,N_890);
and U2101 (N_2101,N_845,N_828);
nor U2102 (N_2102,N_982,N_895);
and U2103 (N_2103,N_1395,N_989);
and U2104 (N_2104,N_1235,N_1175);
or U2105 (N_2105,N_935,N_764);
nor U2106 (N_2106,N_966,N_847);
or U2107 (N_2107,N_1425,N_991);
or U2108 (N_2108,N_1454,N_1265);
nor U2109 (N_2109,N_770,N_1333);
or U2110 (N_2110,N_1354,N_1499);
nand U2111 (N_2111,N_1056,N_1112);
and U2112 (N_2112,N_838,N_794);
xnor U2113 (N_2113,N_1006,N_1465);
or U2114 (N_2114,N_1167,N_928);
and U2115 (N_2115,N_1179,N_785);
and U2116 (N_2116,N_1488,N_965);
and U2117 (N_2117,N_1137,N_868);
nand U2118 (N_2118,N_780,N_1395);
nor U2119 (N_2119,N_939,N_1193);
and U2120 (N_2120,N_1259,N_768);
nand U2121 (N_2121,N_814,N_914);
xnor U2122 (N_2122,N_1100,N_1022);
nor U2123 (N_2123,N_1041,N_1209);
and U2124 (N_2124,N_898,N_1090);
nor U2125 (N_2125,N_1140,N_1447);
or U2126 (N_2126,N_1426,N_1438);
xor U2127 (N_2127,N_1406,N_918);
and U2128 (N_2128,N_1290,N_1421);
xnor U2129 (N_2129,N_861,N_817);
nand U2130 (N_2130,N_954,N_859);
and U2131 (N_2131,N_844,N_1014);
xor U2132 (N_2132,N_1233,N_1442);
or U2133 (N_2133,N_1204,N_1269);
and U2134 (N_2134,N_1049,N_1476);
xor U2135 (N_2135,N_762,N_936);
nor U2136 (N_2136,N_1471,N_832);
xor U2137 (N_2137,N_1087,N_1451);
nor U2138 (N_2138,N_1045,N_997);
nand U2139 (N_2139,N_1028,N_1252);
or U2140 (N_2140,N_1433,N_1081);
and U2141 (N_2141,N_791,N_1428);
and U2142 (N_2142,N_888,N_1488);
xnor U2143 (N_2143,N_1004,N_1165);
nand U2144 (N_2144,N_1377,N_1260);
and U2145 (N_2145,N_1428,N_1052);
nor U2146 (N_2146,N_825,N_1076);
nand U2147 (N_2147,N_1481,N_1375);
nand U2148 (N_2148,N_1330,N_1334);
and U2149 (N_2149,N_1110,N_1202);
nand U2150 (N_2150,N_786,N_1431);
nand U2151 (N_2151,N_811,N_990);
xnor U2152 (N_2152,N_788,N_1236);
xor U2153 (N_2153,N_1455,N_1260);
nor U2154 (N_2154,N_1370,N_1038);
nand U2155 (N_2155,N_1281,N_770);
nand U2156 (N_2156,N_1448,N_1113);
nor U2157 (N_2157,N_752,N_952);
and U2158 (N_2158,N_1295,N_1151);
or U2159 (N_2159,N_1378,N_1252);
nor U2160 (N_2160,N_1362,N_871);
xor U2161 (N_2161,N_875,N_1214);
and U2162 (N_2162,N_1321,N_1186);
nor U2163 (N_2163,N_1227,N_1029);
xnor U2164 (N_2164,N_1211,N_854);
xor U2165 (N_2165,N_828,N_788);
or U2166 (N_2166,N_1397,N_887);
nand U2167 (N_2167,N_1447,N_1353);
or U2168 (N_2168,N_1029,N_1335);
or U2169 (N_2169,N_1063,N_1071);
nor U2170 (N_2170,N_1186,N_1385);
nor U2171 (N_2171,N_1335,N_1097);
xnor U2172 (N_2172,N_1180,N_1254);
and U2173 (N_2173,N_825,N_1237);
or U2174 (N_2174,N_954,N_1091);
and U2175 (N_2175,N_1209,N_1279);
xor U2176 (N_2176,N_814,N_1371);
or U2177 (N_2177,N_1040,N_1282);
xor U2178 (N_2178,N_1390,N_1289);
and U2179 (N_2179,N_1041,N_1487);
nand U2180 (N_2180,N_1169,N_806);
or U2181 (N_2181,N_830,N_775);
xnor U2182 (N_2182,N_1195,N_1213);
or U2183 (N_2183,N_809,N_1402);
nand U2184 (N_2184,N_1128,N_1117);
nand U2185 (N_2185,N_1245,N_1090);
nand U2186 (N_2186,N_786,N_1397);
xor U2187 (N_2187,N_977,N_1469);
or U2188 (N_2188,N_1044,N_1236);
nand U2189 (N_2189,N_1313,N_946);
nor U2190 (N_2190,N_1488,N_1436);
or U2191 (N_2191,N_1315,N_1116);
and U2192 (N_2192,N_1184,N_986);
or U2193 (N_2193,N_783,N_986);
or U2194 (N_2194,N_1374,N_1029);
or U2195 (N_2195,N_1364,N_857);
or U2196 (N_2196,N_1230,N_858);
or U2197 (N_2197,N_1264,N_944);
xnor U2198 (N_2198,N_1319,N_895);
nor U2199 (N_2199,N_973,N_985);
xnor U2200 (N_2200,N_1380,N_802);
or U2201 (N_2201,N_903,N_1084);
nand U2202 (N_2202,N_759,N_1193);
xor U2203 (N_2203,N_1066,N_1337);
nor U2204 (N_2204,N_971,N_1127);
xor U2205 (N_2205,N_896,N_964);
and U2206 (N_2206,N_1023,N_841);
nor U2207 (N_2207,N_1361,N_1498);
nand U2208 (N_2208,N_1140,N_1153);
or U2209 (N_2209,N_1086,N_867);
and U2210 (N_2210,N_1315,N_992);
or U2211 (N_2211,N_849,N_1151);
or U2212 (N_2212,N_814,N_848);
or U2213 (N_2213,N_1231,N_844);
nand U2214 (N_2214,N_827,N_1335);
nor U2215 (N_2215,N_1082,N_903);
or U2216 (N_2216,N_1205,N_1213);
or U2217 (N_2217,N_1191,N_1248);
xnor U2218 (N_2218,N_911,N_1177);
and U2219 (N_2219,N_849,N_919);
or U2220 (N_2220,N_1036,N_1157);
nor U2221 (N_2221,N_985,N_1295);
and U2222 (N_2222,N_842,N_1149);
nand U2223 (N_2223,N_1389,N_770);
and U2224 (N_2224,N_1013,N_1430);
nor U2225 (N_2225,N_1231,N_1093);
nand U2226 (N_2226,N_769,N_901);
nand U2227 (N_2227,N_880,N_1181);
nand U2228 (N_2228,N_1410,N_1213);
xor U2229 (N_2229,N_1345,N_822);
or U2230 (N_2230,N_1343,N_1134);
nand U2231 (N_2231,N_1174,N_1196);
xor U2232 (N_2232,N_1034,N_1053);
or U2233 (N_2233,N_1216,N_1312);
or U2234 (N_2234,N_1143,N_818);
or U2235 (N_2235,N_1251,N_1459);
nand U2236 (N_2236,N_813,N_1078);
xor U2237 (N_2237,N_913,N_860);
nand U2238 (N_2238,N_1225,N_1435);
xnor U2239 (N_2239,N_1249,N_895);
and U2240 (N_2240,N_1435,N_1175);
nor U2241 (N_2241,N_1188,N_1001);
nor U2242 (N_2242,N_1177,N_1001);
nand U2243 (N_2243,N_1265,N_1471);
nor U2244 (N_2244,N_1196,N_1142);
or U2245 (N_2245,N_1051,N_761);
xor U2246 (N_2246,N_1186,N_998);
nor U2247 (N_2247,N_1153,N_1152);
nand U2248 (N_2248,N_887,N_1204);
nand U2249 (N_2249,N_1162,N_1448);
xor U2250 (N_2250,N_1525,N_2060);
or U2251 (N_2251,N_1937,N_1941);
xnor U2252 (N_2252,N_2135,N_2223);
and U2253 (N_2253,N_1575,N_1520);
xnor U2254 (N_2254,N_1701,N_1666);
nor U2255 (N_2255,N_1800,N_2109);
and U2256 (N_2256,N_1566,N_2215);
or U2257 (N_2257,N_2190,N_1567);
and U2258 (N_2258,N_2068,N_1695);
nor U2259 (N_2259,N_2228,N_1549);
nor U2260 (N_2260,N_2176,N_2084);
nand U2261 (N_2261,N_1785,N_1512);
nand U2262 (N_2262,N_2005,N_2094);
or U2263 (N_2263,N_1874,N_1726);
nand U2264 (N_2264,N_1768,N_2170);
or U2265 (N_2265,N_2233,N_2107);
nor U2266 (N_2266,N_2052,N_1594);
and U2267 (N_2267,N_1508,N_1625);
nand U2268 (N_2268,N_1672,N_1585);
and U2269 (N_2269,N_1988,N_2130);
nor U2270 (N_2270,N_2151,N_2159);
or U2271 (N_2271,N_2117,N_1892);
xnor U2272 (N_2272,N_1534,N_1923);
nor U2273 (N_2273,N_1965,N_1600);
nor U2274 (N_2274,N_1572,N_1731);
nor U2275 (N_2275,N_2168,N_1860);
and U2276 (N_2276,N_1806,N_1680);
nor U2277 (N_2277,N_1902,N_2201);
xnor U2278 (N_2278,N_1802,N_1952);
xor U2279 (N_2279,N_2202,N_1515);
xnor U2280 (N_2280,N_1932,N_1839);
nand U2281 (N_2281,N_1691,N_1827);
xnor U2282 (N_2282,N_1503,N_1544);
xor U2283 (N_2283,N_2024,N_2037);
and U2284 (N_2284,N_2186,N_1908);
and U2285 (N_2285,N_1517,N_1976);
or U2286 (N_2286,N_2008,N_1611);
nor U2287 (N_2287,N_1985,N_1776);
nand U2288 (N_2288,N_2081,N_1911);
and U2289 (N_2289,N_1886,N_1794);
nand U2290 (N_2290,N_2053,N_1862);
xnor U2291 (N_2291,N_1852,N_1748);
or U2292 (N_2292,N_2021,N_2067);
nand U2293 (N_2293,N_1917,N_2050);
nor U2294 (N_2294,N_2063,N_1876);
and U2295 (N_2295,N_2129,N_2019);
xor U2296 (N_2296,N_2163,N_2073);
or U2297 (N_2297,N_1675,N_1755);
nand U2298 (N_2298,N_1685,N_1778);
nand U2299 (N_2299,N_2234,N_2072);
or U2300 (N_2300,N_1626,N_1759);
and U2301 (N_2301,N_2022,N_1764);
xnor U2302 (N_2302,N_1717,N_2164);
or U2303 (N_2303,N_2136,N_1724);
or U2304 (N_2304,N_1929,N_1579);
xnor U2305 (N_2305,N_1834,N_1977);
and U2306 (N_2306,N_2016,N_1989);
nand U2307 (N_2307,N_1889,N_1822);
nand U2308 (N_2308,N_1599,N_1820);
nand U2309 (N_2309,N_2230,N_1518);
nor U2310 (N_2310,N_1735,N_2145);
xnor U2311 (N_2311,N_2114,N_1519);
xor U2312 (N_2312,N_1868,N_1938);
or U2313 (N_2313,N_2049,N_1670);
or U2314 (N_2314,N_2115,N_1782);
nor U2315 (N_2315,N_2237,N_1552);
or U2316 (N_2316,N_2142,N_1700);
or U2317 (N_2317,N_1895,N_1578);
nor U2318 (N_2318,N_2134,N_2180);
nand U2319 (N_2319,N_1950,N_2225);
xnor U2320 (N_2320,N_1773,N_1760);
or U2321 (N_2321,N_1931,N_2137);
or U2322 (N_2322,N_1942,N_1875);
or U2323 (N_2323,N_2214,N_1658);
or U2324 (N_2324,N_2108,N_2172);
nor U2325 (N_2325,N_1657,N_2092);
xor U2326 (N_2326,N_2111,N_2040);
or U2327 (N_2327,N_1610,N_2138);
xnor U2328 (N_2328,N_1709,N_2013);
or U2329 (N_2329,N_1619,N_2075);
xnor U2330 (N_2330,N_1509,N_2083);
or U2331 (N_2331,N_1707,N_1817);
or U2332 (N_2332,N_1765,N_1646);
or U2333 (N_2333,N_1713,N_2080);
nor U2334 (N_2334,N_2209,N_1970);
xnor U2335 (N_2335,N_1530,N_1571);
nor U2336 (N_2336,N_1754,N_2061);
xor U2337 (N_2337,N_1510,N_1702);
and U2338 (N_2338,N_2218,N_2112);
and U2339 (N_2339,N_1922,N_1647);
xnor U2340 (N_2340,N_1589,N_1692);
nand U2341 (N_2341,N_2187,N_1537);
xor U2342 (N_2342,N_1655,N_1858);
nand U2343 (N_2343,N_2141,N_1767);
and U2344 (N_2344,N_1752,N_1810);
nor U2345 (N_2345,N_2236,N_1939);
nand U2346 (N_2346,N_1984,N_2222);
or U2347 (N_2347,N_2193,N_1940);
xnor U2348 (N_2348,N_1850,N_1795);
or U2349 (N_2349,N_1677,N_1828);
nor U2350 (N_2350,N_1777,N_1660);
nand U2351 (N_2351,N_1650,N_2227);
nand U2352 (N_2352,N_2113,N_1905);
nand U2353 (N_2353,N_1962,N_1901);
and U2354 (N_2354,N_1704,N_1592);
xor U2355 (N_2355,N_2191,N_1547);
or U2356 (N_2356,N_1705,N_2173);
or U2357 (N_2357,N_1994,N_2248);
or U2358 (N_2358,N_1999,N_1612);
xor U2359 (N_2359,N_2093,N_2125);
or U2360 (N_2360,N_1961,N_1654);
xnor U2361 (N_2361,N_1809,N_1667);
nand U2362 (N_2362,N_1866,N_2192);
xor U2363 (N_2363,N_1881,N_2025);
xor U2364 (N_2364,N_1921,N_1943);
nand U2365 (N_2365,N_1643,N_1811);
nand U2366 (N_2366,N_2028,N_1842);
nand U2367 (N_2367,N_1745,N_1516);
nand U2368 (N_2368,N_1545,N_1887);
xor U2369 (N_2369,N_1521,N_1669);
or U2370 (N_2370,N_2089,N_1927);
and U2371 (N_2371,N_2038,N_1720);
nor U2372 (N_2372,N_1608,N_1631);
xnor U2373 (N_2373,N_1555,N_2247);
or U2374 (N_2374,N_1684,N_1853);
or U2375 (N_2375,N_1529,N_1606);
nand U2376 (N_2376,N_1715,N_2232);
nand U2377 (N_2377,N_1629,N_1980);
nand U2378 (N_2378,N_1668,N_2181);
nor U2379 (N_2379,N_2014,N_1603);
and U2380 (N_2380,N_2047,N_1770);
nor U2381 (N_2381,N_2212,N_2090);
nor U2382 (N_2382,N_1974,N_1873);
or U2383 (N_2383,N_1601,N_2179);
xor U2384 (N_2384,N_2221,N_2224);
nand U2385 (N_2385,N_1664,N_2206);
nand U2386 (N_2386,N_1807,N_1779);
and U2387 (N_2387,N_1659,N_2103);
xnor U2388 (N_2388,N_2045,N_1727);
or U2389 (N_2389,N_1632,N_2189);
and U2390 (N_2390,N_1826,N_1930);
or U2391 (N_2391,N_2204,N_1662);
xor U2392 (N_2392,N_1762,N_2043);
nor U2393 (N_2393,N_2213,N_1651);
nand U2394 (N_2394,N_1910,N_1628);
nor U2395 (N_2395,N_1992,N_1689);
and U2396 (N_2396,N_1502,N_1602);
nand U2397 (N_2397,N_2100,N_1898);
nor U2398 (N_2398,N_2160,N_2182);
nor U2399 (N_2399,N_1661,N_2018);
xnor U2400 (N_2400,N_1627,N_1694);
xor U2401 (N_2401,N_1832,N_2033);
or U2402 (N_2402,N_1590,N_1972);
nand U2403 (N_2403,N_1569,N_1871);
xor U2404 (N_2404,N_2238,N_1904);
or U2405 (N_2405,N_1686,N_2184);
or U2406 (N_2406,N_1856,N_2069);
and U2407 (N_2407,N_1751,N_1725);
or U2408 (N_2408,N_2231,N_2010);
and U2409 (N_2409,N_1722,N_2183);
xnor U2410 (N_2410,N_2102,N_1531);
nand U2411 (N_2411,N_2088,N_1591);
nand U2412 (N_2412,N_2133,N_1738);
or U2413 (N_2413,N_1987,N_1918);
or U2414 (N_2414,N_1674,N_1635);
or U2415 (N_2415,N_2096,N_1814);
nand U2416 (N_2416,N_1574,N_2099);
xnor U2417 (N_2417,N_1582,N_2098);
nor U2418 (N_2418,N_1926,N_1774);
and U2419 (N_2419,N_2119,N_1682);
nor U2420 (N_2420,N_1966,N_1840);
xor U2421 (N_2421,N_2106,N_2044);
or U2422 (N_2422,N_1763,N_2178);
or U2423 (N_2423,N_1830,N_1893);
nand U2424 (N_2424,N_2062,N_1818);
nand U2425 (N_2425,N_1696,N_2007);
xnor U2426 (N_2426,N_1812,N_2120);
xor U2427 (N_2427,N_2001,N_2166);
nor U2428 (N_2428,N_2101,N_1747);
and U2429 (N_2429,N_1882,N_1679);
nor U2430 (N_2430,N_1789,N_2023);
and U2431 (N_2431,N_2076,N_1706);
nand U2432 (N_2432,N_1993,N_1780);
nand U2433 (N_2433,N_2150,N_2065);
nand U2434 (N_2434,N_1618,N_1857);
nor U2435 (N_2435,N_1546,N_1824);
nor U2436 (N_2436,N_1639,N_1522);
and U2437 (N_2437,N_2144,N_1878);
xnor U2438 (N_2438,N_2059,N_1741);
xnor U2439 (N_2439,N_2104,N_2165);
or U2440 (N_2440,N_1753,N_1843);
or U2441 (N_2441,N_1796,N_2105);
nand U2442 (N_2442,N_1855,N_1836);
nand U2443 (N_2443,N_1803,N_2064);
nor U2444 (N_2444,N_1597,N_1790);
nor U2445 (N_2445,N_1543,N_1900);
or U2446 (N_2446,N_2097,N_1924);
or U2447 (N_2447,N_1982,N_2203);
and U2448 (N_2448,N_1699,N_1728);
or U2449 (N_2449,N_2154,N_1757);
and U2450 (N_2450,N_2155,N_1528);
xor U2451 (N_2451,N_1955,N_1527);
xor U2452 (N_2452,N_2077,N_2070);
nor U2453 (N_2453,N_1959,N_1548);
nand U2454 (N_2454,N_1514,N_2085);
xnor U2455 (N_2455,N_2127,N_1894);
nand U2456 (N_2456,N_2199,N_1678);
and U2457 (N_2457,N_1645,N_2175);
nor U2458 (N_2458,N_1864,N_1698);
nand U2459 (N_2459,N_2051,N_2058);
and U2460 (N_2460,N_1671,N_1663);
xor U2461 (N_2461,N_1787,N_1554);
and U2462 (N_2462,N_1504,N_2132);
and U2463 (N_2463,N_1885,N_2095);
nor U2464 (N_2464,N_1511,N_2210);
nor U2465 (N_2465,N_1732,N_1799);
nand U2466 (N_2466,N_2011,N_1622);
nor U2467 (N_2467,N_1958,N_1983);
xor U2468 (N_2468,N_1580,N_1936);
and U2469 (N_2469,N_1890,N_2032);
xor U2470 (N_2470,N_1960,N_1690);
or U2471 (N_2471,N_1729,N_2009);
nor U2472 (N_2472,N_1532,N_2169);
or U2473 (N_2473,N_2217,N_1808);
xor U2474 (N_2474,N_1888,N_1621);
xor U2475 (N_2475,N_2071,N_1605);
nor U2476 (N_2476,N_2004,N_2177);
xnor U2477 (N_2477,N_2148,N_1733);
nand U2478 (N_2478,N_1956,N_1542);
or U2479 (N_2479,N_2091,N_1640);
and U2480 (N_2480,N_1833,N_2118);
and U2481 (N_2481,N_1793,N_1906);
nor U2482 (N_2482,N_2039,N_1872);
and U2483 (N_2483,N_1615,N_2029);
nand U2484 (N_2484,N_1501,N_2207);
and U2485 (N_2485,N_2239,N_1772);
or U2486 (N_2486,N_1859,N_1869);
xnor U2487 (N_2487,N_1756,N_1581);
xnor U2488 (N_2488,N_1607,N_1624);
nand U2489 (N_2489,N_1513,N_1734);
nand U2490 (N_2490,N_1865,N_1642);
xnor U2491 (N_2491,N_1633,N_1617);
xor U2492 (N_2492,N_1573,N_2015);
nand U2493 (N_2493,N_1596,N_1712);
nor U2494 (N_2494,N_2194,N_1584);
and U2495 (N_2495,N_1740,N_1953);
nor U2496 (N_2496,N_2140,N_1653);
nor U2497 (N_2497,N_2031,N_1714);
nor U2498 (N_2498,N_1746,N_1844);
or U2499 (N_2499,N_1766,N_1649);
and U2500 (N_2500,N_1879,N_2124);
xnor U2501 (N_2501,N_1903,N_1831);
nor U2502 (N_2502,N_1791,N_1681);
nand U2503 (N_2503,N_2152,N_2122);
nor U2504 (N_2504,N_1816,N_1576);
or U2505 (N_2505,N_1570,N_1560);
xnor U2506 (N_2506,N_1897,N_1801);
xor U2507 (N_2507,N_1586,N_1673);
and U2508 (N_2508,N_1971,N_1825);
xnor U2509 (N_2509,N_2055,N_1915);
nor U2510 (N_2510,N_1996,N_1963);
nor U2511 (N_2511,N_2042,N_2017);
xor U2512 (N_2512,N_1783,N_1703);
xnor U2513 (N_2513,N_2245,N_1784);
xnor U2514 (N_2514,N_1750,N_1688);
nor U2515 (N_2515,N_2185,N_1620);
nor U2516 (N_2516,N_1946,N_2035);
or U2517 (N_2517,N_1523,N_1861);
nor U2518 (N_2518,N_2048,N_2147);
xor U2519 (N_2519,N_2219,N_2027);
nor U2520 (N_2520,N_1634,N_1805);
nand U2521 (N_2521,N_1835,N_1870);
nor U2522 (N_2522,N_1693,N_2216);
or U2523 (N_2523,N_1708,N_2078);
and U2524 (N_2524,N_1550,N_1697);
xnor U2525 (N_2525,N_1914,N_2034);
and U2526 (N_2526,N_2161,N_1539);
xor U2527 (N_2527,N_1710,N_1979);
or U2528 (N_2528,N_2205,N_1909);
and U2529 (N_2529,N_1829,N_2188);
nor U2530 (N_2530,N_1742,N_1716);
and U2531 (N_2531,N_1577,N_1614);
nand U2532 (N_2532,N_1925,N_1736);
nor U2533 (N_2533,N_2157,N_1786);
and U2534 (N_2534,N_1761,N_2030);
xnor U2535 (N_2535,N_2229,N_2123);
nor U2536 (N_2536,N_1583,N_1846);
and U2537 (N_2537,N_2087,N_2149);
nor U2538 (N_2538,N_1907,N_1973);
or U2539 (N_2539,N_1838,N_1967);
xnor U2540 (N_2540,N_2041,N_1975);
or U2541 (N_2541,N_1919,N_2167);
or U2542 (N_2542,N_1863,N_1991);
xnor U2543 (N_2543,N_1851,N_1758);
xnor U2544 (N_2544,N_1781,N_1562);
nand U2545 (N_2545,N_1719,N_1553);
nand U2546 (N_2546,N_1848,N_2158);
nor U2547 (N_2547,N_2208,N_2195);
nand U2548 (N_2548,N_2153,N_1536);
or U2549 (N_2549,N_2003,N_1813);
and U2550 (N_2550,N_1638,N_1636);
nor U2551 (N_2551,N_1609,N_1947);
xnor U2552 (N_2552,N_1588,N_1899);
xor U2553 (N_2553,N_2243,N_1997);
or U2554 (N_2554,N_1986,N_2156);
nand U2555 (N_2555,N_1564,N_2082);
or U2556 (N_2556,N_1556,N_1644);
nand U2557 (N_2557,N_1557,N_1718);
xnor U2558 (N_2558,N_1526,N_2139);
nand U2559 (N_2559,N_2131,N_2046);
xor U2560 (N_2560,N_1815,N_1823);
nor U2561 (N_2561,N_2057,N_2249);
xnor U2562 (N_2562,N_1683,N_1500);
nor U2563 (N_2563,N_1721,N_1934);
and U2564 (N_2564,N_1598,N_1623);
nand U2565 (N_2565,N_1559,N_1837);
xnor U2566 (N_2566,N_1849,N_1944);
or U2567 (N_2567,N_1804,N_1558);
and U2568 (N_2568,N_2074,N_1995);
or U2569 (N_2569,N_2240,N_2211);
xor U2570 (N_2570,N_2116,N_1769);
nand U2571 (N_2571,N_1896,N_1506);
nor U2572 (N_2572,N_1916,N_1613);
or U2573 (N_2573,N_2036,N_1792);
nor U2574 (N_2574,N_2244,N_1891);
or U2575 (N_2575,N_2241,N_1883);
and U2576 (N_2576,N_1788,N_2056);
and U2577 (N_2577,N_2220,N_2066);
xor U2578 (N_2578,N_2126,N_2174);
and U2579 (N_2579,N_1630,N_1637);
xor U2580 (N_2580,N_1541,N_2235);
nor U2581 (N_2581,N_1648,N_1730);
and U2582 (N_2582,N_1819,N_2128);
xor U2583 (N_2583,N_1998,N_1945);
and U2584 (N_2584,N_2054,N_1676);
nand U2585 (N_2585,N_1884,N_2086);
nand U2586 (N_2586,N_1797,N_2121);
and U2587 (N_2587,N_2006,N_2026);
and U2588 (N_2588,N_2000,N_1968);
xnor U2589 (N_2589,N_1954,N_1563);
nand U2590 (N_2590,N_1951,N_1641);
nor U2591 (N_2591,N_1665,N_1593);
nor U2592 (N_2592,N_1565,N_1775);
and U2593 (N_2593,N_2171,N_1744);
or U2594 (N_2594,N_1561,N_1847);
nand U2595 (N_2595,N_2110,N_1771);
xnor U2596 (N_2596,N_1841,N_1505);
nand U2597 (N_2597,N_2246,N_1845);
or U2598 (N_2598,N_1978,N_2079);
xor U2599 (N_2599,N_1535,N_2143);
xnor U2600 (N_2600,N_1749,N_2020);
xnor U2601 (N_2601,N_1935,N_1933);
or U2602 (N_2602,N_1969,N_1568);
nor U2603 (N_2603,N_2196,N_2198);
and U2604 (N_2604,N_1538,N_1507);
nand U2605 (N_2605,N_1913,N_1948);
or U2606 (N_2606,N_1524,N_1798);
and U2607 (N_2607,N_1739,N_1957);
xor U2608 (N_2608,N_1656,N_1920);
or U2609 (N_2609,N_1723,N_2226);
or U2610 (N_2610,N_1551,N_1595);
xnor U2611 (N_2611,N_1981,N_1711);
nand U2612 (N_2612,N_1880,N_2146);
xor U2613 (N_2613,N_1867,N_1928);
or U2614 (N_2614,N_2162,N_1743);
or U2615 (N_2615,N_2197,N_2002);
and U2616 (N_2616,N_2012,N_1854);
nor U2617 (N_2617,N_1533,N_1964);
xnor U2618 (N_2618,N_1821,N_1616);
nand U2619 (N_2619,N_1912,N_1540);
nor U2620 (N_2620,N_1877,N_2242);
xnor U2621 (N_2621,N_1687,N_1949);
or U2622 (N_2622,N_1990,N_1737);
or U2623 (N_2623,N_1652,N_1587);
or U2624 (N_2624,N_1604,N_2200);
xor U2625 (N_2625,N_1505,N_1946);
xnor U2626 (N_2626,N_1767,N_1687);
or U2627 (N_2627,N_1730,N_1640);
or U2628 (N_2628,N_1605,N_1597);
xnor U2629 (N_2629,N_1661,N_1519);
or U2630 (N_2630,N_2088,N_1716);
nor U2631 (N_2631,N_1786,N_2179);
and U2632 (N_2632,N_1912,N_1678);
nand U2633 (N_2633,N_2148,N_2011);
or U2634 (N_2634,N_1887,N_2112);
and U2635 (N_2635,N_1751,N_1697);
nand U2636 (N_2636,N_2112,N_2060);
xnor U2637 (N_2637,N_1994,N_1771);
nand U2638 (N_2638,N_1811,N_1637);
or U2639 (N_2639,N_1630,N_1901);
and U2640 (N_2640,N_2168,N_1896);
xor U2641 (N_2641,N_1562,N_1881);
xor U2642 (N_2642,N_1985,N_2223);
nand U2643 (N_2643,N_1685,N_1682);
xnor U2644 (N_2644,N_2220,N_1925);
xor U2645 (N_2645,N_1846,N_2236);
xnor U2646 (N_2646,N_1532,N_2036);
nand U2647 (N_2647,N_1553,N_1967);
and U2648 (N_2648,N_1869,N_1768);
xor U2649 (N_2649,N_2122,N_1831);
xnor U2650 (N_2650,N_2206,N_1626);
and U2651 (N_2651,N_1912,N_2170);
nand U2652 (N_2652,N_1839,N_1749);
and U2653 (N_2653,N_1728,N_1686);
or U2654 (N_2654,N_1726,N_1760);
nand U2655 (N_2655,N_2005,N_1922);
nor U2656 (N_2656,N_1643,N_1869);
or U2657 (N_2657,N_1718,N_2046);
and U2658 (N_2658,N_1867,N_1904);
xnor U2659 (N_2659,N_1937,N_1544);
and U2660 (N_2660,N_1829,N_1852);
or U2661 (N_2661,N_1603,N_2041);
and U2662 (N_2662,N_2206,N_2101);
xnor U2663 (N_2663,N_1758,N_1879);
nand U2664 (N_2664,N_1608,N_2245);
nor U2665 (N_2665,N_1977,N_1686);
nand U2666 (N_2666,N_1524,N_1572);
xnor U2667 (N_2667,N_1586,N_1786);
nand U2668 (N_2668,N_1562,N_1891);
nand U2669 (N_2669,N_1559,N_1658);
or U2670 (N_2670,N_1784,N_2249);
nand U2671 (N_2671,N_1759,N_2154);
xor U2672 (N_2672,N_1625,N_1635);
nor U2673 (N_2673,N_1763,N_2004);
nor U2674 (N_2674,N_2058,N_2159);
xor U2675 (N_2675,N_1573,N_2217);
or U2676 (N_2676,N_1621,N_2237);
nand U2677 (N_2677,N_1735,N_1619);
nand U2678 (N_2678,N_1666,N_1990);
xnor U2679 (N_2679,N_1782,N_1814);
xnor U2680 (N_2680,N_1824,N_1636);
nand U2681 (N_2681,N_1694,N_1813);
nor U2682 (N_2682,N_1555,N_2146);
and U2683 (N_2683,N_1567,N_1792);
nor U2684 (N_2684,N_2229,N_1708);
or U2685 (N_2685,N_1825,N_1722);
nor U2686 (N_2686,N_1532,N_1852);
xnor U2687 (N_2687,N_2000,N_1606);
or U2688 (N_2688,N_2102,N_1967);
nand U2689 (N_2689,N_1688,N_2195);
and U2690 (N_2690,N_1745,N_2078);
and U2691 (N_2691,N_1565,N_2064);
or U2692 (N_2692,N_2234,N_1772);
or U2693 (N_2693,N_1861,N_2122);
xnor U2694 (N_2694,N_1773,N_1551);
nand U2695 (N_2695,N_1598,N_1865);
and U2696 (N_2696,N_2082,N_1966);
and U2697 (N_2697,N_2220,N_1929);
nor U2698 (N_2698,N_2000,N_2074);
or U2699 (N_2699,N_1718,N_1763);
or U2700 (N_2700,N_1597,N_2147);
and U2701 (N_2701,N_1951,N_1958);
xor U2702 (N_2702,N_1891,N_2179);
xor U2703 (N_2703,N_1885,N_1681);
and U2704 (N_2704,N_1869,N_1876);
nor U2705 (N_2705,N_1573,N_1518);
xor U2706 (N_2706,N_1944,N_2110);
nand U2707 (N_2707,N_1759,N_1683);
nor U2708 (N_2708,N_1648,N_1985);
and U2709 (N_2709,N_1959,N_2200);
nor U2710 (N_2710,N_1585,N_2050);
nor U2711 (N_2711,N_1823,N_1973);
xor U2712 (N_2712,N_1833,N_2094);
xor U2713 (N_2713,N_1782,N_1917);
or U2714 (N_2714,N_2133,N_1550);
and U2715 (N_2715,N_2107,N_2139);
and U2716 (N_2716,N_1904,N_2013);
and U2717 (N_2717,N_2205,N_1996);
or U2718 (N_2718,N_1825,N_2240);
and U2719 (N_2719,N_1722,N_1754);
nand U2720 (N_2720,N_1516,N_2179);
xnor U2721 (N_2721,N_1811,N_1503);
xor U2722 (N_2722,N_1945,N_2227);
xnor U2723 (N_2723,N_1979,N_2201);
and U2724 (N_2724,N_2133,N_1711);
nand U2725 (N_2725,N_2005,N_2124);
xor U2726 (N_2726,N_2090,N_1841);
and U2727 (N_2727,N_1874,N_2097);
xnor U2728 (N_2728,N_1517,N_1565);
nor U2729 (N_2729,N_1915,N_2008);
nand U2730 (N_2730,N_1702,N_1557);
nor U2731 (N_2731,N_1785,N_2024);
nor U2732 (N_2732,N_1608,N_1757);
and U2733 (N_2733,N_1871,N_1996);
or U2734 (N_2734,N_1600,N_1814);
and U2735 (N_2735,N_2196,N_2050);
xnor U2736 (N_2736,N_1853,N_1904);
xnor U2737 (N_2737,N_1761,N_1801);
xor U2738 (N_2738,N_1611,N_1785);
nor U2739 (N_2739,N_1517,N_2131);
xor U2740 (N_2740,N_1861,N_1781);
or U2741 (N_2741,N_1643,N_1525);
nand U2742 (N_2742,N_1760,N_1916);
nand U2743 (N_2743,N_2098,N_1590);
nand U2744 (N_2744,N_1527,N_1751);
and U2745 (N_2745,N_1835,N_1560);
and U2746 (N_2746,N_1853,N_1681);
xnor U2747 (N_2747,N_1902,N_1821);
nand U2748 (N_2748,N_1943,N_1536);
nand U2749 (N_2749,N_2083,N_1867);
xor U2750 (N_2750,N_2042,N_1790);
and U2751 (N_2751,N_1667,N_2086);
nand U2752 (N_2752,N_2014,N_1848);
or U2753 (N_2753,N_2107,N_1575);
xnor U2754 (N_2754,N_1775,N_1568);
or U2755 (N_2755,N_1895,N_1892);
nand U2756 (N_2756,N_1843,N_2132);
nor U2757 (N_2757,N_2148,N_1936);
nor U2758 (N_2758,N_1583,N_1789);
nor U2759 (N_2759,N_2083,N_2063);
and U2760 (N_2760,N_1740,N_2126);
or U2761 (N_2761,N_1903,N_1884);
nand U2762 (N_2762,N_1752,N_1927);
xor U2763 (N_2763,N_2145,N_2114);
nand U2764 (N_2764,N_1768,N_1628);
and U2765 (N_2765,N_1884,N_1885);
nand U2766 (N_2766,N_2203,N_2167);
xnor U2767 (N_2767,N_2040,N_1705);
nor U2768 (N_2768,N_1770,N_1672);
and U2769 (N_2769,N_1759,N_2003);
nand U2770 (N_2770,N_1556,N_1755);
nand U2771 (N_2771,N_1755,N_1906);
and U2772 (N_2772,N_1868,N_1855);
xor U2773 (N_2773,N_1748,N_1704);
or U2774 (N_2774,N_1697,N_1846);
nand U2775 (N_2775,N_1727,N_1544);
nor U2776 (N_2776,N_2181,N_1512);
or U2777 (N_2777,N_1860,N_2043);
nand U2778 (N_2778,N_1659,N_1539);
or U2779 (N_2779,N_1591,N_1803);
xnor U2780 (N_2780,N_1928,N_1936);
nand U2781 (N_2781,N_1591,N_1750);
nor U2782 (N_2782,N_1881,N_2194);
xor U2783 (N_2783,N_1746,N_1627);
xor U2784 (N_2784,N_1743,N_1537);
nor U2785 (N_2785,N_2136,N_2217);
nor U2786 (N_2786,N_1998,N_1659);
and U2787 (N_2787,N_1835,N_1933);
and U2788 (N_2788,N_1810,N_2218);
nand U2789 (N_2789,N_1527,N_1892);
and U2790 (N_2790,N_1960,N_2163);
nand U2791 (N_2791,N_2034,N_1870);
nor U2792 (N_2792,N_1925,N_1801);
nand U2793 (N_2793,N_1732,N_1754);
and U2794 (N_2794,N_1934,N_1564);
or U2795 (N_2795,N_1925,N_2104);
xnor U2796 (N_2796,N_1744,N_1949);
and U2797 (N_2797,N_2119,N_1820);
or U2798 (N_2798,N_2011,N_1930);
nand U2799 (N_2799,N_2104,N_1785);
and U2800 (N_2800,N_1841,N_1517);
or U2801 (N_2801,N_1683,N_2243);
nor U2802 (N_2802,N_1686,N_1926);
nand U2803 (N_2803,N_2101,N_1764);
nor U2804 (N_2804,N_1742,N_1721);
or U2805 (N_2805,N_2096,N_2230);
and U2806 (N_2806,N_1708,N_2065);
xnor U2807 (N_2807,N_1645,N_1787);
nor U2808 (N_2808,N_1682,N_1793);
or U2809 (N_2809,N_1815,N_1572);
nor U2810 (N_2810,N_1560,N_1736);
xnor U2811 (N_2811,N_2228,N_2081);
nand U2812 (N_2812,N_1729,N_1604);
nor U2813 (N_2813,N_1952,N_2177);
nand U2814 (N_2814,N_2146,N_1936);
or U2815 (N_2815,N_2135,N_1600);
and U2816 (N_2816,N_2018,N_1617);
and U2817 (N_2817,N_2051,N_2108);
or U2818 (N_2818,N_1649,N_1751);
nand U2819 (N_2819,N_1909,N_2037);
nor U2820 (N_2820,N_2204,N_1683);
xnor U2821 (N_2821,N_1730,N_1972);
nor U2822 (N_2822,N_1636,N_1734);
xor U2823 (N_2823,N_1685,N_2104);
nor U2824 (N_2824,N_2047,N_1894);
nor U2825 (N_2825,N_2133,N_2181);
and U2826 (N_2826,N_1627,N_1597);
or U2827 (N_2827,N_1603,N_1696);
xor U2828 (N_2828,N_1889,N_1558);
and U2829 (N_2829,N_1909,N_2103);
or U2830 (N_2830,N_2175,N_1905);
nand U2831 (N_2831,N_2197,N_1745);
or U2832 (N_2832,N_1502,N_1909);
nand U2833 (N_2833,N_1811,N_1977);
or U2834 (N_2834,N_1959,N_2003);
and U2835 (N_2835,N_1826,N_1519);
or U2836 (N_2836,N_1535,N_1919);
and U2837 (N_2837,N_1589,N_1764);
xnor U2838 (N_2838,N_1676,N_1806);
nand U2839 (N_2839,N_2189,N_1758);
or U2840 (N_2840,N_1694,N_1876);
and U2841 (N_2841,N_1879,N_1904);
nor U2842 (N_2842,N_1988,N_1714);
xor U2843 (N_2843,N_1844,N_2069);
xor U2844 (N_2844,N_1687,N_2101);
and U2845 (N_2845,N_1820,N_2181);
nor U2846 (N_2846,N_1590,N_2230);
nand U2847 (N_2847,N_1805,N_2016);
nor U2848 (N_2848,N_1706,N_1816);
and U2849 (N_2849,N_1833,N_1866);
nor U2850 (N_2850,N_1939,N_1893);
xor U2851 (N_2851,N_1569,N_1819);
xor U2852 (N_2852,N_2061,N_2007);
or U2853 (N_2853,N_1511,N_1696);
nand U2854 (N_2854,N_2094,N_1529);
and U2855 (N_2855,N_1739,N_2104);
and U2856 (N_2856,N_1991,N_1975);
or U2857 (N_2857,N_2243,N_1645);
nor U2858 (N_2858,N_2078,N_1926);
nor U2859 (N_2859,N_1922,N_1752);
or U2860 (N_2860,N_1733,N_1903);
nor U2861 (N_2861,N_1754,N_1892);
or U2862 (N_2862,N_2183,N_2125);
or U2863 (N_2863,N_1915,N_1823);
and U2864 (N_2864,N_2169,N_1523);
nand U2865 (N_2865,N_2080,N_1585);
or U2866 (N_2866,N_2240,N_1518);
xnor U2867 (N_2867,N_2197,N_1934);
and U2868 (N_2868,N_1954,N_2118);
nor U2869 (N_2869,N_1617,N_2226);
nand U2870 (N_2870,N_1778,N_1933);
xor U2871 (N_2871,N_1986,N_2147);
and U2872 (N_2872,N_1827,N_1530);
nor U2873 (N_2873,N_1675,N_2182);
and U2874 (N_2874,N_2040,N_1672);
or U2875 (N_2875,N_1677,N_2114);
and U2876 (N_2876,N_2159,N_1899);
xnor U2877 (N_2877,N_2193,N_1975);
and U2878 (N_2878,N_1827,N_1994);
xnor U2879 (N_2879,N_1554,N_1976);
xor U2880 (N_2880,N_1503,N_1919);
xor U2881 (N_2881,N_2024,N_1816);
nand U2882 (N_2882,N_1739,N_2089);
nor U2883 (N_2883,N_2174,N_2064);
nand U2884 (N_2884,N_2138,N_2183);
nand U2885 (N_2885,N_1723,N_1519);
or U2886 (N_2886,N_2227,N_1842);
and U2887 (N_2887,N_1528,N_2024);
nand U2888 (N_2888,N_1952,N_1959);
and U2889 (N_2889,N_1978,N_2179);
nand U2890 (N_2890,N_1771,N_2206);
and U2891 (N_2891,N_2146,N_1719);
nor U2892 (N_2892,N_1866,N_1935);
and U2893 (N_2893,N_1605,N_2198);
nor U2894 (N_2894,N_2073,N_1855);
or U2895 (N_2895,N_1988,N_1711);
nand U2896 (N_2896,N_2049,N_1625);
and U2897 (N_2897,N_1787,N_1712);
nor U2898 (N_2898,N_1834,N_1948);
xor U2899 (N_2899,N_1588,N_1796);
and U2900 (N_2900,N_1634,N_1746);
or U2901 (N_2901,N_1987,N_2028);
or U2902 (N_2902,N_1624,N_2049);
nor U2903 (N_2903,N_1568,N_1911);
or U2904 (N_2904,N_1522,N_2214);
xor U2905 (N_2905,N_1853,N_1602);
or U2906 (N_2906,N_1780,N_1826);
or U2907 (N_2907,N_2122,N_1995);
nor U2908 (N_2908,N_1872,N_2133);
and U2909 (N_2909,N_2138,N_1917);
or U2910 (N_2910,N_1810,N_1532);
xor U2911 (N_2911,N_1933,N_1508);
or U2912 (N_2912,N_2192,N_1846);
nor U2913 (N_2913,N_1775,N_1579);
or U2914 (N_2914,N_1709,N_1762);
or U2915 (N_2915,N_1675,N_2138);
or U2916 (N_2916,N_1575,N_1625);
nor U2917 (N_2917,N_2048,N_2027);
and U2918 (N_2918,N_1607,N_1719);
nor U2919 (N_2919,N_1633,N_1952);
nand U2920 (N_2920,N_1589,N_1549);
nor U2921 (N_2921,N_1982,N_2056);
or U2922 (N_2922,N_1567,N_1955);
xor U2923 (N_2923,N_2223,N_1752);
or U2924 (N_2924,N_2107,N_2222);
or U2925 (N_2925,N_1978,N_1917);
and U2926 (N_2926,N_1865,N_2042);
nor U2927 (N_2927,N_2207,N_1660);
xor U2928 (N_2928,N_2227,N_1854);
and U2929 (N_2929,N_1928,N_1580);
nor U2930 (N_2930,N_1770,N_1938);
or U2931 (N_2931,N_1671,N_2187);
nand U2932 (N_2932,N_2120,N_1769);
or U2933 (N_2933,N_1518,N_2131);
nand U2934 (N_2934,N_2133,N_1661);
and U2935 (N_2935,N_1701,N_1928);
nor U2936 (N_2936,N_1825,N_2103);
nand U2937 (N_2937,N_1994,N_1556);
xor U2938 (N_2938,N_1558,N_1836);
and U2939 (N_2939,N_2190,N_1673);
xnor U2940 (N_2940,N_2030,N_1836);
nand U2941 (N_2941,N_1698,N_2109);
nor U2942 (N_2942,N_2179,N_1688);
nand U2943 (N_2943,N_1503,N_1914);
nor U2944 (N_2944,N_1601,N_2089);
xor U2945 (N_2945,N_1880,N_1983);
xor U2946 (N_2946,N_1947,N_2164);
nor U2947 (N_2947,N_1819,N_2076);
nand U2948 (N_2948,N_1621,N_2203);
xor U2949 (N_2949,N_1785,N_1549);
or U2950 (N_2950,N_2074,N_1899);
or U2951 (N_2951,N_2054,N_1576);
and U2952 (N_2952,N_1552,N_2028);
nand U2953 (N_2953,N_2052,N_1867);
xnor U2954 (N_2954,N_2194,N_1580);
or U2955 (N_2955,N_1556,N_2118);
or U2956 (N_2956,N_1811,N_2006);
nand U2957 (N_2957,N_1910,N_1699);
and U2958 (N_2958,N_1759,N_1896);
and U2959 (N_2959,N_1940,N_1591);
or U2960 (N_2960,N_2038,N_1985);
xnor U2961 (N_2961,N_1979,N_1522);
nand U2962 (N_2962,N_2228,N_1766);
nor U2963 (N_2963,N_1628,N_1907);
or U2964 (N_2964,N_2217,N_1898);
nand U2965 (N_2965,N_2153,N_1893);
or U2966 (N_2966,N_1715,N_1793);
nand U2967 (N_2967,N_2110,N_1700);
nor U2968 (N_2968,N_1822,N_1930);
xor U2969 (N_2969,N_1537,N_2120);
xnor U2970 (N_2970,N_2095,N_1797);
or U2971 (N_2971,N_1737,N_1770);
nand U2972 (N_2972,N_1505,N_1780);
nand U2973 (N_2973,N_1627,N_1970);
xor U2974 (N_2974,N_2074,N_1745);
xnor U2975 (N_2975,N_1878,N_1823);
nand U2976 (N_2976,N_2195,N_1800);
and U2977 (N_2977,N_1548,N_1950);
xnor U2978 (N_2978,N_2091,N_1997);
xnor U2979 (N_2979,N_1819,N_2096);
nand U2980 (N_2980,N_2150,N_2089);
xor U2981 (N_2981,N_1546,N_2238);
and U2982 (N_2982,N_1541,N_1676);
or U2983 (N_2983,N_2080,N_1525);
or U2984 (N_2984,N_2018,N_1874);
nand U2985 (N_2985,N_2152,N_1911);
nor U2986 (N_2986,N_1769,N_1625);
xor U2987 (N_2987,N_1789,N_2241);
and U2988 (N_2988,N_2211,N_1914);
nand U2989 (N_2989,N_1912,N_1570);
or U2990 (N_2990,N_2109,N_2248);
or U2991 (N_2991,N_1628,N_1641);
or U2992 (N_2992,N_2187,N_1575);
xor U2993 (N_2993,N_1923,N_1638);
and U2994 (N_2994,N_1599,N_1501);
nor U2995 (N_2995,N_1713,N_1548);
and U2996 (N_2996,N_1779,N_1735);
nand U2997 (N_2997,N_1909,N_2112);
nor U2998 (N_2998,N_2058,N_1764);
and U2999 (N_2999,N_2187,N_1571);
nor U3000 (N_3000,N_2363,N_2545);
nor U3001 (N_3001,N_2462,N_2272);
nor U3002 (N_3002,N_2427,N_2437);
or U3003 (N_3003,N_2292,N_2274);
xor U3004 (N_3004,N_2326,N_2617);
or U3005 (N_3005,N_2702,N_2487);
xnor U3006 (N_3006,N_2743,N_2745);
and U3007 (N_3007,N_2656,N_2932);
nand U3008 (N_3008,N_2468,N_2341);
xor U3009 (N_3009,N_2293,N_2831);
or U3010 (N_3010,N_2931,N_2692);
xor U3011 (N_3011,N_2637,N_2935);
and U3012 (N_3012,N_2420,N_2886);
or U3013 (N_3013,N_2898,N_2498);
xor U3014 (N_3014,N_2378,N_2574);
or U3015 (N_3015,N_2540,N_2747);
or U3016 (N_3016,N_2984,N_2955);
or U3017 (N_3017,N_2786,N_2628);
nor U3018 (N_3018,N_2734,N_2944);
xor U3019 (N_3019,N_2920,N_2839);
nor U3020 (N_3020,N_2602,N_2391);
xor U3021 (N_3021,N_2787,N_2871);
nand U3022 (N_3022,N_2549,N_2903);
nor U3023 (N_3023,N_2445,N_2496);
or U3024 (N_3024,N_2707,N_2968);
nand U3025 (N_3025,N_2926,N_2298);
nor U3026 (N_3026,N_2647,N_2824);
nand U3027 (N_3027,N_2946,N_2979);
and U3028 (N_3028,N_2792,N_2851);
xor U3029 (N_3029,N_2428,N_2603);
or U3030 (N_3030,N_2418,N_2362);
nor U3031 (N_3031,N_2845,N_2671);
nand U3032 (N_3032,N_2703,N_2969);
or U3033 (N_3033,N_2696,N_2648);
xor U3034 (N_3034,N_2957,N_2364);
nand U3035 (N_3035,N_2897,N_2535);
and U3036 (N_3036,N_2904,N_2988);
and U3037 (N_3037,N_2766,N_2520);
nor U3038 (N_3038,N_2728,N_2780);
and U3039 (N_3039,N_2515,N_2841);
or U3040 (N_3040,N_2982,N_2863);
xnor U3041 (N_3041,N_2365,N_2666);
xnor U3042 (N_3042,N_2807,N_2318);
nand U3043 (N_3043,N_2527,N_2473);
and U3044 (N_3044,N_2634,N_2736);
nand U3045 (N_3045,N_2694,N_2461);
or U3046 (N_3046,N_2853,N_2757);
nand U3047 (N_3047,N_2481,N_2429);
nand U3048 (N_3048,N_2361,N_2950);
or U3049 (N_3049,N_2679,N_2783);
or U3050 (N_3050,N_2744,N_2876);
and U3051 (N_3051,N_2608,N_2701);
nand U3052 (N_3052,N_2494,N_2353);
nand U3053 (N_3053,N_2902,N_2590);
nor U3054 (N_3054,N_2482,N_2392);
and U3055 (N_3055,N_2676,N_2887);
or U3056 (N_3056,N_2951,N_2870);
and U3057 (N_3057,N_2875,N_2862);
nand U3058 (N_3058,N_2421,N_2533);
and U3059 (N_3059,N_2251,N_2606);
or U3060 (N_3060,N_2463,N_2645);
and U3061 (N_3061,N_2624,N_2765);
or U3062 (N_3062,N_2397,N_2912);
or U3063 (N_3063,N_2328,N_2891);
xnor U3064 (N_3064,N_2594,N_2580);
or U3065 (N_3065,N_2877,N_2607);
and U3066 (N_3066,N_2819,N_2396);
nand U3067 (N_3067,N_2796,N_2682);
or U3068 (N_3068,N_2478,N_2906);
and U3069 (N_3069,N_2929,N_2779);
and U3070 (N_3070,N_2347,N_2416);
and U3071 (N_3071,N_2625,N_2714);
xnor U3072 (N_3072,N_2889,N_2384);
nor U3073 (N_3073,N_2810,N_2585);
nor U3074 (N_3074,N_2447,N_2812);
or U3075 (N_3075,N_2281,N_2453);
or U3076 (N_3076,N_2635,N_2699);
nand U3077 (N_3077,N_2866,N_2954);
nand U3078 (N_3078,N_2284,N_2333);
xor U3079 (N_3079,N_2826,N_2681);
and U3080 (N_3080,N_2630,N_2554);
xor U3081 (N_3081,N_2591,N_2941);
or U3082 (N_3082,N_2930,N_2458);
or U3083 (N_3083,N_2697,N_2961);
nor U3084 (N_3084,N_2509,N_2934);
xor U3085 (N_3085,N_2772,N_2868);
nor U3086 (N_3086,N_2255,N_2577);
xnor U3087 (N_3087,N_2755,N_2621);
nor U3088 (N_3088,N_2537,N_2507);
or U3089 (N_3089,N_2956,N_2578);
nor U3090 (N_3090,N_2704,N_2962);
or U3091 (N_3091,N_2252,N_2677);
nand U3092 (N_3092,N_2560,N_2389);
or U3093 (N_3093,N_2782,N_2813);
or U3094 (N_3094,N_2569,N_2484);
xor U3095 (N_3095,N_2804,N_2917);
nor U3096 (N_3096,N_2316,N_2282);
nor U3097 (N_3097,N_2401,N_2471);
and U3098 (N_3098,N_2500,N_2894);
or U3099 (N_3099,N_2966,N_2994);
nor U3100 (N_3100,N_2777,N_2631);
and U3101 (N_3101,N_2953,N_2357);
nor U3102 (N_3102,N_2583,N_2778);
nand U3103 (N_3103,N_2797,N_2505);
or U3104 (N_3104,N_2415,N_2693);
xnor U3105 (N_3105,N_2449,N_2752);
or U3106 (N_3106,N_2290,N_2352);
or U3107 (N_3107,N_2670,N_2986);
xor U3108 (N_3108,N_2869,N_2726);
nor U3109 (N_3109,N_2983,N_2687);
nor U3110 (N_3110,N_2469,N_2791);
nor U3111 (N_3111,N_2678,N_2618);
xor U3112 (N_3112,N_2366,N_2715);
nand U3113 (N_3113,N_2924,N_2788);
nand U3114 (N_3114,N_2426,N_2532);
xor U3115 (N_3115,N_2847,N_2856);
or U3116 (N_3116,N_2908,N_2399);
nand U3117 (N_3117,N_2651,N_2258);
xor U3118 (N_3118,N_2411,N_2980);
nand U3119 (N_3119,N_2900,N_2315);
nor U3120 (N_3120,N_2938,N_2673);
nand U3121 (N_3121,N_2838,N_2636);
or U3122 (N_3122,N_2661,N_2300);
or U3123 (N_3123,N_2700,N_2905);
xor U3124 (N_3124,N_2593,N_2754);
nand U3125 (N_3125,N_2414,N_2892);
nor U3126 (N_3126,N_2448,N_2288);
nor U3127 (N_3127,N_2959,N_2864);
xnor U3128 (N_3128,N_2561,N_2403);
nand U3129 (N_3129,N_2425,N_2525);
xor U3130 (N_3130,N_2340,N_2718);
or U3131 (N_3131,N_2417,N_2450);
and U3132 (N_3132,N_2762,N_2833);
or U3133 (N_3133,N_2658,N_2741);
nand U3134 (N_3134,N_2344,N_2665);
and U3135 (N_3135,N_2739,N_2512);
nand U3136 (N_3136,N_2301,N_2776);
and U3137 (N_3137,N_2719,N_2947);
nand U3138 (N_3138,N_2495,N_2354);
nand U3139 (N_3139,N_2873,N_2922);
nand U3140 (N_3140,N_2614,N_2332);
or U3141 (N_3141,N_2388,N_2250);
and U3142 (N_3142,N_2489,N_2963);
xor U3143 (N_3143,N_2269,N_2558);
and U3144 (N_3144,N_2570,N_2381);
xnor U3145 (N_3145,N_2668,N_2995);
xnor U3146 (N_3146,N_2749,N_2789);
and U3147 (N_3147,N_2914,N_2893);
or U3148 (N_3148,N_2557,N_2901);
or U3149 (N_3149,N_2441,N_2406);
xor U3150 (N_3150,N_2393,N_2548);
nand U3151 (N_3151,N_2379,N_2485);
nor U3152 (N_3152,N_2985,N_2708);
xor U3153 (N_3153,N_2620,N_2937);
or U3154 (N_3154,N_2395,N_2567);
and U3155 (N_3155,N_2475,N_2860);
nand U3156 (N_3156,N_2488,N_2992);
and U3157 (N_3157,N_2861,N_2918);
and U3158 (N_3158,N_2289,N_2433);
nor U3159 (N_3159,N_2576,N_2622);
nor U3160 (N_3160,N_2910,N_2773);
nand U3161 (N_3161,N_2802,N_2742);
xor U3162 (N_3162,N_2541,N_2880);
and U3163 (N_3163,N_2854,N_2817);
and U3164 (N_3164,N_2706,N_2711);
xor U3165 (N_3165,N_2402,N_2562);
or U3166 (N_3166,N_2615,N_2386);
xnor U3167 (N_3167,N_2977,N_2435);
or U3168 (N_3168,N_2368,N_2327);
nand U3169 (N_3169,N_2638,N_2836);
and U3170 (N_3170,N_2993,N_2827);
xnor U3171 (N_3171,N_2431,N_2360);
nor U3172 (N_3172,N_2837,N_2526);
xnor U3173 (N_3173,N_2952,N_2867);
nor U3174 (N_3174,N_2657,N_2476);
and U3175 (N_3175,N_2799,N_2271);
and U3176 (N_3176,N_2349,N_2551);
or U3177 (N_3177,N_2592,N_2304);
xnor U3178 (N_3178,N_2446,N_2305);
or U3179 (N_3179,N_2550,N_2434);
or U3180 (N_3180,N_2596,N_2502);
and U3181 (N_3181,N_2564,N_2555);
nand U3182 (N_3182,N_2848,N_2270);
and U3183 (N_3183,N_2948,N_2599);
nand U3184 (N_3184,N_2534,N_2474);
and U3185 (N_3185,N_2313,N_2419);
xor U3186 (N_3186,N_2761,N_2794);
nor U3187 (N_3187,N_2829,N_2283);
and U3188 (N_3188,N_2975,N_2663);
and U3189 (N_3189,N_2972,N_2949);
xor U3190 (N_3190,N_2430,N_2444);
xor U3191 (N_3191,N_2513,N_2933);
or U3192 (N_3192,N_2552,N_2286);
and U3193 (N_3193,N_2970,N_2543);
nor U3194 (N_3194,N_2523,N_2698);
xor U3195 (N_3195,N_2818,N_2565);
or U3196 (N_3196,N_2524,N_2964);
and U3197 (N_3197,N_2769,N_2273);
nor U3198 (N_3198,N_2967,N_2491);
and U3199 (N_3199,N_2840,N_2456);
and U3200 (N_3200,N_2413,N_2508);
xor U3201 (N_3201,N_2976,N_2639);
nand U3202 (N_3202,N_2601,N_2690);
xnor U3203 (N_3203,N_2990,N_2338);
and U3204 (N_3204,N_2834,N_2683);
nand U3205 (N_3205,N_2409,N_2732);
nor U3206 (N_3206,N_2531,N_2881);
nor U3207 (N_3207,N_2499,N_2811);
xor U3208 (N_3208,N_2613,N_2724);
and U3209 (N_3209,N_2459,N_2923);
and U3210 (N_3210,N_2303,N_2350);
nor U3211 (N_3211,N_2568,N_2571);
xnor U3212 (N_3212,N_2936,N_2597);
nand U3213 (N_3213,N_2264,N_2717);
and U3214 (N_3214,N_2644,N_2852);
nand U3215 (N_3215,N_2916,N_2586);
nor U3216 (N_3216,N_2844,N_2723);
nand U3217 (N_3217,N_2735,N_2521);
nor U3218 (N_3218,N_2722,N_2467);
xnor U3219 (N_3219,N_2510,N_2302);
xnor U3220 (N_3220,N_2928,N_2308);
and U3221 (N_3221,N_2945,N_2493);
nor U3222 (N_3222,N_2346,N_2314);
or U3223 (N_3223,N_2865,N_2254);
nand U3224 (N_3224,N_2942,N_2731);
and U3225 (N_3225,N_2958,N_2733);
nand U3226 (N_3226,N_2815,N_2774);
and U3227 (N_3227,N_2598,N_2767);
and U3228 (N_3228,N_2497,N_2784);
nor U3229 (N_3229,N_2334,N_2432);
or U3230 (N_3230,N_2842,N_2760);
nand U3231 (N_3231,N_2374,N_2859);
nand U3232 (N_3232,N_2530,N_2960);
xnor U3233 (N_3233,N_2372,N_2595);
or U3234 (N_3234,N_2654,N_2649);
nor U3235 (N_3235,N_2604,N_2987);
nand U3236 (N_3236,N_2351,N_2294);
or U3237 (N_3237,N_2822,N_2309);
nor U3238 (N_3238,N_2650,N_2331);
nor U3239 (N_3239,N_2600,N_2342);
or U3240 (N_3240,N_2609,N_2884);
nor U3241 (N_3241,N_2795,N_2882);
or U3242 (N_3242,N_2764,N_2472);
and U3243 (N_3243,N_2611,N_2311);
xnor U3244 (N_3244,N_2641,N_2801);
nand U3245 (N_3245,N_2410,N_2939);
nand U3246 (N_3246,N_2380,N_2684);
and U3247 (N_3247,N_2559,N_2816);
or U3248 (N_3248,N_2412,N_2720);
or U3249 (N_3249,N_2263,N_2763);
and U3250 (N_3250,N_2925,N_2490);
nand U3251 (N_3251,N_2883,N_2584);
nand U3252 (N_3252,N_2394,N_2878);
xor U3253 (N_3253,N_2820,N_2758);
nand U3254 (N_3254,N_2675,N_2846);
and U3255 (N_3255,N_2279,N_2291);
and U3256 (N_3256,N_2680,N_2642);
nand U3257 (N_3257,N_2909,N_2991);
xnor U3258 (N_3258,N_2632,N_2626);
and U3259 (N_3259,N_2573,N_2377);
nor U3260 (N_3260,N_2438,N_2770);
nand U3261 (N_3261,N_2973,N_2479);
or U3262 (N_3262,N_2927,N_2369);
xnor U3263 (N_3263,N_2287,N_2582);
or U3264 (N_3264,N_2725,N_2330);
xor U3265 (N_3265,N_2798,N_2756);
or U3266 (N_3266,N_2501,N_2268);
nor U3267 (N_3267,N_2655,N_2667);
xnor U3268 (N_3268,N_2439,N_2424);
and U3269 (N_3269,N_2506,N_2895);
and U3270 (N_3270,N_2809,N_2516);
nor U3271 (N_3271,N_2358,N_2771);
nand U3272 (N_3272,N_2662,N_2296);
xor U3273 (N_3273,N_2849,N_2610);
nand U3274 (N_3274,N_2278,N_2348);
and U3275 (N_3275,N_2581,N_2627);
xor U3276 (N_3276,N_2319,N_2996);
and U3277 (N_3277,N_2466,N_2913);
nand U3278 (N_3278,N_2383,N_2896);
nand U3279 (N_3279,N_2436,N_2262);
and U3280 (N_3280,N_2400,N_2978);
nand U3281 (N_3281,N_2835,N_2589);
nand U3282 (N_3282,N_2775,N_2404);
nor U3283 (N_3283,N_2814,N_2850);
and U3284 (N_3284,N_2710,N_2325);
nor U3285 (N_3285,N_2566,N_2919);
or U3286 (N_3286,N_2705,N_2253);
xor U3287 (N_3287,N_2750,N_2981);
xnor U3288 (N_3288,N_2669,N_2843);
nand U3289 (N_3289,N_2544,N_2518);
nand U3290 (N_3290,N_2423,N_2738);
nand U3291 (N_3291,N_2572,N_2806);
and U3292 (N_3292,N_2746,N_2373);
nand U3293 (N_3293,N_2385,N_2729);
xnor U3294 (N_3294,N_2921,N_2686);
and U3295 (N_3295,N_2874,N_2716);
nand U3296 (N_3296,N_2793,N_2538);
nor U3297 (N_3297,N_2260,N_2800);
xnor U3298 (N_3298,N_2299,N_2276);
xnor U3299 (N_3299,N_2588,N_2652);
xnor U3300 (N_3300,N_2387,N_2768);
nor U3301 (N_3301,N_2440,N_2971);
nand U3302 (N_3302,N_2587,N_2546);
nor U3303 (N_3303,N_2828,N_2256);
nand U3304 (N_3304,N_2257,N_2879);
or U3305 (N_3305,N_2336,N_2265);
xor U3306 (N_3306,N_2858,N_2748);
nor U3307 (N_3307,N_2989,N_2547);
and U3308 (N_3308,N_2855,N_2727);
nand U3309 (N_3309,N_2563,N_2371);
nand U3310 (N_3310,N_2522,N_2539);
nor U3311 (N_3311,N_2674,N_2266);
nand U3312 (N_3312,N_2899,N_2803);
and U3313 (N_3313,N_2872,N_2285);
xnor U3314 (N_3314,N_2261,N_2685);
nor U3315 (N_3315,N_2503,N_2721);
xnor U3316 (N_3316,N_2888,N_2355);
nand U3317 (N_3317,N_2633,N_2709);
nand U3318 (N_3318,N_2688,N_2823);
or U3319 (N_3319,N_2691,N_2825);
and U3320 (N_3320,N_2465,N_2443);
nor U3321 (N_3321,N_2375,N_2616);
and U3322 (N_3322,N_2343,N_2885);
nor U3323 (N_3323,N_2643,N_2422);
xnor U3324 (N_3324,N_2689,N_2297);
and U3325 (N_3325,N_2999,N_2275);
and U3326 (N_3326,N_2712,N_2464);
nand U3327 (N_3327,N_2277,N_2857);
nor U3328 (N_3328,N_2337,N_2259);
nor U3329 (N_3329,N_2907,N_2329);
nand U3330 (N_3330,N_2528,N_2367);
xor U3331 (N_3331,N_2821,N_2320);
or U3332 (N_3332,N_2306,N_2659);
and U3333 (N_3333,N_2805,N_2511);
and U3334 (N_3334,N_2408,N_2974);
nor U3335 (N_3335,N_2267,N_2890);
nand U3336 (N_3336,N_2830,N_2451);
and U3337 (N_3337,N_2519,N_2339);
nor U3338 (N_3338,N_2517,N_2660);
or U3339 (N_3339,N_2382,N_2442);
nor U3340 (N_3340,N_2737,N_2307);
nor U3341 (N_3341,N_2997,N_2321);
and U3342 (N_3342,N_2629,N_2943);
nand U3343 (N_3343,N_2529,N_2359);
and U3344 (N_3344,N_2457,N_2514);
nor U3345 (N_3345,N_2295,N_2455);
or U3346 (N_3346,N_2759,N_2965);
nand U3347 (N_3347,N_2713,N_2832);
xor U3348 (N_3348,N_2405,N_2390);
nand U3349 (N_3349,N_2730,N_2323);
and U3350 (N_3350,N_2407,N_2345);
xnor U3351 (N_3351,N_2480,N_2460);
nor U3352 (N_3352,N_2605,N_2751);
xor U3353 (N_3353,N_2317,N_2280);
nor U3354 (N_3354,N_2998,N_2612);
xor U3355 (N_3355,N_2483,N_2504);
nor U3356 (N_3356,N_2911,N_2623);
nand U3357 (N_3357,N_2370,N_2470);
xor U3358 (N_3358,N_2672,N_2322);
nor U3359 (N_3359,N_2398,N_2376);
and U3360 (N_3360,N_2790,N_2781);
or U3361 (N_3361,N_2356,N_2664);
and U3362 (N_3362,N_2575,N_2492);
and U3363 (N_3363,N_2653,N_2619);
and U3364 (N_3364,N_2753,N_2940);
xor U3365 (N_3365,N_2486,N_2646);
xor U3366 (N_3366,N_2312,N_2310);
xnor U3367 (N_3367,N_2785,N_2640);
or U3368 (N_3368,N_2542,N_2556);
xnor U3369 (N_3369,N_2454,N_2915);
nor U3370 (N_3370,N_2324,N_2477);
xnor U3371 (N_3371,N_2740,N_2695);
and U3372 (N_3372,N_2536,N_2335);
or U3373 (N_3373,N_2553,N_2452);
xor U3374 (N_3374,N_2808,N_2579);
xnor U3375 (N_3375,N_2840,N_2817);
and U3376 (N_3376,N_2883,N_2314);
nand U3377 (N_3377,N_2792,N_2904);
or U3378 (N_3378,N_2675,N_2554);
and U3379 (N_3379,N_2660,N_2931);
nor U3380 (N_3380,N_2493,N_2530);
nor U3381 (N_3381,N_2754,N_2636);
xor U3382 (N_3382,N_2940,N_2672);
nor U3383 (N_3383,N_2877,N_2968);
and U3384 (N_3384,N_2953,N_2446);
nand U3385 (N_3385,N_2700,N_2629);
nor U3386 (N_3386,N_2941,N_2304);
and U3387 (N_3387,N_2501,N_2689);
nor U3388 (N_3388,N_2723,N_2278);
nor U3389 (N_3389,N_2353,N_2822);
nor U3390 (N_3390,N_2369,N_2550);
nand U3391 (N_3391,N_2870,N_2794);
nor U3392 (N_3392,N_2893,N_2276);
and U3393 (N_3393,N_2476,N_2573);
and U3394 (N_3394,N_2523,N_2988);
xnor U3395 (N_3395,N_2319,N_2263);
nand U3396 (N_3396,N_2847,N_2457);
and U3397 (N_3397,N_2705,N_2793);
and U3398 (N_3398,N_2401,N_2669);
or U3399 (N_3399,N_2860,N_2932);
and U3400 (N_3400,N_2603,N_2323);
nor U3401 (N_3401,N_2598,N_2394);
and U3402 (N_3402,N_2866,N_2731);
nand U3403 (N_3403,N_2470,N_2560);
nor U3404 (N_3404,N_2486,N_2286);
or U3405 (N_3405,N_2370,N_2856);
xnor U3406 (N_3406,N_2801,N_2975);
and U3407 (N_3407,N_2583,N_2273);
or U3408 (N_3408,N_2592,N_2673);
nand U3409 (N_3409,N_2989,N_2978);
xor U3410 (N_3410,N_2949,N_2738);
or U3411 (N_3411,N_2272,N_2388);
nor U3412 (N_3412,N_2618,N_2278);
or U3413 (N_3413,N_2552,N_2962);
nand U3414 (N_3414,N_2693,N_2918);
nor U3415 (N_3415,N_2762,N_2690);
or U3416 (N_3416,N_2660,N_2984);
xnor U3417 (N_3417,N_2779,N_2558);
or U3418 (N_3418,N_2796,N_2714);
or U3419 (N_3419,N_2630,N_2827);
nand U3420 (N_3420,N_2289,N_2599);
or U3421 (N_3421,N_2421,N_2785);
and U3422 (N_3422,N_2449,N_2313);
xor U3423 (N_3423,N_2526,N_2772);
xnor U3424 (N_3424,N_2975,N_2768);
and U3425 (N_3425,N_2325,N_2250);
nor U3426 (N_3426,N_2797,N_2600);
nor U3427 (N_3427,N_2480,N_2604);
or U3428 (N_3428,N_2529,N_2900);
or U3429 (N_3429,N_2578,N_2320);
xor U3430 (N_3430,N_2326,N_2910);
xnor U3431 (N_3431,N_2569,N_2509);
and U3432 (N_3432,N_2326,N_2700);
and U3433 (N_3433,N_2732,N_2905);
nand U3434 (N_3434,N_2909,N_2919);
nor U3435 (N_3435,N_2435,N_2911);
or U3436 (N_3436,N_2899,N_2663);
and U3437 (N_3437,N_2868,N_2354);
and U3438 (N_3438,N_2987,N_2273);
nand U3439 (N_3439,N_2601,N_2517);
or U3440 (N_3440,N_2908,N_2299);
xnor U3441 (N_3441,N_2301,N_2285);
and U3442 (N_3442,N_2818,N_2400);
or U3443 (N_3443,N_2893,N_2387);
or U3444 (N_3444,N_2530,N_2848);
xnor U3445 (N_3445,N_2563,N_2693);
xnor U3446 (N_3446,N_2948,N_2804);
nor U3447 (N_3447,N_2745,N_2318);
or U3448 (N_3448,N_2645,N_2260);
nand U3449 (N_3449,N_2874,N_2697);
nand U3450 (N_3450,N_2918,N_2973);
or U3451 (N_3451,N_2895,N_2476);
and U3452 (N_3452,N_2337,N_2492);
xnor U3453 (N_3453,N_2929,N_2706);
or U3454 (N_3454,N_2305,N_2634);
or U3455 (N_3455,N_2617,N_2524);
xnor U3456 (N_3456,N_2652,N_2720);
or U3457 (N_3457,N_2785,N_2325);
xor U3458 (N_3458,N_2547,N_2798);
and U3459 (N_3459,N_2252,N_2721);
or U3460 (N_3460,N_2546,N_2837);
nand U3461 (N_3461,N_2928,N_2326);
or U3462 (N_3462,N_2400,N_2759);
nand U3463 (N_3463,N_2377,N_2596);
nand U3464 (N_3464,N_2610,N_2673);
nor U3465 (N_3465,N_2333,N_2849);
xor U3466 (N_3466,N_2419,N_2499);
nor U3467 (N_3467,N_2391,N_2316);
xnor U3468 (N_3468,N_2637,N_2518);
xnor U3469 (N_3469,N_2622,N_2818);
and U3470 (N_3470,N_2271,N_2813);
and U3471 (N_3471,N_2898,N_2662);
nor U3472 (N_3472,N_2798,N_2427);
xnor U3473 (N_3473,N_2697,N_2314);
xor U3474 (N_3474,N_2683,N_2984);
nand U3475 (N_3475,N_2985,N_2354);
or U3476 (N_3476,N_2360,N_2462);
xnor U3477 (N_3477,N_2536,N_2569);
nor U3478 (N_3478,N_2436,N_2470);
nor U3479 (N_3479,N_2946,N_2942);
nand U3480 (N_3480,N_2910,N_2735);
and U3481 (N_3481,N_2765,N_2502);
nand U3482 (N_3482,N_2573,N_2295);
and U3483 (N_3483,N_2998,N_2846);
xnor U3484 (N_3484,N_2963,N_2613);
xnor U3485 (N_3485,N_2587,N_2326);
nand U3486 (N_3486,N_2534,N_2579);
nand U3487 (N_3487,N_2522,N_2777);
or U3488 (N_3488,N_2861,N_2546);
or U3489 (N_3489,N_2599,N_2574);
and U3490 (N_3490,N_2305,N_2739);
and U3491 (N_3491,N_2743,N_2977);
and U3492 (N_3492,N_2852,N_2449);
and U3493 (N_3493,N_2889,N_2662);
or U3494 (N_3494,N_2884,N_2450);
and U3495 (N_3495,N_2896,N_2970);
and U3496 (N_3496,N_2877,N_2424);
nor U3497 (N_3497,N_2478,N_2986);
and U3498 (N_3498,N_2376,N_2886);
xnor U3499 (N_3499,N_2826,N_2571);
or U3500 (N_3500,N_2488,N_2395);
nand U3501 (N_3501,N_2343,N_2909);
nand U3502 (N_3502,N_2417,N_2529);
or U3503 (N_3503,N_2525,N_2271);
or U3504 (N_3504,N_2683,N_2958);
nand U3505 (N_3505,N_2762,N_2921);
nor U3506 (N_3506,N_2281,N_2674);
or U3507 (N_3507,N_2468,N_2451);
nor U3508 (N_3508,N_2500,N_2779);
xor U3509 (N_3509,N_2824,N_2462);
nor U3510 (N_3510,N_2828,N_2502);
xor U3511 (N_3511,N_2263,N_2377);
or U3512 (N_3512,N_2332,N_2481);
nand U3513 (N_3513,N_2596,N_2630);
or U3514 (N_3514,N_2794,N_2957);
nor U3515 (N_3515,N_2333,N_2900);
nor U3516 (N_3516,N_2387,N_2780);
nor U3517 (N_3517,N_2873,N_2811);
nand U3518 (N_3518,N_2400,N_2830);
nand U3519 (N_3519,N_2319,N_2391);
or U3520 (N_3520,N_2617,N_2710);
xor U3521 (N_3521,N_2350,N_2396);
or U3522 (N_3522,N_2454,N_2578);
and U3523 (N_3523,N_2922,N_2842);
or U3524 (N_3524,N_2458,N_2454);
nor U3525 (N_3525,N_2544,N_2395);
xnor U3526 (N_3526,N_2764,N_2536);
and U3527 (N_3527,N_2989,N_2788);
nor U3528 (N_3528,N_2492,N_2564);
nor U3529 (N_3529,N_2992,N_2558);
or U3530 (N_3530,N_2923,N_2770);
or U3531 (N_3531,N_2591,N_2409);
and U3532 (N_3532,N_2894,N_2743);
and U3533 (N_3533,N_2411,N_2848);
nor U3534 (N_3534,N_2446,N_2835);
xor U3535 (N_3535,N_2914,N_2543);
xnor U3536 (N_3536,N_2991,N_2630);
or U3537 (N_3537,N_2733,N_2663);
nand U3538 (N_3538,N_2828,N_2313);
nand U3539 (N_3539,N_2911,N_2644);
and U3540 (N_3540,N_2456,N_2366);
and U3541 (N_3541,N_2731,N_2839);
xor U3542 (N_3542,N_2910,N_2333);
nor U3543 (N_3543,N_2937,N_2405);
xor U3544 (N_3544,N_2283,N_2768);
nand U3545 (N_3545,N_2548,N_2727);
and U3546 (N_3546,N_2811,N_2641);
nor U3547 (N_3547,N_2759,N_2343);
and U3548 (N_3548,N_2483,N_2262);
nand U3549 (N_3549,N_2380,N_2359);
and U3550 (N_3550,N_2468,N_2669);
or U3551 (N_3551,N_2836,N_2888);
or U3552 (N_3552,N_2733,N_2776);
and U3553 (N_3553,N_2719,N_2552);
or U3554 (N_3554,N_2527,N_2420);
or U3555 (N_3555,N_2809,N_2333);
xnor U3556 (N_3556,N_2927,N_2763);
and U3557 (N_3557,N_2969,N_2796);
nand U3558 (N_3558,N_2284,N_2428);
and U3559 (N_3559,N_2385,N_2944);
and U3560 (N_3560,N_2792,N_2304);
nand U3561 (N_3561,N_2395,N_2965);
and U3562 (N_3562,N_2521,N_2379);
and U3563 (N_3563,N_2792,N_2295);
or U3564 (N_3564,N_2495,N_2855);
or U3565 (N_3565,N_2407,N_2986);
nor U3566 (N_3566,N_2912,N_2311);
nor U3567 (N_3567,N_2938,N_2806);
nand U3568 (N_3568,N_2351,N_2797);
and U3569 (N_3569,N_2396,N_2397);
and U3570 (N_3570,N_2684,N_2321);
or U3571 (N_3571,N_2463,N_2346);
or U3572 (N_3572,N_2782,N_2908);
xnor U3573 (N_3573,N_2940,N_2553);
and U3574 (N_3574,N_2565,N_2745);
xor U3575 (N_3575,N_2793,N_2653);
or U3576 (N_3576,N_2474,N_2699);
or U3577 (N_3577,N_2498,N_2710);
xor U3578 (N_3578,N_2954,N_2727);
nand U3579 (N_3579,N_2394,N_2872);
nor U3580 (N_3580,N_2305,N_2328);
or U3581 (N_3581,N_2335,N_2469);
nor U3582 (N_3582,N_2837,N_2701);
xnor U3583 (N_3583,N_2322,N_2880);
nor U3584 (N_3584,N_2437,N_2733);
nor U3585 (N_3585,N_2937,N_2501);
xnor U3586 (N_3586,N_2451,N_2307);
and U3587 (N_3587,N_2471,N_2388);
nor U3588 (N_3588,N_2982,N_2542);
nand U3589 (N_3589,N_2379,N_2939);
xnor U3590 (N_3590,N_2322,N_2312);
xor U3591 (N_3591,N_2811,N_2952);
xor U3592 (N_3592,N_2351,N_2302);
nor U3593 (N_3593,N_2258,N_2787);
and U3594 (N_3594,N_2914,N_2763);
nor U3595 (N_3595,N_2640,N_2838);
and U3596 (N_3596,N_2872,N_2463);
and U3597 (N_3597,N_2913,N_2865);
and U3598 (N_3598,N_2957,N_2608);
nor U3599 (N_3599,N_2370,N_2515);
or U3600 (N_3600,N_2383,N_2702);
nor U3601 (N_3601,N_2556,N_2614);
xnor U3602 (N_3602,N_2970,N_2462);
or U3603 (N_3603,N_2459,N_2627);
nand U3604 (N_3604,N_2786,N_2329);
and U3605 (N_3605,N_2371,N_2768);
and U3606 (N_3606,N_2504,N_2955);
nand U3607 (N_3607,N_2377,N_2457);
nand U3608 (N_3608,N_2799,N_2514);
and U3609 (N_3609,N_2921,N_2637);
and U3610 (N_3610,N_2884,N_2483);
nand U3611 (N_3611,N_2261,N_2970);
and U3612 (N_3612,N_2551,N_2698);
nand U3613 (N_3613,N_2331,N_2346);
xnor U3614 (N_3614,N_2308,N_2545);
xor U3615 (N_3615,N_2918,N_2964);
xor U3616 (N_3616,N_2838,N_2599);
xnor U3617 (N_3617,N_2857,N_2768);
or U3618 (N_3618,N_2565,N_2774);
or U3619 (N_3619,N_2328,N_2485);
nor U3620 (N_3620,N_2969,N_2486);
nand U3621 (N_3621,N_2459,N_2477);
xor U3622 (N_3622,N_2901,N_2645);
or U3623 (N_3623,N_2724,N_2311);
nand U3624 (N_3624,N_2968,N_2381);
or U3625 (N_3625,N_2347,N_2329);
xor U3626 (N_3626,N_2835,N_2814);
nand U3627 (N_3627,N_2479,N_2832);
nand U3628 (N_3628,N_2455,N_2641);
xnor U3629 (N_3629,N_2993,N_2639);
xnor U3630 (N_3630,N_2719,N_2266);
nand U3631 (N_3631,N_2542,N_2510);
nand U3632 (N_3632,N_2467,N_2841);
and U3633 (N_3633,N_2470,N_2771);
and U3634 (N_3634,N_2880,N_2864);
and U3635 (N_3635,N_2689,N_2290);
nor U3636 (N_3636,N_2968,N_2579);
or U3637 (N_3637,N_2519,N_2564);
and U3638 (N_3638,N_2757,N_2639);
and U3639 (N_3639,N_2268,N_2796);
and U3640 (N_3640,N_2634,N_2414);
nand U3641 (N_3641,N_2845,N_2868);
nand U3642 (N_3642,N_2818,N_2654);
nor U3643 (N_3643,N_2676,N_2712);
and U3644 (N_3644,N_2596,N_2296);
nand U3645 (N_3645,N_2558,N_2787);
or U3646 (N_3646,N_2299,N_2565);
xor U3647 (N_3647,N_2555,N_2884);
and U3648 (N_3648,N_2326,N_2793);
or U3649 (N_3649,N_2263,N_2389);
or U3650 (N_3650,N_2448,N_2773);
nor U3651 (N_3651,N_2488,N_2849);
nand U3652 (N_3652,N_2991,N_2775);
and U3653 (N_3653,N_2740,N_2848);
xnor U3654 (N_3654,N_2958,N_2508);
or U3655 (N_3655,N_2868,N_2886);
nand U3656 (N_3656,N_2899,N_2522);
nand U3657 (N_3657,N_2516,N_2337);
or U3658 (N_3658,N_2929,N_2917);
and U3659 (N_3659,N_2631,N_2643);
or U3660 (N_3660,N_2312,N_2635);
or U3661 (N_3661,N_2944,N_2572);
xnor U3662 (N_3662,N_2634,N_2894);
nand U3663 (N_3663,N_2489,N_2593);
nor U3664 (N_3664,N_2437,N_2320);
nor U3665 (N_3665,N_2553,N_2360);
and U3666 (N_3666,N_2416,N_2570);
or U3667 (N_3667,N_2271,N_2743);
or U3668 (N_3668,N_2554,N_2264);
nand U3669 (N_3669,N_2780,N_2863);
xnor U3670 (N_3670,N_2531,N_2258);
nand U3671 (N_3671,N_2991,N_2740);
nor U3672 (N_3672,N_2773,N_2964);
xnor U3673 (N_3673,N_2832,N_2391);
or U3674 (N_3674,N_2692,N_2581);
or U3675 (N_3675,N_2777,N_2491);
nor U3676 (N_3676,N_2537,N_2877);
and U3677 (N_3677,N_2267,N_2429);
nand U3678 (N_3678,N_2608,N_2402);
nor U3679 (N_3679,N_2259,N_2975);
nand U3680 (N_3680,N_2973,N_2688);
nor U3681 (N_3681,N_2553,N_2362);
or U3682 (N_3682,N_2960,N_2665);
or U3683 (N_3683,N_2530,N_2648);
nor U3684 (N_3684,N_2705,N_2840);
nand U3685 (N_3685,N_2511,N_2521);
nor U3686 (N_3686,N_2718,N_2286);
and U3687 (N_3687,N_2951,N_2918);
nand U3688 (N_3688,N_2859,N_2695);
nand U3689 (N_3689,N_2641,N_2322);
or U3690 (N_3690,N_2524,N_2369);
or U3691 (N_3691,N_2662,N_2908);
nand U3692 (N_3692,N_2509,N_2789);
nand U3693 (N_3693,N_2869,N_2731);
or U3694 (N_3694,N_2702,N_2679);
or U3695 (N_3695,N_2280,N_2713);
xor U3696 (N_3696,N_2664,N_2679);
and U3697 (N_3697,N_2709,N_2410);
or U3698 (N_3698,N_2593,N_2938);
or U3699 (N_3699,N_2952,N_2565);
nor U3700 (N_3700,N_2953,N_2376);
nand U3701 (N_3701,N_2910,N_2922);
nand U3702 (N_3702,N_2536,N_2334);
nor U3703 (N_3703,N_2783,N_2509);
nor U3704 (N_3704,N_2669,N_2760);
nand U3705 (N_3705,N_2963,N_2530);
xnor U3706 (N_3706,N_2434,N_2956);
nor U3707 (N_3707,N_2275,N_2666);
or U3708 (N_3708,N_2976,N_2978);
xor U3709 (N_3709,N_2864,N_2458);
nand U3710 (N_3710,N_2427,N_2396);
and U3711 (N_3711,N_2480,N_2340);
nor U3712 (N_3712,N_2589,N_2451);
and U3713 (N_3713,N_2525,N_2899);
nor U3714 (N_3714,N_2869,N_2997);
xnor U3715 (N_3715,N_2969,N_2645);
xor U3716 (N_3716,N_2586,N_2408);
or U3717 (N_3717,N_2608,N_2984);
nand U3718 (N_3718,N_2987,N_2785);
or U3719 (N_3719,N_2901,N_2579);
or U3720 (N_3720,N_2489,N_2454);
xnor U3721 (N_3721,N_2577,N_2446);
and U3722 (N_3722,N_2494,N_2394);
nand U3723 (N_3723,N_2313,N_2381);
nor U3724 (N_3724,N_2688,N_2723);
nor U3725 (N_3725,N_2392,N_2977);
xnor U3726 (N_3726,N_2361,N_2984);
nand U3727 (N_3727,N_2659,N_2549);
or U3728 (N_3728,N_2253,N_2493);
nand U3729 (N_3729,N_2740,N_2714);
and U3730 (N_3730,N_2274,N_2636);
nor U3731 (N_3731,N_2875,N_2826);
nand U3732 (N_3732,N_2253,N_2615);
and U3733 (N_3733,N_2417,N_2526);
xor U3734 (N_3734,N_2902,N_2289);
nand U3735 (N_3735,N_2415,N_2819);
and U3736 (N_3736,N_2393,N_2458);
nand U3737 (N_3737,N_2575,N_2426);
xnor U3738 (N_3738,N_2603,N_2661);
or U3739 (N_3739,N_2931,N_2314);
and U3740 (N_3740,N_2827,N_2932);
nand U3741 (N_3741,N_2776,N_2404);
and U3742 (N_3742,N_2413,N_2831);
xnor U3743 (N_3743,N_2830,N_2394);
nor U3744 (N_3744,N_2287,N_2609);
xor U3745 (N_3745,N_2342,N_2539);
or U3746 (N_3746,N_2524,N_2615);
and U3747 (N_3747,N_2659,N_2607);
and U3748 (N_3748,N_2826,N_2300);
nor U3749 (N_3749,N_2313,N_2543);
and U3750 (N_3750,N_3408,N_3708);
and U3751 (N_3751,N_3463,N_3658);
xnor U3752 (N_3752,N_3284,N_3088);
nor U3753 (N_3753,N_3069,N_3421);
or U3754 (N_3754,N_3445,N_3737);
nand U3755 (N_3755,N_3315,N_3612);
or U3756 (N_3756,N_3355,N_3185);
or U3757 (N_3757,N_3164,N_3034);
nand U3758 (N_3758,N_3079,N_3015);
nor U3759 (N_3759,N_3193,N_3622);
and U3760 (N_3760,N_3092,N_3167);
and U3761 (N_3761,N_3276,N_3738);
xnor U3762 (N_3762,N_3594,N_3639);
and U3763 (N_3763,N_3121,N_3110);
nor U3764 (N_3764,N_3203,N_3732);
nor U3765 (N_3765,N_3183,N_3000);
and U3766 (N_3766,N_3261,N_3649);
nor U3767 (N_3767,N_3288,N_3598);
nor U3768 (N_3768,N_3487,N_3652);
xor U3769 (N_3769,N_3456,N_3647);
xnor U3770 (N_3770,N_3389,N_3734);
xor U3771 (N_3771,N_3106,N_3506);
nand U3772 (N_3772,N_3483,N_3661);
nand U3773 (N_3773,N_3132,N_3250);
nor U3774 (N_3774,N_3429,N_3311);
or U3775 (N_3775,N_3577,N_3065);
or U3776 (N_3776,N_3716,N_3613);
xor U3777 (N_3777,N_3295,N_3749);
nand U3778 (N_3778,N_3631,N_3148);
or U3779 (N_3779,N_3133,N_3730);
xor U3780 (N_3780,N_3246,N_3702);
xor U3781 (N_3781,N_3144,N_3310);
nand U3782 (N_3782,N_3351,N_3266);
and U3783 (N_3783,N_3466,N_3071);
or U3784 (N_3784,N_3413,N_3275);
or U3785 (N_3785,N_3384,N_3517);
and U3786 (N_3786,N_3401,N_3255);
nand U3787 (N_3787,N_3320,N_3035);
nand U3788 (N_3788,N_3717,N_3538);
or U3789 (N_3789,N_3136,N_3012);
or U3790 (N_3790,N_3667,N_3592);
and U3791 (N_3791,N_3710,N_3509);
nand U3792 (N_3792,N_3201,N_3465);
or U3793 (N_3793,N_3241,N_3607);
nand U3794 (N_3794,N_3500,N_3321);
or U3795 (N_3795,N_3151,N_3655);
nand U3796 (N_3796,N_3686,N_3270);
or U3797 (N_3797,N_3377,N_3202);
or U3798 (N_3798,N_3245,N_3546);
xor U3799 (N_3799,N_3054,N_3388);
nand U3800 (N_3800,N_3265,N_3197);
or U3801 (N_3801,N_3171,N_3157);
or U3802 (N_3802,N_3214,N_3117);
nor U3803 (N_3803,N_3650,N_3539);
and U3804 (N_3804,N_3031,N_3172);
or U3805 (N_3805,N_3227,N_3610);
nand U3806 (N_3806,N_3623,N_3568);
nand U3807 (N_3807,N_3381,N_3282);
nand U3808 (N_3808,N_3478,N_3318);
nand U3809 (N_3809,N_3533,N_3238);
or U3810 (N_3810,N_3481,N_3375);
nor U3811 (N_3811,N_3343,N_3143);
nor U3812 (N_3812,N_3398,N_3096);
xnor U3813 (N_3813,N_3049,N_3208);
xor U3814 (N_3814,N_3097,N_3178);
or U3815 (N_3815,N_3490,N_3342);
or U3816 (N_3816,N_3672,N_3001);
nand U3817 (N_3817,N_3699,N_3244);
or U3818 (N_3818,N_3135,N_3109);
nand U3819 (N_3819,N_3234,N_3588);
and U3820 (N_3820,N_3681,N_3156);
nand U3821 (N_3821,N_3495,N_3551);
xnor U3822 (N_3822,N_3556,N_3047);
nor U3823 (N_3823,N_3552,N_3419);
or U3824 (N_3824,N_3298,N_3112);
and U3825 (N_3825,N_3361,N_3677);
xor U3826 (N_3826,N_3174,N_3119);
or U3827 (N_3827,N_3308,N_3187);
nor U3828 (N_3828,N_3573,N_3642);
nand U3829 (N_3829,N_3479,N_3258);
or U3830 (N_3830,N_3654,N_3070);
nand U3831 (N_3831,N_3532,N_3718);
xor U3832 (N_3832,N_3231,N_3470);
nand U3833 (N_3833,N_3285,N_3122);
or U3834 (N_3834,N_3491,N_3140);
xnor U3835 (N_3835,N_3191,N_3010);
or U3836 (N_3836,N_3476,N_3524);
or U3837 (N_3837,N_3528,N_3003);
nor U3838 (N_3838,N_3508,N_3219);
or U3839 (N_3839,N_3155,N_3640);
or U3840 (N_3840,N_3145,N_3141);
nand U3841 (N_3841,N_3198,N_3510);
and U3842 (N_3842,N_3370,N_3416);
xnor U3843 (N_3843,N_3696,N_3379);
nor U3844 (N_3844,N_3263,N_3606);
xor U3845 (N_3845,N_3366,N_3196);
nand U3846 (N_3846,N_3085,N_3303);
xor U3847 (N_3847,N_3582,N_3262);
and U3848 (N_3848,N_3345,N_3525);
and U3849 (N_3849,N_3444,N_3504);
nand U3850 (N_3850,N_3057,N_3259);
and U3851 (N_3851,N_3521,N_3352);
nand U3852 (N_3852,N_3492,N_3053);
and U3853 (N_3853,N_3014,N_3645);
and U3854 (N_3854,N_3382,N_3281);
nor U3855 (N_3855,N_3189,N_3665);
or U3856 (N_3856,N_3373,N_3216);
nand U3857 (N_3857,N_3104,N_3215);
and U3858 (N_3858,N_3602,N_3678);
nor U3859 (N_3859,N_3545,N_3499);
and U3860 (N_3860,N_3089,N_3073);
nand U3861 (N_3861,N_3460,N_3002);
xnor U3862 (N_3862,N_3022,N_3742);
nand U3863 (N_3863,N_3072,N_3101);
or U3864 (N_3864,N_3691,N_3411);
and U3865 (N_3865,N_3629,N_3357);
nand U3866 (N_3866,N_3032,N_3572);
or U3867 (N_3867,N_3668,N_3624);
or U3868 (N_3868,N_3591,N_3468);
xnor U3869 (N_3869,N_3125,N_3486);
nor U3870 (N_3870,N_3199,N_3387);
or U3871 (N_3871,N_3368,N_3605);
or U3872 (N_3872,N_3365,N_3230);
and U3873 (N_3873,N_3319,N_3192);
or U3874 (N_3874,N_3074,N_3697);
xor U3875 (N_3875,N_3596,N_3268);
xnor U3876 (N_3876,N_3426,N_3733);
nor U3877 (N_3877,N_3542,N_3673);
and U3878 (N_3878,N_3160,N_3360);
nor U3879 (N_3879,N_3098,N_3446);
xor U3880 (N_3880,N_3497,N_3676);
or U3881 (N_3881,N_3402,N_3438);
nor U3882 (N_3882,N_3496,N_3656);
or U3883 (N_3883,N_3204,N_3559);
or U3884 (N_3884,N_3693,N_3515);
xnor U3885 (N_3885,N_3522,N_3323);
nor U3886 (N_3886,N_3165,N_3128);
and U3887 (N_3887,N_3344,N_3747);
or U3888 (N_3888,N_3743,N_3184);
xnor U3889 (N_3889,N_3518,N_3130);
and U3890 (N_3890,N_3118,N_3564);
nand U3891 (N_3891,N_3217,N_3218);
and U3892 (N_3892,N_3584,N_3236);
nand U3893 (N_3893,N_3333,N_3286);
xor U3894 (N_3894,N_3166,N_3369);
and U3895 (N_3895,N_3719,N_3004);
and U3896 (N_3896,N_3213,N_3170);
and U3897 (N_3897,N_3207,N_3297);
xnor U3898 (N_3898,N_3735,N_3485);
or U3899 (N_3899,N_3279,N_3400);
nor U3900 (N_3900,N_3221,N_3086);
nor U3901 (N_3901,N_3038,N_3585);
nor U3902 (N_3902,N_3417,N_3701);
nand U3903 (N_3903,N_3626,N_3300);
or U3904 (N_3904,N_3354,N_3741);
nand U3905 (N_3905,N_3348,N_3048);
nand U3906 (N_3906,N_3461,N_3569);
nand U3907 (N_3907,N_3670,N_3115);
or U3908 (N_3908,N_3537,N_3636);
and U3909 (N_3909,N_3364,N_3008);
nor U3910 (N_3910,N_3340,N_3583);
nor U3911 (N_3911,N_3412,N_3181);
nand U3912 (N_3912,N_3042,N_3450);
nor U3913 (N_3913,N_3120,N_3422);
xnor U3914 (N_3914,N_3601,N_3313);
nand U3915 (N_3915,N_3587,N_3105);
nor U3916 (N_3916,N_3334,N_3484);
nand U3917 (N_3917,N_3036,N_3457);
and U3918 (N_3918,N_3494,N_3278);
or U3919 (N_3919,N_3580,N_3280);
and U3920 (N_3920,N_3359,N_3102);
or U3921 (N_3921,N_3025,N_3149);
nor U3922 (N_3922,N_3516,N_3033);
xnor U3923 (N_3923,N_3621,N_3688);
and U3924 (N_3924,N_3363,N_3332);
and U3925 (N_3925,N_3597,N_3062);
nand U3926 (N_3926,N_3338,N_3563);
or U3927 (N_3927,N_3698,N_3498);
and U3928 (N_3928,N_3414,N_3287);
or U3929 (N_3929,N_3346,N_3728);
xnor U3930 (N_3930,N_3253,N_3081);
and U3931 (N_3931,N_3627,N_3200);
nand U3932 (N_3932,N_3535,N_3099);
nor U3933 (N_3933,N_3409,N_3224);
xnor U3934 (N_3934,N_3644,N_3442);
nand U3935 (N_3935,N_3455,N_3740);
nand U3936 (N_3936,N_3195,N_3322);
nand U3937 (N_3937,N_3209,N_3159);
xnor U3938 (N_3938,N_3277,N_3679);
xor U3939 (N_3939,N_3653,N_3714);
and U3940 (N_3940,N_3557,N_3523);
nor U3941 (N_3941,N_3009,N_3043);
and U3942 (N_3942,N_3560,N_3242);
xnor U3943 (N_3943,N_3080,N_3294);
nand U3944 (N_3944,N_3558,N_3663);
and U3945 (N_3945,N_3383,N_3620);
nor U3946 (N_3946,N_3090,N_3152);
or U3947 (N_3947,N_3046,N_3020);
and U3948 (N_3948,N_3243,N_3076);
xor U3949 (N_3949,N_3643,N_3531);
xor U3950 (N_3950,N_3632,N_3571);
nand U3951 (N_3951,N_3177,N_3339);
nand U3952 (N_3952,N_3147,N_3347);
xor U3953 (N_3953,N_3611,N_3324);
nand U3954 (N_3954,N_3030,N_3599);
nor U3955 (N_3955,N_3452,N_3314);
and U3956 (N_3956,N_3595,N_3635);
nor U3957 (N_3957,N_3529,N_3252);
nor U3958 (N_3958,N_3007,N_3251);
xnor U3959 (N_3959,N_3700,N_3634);
nor U3960 (N_3960,N_3674,N_3427);
or U3961 (N_3961,N_3283,N_3331);
or U3962 (N_3962,N_3233,N_3307);
and U3963 (N_3963,N_3660,N_3436);
and U3964 (N_3964,N_3095,N_3739);
xnor U3965 (N_3965,N_3662,N_3441);
and U3966 (N_3966,N_3039,N_3059);
or U3967 (N_3967,N_3248,N_3330);
or U3968 (N_3968,N_3567,N_3619);
xor U3969 (N_3969,N_3256,N_3684);
nor U3970 (N_3970,N_3589,N_3378);
or U3971 (N_3971,N_3350,N_3091);
nand U3972 (N_3972,N_3296,N_3094);
or U3973 (N_3973,N_3513,N_3579);
or U3974 (N_3974,N_3267,N_3273);
nand U3975 (N_3975,N_3473,N_3705);
nand U3976 (N_3976,N_3407,N_3431);
nor U3977 (N_3977,N_3162,N_3045);
nor U3978 (N_3978,N_3325,N_3041);
or U3979 (N_3979,N_3188,N_3113);
or U3980 (N_3980,N_3464,N_3190);
xnor U3981 (N_3981,N_3423,N_3608);
nor U3982 (N_3982,N_3274,N_3169);
xor U3983 (N_3983,N_3711,N_3372);
xnor U3984 (N_3984,N_3664,N_3312);
and U3985 (N_3985,N_3462,N_3114);
or U3986 (N_3986,N_3194,N_3453);
and U3987 (N_3987,N_3058,N_3005);
xor U3988 (N_3988,N_3055,N_3428);
or U3989 (N_3989,N_3689,N_3139);
or U3990 (N_3990,N_3028,N_3129);
or U3991 (N_3991,N_3722,N_3240);
or U3992 (N_3992,N_3103,N_3126);
xnor U3993 (N_3993,N_3064,N_3385);
nor U3994 (N_3994,N_3353,N_3309);
and U3995 (N_3995,N_3482,N_3084);
and U3996 (N_3996,N_3182,N_3540);
nand U3997 (N_3997,N_3725,N_3707);
xor U3998 (N_3998,N_3328,N_3748);
or U3999 (N_3999,N_3430,N_3037);
nand U4000 (N_4000,N_3306,N_3618);
or U4001 (N_4001,N_3555,N_3726);
xor U4002 (N_4002,N_3023,N_3615);
or U4003 (N_4003,N_3593,N_3358);
and U4004 (N_4004,N_3335,N_3154);
and U4005 (N_4005,N_3530,N_3021);
and U4006 (N_4006,N_3396,N_3472);
nor U4007 (N_4007,N_3044,N_3637);
xnor U4008 (N_4008,N_3225,N_3474);
xnor U4009 (N_4009,N_3553,N_3675);
nor U4010 (N_4010,N_3503,N_3603);
nand U4011 (N_4011,N_3289,N_3405);
or U4012 (N_4012,N_3434,N_3056);
xor U4013 (N_4013,N_3609,N_3501);
or U4014 (N_4014,N_3235,N_3158);
nand U4015 (N_4015,N_3386,N_3488);
nand U4016 (N_4016,N_3168,N_3581);
xor U4017 (N_4017,N_3690,N_3349);
nand U4018 (N_4018,N_3443,N_3391);
nor U4019 (N_4019,N_3727,N_3514);
xor U4020 (N_4020,N_3301,N_3393);
xnor U4021 (N_4021,N_3570,N_3292);
and U4022 (N_4022,N_3052,N_3367);
and U4023 (N_4023,N_3083,N_3683);
xnor U4024 (N_4024,N_3247,N_3337);
xnor U4025 (N_4025,N_3223,N_3212);
xnor U4026 (N_4026,N_3692,N_3534);
or U4027 (N_4027,N_3406,N_3380);
nand U4028 (N_4028,N_3067,N_3019);
nor U4029 (N_4029,N_3415,N_3469);
nand U4030 (N_4030,N_3271,N_3590);
nand U4031 (N_4031,N_3399,N_3017);
and U4032 (N_4032,N_3574,N_3374);
xnor U4033 (N_4033,N_3395,N_3519);
nor U4034 (N_4034,N_3257,N_3228);
and U4035 (N_4035,N_3520,N_3024);
and U4036 (N_4036,N_3410,N_3075);
xor U4037 (N_4037,N_3467,N_3173);
xor U4038 (N_4038,N_3107,N_3006);
xnor U4039 (N_4039,N_3027,N_3543);
nor U4040 (N_4040,N_3682,N_3205);
and U4041 (N_4041,N_3186,N_3336);
and U4042 (N_4042,N_3418,N_3651);
or U4043 (N_4043,N_3299,N_3305);
xnor U4044 (N_4044,N_3249,N_3226);
and U4045 (N_4045,N_3694,N_3666);
nand U4046 (N_4046,N_3659,N_3736);
nor U4047 (N_4047,N_3695,N_3746);
nand U4048 (N_4048,N_3712,N_3329);
nand U4049 (N_4049,N_3146,N_3161);
or U4050 (N_4050,N_3512,N_3237);
or U4051 (N_4051,N_3548,N_3720);
nand U4052 (N_4052,N_3459,N_3142);
nand U4053 (N_4053,N_3745,N_3458);
or U4054 (N_4054,N_3327,N_3078);
or U4055 (N_4055,N_3051,N_3082);
nor U4056 (N_4056,N_3454,N_3547);
xnor U4057 (N_4057,N_3063,N_3575);
and U4058 (N_4058,N_3550,N_3554);
nand U4059 (N_4059,N_3604,N_3163);
and U4060 (N_4060,N_3424,N_3293);
nor U4061 (N_4061,N_3018,N_3511);
nor U4062 (N_4062,N_3404,N_3638);
nor U4063 (N_4063,N_3704,N_3437);
xnor U4064 (N_4064,N_3440,N_3077);
xor U4065 (N_4065,N_3527,N_3403);
and U4066 (N_4066,N_3180,N_3390);
nand U4067 (N_4067,N_3179,N_3526);
nor U4068 (N_4068,N_3290,N_3447);
and U4069 (N_4069,N_3600,N_3026);
nor U4070 (N_4070,N_3435,N_3502);
nor U4071 (N_4071,N_3731,N_3536);
nor U4072 (N_4072,N_3578,N_3721);
nand U4073 (N_4073,N_3123,N_3220);
nand U4074 (N_4074,N_3628,N_3229);
nor U4075 (N_4075,N_3232,N_3724);
xnor U4076 (N_4076,N_3566,N_3433);
or U4077 (N_4077,N_3657,N_3050);
nand U4078 (N_4078,N_3723,N_3100);
nand U4079 (N_4079,N_3371,N_3116);
xnor U4080 (N_4080,N_3493,N_3138);
nor U4081 (N_4081,N_3211,N_3068);
xor U4082 (N_4082,N_3124,N_3576);
or U4083 (N_4083,N_3477,N_3565);
and U4084 (N_4084,N_3254,N_3394);
and U4085 (N_4085,N_3210,N_3451);
or U4086 (N_4086,N_3304,N_3137);
or U4087 (N_4087,N_3016,N_3562);
nor U4088 (N_4088,N_3706,N_3641);
nor U4089 (N_4089,N_3561,N_3425);
nor U4090 (N_4090,N_3392,N_3013);
or U4091 (N_4091,N_3111,N_3449);
xnor U4092 (N_4092,N_3131,N_3029);
nor U4093 (N_4093,N_3630,N_3541);
nand U4094 (N_4094,N_3648,N_3397);
or U4095 (N_4095,N_3448,N_3087);
nand U4096 (N_4096,N_3544,N_3669);
or U4097 (N_4097,N_3264,N_3480);
nand U4098 (N_4098,N_3206,N_3150);
and U4099 (N_4099,N_3175,N_3376);
xor U4100 (N_4100,N_3685,N_3614);
and U4101 (N_4101,N_3066,N_3222);
nand U4102 (N_4102,N_3671,N_3471);
or U4103 (N_4103,N_3134,N_3439);
or U4104 (N_4104,N_3646,N_3302);
and U4105 (N_4105,N_3703,N_3633);
or U4106 (N_4106,N_3616,N_3729);
nand U4107 (N_4107,N_3617,N_3687);
or U4108 (N_4108,N_3420,N_3011);
xor U4109 (N_4109,N_3260,N_3127);
nor U4110 (N_4110,N_3680,N_3715);
xor U4111 (N_4111,N_3713,N_3176);
and U4112 (N_4112,N_3317,N_3326);
nor U4113 (N_4113,N_3061,N_3549);
nor U4114 (N_4114,N_3505,N_3709);
or U4115 (N_4115,N_3060,N_3316);
xnor U4116 (N_4116,N_3586,N_3341);
and U4117 (N_4117,N_3362,N_3291);
nand U4118 (N_4118,N_3239,N_3269);
or U4119 (N_4119,N_3153,N_3040);
nor U4120 (N_4120,N_3108,N_3272);
nor U4121 (N_4121,N_3507,N_3489);
nand U4122 (N_4122,N_3744,N_3356);
nand U4123 (N_4123,N_3432,N_3093);
nand U4124 (N_4124,N_3625,N_3475);
nand U4125 (N_4125,N_3232,N_3580);
xor U4126 (N_4126,N_3457,N_3465);
or U4127 (N_4127,N_3126,N_3355);
nor U4128 (N_4128,N_3063,N_3019);
or U4129 (N_4129,N_3200,N_3609);
or U4130 (N_4130,N_3614,N_3130);
xnor U4131 (N_4131,N_3022,N_3315);
nand U4132 (N_4132,N_3376,N_3543);
xnor U4133 (N_4133,N_3217,N_3538);
xor U4134 (N_4134,N_3596,N_3365);
and U4135 (N_4135,N_3205,N_3382);
and U4136 (N_4136,N_3612,N_3335);
nand U4137 (N_4137,N_3702,N_3714);
and U4138 (N_4138,N_3624,N_3529);
nor U4139 (N_4139,N_3679,N_3271);
or U4140 (N_4140,N_3267,N_3107);
or U4141 (N_4141,N_3002,N_3163);
xor U4142 (N_4142,N_3644,N_3524);
or U4143 (N_4143,N_3304,N_3651);
nor U4144 (N_4144,N_3065,N_3746);
nand U4145 (N_4145,N_3000,N_3693);
and U4146 (N_4146,N_3034,N_3274);
nor U4147 (N_4147,N_3223,N_3202);
xor U4148 (N_4148,N_3149,N_3544);
xnor U4149 (N_4149,N_3376,N_3636);
nand U4150 (N_4150,N_3397,N_3135);
nor U4151 (N_4151,N_3194,N_3703);
and U4152 (N_4152,N_3602,N_3277);
and U4153 (N_4153,N_3586,N_3215);
nand U4154 (N_4154,N_3019,N_3625);
xor U4155 (N_4155,N_3320,N_3117);
nand U4156 (N_4156,N_3276,N_3347);
or U4157 (N_4157,N_3534,N_3225);
nand U4158 (N_4158,N_3338,N_3038);
nor U4159 (N_4159,N_3224,N_3625);
xor U4160 (N_4160,N_3034,N_3698);
or U4161 (N_4161,N_3147,N_3340);
nand U4162 (N_4162,N_3289,N_3745);
and U4163 (N_4163,N_3027,N_3560);
and U4164 (N_4164,N_3162,N_3033);
nor U4165 (N_4165,N_3431,N_3509);
nand U4166 (N_4166,N_3528,N_3554);
xnor U4167 (N_4167,N_3521,N_3632);
xor U4168 (N_4168,N_3438,N_3506);
nand U4169 (N_4169,N_3464,N_3738);
or U4170 (N_4170,N_3165,N_3178);
or U4171 (N_4171,N_3110,N_3202);
nor U4172 (N_4172,N_3726,N_3205);
nor U4173 (N_4173,N_3071,N_3531);
nand U4174 (N_4174,N_3499,N_3491);
nand U4175 (N_4175,N_3747,N_3354);
or U4176 (N_4176,N_3707,N_3494);
nor U4177 (N_4177,N_3028,N_3714);
xor U4178 (N_4178,N_3409,N_3683);
nand U4179 (N_4179,N_3148,N_3336);
or U4180 (N_4180,N_3506,N_3465);
nand U4181 (N_4181,N_3437,N_3277);
nand U4182 (N_4182,N_3601,N_3061);
or U4183 (N_4183,N_3086,N_3441);
xor U4184 (N_4184,N_3121,N_3549);
xnor U4185 (N_4185,N_3474,N_3312);
nand U4186 (N_4186,N_3577,N_3253);
nand U4187 (N_4187,N_3469,N_3640);
nand U4188 (N_4188,N_3663,N_3194);
xnor U4189 (N_4189,N_3160,N_3140);
or U4190 (N_4190,N_3276,N_3504);
nor U4191 (N_4191,N_3615,N_3382);
nor U4192 (N_4192,N_3584,N_3544);
and U4193 (N_4193,N_3050,N_3242);
or U4194 (N_4194,N_3201,N_3236);
nor U4195 (N_4195,N_3576,N_3095);
and U4196 (N_4196,N_3417,N_3357);
and U4197 (N_4197,N_3032,N_3017);
nor U4198 (N_4198,N_3721,N_3673);
xor U4199 (N_4199,N_3266,N_3055);
or U4200 (N_4200,N_3117,N_3193);
nor U4201 (N_4201,N_3321,N_3607);
nand U4202 (N_4202,N_3465,N_3212);
and U4203 (N_4203,N_3670,N_3710);
nor U4204 (N_4204,N_3264,N_3417);
xor U4205 (N_4205,N_3444,N_3501);
and U4206 (N_4206,N_3035,N_3529);
and U4207 (N_4207,N_3023,N_3470);
nand U4208 (N_4208,N_3372,N_3564);
or U4209 (N_4209,N_3704,N_3527);
nor U4210 (N_4210,N_3004,N_3148);
or U4211 (N_4211,N_3291,N_3435);
nor U4212 (N_4212,N_3406,N_3091);
xnor U4213 (N_4213,N_3734,N_3694);
nor U4214 (N_4214,N_3674,N_3599);
nor U4215 (N_4215,N_3618,N_3520);
nand U4216 (N_4216,N_3330,N_3720);
xnor U4217 (N_4217,N_3270,N_3122);
and U4218 (N_4218,N_3481,N_3147);
nand U4219 (N_4219,N_3268,N_3162);
xor U4220 (N_4220,N_3422,N_3227);
or U4221 (N_4221,N_3249,N_3182);
nor U4222 (N_4222,N_3637,N_3457);
xnor U4223 (N_4223,N_3059,N_3470);
nand U4224 (N_4224,N_3133,N_3303);
and U4225 (N_4225,N_3102,N_3054);
and U4226 (N_4226,N_3331,N_3417);
xor U4227 (N_4227,N_3662,N_3448);
and U4228 (N_4228,N_3275,N_3148);
or U4229 (N_4229,N_3420,N_3351);
or U4230 (N_4230,N_3739,N_3610);
and U4231 (N_4231,N_3477,N_3272);
or U4232 (N_4232,N_3384,N_3074);
and U4233 (N_4233,N_3166,N_3201);
and U4234 (N_4234,N_3422,N_3611);
nor U4235 (N_4235,N_3696,N_3113);
and U4236 (N_4236,N_3600,N_3575);
and U4237 (N_4237,N_3392,N_3678);
and U4238 (N_4238,N_3248,N_3006);
xor U4239 (N_4239,N_3630,N_3669);
nor U4240 (N_4240,N_3539,N_3383);
nor U4241 (N_4241,N_3604,N_3164);
and U4242 (N_4242,N_3001,N_3104);
xor U4243 (N_4243,N_3029,N_3203);
nor U4244 (N_4244,N_3327,N_3095);
xor U4245 (N_4245,N_3628,N_3651);
nand U4246 (N_4246,N_3588,N_3321);
nand U4247 (N_4247,N_3202,N_3050);
or U4248 (N_4248,N_3664,N_3187);
nand U4249 (N_4249,N_3440,N_3677);
or U4250 (N_4250,N_3028,N_3671);
nand U4251 (N_4251,N_3715,N_3145);
and U4252 (N_4252,N_3620,N_3152);
nand U4253 (N_4253,N_3412,N_3232);
nand U4254 (N_4254,N_3569,N_3617);
and U4255 (N_4255,N_3035,N_3329);
nor U4256 (N_4256,N_3235,N_3511);
and U4257 (N_4257,N_3253,N_3535);
nor U4258 (N_4258,N_3090,N_3610);
nand U4259 (N_4259,N_3143,N_3372);
and U4260 (N_4260,N_3507,N_3134);
xnor U4261 (N_4261,N_3152,N_3676);
or U4262 (N_4262,N_3537,N_3695);
nand U4263 (N_4263,N_3429,N_3198);
and U4264 (N_4264,N_3474,N_3483);
xor U4265 (N_4265,N_3652,N_3111);
nor U4266 (N_4266,N_3102,N_3175);
nor U4267 (N_4267,N_3013,N_3722);
or U4268 (N_4268,N_3645,N_3056);
or U4269 (N_4269,N_3276,N_3432);
nand U4270 (N_4270,N_3523,N_3592);
nand U4271 (N_4271,N_3038,N_3399);
nor U4272 (N_4272,N_3123,N_3064);
and U4273 (N_4273,N_3052,N_3168);
or U4274 (N_4274,N_3122,N_3589);
nand U4275 (N_4275,N_3599,N_3726);
or U4276 (N_4276,N_3354,N_3247);
or U4277 (N_4277,N_3466,N_3536);
xor U4278 (N_4278,N_3673,N_3159);
and U4279 (N_4279,N_3056,N_3095);
or U4280 (N_4280,N_3493,N_3026);
or U4281 (N_4281,N_3378,N_3053);
nand U4282 (N_4282,N_3132,N_3209);
nand U4283 (N_4283,N_3011,N_3702);
nand U4284 (N_4284,N_3467,N_3409);
nand U4285 (N_4285,N_3201,N_3701);
nor U4286 (N_4286,N_3454,N_3382);
and U4287 (N_4287,N_3440,N_3141);
or U4288 (N_4288,N_3612,N_3046);
nor U4289 (N_4289,N_3336,N_3509);
xor U4290 (N_4290,N_3620,N_3281);
xnor U4291 (N_4291,N_3700,N_3527);
nand U4292 (N_4292,N_3722,N_3212);
nor U4293 (N_4293,N_3460,N_3655);
or U4294 (N_4294,N_3747,N_3462);
nor U4295 (N_4295,N_3010,N_3664);
nand U4296 (N_4296,N_3072,N_3331);
or U4297 (N_4297,N_3615,N_3276);
nor U4298 (N_4298,N_3547,N_3556);
nor U4299 (N_4299,N_3375,N_3004);
nor U4300 (N_4300,N_3504,N_3435);
and U4301 (N_4301,N_3509,N_3227);
xor U4302 (N_4302,N_3571,N_3372);
nand U4303 (N_4303,N_3557,N_3748);
xnor U4304 (N_4304,N_3662,N_3537);
and U4305 (N_4305,N_3193,N_3517);
xnor U4306 (N_4306,N_3607,N_3260);
or U4307 (N_4307,N_3389,N_3192);
and U4308 (N_4308,N_3112,N_3187);
or U4309 (N_4309,N_3701,N_3526);
nand U4310 (N_4310,N_3728,N_3663);
nor U4311 (N_4311,N_3287,N_3283);
nor U4312 (N_4312,N_3328,N_3429);
and U4313 (N_4313,N_3002,N_3215);
nor U4314 (N_4314,N_3033,N_3153);
nand U4315 (N_4315,N_3722,N_3667);
nand U4316 (N_4316,N_3296,N_3051);
nor U4317 (N_4317,N_3693,N_3092);
nor U4318 (N_4318,N_3646,N_3012);
and U4319 (N_4319,N_3718,N_3568);
or U4320 (N_4320,N_3519,N_3641);
nor U4321 (N_4321,N_3371,N_3561);
nand U4322 (N_4322,N_3014,N_3401);
nor U4323 (N_4323,N_3201,N_3242);
and U4324 (N_4324,N_3372,N_3240);
and U4325 (N_4325,N_3421,N_3740);
xor U4326 (N_4326,N_3121,N_3732);
xor U4327 (N_4327,N_3410,N_3659);
xor U4328 (N_4328,N_3370,N_3316);
nand U4329 (N_4329,N_3657,N_3683);
and U4330 (N_4330,N_3478,N_3747);
and U4331 (N_4331,N_3416,N_3413);
and U4332 (N_4332,N_3247,N_3529);
xnor U4333 (N_4333,N_3699,N_3243);
or U4334 (N_4334,N_3018,N_3455);
nand U4335 (N_4335,N_3331,N_3419);
and U4336 (N_4336,N_3462,N_3085);
or U4337 (N_4337,N_3262,N_3498);
nor U4338 (N_4338,N_3742,N_3505);
or U4339 (N_4339,N_3050,N_3514);
nand U4340 (N_4340,N_3163,N_3031);
xor U4341 (N_4341,N_3669,N_3587);
and U4342 (N_4342,N_3528,N_3230);
nand U4343 (N_4343,N_3022,N_3565);
and U4344 (N_4344,N_3199,N_3061);
nor U4345 (N_4345,N_3423,N_3164);
or U4346 (N_4346,N_3682,N_3706);
nor U4347 (N_4347,N_3463,N_3498);
or U4348 (N_4348,N_3006,N_3227);
nor U4349 (N_4349,N_3513,N_3148);
or U4350 (N_4350,N_3248,N_3478);
and U4351 (N_4351,N_3546,N_3164);
xnor U4352 (N_4352,N_3601,N_3475);
xor U4353 (N_4353,N_3388,N_3376);
xnor U4354 (N_4354,N_3250,N_3074);
nand U4355 (N_4355,N_3718,N_3075);
or U4356 (N_4356,N_3506,N_3246);
nor U4357 (N_4357,N_3735,N_3744);
nand U4358 (N_4358,N_3194,N_3030);
nand U4359 (N_4359,N_3016,N_3008);
nand U4360 (N_4360,N_3394,N_3551);
nand U4361 (N_4361,N_3574,N_3376);
and U4362 (N_4362,N_3081,N_3547);
nand U4363 (N_4363,N_3154,N_3023);
xor U4364 (N_4364,N_3590,N_3037);
and U4365 (N_4365,N_3106,N_3726);
xnor U4366 (N_4366,N_3384,N_3493);
and U4367 (N_4367,N_3194,N_3740);
and U4368 (N_4368,N_3333,N_3152);
nand U4369 (N_4369,N_3327,N_3117);
nor U4370 (N_4370,N_3113,N_3620);
xnor U4371 (N_4371,N_3469,N_3287);
or U4372 (N_4372,N_3539,N_3150);
xnor U4373 (N_4373,N_3012,N_3280);
nand U4374 (N_4374,N_3304,N_3162);
nand U4375 (N_4375,N_3041,N_3147);
or U4376 (N_4376,N_3366,N_3125);
xor U4377 (N_4377,N_3507,N_3260);
and U4378 (N_4378,N_3358,N_3504);
or U4379 (N_4379,N_3611,N_3452);
or U4380 (N_4380,N_3353,N_3479);
or U4381 (N_4381,N_3360,N_3712);
nand U4382 (N_4382,N_3694,N_3171);
xnor U4383 (N_4383,N_3402,N_3284);
nor U4384 (N_4384,N_3464,N_3006);
and U4385 (N_4385,N_3482,N_3515);
and U4386 (N_4386,N_3677,N_3194);
nor U4387 (N_4387,N_3429,N_3269);
and U4388 (N_4388,N_3526,N_3138);
nand U4389 (N_4389,N_3071,N_3705);
nor U4390 (N_4390,N_3279,N_3150);
or U4391 (N_4391,N_3347,N_3694);
xor U4392 (N_4392,N_3559,N_3602);
and U4393 (N_4393,N_3422,N_3519);
and U4394 (N_4394,N_3234,N_3653);
or U4395 (N_4395,N_3213,N_3105);
xnor U4396 (N_4396,N_3016,N_3234);
nand U4397 (N_4397,N_3152,N_3047);
nor U4398 (N_4398,N_3575,N_3080);
nand U4399 (N_4399,N_3540,N_3453);
nor U4400 (N_4400,N_3099,N_3202);
nor U4401 (N_4401,N_3081,N_3461);
xnor U4402 (N_4402,N_3741,N_3568);
nor U4403 (N_4403,N_3531,N_3642);
nor U4404 (N_4404,N_3271,N_3163);
and U4405 (N_4405,N_3306,N_3659);
and U4406 (N_4406,N_3408,N_3681);
and U4407 (N_4407,N_3430,N_3537);
xor U4408 (N_4408,N_3733,N_3410);
or U4409 (N_4409,N_3444,N_3040);
xor U4410 (N_4410,N_3121,N_3578);
or U4411 (N_4411,N_3330,N_3041);
nor U4412 (N_4412,N_3250,N_3147);
nand U4413 (N_4413,N_3557,N_3566);
nand U4414 (N_4414,N_3250,N_3653);
nor U4415 (N_4415,N_3105,N_3550);
nand U4416 (N_4416,N_3571,N_3218);
and U4417 (N_4417,N_3509,N_3391);
nand U4418 (N_4418,N_3465,N_3214);
nand U4419 (N_4419,N_3470,N_3578);
nor U4420 (N_4420,N_3729,N_3741);
xor U4421 (N_4421,N_3099,N_3741);
or U4422 (N_4422,N_3522,N_3507);
or U4423 (N_4423,N_3266,N_3224);
and U4424 (N_4424,N_3607,N_3614);
xor U4425 (N_4425,N_3233,N_3021);
nand U4426 (N_4426,N_3551,N_3736);
nor U4427 (N_4427,N_3040,N_3339);
nor U4428 (N_4428,N_3603,N_3167);
nand U4429 (N_4429,N_3124,N_3257);
and U4430 (N_4430,N_3689,N_3043);
xnor U4431 (N_4431,N_3453,N_3407);
nor U4432 (N_4432,N_3625,N_3330);
and U4433 (N_4433,N_3132,N_3155);
or U4434 (N_4434,N_3452,N_3675);
or U4435 (N_4435,N_3145,N_3004);
nand U4436 (N_4436,N_3193,N_3417);
and U4437 (N_4437,N_3198,N_3341);
or U4438 (N_4438,N_3082,N_3449);
or U4439 (N_4439,N_3143,N_3469);
or U4440 (N_4440,N_3476,N_3671);
xor U4441 (N_4441,N_3001,N_3581);
nor U4442 (N_4442,N_3705,N_3698);
nor U4443 (N_4443,N_3532,N_3430);
nor U4444 (N_4444,N_3554,N_3613);
nand U4445 (N_4445,N_3533,N_3346);
and U4446 (N_4446,N_3029,N_3212);
nand U4447 (N_4447,N_3338,N_3578);
nand U4448 (N_4448,N_3691,N_3291);
and U4449 (N_4449,N_3514,N_3594);
nor U4450 (N_4450,N_3378,N_3398);
or U4451 (N_4451,N_3485,N_3604);
or U4452 (N_4452,N_3491,N_3142);
and U4453 (N_4453,N_3624,N_3384);
or U4454 (N_4454,N_3006,N_3268);
or U4455 (N_4455,N_3694,N_3250);
and U4456 (N_4456,N_3721,N_3068);
nand U4457 (N_4457,N_3604,N_3267);
nor U4458 (N_4458,N_3208,N_3206);
xnor U4459 (N_4459,N_3229,N_3425);
or U4460 (N_4460,N_3035,N_3031);
xor U4461 (N_4461,N_3495,N_3395);
and U4462 (N_4462,N_3346,N_3241);
nor U4463 (N_4463,N_3123,N_3748);
xnor U4464 (N_4464,N_3357,N_3203);
or U4465 (N_4465,N_3453,N_3604);
or U4466 (N_4466,N_3077,N_3695);
nor U4467 (N_4467,N_3225,N_3429);
and U4468 (N_4468,N_3166,N_3630);
and U4469 (N_4469,N_3608,N_3027);
or U4470 (N_4470,N_3626,N_3732);
xnor U4471 (N_4471,N_3727,N_3128);
nor U4472 (N_4472,N_3666,N_3445);
and U4473 (N_4473,N_3659,N_3364);
xor U4474 (N_4474,N_3656,N_3226);
or U4475 (N_4475,N_3028,N_3292);
and U4476 (N_4476,N_3173,N_3497);
nand U4477 (N_4477,N_3632,N_3593);
and U4478 (N_4478,N_3284,N_3368);
xor U4479 (N_4479,N_3544,N_3670);
or U4480 (N_4480,N_3404,N_3744);
and U4481 (N_4481,N_3180,N_3113);
or U4482 (N_4482,N_3702,N_3449);
nor U4483 (N_4483,N_3531,N_3074);
and U4484 (N_4484,N_3212,N_3648);
nand U4485 (N_4485,N_3223,N_3114);
or U4486 (N_4486,N_3322,N_3449);
and U4487 (N_4487,N_3096,N_3081);
or U4488 (N_4488,N_3499,N_3182);
and U4489 (N_4489,N_3385,N_3209);
or U4490 (N_4490,N_3050,N_3627);
and U4491 (N_4491,N_3341,N_3688);
nand U4492 (N_4492,N_3564,N_3190);
or U4493 (N_4493,N_3245,N_3345);
and U4494 (N_4494,N_3178,N_3361);
or U4495 (N_4495,N_3227,N_3223);
xor U4496 (N_4496,N_3408,N_3039);
nand U4497 (N_4497,N_3287,N_3607);
xor U4498 (N_4498,N_3094,N_3112);
xor U4499 (N_4499,N_3714,N_3693);
xnor U4500 (N_4500,N_3821,N_3766);
xor U4501 (N_4501,N_4157,N_4192);
and U4502 (N_4502,N_4374,N_4450);
nor U4503 (N_4503,N_4480,N_4289);
and U4504 (N_4504,N_3830,N_4318);
or U4505 (N_4505,N_4412,N_4092);
xnor U4506 (N_4506,N_4376,N_4275);
nor U4507 (N_4507,N_4199,N_4257);
or U4508 (N_4508,N_4224,N_4000);
nand U4509 (N_4509,N_4117,N_3814);
or U4510 (N_4510,N_4410,N_3998);
nor U4511 (N_4511,N_3771,N_4097);
or U4512 (N_4512,N_4016,N_4398);
and U4513 (N_4513,N_4163,N_4212);
nor U4514 (N_4514,N_4035,N_4047);
xor U4515 (N_4515,N_4351,N_4428);
nand U4516 (N_4516,N_4330,N_4386);
xor U4517 (N_4517,N_3898,N_3990);
nor U4518 (N_4518,N_4265,N_4422);
or U4519 (N_4519,N_3989,N_4134);
nor U4520 (N_4520,N_4286,N_4401);
nor U4521 (N_4521,N_3865,N_4038);
or U4522 (N_4522,N_3957,N_3920);
nor U4523 (N_4523,N_4080,N_3863);
and U4524 (N_4524,N_4417,N_3869);
or U4525 (N_4525,N_4111,N_3803);
or U4526 (N_4526,N_3981,N_4497);
nand U4527 (N_4527,N_3904,N_3820);
and U4528 (N_4528,N_4104,N_4331);
or U4529 (N_4529,N_4392,N_4481);
and U4530 (N_4530,N_4456,N_3905);
or U4531 (N_4531,N_4358,N_4033);
or U4532 (N_4532,N_4053,N_3802);
nor U4533 (N_4533,N_4147,N_3975);
xor U4534 (N_4534,N_4050,N_3809);
or U4535 (N_4535,N_3983,N_3954);
or U4536 (N_4536,N_4446,N_4449);
nor U4537 (N_4537,N_3857,N_4415);
xnor U4538 (N_4538,N_3834,N_3938);
or U4539 (N_4539,N_3811,N_4030);
nand U4540 (N_4540,N_4360,N_4373);
nand U4541 (N_4541,N_4462,N_4332);
xnor U4542 (N_4542,N_3858,N_4442);
and U4543 (N_4543,N_4088,N_3844);
and U4544 (N_4544,N_3915,N_3936);
nand U4545 (N_4545,N_3856,N_4077);
and U4546 (N_4546,N_4178,N_4407);
nor U4547 (N_4547,N_4175,N_4208);
nor U4548 (N_4548,N_4089,N_3781);
nor U4549 (N_4549,N_3808,N_4433);
and U4550 (N_4550,N_3838,N_3779);
nand U4551 (N_4551,N_4206,N_4102);
xnor U4552 (N_4552,N_4362,N_3943);
xnor U4553 (N_4553,N_4315,N_4153);
nor U4554 (N_4554,N_4109,N_3966);
and U4555 (N_4555,N_3890,N_3992);
nand U4556 (N_4556,N_4034,N_4090);
xnor U4557 (N_4557,N_3884,N_3980);
xor U4558 (N_4558,N_4339,N_4486);
xnor U4559 (N_4559,N_4294,N_4059);
nor U4560 (N_4560,N_4384,N_4002);
xnor U4561 (N_4561,N_3796,N_4083);
nand U4562 (N_4562,N_3775,N_4343);
nand U4563 (N_4563,N_4226,N_4353);
nand U4564 (N_4564,N_3942,N_4124);
nor U4565 (N_4565,N_4133,N_4119);
or U4566 (N_4566,N_4247,N_3843);
nor U4567 (N_4567,N_4468,N_4141);
nor U4568 (N_4568,N_4440,N_4411);
and U4569 (N_4569,N_4186,N_4281);
nor U4570 (N_4570,N_4302,N_3845);
nand U4571 (N_4571,N_3793,N_4209);
nor U4572 (N_4572,N_4348,N_4130);
nor U4573 (N_4573,N_4240,N_4015);
xnor U4574 (N_4574,N_4202,N_4017);
nor U4575 (N_4575,N_3790,N_3841);
or U4576 (N_4576,N_4382,N_4120);
nand U4577 (N_4577,N_3977,N_4372);
xnor U4578 (N_4578,N_4094,N_4258);
or U4579 (N_4579,N_4046,N_4181);
xor U4580 (N_4580,N_3787,N_3764);
xnor U4581 (N_4581,N_3991,N_4363);
xnor U4582 (N_4582,N_4167,N_3870);
nor U4583 (N_4583,N_3886,N_4222);
nor U4584 (N_4584,N_4293,N_3799);
or U4585 (N_4585,N_4032,N_3995);
xnor U4586 (N_4586,N_3859,N_4052);
and U4587 (N_4587,N_4327,N_4408);
nor U4588 (N_4588,N_4036,N_4009);
nand U4589 (N_4589,N_4270,N_3924);
nand U4590 (N_4590,N_4314,N_3907);
and U4591 (N_4591,N_4283,N_4100);
xor U4592 (N_4592,N_4326,N_4397);
and U4593 (N_4593,N_3916,N_4498);
or U4594 (N_4594,N_4255,N_4333);
xor U4595 (N_4595,N_4164,N_3911);
or U4596 (N_4596,N_3829,N_3759);
or U4597 (N_4597,N_4288,N_4424);
nor U4598 (N_4598,N_4085,N_4154);
or U4599 (N_4599,N_3988,N_3867);
xnor U4600 (N_4600,N_3947,N_3824);
xor U4601 (N_4601,N_4214,N_4414);
nand U4602 (N_4602,N_4474,N_4023);
xnor U4603 (N_4603,N_4345,N_4253);
or U4604 (N_4604,N_4285,N_4470);
nand U4605 (N_4605,N_4352,N_4118);
nand U4606 (N_4606,N_3922,N_4284);
nor U4607 (N_4607,N_3940,N_4070);
or U4608 (N_4608,N_4403,N_3917);
xor U4609 (N_4609,N_4368,N_4211);
and U4610 (N_4610,N_4146,N_4031);
and U4611 (N_4611,N_4381,N_4241);
xnor U4612 (N_4612,N_4194,N_4019);
nor U4613 (N_4613,N_4168,N_3847);
nand U4614 (N_4614,N_4385,N_4229);
xor U4615 (N_4615,N_3930,N_3819);
nand U4616 (N_4616,N_4074,N_4313);
xor U4617 (N_4617,N_4081,N_3948);
xnor U4618 (N_4618,N_4290,N_3851);
nand U4619 (N_4619,N_3984,N_4320);
nand U4620 (N_4620,N_3773,N_4479);
and U4621 (N_4621,N_3763,N_3906);
or U4622 (N_4622,N_3927,N_3953);
and U4623 (N_4623,N_4370,N_3769);
and U4624 (N_4624,N_4066,N_3950);
nand U4625 (N_4625,N_3831,N_3908);
or U4626 (N_4626,N_4068,N_3864);
and U4627 (N_4627,N_4394,N_4075);
and U4628 (N_4628,N_4048,N_4453);
xnor U4629 (N_4629,N_4344,N_4129);
xor U4630 (N_4630,N_4045,N_4177);
or U4631 (N_4631,N_3903,N_4267);
nand U4632 (N_4632,N_4227,N_3997);
xor U4633 (N_4633,N_3923,N_4135);
nor U4634 (N_4634,N_4391,N_4277);
nor U4635 (N_4635,N_4165,N_4499);
or U4636 (N_4636,N_4496,N_4022);
xnor U4637 (N_4637,N_4242,N_4145);
nor U4638 (N_4638,N_4445,N_3823);
or U4639 (N_4639,N_3879,N_3913);
nor U4640 (N_4640,N_4357,N_3797);
and U4641 (N_4641,N_3946,N_4375);
or U4642 (N_4642,N_4488,N_3918);
nand U4643 (N_4643,N_4413,N_3939);
or U4644 (N_4644,N_4276,N_3952);
nand U4645 (N_4645,N_3852,N_4323);
or U4646 (N_4646,N_4159,N_4107);
nor U4647 (N_4647,N_3817,N_3971);
nand U4648 (N_4648,N_3810,N_4219);
xor U4649 (N_4649,N_4004,N_4179);
nand U4650 (N_4650,N_3816,N_4020);
or U4651 (N_4651,N_4467,N_3806);
or U4652 (N_4652,N_4452,N_3889);
and U4653 (N_4653,N_4426,N_4099);
nor U4654 (N_4654,N_3842,N_4055);
and U4655 (N_4655,N_3887,N_4336);
xor U4656 (N_4656,N_3866,N_3963);
nor U4657 (N_4657,N_4105,N_3926);
or U4658 (N_4658,N_4005,N_3951);
and U4659 (N_4659,N_4093,N_3875);
and U4660 (N_4660,N_4395,N_4063);
or U4661 (N_4661,N_4098,N_4379);
and U4662 (N_4662,N_3780,N_4162);
or U4663 (N_4663,N_3840,N_4245);
and U4664 (N_4664,N_4296,N_4292);
nor U4665 (N_4665,N_3985,N_3969);
nand U4666 (N_4666,N_3825,N_3760);
and U4667 (N_4667,N_4471,N_4328);
nand U4668 (N_4668,N_4136,N_3798);
xor U4669 (N_4669,N_4044,N_3928);
xnor U4670 (N_4670,N_4278,N_3999);
and U4671 (N_4671,N_4246,N_3826);
nor U4672 (N_4672,N_4171,N_3805);
xnor U4673 (N_4673,N_4218,N_4489);
nand U4674 (N_4674,N_4125,N_4239);
nand U4675 (N_4675,N_3935,N_3762);
nor U4676 (N_4676,N_4325,N_4256);
nor U4677 (N_4677,N_3822,N_4155);
or U4678 (N_4678,N_4076,N_3978);
nand U4679 (N_4679,N_4291,N_4233);
and U4680 (N_4680,N_4060,N_4174);
or U4681 (N_4681,N_4176,N_4029);
nor U4682 (N_4682,N_3897,N_3789);
and U4683 (N_4683,N_3751,N_3962);
nand U4684 (N_4684,N_3770,N_4260);
nor U4685 (N_4685,N_4367,N_4039);
nor U4686 (N_4686,N_3986,N_3993);
or U4687 (N_4687,N_4169,N_4065);
nor U4688 (N_4688,N_4185,N_4365);
or U4689 (N_4689,N_3909,N_4454);
and U4690 (N_4690,N_4478,N_4149);
or U4691 (N_4691,N_3833,N_3955);
and U4692 (N_4692,N_4427,N_4429);
or U4693 (N_4693,N_4116,N_3956);
or U4694 (N_4694,N_4364,N_4001);
xor U4695 (N_4695,N_4409,N_4123);
xnor U4696 (N_4696,N_4436,N_3794);
or U4697 (N_4697,N_3827,N_4101);
xnor U4698 (N_4698,N_4091,N_4161);
nor U4699 (N_4699,N_4018,N_4252);
nand U4700 (N_4700,N_4444,N_3848);
nor U4701 (N_4701,N_4355,N_3872);
nor U4702 (N_4702,N_3960,N_3786);
nor U4703 (N_4703,N_4197,N_3895);
nor U4704 (N_4704,N_4354,N_3941);
nand U4705 (N_4705,N_4152,N_3774);
and U4706 (N_4706,N_3944,N_4062);
nand U4707 (N_4707,N_3945,N_4028);
nor U4708 (N_4708,N_3784,N_4347);
xor U4709 (N_4709,N_4151,N_4319);
or U4710 (N_4710,N_4180,N_3788);
nand U4711 (N_4711,N_4191,N_4231);
or U4712 (N_4712,N_3929,N_4447);
nand U4713 (N_4713,N_4073,N_4459);
nand U4714 (N_4714,N_3862,N_3933);
xor U4715 (N_4715,N_4477,N_4448);
and U4716 (N_4716,N_4166,N_4305);
nor U4717 (N_4717,N_4324,N_3934);
xor U4718 (N_4718,N_4232,N_3772);
nor U4719 (N_4719,N_3901,N_4108);
xnor U4720 (N_4720,N_3925,N_3894);
or U4721 (N_4721,N_3880,N_4078);
nor U4722 (N_4722,N_3888,N_4297);
xor U4723 (N_4723,N_4322,N_3987);
nand U4724 (N_4724,N_4484,N_4220);
nor U4725 (N_4725,N_4312,N_3785);
or U4726 (N_4726,N_3767,N_4487);
xor U4727 (N_4727,N_3758,N_4087);
nor U4728 (N_4728,N_3849,N_4306);
or U4729 (N_4729,N_4430,N_4377);
nor U4730 (N_4730,N_3932,N_4303);
xnor U4731 (N_4731,N_4056,N_4172);
nand U4732 (N_4732,N_4140,N_4216);
or U4733 (N_4733,N_4184,N_4485);
and U4734 (N_4734,N_3753,N_4337);
and U4735 (N_4735,N_4201,N_3777);
nor U4736 (N_4736,N_4269,N_3914);
nand U4737 (N_4737,N_4095,N_4432);
or U4738 (N_4738,N_4434,N_4126);
xnor U4739 (N_4739,N_4061,N_4148);
nor U4740 (N_4740,N_4380,N_4158);
or U4741 (N_4741,N_4236,N_3976);
xor U4742 (N_4742,N_4301,N_4210);
xor U4743 (N_4743,N_4193,N_4321);
or U4744 (N_4744,N_4112,N_3937);
and U4745 (N_4745,N_4086,N_4128);
nand U4746 (N_4746,N_4122,N_4213);
nor U4747 (N_4747,N_4304,N_3949);
or U4748 (N_4748,N_3979,N_4404);
nor U4749 (N_4749,N_4494,N_4466);
nand U4750 (N_4750,N_3912,N_3899);
and U4751 (N_4751,N_3967,N_3994);
nor U4752 (N_4752,N_4008,N_4234);
and U4753 (N_4753,N_3959,N_3791);
and U4754 (N_4754,N_4476,N_4188);
nor U4755 (N_4755,N_4225,N_4238);
nor U4756 (N_4756,N_4150,N_4420);
nand U4757 (N_4757,N_4469,N_3973);
xnor U4758 (N_4758,N_4071,N_4113);
nor U4759 (N_4759,N_3972,N_3855);
and U4760 (N_4760,N_3902,N_4402);
or U4761 (N_4761,N_3982,N_4492);
or U4762 (N_4762,N_4472,N_4144);
and U4763 (N_4763,N_4457,N_4121);
nand U4764 (N_4764,N_4183,N_4416);
and U4765 (N_4765,N_4223,N_4244);
and U4766 (N_4766,N_4338,N_3783);
nor U4767 (N_4767,N_4350,N_4040);
or U4768 (N_4768,N_4317,N_4132);
and U4769 (N_4769,N_4106,N_4013);
xnor U4770 (N_4770,N_3804,N_3846);
or U4771 (N_4771,N_4308,N_4007);
xnor U4772 (N_4772,N_4419,N_4139);
nor U4773 (N_4773,N_4263,N_4259);
nand U4774 (N_4774,N_4279,N_4369);
nor U4775 (N_4775,N_4170,N_3996);
xor U4776 (N_4776,N_3815,N_4243);
nand U4777 (N_4777,N_4274,N_4110);
xor U4778 (N_4778,N_4311,N_4437);
nand U4779 (N_4779,N_4042,N_4491);
or U4780 (N_4780,N_3893,N_3800);
nand U4781 (N_4781,N_4156,N_4058);
nand U4782 (N_4782,N_4349,N_4388);
nor U4783 (N_4783,N_4359,N_4435);
xor U4784 (N_4784,N_3853,N_3896);
xor U4785 (N_4785,N_4387,N_4069);
nor U4786 (N_4786,N_3813,N_4431);
nand U4787 (N_4787,N_4406,N_4235);
nor U4788 (N_4788,N_4287,N_4248);
and U4789 (N_4789,N_4182,N_4025);
nand U4790 (N_4790,N_4041,N_4237);
xor U4791 (N_4791,N_4483,N_4014);
or U4792 (N_4792,N_3765,N_4316);
and U4793 (N_4793,N_3881,N_4079);
nor U4794 (N_4794,N_4393,N_4003);
nand U4795 (N_4795,N_3968,N_3836);
or U4796 (N_4796,N_4399,N_4307);
and U4797 (N_4797,N_4441,N_4309);
nor U4798 (N_4798,N_4160,N_4493);
or U4799 (N_4799,N_4037,N_4057);
nand U4800 (N_4800,N_4421,N_4251);
or U4801 (N_4801,N_3910,N_4142);
nor U4802 (N_4802,N_3900,N_4064);
and U4803 (N_4803,N_4187,N_3795);
nor U4804 (N_4804,N_4072,N_3818);
and U4805 (N_4805,N_4299,N_4249);
or U4806 (N_4806,N_4012,N_4371);
or U4807 (N_4807,N_4131,N_3792);
nand U4808 (N_4808,N_4378,N_3768);
xor U4809 (N_4809,N_4204,N_3756);
nor U4810 (N_4810,N_3854,N_3877);
xor U4811 (N_4811,N_3812,N_4400);
or U4812 (N_4812,N_4295,N_4173);
nand U4813 (N_4813,N_3874,N_4340);
xor U4814 (N_4814,N_4011,N_3778);
nor U4815 (N_4815,N_4024,N_4027);
nor U4816 (N_4816,N_4262,N_4458);
nand U4817 (N_4817,N_4361,N_3754);
xor U4818 (N_4818,N_4425,N_4200);
xor U4819 (N_4819,N_4346,N_4298);
xnor U4820 (N_4820,N_4043,N_4084);
or U4821 (N_4821,N_4473,N_4396);
nand U4822 (N_4822,N_4021,N_3750);
xnor U4823 (N_4823,N_4195,N_4221);
and U4824 (N_4824,N_4006,N_4366);
xor U4825 (N_4825,N_3782,N_3885);
and U4826 (N_4826,N_4115,N_3876);
and U4827 (N_4827,N_4230,N_3882);
xor U4828 (N_4828,N_4495,N_4096);
nor U4829 (N_4829,N_4390,N_3871);
nor U4830 (N_4830,N_4051,N_4389);
or U4831 (N_4831,N_4464,N_4439);
xnor U4832 (N_4832,N_4460,N_3873);
xor U4833 (N_4833,N_4438,N_3883);
or U4834 (N_4834,N_4198,N_4423);
and U4835 (N_4835,N_3752,N_4261);
xnor U4836 (N_4836,N_4329,N_4254);
xnor U4837 (N_4837,N_4280,N_4418);
nand U4838 (N_4838,N_4207,N_4143);
nor U4839 (N_4839,N_4273,N_4300);
xor U4840 (N_4840,N_4217,N_4082);
nand U4841 (N_4841,N_4335,N_3965);
nand U4842 (N_4842,N_3931,N_4310);
nand U4843 (N_4843,N_4189,N_4282);
and U4844 (N_4844,N_3974,N_3761);
xor U4845 (N_4845,N_4342,N_4103);
xor U4846 (N_4846,N_3776,N_3878);
and U4847 (N_4847,N_4383,N_4272);
and U4848 (N_4848,N_3757,N_4482);
nor U4849 (N_4849,N_3860,N_3861);
or U4850 (N_4850,N_4264,N_3837);
nand U4851 (N_4851,N_4127,N_4205);
nand U4852 (N_4852,N_3961,N_4455);
xor U4853 (N_4853,N_4271,N_4138);
nor U4854 (N_4854,N_4356,N_4250);
and U4855 (N_4855,N_4266,N_4010);
nor U4856 (N_4856,N_4137,N_4054);
nand U4857 (N_4857,N_3921,N_3958);
or U4858 (N_4858,N_3835,N_4475);
and U4859 (N_4859,N_4334,N_4405);
or U4860 (N_4860,N_4196,N_4451);
or U4861 (N_4861,N_4067,N_3892);
or U4862 (N_4862,N_4490,N_4114);
xnor U4863 (N_4863,N_3755,N_3891);
nor U4864 (N_4864,N_4203,N_3970);
and U4865 (N_4865,N_3801,N_4228);
and U4866 (N_4866,N_4268,N_4190);
xor U4867 (N_4867,N_3832,N_3919);
xor U4868 (N_4868,N_3807,N_3850);
nand U4869 (N_4869,N_4341,N_4461);
nand U4870 (N_4870,N_3839,N_4443);
or U4871 (N_4871,N_3868,N_4463);
and U4872 (N_4872,N_4026,N_4215);
and U4873 (N_4873,N_4465,N_3828);
and U4874 (N_4874,N_4049,N_3964);
xor U4875 (N_4875,N_4023,N_4007);
and U4876 (N_4876,N_4105,N_4301);
or U4877 (N_4877,N_4425,N_4176);
nor U4878 (N_4878,N_4123,N_4055);
xor U4879 (N_4879,N_4176,N_3904);
or U4880 (N_4880,N_3871,N_4327);
xnor U4881 (N_4881,N_4195,N_4013);
nor U4882 (N_4882,N_4280,N_4478);
or U4883 (N_4883,N_3777,N_4131);
nand U4884 (N_4884,N_4397,N_4049);
or U4885 (N_4885,N_4360,N_3808);
xnor U4886 (N_4886,N_4312,N_3898);
and U4887 (N_4887,N_4042,N_4194);
nor U4888 (N_4888,N_3977,N_4428);
xor U4889 (N_4889,N_4487,N_3813);
and U4890 (N_4890,N_4173,N_4298);
xnor U4891 (N_4891,N_4264,N_4260);
and U4892 (N_4892,N_3773,N_3990);
or U4893 (N_4893,N_3873,N_3763);
xor U4894 (N_4894,N_3880,N_4278);
or U4895 (N_4895,N_3755,N_4221);
and U4896 (N_4896,N_4162,N_3954);
nand U4897 (N_4897,N_4135,N_4336);
or U4898 (N_4898,N_4308,N_4252);
or U4899 (N_4899,N_4267,N_4095);
nand U4900 (N_4900,N_4334,N_4225);
xor U4901 (N_4901,N_3851,N_4104);
xor U4902 (N_4902,N_3851,N_4251);
or U4903 (N_4903,N_4025,N_3935);
and U4904 (N_4904,N_4411,N_4375);
or U4905 (N_4905,N_3755,N_3805);
nor U4906 (N_4906,N_4198,N_4230);
and U4907 (N_4907,N_3945,N_3842);
nand U4908 (N_4908,N_3855,N_4236);
or U4909 (N_4909,N_3863,N_4104);
nand U4910 (N_4910,N_4346,N_3868);
and U4911 (N_4911,N_4347,N_4293);
nor U4912 (N_4912,N_3930,N_3807);
and U4913 (N_4913,N_4158,N_4335);
nor U4914 (N_4914,N_4115,N_4246);
or U4915 (N_4915,N_4466,N_3985);
xor U4916 (N_4916,N_4448,N_4270);
and U4917 (N_4917,N_4497,N_4174);
and U4918 (N_4918,N_3865,N_4113);
nor U4919 (N_4919,N_4160,N_4045);
nor U4920 (N_4920,N_4331,N_4356);
and U4921 (N_4921,N_3774,N_4379);
nand U4922 (N_4922,N_3944,N_3930);
and U4923 (N_4923,N_4424,N_4334);
xnor U4924 (N_4924,N_4338,N_4459);
nor U4925 (N_4925,N_4490,N_3927);
or U4926 (N_4926,N_4327,N_3965);
nand U4927 (N_4927,N_4078,N_3902);
or U4928 (N_4928,N_4051,N_4497);
xnor U4929 (N_4929,N_3961,N_3796);
or U4930 (N_4930,N_4494,N_4003);
and U4931 (N_4931,N_4166,N_4365);
nand U4932 (N_4932,N_4441,N_4221);
or U4933 (N_4933,N_3766,N_4466);
nor U4934 (N_4934,N_3999,N_3752);
or U4935 (N_4935,N_4451,N_3979);
nor U4936 (N_4936,N_4450,N_3866);
xnor U4937 (N_4937,N_3920,N_3787);
or U4938 (N_4938,N_3809,N_3951);
or U4939 (N_4939,N_3770,N_4299);
nor U4940 (N_4940,N_4396,N_3818);
and U4941 (N_4941,N_4200,N_4432);
nand U4942 (N_4942,N_4284,N_4476);
nand U4943 (N_4943,N_4276,N_3942);
and U4944 (N_4944,N_3853,N_4271);
nor U4945 (N_4945,N_3831,N_4020);
nand U4946 (N_4946,N_3851,N_3890);
nor U4947 (N_4947,N_4216,N_3783);
xnor U4948 (N_4948,N_3814,N_4076);
and U4949 (N_4949,N_3933,N_4340);
and U4950 (N_4950,N_4480,N_4474);
nor U4951 (N_4951,N_4367,N_4471);
xor U4952 (N_4952,N_3976,N_3827);
or U4953 (N_4953,N_4245,N_4272);
xnor U4954 (N_4954,N_3829,N_3768);
or U4955 (N_4955,N_3864,N_4213);
nand U4956 (N_4956,N_4124,N_3751);
and U4957 (N_4957,N_4290,N_4088);
nor U4958 (N_4958,N_4102,N_4129);
or U4959 (N_4959,N_4132,N_4316);
nand U4960 (N_4960,N_4089,N_3838);
nand U4961 (N_4961,N_3942,N_3958);
or U4962 (N_4962,N_4312,N_4359);
nand U4963 (N_4963,N_4037,N_3760);
nand U4964 (N_4964,N_4113,N_4036);
nand U4965 (N_4965,N_4113,N_4019);
xor U4966 (N_4966,N_4015,N_3858);
xnor U4967 (N_4967,N_4194,N_3916);
nor U4968 (N_4968,N_3766,N_4387);
nor U4969 (N_4969,N_3798,N_4289);
nor U4970 (N_4970,N_4256,N_3907);
xnor U4971 (N_4971,N_3946,N_3893);
xor U4972 (N_4972,N_4462,N_4108);
xor U4973 (N_4973,N_3876,N_3840);
nand U4974 (N_4974,N_4378,N_4422);
nor U4975 (N_4975,N_4037,N_3785);
and U4976 (N_4976,N_3947,N_4483);
or U4977 (N_4977,N_4125,N_4364);
nor U4978 (N_4978,N_4363,N_4185);
xor U4979 (N_4979,N_4179,N_4326);
nand U4980 (N_4980,N_4474,N_3856);
xor U4981 (N_4981,N_4390,N_3814);
nand U4982 (N_4982,N_4173,N_4347);
and U4983 (N_4983,N_3781,N_4450);
nor U4984 (N_4984,N_4293,N_3936);
or U4985 (N_4985,N_4038,N_3959);
and U4986 (N_4986,N_4212,N_3965);
or U4987 (N_4987,N_3888,N_4325);
xnor U4988 (N_4988,N_4294,N_3839);
nor U4989 (N_4989,N_3779,N_4040);
nand U4990 (N_4990,N_4111,N_4116);
or U4991 (N_4991,N_3815,N_4033);
nor U4992 (N_4992,N_4154,N_4155);
xnor U4993 (N_4993,N_4479,N_4384);
or U4994 (N_4994,N_4470,N_4388);
and U4995 (N_4995,N_3779,N_4073);
nor U4996 (N_4996,N_3945,N_4059);
and U4997 (N_4997,N_3900,N_4387);
xor U4998 (N_4998,N_4233,N_4184);
xor U4999 (N_4999,N_4488,N_4322);
and U5000 (N_5000,N_3787,N_4085);
nand U5001 (N_5001,N_4078,N_3963);
xnor U5002 (N_5002,N_3885,N_3973);
and U5003 (N_5003,N_3789,N_3975);
xnor U5004 (N_5004,N_4056,N_4352);
xnor U5005 (N_5005,N_3943,N_4209);
and U5006 (N_5006,N_4434,N_4295);
and U5007 (N_5007,N_3899,N_4155);
nor U5008 (N_5008,N_3962,N_3759);
or U5009 (N_5009,N_4140,N_4226);
and U5010 (N_5010,N_4121,N_3783);
xor U5011 (N_5011,N_4080,N_3955);
xor U5012 (N_5012,N_3851,N_4179);
nand U5013 (N_5013,N_4315,N_4106);
xnor U5014 (N_5014,N_3882,N_4031);
xor U5015 (N_5015,N_3955,N_4240);
or U5016 (N_5016,N_4373,N_4318);
nand U5017 (N_5017,N_4345,N_4055);
nor U5018 (N_5018,N_3955,N_3750);
and U5019 (N_5019,N_3804,N_3781);
or U5020 (N_5020,N_4280,N_4446);
xor U5021 (N_5021,N_4031,N_4272);
or U5022 (N_5022,N_4193,N_3970);
nand U5023 (N_5023,N_4085,N_4052);
nand U5024 (N_5024,N_4212,N_3949);
and U5025 (N_5025,N_4342,N_4256);
or U5026 (N_5026,N_3871,N_4049);
and U5027 (N_5027,N_3966,N_3886);
or U5028 (N_5028,N_3779,N_3896);
nand U5029 (N_5029,N_4108,N_3982);
xnor U5030 (N_5030,N_4417,N_4395);
nor U5031 (N_5031,N_4039,N_3875);
nor U5032 (N_5032,N_3826,N_4461);
and U5033 (N_5033,N_3836,N_4270);
nand U5034 (N_5034,N_3888,N_3853);
nand U5035 (N_5035,N_4388,N_4357);
xor U5036 (N_5036,N_4205,N_3932);
xor U5037 (N_5037,N_3764,N_4298);
or U5038 (N_5038,N_4139,N_3834);
and U5039 (N_5039,N_4055,N_4426);
nand U5040 (N_5040,N_4038,N_4168);
xor U5041 (N_5041,N_4270,N_4384);
nor U5042 (N_5042,N_4290,N_3924);
and U5043 (N_5043,N_3915,N_3856);
or U5044 (N_5044,N_3976,N_3983);
nor U5045 (N_5045,N_3786,N_3952);
nand U5046 (N_5046,N_4201,N_4202);
nor U5047 (N_5047,N_3876,N_4048);
nor U5048 (N_5048,N_3774,N_4326);
and U5049 (N_5049,N_4198,N_3907);
or U5050 (N_5050,N_4299,N_4149);
nand U5051 (N_5051,N_4489,N_4328);
nor U5052 (N_5052,N_4314,N_4253);
nor U5053 (N_5053,N_3876,N_3918);
xnor U5054 (N_5054,N_3799,N_4194);
and U5055 (N_5055,N_4078,N_4145);
xnor U5056 (N_5056,N_4036,N_4337);
or U5057 (N_5057,N_4240,N_3917);
and U5058 (N_5058,N_4495,N_3971);
and U5059 (N_5059,N_3763,N_4293);
nor U5060 (N_5060,N_4116,N_3961);
or U5061 (N_5061,N_4360,N_4193);
nand U5062 (N_5062,N_4365,N_4285);
xor U5063 (N_5063,N_4075,N_4047);
xnor U5064 (N_5064,N_4013,N_4018);
and U5065 (N_5065,N_4456,N_4330);
or U5066 (N_5066,N_4441,N_4292);
nand U5067 (N_5067,N_4092,N_3942);
nor U5068 (N_5068,N_3878,N_4340);
nand U5069 (N_5069,N_3919,N_3794);
or U5070 (N_5070,N_4229,N_3894);
or U5071 (N_5071,N_3779,N_4423);
xor U5072 (N_5072,N_3892,N_3928);
and U5073 (N_5073,N_3827,N_4128);
nor U5074 (N_5074,N_4086,N_4020);
nand U5075 (N_5075,N_4444,N_3997);
or U5076 (N_5076,N_4235,N_4422);
or U5077 (N_5077,N_3780,N_4109);
and U5078 (N_5078,N_4454,N_3948);
xnor U5079 (N_5079,N_3948,N_4463);
nor U5080 (N_5080,N_4366,N_4034);
xor U5081 (N_5081,N_3787,N_4436);
or U5082 (N_5082,N_4034,N_4445);
or U5083 (N_5083,N_4353,N_4428);
or U5084 (N_5084,N_4085,N_4211);
nand U5085 (N_5085,N_3972,N_4092);
and U5086 (N_5086,N_4463,N_4369);
nor U5087 (N_5087,N_4240,N_4373);
nor U5088 (N_5088,N_3767,N_3804);
xnor U5089 (N_5089,N_3918,N_4492);
nand U5090 (N_5090,N_3962,N_3830);
xor U5091 (N_5091,N_4133,N_3773);
nand U5092 (N_5092,N_4112,N_3841);
xor U5093 (N_5093,N_4188,N_4267);
nor U5094 (N_5094,N_4151,N_4431);
xor U5095 (N_5095,N_4263,N_4311);
nor U5096 (N_5096,N_4053,N_3925);
or U5097 (N_5097,N_4109,N_4427);
and U5098 (N_5098,N_4288,N_4041);
and U5099 (N_5099,N_4018,N_4048);
nand U5100 (N_5100,N_3861,N_4419);
xor U5101 (N_5101,N_3804,N_4143);
and U5102 (N_5102,N_4093,N_4098);
nor U5103 (N_5103,N_4061,N_4097);
or U5104 (N_5104,N_4103,N_4434);
nor U5105 (N_5105,N_4088,N_4387);
xor U5106 (N_5106,N_4224,N_4297);
or U5107 (N_5107,N_4197,N_3953);
or U5108 (N_5108,N_4426,N_4128);
nor U5109 (N_5109,N_4099,N_4023);
xnor U5110 (N_5110,N_4226,N_4162);
nor U5111 (N_5111,N_3879,N_4282);
nor U5112 (N_5112,N_4088,N_4202);
and U5113 (N_5113,N_4157,N_4294);
or U5114 (N_5114,N_4461,N_4187);
xnor U5115 (N_5115,N_4072,N_4031);
nand U5116 (N_5116,N_4358,N_3759);
and U5117 (N_5117,N_4491,N_4016);
and U5118 (N_5118,N_4438,N_3904);
nand U5119 (N_5119,N_4291,N_4168);
xnor U5120 (N_5120,N_4409,N_3786);
nand U5121 (N_5121,N_4345,N_4341);
xnor U5122 (N_5122,N_4107,N_4291);
and U5123 (N_5123,N_4491,N_4372);
xnor U5124 (N_5124,N_3955,N_4053);
xnor U5125 (N_5125,N_4298,N_4242);
nand U5126 (N_5126,N_3999,N_4330);
nor U5127 (N_5127,N_3867,N_3968);
and U5128 (N_5128,N_4236,N_3800);
or U5129 (N_5129,N_3867,N_4277);
nand U5130 (N_5130,N_4376,N_4217);
xnor U5131 (N_5131,N_4320,N_4267);
nand U5132 (N_5132,N_4485,N_4261);
xor U5133 (N_5133,N_4489,N_4406);
nor U5134 (N_5134,N_4486,N_4415);
or U5135 (N_5135,N_4012,N_4388);
or U5136 (N_5136,N_4273,N_4191);
or U5137 (N_5137,N_4381,N_3899);
xnor U5138 (N_5138,N_4424,N_3983);
or U5139 (N_5139,N_4449,N_4257);
xnor U5140 (N_5140,N_4007,N_3773);
nor U5141 (N_5141,N_4242,N_3971);
xor U5142 (N_5142,N_4150,N_4470);
and U5143 (N_5143,N_4362,N_4056);
and U5144 (N_5144,N_4178,N_4317);
or U5145 (N_5145,N_4457,N_3946);
nand U5146 (N_5146,N_4118,N_3960);
and U5147 (N_5147,N_4290,N_3872);
or U5148 (N_5148,N_3934,N_4288);
or U5149 (N_5149,N_4192,N_4251);
xnor U5150 (N_5150,N_4116,N_4002);
nand U5151 (N_5151,N_4037,N_4047);
or U5152 (N_5152,N_4355,N_3902);
nand U5153 (N_5153,N_4164,N_4493);
nand U5154 (N_5154,N_4169,N_4428);
nor U5155 (N_5155,N_3935,N_4483);
and U5156 (N_5156,N_4293,N_4486);
nor U5157 (N_5157,N_3841,N_4011);
and U5158 (N_5158,N_4181,N_3903);
nor U5159 (N_5159,N_3883,N_4482);
nor U5160 (N_5160,N_4291,N_4436);
nand U5161 (N_5161,N_4213,N_3914);
nor U5162 (N_5162,N_4349,N_4266);
and U5163 (N_5163,N_4201,N_4161);
xor U5164 (N_5164,N_4116,N_3892);
nand U5165 (N_5165,N_4091,N_3960);
nand U5166 (N_5166,N_4256,N_4182);
nand U5167 (N_5167,N_4369,N_3963);
and U5168 (N_5168,N_4135,N_4485);
xnor U5169 (N_5169,N_4106,N_4362);
or U5170 (N_5170,N_4164,N_3806);
and U5171 (N_5171,N_4308,N_4110);
nor U5172 (N_5172,N_3913,N_4311);
or U5173 (N_5173,N_3888,N_4024);
nand U5174 (N_5174,N_4209,N_4208);
xnor U5175 (N_5175,N_3778,N_4304);
nand U5176 (N_5176,N_3886,N_4176);
nand U5177 (N_5177,N_4461,N_4039);
nor U5178 (N_5178,N_4196,N_4031);
xor U5179 (N_5179,N_4285,N_4098);
nand U5180 (N_5180,N_3815,N_4022);
nor U5181 (N_5181,N_3975,N_3831);
and U5182 (N_5182,N_3949,N_4392);
xor U5183 (N_5183,N_4127,N_4238);
nor U5184 (N_5184,N_3812,N_3789);
nor U5185 (N_5185,N_3885,N_4490);
and U5186 (N_5186,N_4234,N_4343);
and U5187 (N_5187,N_3979,N_3905);
nand U5188 (N_5188,N_4492,N_3939);
or U5189 (N_5189,N_4482,N_4120);
and U5190 (N_5190,N_4120,N_4421);
or U5191 (N_5191,N_4383,N_3940);
or U5192 (N_5192,N_4349,N_3773);
or U5193 (N_5193,N_3764,N_4291);
or U5194 (N_5194,N_4198,N_3838);
nor U5195 (N_5195,N_4490,N_3877);
nand U5196 (N_5196,N_3798,N_4070);
xnor U5197 (N_5197,N_3752,N_3933);
xnor U5198 (N_5198,N_4096,N_4432);
nor U5199 (N_5199,N_4404,N_3853);
nor U5200 (N_5200,N_4354,N_4245);
and U5201 (N_5201,N_3815,N_4269);
nand U5202 (N_5202,N_3880,N_4082);
or U5203 (N_5203,N_3924,N_4170);
xor U5204 (N_5204,N_4368,N_3951);
and U5205 (N_5205,N_4355,N_4489);
nand U5206 (N_5206,N_4325,N_3931);
nand U5207 (N_5207,N_4147,N_4274);
nor U5208 (N_5208,N_3892,N_3900);
xor U5209 (N_5209,N_4179,N_4368);
and U5210 (N_5210,N_4016,N_4062);
nor U5211 (N_5211,N_4122,N_4445);
or U5212 (N_5212,N_4453,N_3804);
and U5213 (N_5213,N_4415,N_3876);
and U5214 (N_5214,N_3854,N_4311);
and U5215 (N_5215,N_4242,N_3942);
xor U5216 (N_5216,N_4210,N_3763);
nand U5217 (N_5217,N_3880,N_4430);
nand U5218 (N_5218,N_3986,N_4140);
nand U5219 (N_5219,N_4346,N_4102);
nor U5220 (N_5220,N_4387,N_3909);
nand U5221 (N_5221,N_4319,N_4362);
or U5222 (N_5222,N_4069,N_3920);
nor U5223 (N_5223,N_4331,N_4115);
xnor U5224 (N_5224,N_4047,N_3910);
or U5225 (N_5225,N_4008,N_3843);
xor U5226 (N_5226,N_4247,N_4049);
and U5227 (N_5227,N_4486,N_4268);
nor U5228 (N_5228,N_4423,N_4228);
nand U5229 (N_5229,N_3921,N_4037);
or U5230 (N_5230,N_4438,N_4240);
and U5231 (N_5231,N_3896,N_4179);
or U5232 (N_5232,N_4101,N_4205);
or U5233 (N_5233,N_3935,N_4038);
or U5234 (N_5234,N_4435,N_4457);
or U5235 (N_5235,N_4002,N_4382);
nand U5236 (N_5236,N_4331,N_4296);
or U5237 (N_5237,N_3919,N_3770);
xor U5238 (N_5238,N_3848,N_3844);
nor U5239 (N_5239,N_4213,N_3910);
and U5240 (N_5240,N_3810,N_3836);
xnor U5241 (N_5241,N_3969,N_3763);
nand U5242 (N_5242,N_4171,N_4094);
nand U5243 (N_5243,N_4408,N_3879);
or U5244 (N_5244,N_3836,N_4221);
and U5245 (N_5245,N_4213,N_4206);
nor U5246 (N_5246,N_4139,N_3752);
nor U5247 (N_5247,N_3756,N_4461);
nand U5248 (N_5248,N_4112,N_4012);
nand U5249 (N_5249,N_3813,N_4355);
xor U5250 (N_5250,N_4800,N_4945);
nand U5251 (N_5251,N_5007,N_4781);
or U5252 (N_5252,N_4757,N_5067);
and U5253 (N_5253,N_5231,N_4891);
xor U5254 (N_5254,N_4782,N_4563);
nor U5255 (N_5255,N_4566,N_4558);
xor U5256 (N_5256,N_4934,N_4517);
xnor U5257 (N_5257,N_5013,N_5004);
nor U5258 (N_5258,N_4737,N_5235);
nand U5259 (N_5259,N_4553,N_4805);
or U5260 (N_5260,N_4920,N_4613);
or U5261 (N_5261,N_4612,N_5200);
nand U5262 (N_5262,N_4738,N_5017);
or U5263 (N_5263,N_5003,N_5071);
xnor U5264 (N_5264,N_4617,N_4573);
nor U5265 (N_5265,N_5210,N_5236);
nand U5266 (N_5266,N_4971,N_4864);
and U5267 (N_5267,N_4731,N_5065);
nor U5268 (N_5268,N_4895,N_4967);
and U5269 (N_5269,N_4594,N_5153);
or U5270 (N_5270,N_4537,N_4548);
or U5271 (N_5271,N_5196,N_5179);
and U5272 (N_5272,N_4858,N_4640);
nor U5273 (N_5273,N_5193,N_4669);
or U5274 (N_5274,N_5203,N_4774);
nand U5275 (N_5275,N_5000,N_4515);
and U5276 (N_5276,N_4648,N_4838);
or U5277 (N_5277,N_4646,N_4939);
xor U5278 (N_5278,N_5039,N_4751);
nor U5279 (N_5279,N_4922,N_5151);
xnor U5280 (N_5280,N_5111,N_4629);
and U5281 (N_5281,N_4596,N_4765);
or U5282 (N_5282,N_4961,N_5030);
xnor U5283 (N_5283,N_5227,N_5079);
nor U5284 (N_5284,N_5016,N_5057);
and U5285 (N_5285,N_4835,N_4874);
xnor U5286 (N_5286,N_5248,N_4704);
or U5287 (N_5287,N_4758,N_5206);
and U5288 (N_5288,N_4813,N_4626);
nand U5289 (N_5289,N_5220,N_4501);
or U5290 (N_5290,N_4621,N_4723);
or U5291 (N_5291,N_4993,N_4830);
and U5292 (N_5292,N_4930,N_5012);
and U5293 (N_5293,N_4590,N_4820);
or U5294 (N_5294,N_4968,N_4959);
nor U5295 (N_5295,N_5122,N_5062);
or U5296 (N_5296,N_4714,N_5087);
nand U5297 (N_5297,N_5105,N_4915);
nand U5298 (N_5298,N_4510,N_4887);
nor U5299 (N_5299,N_5008,N_4883);
xor U5300 (N_5300,N_5136,N_4983);
and U5301 (N_5301,N_5116,N_4581);
nand U5302 (N_5302,N_4685,N_5126);
xnor U5303 (N_5303,N_4651,N_4734);
and U5304 (N_5304,N_4671,N_4933);
and U5305 (N_5305,N_5212,N_4745);
xnor U5306 (N_5306,N_5186,N_5046);
or U5307 (N_5307,N_4914,N_5225);
nand U5308 (N_5308,N_4787,N_4546);
xor U5309 (N_5309,N_5246,N_4942);
or U5310 (N_5310,N_4851,N_5052);
xor U5311 (N_5311,N_4703,N_4588);
or U5312 (N_5312,N_4618,N_4882);
nor U5313 (N_5313,N_5115,N_4752);
nand U5314 (N_5314,N_4688,N_5041);
xor U5315 (N_5315,N_5102,N_4762);
nor U5316 (N_5316,N_5029,N_4916);
and U5317 (N_5317,N_4861,N_5158);
xnor U5318 (N_5318,N_4520,N_4698);
and U5319 (N_5319,N_4866,N_5174);
xnor U5320 (N_5320,N_4700,N_4630);
xor U5321 (N_5321,N_5019,N_5106);
xor U5322 (N_5322,N_5051,N_4913);
xor U5323 (N_5323,N_4662,N_4844);
xnor U5324 (N_5324,N_4921,N_4592);
and U5325 (N_5325,N_5036,N_4832);
nand U5326 (N_5326,N_4719,N_4972);
nor U5327 (N_5327,N_4994,N_4759);
xnor U5328 (N_5328,N_5092,N_5168);
or U5329 (N_5329,N_5217,N_5124);
nor U5330 (N_5330,N_4725,N_5077);
or U5331 (N_5331,N_4801,N_5159);
nand U5332 (N_5332,N_4579,N_5219);
and U5333 (N_5333,N_5025,N_4504);
xor U5334 (N_5334,N_5035,N_4753);
nand U5335 (N_5335,N_4599,N_4679);
nor U5336 (N_5336,N_5044,N_5090);
nor U5337 (N_5337,N_4608,N_4947);
nand U5338 (N_5338,N_4733,N_4954);
or U5339 (N_5339,N_4681,N_4855);
nor U5340 (N_5340,N_5024,N_4761);
or U5341 (N_5341,N_4978,N_4935);
nor U5342 (N_5342,N_4710,N_5249);
nand U5343 (N_5343,N_5050,N_4513);
and U5344 (N_5344,N_4760,N_4996);
xnor U5345 (N_5345,N_4890,N_4728);
nor U5346 (N_5346,N_4684,N_5089);
xnor U5347 (N_5347,N_4951,N_4777);
and U5348 (N_5348,N_4969,N_4525);
nor U5349 (N_5349,N_4840,N_4899);
xor U5350 (N_5350,N_4503,N_4834);
nand U5351 (N_5351,N_5107,N_4905);
and U5352 (N_5352,N_5084,N_5207);
xnor U5353 (N_5353,N_4817,N_4673);
nor U5354 (N_5354,N_5209,N_5202);
nand U5355 (N_5355,N_5185,N_5183);
xnor U5356 (N_5356,N_4987,N_4902);
nand U5357 (N_5357,N_5023,N_5245);
and U5358 (N_5358,N_4661,N_4876);
and U5359 (N_5359,N_4824,N_4664);
nand U5360 (N_5360,N_4849,N_4683);
nor U5361 (N_5361,N_4543,N_4816);
xnor U5362 (N_5362,N_5088,N_4929);
nor U5363 (N_5363,N_5164,N_4649);
nor U5364 (N_5364,N_4518,N_5154);
nand U5365 (N_5365,N_4955,N_4607);
xor U5366 (N_5366,N_5061,N_5130);
or U5367 (N_5367,N_4539,N_4638);
nand U5368 (N_5368,N_4790,N_5074);
xor U5369 (N_5369,N_4549,N_4524);
and U5370 (N_5370,N_4709,N_4586);
and U5371 (N_5371,N_5011,N_5038);
nor U5372 (N_5372,N_5201,N_4949);
nor U5373 (N_5373,N_4544,N_4878);
nor U5374 (N_5374,N_4692,N_5161);
or U5375 (N_5375,N_4516,N_4880);
and U5376 (N_5376,N_5001,N_5134);
xor U5377 (N_5377,N_4602,N_5045);
nor U5378 (N_5378,N_4953,N_4944);
nand U5379 (N_5379,N_5173,N_4636);
nand U5380 (N_5380,N_4846,N_5028);
and U5381 (N_5381,N_5226,N_5175);
nor U5382 (N_5382,N_4742,N_5195);
nand U5383 (N_5383,N_5109,N_4940);
or U5384 (N_5384,N_5123,N_4655);
and U5385 (N_5385,N_4889,N_5176);
xor U5386 (N_5386,N_4672,N_5172);
xnor U5387 (N_5387,N_5223,N_4932);
or U5388 (N_5388,N_5241,N_5101);
nand U5389 (N_5389,N_5110,N_5103);
nand U5390 (N_5390,N_4918,N_4614);
xnor U5391 (N_5391,N_5027,N_5006);
nand U5392 (N_5392,N_4687,N_5069);
and U5393 (N_5393,N_4829,N_5234);
xor U5394 (N_5394,N_4561,N_4875);
and U5395 (N_5395,N_5190,N_5137);
and U5396 (N_5396,N_4810,N_4606);
xor U5397 (N_5397,N_4901,N_4507);
and U5398 (N_5398,N_4711,N_4619);
and U5399 (N_5399,N_4767,N_4966);
xor U5400 (N_5400,N_4772,N_4724);
nor U5401 (N_5401,N_4552,N_4917);
nor U5402 (N_5402,N_4925,N_5140);
and U5403 (N_5403,N_4946,N_4666);
nor U5404 (N_5404,N_5118,N_4668);
xor U5405 (N_5405,N_4744,N_4826);
nor U5406 (N_5406,N_4756,N_5177);
nor U5407 (N_5407,N_5198,N_4506);
and U5408 (N_5408,N_4706,N_4909);
nand U5409 (N_5409,N_4770,N_4884);
nor U5410 (N_5410,N_4936,N_4535);
xor U5411 (N_5411,N_5139,N_5213);
and U5412 (N_5412,N_4522,N_4989);
xnor U5413 (N_5413,N_5064,N_5078);
or U5414 (N_5414,N_4604,N_5184);
and U5415 (N_5415,N_4642,N_4786);
nand U5416 (N_5416,N_4697,N_5053);
or U5417 (N_5417,N_4641,N_4582);
nand U5418 (N_5418,N_4847,N_4521);
or U5419 (N_5419,N_4637,N_4635);
nor U5420 (N_5420,N_4567,N_4571);
and U5421 (N_5421,N_4659,N_5211);
xor U5422 (N_5422,N_5020,N_4812);
nand U5423 (N_5423,N_4593,N_5002);
and U5424 (N_5424,N_4721,N_4540);
xor U5425 (N_5425,N_4665,N_4990);
nand U5426 (N_5426,N_4647,N_5034);
xor U5427 (N_5427,N_4514,N_4633);
nand U5428 (N_5428,N_4928,N_4803);
and U5429 (N_5429,N_5119,N_4695);
nand U5430 (N_5430,N_4746,N_4792);
nand U5431 (N_5431,N_4974,N_4938);
nor U5432 (N_5432,N_5143,N_4825);
nand U5433 (N_5433,N_5049,N_4699);
xnor U5434 (N_5434,N_4653,N_4892);
nor U5435 (N_5435,N_4644,N_5117);
nor U5436 (N_5436,N_5129,N_4982);
and U5437 (N_5437,N_4857,N_4739);
nor U5438 (N_5438,N_4986,N_4715);
nor U5439 (N_5439,N_4568,N_4625);
nor U5440 (N_5440,N_4559,N_4799);
and U5441 (N_5441,N_4754,N_5128);
or U5442 (N_5442,N_4984,N_5162);
nand U5443 (N_5443,N_4574,N_4554);
and U5444 (N_5444,N_5026,N_4511);
and U5445 (N_5445,N_5189,N_4536);
xnor U5446 (N_5446,N_4776,N_5205);
nor U5447 (N_5447,N_4798,N_4763);
nand U5448 (N_5448,N_5135,N_4735);
nor U5449 (N_5449,N_4631,N_5085);
or U5450 (N_5450,N_4707,N_5108);
xnor U5451 (N_5451,N_4839,N_5171);
nor U5452 (N_5452,N_4736,N_4660);
nand U5453 (N_5453,N_4557,N_4815);
nand U5454 (N_5454,N_4718,N_5066);
and U5455 (N_5455,N_4624,N_5099);
or U5456 (N_5456,N_4999,N_4980);
nor U5457 (N_5457,N_5033,N_4863);
xor U5458 (N_5458,N_4551,N_5147);
nor U5459 (N_5459,N_4712,N_5091);
nor U5460 (N_5460,N_4676,N_4585);
nor U5461 (N_5461,N_4663,N_5040);
nand U5462 (N_5462,N_4868,N_5178);
nand U5463 (N_5463,N_4750,N_4981);
or U5464 (N_5464,N_4927,N_5145);
xor U5465 (N_5465,N_4527,N_5022);
and U5466 (N_5466,N_5197,N_4900);
and U5467 (N_5467,N_4879,N_4937);
xor U5468 (N_5468,N_4598,N_4605);
or U5469 (N_5469,N_4717,N_4541);
nor U5470 (N_5470,N_4912,N_5192);
or U5471 (N_5471,N_5100,N_4730);
xnor U5472 (N_5472,N_5215,N_4747);
or U5473 (N_5473,N_4941,N_4806);
xor U5474 (N_5474,N_5054,N_4870);
and U5475 (N_5475,N_4542,N_4862);
or U5476 (N_5476,N_4797,N_5042);
nor U5477 (N_5477,N_5242,N_4841);
and U5478 (N_5478,N_4965,N_5113);
or U5479 (N_5479,N_5005,N_5208);
nand U5480 (N_5480,N_4906,N_4804);
xor U5481 (N_5481,N_4526,N_5237);
or U5482 (N_5482,N_4500,N_4578);
xnor U5483 (N_5483,N_4995,N_4822);
and U5484 (N_5484,N_4611,N_5238);
or U5485 (N_5485,N_4562,N_4924);
nor U5486 (N_5486,N_4809,N_4992);
xnor U5487 (N_5487,N_4645,N_5180);
and U5488 (N_5488,N_5056,N_4694);
or U5489 (N_5489,N_5156,N_4819);
nand U5490 (N_5490,N_4689,N_4764);
nor U5491 (N_5491,N_4885,N_4779);
and U5492 (N_5492,N_4894,N_4749);
xor U5493 (N_5493,N_4748,N_4977);
or U5494 (N_5494,N_5010,N_5127);
and U5495 (N_5495,N_4869,N_4702);
or U5496 (N_5496,N_5094,N_4818);
nor U5497 (N_5497,N_5247,N_5121);
or U5498 (N_5498,N_4888,N_4877);
xnor U5499 (N_5499,N_4852,N_4505);
or U5500 (N_5500,N_5093,N_4896);
and U5501 (N_5501,N_4991,N_4956);
nand U5502 (N_5502,N_4538,N_4519);
nand U5503 (N_5503,N_5232,N_5239);
and U5504 (N_5504,N_5167,N_4973);
xnor U5505 (N_5505,N_4677,N_4555);
nand U5506 (N_5506,N_5229,N_4976);
nor U5507 (N_5507,N_4584,N_4623);
or U5508 (N_5508,N_4794,N_5095);
or U5509 (N_5509,N_4886,N_4670);
nor U5510 (N_5510,N_4589,N_4910);
nand U5511 (N_5511,N_4893,N_5204);
or U5512 (N_5512,N_5080,N_4727);
nand U5513 (N_5513,N_5015,N_5097);
and U5514 (N_5514,N_4867,N_5014);
and U5515 (N_5515,N_4997,N_4778);
xor U5516 (N_5516,N_4674,N_4690);
or U5517 (N_5517,N_4678,N_4530);
and U5518 (N_5518,N_4656,N_5216);
xor U5519 (N_5519,N_4620,N_4523);
nor U5520 (N_5520,N_5141,N_4768);
nand U5521 (N_5521,N_4881,N_4771);
nand U5522 (N_5522,N_4854,N_4907);
or U5523 (N_5523,N_4696,N_5160);
nor U5524 (N_5524,N_5222,N_4837);
nand U5525 (N_5525,N_5075,N_4964);
xnor U5526 (N_5526,N_4686,N_4823);
nor U5527 (N_5527,N_5047,N_4872);
nor U5528 (N_5528,N_5221,N_5138);
xor U5529 (N_5529,N_4873,N_4693);
and U5530 (N_5530,N_4722,N_4897);
nand U5531 (N_5531,N_5073,N_5240);
nor U5532 (N_5532,N_4565,N_5181);
nor U5533 (N_5533,N_4821,N_4743);
xor U5534 (N_5534,N_4975,N_4831);
or U5535 (N_5535,N_4962,N_4708);
nand U5536 (N_5536,N_5170,N_4658);
xnor U5537 (N_5537,N_5112,N_4691);
or U5538 (N_5538,N_4572,N_4643);
or U5539 (N_5539,N_5132,N_5021);
nand U5540 (N_5540,N_4931,N_4560);
and U5541 (N_5541,N_4836,N_4843);
xor U5542 (N_5542,N_5037,N_4948);
and U5543 (N_5543,N_5182,N_4769);
nand U5544 (N_5544,N_5230,N_4904);
xnor U5545 (N_5545,N_4963,N_4632);
or U5546 (N_5546,N_4908,N_5125);
and U5547 (N_5547,N_5244,N_4952);
nand U5548 (N_5548,N_4985,N_5133);
nand U5549 (N_5549,N_4853,N_4957);
xor U5550 (N_5550,N_5048,N_5018);
nand U5551 (N_5551,N_4680,N_4788);
xnor U5552 (N_5552,N_4755,N_4903);
xor U5553 (N_5553,N_5086,N_4808);
and U5554 (N_5554,N_5114,N_4595);
xnor U5555 (N_5555,N_4911,N_4528);
xnor U5556 (N_5556,N_5063,N_4654);
nand U5557 (N_5557,N_5157,N_4600);
or U5558 (N_5558,N_5144,N_4783);
and U5559 (N_5559,N_4729,N_5149);
nor U5560 (N_5560,N_4508,N_4848);
nand U5561 (N_5561,N_5148,N_4785);
xnor U5562 (N_5562,N_5228,N_5081);
and U5563 (N_5563,N_5233,N_4766);
or U5564 (N_5564,N_4701,N_5142);
and U5565 (N_5565,N_5055,N_4576);
nand U5566 (N_5566,N_4705,N_4811);
and U5567 (N_5567,N_4531,N_4827);
and U5568 (N_5568,N_4570,N_5188);
xnor U5569 (N_5569,N_4550,N_4780);
xnor U5570 (N_5570,N_4634,N_5072);
or U5571 (N_5571,N_5165,N_5083);
nor U5572 (N_5572,N_5098,N_5152);
or U5573 (N_5573,N_4533,N_5070);
xnor U5574 (N_5574,N_5146,N_4720);
nand U5575 (N_5575,N_4682,N_5224);
or U5576 (N_5576,N_4587,N_5218);
nand U5577 (N_5577,N_5199,N_5059);
or U5578 (N_5578,N_4795,N_4860);
nor U5579 (N_5579,N_4628,N_5043);
and U5580 (N_5580,N_5031,N_4773);
and U5581 (N_5581,N_4950,N_4580);
nand U5582 (N_5582,N_4740,N_5191);
nor U5583 (N_5583,N_4845,N_5009);
and U5584 (N_5584,N_4597,N_4601);
or U5585 (N_5585,N_4603,N_4616);
and U5586 (N_5586,N_4898,N_4988);
nand U5587 (N_5587,N_4842,N_5076);
nor U5588 (N_5588,N_4564,N_4627);
and U5589 (N_5589,N_4784,N_4970);
nor U5590 (N_5590,N_4789,N_4958);
nand U5591 (N_5591,N_4802,N_4577);
or U5592 (N_5592,N_5194,N_4791);
and U5593 (N_5593,N_4675,N_4667);
xnor U5594 (N_5594,N_5032,N_4609);
nor U5595 (N_5595,N_4859,N_4583);
nand U5596 (N_5596,N_4871,N_4652);
nand U5597 (N_5597,N_4741,N_5163);
xor U5598 (N_5598,N_4502,N_4732);
nand U5599 (N_5599,N_5104,N_4793);
nand U5600 (N_5600,N_4512,N_5058);
or U5601 (N_5601,N_4639,N_4532);
nand U5602 (N_5602,N_5155,N_4865);
nand U5603 (N_5603,N_4547,N_4919);
nand U5604 (N_5604,N_4529,N_4650);
and U5605 (N_5605,N_4807,N_4509);
and U5606 (N_5606,N_4828,N_5120);
xor U5607 (N_5607,N_4657,N_5060);
or U5608 (N_5608,N_5131,N_5096);
nor U5609 (N_5609,N_5169,N_5214);
nand U5610 (N_5610,N_4622,N_5243);
nor U5611 (N_5611,N_4569,N_4610);
nand U5612 (N_5612,N_4833,N_4943);
xor U5613 (N_5613,N_5187,N_4856);
xnor U5614 (N_5614,N_5150,N_4534);
nand U5615 (N_5615,N_4575,N_4960);
nor U5616 (N_5616,N_4545,N_4796);
nor U5617 (N_5617,N_4615,N_4923);
nor U5618 (N_5618,N_5082,N_5068);
nand U5619 (N_5619,N_4998,N_4591);
or U5620 (N_5620,N_4814,N_4713);
and U5621 (N_5621,N_4556,N_4979);
nand U5622 (N_5622,N_4726,N_5166);
and U5623 (N_5623,N_4716,N_4926);
and U5624 (N_5624,N_4775,N_4850);
xor U5625 (N_5625,N_4575,N_4628);
or U5626 (N_5626,N_4539,N_5008);
nand U5627 (N_5627,N_4853,N_4977);
nor U5628 (N_5628,N_4912,N_4902);
or U5629 (N_5629,N_5127,N_4563);
and U5630 (N_5630,N_4634,N_4771);
or U5631 (N_5631,N_4811,N_5022);
or U5632 (N_5632,N_4907,N_4651);
nor U5633 (N_5633,N_4991,N_4505);
or U5634 (N_5634,N_4764,N_4567);
nand U5635 (N_5635,N_4833,N_4962);
and U5636 (N_5636,N_5144,N_5032);
nand U5637 (N_5637,N_4619,N_5044);
nand U5638 (N_5638,N_5187,N_4977);
and U5639 (N_5639,N_4881,N_4918);
and U5640 (N_5640,N_5058,N_4833);
or U5641 (N_5641,N_5119,N_4681);
xor U5642 (N_5642,N_4651,N_5169);
and U5643 (N_5643,N_4652,N_4639);
nor U5644 (N_5644,N_4549,N_5249);
xnor U5645 (N_5645,N_5247,N_4524);
or U5646 (N_5646,N_5228,N_4968);
nor U5647 (N_5647,N_4865,N_4850);
nor U5648 (N_5648,N_4501,N_5099);
or U5649 (N_5649,N_4924,N_4574);
xor U5650 (N_5650,N_4728,N_5029);
nand U5651 (N_5651,N_4540,N_5076);
xnor U5652 (N_5652,N_4757,N_4621);
and U5653 (N_5653,N_4602,N_4827);
xnor U5654 (N_5654,N_4795,N_4601);
nand U5655 (N_5655,N_4698,N_5231);
or U5656 (N_5656,N_5143,N_4766);
xnor U5657 (N_5657,N_4944,N_5138);
nand U5658 (N_5658,N_4958,N_5021);
nor U5659 (N_5659,N_4706,N_4811);
nor U5660 (N_5660,N_4549,N_4838);
xor U5661 (N_5661,N_5198,N_5008);
xnor U5662 (N_5662,N_4969,N_4738);
nand U5663 (N_5663,N_4613,N_5085);
and U5664 (N_5664,N_4573,N_4914);
nor U5665 (N_5665,N_5128,N_5075);
nand U5666 (N_5666,N_4785,N_4846);
nand U5667 (N_5667,N_4678,N_5083);
nand U5668 (N_5668,N_4741,N_4506);
nand U5669 (N_5669,N_4564,N_4646);
xor U5670 (N_5670,N_5055,N_4503);
xor U5671 (N_5671,N_4985,N_5166);
xnor U5672 (N_5672,N_4964,N_4583);
or U5673 (N_5673,N_4737,N_5218);
and U5674 (N_5674,N_4893,N_5176);
or U5675 (N_5675,N_5012,N_5118);
xnor U5676 (N_5676,N_4814,N_4763);
or U5677 (N_5677,N_5141,N_5072);
nand U5678 (N_5678,N_4696,N_4957);
and U5679 (N_5679,N_4527,N_4637);
nand U5680 (N_5680,N_4691,N_5005);
nor U5681 (N_5681,N_4807,N_5146);
nor U5682 (N_5682,N_5010,N_4664);
nor U5683 (N_5683,N_4564,N_5082);
nor U5684 (N_5684,N_4980,N_5212);
and U5685 (N_5685,N_5241,N_4645);
and U5686 (N_5686,N_4618,N_4947);
xnor U5687 (N_5687,N_4637,N_5211);
xnor U5688 (N_5688,N_5090,N_4669);
xnor U5689 (N_5689,N_5215,N_4556);
nand U5690 (N_5690,N_5192,N_5064);
nor U5691 (N_5691,N_5152,N_4709);
xnor U5692 (N_5692,N_4972,N_4578);
nor U5693 (N_5693,N_4554,N_4930);
or U5694 (N_5694,N_4744,N_4929);
or U5695 (N_5695,N_5122,N_5022);
or U5696 (N_5696,N_4925,N_4868);
nor U5697 (N_5697,N_5126,N_4730);
nand U5698 (N_5698,N_4962,N_4993);
and U5699 (N_5699,N_5057,N_4522);
and U5700 (N_5700,N_4954,N_4537);
nand U5701 (N_5701,N_4610,N_5221);
xnor U5702 (N_5702,N_4976,N_4539);
xnor U5703 (N_5703,N_4931,N_4868);
nor U5704 (N_5704,N_5208,N_4778);
nand U5705 (N_5705,N_5056,N_4804);
or U5706 (N_5706,N_4676,N_4545);
and U5707 (N_5707,N_5230,N_5233);
and U5708 (N_5708,N_5046,N_4621);
nor U5709 (N_5709,N_5109,N_4882);
and U5710 (N_5710,N_4997,N_4786);
nor U5711 (N_5711,N_4606,N_4850);
and U5712 (N_5712,N_4509,N_4613);
xor U5713 (N_5713,N_5148,N_5214);
or U5714 (N_5714,N_5237,N_5040);
or U5715 (N_5715,N_4823,N_4613);
and U5716 (N_5716,N_5206,N_4612);
nand U5717 (N_5717,N_4906,N_5105);
and U5718 (N_5718,N_5005,N_4986);
and U5719 (N_5719,N_4855,N_4858);
nor U5720 (N_5720,N_4967,N_4957);
xnor U5721 (N_5721,N_4855,N_4946);
nand U5722 (N_5722,N_4857,N_4766);
and U5723 (N_5723,N_4510,N_4573);
nand U5724 (N_5724,N_5202,N_5123);
or U5725 (N_5725,N_4599,N_4596);
nand U5726 (N_5726,N_4749,N_4804);
or U5727 (N_5727,N_4594,N_4524);
or U5728 (N_5728,N_5010,N_5081);
xor U5729 (N_5729,N_4841,N_4810);
or U5730 (N_5730,N_4540,N_4974);
nand U5731 (N_5731,N_4826,N_4989);
xnor U5732 (N_5732,N_4505,N_4614);
nor U5733 (N_5733,N_4610,N_4780);
xor U5734 (N_5734,N_4582,N_4773);
nor U5735 (N_5735,N_5047,N_5145);
or U5736 (N_5736,N_4743,N_4735);
xor U5737 (N_5737,N_4534,N_4946);
nor U5738 (N_5738,N_4805,N_4759);
nor U5739 (N_5739,N_4570,N_5143);
and U5740 (N_5740,N_4700,N_4936);
or U5741 (N_5741,N_4921,N_4961);
nor U5742 (N_5742,N_5163,N_4561);
xor U5743 (N_5743,N_4706,N_4548);
or U5744 (N_5744,N_4772,N_5044);
and U5745 (N_5745,N_4782,N_4761);
and U5746 (N_5746,N_4983,N_4812);
or U5747 (N_5747,N_4587,N_4679);
nand U5748 (N_5748,N_4890,N_5020);
or U5749 (N_5749,N_5120,N_4616);
xnor U5750 (N_5750,N_5201,N_4639);
nand U5751 (N_5751,N_4506,N_4768);
and U5752 (N_5752,N_5176,N_4998);
xnor U5753 (N_5753,N_4754,N_4595);
nand U5754 (N_5754,N_4873,N_4671);
and U5755 (N_5755,N_5044,N_4999);
xor U5756 (N_5756,N_4927,N_4966);
and U5757 (N_5757,N_4679,N_4928);
or U5758 (N_5758,N_4857,N_5206);
or U5759 (N_5759,N_4860,N_4715);
and U5760 (N_5760,N_5226,N_5133);
nor U5761 (N_5761,N_4638,N_5248);
or U5762 (N_5762,N_4676,N_4673);
xor U5763 (N_5763,N_5073,N_4983);
nand U5764 (N_5764,N_5017,N_4919);
nand U5765 (N_5765,N_4854,N_4701);
or U5766 (N_5766,N_4727,N_5246);
and U5767 (N_5767,N_5117,N_5027);
nor U5768 (N_5768,N_4767,N_4583);
nand U5769 (N_5769,N_4902,N_5071);
xor U5770 (N_5770,N_5192,N_4821);
and U5771 (N_5771,N_4990,N_4586);
nor U5772 (N_5772,N_5128,N_4587);
or U5773 (N_5773,N_4588,N_4960);
nand U5774 (N_5774,N_4560,N_4905);
xnor U5775 (N_5775,N_4608,N_5249);
or U5776 (N_5776,N_4820,N_4503);
and U5777 (N_5777,N_5165,N_4732);
or U5778 (N_5778,N_5147,N_4583);
nand U5779 (N_5779,N_5043,N_5168);
xnor U5780 (N_5780,N_4962,N_5002);
nor U5781 (N_5781,N_4816,N_4520);
and U5782 (N_5782,N_4570,N_5187);
nor U5783 (N_5783,N_4839,N_4939);
and U5784 (N_5784,N_4710,N_5057);
or U5785 (N_5785,N_5214,N_4777);
or U5786 (N_5786,N_4689,N_4564);
nor U5787 (N_5787,N_4601,N_4572);
or U5788 (N_5788,N_5180,N_4827);
or U5789 (N_5789,N_5035,N_4876);
xor U5790 (N_5790,N_4664,N_4604);
and U5791 (N_5791,N_4898,N_4524);
and U5792 (N_5792,N_4869,N_4714);
or U5793 (N_5793,N_5029,N_5173);
nor U5794 (N_5794,N_5163,N_4918);
and U5795 (N_5795,N_4689,N_4656);
or U5796 (N_5796,N_4868,N_4917);
or U5797 (N_5797,N_4573,N_5032);
nor U5798 (N_5798,N_4970,N_4701);
xnor U5799 (N_5799,N_5245,N_5055);
nor U5800 (N_5800,N_5151,N_4764);
or U5801 (N_5801,N_5192,N_5205);
nor U5802 (N_5802,N_4767,N_4875);
xnor U5803 (N_5803,N_4909,N_4619);
and U5804 (N_5804,N_4818,N_4868);
nor U5805 (N_5805,N_5055,N_4969);
nor U5806 (N_5806,N_4869,N_4533);
nand U5807 (N_5807,N_4519,N_4723);
xor U5808 (N_5808,N_5125,N_4868);
xor U5809 (N_5809,N_5222,N_5161);
or U5810 (N_5810,N_4880,N_4718);
or U5811 (N_5811,N_4778,N_4866);
nand U5812 (N_5812,N_4816,N_5231);
nor U5813 (N_5813,N_5040,N_4766);
nor U5814 (N_5814,N_4902,N_4988);
nand U5815 (N_5815,N_4732,N_5189);
or U5816 (N_5816,N_5153,N_4780);
and U5817 (N_5817,N_5114,N_5063);
nand U5818 (N_5818,N_4963,N_5067);
and U5819 (N_5819,N_4761,N_5001);
or U5820 (N_5820,N_4529,N_4990);
xnor U5821 (N_5821,N_4857,N_5184);
nand U5822 (N_5822,N_4701,N_5088);
nor U5823 (N_5823,N_4814,N_4858);
xnor U5824 (N_5824,N_4839,N_5035);
xor U5825 (N_5825,N_4755,N_4758);
nand U5826 (N_5826,N_4806,N_4705);
nand U5827 (N_5827,N_4513,N_4540);
nor U5828 (N_5828,N_5220,N_4908);
nand U5829 (N_5829,N_5127,N_4900);
or U5830 (N_5830,N_5010,N_4712);
or U5831 (N_5831,N_5101,N_5084);
and U5832 (N_5832,N_5109,N_5020);
xnor U5833 (N_5833,N_4794,N_5143);
nand U5834 (N_5834,N_4854,N_4757);
and U5835 (N_5835,N_4909,N_4663);
and U5836 (N_5836,N_4615,N_5080);
nand U5837 (N_5837,N_4821,N_5043);
nand U5838 (N_5838,N_4542,N_4629);
xnor U5839 (N_5839,N_4866,N_5122);
nand U5840 (N_5840,N_4888,N_5248);
xor U5841 (N_5841,N_4956,N_5172);
or U5842 (N_5842,N_4628,N_4894);
and U5843 (N_5843,N_5063,N_5104);
and U5844 (N_5844,N_4549,N_5089);
and U5845 (N_5845,N_4702,N_4579);
and U5846 (N_5846,N_4630,N_4906);
nand U5847 (N_5847,N_4785,N_5122);
and U5848 (N_5848,N_4881,N_4519);
xnor U5849 (N_5849,N_5230,N_4535);
or U5850 (N_5850,N_4582,N_4793);
nand U5851 (N_5851,N_4531,N_5189);
nor U5852 (N_5852,N_4931,N_5125);
nor U5853 (N_5853,N_4742,N_4673);
or U5854 (N_5854,N_5142,N_4985);
xnor U5855 (N_5855,N_4894,N_5220);
and U5856 (N_5856,N_5043,N_4566);
and U5857 (N_5857,N_4903,N_4943);
nor U5858 (N_5858,N_4794,N_5111);
and U5859 (N_5859,N_4684,N_4773);
or U5860 (N_5860,N_4619,N_4767);
nand U5861 (N_5861,N_4640,N_4700);
or U5862 (N_5862,N_4702,N_5026);
nor U5863 (N_5863,N_4731,N_5166);
xnor U5864 (N_5864,N_4601,N_4893);
and U5865 (N_5865,N_5211,N_4813);
and U5866 (N_5866,N_4541,N_4985);
xor U5867 (N_5867,N_4810,N_5137);
nand U5868 (N_5868,N_5237,N_4814);
xor U5869 (N_5869,N_4717,N_4501);
xor U5870 (N_5870,N_4893,N_4932);
and U5871 (N_5871,N_4908,N_5167);
and U5872 (N_5872,N_5144,N_5025);
nand U5873 (N_5873,N_4744,N_4932);
or U5874 (N_5874,N_5194,N_5226);
nor U5875 (N_5875,N_5115,N_5033);
nand U5876 (N_5876,N_5210,N_5038);
nand U5877 (N_5877,N_5004,N_4541);
or U5878 (N_5878,N_4768,N_4718);
nor U5879 (N_5879,N_5059,N_5169);
and U5880 (N_5880,N_4701,N_4561);
xor U5881 (N_5881,N_5117,N_5042);
xor U5882 (N_5882,N_4979,N_4783);
nor U5883 (N_5883,N_5036,N_4944);
xnor U5884 (N_5884,N_5012,N_4793);
and U5885 (N_5885,N_4810,N_5242);
or U5886 (N_5886,N_4784,N_4763);
nor U5887 (N_5887,N_4961,N_4627);
or U5888 (N_5888,N_4541,N_4780);
nand U5889 (N_5889,N_4955,N_4626);
xnor U5890 (N_5890,N_4671,N_4644);
nand U5891 (N_5891,N_4503,N_5182);
and U5892 (N_5892,N_4858,N_4619);
nor U5893 (N_5893,N_4993,N_4813);
or U5894 (N_5894,N_5189,N_4786);
nor U5895 (N_5895,N_4821,N_5112);
xnor U5896 (N_5896,N_4907,N_4898);
and U5897 (N_5897,N_4506,N_4875);
xor U5898 (N_5898,N_4828,N_4662);
xor U5899 (N_5899,N_4553,N_4793);
xor U5900 (N_5900,N_5210,N_5186);
nand U5901 (N_5901,N_4630,N_5086);
and U5902 (N_5902,N_4639,N_4744);
nor U5903 (N_5903,N_5214,N_4715);
and U5904 (N_5904,N_4777,N_4815);
or U5905 (N_5905,N_5015,N_4842);
and U5906 (N_5906,N_4804,N_4969);
nor U5907 (N_5907,N_4795,N_4661);
xor U5908 (N_5908,N_5140,N_4847);
or U5909 (N_5909,N_4782,N_5052);
nand U5910 (N_5910,N_4541,N_5061);
or U5911 (N_5911,N_4581,N_4645);
nor U5912 (N_5912,N_4529,N_4880);
nand U5913 (N_5913,N_4961,N_4538);
or U5914 (N_5914,N_5118,N_4779);
xnor U5915 (N_5915,N_4877,N_4614);
xor U5916 (N_5916,N_5113,N_4655);
and U5917 (N_5917,N_4539,N_4985);
nor U5918 (N_5918,N_4757,N_5189);
nand U5919 (N_5919,N_4565,N_4819);
nand U5920 (N_5920,N_4505,N_4582);
xor U5921 (N_5921,N_4626,N_4810);
and U5922 (N_5922,N_5239,N_4899);
xnor U5923 (N_5923,N_4806,N_5185);
nand U5924 (N_5924,N_5203,N_5020);
xnor U5925 (N_5925,N_5107,N_4721);
nand U5926 (N_5926,N_5056,N_4692);
and U5927 (N_5927,N_4971,N_4589);
nor U5928 (N_5928,N_5042,N_4837);
nor U5929 (N_5929,N_4905,N_4554);
xnor U5930 (N_5930,N_5230,N_4767);
or U5931 (N_5931,N_4736,N_4877);
nand U5932 (N_5932,N_4596,N_4594);
or U5933 (N_5933,N_4764,N_5118);
and U5934 (N_5934,N_5100,N_4897);
xor U5935 (N_5935,N_5027,N_5243);
or U5936 (N_5936,N_4818,N_4731);
and U5937 (N_5937,N_4927,N_4742);
and U5938 (N_5938,N_4942,N_4956);
xnor U5939 (N_5939,N_4666,N_4739);
or U5940 (N_5940,N_4979,N_4688);
nand U5941 (N_5941,N_5126,N_5034);
nor U5942 (N_5942,N_4849,N_5003);
nand U5943 (N_5943,N_5137,N_4795);
or U5944 (N_5944,N_5189,N_4709);
nand U5945 (N_5945,N_5034,N_5210);
or U5946 (N_5946,N_5041,N_5079);
and U5947 (N_5947,N_5052,N_4775);
or U5948 (N_5948,N_5150,N_4743);
xnor U5949 (N_5949,N_4825,N_4949);
xnor U5950 (N_5950,N_4959,N_5225);
xnor U5951 (N_5951,N_5249,N_4557);
or U5952 (N_5952,N_4629,N_4860);
or U5953 (N_5953,N_4524,N_4644);
or U5954 (N_5954,N_4963,N_5199);
nand U5955 (N_5955,N_4564,N_4600);
nor U5956 (N_5956,N_5220,N_4745);
or U5957 (N_5957,N_4679,N_4961);
and U5958 (N_5958,N_5096,N_5048);
nand U5959 (N_5959,N_5107,N_5191);
nor U5960 (N_5960,N_4865,N_5020);
xnor U5961 (N_5961,N_4709,N_4757);
xnor U5962 (N_5962,N_5143,N_4803);
and U5963 (N_5963,N_4610,N_4615);
nor U5964 (N_5964,N_4641,N_5143);
nand U5965 (N_5965,N_4850,N_5045);
nor U5966 (N_5966,N_5117,N_4562);
nand U5967 (N_5967,N_4864,N_4555);
or U5968 (N_5968,N_4801,N_4959);
or U5969 (N_5969,N_4517,N_5027);
and U5970 (N_5970,N_4755,N_5163);
nor U5971 (N_5971,N_4999,N_4833);
nor U5972 (N_5972,N_4894,N_5233);
nor U5973 (N_5973,N_5227,N_5228);
and U5974 (N_5974,N_4693,N_4582);
nor U5975 (N_5975,N_4738,N_5019);
nor U5976 (N_5976,N_4932,N_4729);
xnor U5977 (N_5977,N_4575,N_4521);
nand U5978 (N_5978,N_4895,N_4903);
nor U5979 (N_5979,N_4523,N_4743);
and U5980 (N_5980,N_5128,N_4990);
nor U5981 (N_5981,N_4980,N_5136);
xnor U5982 (N_5982,N_4969,N_5069);
nor U5983 (N_5983,N_4767,N_5063);
nor U5984 (N_5984,N_5196,N_4616);
nand U5985 (N_5985,N_5029,N_4660);
nand U5986 (N_5986,N_4509,N_4840);
and U5987 (N_5987,N_5233,N_4927);
and U5988 (N_5988,N_4880,N_4891);
nor U5989 (N_5989,N_5059,N_4773);
or U5990 (N_5990,N_4650,N_4727);
or U5991 (N_5991,N_4882,N_4521);
nand U5992 (N_5992,N_4725,N_4818);
xor U5993 (N_5993,N_4631,N_4667);
nand U5994 (N_5994,N_4534,N_4732);
xor U5995 (N_5995,N_5185,N_4618);
nor U5996 (N_5996,N_4600,N_4901);
nor U5997 (N_5997,N_4974,N_4959);
xnor U5998 (N_5998,N_4659,N_5095);
nor U5999 (N_5999,N_5023,N_4591);
nand U6000 (N_6000,N_5820,N_5695);
and U6001 (N_6001,N_5311,N_5964);
nor U6002 (N_6002,N_5752,N_5434);
nand U6003 (N_6003,N_5508,N_5324);
nand U6004 (N_6004,N_5488,N_5347);
nand U6005 (N_6005,N_5750,N_5720);
nand U6006 (N_6006,N_5559,N_5393);
nand U6007 (N_6007,N_5723,N_5575);
xnor U6008 (N_6008,N_5682,N_5277);
and U6009 (N_6009,N_5388,N_5961);
nor U6010 (N_6010,N_5350,N_5638);
or U6011 (N_6011,N_5477,N_5300);
nand U6012 (N_6012,N_5813,N_5557);
nand U6013 (N_6013,N_5704,N_5965);
nand U6014 (N_6014,N_5810,N_5861);
nand U6015 (N_6015,N_5370,N_5514);
nor U6016 (N_6016,N_5394,N_5613);
xor U6017 (N_6017,N_5743,N_5878);
and U6018 (N_6018,N_5670,N_5609);
or U6019 (N_6019,N_5969,N_5472);
nand U6020 (N_6020,N_5864,N_5710);
or U6021 (N_6021,N_5905,N_5569);
and U6022 (N_6022,N_5732,N_5921);
nor U6023 (N_6023,N_5698,N_5286);
or U6024 (N_6024,N_5322,N_5589);
nand U6025 (N_6025,N_5292,N_5503);
nor U6026 (N_6026,N_5594,N_5500);
nor U6027 (N_6027,N_5680,N_5600);
nor U6028 (N_6028,N_5577,N_5928);
xnor U6029 (N_6029,N_5829,N_5886);
xor U6030 (N_6030,N_5741,N_5789);
nor U6031 (N_6031,N_5769,N_5954);
or U6032 (N_6032,N_5296,N_5615);
or U6033 (N_6033,N_5592,N_5858);
or U6034 (N_6034,N_5812,N_5379);
and U6035 (N_6035,N_5733,N_5661);
or U6036 (N_6036,N_5908,N_5840);
nand U6037 (N_6037,N_5546,N_5626);
nand U6038 (N_6038,N_5448,N_5711);
nor U6039 (N_6039,N_5304,N_5360);
nor U6040 (N_6040,N_5293,N_5980);
nor U6041 (N_6041,N_5250,N_5894);
nor U6042 (N_6042,N_5962,N_5562);
xnor U6043 (N_6043,N_5409,N_5618);
nand U6044 (N_6044,N_5631,N_5993);
nor U6045 (N_6045,N_5355,N_5767);
nand U6046 (N_6046,N_5456,N_5391);
nand U6047 (N_6047,N_5702,N_5268);
xor U6048 (N_6048,N_5591,N_5349);
or U6049 (N_6049,N_5478,N_5623);
nor U6050 (N_6050,N_5313,N_5992);
and U6051 (N_6051,N_5329,N_5653);
and U6052 (N_6052,N_5650,N_5932);
or U6053 (N_6053,N_5648,N_5983);
and U6054 (N_6054,N_5298,N_5404);
and U6055 (N_6055,N_5490,N_5299);
and U6056 (N_6056,N_5572,N_5947);
nand U6057 (N_6057,N_5454,N_5558);
and U6058 (N_6058,N_5553,N_5466);
xnor U6059 (N_6059,N_5551,N_5328);
nor U6060 (N_6060,N_5746,N_5302);
nand U6061 (N_6061,N_5869,N_5392);
xor U6062 (N_6062,N_5889,N_5629);
and U6063 (N_6063,N_5607,N_5441);
or U6064 (N_6064,N_5469,N_5593);
nand U6065 (N_6065,N_5757,N_5474);
and U6066 (N_6066,N_5522,N_5865);
xor U6067 (N_6067,N_5571,N_5678);
nor U6068 (N_6068,N_5532,N_5544);
and U6069 (N_6069,N_5978,N_5616);
nand U6070 (N_6070,N_5307,N_5586);
and U6071 (N_6071,N_5990,N_5420);
xnor U6072 (N_6072,N_5914,N_5449);
nor U6073 (N_6073,N_5495,N_5583);
nand U6074 (N_6074,N_5975,N_5948);
nand U6075 (N_6075,N_5815,N_5418);
or U6076 (N_6076,N_5870,N_5570);
xor U6077 (N_6077,N_5791,N_5367);
nor U6078 (N_6078,N_5554,N_5933);
and U6079 (N_6079,N_5552,N_5854);
and U6080 (N_6080,N_5986,N_5749);
nor U6081 (N_6081,N_5771,N_5816);
or U6082 (N_6082,N_5663,N_5734);
nand U6083 (N_6083,N_5587,N_5867);
nand U6084 (N_6084,N_5874,N_5599);
nor U6085 (N_6085,N_5943,N_5737);
and U6086 (N_6086,N_5502,N_5797);
nand U6087 (N_6087,N_5460,N_5263);
nor U6088 (N_6088,N_5967,N_5691);
or U6089 (N_6089,N_5841,N_5303);
xnor U6090 (N_6090,N_5317,N_5410);
xnor U6091 (N_6091,N_5278,N_5251);
and U6092 (N_6092,N_5727,N_5868);
xor U6093 (N_6093,N_5848,N_5373);
and U6094 (N_6094,N_5540,N_5729);
nor U6095 (N_6095,N_5550,N_5545);
nor U6096 (N_6096,N_5316,N_5288);
nand U6097 (N_6097,N_5622,N_5452);
nand U6098 (N_6098,N_5708,N_5800);
xnor U6099 (N_6099,N_5739,N_5672);
xnor U6100 (N_6100,N_5686,N_5972);
and U6101 (N_6101,N_5651,N_5376);
xor U6102 (N_6102,N_5389,N_5779);
nand U6103 (N_6103,N_5805,N_5337);
and U6104 (N_6104,N_5447,N_5463);
nor U6105 (N_6105,N_5818,N_5758);
or U6106 (N_6106,N_5802,N_5366);
nor U6107 (N_6107,N_5679,N_5542);
xnor U6108 (N_6108,N_5291,N_5639);
xnor U6109 (N_6109,N_5736,N_5910);
and U6110 (N_6110,N_5520,N_5976);
nor U6111 (N_6111,N_5541,N_5768);
nand U6112 (N_6112,N_5276,N_5357);
xor U6113 (N_6113,N_5269,N_5261);
nand U6114 (N_6114,N_5432,N_5926);
and U6115 (N_6115,N_5836,N_5877);
and U6116 (N_6116,N_5517,N_5283);
nand U6117 (N_6117,N_5635,N_5342);
xnor U6118 (N_6118,N_5382,N_5385);
nand U6119 (N_6119,N_5429,N_5735);
and U6120 (N_6120,N_5703,N_5344);
nor U6121 (N_6121,N_5282,N_5774);
or U6122 (N_6122,N_5946,N_5660);
nor U6123 (N_6123,N_5755,N_5989);
or U6124 (N_6124,N_5785,N_5406);
nor U6125 (N_6125,N_5515,N_5970);
or U6126 (N_6126,N_5476,N_5484);
nand U6127 (N_6127,N_5584,N_5333);
and U6128 (N_6128,N_5931,N_5462);
xor U6129 (N_6129,N_5614,N_5369);
nand U6130 (N_6130,N_5362,N_5919);
and U6131 (N_6131,N_5527,N_5359);
xnor U6132 (N_6132,N_5364,N_5999);
nand U6133 (N_6133,N_5753,N_5601);
and U6134 (N_6134,N_5851,N_5904);
and U6135 (N_6135,N_5425,N_5953);
nand U6136 (N_6136,N_5890,N_5819);
nand U6137 (N_6137,N_5352,N_5803);
or U6138 (N_6138,N_5827,N_5808);
xor U6139 (N_6139,N_5879,N_5578);
and U6140 (N_6140,N_5321,N_5984);
or U6141 (N_6141,N_5855,N_5290);
and U6142 (N_6142,N_5795,N_5830);
or U6143 (N_6143,N_5413,N_5852);
xor U6144 (N_6144,N_5777,N_5881);
nor U6145 (N_6145,N_5966,N_5512);
and U6146 (N_6146,N_5788,N_5822);
or U6147 (N_6147,N_5939,N_5900);
nand U6148 (N_6148,N_5880,N_5323);
or U6149 (N_6149,N_5825,N_5973);
and U6150 (N_6150,N_5315,N_5636);
and U6151 (N_6151,N_5343,N_5747);
nor U6152 (N_6152,N_5941,N_5937);
nor U6153 (N_6153,N_5794,N_5977);
nand U6154 (N_6154,N_5690,N_5312);
nor U6155 (N_6155,N_5915,N_5902);
xnor U6156 (N_6156,N_5439,N_5627);
nor U6157 (N_6157,N_5778,N_5776);
and U6158 (N_6158,N_5790,N_5811);
and U6159 (N_6159,N_5624,N_5403);
or U6160 (N_6160,N_5922,N_5923);
xnor U6161 (N_6161,N_5294,N_5445);
nor U6162 (N_6162,N_5763,N_5875);
or U6163 (N_6163,N_5700,N_5421);
nand U6164 (N_6164,N_5668,N_5345);
nor U6165 (N_6165,N_5893,N_5492);
and U6166 (N_6166,N_5309,N_5565);
xor U6167 (N_6167,N_5634,N_5892);
nor U6168 (N_6168,N_5949,N_5386);
xnor U6169 (N_6169,N_5787,N_5356);
or U6170 (N_6170,N_5724,N_5494);
nand U6171 (N_6171,N_5762,N_5659);
xor U6172 (N_6172,N_5516,N_5860);
and U6173 (N_6173,N_5457,N_5399);
or U6174 (N_6174,N_5731,N_5505);
xnor U6175 (N_6175,N_5912,N_5719);
nand U6176 (N_6176,N_5862,N_5598);
nand U6177 (N_6177,N_5524,N_5301);
nor U6178 (N_6178,N_5930,N_5485);
nand U6179 (N_6179,N_5507,N_5574);
and U6180 (N_6180,N_5252,N_5971);
nor U6181 (N_6181,N_5561,N_5433);
nor U6182 (N_6182,N_5845,N_5667);
xnor U6183 (N_6183,N_5467,N_5533);
nand U6184 (N_6184,N_5426,N_5444);
or U6185 (N_6185,N_5612,N_5371);
nand U6186 (N_6186,N_5258,N_5712);
or U6187 (N_6187,N_5674,N_5715);
nand U6188 (N_6188,N_5677,N_5491);
and U6189 (N_6189,N_5279,N_5306);
and U6190 (N_6190,N_5833,N_5450);
and U6191 (N_6191,N_5253,N_5863);
or U6192 (N_6192,N_5260,N_5633);
and U6193 (N_6193,N_5395,N_5468);
nor U6194 (N_6194,N_5821,N_5496);
or U6195 (N_6195,N_5699,N_5871);
or U6196 (N_6196,N_5611,N_5873);
nand U6197 (N_6197,N_5617,N_5459);
and U6198 (N_6198,N_5424,N_5824);
and U6199 (N_6199,N_5435,N_5605);
nand U6200 (N_6200,N_5907,N_5801);
nor U6201 (N_6201,N_5843,N_5740);
nand U6202 (N_6202,N_5722,N_5354);
or U6203 (N_6203,N_5254,N_5866);
and U6204 (N_6204,N_5957,N_5257);
xnor U6205 (N_6205,N_5657,N_5480);
or U6206 (N_6206,N_5806,N_5585);
or U6207 (N_6207,N_5856,N_5645);
and U6208 (N_6208,N_5673,N_5798);
and U6209 (N_6209,N_5835,N_5671);
nor U6210 (N_6210,N_5728,N_5308);
and U6211 (N_6211,N_5455,N_5332);
xor U6212 (N_6212,N_5760,N_5628);
nor U6213 (N_6213,N_5676,N_5267);
xor U6214 (N_6214,N_5272,N_5918);
and U6215 (N_6215,N_5259,N_5473);
or U6216 (N_6216,N_5378,N_5994);
and U6217 (N_6217,N_5264,N_5408);
xnor U6218 (N_6218,N_5506,N_5883);
and U6219 (N_6219,N_5658,N_5952);
or U6220 (N_6220,N_5581,N_5898);
xnor U6221 (N_6221,N_5325,N_5310);
or U6222 (N_6222,N_5925,N_5440);
nor U6223 (N_6223,N_5896,N_5602);
nand U6224 (N_6224,N_5353,N_5265);
nor U6225 (N_6225,N_5956,N_5335);
nor U6226 (N_6226,N_5374,N_5564);
nand U6227 (N_6227,N_5535,N_5887);
nand U6228 (N_6228,N_5847,N_5996);
nand U6229 (N_6229,N_5979,N_5909);
or U6230 (N_6230,N_5475,N_5619);
xor U6231 (N_6231,N_5662,N_5358);
nand U6232 (N_6232,N_5998,N_5513);
and U6233 (N_6233,N_5706,N_5262);
nor U6234 (N_6234,N_5688,N_5529);
nor U6235 (N_6235,N_5375,N_5436);
nand U6236 (N_6236,N_5784,N_5580);
nor U6237 (N_6237,N_5804,N_5765);
nand U6238 (N_6238,N_5511,N_5327);
nand U6239 (N_6239,N_5539,N_5479);
nor U6240 (N_6240,N_5718,N_5786);
nand U6241 (N_6241,N_5643,N_5846);
nor U6242 (N_6242,N_5526,N_5528);
or U6243 (N_6243,N_5709,N_5576);
or U6244 (N_6244,N_5654,N_5701);
nor U6245 (N_6245,N_5536,N_5625);
xnor U6246 (N_6246,N_5920,N_5656);
nand U6247 (N_6247,N_5694,N_5717);
xnor U6248 (N_6248,N_5451,N_5518);
xnor U6249 (N_6249,N_5764,N_5693);
nand U6250 (N_6250,N_5828,N_5772);
or U6251 (N_6251,N_5853,N_5842);
or U6252 (N_6252,N_5481,N_5361);
or U6253 (N_6253,N_5275,N_5510);
and U6254 (N_6254,N_5320,N_5590);
and U6255 (N_6255,N_5761,N_5482);
nand U6256 (N_6256,N_5608,N_5555);
or U6257 (N_6257,N_5281,N_5895);
nand U6258 (N_6258,N_5669,N_5437);
nand U6259 (N_6259,N_5428,N_5716);
xor U6260 (N_6260,N_5443,N_5988);
nor U6261 (N_6261,N_5649,N_5940);
xor U6262 (N_6262,N_5560,N_5521);
or U6263 (N_6263,N_5461,N_5955);
nor U6264 (N_6264,N_5340,N_5547);
nand U6265 (N_6265,N_5446,N_5665);
nor U6266 (N_6266,N_5929,N_5775);
or U6267 (N_6267,N_5280,N_5348);
nand U6268 (N_6268,N_5346,N_5377);
nor U6269 (N_6269,N_5582,N_5568);
xor U6270 (N_6270,N_5341,N_5287);
nor U6271 (N_6271,N_5826,N_5982);
and U6272 (N_6272,N_5796,N_5684);
or U6273 (N_6273,N_5950,N_5334);
nor U6274 (N_6274,N_5738,N_5799);
nand U6275 (N_6275,N_5793,N_5872);
xor U6276 (N_6276,N_5351,N_5483);
and U6277 (N_6277,N_5464,N_5839);
nor U6278 (N_6278,N_5958,N_5405);
xor U6279 (N_6279,N_5255,N_5637);
nand U6280 (N_6280,N_5326,N_5981);
and U6281 (N_6281,N_5390,N_5917);
nor U6282 (N_6282,N_5906,N_5534);
or U6283 (N_6283,N_5604,N_5531);
nand U6284 (N_6284,N_5573,N_5832);
xnor U6285 (N_6285,N_5655,N_5438);
nand U6286 (N_6286,N_5504,N_5632);
and U6287 (N_6287,N_5530,N_5285);
nor U6288 (N_6288,N_5284,N_5543);
xnor U6289 (N_6289,N_5891,N_5620);
xnor U6290 (N_6290,N_5823,N_5417);
or U6291 (N_6291,N_5523,N_5271);
or U6292 (N_6292,N_5330,N_5742);
and U6293 (N_6293,N_5471,N_5899);
xnor U6294 (N_6294,N_5770,N_5336);
nor U6295 (N_6295,N_5882,N_5951);
or U6296 (N_6296,N_5959,N_5411);
nand U6297 (N_6297,N_5945,N_5713);
nor U6298 (N_6298,N_5640,N_5725);
nand U6299 (N_6299,N_5985,N_5419);
and U6300 (N_6300,N_5579,N_5876);
or U6301 (N_6301,N_5423,N_5934);
nor U6302 (N_6302,N_5331,N_5744);
and U6303 (N_6303,N_5487,N_5319);
or U6304 (N_6304,N_5606,N_5696);
nor U6305 (N_6305,N_5465,N_5781);
nor U6306 (N_6306,N_5556,N_5381);
nand U6307 (N_6307,N_5817,N_5901);
nand U6308 (N_6308,N_5519,N_5644);
or U6309 (N_6309,N_5603,N_5596);
xnor U6310 (N_6310,N_5647,N_5549);
nand U6311 (N_6311,N_5453,N_5683);
or U6312 (N_6312,N_5401,N_5857);
or U6313 (N_6313,N_5991,N_5652);
nand U6314 (N_6314,N_5266,N_5630);
or U6315 (N_6315,N_5697,N_5936);
nand U6316 (N_6316,N_5412,N_5563);
nand U6317 (N_6317,N_5498,N_5493);
nand U6318 (N_6318,N_5400,N_5458);
or U6319 (N_6319,N_5338,N_5685);
nor U6320 (N_6320,N_5675,N_5384);
xnor U6321 (N_6321,N_5692,N_5792);
nand U6322 (N_6322,N_5365,N_5814);
nand U6323 (N_6323,N_5916,N_5885);
xor U6324 (N_6324,N_5745,N_5714);
xor U6325 (N_6325,N_5646,N_5689);
nand U6326 (N_6326,N_5807,N_5256);
nand U6327 (N_6327,N_5363,N_5837);
and U6328 (N_6328,N_5809,N_5681);
xor U6329 (N_6329,N_5942,N_5430);
xor U6330 (N_6330,N_5730,N_5995);
and U6331 (N_6331,N_5289,N_5588);
xnor U6332 (N_6332,N_5431,N_5318);
nand U6333 (N_6333,N_5297,N_5759);
or U6334 (N_6334,N_5566,N_5295);
and U6335 (N_6335,N_5525,N_5372);
or U6336 (N_6336,N_5538,N_5913);
nor U6337 (N_6337,N_5402,N_5305);
xnor U6338 (N_6338,N_5497,N_5414);
nor U6339 (N_6339,N_5621,N_5888);
xor U6340 (N_6340,N_5567,N_5831);
and U6341 (N_6341,N_5415,N_5859);
nor U6342 (N_6342,N_5780,N_5968);
or U6343 (N_6343,N_5427,N_5844);
nand U6344 (N_6344,N_5754,N_5748);
and U6345 (N_6345,N_5642,N_5924);
and U6346 (N_6346,N_5610,N_5387);
nor U6347 (N_6347,N_5997,N_5773);
xor U6348 (N_6348,N_5687,N_5963);
nor U6349 (N_6349,N_5396,N_5489);
nand U6350 (N_6350,N_5721,N_5884);
xor U6351 (N_6351,N_5726,N_5903);
nor U6352 (N_6352,N_5897,N_5368);
or U6353 (N_6353,N_5274,N_5783);
nand U6354 (N_6354,N_5756,N_5664);
and U6355 (N_6355,N_5838,N_5849);
xor U6356 (N_6356,N_5442,N_5314);
nor U6357 (N_6357,N_5911,N_5944);
nand U6358 (N_6358,N_5927,N_5499);
and U6359 (N_6359,N_5987,N_5766);
xor U6360 (N_6360,N_5666,N_5850);
xor U6361 (N_6361,N_5974,N_5407);
xnor U6362 (N_6362,N_5537,N_5782);
nand U6363 (N_6363,N_5486,N_5509);
xnor U6364 (N_6364,N_5751,N_5383);
xnor U6365 (N_6365,N_5935,N_5416);
nor U6366 (N_6366,N_5705,N_5597);
nand U6367 (N_6367,N_5595,N_5273);
or U6368 (N_6368,N_5501,N_5270);
nor U6369 (N_6369,N_5422,N_5707);
nor U6370 (N_6370,N_5398,N_5470);
xor U6371 (N_6371,N_5938,N_5641);
nand U6372 (N_6372,N_5339,N_5380);
nor U6373 (N_6373,N_5960,N_5548);
or U6374 (N_6374,N_5834,N_5397);
xor U6375 (N_6375,N_5275,N_5785);
nand U6376 (N_6376,N_5428,N_5327);
xor U6377 (N_6377,N_5715,N_5655);
or U6378 (N_6378,N_5435,N_5592);
nor U6379 (N_6379,N_5879,N_5697);
nand U6380 (N_6380,N_5629,N_5750);
nor U6381 (N_6381,N_5720,N_5458);
and U6382 (N_6382,N_5937,N_5587);
and U6383 (N_6383,N_5641,N_5300);
and U6384 (N_6384,N_5497,N_5808);
xor U6385 (N_6385,N_5693,N_5746);
nor U6386 (N_6386,N_5363,N_5873);
xnor U6387 (N_6387,N_5670,N_5606);
and U6388 (N_6388,N_5318,N_5447);
xnor U6389 (N_6389,N_5929,N_5765);
or U6390 (N_6390,N_5743,N_5951);
nand U6391 (N_6391,N_5633,N_5626);
or U6392 (N_6392,N_5378,N_5896);
xnor U6393 (N_6393,N_5897,N_5384);
or U6394 (N_6394,N_5256,N_5866);
xnor U6395 (N_6395,N_5926,N_5382);
nand U6396 (N_6396,N_5742,N_5373);
or U6397 (N_6397,N_5427,N_5326);
xnor U6398 (N_6398,N_5587,N_5499);
nand U6399 (N_6399,N_5371,N_5848);
or U6400 (N_6400,N_5384,N_5577);
and U6401 (N_6401,N_5765,N_5803);
nand U6402 (N_6402,N_5519,N_5496);
and U6403 (N_6403,N_5623,N_5955);
and U6404 (N_6404,N_5689,N_5290);
nor U6405 (N_6405,N_5468,N_5467);
nor U6406 (N_6406,N_5347,N_5609);
or U6407 (N_6407,N_5533,N_5974);
or U6408 (N_6408,N_5490,N_5286);
nand U6409 (N_6409,N_5641,N_5908);
xnor U6410 (N_6410,N_5827,N_5513);
nor U6411 (N_6411,N_5360,N_5531);
and U6412 (N_6412,N_5371,N_5565);
or U6413 (N_6413,N_5513,N_5379);
xor U6414 (N_6414,N_5680,N_5327);
or U6415 (N_6415,N_5864,N_5915);
nor U6416 (N_6416,N_5458,N_5937);
nand U6417 (N_6417,N_5739,N_5823);
xnor U6418 (N_6418,N_5847,N_5781);
xor U6419 (N_6419,N_5416,N_5970);
xnor U6420 (N_6420,N_5967,N_5356);
or U6421 (N_6421,N_5682,N_5931);
xor U6422 (N_6422,N_5904,N_5863);
and U6423 (N_6423,N_5640,N_5338);
and U6424 (N_6424,N_5625,N_5474);
or U6425 (N_6425,N_5257,N_5568);
or U6426 (N_6426,N_5585,N_5522);
or U6427 (N_6427,N_5774,N_5457);
nor U6428 (N_6428,N_5592,N_5553);
and U6429 (N_6429,N_5395,N_5711);
nand U6430 (N_6430,N_5962,N_5851);
and U6431 (N_6431,N_5572,N_5798);
nor U6432 (N_6432,N_5348,N_5792);
xor U6433 (N_6433,N_5772,N_5480);
xor U6434 (N_6434,N_5326,N_5387);
or U6435 (N_6435,N_5386,N_5508);
nor U6436 (N_6436,N_5436,N_5652);
or U6437 (N_6437,N_5301,N_5557);
xor U6438 (N_6438,N_5457,N_5571);
nor U6439 (N_6439,N_5303,N_5744);
or U6440 (N_6440,N_5461,N_5768);
and U6441 (N_6441,N_5351,N_5650);
nand U6442 (N_6442,N_5476,N_5799);
nand U6443 (N_6443,N_5863,N_5859);
and U6444 (N_6444,N_5561,N_5703);
and U6445 (N_6445,N_5890,N_5687);
or U6446 (N_6446,N_5554,N_5589);
xnor U6447 (N_6447,N_5907,N_5295);
nor U6448 (N_6448,N_5519,N_5648);
xnor U6449 (N_6449,N_5941,N_5343);
xor U6450 (N_6450,N_5344,N_5618);
and U6451 (N_6451,N_5597,N_5679);
xnor U6452 (N_6452,N_5510,N_5953);
xnor U6453 (N_6453,N_5478,N_5754);
xor U6454 (N_6454,N_5897,N_5479);
xnor U6455 (N_6455,N_5279,N_5270);
or U6456 (N_6456,N_5525,N_5631);
or U6457 (N_6457,N_5402,N_5688);
nand U6458 (N_6458,N_5907,N_5474);
or U6459 (N_6459,N_5405,N_5388);
nor U6460 (N_6460,N_5536,N_5968);
or U6461 (N_6461,N_5321,N_5959);
nand U6462 (N_6462,N_5339,N_5773);
and U6463 (N_6463,N_5494,N_5292);
and U6464 (N_6464,N_5565,N_5796);
nor U6465 (N_6465,N_5546,N_5900);
or U6466 (N_6466,N_5996,N_5310);
and U6467 (N_6467,N_5906,N_5278);
nand U6468 (N_6468,N_5649,N_5807);
xnor U6469 (N_6469,N_5370,N_5282);
xor U6470 (N_6470,N_5702,N_5577);
xor U6471 (N_6471,N_5684,N_5611);
nand U6472 (N_6472,N_5758,N_5490);
xnor U6473 (N_6473,N_5449,N_5675);
and U6474 (N_6474,N_5566,N_5356);
and U6475 (N_6475,N_5262,N_5371);
or U6476 (N_6476,N_5374,N_5535);
and U6477 (N_6477,N_5525,N_5355);
or U6478 (N_6478,N_5735,N_5860);
xnor U6479 (N_6479,N_5707,N_5691);
nand U6480 (N_6480,N_5301,N_5713);
nand U6481 (N_6481,N_5516,N_5954);
and U6482 (N_6482,N_5313,N_5275);
and U6483 (N_6483,N_5374,N_5434);
or U6484 (N_6484,N_5337,N_5975);
xor U6485 (N_6485,N_5520,N_5747);
nor U6486 (N_6486,N_5339,N_5962);
and U6487 (N_6487,N_5786,N_5969);
nand U6488 (N_6488,N_5909,N_5305);
nand U6489 (N_6489,N_5624,N_5616);
or U6490 (N_6490,N_5575,N_5961);
nor U6491 (N_6491,N_5620,N_5428);
or U6492 (N_6492,N_5399,N_5577);
or U6493 (N_6493,N_5361,N_5393);
nand U6494 (N_6494,N_5476,N_5471);
nand U6495 (N_6495,N_5924,N_5370);
xnor U6496 (N_6496,N_5462,N_5875);
nor U6497 (N_6497,N_5823,N_5824);
xnor U6498 (N_6498,N_5846,N_5820);
nand U6499 (N_6499,N_5819,N_5888);
nor U6500 (N_6500,N_5531,N_5426);
and U6501 (N_6501,N_5788,N_5659);
nor U6502 (N_6502,N_5562,N_5777);
nor U6503 (N_6503,N_5639,N_5636);
nand U6504 (N_6504,N_5339,N_5348);
nand U6505 (N_6505,N_5569,N_5549);
and U6506 (N_6506,N_5774,N_5761);
xnor U6507 (N_6507,N_5685,N_5572);
and U6508 (N_6508,N_5401,N_5907);
or U6509 (N_6509,N_5874,N_5801);
and U6510 (N_6510,N_5479,N_5644);
and U6511 (N_6511,N_5457,N_5821);
and U6512 (N_6512,N_5323,N_5409);
nor U6513 (N_6513,N_5256,N_5457);
nor U6514 (N_6514,N_5526,N_5937);
nand U6515 (N_6515,N_5640,N_5675);
xor U6516 (N_6516,N_5700,N_5317);
nand U6517 (N_6517,N_5483,N_5279);
nand U6518 (N_6518,N_5402,N_5532);
nor U6519 (N_6519,N_5515,N_5739);
nor U6520 (N_6520,N_5535,N_5526);
or U6521 (N_6521,N_5846,N_5968);
nor U6522 (N_6522,N_5931,N_5965);
nand U6523 (N_6523,N_5360,N_5999);
nor U6524 (N_6524,N_5930,N_5982);
nor U6525 (N_6525,N_5807,N_5946);
and U6526 (N_6526,N_5493,N_5907);
xnor U6527 (N_6527,N_5911,N_5335);
nor U6528 (N_6528,N_5295,N_5706);
and U6529 (N_6529,N_5645,N_5778);
nand U6530 (N_6530,N_5612,N_5786);
nand U6531 (N_6531,N_5953,N_5530);
nand U6532 (N_6532,N_5411,N_5904);
nand U6533 (N_6533,N_5487,N_5364);
and U6534 (N_6534,N_5893,N_5716);
nand U6535 (N_6535,N_5901,N_5689);
xnor U6536 (N_6536,N_5898,N_5597);
nor U6537 (N_6537,N_5393,N_5941);
or U6538 (N_6538,N_5949,N_5562);
and U6539 (N_6539,N_5908,N_5735);
or U6540 (N_6540,N_5845,N_5450);
or U6541 (N_6541,N_5591,N_5690);
nor U6542 (N_6542,N_5867,N_5704);
xnor U6543 (N_6543,N_5677,N_5259);
and U6544 (N_6544,N_5750,N_5653);
or U6545 (N_6545,N_5269,N_5653);
nor U6546 (N_6546,N_5674,N_5454);
nand U6547 (N_6547,N_5419,N_5891);
nor U6548 (N_6548,N_5498,N_5630);
nand U6549 (N_6549,N_5386,N_5345);
xnor U6550 (N_6550,N_5307,N_5990);
or U6551 (N_6551,N_5399,N_5827);
or U6552 (N_6552,N_5401,N_5676);
or U6553 (N_6553,N_5714,N_5877);
and U6554 (N_6554,N_5656,N_5256);
nand U6555 (N_6555,N_5789,N_5950);
and U6556 (N_6556,N_5562,N_5288);
or U6557 (N_6557,N_5382,N_5579);
and U6558 (N_6558,N_5305,N_5631);
xor U6559 (N_6559,N_5713,N_5490);
and U6560 (N_6560,N_5483,N_5983);
and U6561 (N_6561,N_5502,N_5600);
xnor U6562 (N_6562,N_5694,N_5751);
and U6563 (N_6563,N_5840,N_5301);
xor U6564 (N_6564,N_5722,N_5401);
nand U6565 (N_6565,N_5689,N_5357);
nand U6566 (N_6566,N_5700,N_5486);
xor U6567 (N_6567,N_5533,N_5724);
nand U6568 (N_6568,N_5871,N_5605);
nand U6569 (N_6569,N_5361,N_5993);
or U6570 (N_6570,N_5476,N_5732);
xnor U6571 (N_6571,N_5669,N_5655);
and U6572 (N_6572,N_5459,N_5529);
xor U6573 (N_6573,N_5710,N_5857);
and U6574 (N_6574,N_5897,N_5589);
xnor U6575 (N_6575,N_5989,N_5609);
and U6576 (N_6576,N_5535,N_5417);
nor U6577 (N_6577,N_5863,N_5896);
and U6578 (N_6578,N_5484,N_5497);
nand U6579 (N_6579,N_5964,N_5454);
nand U6580 (N_6580,N_5840,N_5395);
nand U6581 (N_6581,N_5824,N_5947);
nand U6582 (N_6582,N_5831,N_5488);
nor U6583 (N_6583,N_5686,N_5297);
or U6584 (N_6584,N_5881,N_5793);
and U6585 (N_6585,N_5985,N_5437);
nand U6586 (N_6586,N_5889,N_5577);
xnor U6587 (N_6587,N_5552,N_5506);
nand U6588 (N_6588,N_5409,N_5501);
nor U6589 (N_6589,N_5506,N_5936);
nand U6590 (N_6590,N_5672,N_5256);
and U6591 (N_6591,N_5727,N_5580);
xor U6592 (N_6592,N_5973,N_5459);
and U6593 (N_6593,N_5487,N_5976);
and U6594 (N_6594,N_5528,N_5858);
nand U6595 (N_6595,N_5988,N_5616);
nand U6596 (N_6596,N_5738,N_5928);
xnor U6597 (N_6597,N_5468,N_5642);
nand U6598 (N_6598,N_5273,N_5684);
xnor U6599 (N_6599,N_5396,N_5694);
xnor U6600 (N_6600,N_5656,N_5977);
nand U6601 (N_6601,N_5600,N_5554);
nor U6602 (N_6602,N_5326,N_5845);
xor U6603 (N_6603,N_5259,N_5842);
nor U6604 (N_6604,N_5982,N_5691);
xor U6605 (N_6605,N_5545,N_5955);
xnor U6606 (N_6606,N_5351,N_5567);
xor U6607 (N_6607,N_5490,N_5834);
nand U6608 (N_6608,N_5449,N_5628);
nand U6609 (N_6609,N_5417,N_5734);
and U6610 (N_6610,N_5560,N_5843);
nor U6611 (N_6611,N_5664,N_5303);
nor U6612 (N_6612,N_5433,N_5642);
xor U6613 (N_6613,N_5377,N_5333);
xnor U6614 (N_6614,N_5786,N_5437);
nor U6615 (N_6615,N_5565,N_5403);
nand U6616 (N_6616,N_5707,N_5702);
and U6617 (N_6617,N_5969,N_5991);
nand U6618 (N_6618,N_5927,N_5298);
xnor U6619 (N_6619,N_5608,N_5705);
or U6620 (N_6620,N_5285,N_5491);
xnor U6621 (N_6621,N_5984,N_5945);
nand U6622 (N_6622,N_5591,N_5398);
and U6623 (N_6623,N_5639,N_5478);
and U6624 (N_6624,N_5623,N_5793);
nand U6625 (N_6625,N_5311,N_5906);
nor U6626 (N_6626,N_5333,N_5308);
nor U6627 (N_6627,N_5253,N_5791);
nand U6628 (N_6628,N_5472,N_5832);
nor U6629 (N_6629,N_5752,N_5993);
and U6630 (N_6630,N_5813,N_5741);
or U6631 (N_6631,N_5983,N_5557);
nor U6632 (N_6632,N_5284,N_5715);
and U6633 (N_6633,N_5342,N_5298);
nand U6634 (N_6634,N_5691,N_5708);
xor U6635 (N_6635,N_5423,N_5504);
or U6636 (N_6636,N_5927,N_5563);
and U6637 (N_6637,N_5884,N_5317);
or U6638 (N_6638,N_5258,N_5329);
or U6639 (N_6639,N_5880,N_5705);
xnor U6640 (N_6640,N_5689,N_5630);
xnor U6641 (N_6641,N_5628,N_5992);
xor U6642 (N_6642,N_5693,N_5268);
nand U6643 (N_6643,N_5250,N_5936);
or U6644 (N_6644,N_5954,N_5764);
or U6645 (N_6645,N_5938,N_5498);
or U6646 (N_6646,N_5370,N_5733);
nor U6647 (N_6647,N_5557,N_5978);
and U6648 (N_6648,N_5816,N_5762);
nor U6649 (N_6649,N_5434,N_5428);
and U6650 (N_6650,N_5595,N_5342);
and U6651 (N_6651,N_5354,N_5814);
xnor U6652 (N_6652,N_5286,N_5416);
and U6653 (N_6653,N_5643,N_5752);
and U6654 (N_6654,N_5302,N_5412);
or U6655 (N_6655,N_5292,N_5769);
xnor U6656 (N_6656,N_5285,N_5566);
nor U6657 (N_6657,N_5769,N_5487);
nor U6658 (N_6658,N_5253,N_5696);
nand U6659 (N_6659,N_5670,N_5413);
or U6660 (N_6660,N_5373,N_5968);
or U6661 (N_6661,N_5821,N_5643);
and U6662 (N_6662,N_5907,N_5965);
nand U6663 (N_6663,N_5545,N_5663);
nand U6664 (N_6664,N_5356,N_5789);
nand U6665 (N_6665,N_5939,N_5688);
xnor U6666 (N_6666,N_5300,N_5396);
nor U6667 (N_6667,N_5517,N_5975);
or U6668 (N_6668,N_5902,N_5605);
xnor U6669 (N_6669,N_5956,N_5823);
and U6670 (N_6670,N_5255,N_5615);
or U6671 (N_6671,N_5780,N_5692);
nor U6672 (N_6672,N_5798,N_5549);
or U6673 (N_6673,N_5550,N_5292);
nor U6674 (N_6674,N_5793,N_5688);
nor U6675 (N_6675,N_5544,N_5472);
nor U6676 (N_6676,N_5265,N_5282);
or U6677 (N_6677,N_5290,N_5288);
and U6678 (N_6678,N_5316,N_5823);
nor U6679 (N_6679,N_5895,N_5715);
xnor U6680 (N_6680,N_5784,N_5945);
nand U6681 (N_6681,N_5280,N_5764);
nand U6682 (N_6682,N_5960,N_5920);
or U6683 (N_6683,N_5712,N_5708);
and U6684 (N_6684,N_5378,N_5443);
nor U6685 (N_6685,N_5654,N_5611);
nand U6686 (N_6686,N_5303,N_5632);
and U6687 (N_6687,N_5889,N_5996);
xnor U6688 (N_6688,N_5425,N_5345);
and U6689 (N_6689,N_5606,N_5406);
and U6690 (N_6690,N_5860,N_5267);
xnor U6691 (N_6691,N_5547,N_5413);
nand U6692 (N_6692,N_5655,N_5664);
xnor U6693 (N_6693,N_5677,N_5566);
or U6694 (N_6694,N_5722,N_5528);
nand U6695 (N_6695,N_5391,N_5406);
or U6696 (N_6696,N_5691,N_5960);
xnor U6697 (N_6697,N_5672,N_5268);
nand U6698 (N_6698,N_5360,N_5930);
xnor U6699 (N_6699,N_5261,N_5759);
or U6700 (N_6700,N_5927,N_5953);
xor U6701 (N_6701,N_5816,N_5655);
or U6702 (N_6702,N_5286,N_5652);
or U6703 (N_6703,N_5665,N_5702);
or U6704 (N_6704,N_5786,N_5522);
and U6705 (N_6705,N_5776,N_5753);
xnor U6706 (N_6706,N_5923,N_5297);
nand U6707 (N_6707,N_5450,N_5283);
xnor U6708 (N_6708,N_5764,N_5738);
xor U6709 (N_6709,N_5518,N_5784);
and U6710 (N_6710,N_5276,N_5274);
and U6711 (N_6711,N_5398,N_5982);
xnor U6712 (N_6712,N_5397,N_5294);
or U6713 (N_6713,N_5377,N_5996);
nor U6714 (N_6714,N_5590,N_5259);
xnor U6715 (N_6715,N_5768,N_5577);
nand U6716 (N_6716,N_5833,N_5367);
xor U6717 (N_6717,N_5620,N_5429);
nor U6718 (N_6718,N_5754,N_5385);
nand U6719 (N_6719,N_5342,N_5594);
nand U6720 (N_6720,N_5948,N_5538);
or U6721 (N_6721,N_5620,N_5342);
nor U6722 (N_6722,N_5279,N_5254);
nand U6723 (N_6723,N_5721,N_5360);
or U6724 (N_6724,N_5821,N_5600);
and U6725 (N_6725,N_5793,N_5830);
nand U6726 (N_6726,N_5437,N_5508);
xnor U6727 (N_6727,N_5346,N_5868);
nand U6728 (N_6728,N_5282,N_5315);
nand U6729 (N_6729,N_5546,N_5872);
nand U6730 (N_6730,N_5615,N_5708);
nor U6731 (N_6731,N_5431,N_5955);
nand U6732 (N_6732,N_5948,N_5928);
nand U6733 (N_6733,N_5682,N_5587);
nor U6734 (N_6734,N_5518,N_5938);
or U6735 (N_6735,N_5963,N_5521);
or U6736 (N_6736,N_5936,N_5981);
nand U6737 (N_6737,N_5772,N_5934);
xor U6738 (N_6738,N_5711,N_5345);
xnor U6739 (N_6739,N_5715,N_5385);
and U6740 (N_6740,N_5717,N_5928);
or U6741 (N_6741,N_5314,N_5969);
or U6742 (N_6742,N_5739,N_5337);
or U6743 (N_6743,N_5606,N_5604);
xnor U6744 (N_6744,N_5601,N_5390);
or U6745 (N_6745,N_5947,N_5382);
xnor U6746 (N_6746,N_5873,N_5452);
nor U6747 (N_6747,N_5477,N_5307);
and U6748 (N_6748,N_5405,N_5903);
nand U6749 (N_6749,N_5326,N_5751);
and U6750 (N_6750,N_6033,N_6204);
xor U6751 (N_6751,N_6741,N_6360);
nor U6752 (N_6752,N_6081,N_6497);
or U6753 (N_6753,N_6233,N_6588);
nor U6754 (N_6754,N_6327,N_6594);
or U6755 (N_6755,N_6282,N_6577);
and U6756 (N_6756,N_6552,N_6135);
nand U6757 (N_6757,N_6133,N_6143);
xor U6758 (N_6758,N_6507,N_6523);
nand U6759 (N_6759,N_6578,N_6165);
and U6760 (N_6760,N_6568,N_6573);
and U6761 (N_6761,N_6628,N_6627);
nor U6762 (N_6762,N_6046,N_6583);
or U6763 (N_6763,N_6698,N_6351);
or U6764 (N_6764,N_6283,N_6430);
or U6765 (N_6765,N_6374,N_6011);
or U6766 (N_6766,N_6224,N_6186);
and U6767 (N_6767,N_6012,N_6307);
or U6768 (N_6768,N_6525,N_6227);
nor U6769 (N_6769,N_6083,N_6301);
nor U6770 (N_6770,N_6671,N_6348);
or U6771 (N_6771,N_6736,N_6484);
nor U6772 (N_6772,N_6388,N_6181);
and U6773 (N_6773,N_6488,N_6633);
and U6774 (N_6774,N_6674,N_6246);
and U6775 (N_6775,N_6547,N_6250);
xnor U6776 (N_6776,N_6061,N_6020);
or U6777 (N_6777,N_6337,N_6220);
xnor U6778 (N_6778,N_6563,N_6343);
and U6779 (N_6779,N_6159,N_6713);
xor U6780 (N_6780,N_6689,N_6412);
nor U6781 (N_6781,N_6666,N_6206);
or U6782 (N_6782,N_6120,N_6403);
nand U6783 (N_6783,N_6253,N_6269);
nor U6784 (N_6784,N_6209,N_6592);
or U6785 (N_6785,N_6580,N_6310);
and U6786 (N_6786,N_6526,N_6570);
or U6787 (N_6787,N_6333,N_6676);
and U6788 (N_6788,N_6432,N_6656);
and U6789 (N_6789,N_6069,N_6571);
xnor U6790 (N_6790,N_6080,N_6223);
and U6791 (N_6791,N_6396,N_6687);
xnor U6792 (N_6792,N_6553,N_6114);
or U6793 (N_6793,N_6302,N_6158);
nand U6794 (N_6794,N_6336,N_6625);
xnor U6795 (N_6795,N_6144,N_6411);
nand U6796 (N_6796,N_6029,N_6028);
and U6797 (N_6797,N_6052,N_6314);
and U6798 (N_6798,N_6362,N_6106);
xor U6799 (N_6799,N_6677,N_6470);
xor U6800 (N_6800,N_6101,N_6476);
nand U6801 (N_6801,N_6541,N_6501);
nand U6802 (N_6802,N_6426,N_6668);
nand U6803 (N_6803,N_6557,N_6460);
xor U6804 (N_6804,N_6611,N_6010);
and U6805 (N_6805,N_6654,N_6174);
nor U6806 (N_6806,N_6705,N_6319);
nor U6807 (N_6807,N_6700,N_6718);
nand U6808 (N_6808,N_6221,N_6520);
nand U6809 (N_6809,N_6024,N_6236);
nor U6810 (N_6810,N_6112,N_6254);
and U6811 (N_6811,N_6167,N_6602);
xor U6812 (N_6812,N_6299,N_6612);
or U6813 (N_6813,N_6038,N_6717);
nor U6814 (N_6814,N_6405,N_6096);
xor U6815 (N_6815,N_6156,N_6322);
and U6816 (N_6816,N_6703,N_6740);
nor U6817 (N_6817,N_6304,N_6289);
nor U6818 (N_6818,N_6421,N_6309);
nor U6819 (N_6819,N_6228,N_6320);
or U6820 (N_6820,N_6329,N_6495);
nor U6821 (N_6821,N_6267,N_6660);
nor U6822 (N_6822,N_6379,N_6161);
nor U6823 (N_6823,N_6118,N_6205);
xor U6824 (N_6824,N_6519,N_6479);
and U6825 (N_6825,N_6431,N_6615);
nand U6826 (N_6826,N_6657,N_6414);
or U6827 (N_6827,N_6672,N_6330);
xor U6828 (N_6828,N_6555,N_6147);
nor U6829 (N_6829,N_6384,N_6017);
nor U6830 (N_6830,N_6528,N_6030);
and U6831 (N_6831,N_6239,N_6579);
xnor U6832 (N_6832,N_6480,N_6638);
or U6833 (N_6833,N_6266,N_6324);
nand U6834 (N_6834,N_6212,N_6632);
xnor U6835 (N_6835,N_6550,N_6447);
or U6836 (N_6836,N_6249,N_6107);
nand U6837 (N_6837,N_6524,N_6164);
xnor U6838 (N_6838,N_6295,N_6462);
nand U6839 (N_6839,N_6076,N_6214);
and U6840 (N_6840,N_6188,N_6591);
nor U6841 (N_6841,N_6091,N_6271);
nor U6842 (N_6842,N_6037,N_6564);
nor U6843 (N_6843,N_6211,N_6108);
xnor U6844 (N_6844,N_6345,N_6688);
nor U6845 (N_6845,N_6665,N_6323);
xor U6846 (N_6846,N_6739,N_6045);
or U6847 (N_6847,N_6260,N_6609);
nor U6848 (N_6848,N_6637,N_6247);
xnor U6849 (N_6849,N_6117,N_6123);
or U6850 (N_6850,N_6461,N_6465);
nand U6851 (N_6851,N_6210,N_6180);
or U6852 (N_6852,N_6605,N_6272);
nor U6853 (N_6853,N_6022,N_6498);
and U6854 (N_6854,N_6134,N_6601);
nand U6855 (N_6855,N_6261,N_6697);
nand U6856 (N_6856,N_6268,N_6086);
nand U6857 (N_6857,N_6715,N_6357);
nor U6858 (N_6858,N_6537,N_6503);
nor U6859 (N_6859,N_6349,N_6724);
nand U6860 (N_6860,N_6401,N_6599);
xnor U6861 (N_6861,N_6130,N_6621);
xor U6862 (N_6862,N_6725,N_6089);
nand U6863 (N_6863,N_6187,N_6155);
nor U6864 (N_6864,N_6222,N_6315);
xnor U6865 (N_6865,N_6006,N_6531);
xnor U6866 (N_6866,N_6148,N_6366);
or U6867 (N_6867,N_6063,N_6370);
xor U6868 (N_6868,N_6039,N_6265);
and U6869 (N_6869,N_6226,N_6367);
xnor U6870 (N_6870,N_6604,N_6482);
nor U6871 (N_6871,N_6191,N_6023);
and U6872 (N_6872,N_6291,N_6473);
or U6873 (N_6873,N_6506,N_6397);
and U6874 (N_6874,N_6567,N_6516);
xor U6875 (N_6875,N_6726,N_6417);
nand U6876 (N_6876,N_6097,N_6297);
and U6877 (N_6877,N_6256,N_6074);
nor U6878 (N_6878,N_6732,N_6551);
nor U6879 (N_6879,N_6669,N_6483);
nand U6880 (N_6880,N_6047,N_6170);
and U6881 (N_6881,N_6049,N_6326);
or U6882 (N_6882,N_6748,N_6733);
xnor U6883 (N_6883,N_6245,N_6098);
nor U6884 (N_6884,N_6105,N_6548);
and U6885 (N_6885,N_6636,N_6229);
nand U6886 (N_6886,N_6590,N_6041);
nand U6887 (N_6887,N_6400,N_6198);
nor U6888 (N_6888,N_6318,N_6175);
nor U6889 (N_6889,N_6054,N_6438);
xor U6890 (N_6890,N_6415,N_6312);
and U6891 (N_6891,N_6189,N_6296);
xnor U6892 (N_6892,N_6257,N_6734);
or U6893 (N_6893,N_6721,N_6331);
or U6894 (N_6894,N_6190,N_6132);
nand U6895 (N_6895,N_6216,N_6100);
nor U6896 (N_6896,N_6486,N_6514);
nand U6897 (N_6897,N_6368,N_6196);
or U6898 (N_6898,N_6509,N_6584);
xor U6899 (N_6899,N_6539,N_6162);
or U6900 (N_6900,N_6452,N_6694);
nand U6901 (N_6901,N_6399,N_6183);
xnor U6902 (N_6902,N_6662,N_6650);
nand U6903 (N_6903,N_6026,N_6693);
nand U6904 (N_6904,N_6682,N_6154);
xnor U6905 (N_6905,N_6463,N_6353);
or U6906 (N_6906,N_6419,N_6667);
and U6907 (N_6907,N_6424,N_6225);
or U6908 (N_6908,N_6018,N_6735);
nand U6909 (N_6909,N_6150,N_6512);
and U6910 (N_6910,N_6115,N_6679);
nor U6911 (N_6911,N_6502,N_6001);
or U6912 (N_6912,N_6325,N_6293);
or U6913 (N_6913,N_6466,N_6004);
xor U6914 (N_6914,N_6496,N_6352);
xnor U6915 (N_6915,N_6005,N_6369);
or U6916 (N_6916,N_6661,N_6371);
nand U6917 (N_6917,N_6651,N_6394);
nand U6918 (N_6918,N_6193,N_6334);
xnor U6919 (N_6919,N_6533,N_6566);
and U6920 (N_6920,N_6746,N_6275);
nor U6921 (N_6921,N_6398,N_6378);
and U6922 (N_6922,N_6203,N_6276);
and U6923 (N_6923,N_6428,N_6259);
or U6924 (N_6924,N_6375,N_6317);
nor U6925 (N_6925,N_6744,N_6243);
nor U6926 (N_6926,N_6104,N_6613);
and U6927 (N_6927,N_6407,N_6234);
and U6928 (N_6928,N_6082,N_6122);
nor U6929 (N_6929,N_6521,N_6681);
and U6930 (N_6930,N_6121,N_6136);
and U6931 (N_6931,N_6192,N_6389);
nand U6932 (N_6932,N_6051,N_6199);
and U6933 (N_6933,N_6042,N_6610);
nor U6934 (N_6934,N_6534,N_6308);
nand U6935 (N_6935,N_6451,N_6284);
xor U6936 (N_6936,N_6708,N_6749);
or U6937 (N_6937,N_6562,N_6386);
and U6938 (N_6938,N_6459,N_6328);
and U6939 (N_6939,N_6034,N_6013);
xor U6940 (N_6940,N_6278,N_6608);
nor U6941 (N_6941,N_6499,N_6738);
or U6942 (N_6942,N_6119,N_6021);
or U6943 (N_6943,N_6434,N_6171);
or U6944 (N_6944,N_6678,N_6339);
or U6945 (N_6945,N_6274,N_6664);
and U6946 (N_6946,N_6290,N_6113);
nand U6947 (N_6947,N_6099,N_6730);
nand U6948 (N_6948,N_6532,N_6712);
nand U6949 (N_6949,N_6313,N_6728);
xor U6950 (N_6950,N_6606,N_6600);
nor U6951 (N_6951,N_6742,N_6648);
xnor U6952 (N_6952,N_6559,N_6391);
and U6953 (N_6953,N_6517,N_6383);
nor U6954 (N_6954,N_6691,N_6543);
nor U6955 (N_6955,N_6218,N_6574);
xnor U6956 (N_6956,N_6634,N_6084);
nor U6957 (N_6957,N_6458,N_6425);
xnor U6958 (N_6958,N_6050,N_6003);
or U6959 (N_6959,N_6178,N_6129);
nand U6960 (N_6960,N_6572,N_6059);
nor U6961 (N_6961,N_6544,N_6607);
nor U6962 (N_6962,N_6535,N_6586);
and U6963 (N_6963,N_6335,N_6485);
nor U6964 (N_6964,N_6545,N_6409);
nand U6965 (N_6965,N_6103,N_6067);
nor U6966 (N_6966,N_6064,N_6440);
xnor U6967 (N_6967,N_6685,N_6653);
xor U6968 (N_6968,N_6072,N_6596);
nor U6969 (N_6969,N_6701,N_6027);
xor U6970 (N_6970,N_6629,N_6217);
nor U6971 (N_6971,N_6663,N_6439);
nor U6972 (N_6972,N_6722,N_6561);
and U6973 (N_6973,N_6087,N_6350);
and U6974 (N_6974,N_6518,N_6303);
nor U6975 (N_6975,N_6589,N_6088);
nand U6976 (N_6976,N_6527,N_6151);
nand U6977 (N_6977,N_6316,N_6009);
xnor U6978 (N_6978,N_6464,N_6508);
nor U6979 (N_6979,N_6670,N_6455);
nor U6980 (N_6980,N_6540,N_6195);
and U6981 (N_6981,N_6255,N_6699);
xnor U6982 (N_6982,N_6095,N_6575);
and U6983 (N_6983,N_6109,N_6442);
or U6984 (N_6984,N_6347,N_6515);
xor U6985 (N_6985,N_6373,N_6235);
xnor U6986 (N_6986,N_6232,N_6264);
xor U6987 (N_6987,N_6281,N_6385);
xnor U6988 (N_6988,N_6043,N_6053);
nand U6989 (N_6989,N_6185,N_6182);
and U6990 (N_6990,N_6704,N_6258);
or U6991 (N_6991,N_6655,N_6449);
or U6992 (N_6992,N_6731,N_6696);
nand U6993 (N_6993,N_6215,N_6102);
or U6994 (N_6994,N_6393,N_6491);
nor U6995 (N_6995,N_6342,N_6230);
nor U6996 (N_6996,N_6437,N_6416);
and U6997 (N_6997,N_6603,N_6380);
or U6998 (N_6998,N_6622,N_6179);
nand U6999 (N_6999,N_6131,N_6341);
or U7000 (N_7000,N_6617,N_6549);
and U7001 (N_7001,N_6585,N_6321);
nand U7002 (N_7002,N_6619,N_6381);
xor U7003 (N_7003,N_6436,N_6450);
xnor U7004 (N_7004,N_6172,N_6090);
nand U7005 (N_7005,N_6593,N_6408);
xnor U7006 (N_7006,N_6435,N_6273);
and U7007 (N_7007,N_6639,N_6598);
nand U7008 (N_7008,N_6361,N_6472);
xor U7009 (N_7009,N_6073,N_6176);
nor U7010 (N_7010,N_6116,N_6040);
nor U7011 (N_7011,N_6390,N_6433);
or U7012 (N_7012,N_6298,N_6300);
xnor U7013 (N_7013,N_6536,N_6032);
and U7014 (N_7014,N_6202,N_6737);
xor U7015 (N_7015,N_6420,N_6031);
nand U7016 (N_7016,N_6075,N_6522);
nor U7017 (N_7017,N_6716,N_6560);
xor U7018 (N_7018,N_6538,N_6631);
nor U7019 (N_7019,N_6492,N_6644);
nor U7020 (N_7020,N_6443,N_6475);
and U7021 (N_7021,N_6048,N_6680);
xnor U7022 (N_7022,N_6556,N_6340);
nand U7023 (N_7023,N_6727,N_6248);
and U7024 (N_7024,N_6646,N_6242);
xnor U7025 (N_7025,N_6138,N_6569);
nand U7026 (N_7026,N_6616,N_6423);
nand U7027 (N_7027,N_6019,N_6481);
xnor U7028 (N_7028,N_6197,N_6618);
nand U7029 (N_7029,N_6092,N_6626);
or U7030 (N_7030,N_6173,N_6231);
nor U7031 (N_7031,N_6055,N_6279);
or U7032 (N_7032,N_6530,N_6376);
nand U7033 (N_7033,N_6025,N_6576);
nand U7034 (N_7034,N_6344,N_6490);
xnor U7035 (N_7035,N_6690,N_6141);
and U7036 (N_7036,N_6529,N_6079);
nor U7037 (N_7037,N_6007,N_6270);
and U7038 (N_7038,N_6015,N_6285);
xnor U7039 (N_7039,N_6542,N_6002);
and U7040 (N_7040,N_6062,N_6377);
xnor U7041 (N_7041,N_6057,N_6044);
nor U7042 (N_7042,N_6474,N_6262);
and U7043 (N_7043,N_6630,N_6510);
xor U7044 (N_7044,N_6453,N_6673);
nand U7045 (N_7045,N_6658,N_6714);
nor U7046 (N_7046,N_6355,N_6358);
nand U7047 (N_7047,N_6127,N_6635);
xor U7048 (N_7048,N_6213,N_6160);
or U7049 (N_7049,N_6710,N_6058);
nor U7050 (N_7050,N_6645,N_6406);
nor U7051 (N_7051,N_6194,N_6707);
and U7052 (N_7052,N_6140,N_6467);
and U7053 (N_7053,N_6036,N_6207);
or U7054 (N_7054,N_6237,N_6153);
or U7055 (N_7055,N_6695,N_6382);
and U7056 (N_7056,N_6184,N_6149);
nor U7057 (N_7057,N_6111,N_6200);
nor U7058 (N_7058,N_6241,N_6146);
nor U7059 (N_7059,N_6354,N_6070);
nand U7060 (N_7060,N_6640,N_6392);
nand U7061 (N_7061,N_6166,N_6287);
xor U7062 (N_7062,N_6706,N_6614);
nor U7063 (N_7063,N_6469,N_6649);
or U7064 (N_7064,N_6471,N_6652);
nand U7065 (N_7065,N_6332,N_6277);
nand U7066 (N_7066,N_6445,N_6000);
xnor U7067 (N_7067,N_6565,N_6511);
or U7068 (N_7068,N_6346,N_6647);
xnor U7069 (N_7069,N_6035,N_6587);
xnor U7070 (N_7070,N_6643,N_6554);
nand U7071 (N_7071,N_6338,N_6624);
xnor U7072 (N_7072,N_6477,N_6395);
or U7073 (N_7073,N_6238,N_6126);
and U7074 (N_7074,N_6404,N_6094);
nor U7075 (N_7075,N_6723,N_6177);
xor U7076 (N_7076,N_6169,N_6219);
and U7077 (N_7077,N_6078,N_6142);
and U7078 (N_7078,N_6145,N_6065);
nor U7079 (N_7079,N_6071,N_6675);
and U7080 (N_7080,N_6014,N_6720);
or U7081 (N_7081,N_6429,N_6427);
nand U7082 (N_7082,N_6157,N_6641);
xor U7083 (N_7083,N_6139,N_6729);
nor U7084 (N_7084,N_6124,N_6686);
or U7085 (N_7085,N_6364,N_6168);
or U7086 (N_7086,N_6110,N_6008);
xor U7087 (N_7087,N_6252,N_6068);
nand U7088 (N_7088,N_6504,N_6747);
nand U7089 (N_7089,N_6201,N_6642);
and U7090 (N_7090,N_6077,N_6413);
and U7091 (N_7091,N_6365,N_6546);
and U7092 (N_7092,N_6582,N_6448);
nor U7093 (N_7093,N_6623,N_6500);
or U7094 (N_7094,N_6240,N_6288);
nand U7095 (N_7095,N_6422,N_6137);
xor U7096 (N_7096,N_6311,N_6745);
or U7097 (N_7097,N_6581,N_6410);
nor U7098 (N_7098,N_6306,N_6387);
nor U7099 (N_7099,N_6294,N_6597);
xor U7100 (N_7100,N_6494,N_6093);
or U7101 (N_7101,N_6478,N_6684);
or U7102 (N_7102,N_6163,N_6456);
or U7103 (N_7103,N_6066,N_6719);
or U7104 (N_7104,N_6595,N_6292);
xnor U7105 (N_7105,N_6244,N_6468);
and U7106 (N_7106,N_6711,N_6558);
and U7107 (N_7107,N_6152,N_6444);
nand U7108 (N_7108,N_6208,N_6446);
and U7109 (N_7109,N_6251,N_6493);
or U7110 (N_7110,N_6709,N_6056);
nand U7111 (N_7111,N_6743,N_6280);
nor U7112 (N_7112,N_6085,N_6402);
nor U7113 (N_7113,N_6305,N_6441);
nand U7114 (N_7114,N_6620,N_6692);
xnor U7115 (N_7115,N_6457,N_6016);
nor U7116 (N_7116,N_6487,N_6659);
or U7117 (N_7117,N_6683,N_6418);
nand U7118 (N_7118,N_6372,N_6060);
nand U7119 (N_7119,N_6356,N_6359);
and U7120 (N_7120,N_6454,N_6263);
nor U7121 (N_7121,N_6128,N_6489);
nand U7122 (N_7122,N_6125,N_6513);
nand U7123 (N_7123,N_6505,N_6702);
xnor U7124 (N_7124,N_6363,N_6286);
and U7125 (N_7125,N_6418,N_6157);
xnor U7126 (N_7126,N_6535,N_6560);
xnor U7127 (N_7127,N_6424,N_6190);
nand U7128 (N_7128,N_6644,N_6035);
nor U7129 (N_7129,N_6682,N_6748);
or U7130 (N_7130,N_6430,N_6725);
or U7131 (N_7131,N_6017,N_6344);
nand U7132 (N_7132,N_6029,N_6574);
nor U7133 (N_7133,N_6390,N_6061);
or U7134 (N_7134,N_6388,N_6409);
xnor U7135 (N_7135,N_6271,N_6175);
xor U7136 (N_7136,N_6423,N_6016);
nand U7137 (N_7137,N_6610,N_6668);
or U7138 (N_7138,N_6502,N_6533);
or U7139 (N_7139,N_6012,N_6058);
xor U7140 (N_7140,N_6100,N_6495);
or U7141 (N_7141,N_6082,N_6126);
nor U7142 (N_7142,N_6128,N_6192);
nor U7143 (N_7143,N_6728,N_6491);
or U7144 (N_7144,N_6403,N_6072);
xor U7145 (N_7145,N_6391,N_6499);
and U7146 (N_7146,N_6228,N_6069);
nand U7147 (N_7147,N_6102,N_6436);
nand U7148 (N_7148,N_6227,N_6455);
nor U7149 (N_7149,N_6097,N_6629);
nor U7150 (N_7150,N_6196,N_6700);
nor U7151 (N_7151,N_6502,N_6144);
nand U7152 (N_7152,N_6531,N_6502);
nand U7153 (N_7153,N_6601,N_6243);
nand U7154 (N_7154,N_6189,N_6254);
nor U7155 (N_7155,N_6669,N_6440);
nand U7156 (N_7156,N_6711,N_6121);
nand U7157 (N_7157,N_6588,N_6256);
nand U7158 (N_7158,N_6603,N_6588);
nand U7159 (N_7159,N_6218,N_6515);
or U7160 (N_7160,N_6184,N_6177);
xor U7161 (N_7161,N_6071,N_6399);
or U7162 (N_7162,N_6609,N_6490);
xnor U7163 (N_7163,N_6002,N_6381);
or U7164 (N_7164,N_6375,N_6458);
and U7165 (N_7165,N_6749,N_6138);
nor U7166 (N_7166,N_6182,N_6156);
nand U7167 (N_7167,N_6736,N_6233);
and U7168 (N_7168,N_6301,N_6244);
nor U7169 (N_7169,N_6015,N_6124);
or U7170 (N_7170,N_6486,N_6185);
or U7171 (N_7171,N_6398,N_6606);
and U7172 (N_7172,N_6275,N_6240);
xnor U7173 (N_7173,N_6287,N_6076);
or U7174 (N_7174,N_6494,N_6440);
and U7175 (N_7175,N_6191,N_6481);
nand U7176 (N_7176,N_6221,N_6656);
or U7177 (N_7177,N_6349,N_6510);
and U7178 (N_7178,N_6088,N_6329);
or U7179 (N_7179,N_6111,N_6739);
xnor U7180 (N_7180,N_6522,N_6438);
nor U7181 (N_7181,N_6459,N_6016);
nor U7182 (N_7182,N_6371,N_6341);
xor U7183 (N_7183,N_6013,N_6746);
nand U7184 (N_7184,N_6044,N_6020);
nor U7185 (N_7185,N_6545,N_6372);
nand U7186 (N_7186,N_6423,N_6058);
nand U7187 (N_7187,N_6570,N_6191);
nand U7188 (N_7188,N_6682,N_6006);
and U7189 (N_7189,N_6289,N_6334);
xnor U7190 (N_7190,N_6373,N_6581);
or U7191 (N_7191,N_6298,N_6000);
nor U7192 (N_7192,N_6567,N_6225);
nor U7193 (N_7193,N_6153,N_6698);
nand U7194 (N_7194,N_6183,N_6259);
and U7195 (N_7195,N_6644,N_6716);
and U7196 (N_7196,N_6617,N_6167);
xnor U7197 (N_7197,N_6701,N_6602);
nor U7198 (N_7198,N_6082,N_6433);
or U7199 (N_7199,N_6268,N_6137);
xnor U7200 (N_7200,N_6607,N_6472);
and U7201 (N_7201,N_6740,N_6064);
or U7202 (N_7202,N_6467,N_6204);
nor U7203 (N_7203,N_6441,N_6531);
and U7204 (N_7204,N_6739,N_6196);
xor U7205 (N_7205,N_6577,N_6251);
nand U7206 (N_7206,N_6069,N_6313);
nand U7207 (N_7207,N_6545,N_6615);
and U7208 (N_7208,N_6592,N_6572);
xnor U7209 (N_7209,N_6288,N_6567);
or U7210 (N_7210,N_6384,N_6642);
xor U7211 (N_7211,N_6139,N_6408);
nor U7212 (N_7212,N_6506,N_6349);
and U7213 (N_7213,N_6300,N_6176);
and U7214 (N_7214,N_6281,N_6058);
nand U7215 (N_7215,N_6155,N_6655);
or U7216 (N_7216,N_6443,N_6686);
or U7217 (N_7217,N_6220,N_6219);
and U7218 (N_7218,N_6674,N_6155);
and U7219 (N_7219,N_6312,N_6215);
or U7220 (N_7220,N_6354,N_6492);
or U7221 (N_7221,N_6564,N_6436);
and U7222 (N_7222,N_6112,N_6446);
and U7223 (N_7223,N_6327,N_6657);
nand U7224 (N_7224,N_6663,N_6065);
xnor U7225 (N_7225,N_6526,N_6357);
or U7226 (N_7226,N_6338,N_6361);
xnor U7227 (N_7227,N_6104,N_6566);
nand U7228 (N_7228,N_6350,N_6501);
nor U7229 (N_7229,N_6543,N_6636);
or U7230 (N_7230,N_6555,N_6016);
xnor U7231 (N_7231,N_6336,N_6026);
nand U7232 (N_7232,N_6182,N_6193);
nand U7233 (N_7233,N_6740,N_6518);
or U7234 (N_7234,N_6590,N_6625);
nand U7235 (N_7235,N_6220,N_6371);
nand U7236 (N_7236,N_6069,N_6214);
or U7237 (N_7237,N_6008,N_6713);
xor U7238 (N_7238,N_6573,N_6530);
xor U7239 (N_7239,N_6171,N_6234);
xor U7240 (N_7240,N_6315,N_6240);
nor U7241 (N_7241,N_6200,N_6623);
and U7242 (N_7242,N_6137,N_6565);
nor U7243 (N_7243,N_6022,N_6415);
or U7244 (N_7244,N_6240,N_6389);
and U7245 (N_7245,N_6371,N_6592);
nor U7246 (N_7246,N_6648,N_6048);
nor U7247 (N_7247,N_6409,N_6642);
nor U7248 (N_7248,N_6292,N_6425);
or U7249 (N_7249,N_6516,N_6049);
and U7250 (N_7250,N_6536,N_6182);
and U7251 (N_7251,N_6147,N_6594);
nor U7252 (N_7252,N_6739,N_6718);
nor U7253 (N_7253,N_6509,N_6438);
nand U7254 (N_7254,N_6126,N_6013);
xnor U7255 (N_7255,N_6622,N_6569);
and U7256 (N_7256,N_6592,N_6506);
xor U7257 (N_7257,N_6075,N_6597);
or U7258 (N_7258,N_6477,N_6670);
and U7259 (N_7259,N_6057,N_6281);
and U7260 (N_7260,N_6691,N_6647);
nor U7261 (N_7261,N_6682,N_6399);
nand U7262 (N_7262,N_6145,N_6147);
nor U7263 (N_7263,N_6013,N_6308);
or U7264 (N_7264,N_6560,N_6414);
xnor U7265 (N_7265,N_6232,N_6013);
and U7266 (N_7266,N_6221,N_6486);
and U7267 (N_7267,N_6191,N_6718);
and U7268 (N_7268,N_6715,N_6280);
xor U7269 (N_7269,N_6322,N_6269);
nand U7270 (N_7270,N_6704,N_6309);
nand U7271 (N_7271,N_6498,N_6230);
nand U7272 (N_7272,N_6184,N_6040);
nor U7273 (N_7273,N_6313,N_6287);
nor U7274 (N_7274,N_6367,N_6457);
nand U7275 (N_7275,N_6608,N_6664);
and U7276 (N_7276,N_6294,N_6543);
nand U7277 (N_7277,N_6689,N_6474);
nor U7278 (N_7278,N_6393,N_6528);
or U7279 (N_7279,N_6689,N_6191);
and U7280 (N_7280,N_6557,N_6119);
and U7281 (N_7281,N_6026,N_6514);
nor U7282 (N_7282,N_6012,N_6382);
nand U7283 (N_7283,N_6745,N_6611);
nor U7284 (N_7284,N_6080,N_6642);
nand U7285 (N_7285,N_6399,N_6046);
nand U7286 (N_7286,N_6069,N_6083);
xnor U7287 (N_7287,N_6437,N_6611);
nor U7288 (N_7288,N_6553,N_6631);
nand U7289 (N_7289,N_6395,N_6166);
or U7290 (N_7290,N_6374,N_6580);
or U7291 (N_7291,N_6082,N_6666);
and U7292 (N_7292,N_6519,N_6041);
nor U7293 (N_7293,N_6529,N_6019);
xor U7294 (N_7294,N_6509,N_6053);
or U7295 (N_7295,N_6504,N_6701);
xnor U7296 (N_7296,N_6478,N_6582);
xnor U7297 (N_7297,N_6605,N_6743);
xnor U7298 (N_7298,N_6509,N_6664);
and U7299 (N_7299,N_6286,N_6459);
nand U7300 (N_7300,N_6657,N_6326);
xor U7301 (N_7301,N_6410,N_6359);
xor U7302 (N_7302,N_6514,N_6484);
xor U7303 (N_7303,N_6143,N_6296);
xor U7304 (N_7304,N_6635,N_6011);
and U7305 (N_7305,N_6440,N_6593);
nand U7306 (N_7306,N_6491,N_6454);
xnor U7307 (N_7307,N_6067,N_6138);
or U7308 (N_7308,N_6199,N_6300);
nand U7309 (N_7309,N_6678,N_6149);
and U7310 (N_7310,N_6046,N_6364);
nand U7311 (N_7311,N_6549,N_6076);
nor U7312 (N_7312,N_6695,N_6689);
or U7313 (N_7313,N_6092,N_6077);
xor U7314 (N_7314,N_6649,N_6366);
or U7315 (N_7315,N_6319,N_6044);
xor U7316 (N_7316,N_6437,N_6519);
nand U7317 (N_7317,N_6307,N_6197);
or U7318 (N_7318,N_6203,N_6738);
xnor U7319 (N_7319,N_6309,N_6529);
nand U7320 (N_7320,N_6364,N_6459);
xor U7321 (N_7321,N_6288,N_6080);
xor U7322 (N_7322,N_6311,N_6644);
nor U7323 (N_7323,N_6218,N_6372);
or U7324 (N_7324,N_6173,N_6423);
or U7325 (N_7325,N_6401,N_6681);
nor U7326 (N_7326,N_6286,N_6083);
or U7327 (N_7327,N_6708,N_6496);
and U7328 (N_7328,N_6733,N_6209);
or U7329 (N_7329,N_6615,N_6393);
nand U7330 (N_7330,N_6355,N_6291);
and U7331 (N_7331,N_6338,N_6600);
or U7332 (N_7332,N_6402,N_6226);
nand U7333 (N_7333,N_6690,N_6005);
nor U7334 (N_7334,N_6436,N_6237);
or U7335 (N_7335,N_6213,N_6572);
nor U7336 (N_7336,N_6334,N_6659);
nor U7337 (N_7337,N_6031,N_6612);
xnor U7338 (N_7338,N_6057,N_6280);
nor U7339 (N_7339,N_6419,N_6000);
or U7340 (N_7340,N_6410,N_6488);
nor U7341 (N_7341,N_6429,N_6437);
xor U7342 (N_7342,N_6276,N_6403);
nand U7343 (N_7343,N_6524,N_6322);
and U7344 (N_7344,N_6708,N_6520);
or U7345 (N_7345,N_6290,N_6453);
and U7346 (N_7346,N_6008,N_6346);
or U7347 (N_7347,N_6024,N_6529);
and U7348 (N_7348,N_6519,N_6076);
nand U7349 (N_7349,N_6427,N_6644);
xor U7350 (N_7350,N_6684,N_6542);
xnor U7351 (N_7351,N_6545,N_6115);
xnor U7352 (N_7352,N_6594,N_6131);
nand U7353 (N_7353,N_6285,N_6142);
xnor U7354 (N_7354,N_6198,N_6098);
nand U7355 (N_7355,N_6514,N_6376);
or U7356 (N_7356,N_6057,N_6222);
xor U7357 (N_7357,N_6330,N_6245);
and U7358 (N_7358,N_6677,N_6642);
xor U7359 (N_7359,N_6432,N_6175);
and U7360 (N_7360,N_6595,N_6351);
or U7361 (N_7361,N_6165,N_6132);
and U7362 (N_7362,N_6683,N_6503);
or U7363 (N_7363,N_6196,N_6241);
xor U7364 (N_7364,N_6443,N_6042);
and U7365 (N_7365,N_6611,N_6614);
nand U7366 (N_7366,N_6704,N_6515);
or U7367 (N_7367,N_6101,N_6600);
or U7368 (N_7368,N_6076,N_6725);
and U7369 (N_7369,N_6466,N_6098);
xnor U7370 (N_7370,N_6725,N_6656);
or U7371 (N_7371,N_6361,N_6134);
or U7372 (N_7372,N_6379,N_6611);
and U7373 (N_7373,N_6075,N_6715);
or U7374 (N_7374,N_6350,N_6420);
and U7375 (N_7375,N_6549,N_6306);
nand U7376 (N_7376,N_6141,N_6189);
or U7377 (N_7377,N_6131,N_6236);
xnor U7378 (N_7378,N_6669,N_6649);
xnor U7379 (N_7379,N_6709,N_6626);
nand U7380 (N_7380,N_6235,N_6090);
or U7381 (N_7381,N_6352,N_6458);
nor U7382 (N_7382,N_6306,N_6694);
nor U7383 (N_7383,N_6032,N_6743);
xnor U7384 (N_7384,N_6456,N_6186);
xor U7385 (N_7385,N_6090,N_6543);
or U7386 (N_7386,N_6479,N_6659);
nor U7387 (N_7387,N_6687,N_6242);
and U7388 (N_7388,N_6461,N_6253);
or U7389 (N_7389,N_6599,N_6219);
xnor U7390 (N_7390,N_6318,N_6748);
and U7391 (N_7391,N_6581,N_6112);
and U7392 (N_7392,N_6257,N_6703);
and U7393 (N_7393,N_6739,N_6205);
nor U7394 (N_7394,N_6185,N_6699);
or U7395 (N_7395,N_6370,N_6712);
and U7396 (N_7396,N_6716,N_6040);
nand U7397 (N_7397,N_6581,N_6233);
or U7398 (N_7398,N_6374,N_6202);
nor U7399 (N_7399,N_6490,N_6714);
xnor U7400 (N_7400,N_6127,N_6068);
or U7401 (N_7401,N_6099,N_6218);
xor U7402 (N_7402,N_6096,N_6284);
or U7403 (N_7403,N_6306,N_6452);
and U7404 (N_7404,N_6187,N_6548);
and U7405 (N_7405,N_6180,N_6297);
nor U7406 (N_7406,N_6184,N_6603);
and U7407 (N_7407,N_6630,N_6500);
or U7408 (N_7408,N_6325,N_6195);
xor U7409 (N_7409,N_6719,N_6222);
or U7410 (N_7410,N_6345,N_6289);
xor U7411 (N_7411,N_6038,N_6626);
nor U7412 (N_7412,N_6137,N_6430);
and U7413 (N_7413,N_6437,N_6118);
or U7414 (N_7414,N_6350,N_6446);
nor U7415 (N_7415,N_6480,N_6346);
or U7416 (N_7416,N_6143,N_6437);
xnor U7417 (N_7417,N_6670,N_6493);
nand U7418 (N_7418,N_6190,N_6542);
xnor U7419 (N_7419,N_6095,N_6625);
nor U7420 (N_7420,N_6151,N_6382);
nor U7421 (N_7421,N_6138,N_6456);
or U7422 (N_7422,N_6575,N_6396);
nand U7423 (N_7423,N_6327,N_6532);
or U7424 (N_7424,N_6385,N_6326);
xnor U7425 (N_7425,N_6369,N_6607);
nor U7426 (N_7426,N_6137,N_6637);
and U7427 (N_7427,N_6342,N_6207);
nor U7428 (N_7428,N_6644,N_6720);
or U7429 (N_7429,N_6484,N_6392);
nand U7430 (N_7430,N_6516,N_6071);
xnor U7431 (N_7431,N_6419,N_6085);
nand U7432 (N_7432,N_6054,N_6210);
nand U7433 (N_7433,N_6287,N_6738);
xnor U7434 (N_7434,N_6669,N_6454);
nand U7435 (N_7435,N_6147,N_6459);
xnor U7436 (N_7436,N_6175,N_6532);
nand U7437 (N_7437,N_6454,N_6066);
or U7438 (N_7438,N_6358,N_6636);
or U7439 (N_7439,N_6707,N_6291);
and U7440 (N_7440,N_6580,N_6713);
xnor U7441 (N_7441,N_6650,N_6651);
and U7442 (N_7442,N_6133,N_6257);
nand U7443 (N_7443,N_6507,N_6185);
nor U7444 (N_7444,N_6286,N_6485);
xor U7445 (N_7445,N_6719,N_6723);
nor U7446 (N_7446,N_6007,N_6736);
nor U7447 (N_7447,N_6172,N_6218);
xnor U7448 (N_7448,N_6248,N_6001);
nand U7449 (N_7449,N_6347,N_6432);
and U7450 (N_7450,N_6196,N_6316);
xnor U7451 (N_7451,N_6479,N_6624);
or U7452 (N_7452,N_6178,N_6411);
or U7453 (N_7453,N_6176,N_6737);
nor U7454 (N_7454,N_6173,N_6188);
nand U7455 (N_7455,N_6125,N_6022);
and U7456 (N_7456,N_6321,N_6538);
and U7457 (N_7457,N_6711,N_6691);
xnor U7458 (N_7458,N_6437,N_6295);
nor U7459 (N_7459,N_6278,N_6595);
nand U7460 (N_7460,N_6629,N_6159);
or U7461 (N_7461,N_6071,N_6336);
or U7462 (N_7462,N_6306,N_6263);
nor U7463 (N_7463,N_6686,N_6531);
nor U7464 (N_7464,N_6607,N_6243);
xnor U7465 (N_7465,N_6569,N_6372);
xor U7466 (N_7466,N_6380,N_6441);
or U7467 (N_7467,N_6690,N_6123);
nand U7468 (N_7468,N_6038,N_6034);
nor U7469 (N_7469,N_6031,N_6559);
or U7470 (N_7470,N_6111,N_6020);
nand U7471 (N_7471,N_6175,N_6593);
nor U7472 (N_7472,N_6166,N_6576);
or U7473 (N_7473,N_6474,N_6579);
nor U7474 (N_7474,N_6106,N_6213);
xor U7475 (N_7475,N_6583,N_6461);
xnor U7476 (N_7476,N_6122,N_6534);
and U7477 (N_7477,N_6178,N_6016);
nor U7478 (N_7478,N_6154,N_6595);
and U7479 (N_7479,N_6355,N_6040);
nand U7480 (N_7480,N_6071,N_6673);
nand U7481 (N_7481,N_6727,N_6055);
nor U7482 (N_7482,N_6075,N_6030);
nor U7483 (N_7483,N_6614,N_6700);
nand U7484 (N_7484,N_6609,N_6633);
xnor U7485 (N_7485,N_6033,N_6501);
and U7486 (N_7486,N_6325,N_6492);
and U7487 (N_7487,N_6238,N_6702);
and U7488 (N_7488,N_6239,N_6016);
nand U7489 (N_7489,N_6279,N_6346);
and U7490 (N_7490,N_6047,N_6727);
nand U7491 (N_7491,N_6631,N_6690);
or U7492 (N_7492,N_6192,N_6042);
and U7493 (N_7493,N_6126,N_6229);
nand U7494 (N_7494,N_6740,N_6345);
xor U7495 (N_7495,N_6179,N_6079);
or U7496 (N_7496,N_6584,N_6424);
xor U7497 (N_7497,N_6138,N_6498);
and U7498 (N_7498,N_6058,N_6709);
or U7499 (N_7499,N_6551,N_6274);
xnor U7500 (N_7500,N_7282,N_7273);
nor U7501 (N_7501,N_7358,N_7387);
nand U7502 (N_7502,N_7263,N_7042);
nand U7503 (N_7503,N_7089,N_6892);
nand U7504 (N_7504,N_7439,N_7007);
nor U7505 (N_7505,N_7253,N_6985);
nand U7506 (N_7506,N_7090,N_7385);
and U7507 (N_7507,N_7362,N_7075);
or U7508 (N_7508,N_7404,N_6866);
and U7509 (N_7509,N_6889,N_7411);
or U7510 (N_7510,N_6934,N_6851);
and U7511 (N_7511,N_7058,N_7419);
and U7512 (N_7512,N_7400,N_6990);
or U7513 (N_7513,N_6793,N_7196);
nor U7514 (N_7514,N_7124,N_6905);
xor U7515 (N_7515,N_7107,N_7014);
xor U7516 (N_7516,N_6893,N_6918);
xnor U7517 (N_7517,N_6858,N_7488);
xnor U7518 (N_7518,N_7159,N_6783);
nor U7519 (N_7519,N_6843,N_6844);
nor U7520 (N_7520,N_6827,N_6862);
nand U7521 (N_7521,N_7079,N_7341);
xor U7522 (N_7522,N_7366,N_6823);
nor U7523 (N_7523,N_7451,N_7175);
or U7524 (N_7524,N_6886,N_6838);
nand U7525 (N_7525,N_6845,N_7053);
or U7526 (N_7526,N_6920,N_6933);
nand U7527 (N_7527,N_7199,N_6829);
and U7528 (N_7528,N_7453,N_7417);
xor U7529 (N_7529,N_7349,N_7035);
or U7530 (N_7530,N_7003,N_7134);
nand U7531 (N_7531,N_7347,N_7470);
and U7532 (N_7532,N_7157,N_7493);
nor U7533 (N_7533,N_6774,N_6841);
and U7534 (N_7534,N_7085,N_6804);
or U7535 (N_7535,N_7467,N_7337);
nand U7536 (N_7536,N_6812,N_7006);
nor U7537 (N_7537,N_7350,N_7184);
nand U7538 (N_7538,N_7285,N_7128);
and U7539 (N_7539,N_7428,N_7211);
and U7540 (N_7540,N_6924,N_7067);
xnor U7541 (N_7541,N_7235,N_6971);
nand U7542 (N_7542,N_7438,N_7275);
xnor U7543 (N_7543,N_7179,N_6825);
and U7544 (N_7544,N_7143,N_7297);
and U7545 (N_7545,N_7495,N_6782);
xor U7546 (N_7546,N_6968,N_7474);
and U7547 (N_7547,N_6813,N_7078);
nor U7548 (N_7548,N_7039,N_6805);
nand U7549 (N_7549,N_7312,N_7048);
or U7550 (N_7550,N_6810,N_6904);
nand U7551 (N_7551,N_7455,N_7471);
nor U7552 (N_7552,N_7046,N_6945);
nor U7553 (N_7553,N_6791,N_7038);
nor U7554 (N_7554,N_7325,N_6751);
nand U7555 (N_7555,N_7348,N_7465);
and U7556 (N_7556,N_6943,N_7205);
or U7557 (N_7557,N_6761,N_7413);
nand U7558 (N_7558,N_6980,N_7340);
nand U7559 (N_7559,N_7497,N_7204);
xor U7560 (N_7560,N_7069,N_6779);
nand U7561 (N_7561,N_6868,N_7146);
nor U7562 (N_7562,N_7167,N_7278);
and U7563 (N_7563,N_7437,N_6969);
or U7564 (N_7564,N_7216,N_7005);
and U7565 (N_7565,N_7448,N_6898);
xnor U7566 (N_7566,N_6954,N_7298);
or U7567 (N_7567,N_7310,N_7445);
and U7568 (N_7568,N_6917,N_6788);
nand U7569 (N_7569,N_7363,N_6972);
xor U7570 (N_7570,N_7082,N_6789);
and U7571 (N_7571,N_7255,N_7441);
nand U7572 (N_7572,N_6887,N_6847);
nor U7573 (N_7573,N_7477,N_7252);
or U7574 (N_7574,N_6902,N_7209);
nand U7575 (N_7575,N_6808,N_7080);
or U7576 (N_7576,N_7262,N_7496);
and U7577 (N_7577,N_7197,N_6894);
or U7578 (N_7578,N_7045,N_7489);
or U7579 (N_7579,N_7420,N_7449);
nand U7580 (N_7580,N_6869,N_7102);
and U7581 (N_7581,N_7326,N_7190);
nand U7582 (N_7582,N_7403,N_7304);
or U7583 (N_7583,N_6901,N_6935);
and U7584 (N_7584,N_6867,N_7025);
xor U7585 (N_7585,N_7145,N_7333);
or U7586 (N_7586,N_7207,N_7189);
nor U7587 (N_7587,N_6981,N_7029);
nand U7588 (N_7588,N_7414,N_6773);
or U7589 (N_7589,N_7081,N_7402);
nor U7590 (N_7590,N_7461,N_7137);
or U7591 (N_7591,N_6883,N_6856);
xor U7592 (N_7592,N_7138,N_6932);
xor U7593 (N_7593,N_6993,N_7068);
or U7594 (N_7594,N_6963,N_7126);
nor U7595 (N_7595,N_7231,N_7458);
or U7596 (N_7596,N_7462,N_6854);
xnor U7597 (N_7597,N_7247,N_7321);
nor U7598 (N_7598,N_7418,N_7222);
nor U7599 (N_7599,N_6996,N_7272);
or U7600 (N_7600,N_7338,N_7036);
xor U7601 (N_7601,N_7425,N_7074);
xor U7602 (N_7602,N_6863,N_7044);
or U7603 (N_7603,N_7062,N_7352);
nor U7604 (N_7604,N_7299,N_6978);
and U7605 (N_7605,N_7371,N_7239);
or U7606 (N_7606,N_7416,N_7236);
nand U7607 (N_7607,N_6872,N_6919);
xnor U7608 (N_7608,N_6938,N_7113);
and U7609 (N_7609,N_7457,N_7423);
xnor U7610 (N_7610,N_7379,N_6873);
nor U7611 (N_7611,N_6766,N_7181);
nor U7612 (N_7612,N_7040,N_7095);
nor U7613 (N_7613,N_6835,N_7215);
nor U7614 (N_7614,N_7330,N_7319);
nor U7615 (N_7615,N_7224,N_7193);
xnor U7616 (N_7616,N_6786,N_7469);
nand U7617 (N_7617,N_7478,N_6819);
and U7618 (N_7618,N_7206,N_7452);
nand U7619 (N_7619,N_7233,N_6907);
xor U7620 (N_7620,N_7315,N_6961);
or U7621 (N_7621,N_7261,N_6994);
or U7622 (N_7622,N_7234,N_7249);
nand U7623 (N_7623,N_7408,N_6754);
xnor U7624 (N_7624,N_7033,N_7266);
nand U7625 (N_7625,N_7093,N_7480);
xnor U7626 (N_7626,N_6949,N_6794);
xnor U7627 (N_7627,N_7447,N_6846);
nand U7628 (N_7628,N_6855,N_6973);
or U7629 (N_7629,N_6865,N_7001);
xnor U7630 (N_7630,N_6861,N_7066);
xnor U7631 (N_7631,N_6900,N_6952);
nor U7632 (N_7632,N_7208,N_7336);
nor U7633 (N_7633,N_7191,N_7434);
and U7634 (N_7634,N_7294,N_7372);
nand U7635 (N_7635,N_7141,N_7043);
nand U7636 (N_7636,N_7086,N_6914);
or U7637 (N_7637,N_7210,N_7188);
nor U7638 (N_7638,N_7218,N_7361);
nand U7639 (N_7639,N_7169,N_7355);
nor U7640 (N_7640,N_7228,N_6776);
nand U7641 (N_7641,N_6832,N_7246);
xnor U7642 (N_7642,N_7257,N_6908);
and U7643 (N_7643,N_7070,N_7422);
nand U7644 (N_7644,N_7398,N_6840);
and U7645 (N_7645,N_7027,N_7055);
nor U7646 (N_7646,N_7380,N_6822);
nand U7647 (N_7647,N_6770,N_7016);
or U7648 (N_7648,N_7073,N_7407);
or U7649 (N_7649,N_6848,N_7435);
or U7650 (N_7650,N_7083,N_7329);
xor U7651 (N_7651,N_7056,N_6884);
and U7652 (N_7652,N_7251,N_7415);
nand U7653 (N_7653,N_6929,N_7201);
nand U7654 (N_7654,N_7172,N_7032);
and U7655 (N_7655,N_7162,N_6926);
nor U7656 (N_7656,N_6828,N_7443);
and U7657 (N_7657,N_7047,N_7111);
xor U7658 (N_7658,N_7354,N_7308);
xor U7659 (N_7659,N_6801,N_7050);
nand U7660 (N_7660,N_7116,N_7163);
or U7661 (N_7661,N_7060,N_6842);
nor U7662 (N_7662,N_6916,N_7139);
or U7663 (N_7663,N_6906,N_6975);
xor U7664 (N_7664,N_7421,N_6799);
xor U7665 (N_7665,N_7002,N_6998);
xor U7666 (N_7666,N_7314,N_7433);
nand U7667 (N_7667,N_6979,N_6850);
nor U7668 (N_7668,N_7142,N_7287);
and U7669 (N_7669,N_6821,N_7061);
and U7670 (N_7670,N_7316,N_7160);
or U7671 (N_7671,N_7466,N_7270);
xnor U7672 (N_7672,N_6756,N_6957);
nor U7673 (N_7673,N_7374,N_7327);
and U7674 (N_7674,N_6967,N_6922);
nand U7675 (N_7675,N_6896,N_7412);
nand U7676 (N_7676,N_7096,N_7268);
or U7677 (N_7677,N_7401,N_7388);
and U7678 (N_7678,N_7098,N_7094);
and U7679 (N_7679,N_7307,N_7344);
or U7680 (N_7680,N_7490,N_7313);
nand U7681 (N_7681,N_7456,N_7103);
nand U7682 (N_7682,N_6950,N_6798);
nand U7683 (N_7683,N_7010,N_7396);
xnor U7684 (N_7684,N_7147,N_7226);
nand U7685 (N_7685,N_6940,N_6878);
xor U7686 (N_7686,N_7158,N_7265);
nor U7687 (N_7687,N_6765,N_7463);
or U7688 (N_7688,N_7301,N_7243);
and U7689 (N_7689,N_7464,N_7332);
nand U7690 (N_7690,N_6853,N_6925);
xor U7691 (N_7691,N_6942,N_6879);
and U7692 (N_7692,N_7133,N_7108);
xor U7693 (N_7693,N_7009,N_6809);
nand U7694 (N_7694,N_6936,N_6755);
xnor U7695 (N_7695,N_7383,N_7335);
nand U7696 (N_7696,N_6912,N_6830);
or U7697 (N_7697,N_7284,N_7486);
nand U7698 (N_7698,N_7436,N_7409);
nand U7699 (N_7699,N_7072,N_7140);
nor U7700 (N_7700,N_7424,N_7302);
or U7701 (N_7701,N_7250,N_7057);
nand U7702 (N_7702,N_6790,N_6881);
nor U7703 (N_7703,N_7154,N_7394);
or U7704 (N_7704,N_7012,N_7345);
and U7705 (N_7705,N_7034,N_7240);
and U7706 (N_7706,N_6891,N_7019);
or U7707 (N_7707,N_7136,N_6923);
xor U7708 (N_7708,N_6913,N_7386);
xnor U7709 (N_7709,N_6928,N_7306);
nor U7710 (N_7710,N_7018,N_7109);
xnor U7711 (N_7711,N_6882,N_7024);
nor U7712 (N_7712,N_7397,N_7173);
xor U7713 (N_7713,N_7238,N_7125);
and U7714 (N_7714,N_7292,N_7367);
or U7715 (N_7715,N_7256,N_6817);
nor U7716 (N_7716,N_7309,N_7390);
nand U7717 (N_7717,N_7161,N_7318);
nand U7718 (N_7718,N_7473,N_6997);
and U7719 (N_7719,N_6852,N_7377);
xnor U7720 (N_7720,N_7166,N_7324);
or U7721 (N_7721,N_7092,N_7446);
or U7722 (N_7722,N_7264,N_6777);
or U7723 (N_7723,N_7219,N_6947);
nand U7724 (N_7724,N_6834,N_7475);
nand U7725 (N_7725,N_7391,N_7221);
and U7726 (N_7726,N_7015,N_6764);
and U7727 (N_7727,N_7198,N_6989);
nand U7728 (N_7728,N_7130,N_6937);
or U7729 (N_7729,N_7150,N_7339);
xnor U7730 (N_7730,N_7099,N_7353);
nor U7731 (N_7731,N_7481,N_7091);
nor U7732 (N_7732,N_7037,N_6897);
and U7733 (N_7733,N_7454,N_7430);
nand U7734 (N_7734,N_7122,N_6849);
and U7735 (N_7735,N_6955,N_7271);
and U7736 (N_7736,N_7364,N_6910);
or U7737 (N_7737,N_6772,N_7357);
and U7738 (N_7738,N_7176,N_7008);
nor U7739 (N_7739,N_7373,N_7135);
nand U7740 (N_7740,N_7399,N_7063);
or U7741 (N_7741,N_7290,N_6807);
xnor U7742 (N_7742,N_6903,N_7320);
or U7743 (N_7743,N_7245,N_7071);
nor U7744 (N_7744,N_7476,N_7187);
nor U7745 (N_7745,N_6816,N_7180);
or U7746 (N_7746,N_6826,N_6802);
xnor U7747 (N_7747,N_7021,N_6984);
nor U7748 (N_7748,N_7054,N_7123);
and U7749 (N_7749,N_7485,N_6836);
xor U7750 (N_7750,N_7393,N_7195);
nor U7751 (N_7751,N_6800,N_6899);
nor U7752 (N_7752,N_7291,N_6960);
or U7753 (N_7753,N_7186,N_7051);
or U7754 (N_7754,N_7482,N_6871);
nand U7755 (N_7755,N_6760,N_7152);
and U7756 (N_7756,N_6966,N_7498);
and U7757 (N_7757,N_6964,N_7356);
or U7758 (N_7758,N_7227,N_7178);
nor U7759 (N_7759,N_7115,N_7392);
nor U7760 (N_7760,N_7484,N_7431);
nand U7761 (N_7761,N_7028,N_7217);
and U7762 (N_7762,N_7494,N_7395);
nor U7763 (N_7763,N_6987,N_6931);
nor U7764 (N_7764,N_6870,N_7148);
xnor U7765 (N_7765,N_7254,N_7155);
nor U7766 (N_7766,N_6752,N_7279);
nor U7767 (N_7767,N_6885,N_7288);
nor U7768 (N_7768,N_7202,N_6953);
nand U7769 (N_7769,N_7351,N_7293);
and U7770 (N_7770,N_6806,N_7220);
or U7771 (N_7771,N_6860,N_6771);
xor U7772 (N_7772,N_7213,N_6768);
nand U7773 (N_7773,N_6930,N_6875);
nor U7774 (N_7774,N_6757,N_7317);
xnor U7775 (N_7775,N_7479,N_6948);
xnor U7776 (N_7776,N_6767,N_6784);
nand U7777 (N_7777,N_6946,N_6951);
or U7778 (N_7778,N_7328,N_6895);
or U7779 (N_7779,N_7442,N_7346);
or U7780 (N_7780,N_6750,N_7030);
xor U7781 (N_7781,N_7237,N_7011);
or U7782 (N_7782,N_7276,N_6864);
or U7783 (N_7783,N_7017,N_6814);
or U7784 (N_7784,N_7120,N_6956);
nor U7785 (N_7785,N_7472,N_7013);
or U7786 (N_7786,N_7432,N_7118);
xor U7787 (N_7787,N_7440,N_7084);
xnor U7788 (N_7788,N_6837,N_7059);
and U7789 (N_7789,N_7097,N_6965);
nand U7790 (N_7790,N_7381,N_7365);
and U7791 (N_7791,N_7375,N_6758);
nand U7792 (N_7792,N_6983,N_7064);
nor U7793 (N_7793,N_7214,N_6839);
xor U7794 (N_7794,N_6753,N_6921);
xor U7795 (N_7795,N_6763,N_7132);
nand U7796 (N_7796,N_7200,N_7259);
xor U7797 (N_7797,N_7331,N_7104);
xnor U7798 (N_7798,N_7174,N_7376);
nor U7799 (N_7799,N_7444,N_6941);
nand U7800 (N_7800,N_6977,N_6999);
nor U7801 (N_7801,N_7369,N_6857);
nor U7802 (N_7802,N_7323,N_7182);
nand U7803 (N_7803,N_7105,N_6781);
or U7804 (N_7804,N_7170,N_7110);
and U7805 (N_7805,N_7177,N_6991);
nand U7806 (N_7806,N_7242,N_6944);
xnor U7807 (N_7807,N_6803,N_6785);
and U7808 (N_7808,N_6874,N_7119);
xnor U7809 (N_7809,N_6815,N_6769);
and U7810 (N_7810,N_6915,N_6787);
nand U7811 (N_7811,N_7429,N_7280);
nand U7812 (N_7812,N_7131,N_6988);
and U7813 (N_7813,N_7487,N_7129);
and U7814 (N_7814,N_7117,N_7258);
nand U7815 (N_7815,N_7260,N_7343);
or U7816 (N_7816,N_6909,N_7426);
xnor U7817 (N_7817,N_7491,N_6780);
nor U7818 (N_7818,N_6995,N_7168);
nand U7819 (N_7819,N_6796,N_7460);
nor U7820 (N_7820,N_7049,N_7026);
nor U7821 (N_7821,N_7274,N_7322);
nand U7822 (N_7822,N_6974,N_7223);
and U7823 (N_7823,N_7410,N_6890);
xor U7824 (N_7824,N_7165,N_7153);
or U7825 (N_7825,N_6762,N_6959);
nor U7826 (N_7826,N_7241,N_6859);
nand U7827 (N_7827,N_7212,N_7076);
nand U7828 (N_7828,N_6939,N_7359);
nor U7829 (N_7829,N_7267,N_7281);
and U7830 (N_7830,N_7368,N_7450);
and U7831 (N_7831,N_7192,N_6792);
xor U7832 (N_7832,N_6818,N_7334);
xor U7833 (N_7833,N_7000,N_7295);
and U7834 (N_7834,N_7112,N_7031);
or U7835 (N_7835,N_7311,N_7041);
or U7836 (N_7836,N_7203,N_7360);
and U7837 (N_7837,N_7342,N_7406);
and U7838 (N_7838,N_7121,N_7164);
and U7839 (N_7839,N_6976,N_7370);
nor U7840 (N_7840,N_7303,N_7289);
and U7841 (N_7841,N_7185,N_7144);
and U7842 (N_7842,N_7127,N_7244);
nor U7843 (N_7843,N_7468,N_7100);
nor U7844 (N_7844,N_6831,N_7300);
nor U7845 (N_7845,N_7183,N_7225);
nor U7846 (N_7846,N_7101,N_6797);
nand U7847 (N_7847,N_7106,N_7405);
and U7848 (N_7848,N_7384,N_6911);
nand U7849 (N_7849,N_6992,N_7149);
nor U7850 (N_7850,N_7022,N_6876);
or U7851 (N_7851,N_6877,N_7151);
nor U7852 (N_7852,N_7305,N_7427);
nand U7853 (N_7853,N_7194,N_6759);
nor U7854 (N_7854,N_6775,N_6778);
nor U7855 (N_7855,N_7378,N_7020);
xor U7856 (N_7856,N_7077,N_6880);
xnor U7857 (N_7857,N_6820,N_6811);
nand U7858 (N_7858,N_7023,N_7229);
or U7859 (N_7859,N_7277,N_6927);
or U7860 (N_7860,N_7065,N_7296);
and U7861 (N_7861,N_7499,N_7389);
xnor U7862 (N_7862,N_7052,N_7483);
nor U7863 (N_7863,N_6795,N_7088);
or U7864 (N_7864,N_7114,N_7283);
nor U7865 (N_7865,N_7382,N_7232);
xnor U7866 (N_7866,N_6833,N_6958);
and U7867 (N_7867,N_7004,N_7156);
nor U7868 (N_7868,N_7230,N_7286);
or U7869 (N_7869,N_6970,N_6982);
and U7870 (N_7870,N_7087,N_7492);
nor U7871 (N_7871,N_6986,N_6888);
or U7872 (N_7872,N_6962,N_7248);
or U7873 (N_7873,N_6824,N_7269);
or U7874 (N_7874,N_7459,N_7171);
nand U7875 (N_7875,N_7303,N_7264);
or U7876 (N_7876,N_7152,N_6865);
or U7877 (N_7877,N_7422,N_6824);
and U7878 (N_7878,N_7091,N_7486);
xor U7879 (N_7879,N_7388,N_6996);
nand U7880 (N_7880,N_6905,N_7472);
or U7881 (N_7881,N_7480,N_7024);
nor U7882 (N_7882,N_6887,N_7297);
nand U7883 (N_7883,N_7015,N_7168);
xor U7884 (N_7884,N_7000,N_7122);
xor U7885 (N_7885,N_7015,N_7090);
xnor U7886 (N_7886,N_6837,N_6816);
xnor U7887 (N_7887,N_7438,N_7425);
and U7888 (N_7888,N_7478,N_7243);
or U7889 (N_7889,N_7357,N_6987);
nor U7890 (N_7890,N_6915,N_7472);
or U7891 (N_7891,N_6774,N_7422);
nand U7892 (N_7892,N_7127,N_7386);
xor U7893 (N_7893,N_7388,N_7301);
and U7894 (N_7894,N_7155,N_7099);
or U7895 (N_7895,N_7439,N_7020);
xor U7896 (N_7896,N_6778,N_7449);
nand U7897 (N_7897,N_7433,N_7177);
or U7898 (N_7898,N_7372,N_7262);
or U7899 (N_7899,N_7002,N_6966);
nand U7900 (N_7900,N_6767,N_6839);
nor U7901 (N_7901,N_6859,N_7021);
or U7902 (N_7902,N_6972,N_7414);
or U7903 (N_7903,N_6998,N_6887);
nand U7904 (N_7904,N_7126,N_6781);
or U7905 (N_7905,N_7087,N_6865);
or U7906 (N_7906,N_6971,N_6884);
or U7907 (N_7907,N_6887,N_7091);
or U7908 (N_7908,N_7180,N_6974);
xnor U7909 (N_7909,N_7480,N_7092);
nand U7910 (N_7910,N_7388,N_7414);
or U7911 (N_7911,N_6817,N_7191);
and U7912 (N_7912,N_6787,N_7480);
nand U7913 (N_7913,N_6827,N_6891);
nor U7914 (N_7914,N_6934,N_6922);
or U7915 (N_7915,N_7021,N_6946);
or U7916 (N_7916,N_7075,N_7079);
nor U7917 (N_7917,N_6909,N_6866);
nand U7918 (N_7918,N_6756,N_7460);
xnor U7919 (N_7919,N_6788,N_7322);
nand U7920 (N_7920,N_7472,N_6974);
or U7921 (N_7921,N_7407,N_7106);
and U7922 (N_7922,N_7018,N_7023);
nand U7923 (N_7923,N_7247,N_7031);
and U7924 (N_7924,N_6931,N_7153);
xor U7925 (N_7925,N_6941,N_7026);
xor U7926 (N_7926,N_7207,N_7473);
nor U7927 (N_7927,N_7153,N_6841);
nor U7928 (N_7928,N_6797,N_6929);
nor U7929 (N_7929,N_7177,N_7034);
xnor U7930 (N_7930,N_7120,N_7451);
nand U7931 (N_7931,N_6933,N_7283);
nand U7932 (N_7932,N_7328,N_7120);
xnor U7933 (N_7933,N_7435,N_7321);
xnor U7934 (N_7934,N_6971,N_7376);
or U7935 (N_7935,N_6925,N_7226);
xnor U7936 (N_7936,N_7314,N_7019);
nand U7937 (N_7937,N_6786,N_7299);
xor U7938 (N_7938,N_7430,N_7257);
or U7939 (N_7939,N_6751,N_7360);
xnor U7940 (N_7940,N_7249,N_7012);
and U7941 (N_7941,N_6822,N_7327);
nand U7942 (N_7942,N_7065,N_6989);
and U7943 (N_7943,N_7272,N_7266);
xnor U7944 (N_7944,N_6823,N_7087);
nor U7945 (N_7945,N_7380,N_7246);
nand U7946 (N_7946,N_7221,N_6781);
or U7947 (N_7947,N_7400,N_7278);
or U7948 (N_7948,N_7153,N_7475);
nor U7949 (N_7949,N_6980,N_6833);
nand U7950 (N_7950,N_7440,N_6825);
nor U7951 (N_7951,N_6821,N_7283);
and U7952 (N_7952,N_7303,N_7248);
nand U7953 (N_7953,N_6835,N_7165);
nor U7954 (N_7954,N_6874,N_7302);
xor U7955 (N_7955,N_7313,N_7310);
nor U7956 (N_7956,N_7243,N_7015);
nand U7957 (N_7957,N_7322,N_7206);
nand U7958 (N_7958,N_6789,N_6853);
xnor U7959 (N_7959,N_7061,N_7118);
nor U7960 (N_7960,N_7053,N_7150);
nand U7961 (N_7961,N_6752,N_7014);
xor U7962 (N_7962,N_7119,N_7256);
nor U7963 (N_7963,N_7174,N_6857);
nor U7964 (N_7964,N_7257,N_7074);
xnor U7965 (N_7965,N_7160,N_7218);
nand U7966 (N_7966,N_7106,N_6788);
nor U7967 (N_7967,N_7270,N_7262);
nand U7968 (N_7968,N_7313,N_6857);
nand U7969 (N_7969,N_6939,N_6842);
nand U7970 (N_7970,N_6836,N_7395);
and U7971 (N_7971,N_6890,N_7004);
and U7972 (N_7972,N_6767,N_6904);
and U7973 (N_7973,N_7029,N_7306);
xor U7974 (N_7974,N_6844,N_7366);
nand U7975 (N_7975,N_7184,N_6905);
or U7976 (N_7976,N_7249,N_6894);
or U7977 (N_7977,N_6806,N_6766);
xor U7978 (N_7978,N_7031,N_7337);
nand U7979 (N_7979,N_7022,N_7312);
and U7980 (N_7980,N_6942,N_7334);
nand U7981 (N_7981,N_7142,N_7347);
nor U7982 (N_7982,N_7477,N_7391);
nor U7983 (N_7983,N_7077,N_6774);
and U7984 (N_7984,N_7170,N_7264);
nand U7985 (N_7985,N_7014,N_7127);
or U7986 (N_7986,N_7222,N_6909);
nand U7987 (N_7987,N_7352,N_6927);
nand U7988 (N_7988,N_6972,N_7417);
or U7989 (N_7989,N_6846,N_6790);
nand U7990 (N_7990,N_6820,N_6793);
nand U7991 (N_7991,N_6921,N_7493);
or U7992 (N_7992,N_6779,N_6840);
and U7993 (N_7993,N_7262,N_7284);
or U7994 (N_7994,N_7189,N_6876);
and U7995 (N_7995,N_7004,N_6957);
nor U7996 (N_7996,N_6972,N_7152);
nand U7997 (N_7997,N_7410,N_6755);
and U7998 (N_7998,N_7174,N_7111);
xor U7999 (N_7999,N_7316,N_7087);
and U8000 (N_8000,N_7255,N_6773);
nand U8001 (N_8001,N_7305,N_6840);
and U8002 (N_8002,N_7181,N_7417);
xor U8003 (N_8003,N_6980,N_7094);
nor U8004 (N_8004,N_7396,N_7138);
or U8005 (N_8005,N_7160,N_6942);
and U8006 (N_8006,N_6833,N_6829);
nand U8007 (N_8007,N_6948,N_6916);
xnor U8008 (N_8008,N_7179,N_7221);
nor U8009 (N_8009,N_7457,N_6829);
xnor U8010 (N_8010,N_6936,N_7411);
xor U8011 (N_8011,N_7461,N_7130);
xor U8012 (N_8012,N_7023,N_7160);
nand U8013 (N_8013,N_7381,N_7453);
nand U8014 (N_8014,N_7388,N_7015);
and U8015 (N_8015,N_6779,N_7083);
xor U8016 (N_8016,N_7044,N_7092);
and U8017 (N_8017,N_7429,N_7159);
nand U8018 (N_8018,N_7184,N_7098);
xor U8019 (N_8019,N_7295,N_6852);
nand U8020 (N_8020,N_7470,N_7147);
and U8021 (N_8021,N_7091,N_7150);
or U8022 (N_8022,N_7101,N_6904);
or U8023 (N_8023,N_7059,N_7470);
and U8024 (N_8024,N_7250,N_7251);
nor U8025 (N_8025,N_7222,N_7271);
nand U8026 (N_8026,N_7464,N_7305);
xor U8027 (N_8027,N_7359,N_6936);
nand U8028 (N_8028,N_7131,N_7034);
and U8029 (N_8029,N_6798,N_6771);
and U8030 (N_8030,N_7275,N_7091);
or U8031 (N_8031,N_7060,N_7090);
and U8032 (N_8032,N_7240,N_6853);
xor U8033 (N_8033,N_6998,N_7315);
xnor U8034 (N_8034,N_6819,N_7019);
or U8035 (N_8035,N_7470,N_6981);
nor U8036 (N_8036,N_6792,N_6975);
xnor U8037 (N_8037,N_7287,N_7413);
or U8038 (N_8038,N_7225,N_7295);
and U8039 (N_8039,N_7375,N_7049);
xor U8040 (N_8040,N_7378,N_7399);
or U8041 (N_8041,N_7433,N_6968);
nand U8042 (N_8042,N_6870,N_7276);
nor U8043 (N_8043,N_6991,N_7102);
xnor U8044 (N_8044,N_7177,N_7319);
xor U8045 (N_8045,N_7318,N_7061);
or U8046 (N_8046,N_7007,N_7442);
xor U8047 (N_8047,N_7276,N_7417);
and U8048 (N_8048,N_7461,N_6836);
xnor U8049 (N_8049,N_7142,N_6890);
nand U8050 (N_8050,N_7408,N_7440);
nor U8051 (N_8051,N_6870,N_7312);
nor U8052 (N_8052,N_7303,N_7222);
nand U8053 (N_8053,N_7106,N_6986);
or U8054 (N_8054,N_6754,N_7280);
xor U8055 (N_8055,N_6968,N_7140);
nor U8056 (N_8056,N_7296,N_6841);
nand U8057 (N_8057,N_6806,N_7447);
nor U8058 (N_8058,N_7276,N_7126);
xnor U8059 (N_8059,N_7072,N_6900);
xnor U8060 (N_8060,N_7306,N_7309);
or U8061 (N_8061,N_6997,N_7210);
nor U8062 (N_8062,N_7310,N_6828);
nor U8063 (N_8063,N_7347,N_6818);
nor U8064 (N_8064,N_7050,N_7253);
nor U8065 (N_8065,N_7290,N_7407);
or U8066 (N_8066,N_7473,N_7175);
nand U8067 (N_8067,N_7338,N_6917);
nor U8068 (N_8068,N_7251,N_7217);
or U8069 (N_8069,N_7350,N_6910);
xor U8070 (N_8070,N_6896,N_7039);
xnor U8071 (N_8071,N_7203,N_7038);
xor U8072 (N_8072,N_7112,N_7407);
nand U8073 (N_8073,N_7170,N_7108);
nand U8074 (N_8074,N_7362,N_7475);
or U8075 (N_8075,N_7377,N_7088);
or U8076 (N_8076,N_7028,N_6959);
nor U8077 (N_8077,N_7438,N_6934);
nor U8078 (N_8078,N_7092,N_6799);
or U8079 (N_8079,N_6761,N_7325);
or U8080 (N_8080,N_6852,N_7004);
and U8081 (N_8081,N_7437,N_7370);
and U8082 (N_8082,N_7044,N_6839);
nor U8083 (N_8083,N_7098,N_6832);
nand U8084 (N_8084,N_6906,N_7100);
and U8085 (N_8085,N_6852,N_7058);
and U8086 (N_8086,N_7310,N_6873);
nand U8087 (N_8087,N_6854,N_6842);
nand U8088 (N_8088,N_7436,N_6811);
nand U8089 (N_8089,N_7244,N_7032);
and U8090 (N_8090,N_6854,N_7041);
and U8091 (N_8091,N_7299,N_7061);
and U8092 (N_8092,N_7477,N_7452);
or U8093 (N_8093,N_7264,N_6980);
xor U8094 (N_8094,N_7368,N_6954);
nand U8095 (N_8095,N_7218,N_7469);
and U8096 (N_8096,N_7469,N_7266);
nand U8097 (N_8097,N_7431,N_6840);
or U8098 (N_8098,N_6884,N_7389);
nor U8099 (N_8099,N_6952,N_7422);
nand U8100 (N_8100,N_7121,N_6803);
or U8101 (N_8101,N_7307,N_7032);
nand U8102 (N_8102,N_7038,N_7006);
and U8103 (N_8103,N_6985,N_7242);
nor U8104 (N_8104,N_7337,N_6880);
nand U8105 (N_8105,N_6844,N_7124);
nand U8106 (N_8106,N_7260,N_7120);
or U8107 (N_8107,N_6860,N_7455);
or U8108 (N_8108,N_7120,N_7463);
and U8109 (N_8109,N_7258,N_7370);
xor U8110 (N_8110,N_6999,N_7210);
and U8111 (N_8111,N_7099,N_7497);
or U8112 (N_8112,N_7187,N_7497);
nor U8113 (N_8113,N_7014,N_7276);
nor U8114 (N_8114,N_7373,N_7368);
and U8115 (N_8115,N_7198,N_7189);
nand U8116 (N_8116,N_6967,N_7412);
or U8117 (N_8117,N_6936,N_7320);
and U8118 (N_8118,N_7494,N_6796);
nand U8119 (N_8119,N_6896,N_6790);
or U8120 (N_8120,N_7359,N_6833);
nor U8121 (N_8121,N_7195,N_6849);
or U8122 (N_8122,N_7034,N_6829);
or U8123 (N_8123,N_6862,N_6802);
nor U8124 (N_8124,N_7138,N_6835);
nor U8125 (N_8125,N_6817,N_7290);
or U8126 (N_8126,N_6768,N_7341);
nand U8127 (N_8127,N_7035,N_6801);
and U8128 (N_8128,N_7203,N_7477);
xnor U8129 (N_8129,N_7407,N_7235);
nand U8130 (N_8130,N_7260,N_6960);
and U8131 (N_8131,N_7058,N_7076);
or U8132 (N_8132,N_6916,N_7238);
and U8133 (N_8133,N_7436,N_7090);
xor U8134 (N_8134,N_7457,N_7045);
nor U8135 (N_8135,N_6782,N_6842);
nor U8136 (N_8136,N_7027,N_7348);
nand U8137 (N_8137,N_7456,N_7033);
nand U8138 (N_8138,N_6853,N_7104);
xor U8139 (N_8139,N_6824,N_7367);
nand U8140 (N_8140,N_7258,N_7495);
nand U8141 (N_8141,N_6985,N_7155);
or U8142 (N_8142,N_6893,N_7029);
or U8143 (N_8143,N_7351,N_6806);
nor U8144 (N_8144,N_7158,N_7488);
nor U8145 (N_8145,N_6961,N_7086);
or U8146 (N_8146,N_7048,N_6839);
xnor U8147 (N_8147,N_6775,N_7236);
nor U8148 (N_8148,N_6992,N_6984);
xnor U8149 (N_8149,N_7494,N_6922);
and U8150 (N_8150,N_7066,N_7181);
or U8151 (N_8151,N_7289,N_7432);
nand U8152 (N_8152,N_7215,N_7093);
and U8153 (N_8153,N_7101,N_7085);
and U8154 (N_8154,N_7372,N_7155);
and U8155 (N_8155,N_6984,N_6936);
nand U8156 (N_8156,N_7348,N_6893);
or U8157 (N_8157,N_7492,N_7119);
nand U8158 (N_8158,N_7351,N_6983);
and U8159 (N_8159,N_7473,N_7179);
xor U8160 (N_8160,N_6847,N_7433);
xor U8161 (N_8161,N_7294,N_7471);
or U8162 (N_8162,N_7494,N_7371);
xnor U8163 (N_8163,N_6872,N_6892);
nand U8164 (N_8164,N_7286,N_7177);
xor U8165 (N_8165,N_7270,N_6841);
nor U8166 (N_8166,N_7122,N_6933);
nand U8167 (N_8167,N_7195,N_6875);
or U8168 (N_8168,N_7210,N_7390);
nor U8169 (N_8169,N_6884,N_7412);
or U8170 (N_8170,N_7072,N_6955);
nand U8171 (N_8171,N_7181,N_7479);
and U8172 (N_8172,N_7425,N_7034);
nand U8173 (N_8173,N_6855,N_7448);
xnor U8174 (N_8174,N_6883,N_6860);
nor U8175 (N_8175,N_7248,N_7341);
and U8176 (N_8176,N_7397,N_6922);
or U8177 (N_8177,N_7143,N_7201);
or U8178 (N_8178,N_6842,N_6761);
nand U8179 (N_8179,N_7445,N_7301);
or U8180 (N_8180,N_7036,N_6852);
or U8181 (N_8181,N_7156,N_7177);
or U8182 (N_8182,N_6991,N_6758);
nand U8183 (N_8183,N_7012,N_6794);
and U8184 (N_8184,N_7382,N_7419);
or U8185 (N_8185,N_7492,N_6844);
nor U8186 (N_8186,N_6775,N_7193);
nor U8187 (N_8187,N_7391,N_6893);
or U8188 (N_8188,N_7159,N_7091);
nor U8189 (N_8189,N_7479,N_7451);
or U8190 (N_8190,N_7026,N_7134);
nor U8191 (N_8191,N_7008,N_6987);
xor U8192 (N_8192,N_6869,N_7352);
nor U8193 (N_8193,N_6756,N_7185);
nor U8194 (N_8194,N_7405,N_6963);
nor U8195 (N_8195,N_7063,N_6968);
nand U8196 (N_8196,N_7222,N_7106);
xnor U8197 (N_8197,N_7008,N_7408);
nor U8198 (N_8198,N_7473,N_7490);
and U8199 (N_8199,N_7328,N_6959);
nor U8200 (N_8200,N_7462,N_6875);
xnor U8201 (N_8201,N_7058,N_6917);
nor U8202 (N_8202,N_6772,N_7062);
or U8203 (N_8203,N_6823,N_7013);
and U8204 (N_8204,N_7472,N_6926);
nor U8205 (N_8205,N_7482,N_7203);
nor U8206 (N_8206,N_7361,N_6777);
nand U8207 (N_8207,N_6883,N_7263);
or U8208 (N_8208,N_7146,N_7316);
xor U8209 (N_8209,N_7351,N_7070);
and U8210 (N_8210,N_7008,N_7096);
xor U8211 (N_8211,N_7238,N_7024);
nor U8212 (N_8212,N_6918,N_7109);
nand U8213 (N_8213,N_7213,N_7154);
nand U8214 (N_8214,N_7048,N_6812);
or U8215 (N_8215,N_7272,N_7187);
and U8216 (N_8216,N_6835,N_7012);
nand U8217 (N_8217,N_7227,N_7393);
nor U8218 (N_8218,N_6764,N_6805);
nand U8219 (N_8219,N_7398,N_7232);
xnor U8220 (N_8220,N_6822,N_7181);
nand U8221 (N_8221,N_7218,N_7498);
xnor U8222 (N_8222,N_7450,N_7221);
nand U8223 (N_8223,N_6944,N_7454);
and U8224 (N_8224,N_6875,N_6999);
nand U8225 (N_8225,N_7292,N_7277);
nor U8226 (N_8226,N_7178,N_6753);
and U8227 (N_8227,N_7275,N_6788);
or U8228 (N_8228,N_7274,N_7408);
nand U8229 (N_8229,N_7207,N_6912);
and U8230 (N_8230,N_7171,N_6777);
and U8231 (N_8231,N_7329,N_7386);
xor U8232 (N_8232,N_7223,N_7031);
nor U8233 (N_8233,N_7167,N_7015);
or U8234 (N_8234,N_7465,N_7087);
or U8235 (N_8235,N_6917,N_6805);
xnor U8236 (N_8236,N_6919,N_6973);
nor U8237 (N_8237,N_7066,N_7069);
or U8238 (N_8238,N_7326,N_7191);
xor U8239 (N_8239,N_6881,N_7112);
nand U8240 (N_8240,N_6977,N_6866);
or U8241 (N_8241,N_7186,N_7378);
or U8242 (N_8242,N_7082,N_6752);
xor U8243 (N_8243,N_7390,N_6771);
nor U8244 (N_8244,N_6989,N_7478);
and U8245 (N_8245,N_7283,N_7496);
and U8246 (N_8246,N_7448,N_7019);
xnor U8247 (N_8247,N_7104,N_7497);
nor U8248 (N_8248,N_7437,N_6776);
and U8249 (N_8249,N_7218,N_7234);
nor U8250 (N_8250,N_7969,N_7670);
nor U8251 (N_8251,N_8040,N_8139);
and U8252 (N_8252,N_7783,N_7957);
nand U8253 (N_8253,N_7741,N_7620);
or U8254 (N_8254,N_7602,N_7667);
or U8255 (N_8255,N_7572,N_7764);
nand U8256 (N_8256,N_8057,N_8121);
xnor U8257 (N_8257,N_7818,N_7575);
xnor U8258 (N_8258,N_7734,N_8138);
or U8259 (N_8259,N_7862,N_7746);
and U8260 (N_8260,N_8036,N_8095);
nand U8261 (N_8261,N_7593,N_8016);
xor U8262 (N_8262,N_7832,N_7612);
xor U8263 (N_8263,N_7518,N_8226);
nor U8264 (N_8264,N_7562,N_7574);
xor U8265 (N_8265,N_7597,N_8179);
nand U8266 (N_8266,N_7999,N_7683);
nand U8267 (N_8267,N_7504,N_7586);
or U8268 (N_8268,N_7619,N_8010);
or U8269 (N_8269,N_7679,N_7879);
or U8270 (N_8270,N_7827,N_7974);
and U8271 (N_8271,N_7881,N_8155);
nor U8272 (N_8272,N_7585,N_8200);
and U8273 (N_8273,N_7945,N_7660);
or U8274 (N_8274,N_8160,N_7615);
nor U8275 (N_8275,N_7856,N_7591);
nor U8276 (N_8276,N_7692,N_7748);
nor U8277 (N_8277,N_8175,N_7539);
nor U8278 (N_8278,N_7680,N_7896);
nand U8279 (N_8279,N_7942,N_8210);
or U8280 (N_8280,N_8242,N_7738);
nand U8281 (N_8281,N_7844,N_8053);
xnor U8282 (N_8282,N_7808,N_8135);
and U8283 (N_8283,N_7530,N_7689);
or U8284 (N_8284,N_7566,N_8074);
xnor U8285 (N_8285,N_7702,N_7824);
or U8286 (N_8286,N_8034,N_7962);
or U8287 (N_8287,N_7637,N_8117);
nor U8288 (N_8288,N_7907,N_8007);
or U8289 (N_8289,N_8233,N_7654);
nand U8290 (N_8290,N_7920,N_7891);
and U8291 (N_8291,N_7848,N_7737);
nand U8292 (N_8292,N_8174,N_7947);
and U8293 (N_8293,N_7893,N_7977);
or U8294 (N_8294,N_7669,N_7581);
xnor U8295 (N_8295,N_7739,N_8209);
nand U8296 (N_8296,N_7937,N_7554);
and U8297 (N_8297,N_7954,N_7656);
nand U8298 (N_8298,N_7605,N_7727);
or U8299 (N_8299,N_8248,N_7763);
nor U8300 (N_8300,N_7529,N_7772);
nand U8301 (N_8301,N_8140,N_7754);
nand U8302 (N_8302,N_7665,N_8249);
nand U8303 (N_8303,N_7789,N_7646);
nand U8304 (N_8304,N_7743,N_8008);
nand U8305 (N_8305,N_7956,N_7917);
xnor U8306 (N_8306,N_7666,N_7998);
nor U8307 (N_8307,N_7528,N_7625);
nand U8308 (N_8308,N_7798,N_8187);
nand U8309 (N_8309,N_8019,N_7794);
or U8310 (N_8310,N_8212,N_8230);
and U8311 (N_8311,N_8064,N_7836);
nor U8312 (N_8312,N_7671,N_7939);
and U8313 (N_8313,N_7976,N_7521);
or U8314 (N_8314,N_8079,N_7870);
nor U8315 (N_8315,N_7600,N_7613);
nor U8316 (N_8316,N_7708,N_7935);
xnor U8317 (N_8317,N_8213,N_7983);
xnor U8318 (N_8318,N_7551,N_8167);
nor U8319 (N_8319,N_7845,N_7765);
nor U8320 (N_8320,N_8159,N_7672);
xor U8321 (N_8321,N_7548,N_7801);
or U8322 (N_8322,N_7747,N_7797);
and U8323 (N_8323,N_8136,N_8011);
or U8324 (N_8324,N_7880,N_8203);
or U8325 (N_8325,N_8189,N_7690);
or U8326 (N_8326,N_7626,N_8129);
xor U8327 (N_8327,N_7915,N_7547);
nand U8328 (N_8328,N_8003,N_8001);
nor U8329 (N_8329,N_8086,N_7886);
and U8330 (N_8330,N_7859,N_7517);
nand U8331 (N_8331,N_8142,N_7809);
nand U8332 (N_8332,N_7505,N_8055);
nor U8333 (N_8333,N_7614,N_7767);
xnor U8334 (N_8334,N_8090,N_7898);
nor U8335 (N_8335,N_8087,N_7930);
nand U8336 (N_8336,N_7507,N_8130);
or U8337 (N_8337,N_8165,N_7698);
nand U8338 (N_8338,N_7584,N_8024);
xor U8339 (N_8339,N_7636,N_7750);
xnor U8340 (N_8340,N_7780,N_7676);
xnor U8341 (N_8341,N_7972,N_7872);
or U8342 (N_8342,N_8247,N_8186);
xnor U8343 (N_8343,N_8097,N_7904);
and U8344 (N_8344,N_7519,N_7609);
nor U8345 (N_8345,N_8178,N_7580);
nand U8346 (N_8346,N_7569,N_8206);
nor U8347 (N_8347,N_7531,N_8126);
or U8348 (N_8348,N_7823,N_7618);
and U8349 (N_8349,N_7661,N_7647);
or U8350 (N_8350,N_7663,N_7903);
and U8351 (N_8351,N_8150,N_8228);
xnor U8352 (N_8352,N_7892,N_8141);
nor U8353 (N_8353,N_8225,N_7784);
or U8354 (N_8354,N_8050,N_8092);
nand U8355 (N_8355,N_8191,N_8052);
nor U8356 (N_8356,N_7526,N_7802);
xnor U8357 (N_8357,N_8112,N_7653);
xor U8358 (N_8358,N_7829,N_8093);
nor U8359 (N_8359,N_7837,N_7641);
and U8360 (N_8360,N_8182,N_7555);
xor U8361 (N_8361,N_8152,N_7833);
xnor U8362 (N_8362,N_7659,N_7979);
or U8363 (N_8363,N_7697,N_7674);
and U8364 (N_8364,N_7577,N_7851);
or U8365 (N_8365,N_7598,N_7968);
or U8366 (N_8366,N_8239,N_7986);
xor U8367 (N_8367,N_7911,N_7677);
xnor U8368 (N_8368,N_8025,N_7686);
nor U8369 (N_8369,N_8127,N_8176);
nor U8370 (N_8370,N_7673,N_8070);
xor U8371 (N_8371,N_7816,N_8056);
or U8372 (N_8372,N_8188,N_8198);
and U8373 (N_8373,N_7889,N_8113);
nand U8374 (N_8374,N_7715,N_7515);
nand U8375 (N_8375,N_7821,N_8134);
nand U8376 (N_8376,N_8017,N_7616);
and U8377 (N_8377,N_8066,N_7869);
nor U8378 (N_8378,N_7604,N_8207);
nor U8379 (N_8379,N_7759,N_7643);
and U8380 (N_8380,N_8168,N_8161);
nor U8381 (N_8381,N_8243,N_7536);
and U8382 (N_8382,N_8067,N_8035);
xnor U8383 (N_8383,N_8021,N_7792);
nand U8384 (N_8384,N_8109,N_8043);
and U8385 (N_8385,N_8088,N_7556);
nor U8386 (N_8386,N_7768,N_7685);
xnor U8387 (N_8387,N_7963,N_7980);
nand U8388 (N_8388,N_7902,N_8103);
and U8389 (N_8389,N_8098,N_7694);
nand U8390 (N_8390,N_7843,N_7894);
nor U8391 (N_8391,N_8148,N_7941);
and U8392 (N_8392,N_8143,N_7841);
and U8393 (N_8393,N_7776,N_7560);
xor U8394 (N_8394,N_7860,N_7819);
xnor U8395 (N_8395,N_8085,N_8202);
or U8396 (N_8396,N_8221,N_7914);
nor U8397 (N_8397,N_7779,N_7966);
nor U8398 (N_8398,N_7924,N_7693);
nand U8399 (N_8399,N_8089,N_7728);
nor U8400 (N_8400,N_7725,N_7766);
and U8401 (N_8401,N_7731,N_7807);
xor U8402 (N_8402,N_7929,N_8124);
or U8403 (N_8403,N_7944,N_8028);
or U8404 (N_8404,N_7631,N_8125);
nand U8405 (N_8405,N_7813,N_7971);
nor U8406 (N_8406,N_8231,N_7961);
xnor U8407 (N_8407,N_8235,N_8123);
and U8408 (N_8408,N_7897,N_7559);
xnor U8409 (N_8409,N_7687,N_8084);
or U8410 (N_8410,N_8049,N_8119);
nor U8411 (N_8411,N_8022,N_7847);
or U8412 (N_8412,N_7921,N_8193);
and U8413 (N_8413,N_8006,N_7812);
xnor U8414 (N_8414,N_8118,N_7707);
nand U8415 (N_8415,N_8104,N_8208);
and U8416 (N_8416,N_7928,N_8216);
or U8417 (N_8417,N_7988,N_8151);
and U8418 (N_8418,N_7608,N_7740);
nor U8419 (N_8419,N_8059,N_7975);
nand U8420 (N_8420,N_8111,N_7887);
xor U8421 (N_8421,N_7711,N_7934);
nand U8422 (N_8422,N_7714,N_8048);
xor U8423 (N_8423,N_7567,N_8038);
nand U8424 (N_8424,N_7716,N_7542);
and U8425 (N_8425,N_7730,N_8027);
xor U8426 (N_8426,N_7854,N_7884);
nor U8427 (N_8427,N_7733,N_7516);
xnor U8428 (N_8428,N_7868,N_8149);
and U8429 (N_8429,N_8154,N_8180);
nand U8430 (N_8430,N_8169,N_7788);
or U8431 (N_8431,N_7630,N_7997);
xor U8432 (N_8432,N_7781,N_8137);
xor U8433 (N_8433,N_7540,N_7511);
xnor U8434 (N_8434,N_8133,N_8030);
nand U8435 (N_8435,N_7790,N_7564);
nand U8436 (N_8436,N_7503,N_8194);
xor U8437 (N_8437,N_7838,N_7512);
nor U8438 (N_8438,N_7583,N_8100);
nand U8439 (N_8439,N_8181,N_7657);
and U8440 (N_8440,N_7900,N_7861);
xor U8441 (N_8441,N_7965,N_8246);
or U8442 (N_8442,N_7796,N_7610);
or U8443 (N_8443,N_7948,N_7596);
and U8444 (N_8444,N_7927,N_8044);
and U8445 (N_8445,N_8014,N_7640);
nand U8446 (N_8446,N_7918,N_7570);
nor U8447 (N_8447,N_7595,N_8163);
nand U8448 (N_8448,N_8042,N_8238);
nor U8449 (N_8449,N_7546,N_8114);
or U8450 (N_8450,N_8076,N_7946);
nor U8451 (N_8451,N_8241,N_8031);
nor U8452 (N_8452,N_8217,N_7991);
nor U8453 (N_8453,N_7787,N_7960);
xnor U8454 (N_8454,N_8018,N_7949);
and U8455 (N_8455,N_7751,N_7878);
or U8456 (N_8456,N_8106,N_7744);
or U8457 (N_8457,N_7825,N_7658);
and U8458 (N_8458,N_7933,N_8131);
or U8459 (N_8459,N_7502,N_8071);
nand U8460 (N_8460,N_7877,N_7817);
or U8461 (N_8461,N_7905,N_7814);
nand U8462 (N_8462,N_7916,N_7565);
xnor U8463 (N_8463,N_7705,N_7645);
nor U8464 (N_8464,N_8144,N_8156);
xnor U8465 (N_8465,N_7782,N_7840);
nor U8466 (N_8466,N_7664,N_7992);
xnor U8467 (N_8467,N_8062,N_7996);
or U8468 (N_8468,N_8110,N_7508);
and U8469 (N_8469,N_7982,N_7682);
and U8470 (N_8470,N_7799,N_7717);
xnor U8471 (N_8471,N_7770,N_7831);
nor U8472 (N_8472,N_8009,N_7793);
or U8473 (N_8473,N_7883,N_7558);
nand U8474 (N_8474,N_8046,N_7958);
nand U8475 (N_8475,N_7644,N_7775);
nor U8476 (N_8476,N_7650,N_7822);
nor U8477 (N_8477,N_8058,N_7882);
nor U8478 (N_8478,N_8220,N_7745);
and U8479 (N_8479,N_8075,N_8224);
xnor U8480 (N_8480,N_7773,N_7786);
nor U8481 (N_8481,N_7699,N_7970);
or U8482 (N_8482,N_7864,N_7501);
and U8483 (N_8483,N_7795,N_7622);
xnor U8484 (N_8484,N_8211,N_7681);
and U8485 (N_8485,N_7695,N_8177);
xor U8486 (N_8486,N_8013,N_8039);
and U8487 (N_8487,N_8229,N_7756);
nor U8488 (N_8488,N_7815,N_7888);
nand U8489 (N_8489,N_7810,N_7749);
or U8490 (N_8490,N_8236,N_8068);
xor U8491 (N_8491,N_7820,N_8101);
nor U8492 (N_8492,N_8065,N_8195);
xor U8493 (N_8493,N_7729,N_7621);
and U8494 (N_8494,N_7876,N_8227);
nand U8495 (N_8495,N_7774,N_7757);
nor U8496 (N_8496,N_7651,N_7668);
or U8497 (N_8497,N_7603,N_7855);
and U8498 (N_8498,N_7785,N_7599);
xor U8499 (N_8499,N_7696,N_8107);
nor U8500 (N_8500,N_7710,N_7846);
or U8501 (N_8501,N_7722,N_8061);
and U8502 (N_8502,N_8094,N_7828);
and U8503 (N_8503,N_7735,N_8072);
nor U8504 (N_8504,N_7834,N_7761);
and U8505 (N_8505,N_8115,N_8041);
xor U8506 (N_8506,N_8060,N_7912);
nor U8507 (N_8507,N_8015,N_8128);
xnor U8508 (N_8508,N_7811,N_7760);
or U8509 (N_8509,N_7805,N_7901);
nor U8510 (N_8510,N_7525,N_8096);
and U8511 (N_8511,N_7545,N_8120);
and U8512 (N_8512,N_7557,N_7926);
and U8513 (N_8513,N_7849,N_7940);
and U8514 (N_8514,N_7895,N_7753);
nand U8515 (N_8515,N_8215,N_7535);
nor U8516 (N_8516,N_7541,N_7588);
nand U8517 (N_8517,N_7549,N_7842);
nor U8518 (N_8518,N_8020,N_7804);
nor U8519 (N_8519,N_7678,N_7606);
nor U8520 (N_8520,N_7544,N_7987);
or U8521 (N_8521,N_7704,N_8205);
nor U8522 (N_8522,N_7908,N_7628);
and U8523 (N_8523,N_8132,N_7984);
nor U8524 (N_8524,N_7573,N_7919);
nand U8525 (N_8525,N_8077,N_7985);
xor U8526 (N_8526,N_7720,N_8196);
nor U8527 (N_8527,N_7662,N_7524);
xor U8528 (N_8528,N_7839,N_7629);
or U8529 (N_8529,N_7803,N_8172);
and U8530 (N_8530,N_7642,N_7709);
xnor U8531 (N_8531,N_8078,N_7913);
nand U8532 (N_8532,N_7553,N_8170);
xor U8533 (N_8533,N_7527,N_7590);
xor U8534 (N_8534,N_7931,N_7852);
nor U8535 (N_8535,N_8219,N_8045);
nor U8536 (N_8536,N_7552,N_7617);
or U8537 (N_8537,N_7938,N_8051);
xnor U8538 (N_8538,N_8029,N_8237);
or U8539 (N_8539,N_7955,N_8083);
or U8540 (N_8540,N_7624,N_7778);
nand U8541 (N_8541,N_7568,N_7899);
nand U8542 (N_8542,N_7655,N_7726);
and U8543 (N_8543,N_7885,N_7700);
and U8544 (N_8544,N_7995,N_7706);
nand U8545 (N_8545,N_8166,N_8245);
and U8546 (N_8546,N_8012,N_7993);
or U8547 (N_8547,N_7721,N_7874);
xor U8548 (N_8548,N_7967,N_8145);
nor U8549 (N_8549,N_8171,N_7777);
nand U8550 (N_8550,N_7871,N_7830);
nand U8551 (N_8551,N_7943,N_7863);
nor U8552 (N_8552,N_8184,N_7648);
nor U8553 (N_8553,N_7981,N_8232);
and U8554 (N_8554,N_8004,N_7684);
nor U8555 (N_8555,N_7951,N_7762);
xor U8556 (N_8556,N_7910,N_7959);
or U8557 (N_8557,N_8032,N_7533);
nand U8558 (N_8558,N_7712,N_8240);
or U8559 (N_8559,N_7989,N_8037);
or U8560 (N_8560,N_7538,N_8185);
and U8561 (N_8561,N_7755,N_7800);
nor U8562 (N_8562,N_7925,N_7582);
xnor U8563 (N_8563,N_8080,N_8063);
nor U8564 (N_8564,N_7953,N_7537);
nand U8565 (N_8565,N_7649,N_8222);
xor U8566 (N_8566,N_8054,N_7532);
nand U8567 (N_8567,N_7857,N_7994);
nor U8568 (N_8568,N_7623,N_7742);
nand U8569 (N_8569,N_8199,N_7550);
and U8570 (N_8570,N_7506,N_7633);
and U8571 (N_8571,N_8214,N_7858);
and U8572 (N_8572,N_7522,N_7513);
and U8573 (N_8573,N_7736,N_7701);
or U8574 (N_8574,N_8164,N_8192);
nand U8575 (N_8575,N_7688,N_7923);
or U8576 (N_8576,N_7835,N_7826);
nand U8577 (N_8577,N_8023,N_8201);
and U8578 (N_8578,N_8091,N_7634);
nand U8579 (N_8579,N_7732,N_8047);
nor U8580 (N_8580,N_7594,N_7853);
nand U8581 (N_8581,N_7866,N_8069);
or U8582 (N_8582,N_7520,N_8002);
nand U8583 (N_8583,N_8158,N_7769);
nand U8584 (N_8584,N_7713,N_7571);
xnor U8585 (N_8585,N_8146,N_8244);
nor U8586 (N_8586,N_8218,N_7791);
nor U8587 (N_8587,N_8204,N_7638);
nand U8588 (N_8588,N_8122,N_8102);
nor U8589 (N_8589,N_7703,N_7514);
nor U8590 (N_8590,N_7865,N_7964);
or U8591 (N_8591,N_7906,N_8073);
xnor U8592 (N_8592,N_7850,N_7875);
nor U8593 (N_8593,N_7932,N_7867);
nor U8594 (N_8594,N_7607,N_7890);
nor U8595 (N_8595,N_7601,N_8026);
nor U8596 (N_8596,N_7723,N_7509);
and U8597 (N_8597,N_7579,N_8082);
nor U8598 (N_8598,N_7543,N_7936);
nand U8599 (N_8599,N_7627,N_7611);
or U8600 (N_8600,N_7978,N_7578);
nor U8601 (N_8601,N_7752,N_7561);
xnor U8602 (N_8602,N_7510,N_8157);
or U8603 (N_8603,N_8153,N_7952);
and U8604 (N_8604,N_8162,N_7909);
and U8605 (N_8605,N_7652,N_7500);
and U8606 (N_8606,N_7758,N_7806);
nand U8607 (N_8607,N_8005,N_8105);
nand U8608 (N_8608,N_8223,N_8183);
nand U8609 (N_8609,N_7639,N_8116);
nand U8610 (N_8610,N_8081,N_8108);
or U8611 (N_8611,N_7691,N_8190);
and U8612 (N_8612,N_7675,N_7632);
or U8613 (N_8613,N_7563,N_8234);
xnor U8614 (N_8614,N_7950,N_7576);
and U8615 (N_8615,N_7592,N_8197);
nor U8616 (N_8616,N_8147,N_7718);
nand U8617 (N_8617,N_7635,N_7724);
xnor U8618 (N_8618,N_8099,N_7990);
or U8619 (N_8619,N_8173,N_7873);
nand U8620 (N_8620,N_8000,N_7523);
nor U8621 (N_8621,N_7973,N_8033);
and U8622 (N_8622,N_7922,N_7771);
xor U8623 (N_8623,N_7719,N_7587);
or U8624 (N_8624,N_7589,N_7534);
xnor U8625 (N_8625,N_8133,N_7724);
or U8626 (N_8626,N_7674,N_7824);
and U8627 (N_8627,N_8221,N_7917);
nor U8628 (N_8628,N_7692,N_8047);
or U8629 (N_8629,N_7597,N_8121);
and U8630 (N_8630,N_7858,N_7779);
nor U8631 (N_8631,N_7915,N_7563);
nor U8632 (N_8632,N_7531,N_8204);
and U8633 (N_8633,N_8098,N_7520);
xor U8634 (N_8634,N_7903,N_8099);
or U8635 (N_8635,N_7775,N_7716);
xnor U8636 (N_8636,N_7638,N_8106);
nand U8637 (N_8637,N_7857,N_7732);
and U8638 (N_8638,N_7873,N_8100);
nand U8639 (N_8639,N_7882,N_7764);
nand U8640 (N_8640,N_8186,N_7532);
or U8641 (N_8641,N_7969,N_7590);
or U8642 (N_8642,N_7595,N_7670);
xor U8643 (N_8643,N_7900,N_7740);
nand U8644 (N_8644,N_7529,N_7637);
xnor U8645 (N_8645,N_7771,N_8005);
nand U8646 (N_8646,N_8148,N_7551);
xnor U8647 (N_8647,N_8111,N_7845);
nor U8648 (N_8648,N_7895,N_7866);
nor U8649 (N_8649,N_8159,N_7915);
nor U8650 (N_8650,N_7841,N_7660);
or U8651 (N_8651,N_8077,N_7714);
xnor U8652 (N_8652,N_7908,N_8105);
and U8653 (N_8653,N_8218,N_7507);
and U8654 (N_8654,N_7809,N_7979);
nand U8655 (N_8655,N_8142,N_7551);
or U8656 (N_8656,N_7938,N_7982);
or U8657 (N_8657,N_7560,N_7656);
xnor U8658 (N_8658,N_7852,N_8035);
nor U8659 (N_8659,N_7538,N_8124);
xor U8660 (N_8660,N_7558,N_7546);
or U8661 (N_8661,N_7940,N_7617);
xor U8662 (N_8662,N_8193,N_7631);
nor U8663 (N_8663,N_7907,N_7960);
xnor U8664 (N_8664,N_7784,N_7646);
nor U8665 (N_8665,N_7525,N_8084);
xnor U8666 (N_8666,N_8105,N_7942);
or U8667 (N_8667,N_7990,N_7737);
xnor U8668 (N_8668,N_8166,N_7765);
xnor U8669 (N_8669,N_7951,N_7649);
nand U8670 (N_8670,N_7858,N_7624);
xnor U8671 (N_8671,N_8241,N_7899);
and U8672 (N_8672,N_7655,N_7676);
nand U8673 (N_8673,N_7934,N_7873);
or U8674 (N_8674,N_7536,N_7775);
nor U8675 (N_8675,N_7532,N_7903);
and U8676 (N_8676,N_7790,N_7811);
or U8677 (N_8677,N_7632,N_7861);
nor U8678 (N_8678,N_7870,N_8191);
and U8679 (N_8679,N_7705,N_7681);
and U8680 (N_8680,N_7632,N_7794);
and U8681 (N_8681,N_8138,N_7515);
and U8682 (N_8682,N_7750,N_8239);
or U8683 (N_8683,N_7854,N_7687);
and U8684 (N_8684,N_8145,N_8168);
nand U8685 (N_8685,N_7707,N_7961);
and U8686 (N_8686,N_7874,N_8205);
xnor U8687 (N_8687,N_7889,N_7918);
xor U8688 (N_8688,N_7676,N_7897);
xnor U8689 (N_8689,N_7732,N_7962);
xor U8690 (N_8690,N_8053,N_8139);
nor U8691 (N_8691,N_7822,N_7755);
and U8692 (N_8692,N_8051,N_7577);
or U8693 (N_8693,N_7604,N_7617);
nand U8694 (N_8694,N_7527,N_8064);
and U8695 (N_8695,N_7917,N_7669);
and U8696 (N_8696,N_8180,N_7635);
or U8697 (N_8697,N_7943,N_7525);
and U8698 (N_8698,N_7689,N_7521);
and U8699 (N_8699,N_7659,N_7948);
and U8700 (N_8700,N_8097,N_7713);
and U8701 (N_8701,N_7727,N_8033);
nand U8702 (N_8702,N_7695,N_8138);
or U8703 (N_8703,N_8149,N_7768);
nor U8704 (N_8704,N_7568,N_7848);
and U8705 (N_8705,N_7687,N_7690);
nor U8706 (N_8706,N_7649,N_7507);
or U8707 (N_8707,N_8113,N_7643);
and U8708 (N_8708,N_7803,N_7671);
nor U8709 (N_8709,N_8241,N_8128);
nand U8710 (N_8710,N_7562,N_7869);
nand U8711 (N_8711,N_7662,N_8121);
and U8712 (N_8712,N_7749,N_7802);
nor U8713 (N_8713,N_8235,N_8092);
nor U8714 (N_8714,N_7655,N_7869);
nor U8715 (N_8715,N_8149,N_8215);
nand U8716 (N_8716,N_7577,N_7702);
nor U8717 (N_8717,N_7855,N_7551);
xor U8718 (N_8718,N_7925,N_7610);
nor U8719 (N_8719,N_7841,N_7563);
and U8720 (N_8720,N_8063,N_7915);
and U8721 (N_8721,N_7712,N_8142);
xor U8722 (N_8722,N_7547,N_7927);
xnor U8723 (N_8723,N_7773,N_8125);
or U8724 (N_8724,N_7955,N_7901);
xnor U8725 (N_8725,N_7684,N_7961);
or U8726 (N_8726,N_8081,N_7517);
and U8727 (N_8727,N_7522,N_7585);
nor U8728 (N_8728,N_7716,N_8236);
and U8729 (N_8729,N_7814,N_7811);
xor U8730 (N_8730,N_7504,N_8179);
xnor U8731 (N_8731,N_8087,N_7795);
nand U8732 (N_8732,N_7673,N_8024);
xnor U8733 (N_8733,N_8038,N_7955);
or U8734 (N_8734,N_7656,N_7582);
and U8735 (N_8735,N_7986,N_7555);
or U8736 (N_8736,N_8171,N_8015);
xor U8737 (N_8737,N_7796,N_8191);
and U8738 (N_8738,N_7641,N_7584);
and U8739 (N_8739,N_7852,N_7808);
or U8740 (N_8740,N_7702,N_7724);
or U8741 (N_8741,N_7857,N_7684);
nor U8742 (N_8742,N_8098,N_7653);
and U8743 (N_8743,N_7806,N_7589);
nor U8744 (N_8744,N_7991,N_7931);
and U8745 (N_8745,N_8236,N_7746);
nand U8746 (N_8746,N_7946,N_8086);
nor U8747 (N_8747,N_7887,N_7632);
and U8748 (N_8748,N_7681,N_7742);
and U8749 (N_8749,N_7843,N_8065);
and U8750 (N_8750,N_7680,N_7803);
nand U8751 (N_8751,N_7993,N_8028);
xnor U8752 (N_8752,N_8018,N_7841);
nor U8753 (N_8753,N_7859,N_8157);
or U8754 (N_8754,N_7523,N_8150);
or U8755 (N_8755,N_7588,N_8144);
nor U8756 (N_8756,N_8241,N_7907);
xnor U8757 (N_8757,N_8166,N_7960);
nor U8758 (N_8758,N_8105,N_8015);
and U8759 (N_8759,N_7905,N_7626);
and U8760 (N_8760,N_8208,N_7590);
and U8761 (N_8761,N_7899,N_7871);
nand U8762 (N_8762,N_7621,N_7855);
nand U8763 (N_8763,N_8247,N_7911);
and U8764 (N_8764,N_7871,N_7724);
and U8765 (N_8765,N_7662,N_7999);
nand U8766 (N_8766,N_7845,N_8039);
nand U8767 (N_8767,N_7638,N_7737);
and U8768 (N_8768,N_7836,N_8189);
nand U8769 (N_8769,N_8210,N_7648);
xnor U8770 (N_8770,N_8062,N_7715);
nor U8771 (N_8771,N_7650,N_8039);
xor U8772 (N_8772,N_8170,N_7976);
and U8773 (N_8773,N_7541,N_7916);
nor U8774 (N_8774,N_7629,N_7971);
and U8775 (N_8775,N_7675,N_7952);
and U8776 (N_8776,N_7654,N_7650);
and U8777 (N_8777,N_8112,N_7737);
nand U8778 (N_8778,N_8075,N_8161);
xnor U8779 (N_8779,N_8017,N_7813);
nand U8780 (N_8780,N_8128,N_8022);
xor U8781 (N_8781,N_8134,N_8183);
xor U8782 (N_8782,N_7778,N_7621);
xnor U8783 (N_8783,N_8232,N_7640);
nor U8784 (N_8784,N_7571,N_7863);
or U8785 (N_8785,N_8075,N_7676);
and U8786 (N_8786,N_7922,N_7882);
nor U8787 (N_8787,N_8166,N_8039);
or U8788 (N_8788,N_8068,N_7695);
xor U8789 (N_8789,N_7529,N_8041);
or U8790 (N_8790,N_7684,N_7867);
xor U8791 (N_8791,N_8045,N_7816);
or U8792 (N_8792,N_8105,N_8247);
and U8793 (N_8793,N_7986,N_7625);
xnor U8794 (N_8794,N_7502,N_7723);
nand U8795 (N_8795,N_7557,N_7641);
nand U8796 (N_8796,N_7650,N_8048);
xor U8797 (N_8797,N_8031,N_8113);
nor U8798 (N_8798,N_7880,N_8141);
xnor U8799 (N_8799,N_7948,N_7828);
xnor U8800 (N_8800,N_8016,N_7912);
xnor U8801 (N_8801,N_7587,N_7574);
and U8802 (N_8802,N_7510,N_7823);
nor U8803 (N_8803,N_8011,N_7625);
nor U8804 (N_8804,N_7739,N_8110);
xnor U8805 (N_8805,N_8011,N_8096);
or U8806 (N_8806,N_8245,N_8010);
and U8807 (N_8807,N_8072,N_7906);
nand U8808 (N_8808,N_7708,N_7857);
nand U8809 (N_8809,N_8138,N_8071);
or U8810 (N_8810,N_8126,N_7775);
xnor U8811 (N_8811,N_7673,N_8189);
and U8812 (N_8812,N_7664,N_7953);
and U8813 (N_8813,N_7901,N_7510);
nand U8814 (N_8814,N_7956,N_7787);
nor U8815 (N_8815,N_8033,N_7725);
xor U8816 (N_8816,N_8062,N_8054);
xor U8817 (N_8817,N_7904,N_7961);
or U8818 (N_8818,N_7627,N_8023);
and U8819 (N_8819,N_8184,N_7618);
xnor U8820 (N_8820,N_7799,N_8111);
nor U8821 (N_8821,N_7611,N_7874);
xnor U8822 (N_8822,N_7557,N_8110);
xnor U8823 (N_8823,N_7687,N_8094);
and U8824 (N_8824,N_7689,N_7837);
xor U8825 (N_8825,N_7661,N_8191);
nand U8826 (N_8826,N_8196,N_7691);
xor U8827 (N_8827,N_7563,N_7518);
or U8828 (N_8828,N_7883,N_8119);
and U8829 (N_8829,N_7641,N_8179);
nand U8830 (N_8830,N_8155,N_7961);
nand U8831 (N_8831,N_8074,N_8190);
xnor U8832 (N_8832,N_7626,N_7712);
or U8833 (N_8833,N_8125,N_7537);
and U8834 (N_8834,N_7699,N_7670);
xnor U8835 (N_8835,N_7931,N_8049);
and U8836 (N_8836,N_7950,N_7555);
nand U8837 (N_8837,N_8036,N_7525);
xnor U8838 (N_8838,N_8004,N_7832);
and U8839 (N_8839,N_7985,N_7813);
nand U8840 (N_8840,N_8208,N_8154);
or U8841 (N_8841,N_7900,N_7560);
xnor U8842 (N_8842,N_8058,N_7643);
nor U8843 (N_8843,N_8174,N_7678);
and U8844 (N_8844,N_8181,N_7590);
or U8845 (N_8845,N_8043,N_7637);
nor U8846 (N_8846,N_7981,N_8036);
or U8847 (N_8847,N_7822,N_8191);
xnor U8848 (N_8848,N_8185,N_7549);
or U8849 (N_8849,N_7770,N_7726);
or U8850 (N_8850,N_8044,N_8166);
nand U8851 (N_8851,N_7606,N_7668);
or U8852 (N_8852,N_7996,N_7517);
xor U8853 (N_8853,N_7910,N_7525);
or U8854 (N_8854,N_7668,N_8091);
nor U8855 (N_8855,N_7622,N_7791);
nor U8856 (N_8856,N_7543,N_7877);
nand U8857 (N_8857,N_7795,N_7824);
and U8858 (N_8858,N_7675,N_8238);
nand U8859 (N_8859,N_7721,N_7945);
nor U8860 (N_8860,N_8189,N_8016);
or U8861 (N_8861,N_7857,N_7548);
or U8862 (N_8862,N_7627,N_7796);
nand U8863 (N_8863,N_7505,N_7582);
or U8864 (N_8864,N_7544,N_7660);
or U8865 (N_8865,N_8200,N_7890);
nor U8866 (N_8866,N_8239,N_8157);
nor U8867 (N_8867,N_7757,N_7926);
or U8868 (N_8868,N_7577,N_8184);
nand U8869 (N_8869,N_8191,N_7510);
nand U8870 (N_8870,N_7870,N_8077);
or U8871 (N_8871,N_8147,N_8082);
nand U8872 (N_8872,N_7652,N_8057);
nor U8873 (N_8873,N_7885,N_7758);
nand U8874 (N_8874,N_7730,N_8050);
nand U8875 (N_8875,N_8043,N_7872);
nand U8876 (N_8876,N_7954,N_8180);
nand U8877 (N_8877,N_7596,N_7646);
nand U8878 (N_8878,N_7636,N_7710);
or U8879 (N_8879,N_8193,N_7790);
or U8880 (N_8880,N_7857,N_7570);
xnor U8881 (N_8881,N_7782,N_7608);
nand U8882 (N_8882,N_7577,N_7667);
and U8883 (N_8883,N_7603,N_7579);
xor U8884 (N_8884,N_7620,N_8036);
or U8885 (N_8885,N_7535,N_7564);
nor U8886 (N_8886,N_7671,N_7909);
nand U8887 (N_8887,N_8147,N_7919);
nand U8888 (N_8888,N_7807,N_7839);
nor U8889 (N_8889,N_7993,N_7596);
xnor U8890 (N_8890,N_7515,N_7695);
nor U8891 (N_8891,N_8158,N_7792);
nor U8892 (N_8892,N_8055,N_7881);
nor U8893 (N_8893,N_8189,N_8054);
or U8894 (N_8894,N_8059,N_7754);
or U8895 (N_8895,N_8130,N_7652);
xor U8896 (N_8896,N_7503,N_7769);
xor U8897 (N_8897,N_7699,N_8119);
or U8898 (N_8898,N_8133,N_7526);
nor U8899 (N_8899,N_7854,N_8074);
or U8900 (N_8900,N_8041,N_7683);
nand U8901 (N_8901,N_8216,N_7611);
nor U8902 (N_8902,N_7700,N_7926);
nor U8903 (N_8903,N_8146,N_7594);
and U8904 (N_8904,N_7571,N_8027);
or U8905 (N_8905,N_8124,N_7673);
nand U8906 (N_8906,N_7701,N_8002);
xnor U8907 (N_8907,N_7648,N_8134);
nor U8908 (N_8908,N_8161,N_8249);
xnor U8909 (N_8909,N_7530,N_7675);
and U8910 (N_8910,N_8056,N_7858);
nand U8911 (N_8911,N_7862,N_7799);
or U8912 (N_8912,N_7559,N_7851);
nand U8913 (N_8913,N_7586,N_7809);
nor U8914 (N_8914,N_8020,N_7598);
xnor U8915 (N_8915,N_8123,N_7906);
nor U8916 (N_8916,N_7545,N_8116);
nand U8917 (N_8917,N_7508,N_7971);
and U8918 (N_8918,N_8004,N_7942);
or U8919 (N_8919,N_8026,N_7788);
xnor U8920 (N_8920,N_8039,N_7662);
xor U8921 (N_8921,N_7719,N_7505);
and U8922 (N_8922,N_7989,N_7852);
and U8923 (N_8923,N_7668,N_8039);
or U8924 (N_8924,N_7579,N_7697);
nand U8925 (N_8925,N_7633,N_7806);
and U8926 (N_8926,N_7562,N_7884);
nor U8927 (N_8927,N_8221,N_7579);
nand U8928 (N_8928,N_8000,N_8119);
and U8929 (N_8929,N_7874,N_8101);
nand U8930 (N_8930,N_7550,N_8188);
or U8931 (N_8931,N_7735,N_8132);
and U8932 (N_8932,N_8195,N_7968);
nand U8933 (N_8933,N_7910,N_7723);
xnor U8934 (N_8934,N_8163,N_7734);
nand U8935 (N_8935,N_7877,N_8108);
xnor U8936 (N_8936,N_7744,N_8191);
nand U8937 (N_8937,N_7766,N_7765);
xor U8938 (N_8938,N_7563,N_8094);
and U8939 (N_8939,N_7895,N_8187);
nor U8940 (N_8940,N_8022,N_7522);
nand U8941 (N_8941,N_8178,N_8075);
and U8942 (N_8942,N_7624,N_7912);
xor U8943 (N_8943,N_7805,N_7698);
or U8944 (N_8944,N_8050,N_7711);
and U8945 (N_8945,N_7598,N_8169);
or U8946 (N_8946,N_7986,N_7685);
xnor U8947 (N_8947,N_7956,N_8094);
nand U8948 (N_8948,N_8058,N_7504);
nor U8949 (N_8949,N_7776,N_7953);
nand U8950 (N_8950,N_7856,N_8007);
or U8951 (N_8951,N_8000,N_7893);
nor U8952 (N_8952,N_7567,N_7834);
nand U8953 (N_8953,N_8064,N_7925);
nor U8954 (N_8954,N_7969,N_8137);
xnor U8955 (N_8955,N_7759,N_8075);
and U8956 (N_8956,N_8034,N_8107);
nor U8957 (N_8957,N_8027,N_8010);
or U8958 (N_8958,N_8026,N_8202);
and U8959 (N_8959,N_8145,N_7722);
xor U8960 (N_8960,N_7653,N_7709);
or U8961 (N_8961,N_7806,N_8200);
nand U8962 (N_8962,N_7939,N_7974);
nand U8963 (N_8963,N_8165,N_7879);
or U8964 (N_8964,N_7718,N_8178);
nor U8965 (N_8965,N_7588,N_7858);
or U8966 (N_8966,N_7944,N_7733);
and U8967 (N_8967,N_7878,N_7910);
nand U8968 (N_8968,N_7829,N_8037);
nand U8969 (N_8969,N_7729,N_8086);
or U8970 (N_8970,N_7936,N_7984);
nand U8971 (N_8971,N_7685,N_7760);
xor U8972 (N_8972,N_7806,N_8085);
nor U8973 (N_8973,N_8054,N_7848);
and U8974 (N_8974,N_7895,N_7541);
or U8975 (N_8975,N_7941,N_7572);
xnor U8976 (N_8976,N_7532,N_7853);
xnor U8977 (N_8977,N_7842,N_7815);
nand U8978 (N_8978,N_8162,N_8206);
and U8979 (N_8979,N_8008,N_7524);
nor U8980 (N_8980,N_7896,N_7588);
or U8981 (N_8981,N_7565,N_7601);
xnor U8982 (N_8982,N_7630,N_7611);
and U8983 (N_8983,N_8074,N_7690);
and U8984 (N_8984,N_7518,N_7659);
nand U8985 (N_8985,N_7842,N_7743);
xnor U8986 (N_8986,N_7786,N_7859);
xnor U8987 (N_8987,N_7619,N_7796);
nor U8988 (N_8988,N_7893,N_7626);
nand U8989 (N_8989,N_7947,N_7841);
xnor U8990 (N_8990,N_7588,N_7607);
xor U8991 (N_8991,N_7605,N_7847);
nand U8992 (N_8992,N_8171,N_8104);
and U8993 (N_8993,N_8016,N_7583);
nand U8994 (N_8994,N_7504,N_8045);
or U8995 (N_8995,N_7944,N_7545);
nor U8996 (N_8996,N_7505,N_7996);
nand U8997 (N_8997,N_7605,N_7548);
nand U8998 (N_8998,N_7713,N_8160);
or U8999 (N_8999,N_8135,N_7621);
or U9000 (N_9000,N_8737,N_8618);
nor U9001 (N_9001,N_8800,N_8733);
or U9002 (N_9002,N_8823,N_8254);
or U9003 (N_9003,N_8730,N_8720);
xor U9004 (N_9004,N_8373,N_8963);
xnor U9005 (N_9005,N_8485,N_8389);
and U9006 (N_9006,N_8628,N_8554);
or U9007 (N_9007,N_8457,N_8679);
nor U9008 (N_9008,N_8453,N_8399);
and U9009 (N_9009,N_8342,N_8371);
and U9010 (N_9010,N_8321,N_8917);
and U9011 (N_9011,N_8636,N_8571);
nor U9012 (N_9012,N_8986,N_8871);
nand U9013 (N_9013,N_8774,N_8708);
nor U9014 (N_9014,N_8822,N_8319);
xnor U9015 (N_9015,N_8288,N_8690);
nor U9016 (N_9016,N_8482,N_8624);
nor U9017 (N_9017,N_8370,N_8567);
xnor U9018 (N_9018,N_8658,N_8763);
nand U9019 (N_9019,N_8674,N_8810);
and U9020 (N_9020,N_8384,N_8831);
xnor U9021 (N_9021,N_8606,N_8689);
nor U9022 (N_9022,N_8488,N_8285);
or U9023 (N_9023,N_8880,N_8661);
nand U9024 (N_9024,N_8335,N_8356);
or U9025 (N_9025,N_8867,N_8623);
nor U9026 (N_9026,N_8448,N_8887);
nand U9027 (N_9027,N_8341,N_8458);
or U9028 (N_9028,N_8326,N_8374);
or U9029 (N_9029,N_8723,N_8985);
nand U9030 (N_9030,N_8492,N_8475);
or U9031 (N_9031,N_8587,N_8514);
and U9032 (N_9032,N_8578,N_8447);
nor U9033 (N_9033,N_8526,N_8261);
or U9034 (N_9034,N_8836,N_8781);
xor U9035 (N_9035,N_8923,N_8675);
or U9036 (N_9036,N_8480,N_8821);
and U9037 (N_9037,N_8343,N_8385);
or U9038 (N_9038,N_8949,N_8643);
nand U9039 (N_9039,N_8420,N_8642);
and U9040 (N_9040,N_8706,N_8273);
nor U9041 (N_9041,N_8609,N_8602);
xor U9042 (N_9042,N_8264,N_8979);
nand U9043 (N_9043,N_8603,N_8421);
xor U9044 (N_9044,N_8424,N_8667);
nor U9045 (N_9045,N_8517,N_8811);
nand U9046 (N_9046,N_8664,N_8583);
xnor U9047 (N_9047,N_8255,N_8942);
or U9048 (N_9048,N_8407,N_8287);
or U9049 (N_9049,N_8864,N_8995);
nor U9050 (N_9050,N_8777,N_8964);
and U9051 (N_9051,N_8958,N_8778);
and U9052 (N_9052,N_8681,N_8316);
and U9053 (N_9053,N_8666,N_8965);
nand U9054 (N_9054,N_8417,N_8591);
nor U9055 (N_9055,N_8620,N_8750);
nor U9056 (N_9056,N_8691,N_8479);
nand U9057 (N_9057,N_8845,N_8987);
and U9058 (N_9058,N_8592,N_8747);
nor U9059 (N_9059,N_8915,N_8473);
xnor U9060 (N_9060,N_8393,N_8476);
and U9061 (N_9061,N_8994,N_8699);
nor U9062 (N_9062,N_8415,N_8300);
or U9063 (N_9063,N_8413,N_8450);
or U9064 (N_9064,N_8497,N_8773);
xnor U9065 (N_9065,N_8283,N_8700);
nand U9066 (N_9066,N_8632,N_8952);
or U9067 (N_9067,N_8869,N_8862);
or U9068 (N_9068,N_8260,N_8984);
xor U9069 (N_9069,N_8914,N_8516);
nor U9070 (N_9070,N_8329,N_8391);
xor U9071 (N_9071,N_8439,N_8968);
nand U9072 (N_9072,N_8452,N_8962);
xnor U9073 (N_9073,N_8590,N_8900);
or U9074 (N_9074,N_8631,N_8438);
nor U9075 (N_9075,N_8511,N_8835);
or U9076 (N_9076,N_8572,N_8879);
xor U9077 (N_9077,N_8359,N_8368);
or U9078 (N_9078,N_8748,N_8780);
xnor U9079 (N_9079,N_8816,N_8802);
nand U9080 (N_9080,N_8890,N_8815);
nand U9081 (N_9081,N_8464,N_8555);
or U9082 (N_9082,N_8716,N_8328);
or U9083 (N_9083,N_8634,N_8732);
and U9084 (N_9084,N_8755,N_8641);
nand U9085 (N_9085,N_8896,N_8635);
or U9086 (N_9086,N_8712,N_8377);
xnor U9087 (N_9087,N_8537,N_8932);
xnor U9088 (N_9088,N_8752,N_8881);
or U9089 (N_9089,N_8650,N_8433);
nor U9090 (N_9090,N_8509,N_8309);
xnor U9091 (N_9091,N_8895,N_8779);
or U9092 (N_9092,N_8355,N_8375);
nor U9093 (N_9093,N_8615,N_8529);
xnor U9094 (N_9094,N_8336,N_8740);
nand U9095 (N_9095,N_8495,N_8749);
and U9096 (N_9096,N_8813,N_8992);
nor U9097 (N_9097,N_8619,N_8348);
and U9098 (N_9098,N_8627,N_8344);
xor U9099 (N_9099,N_8945,N_8959);
or U9100 (N_9100,N_8698,N_8652);
nor U9101 (N_9101,N_8331,N_8535);
xor U9102 (N_9102,N_8954,N_8597);
nor U9103 (N_9103,N_8943,N_8847);
and U9104 (N_9104,N_8621,N_8607);
nor U9105 (N_9105,N_8367,N_8756);
nand U9106 (N_9106,N_8648,N_8918);
nor U9107 (N_9107,N_8825,N_8988);
xor U9108 (N_9108,N_8649,N_8686);
or U9109 (N_9109,N_8289,N_8882);
nor U9110 (N_9110,N_8852,N_8299);
nand U9111 (N_9111,N_8613,N_8787);
and U9112 (N_9112,N_8454,N_8767);
nand U9113 (N_9113,N_8967,N_8425);
nor U9114 (N_9114,N_8817,N_8558);
and U9115 (N_9115,N_8493,N_8724);
xnor U9116 (N_9116,N_8707,N_8982);
nor U9117 (N_9117,N_8272,N_8501);
nand U9118 (N_9118,N_8494,N_8906);
xnor U9119 (N_9119,N_8429,N_8568);
nand U9120 (N_9120,N_8818,N_8547);
and U9121 (N_9121,N_8585,N_8274);
xnor U9122 (N_9122,N_8539,N_8350);
or U9123 (N_9123,N_8941,N_8463);
xnor U9124 (N_9124,N_8769,N_8382);
or U9125 (N_9125,N_8518,N_8322);
xnor U9126 (N_9126,N_8794,N_8804);
and U9127 (N_9127,N_8792,N_8647);
or U9128 (N_9128,N_8745,N_8569);
and U9129 (N_9129,N_8738,N_8286);
or U9130 (N_9130,N_8386,N_8981);
xor U9131 (N_9131,N_8616,N_8296);
and U9132 (N_9132,N_8604,N_8971);
or U9133 (N_9133,N_8910,N_8874);
and U9134 (N_9134,N_8625,N_8305);
or U9135 (N_9135,N_8540,N_8279);
xnor U9136 (N_9136,N_8496,N_8894);
or U9137 (N_9137,N_8435,N_8937);
or U9138 (N_9138,N_8916,N_8673);
or U9139 (N_9139,N_8710,N_8853);
xor U9140 (N_9140,N_8306,N_8901);
or U9141 (N_9141,N_8731,N_8803);
nand U9142 (N_9142,N_8754,N_8432);
xnor U9143 (N_9143,N_8969,N_8360);
nor U9144 (N_9144,N_8601,N_8793);
or U9145 (N_9145,N_8414,N_8566);
nand U9146 (N_9146,N_8837,N_8303);
nand U9147 (N_9147,N_8653,N_8378);
xnor U9148 (N_9148,N_8766,N_8580);
xor U9149 (N_9149,N_8576,N_8323);
nand U9150 (N_9150,N_8687,N_8795);
xnor U9151 (N_9151,N_8584,N_8519);
and U9152 (N_9152,N_8588,N_8885);
or U9153 (N_9153,N_8873,N_8865);
nor U9154 (N_9154,N_8357,N_8284);
nand U9155 (N_9155,N_8776,N_8428);
xor U9156 (N_9156,N_8304,N_8721);
and U9157 (N_9157,N_8701,N_8861);
or U9158 (N_9158,N_8644,N_8266);
nand U9159 (N_9159,N_8596,N_8528);
nand U9160 (N_9160,N_8256,N_8499);
and U9161 (N_9161,N_8696,N_8437);
nand U9162 (N_9162,N_8352,N_8663);
and U9163 (N_9163,N_8904,N_8970);
nor U9164 (N_9164,N_8291,N_8799);
and U9165 (N_9165,N_8638,N_8310);
nand U9166 (N_9166,N_8934,N_8976);
nand U9167 (N_9167,N_8922,N_8361);
xnor U9168 (N_9168,N_8451,N_8395);
nand U9169 (N_9169,N_8645,N_8599);
and U9170 (N_9170,N_8442,N_8251);
xor U9171 (N_9171,N_8267,N_8997);
nor U9172 (N_9172,N_8277,N_8434);
nand U9173 (N_9173,N_8469,N_8844);
nor U9174 (N_9174,N_8843,N_8376);
nand U9175 (N_9175,N_8411,N_8998);
or U9176 (N_9176,N_8418,N_8388);
or U9177 (N_9177,N_8550,N_8783);
xor U9178 (N_9178,N_8408,N_8751);
and U9179 (N_9179,N_8523,N_8928);
or U9180 (N_9180,N_8722,N_8692);
nor U9181 (N_9181,N_8459,N_8927);
nand U9182 (N_9182,N_8911,N_8472);
xnor U9183 (N_9183,N_8764,N_8925);
and U9184 (N_9184,N_8956,N_8757);
and U9185 (N_9185,N_8579,N_8889);
nand U9186 (N_9186,N_8654,N_8931);
or U9187 (N_9187,N_8884,N_8819);
nand U9188 (N_9188,N_8657,N_8586);
nor U9189 (N_9189,N_8353,N_8974);
nor U9190 (N_9190,N_8610,N_8688);
and U9191 (N_9191,N_8705,N_8468);
nand U9192 (N_9192,N_8301,N_8455);
nor U9193 (N_9193,N_8490,N_8401);
or U9194 (N_9194,N_8728,N_8639);
nand U9195 (N_9195,N_8381,N_8878);
nor U9196 (N_9196,N_8784,N_8717);
nor U9197 (N_9197,N_8899,N_8935);
nand U9198 (N_9198,N_8714,N_8951);
nand U9199 (N_9199,N_8946,N_8630);
nor U9200 (N_9200,N_8403,N_8838);
nor U9201 (N_9201,N_8685,N_8668);
and U9202 (N_9202,N_8947,N_8761);
or U9203 (N_9203,N_8695,N_8791);
or U9204 (N_9204,N_8842,N_8978);
or U9205 (N_9205,N_8702,N_8387);
nand U9206 (N_9206,N_8626,N_8789);
nor U9207 (N_9207,N_8905,N_8912);
nor U9208 (N_9208,N_8358,N_8877);
nor U9209 (N_9209,N_8972,N_8595);
xor U9210 (N_9210,N_8849,N_8546);
nor U9211 (N_9211,N_8725,N_8268);
xor U9212 (N_9212,N_8466,N_8252);
and U9213 (N_9213,N_8308,N_8872);
xor U9214 (N_9214,N_8826,N_8933);
and U9215 (N_9215,N_8858,N_8924);
or U9216 (N_9216,N_8913,N_8735);
nand U9217 (N_9217,N_8500,N_8379);
nand U9218 (N_9218,N_8362,N_8907);
or U9219 (N_9219,N_8727,N_8396);
and U9220 (N_9220,N_8957,N_8562);
and U9221 (N_9221,N_8670,N_8759);
or U9222 (N_9222,N_8281,N_8332);
or U9223 (N_9223,N_8392,N_8504);
and U9224 (N_9224,N_8856,N_8561);
xor U9225 (N_9225,N_8614,N_8990);
or U9226 (N_9226,N_8543,N_8581);
nand U9227 (N_9227,N_8807,N_8851);
and U9228 (N_9228,N_8859,N_8522);
and U9229 (N_9229,N_8444,N_8840);
xor U9230 (N_9230,N_8888,N_8427);
nor U9231 (N_9231,N_8545,N_8505);
and U9232 (N_9232,N_8593,N_8423);
xor U9233 (N_9233,N_8734,N_8406);
or U9234 (N_9234,N_8575,N_8542);
and U9235 (N_9235,N_8345,N_8743);
and U9236 (N_9236,N_8541,N_8398);
and U9237 (N_9237,N_8557,N_8640);
nor U9238 (N_9238,N_8973,N_8833);
nor U9239 (N_9239,N_8953,N_8920);
xnor U9240 (N_9240,N_8897,N_8405);
nor U9241 (N_9241,N_8669,N_8312);
nand U9242 (N_9242,N_8339,N_8848);
and U9243 (N_9243,N_8936,N_8474);
xor U9244 (N_9244,N_8975,N_8665);
nor U9245 (N_9245,N_8498,N_8866);
nor U9246 (N_9246,N_8886,N_8351);
and U9247 (N_9247,N_8520,N_8892);
nor U9248 (N_9248,N_8908,N_8354);
or U9249 (N_9249,N_8314,N_8440);
and U9250 (N_9250,N_8506,N_8416);
xnor U9251 (N_9251,N_8919,N_8676);
xor U9252 (N_9252,N_8646,N_8834);
and U9253 (N_9253,N_8589,N_8655);
or U9254 (N_9254,N_8736,N_8797);
nor U9255 (N_9255,N_8262,N_8883);
nand U9256 (N_9256,N_8533,N_8809);
xor U9257 (N_9257,N_8524,N_8921);
xnor U9258 (N_9258,N_8265,N_8292);
or U9259 (N_9259,N_8903,N_8402);
and U9260 (N_9260,N_8857,N_8828);
xor U9261 (N_9261,N_8366,N_8611);
or U9262 (N_9262,N_8502,N_8678);
nor U9263 (N_9263,N_8536,N_8521);
or U9264 (N_9264,N_8333,N_8684);
xor U9265 (N_9265,N_8788,N_8515);
nand U9266 (N_9266,N_8909,N_8704);
or U9267 (N_9267,N_8713,N_8999);
xor U9268 (N_9268,N_8409,N_8563);
and U9269 (N_9269,N_8659,N_8337);
or U9270 (N_9270,N_8552,N_8746);
nor U9271 (N_9271,N_8608,N_8785);
nand U9272 (N_9272,N_8276,N_8940);
xnor U9273 (N_9273,N_8996,N_8683);
nand U9274 (N_9274,N_8349,N_8446);
or U9275 (N_9275,N_8771,N_8460);
or U9276 (N_9276,N_8311,N_8327);
xnor U9277 (N_9277,N_8570,N_8478);
xnor U9278 (N_9278,N_8307,N_8762);
xor U9279 (N_9279,N_8944,N_8715);
and U9280 (N_9280,N_8422,N_8739);
nor U9281 (N_9281,N_8430,N_8275);
nor U9282 (N_9282,N_8841,N_8577);
nand U9283 (N_9283,N_8617,N_8483);
nor U9284 (N_9284,N_8980,N_8263);
nor U9285 (N_9285,N_8565,N_8948);
nand U9286 (N_9286,N_8259,N_8513);
and U9287 (N_9287,N_8812,N_8955);
nor U9288 (N_9288,N_8938,N_8786);
xor U9289 (N_9289,N_8929,N_8324);
nor U9290 (N_9290,N_8829,N_8693);
nor U9291 (N_9291,N_8718,N_8538);
nand U9292 (N_9292,N_8622,N_8775);
xor U9293 (N_9293,N_8346,N_8313);
nor U9294 (N_9294,N_8445,N_8677);
or U9295 (N_9295,N_8991,N_8902);
or U9296 (N_9296,N_8832,N_8605);
or U9297 (N_9297,N_8598,N_8814);
and U9298 (N_9298,N_8318,N_8855);
nor U9299 (N_9299,N_8893,N_8860);
xnor U9300 (N_9300,N_8489,N_8633);
xnor U9301 (N_9301,N_8983,N_8656);
or U9302 (N_9302,N_8282,N_8600);
and U9303 (N_9303,N_8534,N_8508);
or U9304 (N_9304,N_8250,N_8280);
or U9305 (N_9305,N_8369,N_8875);
nor U9306 (N_9306,N_8487,N_8271);
xor U9307 (N_9307,N_8989,N_8612);
xnor U9308 (N_9308,N_8481,N_8790);
xor U9309 (N_9309,N_8461,N_8347);
and U9310 (N_9310,N_8269,N_8682);
and U9311 (N_9311,N_8364,N_8548);
nand U9312 (N_9312,N_8709,N_8449);
or U9313 (N_9313,N_8768,N_8977);
xnor U9314 (N_9314,N_8966,N_8456);
xor U9315 (N_9315,N_8719,N_8573);
xor U9316 (N_9316,N_8443,N_8560);
or U9317 (N_9317,N_8491,N_8993);
nor U9318 (N_9318,N_8930,N_8486);
or U9319 (N_9319,N_8830,N_8338);
xor U9320 (N_9320,N_8574,N_8380);
or U9321 (N_9321,N_8556,N_8839);
and U9322 (N_9322,N_8412,N_8760);
nor U9323 (N_9323,N_8891,N_8703);
or U9324 (N_9324,N_8824,N_8394);
xnor U9325 (N_9325,N_8671,N_8950);
nor U9326 (N_9326,N_8680,N_8330);
xor U9327 (N_9327,N_8742,N_8436);
xnor U9328 (N_9328,N_8868,N_8637);
xor U9329 (N_9329,N_8808,N_8258);
nand U9330 (N_9330,N_8939,N_8629);
xor U9331 (N_9331,N_8798,N_8582);
or U9332 (N_9332,N_8532,N_8876);
nor U9333 (N_9333,N_8926,N_8470);
nor U9334 (N_9334,N_8302,N_8441);
nand U9335 (N_9335,N_8477,N_8694);
nand U9336 (N_9336,N_8317,N_8298);
or U9337 (N_9337,N_8525,N_8503);
nand U9338 (N_9338,N_8471,N_8253);
xor U9339 (N_9339,N_8961,N_8295);
or U9340 (N_9340,N_8325,N_8293);
nor U9341 (N_9341,N_8257,N_8651);
nor U9342 (N_9342,N_8772,N_8365);
or U9343 (N_9343,N_8531,N_8270);
or U9344 (N_9344,N_8898,N_8960);
nand U9345 (N_9345,N_8465,N_8340);
and U9346 (N_9346,N_8553,N_8870);
nand U9347 (N_9347,N_8431,N_8820);
nor U9348 (N_9348,N_8484,N_8782);
nand U9349 (N_9349,N_8697,N_8315);
nand U9350 (N_9350,N_8549,N_8850);
xnor U9351 (N_9351,N_8320,N_8397);
nor U9352 (N_9352,N_8827,N_8512);
nor U9353 (N_9353,N_8801,N_8510);
or U9354 (N_9354,N_8507,N_8711);
xor U9355 (N_9355,N_8863,N_8741);
and U9356 (N_9356,N_8770,N_8390);
or U9357 (N_9357,N_8726,N_8559);
nor U9358 (N_9358,N_8426,N_8544);
and U9359 (N_9359,N_8551,N_8594);
or U9360 (N_9360,N_8297,N_8729);
nor U9361 (N_9361,N_8334,N_8527);
nand U9362 (N_9362,N_8363,N_8419);
xor U9363 (N_9363,N_8744,N_8660);
nor U9364 (N_9364,N_8278,N_8467);
and U9365 (N_9365,N_8462,N_8753);
xnor U9366 (N_9366,N_8400,N_8662);
or U9367 (N_9367,N_8564,N_8796);
nand U9368 (N_9368,N_8758,N_8372);
nand U9369 (N_9369,N_8383,N_8854);
and U9370 (N_9370,N_8805,N_8806);
and U9371 (N_9371,N_8290,N_8404);
and U9372 (N_9372,N_8765,N_8410);
and U9373 (N_9373,N_8294,N_8672);
nor U9374 (N_9374,N_8530,N_8846);
nand U9375 (N_9375,N_8331,N_8819);
or U9376 (N_9376,N_8359,N_8914);
nand U9377 (N_9377,N_8339,N_8937);
and U9378 (N_9378,N_8394,N_8994);
nand U9379 (N_9379,N_8819,N_8715);
nor U9380 (N_9380,N_8284,N_8878);
and U9381 (N_9381,N_8271,N_8441);
nand U9382 (N_9382,N_8949,N_8625);
xor U9383 (N_9383,N_8460,N_8994);
and U9384 (N_9384,N_8858,N_8970);
nand U9385 (N_9385,N_8880,N_8699);
or U9386 (N_9386,N_8502,N_8743);
xnor U9387 (N_9387,N_8744,N_8341);
and U9388 (N_9388,N_8474,N_8562);
xor U9389 (N_9389,N_8556,N_8531);
xor U9390 (N_9390,N_8867,N_8808);
xor U9391 (N_9391,N_8746,N_8668);
xor U9392 (N_9392,N_8458,N_8587);
nor U9393 (N_9393,N_8719,N_8694);
nor U9394 (N_9394,N_8675,N_8400);
or U9395 (N_9395,N_8446,N_8505);
nand U9396 (N_9396,N_8402,N_8748);
nand U9397 (N_9397,N_8894,N_8548);
nand U9398 (N_9398,N_8353,N_8260);
nand U9399 (N_9399,N_8918,N_8773);
or U9400 (N_9400,N_8950,N_8346);
xnor U9401 (N_9401,N_8517,N_8767);
nand U9402 (N_9402,N_8340,N_8265);
nand U9403 (N_9403,N_8512,N_8560);
or U9404 (N_9404,N_8851,N_8419);
and U9405 (N_9405,N_8714,N_8703);
nand U9406 (N_9406,N_8858,N_8927);
and U9407 (N_9407,N_8265,N_8928);
xnor U9408 (N_9408,N_8326,N_8592);
or U9409 (N_9409,N_8902,N_8942);
xor U9410 (N_9410,N_8498,N_8775);
nand U9411 (N_9411,N_8296,N_8636);
xor U9412 (N_9412,N_8467,N_8955);
or U9413 (N_9413,N_8357,N_8470);
xor U9414 (N_9414,N_8731,N_8602);
and U9415 (N_9415,N_8892,N_8646);
or U9416 (N_9416,N_8577,N_8728);
nand U9417 (N_9417,N_8833,N_8277);
nor U9418 (N_9418,N_8816,N_8722);
xor U9419 (N_9419,N_8648,N_8486);
nand U9420 (N_9420,N_8939,N_8612);
nand U9421 (N_9421,N_8704,N_8508);
or U9422 (N_9422,N_8318,N_8704);
nor U9423 (N_9423,N_8666,N_8519);
or U9424 (N_9424,N_8905,N_8623);
xor U9425 (N_9425,N_8624,N_8492);
and U9426 (N_9426,N_8983,N_8903);
and U9427 (N_9427,N_8929,N_8401);
xnor U9428 (N_9428,N_8936,N_8774);
nor U9429 (N_9429,N_8263,N_8404);
and U9430 (N_9430,N_8336,N_8868);
nand U9431 (N_9431,N_8945,N_8254);
nand U9432 (N_9432,N_8481,N_8623);
or U9433 (N_9433,N_8646,N_8307);
nor U9434 (N_9434,N_8908,N_8559);
or U9435 (N_9435,N_8782,N_8561);
and U9436 (N_9436,N_8954,N_8416);
xnor U9437 (N_9437,N_8623,N_8815);
and U9438 (N_9438,N_8255,N_8699);
xnor U9439 (N_9439,N_8810,N_8467);
and U9440 (N_9440,N_8753,N_8780);
and U9441 (N_9441,N_8908,N_8636);
or U9442 (N_9442,N_8824,N_8377);
nor U9443 (N_9443,N_8537,N_8370);
nand U9444 (N_9444,N_8684,N_8699);
xnor U9445 (N_9445,N_8838,N_8673);
or U9446 (N_9446,N_8254,N_8347);
or U9447 (N_9447,N_8941,N_8878);
and U9448 (N_9448,N_8803,N_8383);
or U9449 (N_9449,N_8436,N_8892);
nor U9450 (N_9450,N_8469,N_8446);
and U9451 (N_9451,N_8557,N_8495);
and U9452 (N_9452,N_8955,N_8790);
nand U9453 (N_9453,N_8645,N_8662);
xor U9454 (N_9454,N_8968,N_8411);
nor U9455 (N_9455,N_8694,N_8738);
xnor U9456 (N_9456,N_8890,N_8673);
nand U9457 (N_9457,N_8275,N_8754);
and U9458 (N_9458,N_8859,N_8265);
nand U9459 (N_9459,N_8636,N_8971);
or U9460 (N_9460,N_8694,N_8637);
or U9461 (N_9461,N_8931,N_8804);
or U9462 (N_9462,N_8649,N_8703);
xnor U9463 (N_9463,N_8667,N_8743);
and U9464 (N_9464,N_8644,N_8546);
or U9465 (N_9465,N_8610,N_8805);
nor U9466 (N_9466,N_8795,N_8779);
xnor U9467 (N_9467,N_8637,N_8884);
or U9468 (N_9468,N_8305,N_8397);
nor U9469 (N_9469,N_8931,N_8664);
nand U9470 (N_9470,N_8520,N_8746);
and U9471 (N_9471,N_8267,N_8583);
nor U9472 (N_9472,N_8758,N_8315);
and U9473 (N_9473,N_8935,N_8295);
nand U9474 (N_9474,N_8437,N_8994);
or U9475 (N_9475,N_8613,N_8505);
nand U9476 (N_9476,N_8543,N_8754);
or U9477 (N_9477,N_8511,N_8715);
or U9478 (N_9478,N_8678,N_8879);
nand U9479 (N_9479,N_8309,N_8907);
and U9480 (N_9480,N_8702,N_8720);
xor U9481 (N_9481,N_8575,N_8639);
and U9482 (N_9482,N_8836,N_8501);
nor U9483 (N_9483,N_8534,N_8309);
or U9484 (N_9484,N_8474,N_8880);
or U9485 (N_9485,N_8426,N_8954);
xnor U9486 (N_9486,N_8882,N_8893);
nor U9487 (N_9487,N_8674,N_8262);
or U9488 (N_9488,N_8307,N_8690);
and U9489 (N_9489,N_8927,N_8437);
and U9490 (N_9490,N_8343,N_8880);
xnor U9491 (N_9491,N_8819,N_8525);
nor U9492 (N_9492,N_8533,N_8650);
and U9493 (N_9493,N_8270,N_8503);
nor U9494 (N_9494,N_8706,N_8777);
nor U9495 (N_9495,N_8619,N_8391);
nor U9496 (N_9496,N_8657,N_8572);
and U9497 (N_9497,N_8959,N_8976);
xor U9498 (N_9498,N_8931,N_8625);
xnor U9499 (N_9499,N_8435,N_8520);
and U9500 (N_9500,N_8577,N_8330);
and U9501 (N_9501,N_8814,N_8643);
nor U9502 (N_9502,N_8497,N_8424);
nor U9503 (N_9503,N_8658,N_8861);
or U9504 (N_9504,N_8983,N_8540);
and U9505 (N_9505,N_8814,N_8667);
nand U9506 (N_9506,N_8649,N_8549);
nor U9507 (N_9507,N_8904,N_8456);
and U9508 (N_9508,N_8880,N_8607);
or U9509 (N_9509,N_8875,N_8427);
nand U9510 (N_9510,N_8410,N_8817);
or U9511 (N_9511,N_8793,N_8358);
or U9512 (N_9512,N_8624,N_8606);
nand U9513 (N_9513,N_8534,N_8431);
and U9514 (N_9514,N_8489,N_8791);
nand U9515 (N_9515,N_8435,N_8270);
and U9516 (N_9516,N_8659,N_8778);
and U9517 (N_9517,N_8432,N_8252);
xor U9518 (N_9518,N_8742,N_8938);
xor U9519 (N_9519,N_8988,N_8625);
nor U9520 (N_9520,N_8782,N_8667);
nand U9521 (N_9521,N_8573,N_8494);
nor U9522 (N_9522,N_8929,N_8630);
or U9523 (N_9523,N_8973,N_8907);
xnor U9524 (N_9524,N_8683,N_8778);
or U9525 (N_9525,N_8255,N_8780);
and U9526 (N_9526,N_8598,N_8439);
or U9527 (N_9527,N_8919,N_8566);
xnor U9528 (N_9528,N_8870,N_8475);
or U9529 (N_9529,N_8836,N_8913);
xnor U9530 (N_9530,N_8858,N_8304);
and U9531 (N_9531,N_8977,N_8422);
or U9532 (N_9532,N_8650,N_8838);
xor U9533 (N_9533,N_8658,N_8999);
nor U9534 (N_9534,N_8705,N_8959);
xnor U9535 (N_9535,N_8331,N_8923);
and U9536 (N_9536,N_8794,N_8608);
or U9537 (N_9537,N_8895,N_8324);
xnor U9538 (N_9538,N_8915,N_8446);
nor U9539 (N_9539,N_8767,N_8482);
and U9540 (N_9540,N_8363,N_8304);
and U9541 (N_9541,N_8332,N_8344);
or U9542 (N_9542,N_8835,N_8794);
nor U9543 (N_9543,N_8607,N_8955);
and U9544 (N_9544,N_8884,N_8394);
and U9545 (N_9545,N_8735,N_8359);
or U9546 (N_9546,N_8313,N_8571);
nand U9547 (N_9547,N_8783,N_8310);
xnor U9548 (N_9548,N_8793,N_8597);
nor U9549 (N_9549,N_8835,N_8690);
and U9550 (N_9550,N_8397,N_8922);
xnor U9551 (N_9551,N_8609,N_8439);
nand U9552 (N_9552,N_8381,N_8670);
nor U9553 (N_9553,N_8829,N_8530);
xor U9554 (N_9554,N_8543,N_8515);
nand U9555 (N_9555,N_8894,N_8561);
nor U9556 (N_9556,N_8702,N_8799);
or U9557 (N_9557,N_8303,N_8305);
or U9558 (N_9558,N_8814,N_8940);
and U9559 (N_9559,N_8898,N_8400);
and U9560 (N_9560,N_8602,N_8622);
and U9561 (N_9561,N_8542,N_8460);
xnor U9562 (N_9562,N_8753,N_8338);
nor U9563 (N_9563,N_8808,N_8614);
nor U9564 (N_9564,N_8538,N_8253);
and U9565 (N_9565,N_8780,N_8974);
nand U9566 (N_9566,N_8769,N_8802);
nand U9567 (N_9567,N_8275,N_8801);
nand U9568 (N_9568,N_8894,N_8307);
xnor U9569 (N_9569,N_8322,N_8462);
and U9570 (N_9570,N_8553,N_8960);
or U9571 (N_9571,N_8934,N_8529);
and U9572 (N_9572,N_8646,N_8886);
xnor U9573 (N_9573,N_8605,N_8850);
xnor U9574 (N_9574,N_8609,N_8331);
nand U9575 (N_9575,N_8768,N_8566);
or U9576 (N_9576,N_8524,N_8804);
or U9577 (N_9577,N_8657,N_8882);
and U9578 (N_9578,N_8762,N_8637);
or U9579 (N_9579,N_8972,N_8355);
xnor U9580 (N_9580,N_8837,N_8297);
and U9581 (N_9581,N_8407,N_8441);
or U9582 (N_9582,N_8343,N_8840);
nor U9583 (N_9583,N_8414,N_8945);
nand U9584 (N_9584,N_8718,N_8896);
or U9585 (N_9585,N_8866,N_8772);
and U9586 (N_9586,N_8671,N_8778);
nor U9587 (N_9587,N_8930,N_8942);
and U9588 (N_9588,N_8658,N_8595);
nor U9589 (N_9589,N_8657,N_8315);
xnor U9590 (N_9590,N_8455,N_8505);
or U9591 (N_9591,N_8948,N_8820);
nand U9592 (N_9592,N_8577,N_8252);
xnor U9593 (N_9593,N_8398,N_8603);
and U9594 (N_9594,N_8506,N_8454);
and U9595 (N_9595,N_8962,N_8269);
nand U9596 (N_9596,N_8398,N_8409);
or U9597 (N_9597,N_8732,N_8622);
nand U9598 (N_9598,N_8933,N_8503);
or U9599 (N_9599,N_8636,N_8255);
xor U9600 (N_9600,N_8678,N_8655);
nand U9601 (N_9601,N_8280,N_8838);
nor U9602 (N_9602,N_8253,N_8616);
xor U9603 (N_9603,N_8756,N_8261);
xnor U9604 (N_9604,N_8596,N_8864);
or U9605 (N_9605,N_8534,N_8852);
nand U9606 (N_9606,N_8383,N_8786);
or U9607 (N_9607,N_8955,N_8769);
nor U9608 (N_9608,N_8309,N_8867);
xor U9609 (N_9609,N_8389,N_8805);
xnor U9610 (N_9610,N_8983,N_8478);
and U9611 (N_9611,N_8299,N_8495);
nand U9612 (N_9612,N_8613,N_8826);
nand U9613 (N_9613,N_8961,N_8877);
xor U9614 (N_9614,N_8773,N_8513);
or U9615 (N_9615,N_8586,N_8452);
and U9616 (N_9616,N_8271,N_8394);
or U9617 (N_9617,N_8359,N_8774);
nand U9618 (N_9618,N_8783,N_8980);
nand U9619 (N_9619,N_8777,N_8612);
nand U9620 (N_9620,N_8760,N_8391);
nor U9621 (N_9621,N_8980,N_8890);
nand U9622 (N_9622,N_8861,N_8525);
nor U9623 (N_9623,N_8297,N_8597);
xor U9624 (N_9624,N_8767,N_8732);
nand U9625 (N_9625,N_8496,N_8480);
and U9626 (N_9626,N_8373,N_8432);
nor U9627 (N_9627,N_8726,N_8374);
or U9628 (N_9628,N_8420,N_8273);
nand U9629 (N_9629,N_8748,N_8323);
nor U9630 (N_9630,N_8375,N_8551);
nor U9631 (N_9631,N_8644,N_8570);
nor U9632 (N_9632,N_8753,N_8729);
nor U9633 (N_9633,N_8585,N_8665);
or U9634 (N_9634,N_8522,N_8929);
xor U9635 (N_9635,N_8918,N_8416);
nand U9636 (N_9636,N_8428,N_8946);
xor U9637 (N_9637,N_8261,N_8831);
nand U9638 (N_9638,N_8870,N_8380);
xnor U9639 (N_9639,N_8427,N_8292);
nor U9640 (N_9640,N_8543,N_8345);
nand U9641 (N_9641,N_8814,N_8697);
nor U9642 (N_9642,N_8395,N_8716);
or U9643 (N_9643,N_8397,N_8418);
or U9644 (N_9644,N_8275,N_8391);
nand U9645 (N_9645,N_8626,N_8741);
xor U9646 (N_9646,N_8686,N_8653);
nor U9647 (N_9647,N_8812,N_8277);
nand U9648 (N_9648,N_8597,N_8266);
and U9649 (N_9649,N_8425,N_8664);
xnor U9650 (N_9650,N_8297,N_8831);
or U9651 (N_9651,N_8376,N_8676);
nor U9652 (N_9652,N_8907,N_8531);
or U9653 (N_9653,N_8965,N_8358);
or U9654 (N_9654,N_8791,N_8938);
or U9655 (N_9655,N_8927,N_8844);
nand U9656 (N_9656,N_8569,N_8331);
nand U9657 (N_9657,N_8463,N_8527);
nor U9658 (N_9658,N_8600,N_8419);
nand U9659 (N_9659,N_8345,N_8828);
or U9660 (N_9660,N_8955,N_8616);
nand U9661 (N_9661,N_8980,N_8914);
nor U9662 (N_9662,N_8819,N_8550);
and U9663 (N_9663,N_8823,N_8367);
nor U9664 (N_9664,N_8625,N_8344);
nand U9665 (N_9665,N_8496,N_8716);
and U9666 (N_9666,N_8701,N_8726);
xor U9667 (N_9667,N_8256,N_8699);
or U9668 (N_9668,N_8758,N_8621);
nor U9669 (N_9669,N_8862,N_8628);
or U9670 (N_9670,N_8357,N_8933);
or U9671 (N_9671,N_8468,N_8767);
or U9672 (N_9672,N_8868,N_8325);
nor U9673 (N_9673,N_8353,N_8429);
nor U9674 (N_9674,N_8657,N_8435);
nand U9675 (N_9675,N_8396,N_8254);
xnor U9676 (N_9676,N_8894,N_8848);
xnor U9677 (N_9677,N_8858,N_8632);
and U9678 (N_9678,N_8619,N_8729);
xor U9679 (N_9679,N_8655,N_8539);
nand U9680 (N_9680,N_8523,N_8746);
or U9681 (N_9681,N_8272,N_8948);
xnor U9682 (N_9682,N_8542,N_8591);
xor U9683 (N_9683,N_8538,N_8515);
nor U9684 (N_9684,N_8701,N_8582);
nor U9685 (N_9685,N_8884,N_8670);
xnor U9686 (N_9686,N_8788,N_8797);
or U9687 (N_9687,N_8455,N_8478);
xnor U9688 (N_9688,N_8355,N_8404);
nor U9689 (N_9689,N_8808,N_8887);
nand U9690 (N_9690,N_8766,N_8344);
nand U9691 (N_9691,N_8897,N_8578);
nor U9692 (N_9692,N_8499,N_8910);
nand U9693 (N_9693,N_8420,N_8325);
and U9694 (N_9694,N_8623,N_8320);
nor U9695 (N_9695,N_8644,N_8977);
nor U9696 (N_9696,N_8533,N_8454);
and U9697 (N_9697,N_8319,N_8701);
or U9698 (N_9698,N_8589,N_8958);
nor U9699 (N_9699,N_8868,N_8369);
or U9700 (N_9700,N_8977,N_8703);
nand U9701 (N_9701,N_8452,N_8679);
nand U9702 (N_9702,N_8399,N_8280);
nor U9703 (N_9703,N_8803,N_8807);
and U9704 (N_9704,N_8508,N_8266);
or U9705 (N_9705,N_8957,N_8297);
nand U9706 (N_9706,N_8866,N_8421);
or U9707 (N_9707,N_8780,N_8655);
and U9708 (N_9708,N_8547,N_8957);
or U9709 (N_9709,N_8915,N_8549);
nor U9710 (N_9710,N_8885,N_8810);
xnor U9711 (N_9711,N_8929,N_8260);
and U9712 (N_9712,N_8619,N_8364);
or U9713 (N_9713,N_8413,N_8310);
xnor U9714 (N_9714,N_8543,N_8266);
and U9715 (N_9715,N_8527,N_8985);
nor U9716 (N_9716,N_8418,N_8386);
nor U9717 (N_9717,N_8559,N_8956);
xor U9718 (N_9718,N_8408,N_8904);
nor U9719 (N_9719,N_8973,N_8629);
nor U9720 (N_9720,N_8683,N_8845);
or U9721 (N_9721,N_8598,N_8595);
or U9722 (N_9722,N_8263,N_8951);
and U9723 (N_9723,N_8764,N_8554);
xnor U9724 (N_9724,N_8984,N_8472);
and U9725 (N_9725,N_8493,N_8400);
or U9726 (N_9726,N_8740,N_8646);
or U9727 (N_9727,N_8558,N_8565);
xor U9728 (N_9728,N_8969,N_8977);
and U9729 (N_9729,N_8529,N_8377);
nand U9730 (N_9730,N_8600,N_8958);
xnor U9731 (N_9731,N_8970,N_8305);
nor U9732 (N_9732,N_8846,N_8368);
xnor U9733 (N_9733,N_8896,N_8429);
nand U9734 (N_9734,N_8771,N_8515);
or U9735 (N_9735,N_8934,N_8726);
nand U9736 (N_9736,N_8413,N_8369);
nor U9737 (N_9737,N_8904,N_8958);
nor U9738 (N_9738,N_8339,N_8985);
nor U9739 (N_9739,N_8499,N_8450);
nor U9740 (N_9740,N_8675,N_8579);
and U9741 (N_9741,N_8423,N_8287);
xnor U9742 (N_9742,N_8493,N_8634);
xor U9743 (N_9743,N_8471,N_8665);
and U9744 (N_9744,N_8638,N_8974);
nand U9745 (N_9745,N_8394,N_8784);
nand U9746 (N_9746,N_8776,N_8835);
and U9747 (N_9747,N_8743,N_8257);
nand U9748 (N_9748,N_8659,N_8417);
xnor U9749 (N_9749,N_8969,N_8964);
nor U9750 (N_9750,N_9443,N_9113);
or U9751 (N_9751,N_9404,N_9579);
or U9752 (N_9752,N_9039,N_9091);
xnor U9753 (N_9753,N_9024,N_9205);
xnor U9754 (N_9754,N_9350,N_9636);
xnor U9755 (N_9755,N_9660,N_9374);
and U9756 (N_9756,N_9232,N_9026);
nor U9757 (N_9757,N_9449,N_9191);
and U9758 (N_9758,N_9440,N_9391);
nand U9759 (N_9759,N_9461,N_9160);
nand U9760 (N_9760,N_9613,N_9500);
or U9761 (N_9761,N_9220,N_9177);
nor U9762 (N_9762,N_9437,N_9467);
nand U9763 (N_9763,N_9485,N_9609);
and U9764 (N_9764,N_9451,N_9158);
nor U9765 (N_9765,N_9325,N_9653);
xnor U9766 (N_9766,N_9625,N_9320);
and U9767 (N_9767,N_9617,N_9706);
nand U9768 (N_9768,N_9596,N_9241);
and U9769 (N_9769,N_9140,N_9086);
or U9770 (N_9770,N_9657,N_9360);
or U9771 (N_9771,N_9628,N_9203);
or U9772 (N_9772,N_9742,N_9152);
nor U9773 (N_9773,N_9080,N_9056);
or U9774 (N_9774,N_9299,N_9604);
nor U9775 (N_9775,N_9690,N_9547);
nand U9776 (N_9776,N_9606,N_9621);
nor U9777 (N_9777,N_9726,N_9081);
nand U9778 (N_9778,N_9531,N_9398);
nor U9779 (N_9779,N_9484,N_9292);
xnor U9780 (N_9780,N_9174,N_9560);
xnor U9781 (N_9781,N_9571,N_9051);
nor U9782 (N_9782,N_9243,N_9058);
or U9783 (N_9783,N_9352,N_9746);
xor U9784 (N_9784,N_9736,N_9458);
nand U9785 (N_9785,N_9704,N_9632);
and U9786 (N_9786,N_9186,N_9365);
xor U9787 (N_9787,N_9240,N_9445);
or U9788 (N_9788,N_9748,N_9734);
and U9789 (N_9789,N_9427,N_9337);
xor U9790 (N_9790,N_9209,N_9361);
or U9791 (N_9791,N_9169,N_9137);
nor U9792 (N_9792,N_9366,N_9647);
nand U9793 (N_9793,N_9099,N_9181);
and U9794 (N_9794,N_9085,N_9249);
and U9795 (N_9795,N_9151,N_9370);
and U9796 (N_9796,N_9127,N_9201);
nand U9797 (N_9797,N_9543,N_9228);
nor U9798 (N_9798,N_9421,N_9576);
nand U9799 (N_9799,N_9568,N_9067);
xor U9800 (N_9800,N_9331,N_9263);
nor U9801 (N_9801,N_9645,N_9117);
nor U9802 (N_9802,N_9256,N_9721);
and U9803 (N_9803,N_9394,N_9426);
and U9804 (N_9804,N_9522,N_9048);
and U9805 (N_9805,N_9372,N_9095);
nand U9806 (N_9806,N_9573,N_9066);
xor U9807 (N_9807,N_9434,N_9304);
or U9808 (N_9808,N_9592,N_9640);
or U9809 (N_9809,N_9428,N_9005);
and U9810 (N_9810,N_9214,N_9495);
xnor U9811 (N_9811,N_9261,N_9655);
nor U9812 (N_9812,N_9709,N_9245);
nand U9813 (N_9813,N_9298,N_9504);
nand U9814 (N_9814,N_9712,N_9676);
nand U9815 (N_9815,N_9662,N_9567);
nor U9816 (N_9816,N_9217,N_9057);
xor U9817 (N_9817,N_9650,N_9247);
or U9818 (N_9818,N_9441,N_9699);
nor U9819 (N_9819,N_9462,N_9120);
nor U9820 (N_9820,N_9025,N_9079);
xor U9821 (N_9821,N_9255,N_9028);
or U9822 (N_9822,N_9224,N_9674);
or U9823 (N_9823,N_9179,N_9727);
and U9824 (N_9824,N_9288,N_9377);
nand U9825 (N_9825,N_9725,N_9110);
xor U9826 (N_9826,N_9431,N_9368);
nand U9827 (N_9827,N_9083,N_9555);
nand U9828 (N_9828,N_9023,N_9591);
and U9829 (N_9829,N_9528,N_9313);
nand U9830 (N_9830,N_9615,N_9733);
and U9831 (N_9831,N_9605,N_9334);
nor U9832 (N_9832,N_9344,N_9001);
or U9833 (N_9833,N_9561,N_9306);
or U9834 (N_9834,N_9143,N_9332);
nand U9835 (N_9835,N_9737,N_9371);
and U9836 (N_9836,N_9652,N_9603);
or U9837 (N_9837,N_9116,N_9622);
xnor U9838 (N_9838,N_9097,N_9167);
nand U9839 (N_9839,N_9040,N_9716);
nand U9840 (N_9840,N_9314,N_9134);
nand U9841 (N_9841,N_9094,N_9506);
xnor U9842 (N_9842,N_9390,N_9651);
xor U9843 (N_9843,N_9045,N_9038);
and U9844 (N_9844,N_9469,N_9385);
nor U9845 (N_9845,N_9614,N_9211);
or U9846 (N_9846,N_9319,N_9121);
or U9847 (N_9847,N_9675,N_9397);
or U9848 (N_9848,N_9358,N_9542);
and U9849 (N_9849,N_9303,N_9698);
xnor U9850 (N_9850,N_9607,N_9087);
xnor U9851 (N_9851,N_9705,N_9339);
or U9852 (N_9852,N_9092,N_9406);
or U9853 (N_9853,N_9523,N_9073);
nand U9854 (N_9854,N_9638,N_9035);
nand U9855 (N_9855,N_9043,N_9700);
nor U9856 (N_9856,N_9257,N_9291);
nor U9857 (N_9857,N_9537,N_9046);
or U9858 (N_9858,N_9264,N_9223);
xor U9859 (N_9859,N_9269,N_9102);
or U9860 (N_9860,N_9150,N_9659);
xnor U9861 (N_9861,N_9107,N_9405);
nand U9862 (N_9862,N_9012,N_9435);
or U9863 (N_9863,N_9007,N_9723);
or U9864 (N_9864,N_9146,N_9741);
or U9865 (N_9865,N_9180,N_9093);
or U9866 (N_9866,N_9558,N_9408);
and U9867 (N_9867,N_9172,N_9731);
nand U9868 (N_9868,N_9600,N_9738);
or U9869 (N_9869,N_9595,N_9271);
or U9870 (N_9870,N_9032,N_9559);
nor U9871 (N_9871,N_9052,N_9598);
or U9872 (N_9872,N_9400,N_9494);
nand U9873 (N_9873,N_9399,N_9572);
nand U9874 (N_9874,N_9487,N_9208);
and U9875 (N_9875,N_9016,N_9381);
and U9876 (N_9876,N_9379,N_9532);
xnor U9877 (N_9877,N_9307,N_9565);
and U9878 (N_9878,N_9135,N_9509);
nand U9879 (N_9879,N_9070,N_9029);
and U9880 (N_9880,N_9378,N_9017);
and U9881 (N_9881,N_9316,N_9281);
nor U9882 (N_9882,N_9597,N_9284);
or U9883 (N_9883,N_9432,N_9589);
and U9884 (N_9884,N_9218,N_9602);
nand U9885 (N_9885,N_9688,N_9646);
or U9886 (N_9886,N_9342,N_9041);
nor U9887 (N_9887,N_9252,N_9594);
nand U9888 (N_9888,N_9586,N_9010);
nand U9889 (N_9889,N_9015,N_9225);
nor U9890 (N_9890,N_9195,N_9265);
and U9891 (N_9891,N_9612,N_9219);
or U9892 (N_9892,N_9315,N_9515);
or U9893 (N_9893,N_9136,N_9680);
or U9894 (N_9894,N_9090,N_9514);
nand U9895 (N_9895,N_9422,N_9419);
nand U9896 (N_9896,N_9412,N_9566);
or U9897 (N_9897,N_9672,N_9683);
or U9898 (N_9898,N_9367,N_9351);
and U9899 (N_9899,N_9335,N_9343);
nor U9900 (N_9900,N_9720,N_9533);
nor U9901 (N_9901,N_9132,N_9004);
nand U9902 (N_9902,N_9037,N_9403);
xnor U9903 (N_9903,N_9587,N_9444);
nor U9904 (N_9904,N_9165,N_9295);
or U9905 (N_9905,N_9154,N_9643);
nand U9906 (N_9906,N_9623,N_9144);
and U9907 (N_9907,N_9138,N_9356);
xnor U9908 (N_9908,N_9329,N_9153);
nand U9909 (N_9909,N_9654,N_9049);
or U9910 (N_9910,N_9664,N_9145);
nor U9911 (N_9911,N_9318,N_9616);
and U9912 (N_9912,N_9354,N_9003);
and U9913 (N_9913,N_9078,N_9108);
nor U9914 (N_9914,N_9216,N_9388);
nor U9915 (N_9915,N_9562,N_9701);
nand U9916 (N_9916,N_9627,N_9266);
nand U9917 (N_9917,N_9418,N_9278);
nor U9918 (N_9918,N_9340,N_9502);
nand U9919 (N_9919,N_9668,N_9710);
nor U9920 (N_9920,N_9302,N_9658);
nor U9921 (N_9921,N_9364,N_9194);
xnor U9922 (N_9922,N_9280,N_9456);
or U9923 (N_9923,N_9473,N_9410);
xnor U9924 (N_9924,N_9088,N_9417);
nor U9925 (N_9925,N_9231,N_9715);
or U9926 (N_9926,N_9103,N_9393);
nand U9927 (N_9927,N_9549,N_9663);
or U9928 (N_9928,N_9062,N_9253);
or U9929 (N_9929,N_9407,N_9348);
or U9930 (N_9930,N_9133,N_9239);
nand U9931 (N_9931,N_9525,N_9577);
nor U9932 (N_9932,N_9115,N_9055);
nand U9933 (N_9933,N_9050,N_9420);
nor U9934 (N_9934,N_9489,N_9262);
nand U9935 (N_9935,N_9250,N_9375);
nand U9936 (N_9936,N_9460,N_9126);
nor U9937 (N_9937,N_9268,N_9207);
or U9938 (N_9938,N_9749,N_9230);
nor U9939 (N_9939,N_9027,N_9020);
and U9940 (N_9940,N_9213,N_9511);
or U9941 (N_9941,N_9745,N_9521);
nor U9942 (N_9942,N_9516,N_9499);
nand U9943 (N_9943,N_9369,N_9535);
nand U9944 (N_9944,N_9197,N_9722);
or U9945 (N_9945,N_9130,N_9582);
and U9946 (N_9946,N_9159,N_9061);
xnor U9947 (N_9947,N_9128,N_9357);
or U9948 (N_9948,N_9242,N_9382);
nand U9949 (N_9949,N_9297,N_9717);
xor U9950 (N_9950,N_9168,N_9554);
xor U9951 (N_9951,N_9327,N_9148);
nand U9952 (N_9952,N_9294,N_9301);
or U9953 (N_9953,N_9321,N_9633);
nor U9954 (N_9954,N_9311,N_9074);
or U9955 (N_9955,N_9258,N_9510);
or U9956 (N_9956,N_9744,N_9411);
nand U9957 (N_9957,N_9682,N_9149);
nor U9958 (N_9958,N_9210,N_9383);
nand U9959 (N_9959,N_9323,N_9122);
and U9960 (N_9960,N_9142,N_9707);
nor U9961 (N_9961,N_9063,N_9059);
and U9962 (N_9962,N_9060,N_9539);
xor U9963 (N_9963,N_9100,N_9109);
or U9964 (N_9964,N_9730,N_9466);
or U9965 (N_9965,N_9488,N_9464);
xnor U9966 (N_9966,N_9260,N_9279);
nand U9967 (N_9967,N_9237,N_9147);
xor U9968 (N_9968,N_9416,N_9082);
or U9969 (N_9969,N_9503,N_9601);
and U9970 (N_9970,N_9719,N_9157);
and U9971 (N_9971,N_9548,N_9305);
nand U9972 (N_9972,N_9696,N_9436);
xor U9973 (N_9973,N_9386,N_9006);
xnor U9974 (N_9974,N_9124,N_9076);
xnor U9975 (N_9975,N_9557,N_9362);
and U9976 (N_9976,N_9282,N_9442);
nor U9977 (N_9977,N_9123,N_9013);
and U9978 (N_9978,N_9501,N_9170);
xor U9979 (N_9979,N_9118,N_9474);
xor U9980 (N_9980,N_9202,N_9183);
nand U9981 (N_9981,N_9105,N_9517);
nor U9982 (N_9982,N_9353,N_9112);
or U9983 (N_9983,N_9275,N_9141);
and U9984 (N_9984,N_9527,N_9328);
and U9985 (N_9985,N_9359,N_9190);
or U9986 (N_9986,N_9656,N_9193);
nor U9987 (N_9987,N_9739,N_9452);
nor U9988 (N_9988,N_9396,N_9491);
or U9989 (N_9989,N_9574,N_9681);
or U9990 (N_9990,N_9175,N_9639);
xor U9991 (N_9991,N_9333,N_9611);
nor U9992 (N_9992,N_9714,N_9564);
nand U9993 (N_9993,N_9187,N_9376);
nor U9994 (N_9994,N_9430,N_9014);
and U9995 (N_9995,N_9054,N_9077);
nand U9996 (N_9996,N_9414,N_9324);
xor U9997 (N_9997,N_9585,N_9139);
or U9998 (N_9998,N_9283,N_9310);
nor U9999 (N_9999,N_9641,N_9273);
and U10000 (N_10000,N_9665,N_9238);
or U10001 (N_10001,N_9630,N_9518);
and U10002 (N_10002,N_9200,N_9008);
and U10003 (N_10003,N_9155,N_9125);
nand U10004 (N_10004,N_9526,N_9096);
nand U10005 (N_10005,N_9317,N_9673);
or U10006 (N_10006,N_9387,N_9729);
xnor U10007 (N_10007,N_9496,N_9098);
nor U10008 (N_10008,N_9735,N_9724);
or U10009 (N_10009,N_9718,N_9234);
nand U10010 (N_10010,N_9669,N_9661);
nand U10011 (N_10011,N_9300,N_9446);
and U10012 (N_10012,N_9610,N_9479);
nand U10013 (N_10013,N_9053,N_9164);
xnor U10014 (N_10014,N_9289,N_9563);
or U10015 (N_10015,N_9246,N_9634);
or U10016 (N_10016,N_9072,N_9593);
and U10017 (N_10017,N_9251,N_9553);
nor U10018 (N_10018,N_9689,N_9580);
xor U10019 (N_10019,N_9171,N_9695);
nor U10020 (N_10020,N_9678,N_9002);
xor U10021 (N_10021,N_9471,N_9244);
nand U10022 (N_10022,N_9740,N_9472);
and U10023 (N_10023,N_9021,N_9270);
xor U10024 (N_10024,N_9009,N_9747);
nor U10025 (N_10025,N_9578,N_9743);
nor U10026 (N_10026,N_9429,N_9693);
nand U10027 (N_10027,N_9454,N_9104);
and U10028 (N_10028,N_9463,N_9274);
nor U10029 (N_10029,N_9166,N_9538);
and U10030 (N_10030,N_9345,N_9308);
xor U10031 (N_10031,N_9570,N_9185);
nand U10032 (N_10032,N_9536,N_9413);
nor U10033 (N_10033,N_9433,N_9544);
or U10034 (N_10034,N_9624,N_9581);
nand U10035 (N_10035,N_9644,N_9034);
nand U10036 (N_10036,N_9330,N_9176);
or U10037 (N_10037,N_9694,N_9030);
or U10038 (N_10038,N_9031,N_9022);
nor U10039 (N_10039,N_9529,N_9524);
nor U10040 (N_10040,N_9507,N_9424);
or U10041 (N_10041,N_9163,N_9033);
xor U10042 (N_10042,N_9119,N_9178);
nor U10043 (N_10043,N_9401,N_9346);
xor U10044 (N_10044,N_9227,N_9161);
xnor U10045 (N_10045,N_9703,N_9044);
xnor U10046 (N_10046,N_9711,N_9728);
and U10047 (N_10047,N_9089,N_9687);
nand U10048 (N_10048,N_9649,N_9392);
xnor U10049 (N_10049,N_9459,N_9453);
and U10050 (N_10050,N_9497,N_9546);
and U10051 (N_10051,N_9423,N_9530);
nand U10052 (N_10052,N_9259,N_9212);
nor U10053 (N_10053,N_9642,N_9620);
and U10054 (N_10054,N_9309,N_9018);
or U10055 (N_10055,N_9409,N_9475);
nor U10056 (N_10056,N_9296,N_9691);
nor U10057 (N_10057,N_9285,N_9222);
nor U10058 (N_10058,N_9713,N_9492);
or U10059 (N_10059,N_9671,N_9189);
nor U10060 (N_10060,N_9267,N_9069);
and U10061 (N_10061,N_9215,N_9584);
nand U10062 (N_10062,N_9448,N_9326);
nand U10063 (N_10063,N_9519,N_9470);
nor U10064 (N_10064,N_9481,N_9498);
and U10065 (N_10065,N_9708,N_9619);
nand U10066 (N_10066,N_9106,N_9512);
nor U10067 (N_10067,N_9483,N_9355);
and U10068 (N_10068,N_9490,N_9482);
and U10069 (N_10069,N_9480,N_9588);
nand U10070 (N_10070,N_9084,N_9156);
and U10071 (N_10071,N_9286,N_9465);
xnor U10072 (N_10072,N_9235,N_9590);
nand U10073 (N_10073,N_9666,N_9686);
xnor U10074 (N_10074,N_9162,N_9635);
or U10075 (N_10075,N_9114,N_9047);
and U10076 (N_10076,N_9534,N_9198);
or U10077 (N_10077,N_9363,N_9425);
or U10078 (N_10078,N_9384,N_9184);
nand U10079 (N_10079,N_9520,N_9447);
nand U10080 (N_10080,N_9293,N_9347);
xnor U10081 (N_10081,N_9287,N_9248);
and U10082 (N_10082,N_9322,N_9575);
or U10083 (N_10083,N_9349,N_9000);
or U10084 (N_10084,N_9276,N_9075);
nor U10085 (N_10085,N_9233,N_9599);
or U10086 (N_10086,N_9648,N_9196);
nor U10087 (N_10087,N_9468,N_9667);
or U10088 (N_10088,N_9131,N_9476);
xor U10089 (N_10089,N_9637,N_9583);
xor U10090 (N_10090,N_9272,N_9290);
xor U10091 (N_10091,N_9556,N_9692);
xor U10092 (N_10092,N_9373,N_9685);
nor U10093 (N_10093,N_9226,N_9415);
or U10094 (N_10094,N_9455,N_9629);
and U10095 (N_10095,N_9540,N_9129);
and U10096 (N_10096,N_9679,N_9702);
nor U10097 (N_10097,N_9402,N_9631);
or U10098 (N_10098,N_9221,N_9486);
nand U10099 (N_10099,N_9341,N_9457);
nand U10100 (N_10100,N_9505,N_9608);
xor U10101 (N_10101,N_9229,N_9732);
nor U10102 (N_10102,N_9101,N_9395);
or U10103 (N_10103,N_9552,N_9618);
and U10104 (N_10104,N_9011,N_9338);
and U10105 (N_10105,N_9312,N_9513);
nor U10106 (N_10106,N_9438,N_9493);
or U10107 (N_10107,N_9277,N_9064);
nand U10108 (N_10108,N_9206,N_9550);
nand U10109 (N_10109,N_9670,N_9478);
xnor U10110 (N_10110,N_9380,N_9182);
nand U10111 (N_10111,N_9569,N_9677);
or U10112 (N_10112,N_9545,N_9439);
nand U10113 (N_10113,N_9236,N_9204);
nand U10114 (N_10114,N_9199,N_9019);
nand U10115 (N_10115,N_9697,N_9071);
or U10116 (N_10116,N_9336,N_9192);
xnor U10117 (N_10117,N_9036,N_9450);
or U10118 (N_10118,N_9188,N_9111);
and U10119 (N_10119,N_9626,N_9173);
or U10120 (N_10120,N_9477,N_9068);
and U10121 (N_10121,N_9389,N_9065);
and U10122 (N_10122,N_9254,N_9684);
nand U10123 (N_10123,N_9541,N_9042);
nand U10124 (N_10124,N_9508,N_9551);
nand U10125 (N_10125,N_9574,N_9258);
nor U10126 (N_10126,N_9385,N_9250);
nand U10127 (N_10127,N_9485,N_9258);
and U10128 (N_10128,N_9397,N_9476);
and U10129 (N_10129,N_9316,N_9680);
xnor U10130 (N_10130,N_9387,N_9291);
and U10131 (N_10131,N_9264,N_9631);
or U10132 (N_10132,N_9389,N_9354);
nor U10133 (N_10133,N_9053,N_9046);
xnor U10134 (N_10134,N_9247,N_9217);
nor U10135 (N_10135,N_9056,N_9648);
nor U10136 (N_10136,N_9200,N_9422);
nand U10137 (N_10137,N_9138,N_9315);
xor U10138 (N_10138,N_9055,N_9696);
and U10139 (N_10139,N_9555,N_9528);
nor U10140 (N_10140,N_9091,N_9348);
nor U10141 (N_10141,N_9720,N_9284);
or U10142 (N_10142,N_9691,N_9628);
nor U10143 (N_10143,N_9704,N_9709);
xnor U10144 (N_10144,N_9639,N_9019);
nand U10145 (N_10145,N_9208,N_9070);
or U10146 (N_10146,N_9478,N_9665);
or U10147 (N_10147,N_9243,N_9596);
nand U10148 (N_10148,N_9275,N_9461);
xor U10149 (N_10149,N_9192,N_9295);
xnor U10150 (N_10150,N_9203,N_9613);
xnor U10151 (N_10151,N_9254,N_9485);
or U10152 (N_10152,N_9088,N_9462);
or U10153 (N_10153,N_9465,N_9017);
and U10154 (N_10154,N_9034,N_9160);
and U10155 (N_10155,N_9649,N_9257);
xnor U10156 (N_10156,N_9294,N_9638);
xor U10157 (N_10157,N_9164,N_9560);
nor U10158 (N_10158,N_9679,N_9295);
nand U10159 (N_10159,N_9501,N_9040);
or U10160 (N_10160,N_9062,N_9574);
nor U10161 (N_10161,N_9654,N_9130);
xor U10162 (N_10162,N_9528,N_9346);
xor U10163 (N_10163,N_9308,N_9605);
and U10164 (N_10164,N_9312,N_9179);
nand U10165 (N_10165,N_9177,N_9551);
nand U10166 (N_10166,N_9069,N_9600);
nor U10167 (N_10167,N_9115,N_9568);
xnor U10168 (N_10168,N_9493,N_9171);
or U10169 (N_10169,N_9673,N_9746);
nand U10170 (N_10170,N_9066,N_9746);
and U10171 (N_10171,N_9022,N_9231);
or U10172 (N_10172,N_9571,N_9453);
nor U10173 (N_10173,N_9392,N_9282);
xnor U10174 (N_10174,N_9157,N_9722);
and U10175 (N_10175,N_9041,N_9241);
and U10176 (N_10176,N_9062,N_9174);
nor U10177 (N_10177,N_9158,N_9585);
nand U10178 (N_10178,N_9422,N_9507);
nand U10179 (N_10179,N_9306,N_9598);
xnor U10180 (N_10180,N_9233,N_9481);
xnor U10181 (N_10181,N_9417,N_9448);
or U10182 (N_10182,N_9015,N_9041);
xnor U10183 (N_10183,N_9144,N_9301);
xor U10184 (N_10184,N_9244,N_9011);
or U10185 (N_10185,N_9280,N_9688);
or U10186 (N_10186,N_9331,N_9648);
or U10187 (N_10187,N_9487,N_9211);
nor U10188 (N_10188,N_9748,N_9596);
nand U10189 (N_10189,N_9619,N_9098);
or U10190 (N_10190,N_9281,N_9456);
and U10191 (N_10191,N_9232,N_9242);
xor U10192 (N_10192,N_9394,N_9040);
nor U10193 (N_10193,N_9305,N_9162);
or U10194 (N_10194,N_9560,N_9382);
nor U10195 (N_10195,N_9006,N_9233);
nor U10196 (N_10196,N_9157,N_9378);
nand U10197 (N_10197,N_9203,N_9571);
or U10198 (N_10198,N_9363,N_9465);
or U10199 (N_10199,N_9369,N_9506);
nor U10200 (N_10200,N_9482,N_9703);
nor U10201 (N_10201,N_9065,N_9554);
and U10202 (N_10202,N_9150,N_9568);
and U10203 (N_10203,N_9501,N_9236);
or U10204 (N_10204,N_9493,N_9702);
or U10205 (N_10205,N_9185,N_9616);
and U10206 (N_10206,N_9009,N_9081);
xnor U10207 (N_10207,N_9599,N_9209);
nand U10208 (N_10208,N_9677,N_9224);
and U10209 (N_10209,N_9215,N_9403);
or U10210 (N_10210,N_9226,N_9116);
xor U10211 (N_10211,N_9369,N_9645);
and U10212 (N_10212,N_9722,N_9360);
and U10213 (N_10213,N_9388,N_9331);
nor U10214 (N_10214,N_9658,N_9379);
xor U10215 (N_10215,N_9578,N_9382);
nor U10216 (N_10216,N_9721,N_9188);
nand U10217 (N_10217,N_9274,N_9113);
xnor U10218 (N_10218,N_9654,N_9607);
or U10219 (N_10219,N_9694,N_9719);
xor U10220 (N_10220,N_9155,N_9285);
xor U10221 (N_10221,N_9720,N_9241);
nor U10222 (N_10222,N_9486,N_9659);
or U10223 (N_10223,N_9210,N_9240);
and U10224 (N_10224,N_9354,N_9037);
nor U10225 (N_10225,N_9556,N_9384);
nor U10226 (N_10226,N_9473,N_9236);
or U10227 (N_10227,N_9289,N_9184);
and U10228 (N_10228,N_9547,N_9579);
and U10229 (N_10229,N_9243,N_9138);
xnor U10230 (N_10230,N_9068,N_9510);
nor U10231 (N_10231,N_9483,N_9343);
and U10232 (N_10232,N_9651,N_9616);
or U10233 (N_10233,N_9666,N_9316);
nor U10234 (N_10234,N_9671,N_9517);
and U10235 (N_10235,N_9525,N_9063);
xnor U10236 (N_10236,N_9202,N_9643);
or U10237 (N_10237,N_9048,N_9224);
or U10238 (N_10238,N_9330,N_9509);
or U10239 (N_10239,N_9173,N_9192);
or U10240 (N_10240,N_9545,N_9337);
xor U10241 (N_10241,N_9721,N_9586);
and U10242 (N_10242,N_9353,N_9081);
nand U10243 (N_10243,N_9007,N_9522);
nand U10244 (N_10244,N_9613,N_9691);
or U10245 (N_10245,N_9244,N_9729);
nand U10246 (N_10246,N_9117,N_9328);
xor U10247 (N_10247,N_9599,N_9468);
and U10248 (N_10248,N_9225,N_9171);
or U10249 (N_10249,N_9467,N_9043);
and U10250 (N_10250,N_9206,N_9544);
or U10251 (N_10251,N_9347,N_9236);
and U10252 (N_10252,N_9560,N_9653);
or U10253 (N_10253,N_9158,N_9690);
nand U10254 (N_10254,N_9581,N_9495);
nor U10255 (N_10255,N_9318,N_9546);
and U10256 (N_10256,N_9478,N_9659);
or U10257 (N_10257,N_9250,N_9666);
and U10258 (N_10258,N_9232,N_9019);
nor U10259 (N_10259,N_9407,N_9419);
nor U10260 (N_10260,N_9521,N_9030);
or U10261 (N_10261,N_9103,N_9326);
or U10262 (N_10262,N_9735,N_9138);
or U10263 (N_10263,N_9532,N_9308);
nor U10264 (N_10264,N_9622,N_9007);
or U10265 (N_10265,N_9212,N_9078);
and U10266 (N_10266,N_9321,N_9185);
and U10267 (N_10267,N_9206,N_9690);
nand U10268 (N_10268,N_9202,N_9629);
nor U10269 (N_10269,N_9383,N_9164);
xnor U10270 (N_10270,N_9003,N_9552);
xor U10271 (N_10271,N_9581,N_9293);
nor U10272 (N_10272,N_9676,N_9018);
xnor U10273 (N_10273,N_9701,N_9397);
xnor U10274 (N_10274,N_9591,N_9561);
xnor U10275 (N_10275,N_9471,N_9643);
or U10276 (N_10276,N_9060,N_9368);
and U10277 (N_10277,N_9655,N_9400);
xnor U10278 (N_10278,N_9735,N_9707);
nor U10279 (N_10279,N_9353,N_9431);
nand U10280 (N_10280,N_9386,N_9547);
or U10281 (N_10281,N_9182,N_9745);
nor U10282 (N_10282,N_9389,N_9721);
and U10283 (N_10283,N_9353,N_9567);
nor U10284 (N_10284,N_9423,N_9333);
xor U10285 (N_10285,N_9723,N_9720);
xor U10286 (N_10286,N_9431,N_9524);
and U10287 (N_10287,N_9637,N_9003);
xnor U10288 (N_10288,N_9734,N_9270);
nor U10289 (N_10289,N_9153,N_9501);
and U10290 (N_10290,N_9570,N_9621);
xor U10291 (N_10291,N_9437,N_9665);
nand U10292 (N_10292,N_9300,N_9423);
nor U10293 (N_10293,N_9388,N_9025);
or U10294 (N_10294,N_9274,N_9071);
nand U10295 (N_10295,N_9016,N_9019);
or U10296 (N_10296,N_9109,N_9086);
nor U10297 (N_10297,N_9420,N_9564);
nor U10298 (N_10298,N_9397,N_9321);
nor U10299 (N_10299,N_9081,N_9101);
nor U10300 (N_10300,N_9028,N_9679);
xnor U10301 (N_10301,N_9712,N_9258);
nor U10302 (N_10302,N_9609,N_9239);
xor U10303 (N_10303,N_9182,N_9441);
nand U10304 (N_10304,N_9277,N_9161);
and U10305 (N_10305,N_9605,N_9043);
nand U10306 (N_10306,N_9421,N_9516);
nor U10307 (N_10307,N_9317,N_9721);
or U10308 (N_10308,N_9743,N_9687);
nand U10309 (N_10309,N_9480,N_9278);
and U10310 (N_10310,N_9417,N_9009);
or U10311 (N_10311,N_9616,N_9552);
xor U10312 (N_10312,N_9645,N_9105);
and U10313 (N_10313,N_9373,N_9123);
nor U10314 (N_10314,N_9734,N_9579);
nor U10315 (N_10315,N_9677,N_9710);
and U10316 (N_10316,N_9747,N_9607);
and U10317 (N_10317,N_9173,N_9226);
or U10318 (N_10318,N_9482,N_9370);
xnor U10319 (N_10319,N_9243,N_9207);
xor U10320 (N_10320,N_9373,N_9678);
xor U10321 (N_10321,N_9532,N_9254);
and U10322 (N_10322,N_9170,N_9112);
and U10323 (N_10323,N_9595,N_9021);
xor U10324 (N_10324,N_9407,N_9249);
nor U10325 (N_10325,N_9585,N_9083);
nand U10326 (N_10326,N_9253,N_9558);
and U10327 (N_10327,N_9574,N_9455);
nand U10328 (N_10328,N_9653,N_9354);
or U10329 (N_10329,N_9130,N_9626);
nand U10330 (N_10330,N_9219,N_9658);
xnor U10331 (N_10331,N_9283,N_9518);
and U10332 (N_10332,N_9414,N_9337);
xor U10333 (N_10333,N_9364,N_9030);
and U10334 (N_10334,N_9445,N_9501);
xor U10335 (N_10335,N_9707,N_9020);
xor U10336 (N_10336,N_9350,N_9321);
nand U10337 (N_10337,N_9401,N_9442);
nor U10338 (N_10338,N_9020,N_9503);
nand U10339 (N_10339,N_9598,N_9180);
nor U10340 (N_10340,N_9265,N_9400);
xnor U10341 (N_10341,N_9508,N_9482);
xnor U10342 (N_10342,N_9458,N_9409);
xor U10343 (N_10343,N_9065,N_9132);
xnor U10344 (N_10344,N_9296,N_9305);
or U10345 (N_10345,N_9204,N_9437);
or U10346 (N_10346,N_9528,N_9255);
nor U10347 (N_10347,N_9125,N_9593);
or U10348 (N_10348,N_9194,N_9516);
nand U10349 (N_10349,N_9146,N_9269);
or U10350 (N_10350,N_9639,N_9141);
nor U10351 (N_10351,N_9274,N_9719);
nand U10352 (N_10352,N_9236,N_9349);
or U10353 (N_10353,N_9057,N_9745);
and U10354 (N_10354,N_9058,N_9264);
or U10355 (N_10355,N_9607,N_9255);
or U10356 (N_10356,N_9220,N_9403);
or U10357 (N_10357,N_9649,N_9532);
and U10358 (N_10358,N_9449,N_9153);
nand U10359 (N_10359,N_9220,N_9410);
xor U10360 (N_10360,N_9287,N_9737);
xnor U10361 (N_10361,N_9088,N_9365);
nand U10362 (N_10362,N_9321,N_9388);
nand U10363 (N_10363,N_9397,N_9120);
xor U10364 (N_10364,N_9664,N_9557);
and U10365 (N_10365,N_9143,N_9286);
xnor U10366 (N_10366,N_9314,N_9696);
xnor U10367 (N_10367,N_9555,N_9447);
xnor U10368 (N_10368,N_9477,N_9283);
and U10369 (N_10369,N_9290,N_9521);
nor U10370 (N_10370,N_9647,N_9185);
nand U10371 (N_10371,N_9747,N_9576);
nor U10372 (N_10372,N_9213,N_9562);
or U10373 (N_10373,N_9105,N_9361);
and U10374 (N_10374,N_9696,N_9394);
or U10375 (N_10375,N_9026,N_9717);
or U10376 (N_10376,N_9411,N_9572);
xnor U10377 (N_10377,N_9374,N_9093);
nor U10378 (N_10378,N_9108,N_9730);
xor U10379 (N_10379,N_9107,N_9421);
xor U10380 (N_10380,N_9214,N_9360);
xnor U10381 (N_10381,N_9473,N_9498);
xor U10382 (N_10382,N_9245,N_9087);
nand U10383 (N_10383,N_9674,N_9361);
or U10384 (N_10384,N_9014,N_9407);
or U10385 (N_10385,N_9384,N_9545);
nor U10386 (N_10386,N_9526,N_9239);
or U10387 (N_10387,N_9177,N_9593);
nand U10388 (N_10388,N_9309,N_9689);
or U10389 (N_10389,N_9583,N_9091);
nor U10390 (N_10390,N_9422,N_9078);
and U10391 (N_10391,N_9528,N_9526);
nand U10392 (N_10392,N_9495,N_9263);
or U10393 (N_10393,N_9212,N_9463);
xor U10394 (N_10394,N_9047,N_9706);
nor U10395 (N_10395,N_9613,N_9673);
or U10396 (N_10396,N_9687,N_9564);
xor U10397 (N_10397,N_9577,N_9382);
xnor U10398 (N_10398,N_9126,N_9026);
or U10399 (N_10399,N_9382,N_9426);
or U10400 (N_10400,N_9263,N_9503);
or U10401 (N_10401,N_9125,N_9500);
and U10402 (N_10402,N_9370,N_9303);
nand U10403 (N_10403,N_9707,N_9357);
xor U10404 (N_10404,N_9669,N_9716);
or U10405 (N_10405,N_9748,N_9244);
and U10406 (N_10406,N_9157,N_9018);
or U10407 (N_10407,N_9498,N_9067);
and U10408 (N_10408,N_9099,N_9079);
and U10409 (N_10409,N_9326,N_9315);
xor U10410 (N_10410,N_9070,N_9028);
and U10411 (N_10411,N_9537,N_9723);
nor U10412 (N_10412,N_9627,N_9539);
nor U10413 (N_10413,N_9007,N_9515);
nor U10414 (N_10414,N_9569,N_9453);
and U10415 (N_10415,N_9022,N_9045);
and U10416 (N_10416,N_9340,N_9178);
or U10417 (N_10417,N_9275,N_9707);
xor U10418 (N_10418,N_9271,N_9520);
xor U10419 (N_10419,N_9641,N_9183);
or U10420 (N_10420,N_9318,N_9527);
and U10421 (N_10421,N_9113,N_9345);
xnor U10422 (N_10422,N_9394,N_9469);
or U10423 (N_10423,N_9235,N_9406);
nand U10424 (N_10424,N_9116,N_9308);
and U10425 (N_10425,N_9666,N_9034);
or U10426 (N_10426,N_9328,N_9485);
and U10427 (N_10427,N_9278,N_9051);
nand U10428 (N_10428,N_9109,N_9525);
nor U10429 (N_10429,N_9118,N_9094);
and U10430 (N_10430,N_9043,N_9257);
nor U10431 (N_10431,N_9048,N_9193);
nand U10432 (N_10432,N_9492,N_9232);
nand U10433 (N_10433,N_9324,N_9196);
nand U10434 (N_10434,N_9483,N_9647);
or U10435 (N_10435,N_9259,N_9390);
and U10436 (N_10436,N_9141,N_9507);
xor U10437 (N_10437,N_9267,N_9091);
and U10438 (N_10438,N_9403,N_9171);
xnor U10439 (N_10439,N_9271,N_9455);
nor U10440 (N_10440,N_9660,N_9140);
xnor U10441 (N_10441,N_9234,N_9040);
and U10442 (N_10442,N_9076,N_9320);
and U10443 (N_10443,N_9673,N_9093);
nor U10444 (N_10444,N_9332,N_9394);
xor U10445 (N_10445,N_9010,N_9056);
nand U10446 (N_10446,N_9004,N_9330);
and U10447 (N_10447,N_9227,N_9608);
or U10448 (N_10448,N_9434,N_9637);
nand U10449 (N_10449,N_9015,N_9632);
or U10450 (N_10450,N_9695,N_9103);
or U10451 (N_10451,N_9023,N_9548);
xnor U10452 (N_10452,N_9431,N_9097);
or U10453 (N_10453,N_9429,N_9057);
nand U10454 (N_10454,N_9492,N_9367);
and U10455 (N_10455,N_9251,N_9022);
nor U10456 (N_10456,N_9698,N_9186);
nor U10457 (N_10457,N_9326,N_9616);
xnor U10458 (N_10458,N_9093,N_9271);
and U10459 (N_10459,N_9017,N_9318);
or U10460 (N_10460,N_9359,N_9069);
nor U10461 (N_10461,N_9443,N_9508);
or U10462 (N_10462,N_9552,N_9279);
or U10463 (N_10463,N_9432,N_9100);
nor U10464 (N_10464,N_9240,N_9304);
nand U10465 (N_10465,N_9689,N_9538);
nand U10466 (N_10466,N_9667,N_9662);
xor U10467 (N_10467,N_9087,N_9509);
xor U10468 (N_10468,N_9032,N_9573);
or U10469 (N_10469,N_9048,N_9276);
xnor U10470 (N_10470,N_9353,N_9086);
or U10471 (N_10471,N_9563,N_9133);
and U10472 (N_10472,N_9090,N_9180);
nor U10473 (N_10473,N_9072,N_9548);
nor U10474 (N_10474,N_9176,N_9510);
nor U10475 (N_10475,N_9354,N_9341);
and U10476 (N_10476,N_9577,N_9593);
nand U10477 (N_10477,N_9605,N_9637);
nand U10478 (N_10478,N_9180,N_9278);
and U10479 (N_10479,N_9383,N_9624);
and U10480 (N_10480,N_9322,N_9557);
or U10481 (N_10481,N_9538,N_9744);
or U10482 (N_10482,N_9213,N_9441);
nand U10483 (N_10483,N_9031,N_9511);
and U10484 (N_10484,N_9318,N_9207);
or U10485 (N_10485,N_9598,N_9411);
xor U10486 (N_10486,N_9011,N_9383);
and U10487 (N_10487,N_9350,N_9559);
or U10488 (N_10488,N_9717,N_9071);
nand U10489 (N_10489,N_9302,N_9559);
nand U10490 (N_10490,N_9237,N_9276);
or U10491 (N_10491,N_9740,N_9569);
nor U10492 (N_10492,N_9553,N_9173);
or U10493 (N_10493,N_9581,N_9029);
or U10494 (N_10494,N_9724,N_9316);
nand U10495 (N_10495,N_9505,N_9185);
or U10496 (N_10496,N_9083,N_9264);
nor U10497 (N_10497,N_9270,N_9032);
nand U10498 (N_10498,N_9383,N_9297);
xnor U10499 (N_10499,N_9533,N_9044);
xnor U10500 (N_10500,N_10446,N_9961);
xnor U10501 (N_10501,N_9990,N_10073);
nand U10502 (N_10502,N_10003,N_10028);
nor U10503 (N_10503,N_10230,N_10475);
xor U10504 (N_10504,N_9837,N_10265);
and U10505 (N_10505,N_10032,N_9822);
nand U10506 (N_10506,N_10306,N_10043);
xor U10507 (N_10507,N_9907,N_10431);
and U10508 (N_10508,N_9908,N_10137);
or U10509 (N_10509,N_10372,N_9888);
or U10510 (N_10510,N_10423,N_10388);
nand U10511 (N_10511,N_9813,N_9835);
xnor U10512 (N_10512,N_9989,N_10232);
nor U10513 (N_10513,N_9899,N_10392);
or U10514 (N_10514,N_10381,N_10396);
nand U10515 (N_10515,N_10052,N_10261);
nor U10516 (N_10516,N_10143,N_10207);
or U10517 (N_10517,N_10377,N_9890);
or U10518 (N_10518,N_10116,N_10068);
or U10519 (N_10519,N_10435,N_10304);
xor U10520 (N_10520,N_9828,N_10309);
nand U10521 (N_10521,N_9911,N_9993);
nand U10522 (N_10522,N_10468,N_10141);
xnor U10523 (N_10523,N_9849,N_10453);
xor U10524 (N_10524,N_10273,N_10194);
and U10525 (N_10525,N_10231,N_10237);
or U10526 (N_10526,N_10411,N_10002);
or U10527 (N_10527,N_10144,N_10358);
xnor U10528 (N_10528,N_9992,N_10177);
or U10529 (N_10529,N_10181,N_9987);
nand U10530 (N_10530,N_10399,N_10338);
nor U10531 (N_10531,N_10121,N_10406);
nor U10532 (N_10532,N_9998,N_10478);
nand U10533 (N_10533,N_10488,N_10152);
xor U10534 (N_10534,N_10375,N_10100);
or U10535 (N_10535,N_9980,N_10397);
nand U10536 (N_10536,N_9824,N_9827);
nand U10537 (N_10537,N_10102,N_9750);
or U10538 (N_10538,N_10015,N_9756);
and U10539 (N_10539,N_9875,N_10366);
or U10540 (N_10540,N_10112,N_10291);
xor U10541 (N_10541,N_9877,N_9859);
and U10542 (N_10542,N_10487,N_10029);
xnor U10543 (N_10543,N_9816,N_9785);
xnor U10544 (N_10544,N_10492,N_9969);
xor U10545 (N_10545,N_10420,N_9767);
nand U10546 (N_10546,N_10202,N_10120);
and U10547 (N_10547,N_10283,N_10184);
nand U10548 (N_10548,N_9820,N_10463);
nand U10549 (N_10549,N_9852,N_10499);
nor U10550 (N_10550,N_10437,N_10038);
nor U10551 (N_10551,N_9838,N_10424);
xnor U10552 (N_10552,N_10319,N_10074);
xor U10553 (N_10553,N_10408,N_10404);
or U10554 (N_10554,N_9800,N_10233);
and U10555 (N_10555,N_10425,N_10157);
nand U10556 (N_10556,N_10327,N_10089);
nand U10557 (N_10557,N_10361,N_10307);
or U10558 (N_10558,N_10215,N_10268);
nor U10559 (N_10559,N_9842,N_10274);
nor U10560 (N_10560,N_10452,N_10042);
xnor U10561 (N_10561,N_10407,N_10403);
or U10562 (N_10562,N_10082,N_9757);
xnor U10563 (N_10563,N_10386,N_10359);
nor U10564 (N_10564,N_9830,N_10454);
nand U10565 (N_10565,N_10337,N_9878);
nor U10566 (N_10566,N_9836,N_10287);
xnor U10567 (N_10567,N_9894,N_10278);
nand U10568 (N_10568,N_10191,N_10033);
or U10569 (N_10569,N_10223,N_9900);
and U10570 (N_10570,N_10438,N_9979);
nand U10571 (N_10571,N_10224,N_10021);
nor U10572 (N_10572,N_10410,N_10115);
and U10573 (N_10573,N_10395,N_9766);
xor U10574 (N_10574,N_9944,N_10227);
xnor U10575 (N_10575,N_9893,N_10185);
or U10576 (N_10576,N_9973,N_10483);
or U10577 (N_10577,N_9862,N_10260);
and U10578 (N_10578,N_9910,N_10365);
xnor U10579 (N_10579,N_10456,N_10014);
nor U10580 (N_10580,N_10040,N_10256);
nand U10581 (N_10581,N_9833,N_9909);
and U10582 (N_10582,N_9886,N_9929);
xor U10583 (N_10583,N_10344,N_10330);
or U10584 (N_10584,N_9755,N_9902);
nor U10585 (N_10585,N_9947,N_9951);
nor U10586 (N_10586,N_10351,N_10302);
nand U10587 (N_10587,N_10443,N_10203);
nor U10588 (N_10588,N_10083,N_10469);
and U10589 (N_10589,N_10432,N_10434);
nor U10590 (N_10590,N_10051,N_10449);
xor U10591 (N_10591,N_9896,N_10091);
and U10592 (N_10592,N_10213,N_10098);
xnor U10593 (N_10593,N_9945,N_10335);
nand U10594 (N_10594,N_10197,N_10336);
nand U10595 (N_10595,N_10226,N_10168);
xnor U10596 (N_10596,N_10229,N_10109);
nor U10597 (N_10597,N_10360,N_9781);
and U10598 (N_10598,N_9866,N_10059);
or U10599 (N_10599,N_9801,N_10315);
nor U10600 (N_10600,N_10228,N_10034);
xnor U10601 (N_10601,N_10379,N_10225);
xor U10602 (N_10602,N_10380,N_9834);
nand U10603 (N_10603,N_10093,N_10142);
or U10604 (N_10604,N_10331,N_9790);
nor U10605 (N_10605,N_9782,N_10371);
xnor U10606 (N_10606,N_10356,N_9794);
nor U10607 (N_10607,N_9791,N_10005);
nor U10608 (N_10608,N_10076,N_9956);
nand U10609 (N_10609,N_9788,N_9832);
or U10610 (N_10610,N_10317,N_10138);
and U10611 (N_10611,N_10297,N_10470);
xnor U10612 (N_10612,N_9936,N_9793);
nor U10613 (N_10613,N_9920,N_9772);
nand U10614 (N_10614,N_10054,N_10201);
nor U10615 (N_10615,N_10486,N_10106);
or U10616 (N_10616,N_9864,N_10087);
nand U10617 (N_10617,N_10279,N_10219);
or U10618 (N_10618,N_10349,N_10390);
or U10619 (N_10619,N_9986,N_9871);
nand U10620 (N_10620,N_10246,N_9943);
nand U10621 (N_10621,N_9759,N_10122);
or U10622 (N_10622,N_10347,N_10192);
and U10623 (N_10623,N_9983,N_10310);
or U10624 (N_10624,N_10345,N_10149);
nor U10625 (N_10625,N_10130,N_9777);
nor U10626 (N_10626,N_10060,N_10174);
nand U10627 (N_10627,N_10162,N_10267);
xnor U10628 (N_10628,N_9839,N_10393);
xor U10629 (N_10629,N_10173,N_10286);
nor U10630 (N_10630,N_10497,N_10333);
xor U10631 (N_10631,N_9985,N_10472);
nor U10632 (N_10632,N_10064,N_10282);
xnor U10633 (N_10633,N_9825,N_10176);
nand U10634 (N_10634,N_10266,N_10164);
nand U10635 (N_10635,N_10293,N_10303);
nor U10636 (N_10636,N_10494,N_9970);
or U10637 (N_10637,N_10113,N_10378);
xor U10638 (N_10638,N_10458,N_10242);
and U10639 (N_10639,N_10257,N_10247);
and U10640 (N_10640,N_10325,N_10264);
and U10641 (N_10641,N_9857,N_10476);
nor U10642 (N_10642,N_10161,N_10128);
xnor U10643 (N_10643,N_10166,N_10394);
nand U10644 (N_10644,N_10180,N_9982);
and U10645 (N_10645,N_10046,N_10323);
and U10646 (N_10646,N_10030,N_9972);
nor U10647 (N_10647,N_9975,N_10415);
nand U10648 (N_10648,N_9991,N_10004);
or U10649 (N_10649,N_9764,N_9974);
nand U10650 (N_10650,N_9758,N_9905);
xor U10651 (N_10651,N_9829,N_9776);
or U10652 (N_10652,N_10471,N_9976);
nand U10653 (N_10653,N_9798,N_10439);
nand U10654 (N_10654,N_9805,N_10474);
nand U10655 (N_10655,N_10295,N_9814);
xor U10656 (N_10656,N_10496,N_10172);
nor U10657 (N_10657,N_10284,N_10117);
and U10658 (N_10658,N_10491,N_10084);
xnor U10659 (N_10659,N_9754,N_10000);
nor U10660 (N_10660,N_10444,N_9809);
and U10661 (N_10661,N_10313,N_10234);
nand U10662 (N_10662,N_10455,N_10036);
or U10663 (N_10663,N_9752,N_10401);
or U10664 (N_10664,N_10460,N_10362);
and U10665 (N_10665,N_10254,N_9901);
or U10666 (N_10666,N_10127,N_10175);
nor U10667 (N_10667,N_10367,N_10158);
nor U10668 (N_10668,N_10037,N_10334);
or U10669 (N_10669,N_10414,N_9846);
and U10670 (N_10670,N_9861,N_10412);
xnor U10671 (N_10671,N_10357,N_9880);
or U10672 (N_10672,N_9796,N_9806);
and U10673 (N_10673,N_9942,N_9760);
or U10674 (N_10674,N_9981,N_9912);
or U10675 (N_10675,N_10096,N_10479);
xnor U10676 (N_10676,N_10305,N_9853);
or U10677 (N_10677,N_9867,N_9803);
nand U10678 (N_10678,N_9950,N_10243);
or U10679 (N_10679,N_10067,N_10277);
or U10680 (N_10680,N_10241,N_9918);
nor U10681 (N_10681,N_9787,N_10457);
nor U10682 (N_10682,N_10238,N_10354);
xnor U10683 (N_10683,N_9784,N_10169);
and U10684 (N_10684,N_10348,N_10353);
nor U10685 (N_10685,N_10222,N_9818);
and U10686 (N_10686,N_10490,N_10035);
nor U10687 (N_10687,N_10342,N_10442);
or U10688 (N_10688,N_9843,N_9921);
nor U10689 (N_10689,N_10465,N_9768);
nand U10690 (N_10690,N_9999,N_10045);
or U10691 (N_10691,N_10298,N_10248);
nor U10692 (N_10692,N_10069,N_9799);
nand U10693 (N_10693,N_10085,N_9812);
nor U10694 (N_10694,N_9962,N_10409);
nand U10695 (N_10695,N_10467,N_10466);
nand U10696 (N_10696,N_9977,N_10332);
or U10697 (N_10697,N_10146,N_10053);
or U10698 (N_10698,N_10462,N_10376);
nand U10699 (N_10699,N_10387,N_10077);
nor U10700 (N_10700,N_9876,N_10016);
xnor U10701 (N_10701,N_10373,N_10339);
and U10702 (N_10702,N_10204,N_10178);
nand U10703 (N_10703,N_10391,N_9939);
or U10704 (N_10704,N_9810,N_9882);
xnor U10705 (N_10705,N_10495,N_9775);
and U10706 (N_10706,N_10405,N_10153);
or U10707 (N_10707,N_9844,N_9953);
or U10708 (N_10708,N_9913,N_9955);
nand U10709 (N_10709,N_10118,N_9994);
or U10710 (N_10710,N_9996,N_10057);
and U10711 (N_10711,N_10114,N_10189);
nor U10712 (N_10712,N_10131,N_10383);
or U10713 (N_10713,N_10272,N_9786);
nor U10714 (N_10714,N_9949,N_10363);
nand U10715 (N_10715,N_10428,N_9968);
xor U10716 (N_10716,N_10433,N_9915);
xnor U10717 (N_10717,N_10062,N_9863);
or U10718 (N_10718,N_10436,N_10123);
or U10719 (N_10719,N_9840,N_9797);
nand U10720 (N_10720,N_10430,N_9940);
xor U10721 (N_10721,N_10159,N_9978);
or U10722 (N_10722,N_10321,N_9897);
and U10723 (N_10723,N_10183,N_10125);
and U10724 (N_10724,N_10165,N_10056);
xnor U10725 (N_10725,N_9826,N_10450);
nand U10726 (N_10726,N_9967,N_10218);
or U10727 (N_10727,N_10111,N_10013);
or U10728 (N_10728,N_10210,N_9763);
or U10729 (N_10729,N_10316,N_10290);
nand U10730 (N_10730,N_10245,N_10417);
nand U10731 (N_10731,N_10079,N_9971);
and U10732 (N_10732,N_9779,N_10018);
or U10733 (N_10733,N_10448,N_10099);
or U10734 (N_10734,N_10092,N_9958);
nor U10735 (N_10735,N_9879,N_10095);
xor U10736 (N_10736,N_9938,N_10097);
xor U10737 (N_10737,N_10292,N_9845);
and U10738 (N_10738,N_10285,N_10044);
nand U10739 (N_10739,N_9895,N_9765);
nand U10740 (N_10740,N_10078,N_9869);
and U10741 (N_10741,N_10101,N_10355);
nand U10742 (N_10742,N_10107,N_10239);
nor U10743 (N_10743,N_9906,N_10413);
nor U10744 (N_10744,N_10384,N_10094);
xor U10745 (N_10745,N_10294,N_10447);
nand U10746 (N_10746,N_10020,N_10048);
and U10747 (N_10747,N_9904,N_10063);
and U10748 (N_10748,N_10271,N_10244);
nor U10749 (N_10749,N_9963,N_10024);
or U10750 (N_10750,N_9817,N_9946);
xnor U10751 (N_10751,N_9925,N_10350);
nand U10752 (N_10752,N_10179,N_10385);
or U10753 (N_10753,N_9934,N_10135);
xnor U10754 (N_10754,N_10459,N_10477);
nor U10755 (N_10755,N_9770,N_10281);
nand U10756 (N_10756,N_9923,N_9995);
or U10757 (N_10757,N_10484,N_10221);
and U10758 (N_10758,N_10429,N_10236);
xor U10759 (N_10759,N_9917,N_10108);
nand U10760 (N_10760,N_10427,N_10012);
nor U10761 (N_10761,N_10193,N_9930);
nand U10762 (N_10762,N_9773,N_10262);
xor U10763 (N_10763,N_10133,N_10498);
and U10764 (N_10764,N_9850,N_10145);
nand U10765 (N_10765,N_10216,N_10163);
nor U10766 (N_10766,N_10217,N_10481);
xnor U10767 (N_10767,N_10352,N_10473);
nand U10768 (N_10768,N_10055,N_10289);
nand U10769 (N_10769,N_10370,N_10081);
nor U10770 (N_10770,N_10017,N_10329);
nand U10771 (N_10771,N_10025,N_10212);
or U10772 (N_10772,N_9965,N_10151);
or U10773 (N_10773,N_9997,N_9960);
or U10774 (N_10774,N_10160,N_9935);
xor U10775 (N_10775,N_9892,N_10209);
or U10776 (N_10776,N_9789,N_9858);
nor U10777 (N_10777,N_9933,N_10341);
nor U10778 (N_10778,N_9924,N_10326);
nand U10779 (N_10779,N_10461,N_10250);
nand U10780 (N_10780,N_10186,N_9881);
xor U10781 (N_10781,N_10312,N_9964);
xnor U10782 (N_10782,N_9780,N_10105);
and U10783 (N_10783,N_10196,N_9762);
xnor U10784 (N_10784,N_9874,N_9870);
nor U10785 (N_10785,N_10010,N_10253);
and U10786 (N_10786,N_10199,N_9926);
or U10787 (N_10787,N_10426,N_10156);
nor U10788 (N_10788,N_10311,N_10322);
and U10789 (N_10789,N_9761,N_10065);
or U10790 (N_10790,N_10182,N_9753);
nand U10791 (N_10791,N_9841,N_9823);
and U10792 (N_10792,N_9804,N_9831);
and U10793 (N_10793,N_10006,N_9855);
nand U10794 (N_10794,N_9966,N_10140);
nand U10795 (N_10795,N_10263,N_10080);
nor U10796 (N_10796,N_9860,N_10270);
xnor U10797 (N_10797,N_10419,N_10255);
nand U10798 (N_10798,N_10314,N_10155);
nand U10799 (N_10799,N_10187,N_9807);
nor U10800 (N_10800,N_10072,N_9815);
and U10801 (N_10801,N_9872,N_9821);
xor U10802 (N_10802,N_9889,N_9811);
nand U10803 (N_10803,N_9922,N_10343);
xnor U10804 (N_10804,N_10061,N_10023);
or U10805 (N_10805,N_9927,N_10464);
xor U10806 (N_10806,N_10009,N_10440);
nand U10807 (N_10807,N_9948,N_9795);
or U10808 (N_10808,N_10208,N_10259);
or U10809 (N_10809,N_9883,N_9819);
or U10810 (N_10810,N_9937,N_10318);
nor U10811 (N_10811,N_10027,N_9916);
nor U10812 (N_10812,N_9984,N_9931);
xor U10813 (N_10813,N_9865,N_9751);
and U10814 (N_10814,N_10480,N_10276);
nor U10815 (N_10815,N_9959,N_10170);
xnor U10816 (N_10816,N_10041,N_10132);
or U10817 (N_10817,N_9988,N_10058);
xnor U10818 (N_10818,N_10301,N_10167);
nand U10819 (N_10819,N_10129,N_9914);
or U10820 (N_10820,N_10139,N_10198);
and U10821 (N_10821,N_9778,N_10019);
and U10822 (N_10822,N_10150,N_10493);
and U10823 (N_10823,N_9847,N_10451);
or U10824 (N_10824,N_10328,N_10240);
nor U10825 (N_10825,N_9941,N_10104);
nor U10826 (N_10826,N_10200,N_9771);
or U10827 (N_10827,N_10489,N_10211);
and U10828 (N_10828,N_9919,N_10007);
and U10829 (N_10829,N_10421,N_10346);
and U10830 (N_10830,N_10258,N_9928);
xor U10831 (N_10831,N_10485,N_10088);
nand U10832 (N_10832,N_10011,N_10280);
nand U10833 (N_10833,N_10206,N_9873);
and U10834 (N_10834,N_10445,N_10374);
xnor U10835 (N_10835,N_10382,N_10368);
or U10836 (N_10836,N_10148,N_10103);
xor U10837 (N_10837,N_10275,N_9898);
nand U10838 (N_10838,N_10075,N_10050);
nand U10839 (N_10839,N_10086,N_10205);
nand U10840 (N_10840,N_10190,N_10220);
nand U10841 (N_10841,N_10369,N_10071);
and U10842 (N_10842,N_9851,N_9903);
or U10843 (N_10843,N_10299,N_10249);
or U10844 (N_10844,N_10235,N_10134);
nor U10845 (N_10845,N_10441,N_9783);
nor U10846 (N_10846,N_10008,N_10214);
and U10847 (N_10847,N_9848,N_9891);
nor U10848 (N_10848,N_9885,N_10300);
and U10849 (N_10849,N_10188,N_10269);
nor U10850 (N_10850,N_10416,N_10022);
xnor U10851 (N_10851,N_10400,N_9868);
or U10852 (N_10852,N_10288,N_10110);
or U10853 (N_10853,N_9854,N_9954);
nand U10854 (N_10854,N_10340,N_9792);
xor U10855 (N_10855,N_10154,N_10171);
nor U10856 (N_10856,N_10389,N_10039);
and U10857 (N_10857,N_9802,N_10001);
xor U10858 (N_10858,N_9884,N_10136);
or U10859 (N_10859,N_9887,N_9774);
nor U10860 (N_10860,N_10026,N_9932);
nor U10861 (N_10861,N_10296,N_9856);
or U10862 (N_10862,N_10126,N_10308);
nor U10863 (N_10863,N_9952,N_9769);
xnor U10864 (N_10864,N_10320,N_10031);
or U10865 (N_10865,N_10147,N_9808);
xnor U10866 (N_10866,N_10324,N_10124);
or U10867 (N_10867,N_10047,N_10195);
or U10868 (N_10868,N_10066,N_10422);
and U10869 (N_10869,N_10049,N_10418);
nor U10870 (N_10870,N_10398,N_10402);
nand U10871 (N_10871,N_10252,N_10090);
nand U10872 (N_10872,N_10251,N_10119);
or U10873 (N_10873,N_9957,N_10364);
nor U10874 (N_10874,N_10070,N_10482);
nand U10875 (N_10875,N_10086,N_10319);
nand U10876 (N_10876,N_10201,N_10358);
nor U10877 (N_10877,N_10043,N_10090);
xnor U10878 (N_10878,N_10390,N_9860);
xor U10879 (N_10879,N_10279,N_10101);
and U10880 (N_10880,N_10260,N_10387);
or U10881 (N_10881,N_10121,N_10090);
xor U10882 (N_10882,N_10418,N_10467);
xor U10883 (N_10883,N_10075,N_10180);
nand U10884 (N_10884,N_10370,N_10009);
or U10885 (N_10885,N_10161,N_9872);
or U10886 (N_10886,N_10176,N_9883);
or U10887 (N_10887,N_10339,N_10455);
and U10888 (N_10888,N_10164,N_10106);
nor U10889 (N_10889,N_10171,N_10378);
xor U10890 (N_10890,N_9759,N_10208);
nor U10891 (N_10891,N_9975,N_9961);
nor U10892 (N_10892,N_10371,N_10227);
xor U10893 (N_10893,N_10219,N_10381);
or U10894 (N_10894,N_9790,N_10189);
nor U10895 (N_10895,N_10453,N_10301);
xor U10896 (N_10896,N_10486,N_10191);
xnor U10897 (N_10897,N_9877,N_10396);
nand U10898 (N_10898,N_10406,N_9963);
and U10899 (N_10899,N_10085,N_10029);
xnor U10900 (N_10900,N_10438,N_10014);
and U10901 (N_10901,N_10364,N_10471);
and U10902 (N_10902,N_10194,N_10150);
and U10903 (N_10903,N_9992,N_9839);
nor U10904 (N_10904,N_10422,N_10369);
nand U10905 (N_10905,N_10176,N_9906);
nand U10906 (N_10906,N_9953,N_9856);
nand U10907 (N_10907,N_10237,N_10013);
nor U10908 (N_10908,N_10204,N_9984);
xnor U10909 (N_10909,N_9914,N_10430);
nand U10910 (N_10910,N_10078,N_10329);
and U10911 (N_10911,N_10482,N_10266);
and U10912 (N_10912,N_9890,N_9795);
xor U10913 (N_10913,N_10060,N_10185);
nor U10914 (N_10914,N_10228,N_10315);
nand U10915 (N_10915,N_10165,N_10175);
or U10916 (N_10916,N_10002,N_10404);
xnor U10917 (N_10917,N_9935,N_10252);
xnor U10918 (N_10918,N_9828,N_10283);
nand U10919 (N_10919,N_10082,N_10168);
or U10920 (N_10920,N_10382,N_10437);
or U10921 (N_10921,N_10437,N_9990);
xor U10922 (N_10922,N_9901,N_10233);
nand U10923 (N_10923,N_9845,N_9897);
xnor U10924 (N_10924,N_9972,N_9752);
nor U10925 (N_10925,N_10443,N_10475);
xnor U10926 (N_10926,N_10015,N_10016);
nor U10927 (N_10927,N_10112,N_10020);
nor U10928 (N_10928,N_10360,N_10353);
nand U10929 (N_10929,N_10432,N_9883);
nor U10930 (N_10930,N_10377,N_10204);
nand U10931 (N_10931,N_10029,N_10431);
xnor U10932 (N_10932,N_10042,N_9819);
xor U10933 (N_10933,N_10043,N_10380);
nor U10934 (N_10934,N_9759,N_9896);
or U10935 (N_10935,N_9930,N_10087);
nand U10936 (N_10936,N_10062,N_9904);
nor U10937 (N_10937,N_10078,N_9908);
and U10938 (N_10938,N_10429,N_10189);
and U10939 (N_10939,N_10365,N_9947);
nand U10940 (N_10940,N_9873,N_10440);
nor U10941 (N_10941,N_9798,N_10192);
and U10942 (N_10942,N_10039,N_10338);
nand U10943 (N_10943,N_9855,N_9815);
or U10944 (N_10944,N_10414,N_9907);
or U10945 (N_10945,N_9942,N_9964);
nand U10946 (N_10946,N_10388,N_10486);
nand U10947 (N_10947,N_10470,N_10458);
nand U10948 (N_10948,N_10080,N_10071);
nand U10949 (N_10949,N_10427,N_10164);
or U10950 (N_10950,N_10303,N_10223);
or U10951 (N_10951,N_9774,N_9915);
nand U10952 (N_10952,N_9935,N_10184);
or U10953 (N_10953,N_10355,N_9982);
or U10954 (N_10954,N_10391,N_9819);
nand U10955 (N_10955,N_10191,N_10335);
nand U10956 (N_10956,N_10254,N_10156);
nor U10957 (N_10957,N_10326,N_10271);
nor U10958 (N_10958,N_10360,N_9863);
or U10959 (N_10959,N_9831,N_10331);
nand U10960 (N_10960,N_10242,N_9837);
or U10961 (N_10961,N_9885,N_10463);
and U10962 (N_10962,N_10218,N_10325);
nor U10963 (N_10963,N_10403,N_10056);
or U10964 (N_10964,N_10278,N_10217);
nand U10965 (N_10965,N_9852,N_10340);
nand U10966 (N_10966,N_9854,N_9959);
and U10967 (N_10967,N_10438,N_10328);
or U10968 (N_10968,N_9899,N_10201);
nand U10969 (N_10969,N_9863,N_10019);
nand U10970 (N_10970,N_10400,N_10218);
nor U10971 (N_10971,N_10111,N_9998);
and U10972 (N_10972,N_9961,N_9884);
and U10973 (N_10973,N_10401,N_10415);
xor U10974 (N_10974,N_10242,N_9782);
and U10975 (N_10975,N_10120,N_10407);
or U10976 (N_10976,N_10381,N_10014);
nand U10977 (N_10977,N_10392,N_10352);
and U10978 (N_10978,N_10157,N_10411);
xnor U10979 (N_10979,N_9987,N_9838);
nor U10980 (N_10980,N_10116,N_9874);
xnor U10981 (N_10981,N_9827,N_10224);
nand U10982 (N_10982,N_10276,N_10320);
or U10983 (N_10983,N_10489,N_9810);
nand U10984 (N_10984,N_10189,N_10356);
nor U10985 (N_10985,N_10147,N_9911);
nor U10986 (N_10986,N_9751,N_10469);
or U10987 (N_10987,N_10004,N_9854);
nand U10988 (N_10988,N_9855,N_10484);
or U10989 (N_10989,N_10336,N_9985);
and U10990 (N_10990,N_10347,N_10289);
xnor U10991 (N_10991,N_9767,N_9759);
and U10992 (N_10992,N_9841,N_10165);
xnor U10993 (N_10993,N_10398,N_10081);
or U10994 (N_10994,N_9898,N_10147);
and U10995 (N_10995,N_10350,N_9856);
nor U10996 (N_10996,N_10346,N_10047);
nor U10997 (N_10997,N_10409,N_9833);
and U10998 (N_10998,N_9972,N_9884);
nand U10999 (N_10999,N_10233,N_9976);
nor U11000 (N_11000,N_10181,N_10022);
and U11001 (N_11001,N_9852,N_9888);
nand U11002 (N_11002,N_10212,N_10147);
nand U11003 (N_11003,N_10397,N_9998);
and U11004 (N_11004,N_10297,N_10362);
nor U11005 (N_11005,N_9877,N_10349);
nand U11006 (N_11006,N_10482,N_10465);
nand U11007 (N_11007,N_9811,N_10176);
and U11008 (N_11008,N_9814,N_10298);
or U11009 (N_11009,N_9793,N_10180);
xnor U11010 (N_11010,N_9972,N_10319);
and U11011 (N_11011,N_10403,N_9802);
nand U11012 (N_11012,N_10431,N_10078);
nand U11013 (N_11013,N_9878,N_9792);
xor U11014 (N_11014,N_10401,N_9766);
nand U11015 (N_11015,N_10411,N_10132);
or U11016 (N_11016,N_10135,N_9781);
or U11017 (N_11017,N_9876,N_10341);
and U11018 (N_11018,N_9878,N_10249);
and U11019 (N_11019,N_10390,N_10054);
or U11020 (N_11020,N_9761,N_10431);
nor U11021 (N_11021,N_9920,N_10068);
nand U11022 (N_11022,N_10442,N_10405);
or U11023 (N_11023,N_9864,N_10461);
and U11024 (N_11024,N_10436,N_10139);
and U11025 (N_11025,N_10174,N_10304);
or U11026 (N_11026,N_9858,N_10242);
and U11027 (N_11027,N_10158,N_10120);
xnor U11028 (N_11028,N_10184,N_9772);
nor U11029 (N_11029,N_10108,N_10356);
xnor U11030 (N_11030,N_9835,N_9801);
and U11031 (N_11031,N_10153,N_10437);
and U11032 (N_11032,N_10258,N_10092);
and U11033 (N_11033,N_9781,N_10388);
xor U11034 (N_11034,N_9875,N_9956);
nand U11035 (N_11035,N_9894,N_9884);
or U11036 (N_11036,N_10121,N_10170);
xor U11037 (N_11037,N_10257,N_9886);
or U11038 (N_11038,N_9821,N_9893);
and U11039 (N_11039,N_10039,N_9836);
nand U11040 (N_11040,N_9911,N_9835);
xnor U11041 (N_11041,N_10138,N_10390);
and U11042 (N_11042,N_9923,N_10407);
xnor U11043 (N_11043,N_10177,N_9930);
nand U11044 (N_11044,N_9765,N_10259);
xnor U11045 (N_11045,N_10026,N_10432);
and U11046 (N_11046,N_10028,N_10460);
nand U11047 (N_11047,N_10175,N_9865);
nor U11048 (N_11048,N_9835,N_10457);
nand U11049 (N_11049,N_9917,N_10449);
xnor U11050 (N_11050,N_10365,N_10438);
and U11051 (N_11051,N_9785,N_9980);
nor U11052 (N_11052,N_10074,N_10143);
or U11053 (N_11053,N_10144,N_10321);
or U11054 (N_11054,N_9955,N_10338);
nand U11055 (N_11055,N_10146,N_9762);
or U11056 (N_11056,N_10201,N_10324);
or U11057 (N_11057,N_10486,N_10473);
nand U11058 (N_11058,N_9750,N_9924);
nand U11059 (N_11059,N_10297,N_10498);
nand U11060 (N_11060,N_10403,N_10128);
nand U11061 (N_11061,N_10477,N_10304);
nor U11062 (N_11062,N_10396,N_10210);
or U11063 (N_11063,N_10084,N_9790);
nand U11064 (N_11064,N_10244,N_9763);
xor U11065 (N_11065,N_10095,N_10060);
and U11066 (N_11066,N_10432,N_9881);
and U11067 (N_11067,N_9826,N_10111);
nand U11068 (N_11068,N_9820,N_10477);
nor U11069 (N_11069,N_9916,N_10250);
and U11070 (N_11070,N_10102,N_9875);
nor U11071 (N_11071,N_10304,N_9997);
nor U11072 (N_11072,N_10442,N_9787);
and U11073 (N_11073,N_10153,N_10033);
and U11074 (N_11074,N_9867,N_10249);
nor U11075 (N_11075,N_10184,N_10298);
xor U11076 (N_11076,N_9963,N_10083);
xor U11077 (N_11077,N_10433,N_10326);
nor U11078 (N_11078,N_9823,N_10122);
or U11079 (N_11079,N_10183,N_9786);
or U11080 (N_11080,N_10494,N_10465);
nand U11081 (N_11081,N_9791,N_10270);
xor U11082 (N_11082,N_9767,N_10329);
xor U11083 (N_11083,N_9834,N_10436);
and U11084 (N_11084,N_10184,N_10463);
and U11085 (N_11085,N_9940,N_10463);
xor U11086 (N_11086,N_10436,N_10021);
nand U11087 (N_11087,N_10416,N_10054);
xnor U11088 (N_11088,N_9794,N_10033);
xnor U11089 (N_11089,N_10332,N_9860);
or U11090 (N_11090,N_10217,N_10311);
nor U11091 (N_11091,N_10055,N_10268);
and U11092 (N_11092,N_10171,N_10168);
nand U11093 (N_11093,N_9844,N_10275);
xor U11094 (N_11094,N_10007,N_9988);
or U11095 (N_11095,N_10233,N_9856);
and U11096 (N_11096,N_10045,N_10018);
or U11097 (N_11097,N_10049,N_10295);
xnor U11098 (N_11098,N_10164,N_10197);
or U11099 (N_11099,N_9847,N_10142);
nand U11100 (N_11100,N_10246,N_10200);
xnor U11101 (N_11101,N_10110,N_9902);
and U11102 (N_11102,N_9951,N_9899);
or U11103 (N_11103,N_10373,N_10199);
xor U11104 (N_11104,N_10348,N_10149);
or U11105 (N_11105,N_9944,N_10189);
or U11106 (N_11106,N_10338,N_10106);
and U11107 (N_11107,N_10478,N_10066);
nor U11108 (N_11108,N_10156,N_10433);
nand U11109 (N_11109,N_9881,N_9936);
xnor U11110 (N_11110,N_10386,N_10275);
xor U11111 (N_11111,N_10058,N_10026);
nand U11112 (N_11112,N_9861,N_9896);
and U11113 (N_11113,N_9850,N_10309);
xnor U11114 (N_11114,N_10011,N_9936);
and U11115 (N_11115,N_9950,N_10099);
nor U11116 (N_11116,N_10189,N_10377);
nand U11117 (N_11117,N_9928,N_9794);
nand U11118 (N_11118,N_10196,N_10265);
xnor U11119 (N_11119,N_10087,N_10030);
nand U11120 (N_11120,N_9848,N_9881);
xor U11121 (N_11121,N_10349,N_10431);
or U11122 (N_11122,N_10229,N_9988);
or U11123 (N_11123,N_10350,N_10258);
nand U11124 (N_11124,N_9916,N_10155);
xnor U11125 (N_11125,N_10088,N_10137);
or U11126 (N_11126,N_10345,N_10157);
nor U11127 (N_11127,N_10406,N_10208);
and U11128 (N_11128,N_9793,N_10209);
or U11129 (N_11129,N_10456,N_9756);
nand U11130 (N_11130,N_10133,N_9974);
xor U11131 (N_11131,N_9805,N_10034);
and U11132 (N_11132,N_10293,N_10067);
nand U11133 (N_11133,N_9768,N_10022);
xnor U11134 (N_11134,N_9824,N_9793);
nor U11135 (N_11135,N_9753,N_10196);
and U11136 (N_11136,N_10255,N_9893);
nand U11137 (N_11137,N_9874,N_10270);
nor U11138 (N_11138,N_9995,N_9761);
xnor U11139 (N_11139,N_10287,N_9777);
nor U11140 (N_11140,N_10232,N_10326);
nor U11141 (N_11141,N_9988,N_9976);
xnor U11142 (N_11142,N_10493,N_10138);
nand U11143 (N_11143,N_10238,N_9983);
nand U11144 (N_11144,N_10246,N_10259);
xor U11145 (N_11145,N_10288,N_10015);
and U11146 (N_11146,N_10235,N_9929);
and U11147 (N_11147,N_9769,N_10471);
xnor U11148 (N_11148,N_9993,N_10286);
nor U11149 (N_11149,N_9832,N_10364);
or U11150 (N_11150,N_10168,N_10159);
nor U11151 (N_11151,N_10375,N_10334);
nor U11152 (N_11152,N_10159,N_9836);
xnor U11153 (N_11153,N_10170,N_10101);
nor U11154 (N_11154,N_10264,N_10159);
and U11155 (N_11155,N_9892,N_10263);
or U11156 (N_11156,N_9757,N_10024);
xnor U11157 (N_11157,N_9934,N_10093);
or U11158 (N_11158,N_10247,N_9992);
xor U11159 (N_11159,N_10475,N_9935);
and U11160 (N_11160,N_10319,N_9813);
and U11161 (N_11161,N_10074,N_10126);
nand U11162 (N_11162,N_10363,N_10285);
xor U11163 (N_11163,N_10375,N_10167);
nor U11164 (N_11164,N_10330,N_10321);
or U11165 (N_11165,N_9875,N_10182);
nor U11166 (N_11166,N_10331,N_9971);
nor U11167 (N_11167,N_10018,N_10484);
or U11168 (N_11168,N_9907,N_10478);
and U11169 (N_11169,N_10003,N_9794);
or U11170 (N_11170,N_9933,N_10236);
or U11171 (N_11171,N_9968,N_9813);
and U11172 (N_11172,N_10321,N_10378);
nor U11173 (N_11173,N_10445,N_10132);
and U11174 (N_11174,N_10065,N_9822);
or U11175 (N_11175,N_10264,N_9845);
nand U11176 (N_11176,N_10320,N_10438);
nor U11177 (N_11177,N_10289,N_10259);
nand U11178 (N_11178,N_10387,N_10285);
and U11179 (N_11179,N_9777,N_10095);
nor U11180 (N_11180,N_9887,N_10324);
xor U11181 (N_11181,N_9956,N_10471);
and U11182 (N_11182,N_10332,N_10047);
nand U11183 (N_11183,N_9984,N_10172);
nand U11184 (N_11184,N_10304,N_10333);
or U11185 (N_11185,N_10339,N_10347);
xnor U11186 (N_11186,N_10171,N_9833);
nand U11187 (N_11187,N_9969,N_10386);
xor U11188 (N_11188,N_9753,N_9860);
or U11189 (N_11189,N_10060,N_9777);
nor U11190 (N_11190,N_9931,N_10216);
nor U11191 (N_11191,N_10132,N_10249);
and U11192 (N_11192,N_9870,N_10121);
nor U11193 (N_11193,N_10052,N_10495);
xnor U11194 (N_11194,N_9770,N_10282);
xor U11195 (N_11195,N_10243,N_9794);
and U11196 (N_11196,N_10046,N_10409);
or U11197 (N_11197,N_10210,N_10031);
nor U11198 (N_11198,N_9950,N_10054);
nor U11199 (N_11199,N_10217,N_10094);
nor U11200 (N_11200,N_10213,N_10318);
or U11201 (N_11201,N_10259,N_10245);
and U11202 (N_11202,N_9846,N_10400);
or U11203 (N_11203,N_10341,N_10396);
and U11204 (N_11204,N_10465,N_9940);
nor U11205 (N_11205,N_9787,N_10193);
nor U11206 (N_11206,N_10499,N_9760);
or U11207 (N_11207,N_9842,N_9925);
nor U11208 (N_11208,N_10453,N_10428);
xnor U11209 (N_11209,N_10353,N_10392);
or U11210 (N_11210,N_10105,N_10357);
or U11211 (N_11211,N_10424,N_10005);
nor U11212 (N_11212,N_10073,N_10259);
nor U11213 (N_11213,N_10485,N_9888);
nand U11214 (N_11214,N_9957,N_10011);
and U11215 (N_11215,N_9753,N_9928);
nor U11216 (N_11216,N_9920,N_10407);
or U11217 (N_11217,N_10292,N_9985);
or U11218 (N_11218,N_9756,N_9953);
nor U11219 (N_11219,N_9788,N_9821);
nand U11220 (N_11220,N_10238,N_10294);
nand U11221 (N_11221,N_9926,N_9997);
and U11222 (N_11222,N_10406,N_10068);
nor U11223 (N_11223,N_10465,N_10469);
and U11224 (N_11224,N_10129,N_9904);
xnor U11225 (N_11225,N_9908,N_10497);
and U11226 (N_11226,N_10290,N_10187);
xnor U11227 (N_11227,N_10130,N_10423);
nand U11228 (N_11228,N_10019,N_9945);
or U11229 (N_11229,N_9770,N_9994);
nor U11230 (N_11230,N_9763,N_9821);
xnor U11231 (N_11231,N_9864,N_9861);
xor U11232 (N_11232,N_10421,N_9845);
xnor U11233 (N_11233,N_10039,N_10017);
nor U11234 (N_11234,N_10360,N_10405);
or U11235 (N_11235,N_9891,N_10432);
nand U11236 (N_11236,N_9861,N_10088);
nor U11237 (N_11237,N_10317,N_9917);
or U11238 (N_11238,N_9998,N_10242);
nand U11239 (N_11239,N_10074,N_9858);
or U11240 (N_11240,N_9755,N_10188);
xnor U11241 (N_11241,N_9967,N_9938);
nor U11242 (N_11242,N_9934,N_10180);
or U11243 (N_11243,N_10206,N_9917);
nand U11244 (N_11244,N_10367,N_9825);
and U11245 (N_11245,N_10140,N_10240);
nand U11246 (N_11246,N_10232,N_9934);
xnor U11247 (N_11247,N_10232,N_10442);
xnor U11248 (N_11248,N_10419,N_10324);
xnor U11249 (N_11249,N_9892,N_10432);
or U11250 (N_11250,N_11042,N_11071);
nor U11251 (N_11251,N_10892,N_10591);
or U11252 (N_11252,N_10769,N_11006);
and U11253 (N_11253,N_10571,N_11084);
nor U11254 (N_11254,N_10614,N_11064);
xnor U11255 (N_11255,N_10874,N_10573);
or U11256 (N_11256,N_10736,N_10574);
nor U11257 (N_11257,N_10524,N_10785);
or U11258 (N_11258,N_11146,N_10692);
or U11259 (N_11259,N_10621,N_10841);
nor U11260 (N_11260,N_10526,N_10963);
nor U11261 (N_11261,N_11182,N_10625);
and U11262 (N_11262,N_10786,N_10965);
nand U11263 (N_11263,N_10779,N_10729);
and U11264 (N_11264,N_10952,N_11175);
xnor U11265 (N_11265,N_10525,N_10985);
nand U11266 (N_11266,N_10734,N_10822);
xor U11267 (N_11267,N_10577,N_11185);
or U11268 (N_11268,N_11072,N_10813);
and U11269 (N_11269,N_11007,N_10540);
or U11270 (N_11270,N_11050,N_10996);
or U11271 (N_11271,N_10661,N_11133);
and U11272 (N_11272,N_10857,N_10776);
nor U11273 (N_11273,N_10935,N_10914);
and U11274 (N_11274,N_10878,N_10703);
nand U11275 (N_11275,N_10659,N_11149);
xor U11276 (N_11276,N_10522,N_10881);
or U11277 (N_11277,N_10856,N_10840);
or U11278 (N_11278,N_10508,N_10981);
or U11279 (N_11279,N_10553,N_10739);
and U11280 (N_11280,N_11016,N_10992);
nor U11281 (N_11281,N_11115,N_10842);
xor U11282 (N_11282,N_10554,N_10937);
nor U11283 (N_11283,N_10720,N_10768);
nand U11284 (N_11284,N_10596,N_10559);
or U11285 (N_11285,N_11210,N_11138);
or U11286 (N_11286,N_10609,N_10607);
xnor U11287 (N_11287,N_11188,N_10610);
or U11288 (N_11288,N_10599,N_10814);
or U11289 (N_11289,N_11011,N_11035);
xor U11290 (N_11290,N_10651,N_10950);
xnor U11291 (N_11291,N_10957,N_10564);
and U11292 (N_11292,N_10618,N_10649);
nor U11293 (N_11293,N_10701,N_10948);
nor U11294 (N_11294,N_10517,N_10839);
or U11295 (N_11295,N_11154,N_10859);
and U11296 (N_11296,N_11039,N_11102);
or U11297 (N_11297,N_10853,N_10897);
and U11298 (N_11298,N_10527,N_11067);
nor U11299 (N_11299,N_10636,N_10654);
or U11300 (N_11300,N_11082,N_10514);
nand U11301 (N_11301,N_11107,N_10560);
nand U11302 (N_11302,N_10794,N_11128);
nor U11303 (N_11303,N_10602,N_10835);
nand U11304 (N_11304,N_10656,N_10975);
nor U11305 (N_11305,N_10576,N_11065);
nand U11306 (N_11306,N_10558,N_11002);
nor U11307 (N_11307,N_10593,N_11096);
xnor U11308 (N_11308,N_10706,N_10851);
nor U11309 (N_11309,N_10657,N_10807);
and U11310 (N_11310,N_11017,N_10547);
nor U11311 (N_11311,N_10708,N_11069);
or U11312 (N_11312,N_11018,N_10848);
nor U11313 (N_11313,N_10579,N_11235);
and U11314 (N_11314,N_10766,N_11086);
and U11315 (N_11315,N_10863,N_10556);
nor U11316 (N_11316,N_11236,N_10974);
and U11317 (N_11317,N_11213,N_10601);
and U11318 (N_11318,N_11159,N_10995);
or U11319 (N_11319,N_10740,N_10541);
xor U11320 (N_11320,N_10660,N_10873);
nand U11321 (N_11321,N_10843,N_10650);
xor U11322 (N_11322,N_10764,N_10689);
nand U11323 (N_11323,N_10888,N_10664);
or U11324 (N_11324,N_10868,N_11156);
xor U11325 (N_11325,N_11066,N_10917);
nor U11326 (N_11326,N_10889,N_10698);
nand U11327 (N_11327,N_11121,N_11075);
nor U11328 (N_11328,N_10772,N_11222);
nand U11329 (N_11329,N_11049,N_10972);
and U11330 (N_11330,N_10630,N_11073);
nor U11331 (N_11331,N_10683,N_11201);
nand U11332 (N_11332,N_10982,N_11012);
xnor U11333 (N_11333,N_10686,N_11215);
or U11334 (N_11334,N_11232,N_10635);
or U11335 (N_11335,N_10936,N_10905);
xnor U11336 (N_11336,N_10767,N_10548);
nor U11337 (N_11337,N_11170,N_10770);
nor U11338 (N_11338,N_11190,N_11151);
xnor U11339 (N_11339,N_10631,N_10969);
or U11340 (N_11340,N_10731,N_10836);
nand U11341 (N_11341,N_10902,N_10688);
xnor U11342 (N_11342,N_10855,N_11090);
nand U11343 (N_11343,N_10871,N_10988);
nor U11344 (N_11344,N_10928,N_11217);
and U11345 (N_11345,N_10805,N_11059);
and U11346 (N_11346,N_10586,N_10940);
and U11347 (N_11347,N_10726,N_10529);
nand U11348 (N_11348,N_11010,N_10763);
or U11349 (N_11349,N_10968,N_10699);
and U11350 (N_11350,N_10815,N_11013);
xor U11351 (N_11351,N_10994,N_10745);
and U11352 (N_11352,N_10641,N_10854);
nand U11353 (N_11353,N_11135,N_11108);
nand U11354 (N_11354,N_10542,N_10959);
nand U11355 (N_11355,N_10738,N_10771);
and U11356 (N_11356,N_11105,N_10746);
or U11357 (N_11357,N_10580,N_11085);
nand U11358 (N_11358,N_10678,N_10569);
or U11359 (N_11359,N_10816,N_10960);
or U11360 (N_11360,N_10826,N_11112);
nor U11361 (N_11361,N_11131,N_10642);
xor U11362 (N_11362,N_10752,N_11089);
xnor U11363 (N_11363,N_10903,N_10949);
nor U11364 (N_11364,N_10684,N_10587);
nand U11365 (N_11365,N_10755,N_10804);
nor U11366 (N_11366,N_10709,N_10846);
nand U11367 (N_11367,N_11098,N_10510);
and U11368 (N_11368,N_11220,N_11172);
nand U11369 (N_11369,N_10674,N_11046);
xor U11370 (N_11370,N_11168,N_10637);
nand U11371 (N_11371,N_11130,N_10557);
nand U11372 (N_11372,N_10906,N_11103);
xor U11373 (N_11373,N_10912,N_10711);
xor U11374 (N_11374,N_10552,N_11228);
and U11375 (N_11375,N_10900,N_10750);
and U11376 (N_11376,N_10612,N_10980);
nor U11377 (N_11377,N_10507,N_10796);
nor U11378 (N_11378,N_10680,N_10644);
or U11379 (N_11379,N_10971,N_11001);
nand U11380 (N_11380,N_10502,N_10943);
xnor U11381 (N_11381,N_10611,N_11126);
xor U11382 (N_11382,N_10531,N_10882);
or U11383 (N_11383,N_11211,N_11184);
xnor U11384 (N_11384,N_10978,N_10789);
xor U11385 (N_11385,N_10597,N_10845);
xnor U11386 (N_11386,N_10781,N_10691);
xnor U11387 (N_11387,N_10964,N_10802);
xor U11388 (N_11388,N_10954,N_11180);
or U11389 (N_11389,N_10808,N_11056);
nand U11390 (N_11390,N_10872,N_11003);
nand U11391 (N_11391,N_11015,N_10676);
nor U11392 (N_11392,N_11019,N_11063);
xor U11393 (N_11393,N_11139,N_10511);
xnor U11394 (N_11394,N_11053,N_11174);
or U11395 (N_11395,N_10667,N_11218);
nor U11396 (N_11396,N_10737,N_10753);
or U11397 (N_11397,N_11078,N_10951);
nand U11398 (N_11398,N_11093,N_10723);
and U11399 (N_11399,N_10617,N_10655);
xor U11400 (N_11400,N_11216,N_10710);
or U11401 (N_11401,N_10918,N_10504);
nor U11402 (N_11402,N_10604,N_11051);
or U11403 (N_11403,N_10645,N_10890);
nand U11404 (N_11404,N_11062,N_10697);
and U11405 (N_11405,N_10622,N_10687);
or U11406 (N_11406,N_10877,N_11153);
or U11407 (N_11407,N_10879,N_10575);
nor U11408 (N_11408,N_10911,N_10880);
or U11409 (N_11409,N_11152,N_10926);
or U11410 (N_11410,N_10800,N_10942);
or U11411 (N_11411,N_10898,N_10665);
nand U11412 (N_11412,N_10501,N_10748);
nand U11413 (N_11413,N_10515,N_10567);
nor U11414 (N_11414,N_10714,N_10572);
nor U11415 (N_11415,N_11036,N_11113);
nand U11416 (N_11416,N_10530,N_11041);
xnor U11417 (N_11417,N_10545,N_10707);
or U11418 (N_11418,N_11045,N_10788);
and U11419 (N_11419,N_11111,N_10973);
xnor U11420 (N_11420,N_11021,N_10820);
nor U11421 (N_11421,N_11148,N_11161);
or U11422 (N_11422,N_11127,N_11114);
xnor U11423 (N_11423,N_10727,N_11000);
or U11424 (N_11424,N_10549,N_10647);
or U11425 (N_11425,N_11077,N_10639);
nor U11426 (N_11426,N_11150,N_10817);
nor U11427 (N_11427,N_10931,N_10941);
xnor U11428 (N_11428,N_10732,N_11141);
or U11429 (N_11429,N_11123,N_10758);
or U11430 (N_11430,N_10884,N_10741);
nand U11431 (N_11431,N_11186,N_10901);
and U11432 (N_11432,N_11239,N_11212);
nor U11433 (N_11433,N_11054,N_10894);
xnor U11434 (N_11434,N_10718,N_10916);
and U11435 (N_11435,N_10929,N_10893);
nor U11436 (N_11436,N_10668,N_10538);
nand U11437 (N_11437,N_11116,N_10934);
or U11438 (N_11438,N_10761,N_10619);
xor U11439 (N_11439,N_10725,N_10722);
nor U11440 (N_11440,N_10953,N_10512);
or U11441 (N_11441,N_10838,N_10589);
or U11442 (N_11442,N_11166,N_10624);
xor U11443 (N_11443,N_10534,N_11118);
nand U11444 (N_11444,N_10883,N_10966);
and U11445 (N_11445,N_10885,N_11206);
and U11446 (N_11446,N_11004,N_10896);
nand U11447 (N_11447,N_11140,N_11047);
nor U11448 (N_11448,N_10719,N_11244);
or U11449 (N_11449,N_11189,N_10773);
or U11450 (N_11450,N_11100,N_11183);
nand U11451 (N_11451,N_10724,N_10673);
nand U11452 (N_11452,N_11162,N_10730);
xor U11453 (N_11453,N_11029,N_10812);
and U11454 (N_11454,N_10821,N_10628);
and U11455 (N_11455,N_11167,N_10595);
or U11456 (N_11456,N_10696,N_10690);
nand U11457 (N_11457,N_11227,N_10682);
nor U11458 (N_11458,N_10565,N_10875);
or U11459 (N_11459,N_11097,N_10747);
and U11460 (N_11460,N_10584,N_11122);
and U11461 (N_11461,N_10946,N_11198);
or U11462 (N_11462,N_11060,N_11230);
xnor U11463 (N_11463,N_10955,N_11038);
or U11464 (N_11464,N_11094,N_11243);
nor U11465 (N_11465,N_11238,N_10915);
and U11466 (N_11466,N_10904,N_10694);
nand U11467 (N_11467,N_11080,N_10551);
nand U11468 (N_11468,N_10503,N_10819);
nand U11469 (N_11469,N_11110,N_11033);
nand U11470 (N_11470,N_11176,N_10570);
nand U11471 (N_11471,N_10793,N_10823);
nor U11472 (N_11472,N_10986,N_10742);
xor U11473 (N_11473,N_10967,N_11024);
or U11474 (N_11474,N_10924,N_10518);
xor U11475 (N_11475,N_11032,N_10891);
nor U11476 (N_11476,N_10716,N_11240);
or U11477 (N_11477,N_11209,N_10864);
nand U11478 (N_11478,N_10590,N_11109);
or U11479 (N_11479,N_10733,N_10827);
and U11480 (N_11480,N_10913,N_10550);
nand U11481 (N_11481,N_10536,N_10632);
nor U11482 (N_11482,N_10832,N_11155);
and U11483 (N_11483,N_10834,N_10850);
or U11484 (N_11484,N_11023,N_10585);
nor U11485 (N_11485,N_11169,N_11225);
or U11486 (N_11486,N_11247,N_11231);
nor U11487 (N_11487,N_11224,N_10970);
or U11488 (N_11488,N_10977,N_11197);
or U11489 (N_11489,N_11202,N_10962);
nand U11490 (N_11490,N_11214,N_11160);
nor U11491 (N_11491,N_10833,N_10790);
and U11492 (N_11492,N_10728,N_10930);
or U11493 (N_11493,N_10824,N_11068);
nor U11494 (N_11494,N_10782,N_11020);
nand U11495 (N_11495,N_10615,N_11091);
and U11496 (N_11496,N_10643,N_10847);
xor U11497 (N_11497,N_11074,N_10700);
xnor U11498 (N_11498,N_11163,N_10671);
xnor U11499 (N_11499,N_10806,N_10945);
nor U11500 (N_11500,N_10870,N_11005);
nand U11501 (N_11501,N_10670,N_10582);
xnor U11502 (N_11502,N_10629,N_10958);
nand U11503 (N_11503,N_10860,N_10606);
nand U11504 (N_11504,N_10563,N_10895);
nand U11505 (N_11505,N_11196,N_11226);
nand U11506 (N_11506,N_10681,N_10605);
nand U11507 (N_11507,N_11014,N_10594);
and U11508 (N_11508,N_10837,N_11079);
nand U11509 (N_11509,N_10997,N_11052);
nand U11510 (N_11510,N_11177,N_11192);
xnor U11511 (N_11511,N_10780,N_11028);
nand U11512 (N_11512,N_10715,N_10533);
xor U11513 (N_11513,N_10712,N_11194);
and U11514 (N_11514,N_10987,N_10791);
or U11515 (N_11515,N_11147,N_10909);
or U11516 (N_11516,N_11233,N_10623);
nand U11517 (N_11517,N_10662,N_11237);
xor U11518 (N_11518,N_11088,N_10634);
or U11519 (N_11519,N_11034,N_10744);
nand U11520 (N_11520,N_10886,N_10505);
nor U11521 (N_11521,N_11125,N_11221);
xor U11522 (N_11522,N_10803,N_10828);
nor U11523 (N_11523,N_10998,N_10713);
nor U11524 (N_11524,N_10798,N_10908);
or U11525 (N_11525,N_10535,N_11219);
xnor U11526 (N_11526,N_11137,N_11101);
xnor U11527 (N_11527,N_10652,N_10638);
and U11528 (N_11528,N_10756,N_11043);
and U11529 (N_11529,N_10976,N_10947);
nand U11530 (N_11530,N_10588,N_11099);
xnor U11531 (N_11531,N_11245,N_10669);
and U11532 (N_11532,N_10562,N_11143);
and U11533 (N_11533,N_10775,N_10869);
or U11534 (N_11534,N_10899,N_11027);
nor U11535 (N_11535,N_11040,N_10944);
nand U11536 (N_11536,N_10993,N_11022);
or U11537 (N_11537,N_11087,N_10513);
nor U11538 (N_11538,N_10537,N_10583);
nand U11539 (N_11539,N_10546,N_10648);
nand U11540 (N_11540,N_11249,N_10633);
and U11541 (N_11541,N_11200,N_10777);
nor U11542 (N_11542,N_10616,N_10925);
or U11543 (N_11543,N_11026,N_10685);
nand U11544 (N_11544,N_11124,N_11142);
or U11545 (N_11545,N_10810,N_11248);
and U11546 (N_11546,N_10760,N_10520);
or U11547 (N_11547,N_10989,N_11187);
nand U11548 (N_11548,N_10543,N_10704);
or U11549 (N_11549,N_11171,N_11165);
xor U11550 (N_11550,N_10910,N_11061);
xor U11551 (N_11551,N_11058,N_11092);
or U11552 (N_11552,N_10825,N_10519);
and U11553 (N_11553,N_11234,N_11246);
and U11554 (N_11554,N_11157,N_10523);
xnor U11555 (N_11555,N_10811,N_10754);
nor U11556 (N_11556,N_10933,N_11076);
xor U11557 (N_11557,N_11048,N_10849);
nor U11558 (N_11558,N_11055,N_10797);
and U11559 (N_11559,N_11030,N_10627);
nor U11560 (N_11560,N_10516,N_11095);
nand U11561 (N_11561,N_10555,N_11205);
nor U11562 (N_11562,N_10561,N_10795);
or U11563 (N_11563,N_10999,N_10867);
or U11564 (N_11564,N_10608,N_11193);
xor U11565 (N_11565,N_11181,N_10663);
and U11566 (N_11566,N_10932,N_11117);
nor U11567 (N_11567,N_10675,N_11129);
or U11568 (N_11568,N_10695,N_10830);
and U11569 (N_11569,N_10865,N_11081);
xnor U11570 (N_11570,N_10749,N_10844);
or U11571 (N_11571,N_11009,N_10658);
or U11572 (N_11572,N_10774,N_10927);
xor U11573 (N_11573,N_11145,N_10979);
or U11574 (N_11574,N_10938,N_11242);
xnor U11575 (N_11575,N_10693,N_10923);
and U11576 (N_11576,N_10702,N_10528);
or U11577 (N_11577,N_11191,N_10818);
nor U11578 (N_11578,N_10876,N_10809);
and U11579 (N_11579,N_10919,N_10603);
xor U11580 (N_11580,N_11179,N_11120);
xnor U11581 (N_11581,N_10509,N_10646);
xor U11582 (N_11582,N_10920,N_10500);
xor U11583 (N_11583,N_10990,N_10626);
xnor U11584 (N_11584,N_10792,N_10672);
xor U11585 (N_11585,N_11207,N_11203);
or U11586 (N_11586,N_10581,N_10598);
xnor U11587 (N_11587,N_10751,N_10620);
nand U11588 (N_11588,N_11199,N_10566);
nor U11589 (N_11589,N_11158,N_10759);
nor U11590 (N_11590,N_10852,N_11208);
and U11591 (N_11591,N_10984,N_10705);
nor U11592 (N_11592,N_10544,N_11223);
nand U11593 (N_11593,N_10757,N_11031);
nand U11594 (N_11594,N_10939,N_10862);
xnor U11595 (N_11595,N_11044,N_11241);
or U11596 (N_11596,N_11204,N_10778);
or U11597 (N_11597,N_11057,N_10743);
nor U11598 (N_11598,N_10539,N_10653);
xor U11599 (N_11599,N_10866,N_11070);
and U11600 (N_11600,N_10991,N_11119);
nor U11601 (N_11601,N_11104,N_10568);
nor U11602 (N_11602,N_11008,N_10640);
or U11603 (N_11603,N_10532,N_10666);
and U11604 (N_11604,N_10961,N_10956);
nand U11605 (N_11605,N_10717,N_11144);
nand U11606 (N_11606,N_10521,N_10784);
xnor U11607 (N_11607,N_10921,N_10922);
nor U11608 (N_11608,N_10578,N_11134);
and U11609 (N_11609,N_10679,N_10765);
nor U11610 (N_11610,N_11132,N_10861);
nand U11611 (N_11611,N_11173,N_10677);
or U11612 (N_11612,N_10506,N_10735);
or U11613 (N_11613,N_10799,N_10787);
or U11614 (N_11614,N_10762,N_11178);
and U11615 (N_11615,N_10600,N_10613);
xnor U11616 (N_11616,N_10801,N_11106);
xor U11617 (N_11617,N_11229,N_11195);
or U11618 (N_11618,N_10858,N_11025);
and U11619 (N_11619,N_11164,N_11136);
and U11620 (N_11620,N_11037,N_10829);
and U11621 (N_11621,N_10907,N_10831);
xor U11622 (N_11622,N_10592,N_11083);
and U11623 (N_11623,N_10721,N_10887);
or U11624 (N_11624,N_10783,N_10983);
nand U11625 (N_11625,N_11056,N_10968);
nor U11626 (N_11626,N_10832,N_11044);
nor U11627 (N_11627,N_11151,N_10837);
and U11628 (N_11628,N_10780,N_11147);
or U11629 (N_11629,N_11126,N_10799);
or U11630 (N_11630,N_11176,N_10513);
nand U11631 (N_11631,N_10831,N_10674);
or U11632 (N_11632,N_10780,N_11186);
and U11633 (N_11633,N_11010,N_11005);
xnor U11634 (N_11634,N_11229,N_10857);
or U11635 (N_11635,N_10909,N_10992);
and U11636 (N_11636,N_10959,N_10964);
and U11637 (N_11637,N_10913,N_10666);
nand U11638 (N_11638,N_10873,N_10803);
and U11639 (N_11639,N_10619,N_11131);
and U11640 (N_11640,N_10836,N_10711);
nand U11641 (N_11641,N_11211,N_10857);
nor U11642 (N_11642,N_11060,N_11221);
or U11643 (N_11643,N_11137,N_10501);
nand U11644 (N_11644,N_10907,N_10896);
and U11645 (N_11645,N_10776,N_10611);
xnor U11646 (N_11646,N_11028,N_10562);
and U11647 (N_11647,N_10777,N_11109);
or U11648 (N_11648,N_11177,N_10967);
nand U11649 (N_11649,N_10774,N_10868);
and U11650 (N_11650,N_10673,N_10752);
or U11651 (N_11651,N_10730,N_10709);
or U11652 (N_11652,N_10652,N_10989);
nand U11653 (N_11653,N_10648,N_11076);
or U11654 (N_11654,N_11011,N_10991);
or U11655 (N_11655,N_10992,N_10734);
nand U11656 (N_11656,N_10654,N_10578);
nor U11657 (N_11657,N_10526,N_11171);
nand U11658 (N_11658,N_10530,N_10794);
or U11659 (N_11659,N_10959,N_10707);
nand U11660 (N_11660,N_10815,N_10509);
and U11661 (N_11661,N_10841,N_11237);
nor U11662 (N_11662,N_11218,N_10783);
nand U11663 (N_11663,N_10587,N_10574);
nor U11664 (N_11664,N_10971,N_10606);
xnor U11665 (N_11665,N_10901,N_10867);
xor U11666 (N_11666,N_10856,N_11169);
or U11667 (N_11667,N_11102,N_10834);
and U11668 (N_11668,N_10622,N_10564);
xnor U11669 (N_11669,N_10594,N_10576);
xor U11670 (N_11670,N_10576,N_10617);
xor U11671 (N_11671,N_10653,N_11161);
nor U11672 (N_11672,N_11032,N_10765);
or U11673 (N_11673,N_10590,N_10987);
nand U11674 (N_11674,N_10730,N_10938);
nand U11675 (N_11675,N_10614,N_11245);
or U11676 (N_11676,N_10701,N_10821);
nor U11677 (N_11677,N_10502,N_10987);
xnor U11678 (N_11678,N_10635,N_10633);
nand U11679 (N_11679,N_10531,N_11185);
nor U11680 (N_11680,N_10700,N_11142);
nand U11681 (N_11681,N_10675,N_10956);
nand U11682 (N_11682,N_10908,N_11081);
nand U11683 (N_11683,N_11051,N_10706);
xnor U11684 (N_11684,N_10618,N_10600);
nand U11685 (N_11685,N_10610,N_11192);
nand U11686 (N_11686,N_10923,N_10849);
or U11687 (N_11687,N_10721,N_11039);
nor U11688 (N_11688,N_10946,N_10598);
or U11689 (N_11689,N_10530,N_10993);
nand U11690 (N_11690,N_11182,N_11003);
and U11691 (N_11691,N_11036,N_10662);
xor U11692 (N_11692,N_10860,N_10631);
xnor U11693 (N_11693,N_11164,N_11241);
or U11694 (N_11694,N_10793,N_10578);
nor U11695 (N_11695,N_11166,N_10636);
nor U11696 (N_11696,N_10616,N_10519);
or U11697 (N_11697,N_10574,N_10977);
nor U11698 (N_11698,N_10756,N_11171);
or U11699 (N_11699,N_11227,N_10956);
xor U11700 (N_11700,N_11195,N_10639);
nand U11701 (N_11701,N_10948,N_10688);
nand U11702 (N_11702,N_10782,N_11123);
xor U11703 (N_11703,N_10983,N_11093);
xnor U11704 (N_11704,N_10693,N_10699);
and U11705 (N_11705,N_11049,N_11081);
nor U11706 (N_11706,N_10650,N_11096);
or U11707 (N_11707,N_10554,N_10880);
nand U11708 (N_11708,N_10923,N_11042);
or U11709 (N_11709,N_10631,N_10831);
nand U11710 (N_11710,N_10802,N_11067);
or U11711 (N_11711,N_10693,N_11085);
xor U11712 (N_11712,N_11173,N_10618);
nor U11713 (N_11713,N_10583,N_10952);
nand U11714 (N_11714,N_11242,N_10720);
and U11715 (N_11715,N_11130,N_11114);
xor U11716 (N_11716,N_10915,N_10551);
and U11717 (N_11717,N_10655,N_10682);
nand U11718 (N_11718,N_10894,N_10938);
or U11719 (N_11719,N_10996,N_10824);
xor U11720 (N_11720,N_10980,N_10572);
xor U11721 (N_11721,N_10629,N_11145);
nor U11722 (N_11722,N_11088,N_11224);
or U11723 (N_11723,N_10645,N_10509);
and U11724 (N_11724,N_11089,N_11138);
xnor U11725 (N_11725,N_11060,N_11143);
or U11726 (N_11726,N_11147,N_11011);
or U11727 (N_11727,N_10629,N_10735);
nor U11728 (N_11728,N_11108,N_11153);
nand U11729 (N_11729,N_10917,N_11178);
or U11730 (N_11730,N_10736,N_10630);
nand U11731 (N_11731,N_11193,N_10764);
xnor U11732 (N_11732,N_10573,N_10791);
nor U11733 (N_11733,N_10979,N_10834);
or U11734 (N_11734,N_10695,N_10704);
nor U11735 (N_11735,N_11247,N_10668);
nand U11736 (N_11736,N_11162,N_10575);
nand U11737 (N_11737,N_10707,N_10634);
and U11738 (N_11738,N_11123,N_11008);
or U11739 (N_11739,N_10918,N_10658);
nor U11740 (N_11740,N_10551,N_10677);
nand U11741 (N_11741,N_10774,N_10557);
nor U11742 (N_11742,N_10515,N_11020);
and U11743 (N_11743,N_11196,N_10740);
nor U11744 (N_11744,N_10800,N_10575);
xor U11745 (N_11745,N_10577,N_10696);
xor U11746 (N_11746,N_10829,N_10857);
or U11747 (N_11747,N_11207,N_11056);
xor U11748 (N_11748,N_10974,N_10531);
nor U11749 (N_11749,N_11008,N_10907);
xor U11750 (N_11750,N_10710,N_10558);
or U11751 (N_11751,N_10658,N_11155);
nand U11752 (N_11752,N_11068,N_10988);
nand U11753 (N_11753,N_11182,N_10521);
and U11754 (N_11754,N_10558,N_10626);
nor U11755 (N_11755,N_10840,N_10862);
and U11756 (N_11756,N_10740,N_10847);
and U11757 (N_11757,N_10790,N_11142);
and U11758 (N_11758,N_10561,N_10616);
xor U11759 (N_11759,N_10671,N_11183);
and U11760 (N_11760,N_10593,N_11156);
xor U11761 (N_11761,N_11161,N_10985);
xnor U11762 (N_11762,N_10978,N_10616);
xnor U11763 (N_11763,N_11197,N_10594);
xor U11764 (N_11764,N_10903,N_11038);
nor U11765 (N_11765,N_11210,N_10751);
or U11766 (N_11766,N_11209,N_11087);
nand U11767 (N_11767,N_10698,N_11092);
and U11768 (N_11768,N_11180,N_10617);
or U11769 (N_11769,N_11129,N_10785);
or U11770 (N_11770,N_10883,N_10505);
nand U11771 (N_11771,N_10598,N_10705);
nand U11772 (N_11772,N_11224,N_11193);
or U11773 (N_11773,N_11196,N_10649);
or U11774 (N_11774,N_10568,N_10990);
or U11775 (N_11775,N_10768,N_11026);
and U11776 (N_11776,N_11005,N_11071);
or U11777 (N_11777,N_11059,N_11043);
nand U11778 (N_11778,N_10958,N_10501);
nand U11779 (N_11779,N_11190,N_10618);
nor U11780 (N_11780,N_11124,N_10639);
xnor U11781 (N_11781,N_10986,N_10864);
nand U11782 (N_11782,N_10646,N_10726);
nand U11783 (N_11783,N_10576,N_10954);
nor U11784 (N_11784,N_11018,N_10867);
or U11785 (N_11785,N_11236,N_10656);
and U11786 (N_11786,N_10995,N_10579);
nor U11787 (N_11787,N_11184,N_10813);
xor U11788 (N_11788,N_10878,N_11146);
or U11789 (N_11789,N_10900,N_10854);
xnor U11790 (N_11790,N_10985,N_10899);
nor U11791 (N_11791,N_10930,N_10632);
nor U11792 (N_11792,N_10528,N_11244);
and U11793 (N_11793,N_10927,N_10909);
nand U11794 (N_11794,N_11189,N_10798);
nor U11795 (N_11795,N_10676,N_10851);
xnor U11796 (N_11796,N_10945,N_10647);
or U11797 (N_11797,N_10573,N_10916);
xnor U11798 (N_11798,N_10536,N_10902);
nand U11799 (N_11799,N_10748,N_11004);
and U11800 (N_11800,N_10504,N_10928);
xor U11801 (N_11801,N_11130,N_11020);
and U11802 (N_11802,N_11080,N_11174);
or U11803 (N_11803,N_10774,N_10521);
nand U11804 (N_11804,N_11182,N_10768);
xnor U11805 (N_11805,N_11119,N_11093);
nor U11806 (N_11806,N_10701,N_10705);
xor U11807 (N_11807,N_11151,N_10823);
nor U11808 (N_11808,N_11129,N_11074);
xnor U11809 (N_11809,N_10513,N_10569);
and U11810 (N_11810,N_11095,N_11068);
xnor U11811 (N_11811,N_10966,N_10947);
or U11812 (N_11812,N_10991,N_11010);
nand U11813 (N_11813,N_10631,N_11135);
and U11814 (N_11814,N_11227,N_10871);
xor U11815 (N_11815,N_10551,N_10739);
nor U11816 (N_11816,N_10925,N_10982);
xnor U11817 (N_11817,N_10729,N_10673);
nand U11818 (N_11818,N_10508,N_10616);
xor U11819 (N_11819,N_10911,N_10591);
and U11820 (N_11820,N_10563,N_10578);
or U11821 (N_11821,N_10907,N_11155);
and U11822 (N_11822,N_10697,N_10659);
nor U11823 (N_11823,N_11182,N_10565);
nand U11824 (N_11824,N_10633,N_10609);
or U11825 (N_11825,N_11118,N_10634);
nor U11826 (N_11826,N_10987,N_11182);
and U11827 (N_11827,N_10507,N_10790);
xnor U11828 (N_11828,N_10602,N_10693);
or U11829 (N_11829,N_10552,N_10696);
and U11830 (N_11830,N_10737,N_11021);
and U11831 (N_11831,N_10866,N_11088);
nand U11832 (N_11832,N_11170,N_11129);
nand U11833 (N_11833,N_10852,N_11058);
nand U11834 (N_11834,N_10842,N_10854);
xor U11835 (N_11835,N_11137,N_10707);
xnor U11836 (N_11836,N_10633,N_11144);
nand U11837 (N_11837,N_10838,N_10930);
and U11838 (N_11838,N_10576,N_10647);
nor U11839 (N_11839,N_10849,N_11097);
xor U11840 (N_11840,N_10774,N_10590);
xnor U11841 (N_11841,N_10782,N_11202);
and U11842 (N_11842,N_10580,N_10745);
nand U11843 (N_11843,N_10509,N_10631);
nand U11844 (N_11844,N_10814,N_11236);
or U11845 (N_11845,N_10684,N_10988);
or U11846 (N_11846,N_10836,N_10875);
nand U11847 (N_11847,N_10616,N_10945);
and U11848 (N_11848,N_11236,N_10526);
xor U11849 (N_11849,N_10917,N_10765);
xor U11850 (N_11850,N_11194,N_10854);
nor U11851 (N_11851,N_10645,N_11228);
and U11852 (N_11852,N_10709,N_10701);
and U11853 (N_11853,N_10697,N_10944);
xor U11854 (N_11854,N_10839,N_10707);
and U11855 (N_11855,N_10914,N_11139);
or U11856 (N_11856,N_11212,N_11093);
nor U11857 (N_11857,N_10761,N_11058);
nor U11858 (N_11858,N_10577,N_11201);
or U11859 (N_11859,N_10959,N_10645);
xor U11860 (N_11860,N_10712,N_11150);
xnor U11861 (N_11861,N_10955,N_10939);
nor U11862 (N_11862,N_11129,N_10550);
nand U11863 (N_11863,N_10740,N_10569);
xnor U11864 (N_11864,N_10922,N_10828);
nand U11865 (N_11865,N_10730,N_11085);
nor U11866 (N_11866,N_10933,N_10562);
nor U11867 (N_11867,N_11146,N_10922);
nor U11868 (N_11868,N_10714,N_10947);
xnor U11869 (N_11869,N_11011,N_10841);
or U11870 (N_11870,N_10629,N_10713);
nor U11871 (N_11871,N_10743,N_10806);
xnor U11872 (N_11872,N_10583,N_11026);
nor U11873 (N_11873,N_10731,N_11135);
xor U11874 (N_11874,N_10645,N_10734);
xor U11875 (N_11875,N_10718,N_10934);
nand U11876 (N_11876,N_10573,N_10545);
nor U11877 (N_11877,N_11225,N_10705);
and U11878 (N_11878,N_10909,N_10889);
xor U11879 (N_11879,N_10929,N_11212);
or U11880 (N_11880,N_10600,N_10521);
or U11881 (N_11881,N_11070,N_10626);
and U11882 (N_11882,N_10857,N_11114);
or U11883 (N_11883,N_10609,N_10831);
xnor U11884 (N_11884,N_10589,N_11074);
nor U11885 (N_11885,N_10564,N_10626);
nor U11886 (N_11886,N_10653,N_11127);
nand U11887 (N_11887,N_11101,N_11177);
nor U11888 (N_11888,N_11014,N_10565);
or U11889 (N_11889,N_11185,N_10561);
or U11890 (N_11890,N_10730,N_10702);
xnor U11891 (N_11891,N_10767,N_11117);
xor U11892 (N_11892,N_10942,N_10992);
or U11893 (N_11893,N_11039,N_11184);
xnor U11894 (N_11894,N_10884,N_10760);
and U11895 (N_11895,N_10866,N_10835);
and U11896 (N_11896,N_11049,N_11032);
and U11897 (N_11897,N_10764,N_11029);
xor U11898 (N_11898,N_10549,N_10974);
xor U11899 (N_11899,N_10525,N_11097);
xnor U11900 (N_11900,N_11202,N_11177);
nor U11901 (N_11901,N_10761,N_10718);
nand U11902 (N_11902,N_10509,N_10785);
and U11903 (N_11903,N_11086,N_11185);
xor U11904 (N_11904,N_11207,N_11173);
nor U11905 (N_11905,N_10563,N_10827);
or U11906 (N_11906,N_10815,N_10658);
and U11907 (N_11907,N_10742,N_11093);
and U11908 (N_11908,N_11053,N_10966);
and U11909 (N_11909,N_10549,N_10874);
nand U11910 (N_11910,N_10831,N_10972);
nand U11911 (N_11911,N_10619,N_10646);
nand U11912 (N_11912,N_10651,N_10869);
and U11913 (N_11913,N_10627,N_11226);
xnor U11914 (N_11914,N_10966,N_11162);
nor U11915 (N_11915,N_10799,N_10715);
and U11916 (N_11916,N_11233,N_10685);
or U11917 (N_11917,N_10957,N_10915);
nand U11918 (N_11918,N_11000,N_10716);
or U11919 (N_11919,N_10822,N_10840);
nor U11920 (N_11920,N_10542,N_11249);
xor U11921 (N_11921,N_10709,N_10600);
xor U11922 (N_11922,N_11057,N_10542);
and U11923 (N_11923,N_11047,N_10921);
nor U11924 (N_11924,N_11078,N_10760);
and U11925 (N_11925,N_10989,N_10580);
xnor U11926 (N_11926,N_11213,N_11171);
xnor U11927 (N_11927,N_11070,N_11099);
nand U11928 (N_11928,N_10653,N_10726);
xor U11929 (N_11929,N_10729,N_10650);
xor U11930 (N_11930,N_10698,N_10742);
xor U11931 (N_11931,N_11157,N_10920);
and U11932 (N_11932,N_10513,N_10936);
and U11933 (N_11933,N_10896,N_10755);
or U11934 (N_11934,N_10913,N_10566);
or U11935 (N_11935,N_10762,N_11133);
nor U11936 (N_11936,N_10696,N_11231);
nor U11937 (N_11937,N_10784,N_11230);
and U11938 (N_11938,N_10941,N_10884);
xnor U11939 (N_11939,N_11174,N_11023);
and U11940 (N_11940,N_10642,N_10928);
or U11941 (N_11941,N_10736,N_11124);
xnor U11942 (N_11942,N_10514,N_10906);
and U11943 (N_11943,N_10866,N_10800);
nor U11944 (N_11944,N_10988,N_11218);
xnor U11945 (N_11945,N_10621,N_10904);
xnor U11946 (N_11946,N_10968,N_11110);
and U11947 (N_11947,N_10718,N_10533);
xor U11948 (N_11948,N_10818,N_10786);
nand U11949 (N_11949,N_11172,N_11011);
xnor U11950 (N_11950,N_11044,N_10598);
xnor U11951 (N_11951,N_10527,N_10686);
or U11952 (N_11952,N_10937,N_10999);
and U11953 (N_11953,N_11033,N_10955);
nand U11954 (N_11954,N_10664,N_10577);
nor U11955 (N_11955,N_10577,N_10901);
and U11956 (N_11956,N_10856,N_10581);
or U11957 (N_11957,N_10999,N_10595);
and U11958 (N_11958,N_10810,N_10841);
or U11959 (N_11959,N_10846,N_10609);
and U11960 (N_11960,N_10852,N_10857);
and U11961 (N_11961,N_10938,N_10701);
and U11962 (N_11962,N_10923,N_10932);
nand U11963 (N_11963,N_10797,N_11003);
and U11964 (N_11964,N_10588,N_11248);
xor U11965 (N_11965,N_10654,N_11046);
nand U11966 (N_11966,N_10718,N_10864);
or U11967 (N_11967,N_11117,N_10501);
and U11968 (N_11968,N_11005,N_10760);
xor U11969 (N_11969,N_10870,N_10701);
or U11970 (N_11970,N_11056,N_10887);
and U11971 (N_11971,N_10620,N_10990);
xor U11972 (N_11972,N_10693,N_11161);
xor U11973 (N_11973,N_10736,N_11159);
xor U11974 (N_11974,N_10684,N_10984);
nor U11975 (N_11975,N_10864,N_10657);
nand U11976 (N_11976,N_10511,N_10847);
nand U11977 (N_11977,N_10837,N_11093);
nor U11978 (N_11978,N_11101,N_10501);
or U11979 (N_11979,N_10636,N_11162);
xnor U11980 (N_11980,N_11062,N_10614);
or U11981 (N_11981,N_11142,N_10534);
nand U11982 (N_11982,N_10700,N_11079);
nand U11983 (N_11983,N_10816,N_11037);
or U11984 (N_11984,N_10660,N_11130);
nor U11985 (N_11985,N_10506,N_11159);
or U11986 (N_11986,N_11215,N_11115);
and U11987 (N_11987,N_11023,N_10584);
nand U11988 (N_11988,N_11065,N_10632);
xnor U11989 (N_11989,N_10583,N_10805);
nand U11990 (N_11990,N_10681,N_10733);
nand U11991 (N_11991,N_10702,N_10986);
xnor U11992 (N_11992,N_10851,N_10734);
nand U11993 (N_11993,N_11177,N_11146);
nor U11994 (N_11994,N_11003,N_10643);
nand U11995 (N_11995,N_10540,N_10780);
nand U11996 (N_11996,N_11189,N_10942);
nor U11997 (N_11997,N_10611,N_11060);
nand U11998 (N_11998,N_10500,N_11150);
xnor U11999 (N_11999,N_11053,N_11182);
nor U12000 (N_12000,N_11471,N_11761);
or U12001 (N_12001,N_11920,N_11676);
nand U12002 (N_12002,N_11685,N_11802);
and U12003 (N_12003,N_11546,N_11704);
nand U12004 (N_12004,N_11492,N_11635);
xor U12005 (N_12005,N_11860,N_11778);
xnor U12006 (N_12006,N_11381,N_11719);
and U12007 (N_12007,N_11942,N_11820);
or U12008 (N_12008,N_11638,N_11564);
and U12009 (N_12009,N_11464,N_11305);
xor U12010 (N_12010,N_11251,N_11895);
xor U12011 (N_12011,N_11536,N_11818);
nand U12012 (N_12012,N_11827,N_11526);
and U12013 (N_12013,N_11801,N_11613);
xor U12014 (N_12014,N_11530,N_11923);
nor U12015 (N_12015,N_11968,N_11750);
nor U12016 (N_12016,N_11290,N_11337);
nand U12017 (N_12017,N_11634,N_11382);
nand U12018 (N_12018,N_11545,N_11787);
nor U12019 (N_12019,N_11569,N_11748);
or U12020 (N_12020,N_11534,N_11419);
xor U12021 (N_12021,N_11854,N_11932);
xor U12022 (N_12022,N_11769,N_11675);
xnor U12023 (N_12023,N_11507,N_11378);
or U12024 (N_12024,N_11570,N_11962);
nor U12025 (N_12025,N_11706,N_11847);
or U12026 (N_12026,N_11799,N_11559);
nand U12027 (N_12027,N_11298,N_11728);
nor U12028 (N_12028,N_11425,N_11652);
xor U12029 (N_12029,N_11605,N_11259);
and U12030 (N_12030,N_11985,N_11404);
xnor U12031 (N_12031,N_11930,N_11292);
or U12032 (N_12032,N_11301,N_11568);
or U12033 (N_12033,N_11928,N_11496);
or U12034 (N_12034,N_11549,N_11880);
nor U12035 (N_12035,N_11308,N_11899);
nor U12036 (N_12036,N_11734,N_11736);
nor U12037 (N_12037,N_11870,N_11966);
nor U12038 (N_12038,N_11480,N_11817);
or U12039 (N_12039,N_11947,N_11868);
and U12040 (N_12040,N_11636,N_11552);
xnor U12041 (N_12041,N_11272,N_11421);
nand U12042 (N_12042,N_11410,N_11918);
nor U12043 (N_12043,N_11285,N_11705);
or U12044 (N_12044,N_11758,N_11729);
xnor U12045 (N_12045,N_11774,N_11806);
and U12046 (N_12046,N_11663,N_11318);
or U12047 (N_12047,N_11535,N_11521);
xor U12048 (N_12048,N_11463,N_11882);
xnor U12049 (N_12049,N_11803,N_11621);
xor U12050 (N_12050,N_11694,N_11789);
nand U12051 (N_12051,N_11885,N_11999);
nand U12052 (N_12052,N_11565,N_11762);
nor U12053 (N_12053,N_11374,N_11629);
nand U12054 (N_12054,N_11493,N_11864);
xor U12055 (N_12055,N_11708,N_11996);
xnor U12056 (N_12056,N_11586,N_11367);
nor U12057 (N_12057,N_11749,N_11357);
xnor U12058 (N_12058,N_11506,N_11261);
or U12059 (N_12059,N_11597,N_11341);
and U12060 (N_12060,N_11435,N_11953);
nor U12061 (N_12061,N_11933,N_11399);
or U12062 (N_12062,N_11366,N_11595);
nand U12063 (N_12063,N_11566,N_11403);
and U12064 (N_12064,N_11945,N_11458);
nor U12065 (N_12065,N_11743,N_11328);
or U12066 (N_12066,N_11361,N_11960);
and U12067 (N_12067,N_11735,N_11585);
and U12068 (N_12068,N_11839,N_11959);
nand U12069 (N_12069,N_11262,N_11335);
xor U12070 (N_12070,N_11865,N_11423);
nor U12071 (N_12071,N_11297,N_11776);
nor U12072 (N_12072,N_11619,N_11445);
or U12073 (N_12073,N_11725,N_11876);
or U12074 (N_12074,N_11352,N_11469);
nor U12075 (N_12075,N_11791,N_11383);
nand U12076 (N_12076,N_11655,N_11974);
and U12077 (N_12077,N_11909,N_11257);
or U12078 (N_12078,N_11772,N_11793);
nand U12079 (N_12079,N_11937,N_11656);
xnor U12080 (N_12080,N_11944,N_11970);
and U12081 (N_12081,N_11353,N_11583);
xnor U12082 (N_12082,N_11726,N_11926);
xnor U12083 (N_12083,N_11805,N_11855);
and U12084 (N_12084,N_11409,N_11911);
and U12085 (N_12085,N_11919,N_11543);
nand U12086 (N_12086,N_11287,N_11714);
or U12087 (N_12087,N_11258,N_11473);
xnor U12088 (N_12088,N_11482,N_11594);
or U12089 (N_12089,N_11830,N_11896);
nor U12090 (N_12090,N_11835,N_11276);
nand U12091 (N_12091,N_11329,N_11338);
xnor U12092 (N_12092,N_11697,N_11266);
xor U12093 (N_12093,N_11336,N_11505);
or U12094 (N_12094,N_11269,N_11551);
xnor U12095 (N_12095,N_11432,N_11498);
or U12096 (N_12096,N_11842,N_11649);
xor U12097 (N_12097,N_11707,N_11304);
or U12098 (N_12098,N_11296,N_11980);
and U12099 (N_12099,N_11373,N_11641);
nor U12100 (N_12100,N_11683,N_11653);
nor U12101 (N_12101,N_11412,N_11288);
and U12102 (N_12102,N_11540,N_11913);
and U12103 (N_12103,N_11742,N_11508);
xor U12104 (N_12104,N_11350,N_11879);
nor U12105 (N_12105,N_11345,N_11912);
or U12106 (N_12106,N_11522,N_11739);
and U12107 (N_12107,N_11533,N_11394);
or U12108 (N_12108,N_11718,N_11836);
and U12109 (N_12109,N_11981,N_11558);
nor U12110 (N_12110,N_11833,N_11686);
and U12111 (N_12111,N_11299,N_11823);
nor U12112 (N_12112,N_11972,N_11364);
nor U12113 (N_12113,N_11733,N_11950);
nand U12114 (N_12114,N_11720,N_11756);
nand U12115 (N_12115,N_11574,N_11989);
nand U12116 (N_12116,N_11388,N_11359);
nor U12117 (N_12117,N_11859,N_11666);
nor U12118 (N_12118,N_11593,N_11914);
nor U12119 (N_12119,N_11523,N_11715);
nand U12120 (N_12120,N_11851,N_11936);
nor U12121 (N_12121,N_11516,N_11282);
xor U12122 (N_12122,N_11503,N_11547);
nor U12123 (N_12123,N_11467,N_11658);
nor U12124 (N_12124,N_11938,N_11598);
or U12125 (N_12125,N_11783,N_11422);
nand U12126 (N_12126,N_11396,N_11407);
and U12127 (N_12127,N_11339,N_11444);
nand U12128 (N_12128,N_11529,N_11518);
nand U12129 (N_12129,N_11307,N_11954);
nor U12130 (N_12130,N_11362,N_11541);
nand U12131 (N_12131,N_11478,N_11963);
and U12132 (N_12132,N_11887,N_11376);
nand U12133 (N_12133,N_11600,N_11810);
nor U12134 (N_12134,N_11692,N_11703);
xnor U12135 (N_12135,N_11838,N_11527);
nor U12136 (N_12136,N_11767,N_11916);
xor U12137 (N_12137,N_11908,N_11857);
nand U12138 (N_12138,N_11948,N_11821);
and U12139 (N_12139,N_11757,N_11456);
nor U12140 (N_12140,N_11796,N_11606);
and U12141 (N_12141,N_11517,N_11389);
nor U12142 (N_12142,N_11866,N_11490);
nand U12143 (N_12143,N_11252,N_11662);
nand U12144 (N_12144,N_11607,N_11271);
nor U12145 (N_12145,N_11939,N_11539);
xor U12146 (N_12146,N_11631,N_11700);
nor U12147 (N_12147,N_11599,N_11524);
nand U12148 (N_12148,N_11609,N_11431);
nor U12149 (N_12149,N_11878,N_11580);
xor U12150 (N_12150,N_11779,N_11455);
nor U12151 (N_12151,N_11843,N_11532);
or U12152 (N_12152,N_11765,N_11380);
nand U12153 (N_12153,N_11509,N_11957);
xnor U12154 (N_12154,N_11964,N_11481);
nand U12155 (N_12155,N_11483,N_11832);
and U12156 (N_12156,N_11804,N_11317);
and U12157 (N_12157,N_11618,N_11512);
and U12158 (N_12158,N_11997,N_11602);
nand U12159 (N_12159,N_11354,N_11905);
or U12160 (N_12160,N_11661,N_11453);
and U12161 (N_12161,N_11608,N_11672);
or U12162 (N_12162,N_11500,N_11751);
nor U12163 (N_12163,N_11753,N_11659);
and U12164 (N_12164,N_11293,N_11253);
nand U12165 (N_12165,N_11592,N_11745);
and U12166 (N_12166,N_11993,N_11616);
or U12167 (N_12167,N_11763,N_11889);
nor U12168 (N_12168,N_11504,N_11371);
or U12169 (N_12169,N_11312,N_11465);
nand U12170 (N_12170,N_11794,N_11554);
xor U12171 (N_12171,N_11561,N_11732);
nor U12172 (N_12172,N_11447,N_11398);
nor U12173 (N_12173,N_11446,N_11320);
and U12174 (N_12174,N_11520,N_11433);
or U12175 (N_12175,N_11768,N_11679);
nor U12176 (N_12176,N_11347,N_11982);
xor U12177 (N_12177,N_11846,N_11844);
nand U12178 (N_12178,N_11956,N_11958);
and U12179 (N_12179,N_11411,N_11440);
nor U12180 (N_12180,N_11395,N_11727);
and U12181 (N_12181,N_11784,N_11510);
nand U12182 (N_12182,N_11610,N_11591);
or U12183 (N_12183,N_11420,N_11901);
nand U12184 (N_12184,N_11850,N_11701);
and U12185 (N_12185,N_11929,N_11265);
and U12186 (N_12186,N_11922,N_11489);
and U12187 (N_12187,N_11548,N_11746);
or U12188 (N_12188,N_11562,N_11589);
and U12189 (N_12189,N_11286,N_11484);
nand U12190 (N_12190,N_11849,N_11623);
and U12191 (N_12191,N_11946,N_11436);
or U12192 (N_12192,N_11990,N_11691);
nand U12193 (N_12193,N_11837,N_11637);
or U12194 (N_12194,N_11978,N_11786);
nor U12195 (N_12195,N_11397,N_11824);
nor U12196 (N_12196,N_11925,N_11760);
nand U12197 (N_12197,N_11906,N_11826);
or U12198 (N_12198,N_11379,N_11319);
or U12199 (N_12199,N_11903,N_11370);
xnor U12200 (N_12200,N_11664,N_11788);
or U12201 (N_12201,N_11684,N_11582);
and U12202 (N_12202,N_11537,N_11441);
and U12203 (N_12203,N_11386,N_11528);
xor U12204 (N_12204,N_11965,N_11759);
or U12205 (N_12205,N_11384,N_11571);
or U12206 (N_12206,N_11501,N_11798);
xor U12207 (N_12207,N_11951,N_11323);
and U12208 (N_12208,N_11375,N_11674);
nand U12209 (N_12209,N_11800,N_11888);
or U12210 (N_12210,N_11983,N_11660);
nand U12211 (N_12211,N_11274,N_11325);
or U12212 (N_12212,N_11315,N_11316);
xnor U12213 (N_12213,N_11741,N_11314);
and U12214 (N_12214,N_11814,N_11256);
and U12215 (N_12215,N_11434,N_11499);
or U12216 (N_12216,N_11356,N_11724);
nor U12217 (N_12217,N_11615,N_11690);
xnor U12218 (N_12218,N_11390,N_11514);
nand U12219 (N_12219,N_11809,N_11563);
or U12220 (N_12220,N_11852,N_11740);
xnor U12221 (N_12221,N_11931,N_11342);
nor U12222 (N_12222,N_11355,N_11416);
nand U12223 (N_12223,N_11576,N_11770);
and U12224 (N_12224,N_11967,N_11639);
xnor U12225 (N_12225,N_11702,N_11494);
xor U12226 (N_12226,N_11330,N_11603);
and U12227 (N_12227,N_11472,N_11834);
xor U12228 (N_12228,N_11327,N_11747);
nor U12229 (N_12229,N_11738,N_11369);
nor U12230 (N_12230,N_11991,N_11579);
nand U12231 (N_12231,N_11813,N_11572);
and U12232 (N_12232,N_11898,N_11525);
nand U12233 (N_12233,N_11979,N_11279);
and U12234 (N_12234,N_11975,N_11477);
and U12235 (N_12235,N_11321,N_11792);
nor U12236 (N_12236,N_11542,N_11622);
or U12237 (N_12237,N_11401,N_11890);
nand U12238 (N_12238,N_11502,N_11437);
or U12239 (N_12239,N_11790,N_11428);
xor U12240 (N_12240,N_11952,N_11577);
nand U12241 (N_12241,N_11267,N_11300);
and U12242 (N_12242,N_11709,N_11450);
and U12243 (N_12243,N_11698,N_11626);
nor U12244 (N_12244,N_11311,N_11557);
and U12245 (N_12245,N_11680,N_11873);
xnor U12246 (N_12246,N_11681,N_11587);
or U12247 (N_12247,N_11448,N_11581);
nor U12248 (N_12248,N_11358,N_11955);
xnor U12249 (N_12249,N_11313,N_11306);
nand U12250 (N_12250,N_11668,N_11977);
or U12251 (N_12251,N_11488,N_11961);
or U12252 (N_12252,N_11984,N_11816);
xnor U12253 (N_12253,N_11877,N_11573);
xnor U12254 (N_12254,N_11567,N_11902);
or U12255 (N_12255,N_11716,N_11822);
and U12256 (N_12256,N_11466,N_11643);
nor U12257 (N_12257,N_11863,N_11949);
nand U12258 (N_12258,N_11487,N_11730);
nand U12259 (N_12259,N_11332,N_11695);
or U12260 (N_12260,N_11644,N_11891);
nor U12261 (N_12261,N_11755,N_11400);
and U12262 (N_12262,N_11413,N_11575);
xor U12263 (N_12263,N_11969,N_11277);
xnor U12264 (N_12264,N_11721,N_11309);
or U12265 (N_12265,N_11874,N_11344);
or U12266 (N_12266,N_11710,N_11302);
nor U12267 (N_12267,N_11976,N_11673);
and U12268 (N_12268,N_11550,N_11722);
and U12269 (N_12269,N_11921,N_11544);
nand U12270 (N_12270,N_11845,N_11775);
nand U12271 (N_12271,N_11712,N_11654);
nand U12272 (N_12272,N_11442,N_11785);
and U12273 (N_12273,N_11867,N_11825);
xnor U12274 (N_12274,N_11333,N_11897);
or U12275 (N_12275,N_11538,N_11491);
or U12276 (N_12276,N_11858,N_11417);
xor U12277 (N_12277,N_11270,N_11987);
nand U12278 (N_12278,N_11689,N_11254);
nor U12279 (N_12279,N_11457,N_11268);
nand U12280 (N_12280,N_11872,N_11360);
and U12281 (N_12281,N_11754,N_11497);
and U12282 (N_12282,N_11351,N_11614);
nor U12283 (N_12283,N_11295,N_11343);
and U12284 (N_12284,N_11828,N_11699);
xor U12285 (N_12285,N_11627,N_11862);
and U12286 (N_12286,N_11829,N_11310);
nand U12287 (N_12287,N_11630,N_11250);
nor U12288 (N_12288,N_11764,N_11515);
nand U12289 (N_12289,N_11531,N_11443);
nand U12290 (N_12290,N_11495,N_11875);
or U12291 (N_12291,N_11640,N_11555);
or U12292 (N_12292,N_11628,N_11596);
nand U12293 (N_12293,N_11625,N_11646);
xnor U12294 (N_12294,N_11284,N_11590);
nand U12295 (N_12295,N_11476,N_11438);
nor U12296 (N_12296,N_11519,N_11841);
nand U12297 (N_12297,N_11263,N_11894);
nand U12298 (N_12298,N_11780,N_11831);
and U12299 (N_12299,N_11781,N_11893);
or U12300 (N_12300,N_11807,N_11475);
xor U12301 (N_12301,N_11853,N_11324);
and U12302 (N_12302,N_11869,N_11795);
nor U12303 (N_12303,N_11449,N_11439);
and U12304 (N_12304,N_11924,N_11424);
or U12305 (N_12305,N_11688,N_11604);
or U12306 (N_12306,N_11943,N_11601);
xnor U12307 (N_12307,N_11459,N_11462);
or U12308 (N_12308,N_11995,N_11647);
nor U12309 (N_12309,N_11348,N_11346);
nand U12310 (N_12310,N_11840,N_11405);
nor U12311 (N_12311,N_11998,N_11886);
or U12312 (N_12312,N_11992,N_11452);
nand U12313 (N_12313,N_11468,N_11340);
nand U12314 (N_12314,N_11915,N_11986);
nor U12315 (N_12315,N_11460,N_11291);
nand U12316 (N_12316,N_11402,N_11486);
xnor U12317 (N_12317,N_11578,N_11273);
nor U12318 (N_12318,N_11940,N_11260);
and U12319 (N_12319,N_11651,N_11892);
or U12320 (N_12320,N_11281,N_11766);
xor U12321 (N_12321,N_11648,N_11331);
nor U12322 (N_12322,N_11612,N_11669);
or U12323 (N_12323,N_11861,N_11665);
and U12324 (N_12324,N_11255,N_11934);
or U12325 (N_12325,N_11624,N_11650);
nor U12326 (N_12326,N_11797,N_11927);
xor U12327 (N_12327,N_11771,N_11904);
nor U12328 (N_12328,N_11811,N_11871);
nand U12329 (N_12329,N_11611,N_11696);
xor U12330 (N_12330,N_11988,N_11429);
xor U12331 (N_12331,N_11556,N_11479);
and U12332 (N_12332,N_11682,N_11645);
nand U12333 (N_12333,N_11819,N_11671);
and U12334 (N_12334,N_11670,N_11617);
nor U12335 (N_12335,N_11667,N_11289);
nor U12336 (N_12336,N_11744,N_11657);
or U12337 (N_12337,N_11884,N_11474);
nand U12338 (N_12338,N_11278,N_11994);
or U12339 (N_12339,N_11264,N_11451);
nand U12340 (N_12340,N_11415,N_11678);
nand U12341 (N_12341,N_11303,N_11368);
xor U12342 (N_12342,N_11426,N_11363);
xnor U12343 (N_12343,N_11454,N_11848);
or U12344 (N_12344,N_11935,N_11385);
nor U12345 (N_12345,N_11427,N_11632);
or U12346 (N_12346,N_11283,N_11275);
xor U12347 (N_12347,N_11377,N_11808);
nor U12348 (N_12348,N_11642,N_11365);
xnor U12349 (N_12349,N_11941,N_11711);
nor U12350 (N_12350,N_11917,N_11971);
or U12351 (N_12351,N_11881,N_11372);
or U12352 (N_12352,N_11815,N_11334);
or U12353 (N_12353,N_11731,N_11633);
nand U12354 (N_12354,N_11470,N_11553);
or U12355 (N_12355,N_11391,N_11883);
xnor U12356 (N_12356,N_11693,N_11687);
nand U12357 (N_12357,N_11737,N_11752);
xor U12358 (N_12358,N_11406,N_11408);
nor U12359 (N_12359,N_11900,N_11584);
and U12360 (N_12360,N_11973,N_11812);
nor U12361 (N_12361,N_11588,N_11717);
and U12362 (N_12362,N_11713,N_11485);
xor U12363 (N_12363,N_11560,N_11387);
and U12364 (N_12364,N_11782,N_11461);
or U12365 (N_12365,N_11910,N_11677);
nand U12366 (N_12366,N_11907,N_11773);
nand U12367 (N_12367,N_11511,N_11393);
nand U12368 (N_12368,N_11326,N_11777);
or U12369 (N_12369,N_11392,N_11414);
or U12370 (N_12370,N_11349,N_11294);
and U12371 (N_12371,N_11430,N_11322);
xnor U12372 (N_12372,N_11620,N_11418);
and U12373 (N_12373,N_11856,N_11513);
nor U12374 (N_12374,N_11723,N_11280);
nand U12375 (N_12375,N_11275,N_11437);
xnor U12376 (N_12376,N_11799,N_11864);
nor U12377 (N_12377,N_11352,N_11423);
and U12378 (N_12378,N_11334,N_11989);
nor U12379 (N_12379,N_11668,N_11917);
xor U12380 (N_12380,N_11416,N_11970);
nand U12381 (N_12381,N_11786,N_11600);
or U12382 (N_12382,N_11465,N_11734);
and U12383 (N_12383,N_11768,N_11570);
or U12384 (N_12384,N_11887,N_11751);
or U12385 (N_12385,N_11979,N_11994);
nor U12386 (N_12386,N_11419,N_11340);
xnor U12387 (N_12387,N_11459,N_11563);
nand U12388 (N_12388,N_11871,N_11762);
and U12389 (N_12389,N_11599,N_11255);
and U12390 (N_12390,N_11783,N_11618);
and U12391 (N_12391,N_11584,N_11565);
or U12392 (N_12392,N_11615,N_11938);
nand U12393 (N_12393,N_11460,N_11650);
nor U12394 (N_12394,N_11658,N_11448);
nor U12395 (N_12395,N_11442,N_11781);
xnor U12396 (N_12396,N_11875,N_11857);
nand U12397 (N_12397,N_11448,N_11424);
or U12398 (N_12398,N_11826,N_11691);
xnor U12399 (N_12399,N_11293,N_11756);
nor U12400 (N_12400,N_11523,N_11252);
nand U12401 (N_12401,N_11281,N_11481);
xor U12402 (N_12402,N_11720,N_11787);
xor U12403 (N_12403,N_11455,N_11351);
and U12404 (N_12404,N_11653,N_11776);
or U12405 (N_12405,N_11860,N_11927);
nor U12406 (N_12406,N_11469,N_11970);
or U12407 (N_12407,N_11348,N_11733);
xnor U12408 (N_12408,N_11494,N_11451);
nand U12409 (N_12409,N_11461,N_11616);
and U12410 (N_12410,N_11330,N_11739);
and U12411 (N_12411,N_11712,N_11649);
and U12412 (N_12412,N_11373,N_11630);
nor U12413 (N_12413,N_11624,N_11466);
nor U12414 (N_12414,N_11921,N_11907);
and U12415 (N_12415,N_11517,N_11509);
nor U12416 (N_12416,N_11650,N_11807);
or U12417 (N_12417,N_11799,N_11694);
nand U12418 (N_12418,N_11720,N_11580);
or U12419 (N_12419,N_11286,N_11618);
nand U12420 (N_12420,N_11355,N_11828);
nand U12421 (N_12421,N_11533,N_11575);
and U12422 (N_12422,N_11892,N_11284);
and U12423 (N_12423,N_11506,N_11526);
xor U12424 (N_12424,N_11278,N_11435);
nand U12425 (N_12425,N_11459,N_11271);
xnor U12426 (N_12426,N_11800,N_11665);
nand U12427 (N_12427,N_11890,N_11425);
xnor U12428 (N_12428,N_11332,N_11590);
nor U12429 (N_12429,N_11680,N_11328);
or U12430 (N_12430,N_11489,N_11562);
or U12431 (N_12431,N_11827,N_11297);
xor U12432 (N_12432,N_11946,N_11755);
xor U12433 (N_12433,N_11871,N_11663);
nor U12434 (N_12434,N_11463,N_11920);
nor U12435 (N_12435,N_11361,N_11672);
or U12436 (N_12436,N_11687,N_11714);
and U12437 (N_12437,N_11894,N_11999);
xor U12438 (N_12438,N_11865,N_11371);
nand U12439 (N_12439,N_11524,N_11614);
nand U12440 (N_12440,N_11378,N_11771);
nor U12441 (N_12441,N_11953,N_11547);
nand U12442 (N_12442,N_11769,N_11410);
and U12443 (N_12443,N_11467,N_11833);
and U12444 (N_12444,N_11965,N_11353);
nand U12445 (N_12445,N_11463,N_11887);
or U12446 (N_12446,N_11316,N_11405);
nand U12447 (N_12447,N_11618,N_11298);
or U12448 (N_12448,N_11262,N_11884);
xnor U12449 (N_12449,N_11548,N_11856);
xor U12450 (N_12450,N_11975,N_11650);
and U12451 (N_12451,N_11506,N_11268);
or U12452 (N_12452,N_11376,N_11495);
nor U12453 (N_12453,N_11422,N_11943);
nand U12454 (N_12454,N_11946,N_11339);
nand U12455 (N_12455,N_11906,N_11441);
nor U12456 (N_12456,N_11868,N_11973);
nand U12457 (N_12457,N_11878,N_11456);
xnor U12458 (N_12458,N_11411,N_11606);
nand U12459 (N_12459,N_11914,N_11771);
nor U12460 (N_12460,N_11924,N_11983);
and U12461 (N_12461,N_11887,N_11337);
xnor U12462 (N_12462,N_11684,N_11348);
xor U12463 (N_12463,N_11578,N_11837);
or U12464 (N_12464,N_11737,N_11789);
or U12465 (N_12465,N_11876,N_11680);
xor U12466 (N_12466,N_11856,N_11454);
nand U12467 (N_12467,N_11722,N_11980);
or U12468 (N_12468,N_11710,N_11642);
and U12469 (N_12469,N_11875,N_11810);
and U12470 (N_12470,N_11583,N_11526);
and U12471 (N_12471,N_11691,N_11993);
nand U12472 (N_12472,N_11537,N_11720);
xor U12473 (N_12473,N_11751,N_11619);
xnor U12474 (N_12474,N_11579,N_11947);
xnor U12475 (N_12475,N_11861,N_11544);
nand U12476 (N_12476,N_11803,N_11796);
nand U12477 (N_12477,N_11707,N_11840);
and U12478 (N_12478,N_11791,N_11452);
and U12479 (N_12479,N_11546,N_11762);
or U12480 (N_12480,N_11891,N_11952);
nor U12481 (N_12481,N_11992,N_11910);
and U12482 (N_12482,N_11298,N_11671);
nor U12483 (N_12483,N_11643,N_11809);
nand U12484 (N_12484,N_11814,N_11832);
nand U12485 (N_12485,N_11621,N_11494);
nand U12486 (N_12486,N_11737,N_11561);
nor U12487 (N_12487,N_11688,N_11390);
and U12488 (N_12488,N_11254,N_11555);
xor U12489 (N_12489,N_11846,N_11516);
nand U12490 (N_12490,N_11427,N_11851);
nand U12491 (N_12491,N_11498,N_11913);
xor U12492 (N_12492,N_11842,N_11357);
nor U12493 (N_12493,N_11492,N_11498);
nand U12494 (N_12494,N_11868,N_11296);
and U12495 (N_12495,N_11321,N_11758);
nor U12496 (N_12496,N_11368,N_11857);
nand U12497 (N_12497,N_11620,N_11816);
or U12498 (N_12498,N_11775,N_11770);
nor U12499 (N_12499,N_11451,N_11689);
xnor U12500 (N_12500,N_11328,N_11513);
xor U12501 (N_12501,N_11339,N_11254);
and U12502 (N_12502,N_11374,N_11746);
xnor U12503 (N_12503,N_11904,N_11394);
or U12504 (N_12504,N_11659,N_11530);
nand U12505 (N_12505,N_11459,N_11266);
xnor U12506 (N_12506,N_11442,N_11617);
nand U12507 (N_12507,N_11374,N_11642);
nor U12508 (N_12508,N_11562,N_11377);
nor U12509 (N_12509,N_11681,N_11450);
or U12510 (N_12510,N_11395,N_11740);
or U12511 (N_12511,N_11523,N_11776);
xor U12512 (N_12512,N_11419,N_11357);
nor U12513 (N_12513,N_11482,N_11763);
nor U12514 (N_12514,N_11718,N_11757);
nand U12515 (N_12515,N_11647,N_11360);
or U12516 (N_12516,N_11959,N_11546);
and U12517 (N_12517,N_11336,N_11862);
xor U12518 (N_12518,N_11420,N_11317);
and U12519 (N_12519,N_11440,N_11424);
nand U12520 (N_12520,N_11709,N_11725);
or U12521 (N_12521,N_11545,N_11899);
xnor U12522 (N_12522,N_11345,N_11968);
nand U12523 (N_12523,N_11387,N_11686);
nand U12524 (N_12524,N_11910,N_11865);
and U12525 (N_12525,N_11454,N_11617);
xor U12526 (N_12526,N_11393,N_11371);
or U12527 (N_12527,N_11888,N_11656);
nor U12528 (N_12528,N_11308,N_11415);
or U12529 (N_12529,N_11663,N_11598);
or U12530 (N_12530,N_11402,N_11460);
nand U12531 (N_12531,N_11735,N_11744);
and U12532 (N_12532,N_11926,N_11813);
and U12533 (N_12533,N_11315,N_11385);
or U12534 (N_12534,N_11535,N_11671);
or U12535 (N_12535,N_11755,N_11345);
nor U12536 (N_12536,N_11751,N_11963);
and U12537 (N_12537,N_11714,N_11407);
or U12538 (N_12538,N_11686,N_11637);
or U12539 (N_12539,N_11495,N_11347);
and U12540 (N_12540,N_11274,N_11256);
nor U12541 (N_12541,N_11624,N_11752);
or U12542 (N_12542,N_11928,N_11924);
nor U12543 (N_12543,N_11647,N_11483);
and U12544 (N_12544,N_11264,N_11487);
nor U12545 (N_12545,N_11737,N_11463);
nor U12546 (N_12546,N_11718,N_11917);
xnor U12547 (N_12547,N_11973,N_11545);
nand U12548 (N_12548,N_11303,N_11764);
or U12549 (N_12549,N_11822,N_11287);
or U12550 (N_12550,N_11265,N_11780);
nand U12551 (N_12551,N_11335,N_11717);
xor U12552 (N_12552,N_11721,N_11512);
xor U12553 (N_12553,N_11986,N_11630);
nand U12554 (N_12554,N_11779,N_11321);
nor U12555 (N_12555,N_11274,N_11962);
xnor U12556 (N_12556,N_11300,N_11626);
xor U12557 (N_12557,N_11820,N_11706);
or U12558 (N_12558,N_11345,N_11898);
or U12559 (N_12559,N_11869,N_11578);
nand U12560 (N_12560,N_11621,N_11721);
nand U12561 (N_12561,N_11977,N_11819);
and U12562 (N_12562,N_11528,N_11909);
xnor U12563 (N_12563,N_11621,N_11847);
and U12564 (N_12564,N_11447,N_11771);
nand U12565 (N_12565,N_11254,N_11872);
and U12566 (N_12566,N_11860,N_11354);
nor U12567 (N_12567,N_11687,N_11331);
nor U12568 (N_12568,N_11413,N_11991);
xnor U12569 (N_12569,N_11648,N_11861);
nor U12570 (N_12570,N_11989,N_11436);
nand U12571 (N_12571,N_11984,N_11894);
or U12572 (N_12572,N_11788,N_11880);
xnor U12573 (N_12573,N_11676,N_11504);
nand U12574 (N_12574,N_11874,N_11441);
xor U12575 (N_12575,N_11604,N_11374);
and U12576 (N_12576,N_11975,N_11718);
xnor U12577 (N_12577,N_11605,N_11373);
nor U12578 (N_12578,N_11623,N_11320);
nand U12579 (N_12579,N_11326,N_11986);
and U12580 (N_12580,N_11818,N_11829);
and U12581 (N_12581,N_11824,N_11688);
and U12582 (N_12582,N_11980,N_11736);
nor U12583 (N_12583,N_11508,N_11974);
or U12584 (N_12584,N_11392,N_11587);
xnor U12585 (N_12585,N_11811,N_11445);
nand U12586 (N_12586,N_11558,N_11330);
nand U12587 (N_12587,N_11883,N_11918);
and U12588 (N_12588,N_11987,N_11791);
and U12589 (N_12589,N_11949,N_11275);
xor U12590 (N_12590,N_11749,N_11732);
and U12591 (N_12591,N_11499,N_11649);
nor U12592 (N_12592,N_11277,N_11573);
nor U12593 (N_12593,N_11569,N_11740);
nor U12594 (N_12594,N_11478,N_11407);
xor U12595 (N_12595,N_11639,N_11685);
nand U12596 (N_12596,N_11616,N_11469);
or U12597 (N_12597,N_11301,N_11970);
nor U12598 (N_12598,N_11451,N_11712);
and U12599 (N_12599,N_11251,N_11734);
and U12600 (N_12600,N_11521,N_11963);
and U12601 (N_12601,N_11704,N_11462);
and U12602 (N_12602,N_11713,N_11665);
nor U12603 (N_12603,N_11299,N_11661);
xnor U12604 (N_12604,N_11395,N_11530);
and U12605 (N_12605,N_11606,N_11960);
and U12606 (N_12606,N_11680,N_11493);
and U12607 (N_12607,N_11595,N_11636);
and U12608 (N_12608,N_11924,N_11514);
or U12609 (N_12609,N_11978,N_11424);
and U12610 (N_12610,N_11443,N_11824);
or U12611 (N_12611,N_11732,N_11584);
nor U12612 (N_12612,N_11445,N_11829);
and U12613 (N_12613,N_11569,N_11793);
nor U12614 (N_12614,N_11291,N_11968);
nand U12615 (N_12615,N_11979,N_11569);
nor U12616 (N_12616,N_11426,N_11663);
or U12617 (N_12617,N_11295,N_11495);
and U12618 (N_12618,N_11956,N_11311);
nand U12619 (N_12619,N_11313,N_11858);
or U12620 (N_12620,N_11274,N_11698);
nand U12621 (N_12621,N_11941,N_11251);
or U12622 (N_12622,N_11610,N_11529);
nand U12623 (N_12623,N_11814,N_11792);
xor U12624 (N_12624,N_11937,N_11955);
xnor U12625 (N_12625,N_11969,N_11998);
or U12626 (N_12626,N_11724,N_11343);
nor U12627 (N_12627,N_11485,N_11860);
xor U12628 (N_12628,N_11452,N_11310);
nand U12629 (N_12629,N_11293,N_11273);
nand U12630 (N_12630,N_11415,N_11680);
or U12631 (N_12631,N_11753,N_11346);
or U12632 (N_12632,N_11502,N_11303);
nor U12633 (N_12633,N_11855,N_11296);
xor U12634 (N_12634,N_11853,N_11526);
or U12635 (N_12635,N_11554,N_11388);
nand U12636 (N_12636,N_11303,N_11914);
and U12637 (N_12637,N_11604,N_11641);
nor U12638 (N_12638,N_11794,N_11872);
xnor U12639 (N_12639,N_11784,N_11839);
nand U12640 (N_12640,N_11283,N_11258);
xor U12641 (N_12641,N_11729,N_11673);
and U12642 (N_12642,N_11428,N_11599);
nand U12643 (N_12643,N_11299,N_11608);
or U12644 (N_12644,N_11600,N_11760);
xnor U12645 (N_12645,N_11868,N_11585);
or U12646 (N_12646,N_11697,N_11396);
xnor U12647 (N_12647,N_11370,N_11491);
and U12648 (N_12648,N_11671,N_11880);
or U12649 (N_12649,N_11951,N_11887);
nand U12650 (N_12650,N_11786,N_11968);
or U12651 (N_12651,N_11847,N_11412);
xor U12652 (N_12652,N_11491,N_11832);
and U12653 (N_12653,N_11447,N_11601);
nand U12654 (N_12654,N_11538,N_11326);
nor U12655 (N_12655,N_11434,N_11276);
nand U12656 (N_12656,N_11253,N_11768);
xor U12657 (N_12657,N_11869,N_11750);
and U12658 (N_12658,N_11636,N_11740);
nor U12659 (N_12659,N_11607,N_11658);
nand U12660 (N_12660,N_11619,N_11899);
nor U12661 (N_12661,N_11558,N_11585);
xnor U12662 (N_12662,N_11393,N_11611);
or U12663 (N_12663,N_11755,N_11262);
or U12664 (N_12664,N_11403,N_11815);
nand U12665 (N_12665,N_11927,N_11783);
nor U12666 (N_12666,N_11664,N_11976);
nand U12667 (N_12667,N_11646,N_11321);
or U12668 (N_12668,N_11285,N_11424);
or U12669 (N_12669,N_11524,N_11813);
xor U12670 (N_12670,N_11400,N_11820);
xnor U12671 (N_12671,N_11412,N_11334);
nand U12672 (N_12672,N_11986,N_11997);
and U12673 (N_12673,N_11861,N_11479);
and U12674 (N_12674,N_11324,N_11972);
nand U12675 (N_12675,N_11865,N_11850);
nand U12676 (N_12676,N_11867,N_11934);
or U12677 (N_12677,N_11873,N_11798);
xor U12678 (N_12678,N_11951,N_11396);
nand U12679 (N_12679,N_11941,N_11813);
or U12680 (N_12680,N_11924,N_11299);
nor U12681 (N_12681,N_11442,N_11336);
and U12682 (N_12682,N_11825,N_11540);
and U12683 (N_12683,N_11524,N_11991);
or U12684 (N_12684,N_11656,N_11595);
nor U12685 (N_12685,N_11844,N_11838);
nand U12686 (N_12686,N_11850,N_11577);
and U12687 (N_12687,N_11339,N_11472);
or U12688 (N_12688,N_11828,N_11901);
nand U12689 (N_12689,N_11906,N_11498);
nand U12690 (N_12690,N_11572,N_11427);
nor U12691 (N_12691,N_11471,N_11947);
or U12692 (N_12692,N_11446,N_11673);
or U12693 (N_12693,N_11885,N_11553);
and U12694 (N_12694,N_11997,N_11701);
xnor U12695 (N_12695,N_11312,N_11667);
or U12696 (N_12696,N_11614,N_11789);
or U12697 (N_12697,N_11818,N_11379);
nand U12698 (N_12698,N_11689,N_11562);
nand U12699 (N_12699,N_11397,N_11871);
xor U12700 (N_12700,N_11464,N_11526);
or U12701 (N_12701,N_11970,N_11474);
and U12702 (N_12702,N_11645,N_11278);
and U12703 (N_12703,N_11885,N_11933);
nand U12704 (N_12704,N_11663,N_11280);
and U12705 (N_12705,N_11777,N_11607);
nand U12706 (N_12706,N_11748,N_11540);
nor U12707 (N_12707,N_11542,N_11719);
nor U12708 (N_12708,N_11390,N_11681);
or U12709 (N_12709,N_11880,N_11492);
nand U12710 (N_12710,N_11737,N_11813);
nor U12711 (N_12711,N_11550,N_11809);
xor U12712 (N_12712,N_11721,N_11491);
xnor U12713 (N_12713,N_11834,N_11776);
nand U12714 (N_12714,N_11753,N_11561);
nor U12715 (N_12715,N_11526,N_11685);
nand U12716 (N_12716,N_11719,N_11422);
xnor U12717 (N_12717,N_11523,N_11477);
xor U12718 (N_12718,N_11967,N_11643);
nor U12719 (N_12719,N_11345,N_11375);
and U12720 (N_12720,N_11379,N_11301);
xnor U12721 (N_12721,N_11837,N_11903);
or U12722 (N_12722,N_11606,N_11269);
or U12723 (N_12723,N_11773,N_11558);
nand U12724 (N_12724,N_11699,N_11693);
and U12725 (N_12725,N_11979,N_11494);
and U12726 (N_12726,N_11779,N_11388);
or U12727 (N_12727,N_11295,N_11844);
and U12728 (N_12728,N_11332,N_11267);
nand U12729 (N_12729,N_11317,N_11411);
or U12730 (N_12730,N_11820,N_11488);
nor U12731 (N_12731,N_11923,N_11876);
nor U12732 (N_12732,N_11649,N_11404);
nand U12733 (N_12733,N_11974,N_11985);
and U12734 (N_12734,N_11595,N_11549);
nor U12735 (N_12735,N_11552,N_11393);
or U12736 (N_12736,N_11888,N_11940);
nor U12737 (N_12737,N_11962,N_11571);
nand U12738 (N_12738,N_11870,N_11804);
nand U12739 (N_12739,N_11686,N_11458);
nor U12740 (N_12740,N_11888,N_11949);
xnor U12741 (N_12741,N_11614,N_11689);
and U12742 (N_12742,N_11763,N_11850);
or U12743 (N_12743,N_11815,N_11879);
nor U12744 (N_12744,N_11953,N_11772);
nor U12745 (N_12745,N_11964,N_11679);
nor U12746 (N_12746,N_11336,N_11985);
xnor U12747 (N_12747,N_11870,N_11909);
nor U12748 (N_12748,N_11810,N_11491);
nand U12749 (N_12749,N_11871,N_11890);
nand U12750 (N_12750,N_12403,N_12276);
xor U12751 (N_12751,N_12261,N_12561);
xnor U12752 (N_12752,N_12135,N_12225);
and U12753 (N_12753,N_12603,N_12482);
xnor U12754 (N_12754,N_12450,N_12352);
or U12755 (N_12755,N_12480,N_12004);
or U12756 (N_12756,N_12055,N_12653);
nand U12757 (N_12757,N_12385,N_12686);
nor U12758 (N_12758,N_12436,N_12151);
or U12759 (N_12759,N_12437,N_12623);
nor U12760 (N_12760,N_12066,N_12416);
xnor U12761 (N_12761,N_12470,N_12419);
and U12762 (N_12762,N_12389,N_12089);
xnor U12763 (N_12763,N_12246,N_12645);
xor U12764 (N_12764,N_12071,N_12616);
nand U12765 (N_12765,N_12165,N_12149);
nand U12766 (N_12766,N_12621,N_12119);
xor U12767 (N_12767,N_12493,N_12425);
nand U12768 (N_12768,N_12639,N_12682);
or U12769 (N_12769,N_12001,N_12034);
nor U12770 (N_12770,N_12594,N_12669);
and U12771 (N_12771,N_12449,N_12635);
nand U12772 (N_12772,N_12063,N_12008);
or U12773 (N_12773,N_12665,N_12137);
and U12774 (N_12774,N_12680,N_12115);
nor U12775 (N_12775,N_12729,N_12249);
or U12776 (N_12776,N_12585,N_12534);
xor U12777 (N_12777,N_12117,N_12345);
or U12778 (N_12778,N_12229,N_12703);
or U12779 (N_12779,N_12587,N_12530);
nand U12780 (N_12780,N_12502,N_12606);
nand U12781 (N_12781,N_12576,N_12304);
nand U12782 (N_12782,N_12365,N_12180);
or U12783 (N_12783,N_12218,N_12347);
xor U12784 (N_12784,N_12191,N_12068);
xor U12785 (N_12785,N_12663,N_12633);
and U12786 (N_12786,N_12279,N_12111);
nand U12787 (N_12787,N_12118,N_12146);
nor U12788 (N_12788,N_12013,N_12208);
nand U12789 (N_12789,N_12062,N_12492);
nand U12790 (N_12790,N_12592,N_12746);
nand U12791 (N_12791,N_12473,N_12438);
nor U12792 (N_12792,N_12692,N_12448);
nand U12793 (N_12793,N_12145,N_12679);
and U12794 (N_12794,N_12659,N_12608);
nor U12795 (N_12795,N_12120,N_12409);
or U12796 (N_12796,N_12346,N_12017);
nor U12797 (N_12797,N_12007,N_12735);
xor U12798 (N_12798,N_12718,N_12320);
or U12799 (N_12799,N_12081,N_12490);
or U12800 (N_12800,N_12581,N_12141);
or U12801 (N_12801,N_12460,N_12230);
nor U12802 (N_12802,N_12381,N_12084);
and U12803 (N_12803,N_12205,N_12725);
or U12804 (N_12804,N_12139,N_12029);
and U12805 (N_12805,N_12021,N_12289);
nand U12806 (N_12806,N_12248,N_12016);
or U12807 (N_12807,N_12324,N_12395);
and U12808 (N_12808,N_12393,N_12681);
nor U12809 (N_12809,N_12307,N_12426);
or U12810 (N_12810,N_12267,N_12458);
or U12811 (N_12811,N_12599,N_12006);
xor U12812 (N_12812,N_12337,N_12150);
and U12813 (N_12813,N_12446,N_12714);
xnor U12814 (N_12814,N_12420,N_12424);
nor U12815 (N_12815,N_12356,N_12049);
nor U12816 (N_12816,N_12154,N_12491);
xnor U12817 (N_12817,N_12190,N_12025);
xnor U12818 (N_12818,N_12051,N_12106);
and U12819 (N_12819,N_12100,N_12042);
and U12820 (N_12820,N_12495,N_12577);
xor U12821 (N_12821,N_12690,N_12551);
xnor U12822 (N_12822,N_12309,N_12565);
and U12823 (N_12823,N_12125,N_12711);
xnor U12824 (N_12824,N_12109,N_12739);
xor U12825 (N_12825,N_12262,N_12281);
or U12826 (N_12826,N_12227,N_12173);
nand U12827 (N_12827,N_12092,N_12694);
nor U12828 (N_12828,N_12722,N_12133);
nand U12829 (N_12829,N_12504,N_12521);
and U12830 (N_12830,N_12011,N_12539);
and U12831 (N_12831,N_12039,N_12287);
and U12832 (N_12832,N_12415,N_12434);
nand U12833 (N_12833,N_12743,N_12142);
nor U12834 (N_12834,N_12405,N_12728);
nand U12835 (N_12835,N_12048,N_12310);
nand U12836 (N_12836,N_12043,N_12384);
nand U12837 (N_12837,N_12342,N_12000);
or U12838 (N_12838,N_12536,N_12358);
or U12839 (N_12839,N_12721,N_12411);
xnor U12840 (N_12840,N_12265,N_12073);
nor U12841 (N_12841,N_12077,N_12516);
or U12842 (N_12842,N_12741,N_12651);
and U12843 (N_12843,N_12467,N_12745);
xnor U12844 (N_12844,N_12041,N_12510);
nand U12845 (N_12845,N_12734,N_12367);
nand U12846 (N_12846,N_12010,N_12563);
and U12847 (N_12847,N_12442,N_12642);
xnor U12848 (N_12848,N_12147,N_12598);
nand U12849 (N_12849,N_12252,N_12290);
nor U12850 (N_12850,N_12638,N_12580);
or U12851 (N_12851,N_12589,N_12666);
nand U12852 (N_12852,N_12527,N_12654);
xnor U12853 (N_12853,N_12184,N_12501);
or U12854 (N_12854,N_12479,N_12296);
xor U12855 (N_12855,N_12387,N_12263);
nor U12856 (N_12856,N_12670,N_12541);
nand U12857 (N_12857,N_12543,N_12588);
xor U12858 (N_12858,N_12259,N_12514);
xnor U12859 (N_12859,N_12167,N_12702);
nor U12860 (N_12860,N_12097,N_12206);
or U12861 (N_12861,N_12518,N_12047);
or U12862 (N_12862,N_12056,N_12103);
and U12863 (N_12863,N_12648,N_12338);
and U12864 (N_12864,N_12602,N_12005);
nor U12865 (N_12865,N_12303,N_12275);
nand U12866 (N_12866,N_12212,N_12369);
nand U12867 (N_12867,N_12171,N_12520);
or U12868 (N_12868,N_12020,N_12193);
and U12869 (N_12869,N_12175,N_12571);
and U12870 (N_12870,N_12629,N_12045);
nor U12871 (N_12871,N_12240,N_12114);
xor U12872 (N_12872,N_12363,N_12214);
nand U12873 (N_12873,N_12636,N_12003);
nor U12874 (N_12874,N_12559,N_12698);
and U12875 (N_12875,N_12090,N_12590);
and U12876 (N_12876,N_12209,N_12391);
nor U12877 (N_12877,N_12236,N_12494);
nand U12878 (N_12878,N_12144,N_12583);
nor U12879 (N_12879,N_12412,N_12658);
or U12880 (N_12880,N_12455,N_12254);
and U12881 (N_12881,N_12700,N_12286);
or U12882 (N_12882,N_12153,N_12037);
nor U12883 (N_12883,N_12738,N_12194);
nand U12884 (N_12884,N_12484,N_12328);
nand U12885 (N_12885,N_12497,N_12406);
nor U12886 (N_12886,N_12657,N_12258);
and U12887 (N_12887,N_12186,N_12123);
or U12888 (N_12888,N_12707,N_12339);
or U12889 (N_12889,N_12508,N_12222);
nand U12890 (N_12890,N_12532,N_12523);
nand U12891 (N_12891,N_12321,N_12368);
nand U12892 (N_12892,N_12087,N_12285);
xor U12893 (N_12893,N_12019,N_12121);
nand U12894 (N_12894,N_12675,N_12268);
and U12895 (N_12895,N_12742,N_12529);
or U12896 (N_12896,N_12428,N_12231);
nand U12897 (N_12897,N_12294,N_12127);
xnor U12898 (N_12898,N_12274,N_12535);
nor U12899 (N_12899,N_12512,N_12716);
nor U12900 (N_12900,N_12672,N_12207);
xor U12901 (N_12901,N_12749,N_12649);
nor U12902 (N_12902,N_12288,N_12132);
nor U12903 (N_12903,N_12542,N_12018);
nand U12904 (N_12904,N_12223,N_12628);
xor U12905 (N_12905,N_12065,N_12401);
nand U12906 (N_12906,N_12238,N_12197);
nor U12907 (N_12907,N_12600,N_12509);
or U12908 (N_12908,N_12113,N_12414);
and U12909 (N_12909,N_12015,N_12567);
and U12910 (N_12910,N_12404,N_12457);
xnor U12911 (N_12911,N_12370,N_12101);
or U12912 (N_12912,N_12189,N_12421);
or U12913 (N_12913,N_12334,N_12394);
and U12914 (N_12914,N_12323,N_12713);
nand U12915 (N_12915,N_12605,N_12162);
nand U12916 (N_12916,N_12496,N_12632);
xor U12917 (N_12917,N_12643,N_12574);
xnor U12918 (N_12918,N_12374,N_12641);
nand U12919 (N_12919,N_12256,N_12255);
or U12920 (N_12920,N_12687,N_12456);
and U12921 (N_12921,N_12105,N_12022);
nand U12922 (N_12922,N_12744,N_12388);
and U12923 (N_12923,N_12531,N_12203);
nor U12924 (N_12924,N_12292,N_12736);
nand U12925 (N_12925,N_12366,N_12554);
nor U12926 (N_12926,N_12319,N_12474);
nor U12927 (N_12927,N_12176,N_12283);
xor U12928 (N_12928,N_12245,N_12382);
xnor U12929 (N_12929,N_12177,N_12549);
nor U12930 (N_12930,N_12349,N_12201);
nand U12931 (N_12931,N_12110,N_12232);
xor U12932 (N_12932,N_12607,N_12211);
nand U12933 (N_12933,N_12555,N_12584);
or U12934 (N_12934,N_12044,N_12515);
xnor U12935 (N_12935,N_12652,N_12159);
nor U12936 (N_12936,N_12701,N_12631);
nor U12937 (N_12937,N_12272,N_12586);
nor U12938 (N_12938,N_12647,N_12575);
xnor U12939 (N_12939,N_12213,N_12557);
and U12940 (N_12940,N_12182,N_12688);
xnor U12941 (N_12941,N_12183,N_12336);
nor U12942 (N_12942,N_12174,N_12610);
nand U12943 (N_12943,N_12499,N_12485);
xnor U12944 (N_12944,N_12348,N_12046);
or U12945 (N_12945,N_12312,N_12462);
xnor U12946 (N_12946,N_12335,N_12002);
xnor U12947 (N_12947,N_12095,N_12298);
and U12948 (N_12948,N_12553,N_12390);
xor U12949 (N_12949,N_12085,N_12228);
and U12950 (N_12950,N_12400,N_12126);
nor U12951 (N_12951,N_12295,N_12568);
nor U12952 (N_12952,N_12094,N_12244);
and U12953 (N_12953,N_12566,N_12082);
and U12954 (N_12954,N_12313,N_12724);
nand U12955 (N_12955,N_12656,N_12644);
and U12956 (N_12956,N_12737,N_12273);
nand U12957 (N_12957,N_12548,N_12134);
nor U12958 (N_12958,N_12293,N_12614);
or U12959 (N_12959,N_12234,N_12253);
and U12960 (N_12960,N_12064,N_12699);
nand U12961 (N_12961,N_12591,N_12096);
nand U12962 (N_12962,N_12200,N_12427);
or U12963 (N_12963,N_12612,N_12488);
nor U12964 (N_12964,N_12251,N_12210);
and U12965 (N_12965,N_12706,N_12524);
or U12966 (N_12966,N_12216,N_12302);
nand U12967 (N_12967,N_12300,N_12188);
or U12968 (N_12968,N_12032,N_12650);
or U12969 (N_12969,N_12560,N_12624);
nor U12970 (N_12970,N_12152,N_12379);
nor U12971 (N_12971,N_12318,N_12451);
xnor U12972 (N_12972,N_12486,N_12489);
and U12973 (N_12973,N_12550,N_12471);
and U12974 (N_12974,N_12627,N_12078);
and U12975 (N_12975,N_12195,N_12572);
xor U12976 (N_12976,N_12361,N_12477);
xor U12977 (N_12977,N_12684,N_12333);
and U12978 (N_12978,N_12717,N_12454);
nand U12979 (N_12979,N_12517,N_12564);
and U12980 (N_12980,N_12076,N_12615);
xnor U12981 (N_12981,N_12693,N_12314);
or U12982 (N_12982,N_12012,N_12116);
nor U12983 (N_12983,N_12464,N_12422);
nor U12984 (N_12984,N_12074,N_12060);
nand U12985 (N_12985,N_12140,N_12511);
nor U12986 (N_12986,N_12498,N_12447);
nand U12987 (N_12987,N_12164,N_12556);
xor U12988 (N_12988,N_12468,N_12306);
or U12989 (N_12989,N_12122,N_12239);
nand U12990 (N_12990,N_12423,N_12432);
nor U12991 (N_12991,N_12161,N_12646);
and U12992 (N_12992,N_12500,N_12579);
and U12993 (N_12993,N_12377,N_12311);
nor U12994 (N_12994,N_12102,N_12673);
and U12995 (N_12995,N_12226,N_12397);
nor U12996 (N_12996,N_12067,N_12266);
and U12997 (N_12997,N_12330,N_12430);
nor U12998 (N_12998,N_12676,N_12506);
xor U12999 (N_12999,N_12315,N_12091);
and U13000 (N_13000,N_12655,N_12027);
xor U13001 (N_13001,N_12155,N_12748);
nand U13002 (N_13002,N_12098,N_12476);
xor U13003 (N_13003,N_12630,N_12383);
nor U13004 (N_13004,N_12260,N_12596);
nor U13005 (N_13005,N_12380,N_12291);
nor U13006 (N_13006,N_12083,N_12179);
or U13007 (N_13007,N_12247,N_12689);
and U13008 (N_13008,N_12407,N_12198);
nand U13009 (N_13009,N_12507,N_12278);
and U13010 (N_13010,N_12661,N_12696);
xor U13011 (N_13011,N_12031,N_12505);
or U13012 (N_13012,N_12709,N_12481);
nand U13013 (N_13013,N_12353,N_12086);
xor U13014 (N_13014,N_12220,N_12622);
xnor U13015 (N_13015,N_12376,N_12129);
or U13016 (N_13016,N_12217,N_12710);
nand U13017 (N_13017,N_12625,N_12344);
xor U13018 (N_13018,N_12640,N_12715);
nor U13019 (N_13019,N_12704,N_12440);
nor U13020 (N_13020,N_12157,N_12578);
nor U13021 (N_13021,N_12070,N_12269);
nand U13022 (N_13022,N_12326,N_12611);
xnor U13023 (N_13023,N_12172,N_12727);
nand U13024 (N_13024,N_12595,N_12257);
and U13025 (N_13025,N_12237,N_12163);
xnor U13026 (N_13026,N_12329,N_12634);
and U13027 (N_13027,N_12112,N_12350);
or U13028 (N_13028,N_12340,N_12136);
xnor U13029 (N_13029,N_12343,N_12604);
and U13030 (N_13030,N_12413,N_12726);
xnor U13031 (N_13031,N_12053,N_12429);
nor U13032 (N_13032,N_12683,N_12196);
nor U13033 (N_13033,N_12463,N_12325);
xnor U13034 (N_13034,N_12540,N_12023);
and U13035 (N_13035,N_12459,N_12399);
and U13036 (N_13036,N_12124,N_12372);
xor U13037 (N_13037,N_12204,N_12075);
and U13038 (N_13038,N_12028,N_12143);
nand U13039 (N_13039,N_12264,N_12619);
nor U13040 (N_13040,N_12732,N_12410);
nor U13041 (N_13041,N_12674,N_12322);
nor U13042 (N_13042,N_12277,N_12362);
and U13043 (N_13043,N_12138,N_12280);
xnor U13044 (N_13044,N_12417,N_12316);
or U13045 (N_13045,N_12441,N_12284);
xor U13046 (N_13046,N_12487,N_12371);
or U13047 (N_13047,N_12691,N_12079);
xnor U13048 (N_13048,N_12355,N_12452);
or U13049 (N_13049,N_12351,N_12620);
nor U13050 (N_13050,N_12733,N_12618);
nor U13051 (N_13051,N_12522,N_12192);
or U13052 (N_13052,N_12705,N_12364);
or U13053 (N_13053,N_12398,N_12243);
nor U13054 (N_13054,N_12617,N_12088);
nor U13055 (N_13055,N_12009,N_12545);
nand U13056 (N_13056,N_12219,N_12533);
and U13057 (N_13057,N_12720,N_12059);
and U13058 (N_13058,N_12723,N_12433);
nor U13059 (N_13059,N_12354,N_12202);
xor U13060 (N_13060,N_12026,N_12731);
xor U13061 (N_13061,N_12569,N_12740);
and U13062 (N_13062,N_12626,N_12317);
or U13063 (N_13063,N_12107,N_12478);
or U13064 (N_13064,N_12271,N_12301);
nand U13065 (N_13065,N_12038,N_12169);
or U13066 (N_13066,N_12461,N_12052);
nor U13067 (N_13067,N_12475,N_12695);
or U13068 (N_13068,N_12050,N_12668);
or U13069 (N_13069,N_12308,N_12519);
or U13070 (N_13070,N_12538,N_12408);
or U13071 (N_13071,N_12453,N_12503);
nor U13072 (N_13072,N_12719,N_12678);
nor U13073 (N_13073,N_12187,N_12558);
or U13074 (N_13074,N_12199,N_12221);
nor U13075 (N_13075,N_12667,N_12297);
xnor U13076 (N_13076,N_12360,N_12375);
xnor U13077 (N_13077,N_12697,N_12537);
xor U13078 (N_13078,N_12130,N_12242);
nand U13079 (N_13079,N_12181,N_12662);
and U13080 (N_13080,N_12443,N_12593);
xnor U13081 (N_13081,N_12708,N_12040);
nor U13082 (N_13082,N_12712,N_12158);
xnor U13083 (N_13083,N_12061,N_12677);
nor U13084 (N_13084,N_12185,N_12472);
and U13085 (N_13085,N_12166,N_12250);
nand U13086 (N_13086,N_12373,N_12546);
and U13087 (N_13087,N_12160,N_12058);
nor U13088 (N_13088,N_12386,N_12331);
and U13089 (N_13089,N_12024,N_12270);
xnor U13090 (N_13090,N_12469,N_12525);
nand U13091 (N_13091,N_12104,N_12033);
or U13092 (N_13092,N_12215,N_12392);
xor U13093 (N_13093,N_12402,N_12418);
nand U13094 (N_13094,N_12378,N_12168);
and U13095 (N_13095,N_12233,N_12613);
and U13096 (N_13096,N_12664,N_12072);
nor U13097 (N_13097,N_12547,N_12685);
nor U13098 (N_13098,N_12054,N_12080);
nand U13099 (N_13099,N_12131,N_12466);
or U13100 (N_13100,N_12483,N_12562);
and U13101 (N_13101,N_12570,N_12582);
nor U13102 (N_13102,N_12093,N_12359);
xnor U13103 (N_13103,N_12444,N_12396);
xor U13104 (N_13104,N_12069,N_12445);
and U13105 (N_13105,N_12030,N_12660);
nor U13106 (N_13106,N_12332,N_12439);
nor U13107 (N_13107,N_12148,N_12282);
nor U13108 (N_13108,N_12601,N_12099);
nand U13109 (N_13109,N_12597,N_12357);
nor U13110 (N_13110,N_12465,N_12178);
and U13111 (N_13111,N_12526,N_12637);
nor U13112 (N_13112,N_12435,N_12235);
or U13113 (N_13113,N_12108,N_12671);
and U13114 (N_13114,N_12156,N_12036);
nand U13115 (N_13115,N_12327,N_12528);
or U13116 (N_13116,N_12609,N_12014);
xor U13117 (N_13117,N_12513,N_12544);
nor U13118 (N_13118,N_12747,N_12552);
or U13119 (N_13119,N_12730,N_12341);
nand U13120 (N_13120,N_12170,N_12305);
xor U13121 (N_13121,N_12057,N_12035);
and U13122 (N_13122,N_12224,N_12299);
nor U13123 (N_13123,N_12573,N_12431);
nand U13124 (N_13124,N_12128,N_12241);
xor U13125 (N_13125,N_12471,N_12626);
nor U13126 (N_13126,N_12705,N_12067);
nand U13127 (N_13127,N_12078,N_12468);
nor U13128 (N_13128,N_12003,N_12166);
nand U13129 (N_13129,N_12495,N_12457);
xnor U13130 (N_13130,N_12332,N_12200);
xnor U13131 (N_13131,N_12220,N_12529);
nand U13132 (N_13132,N_12673,N_12403);
and U13133 (N_13133,N_12019,N_12347);
nor U13134 (N_13134,N_12142,N_12078);
or U13135 (N_13135,N_12053,N_12721);
nand U13136 (N_13136,N_12678,N_12601);
or U13137 (N_13137,N_12421,N_12470);
and U13138 (N_13138,N_12502,N_12591);
nand U13139 (N_13139,N_12658,N_12252);
nand U13140 (N_13140,N_12669,N_12734);
xnor U13141 (N_13141,N_12669,N_12562);
nor U13142 (N_13142,N_12210,N_12642);
nand U13143 (N_13143,N_12486,N_12418);
xnor U13144 (N_13144,N_12363,N_12193);
or U13145 (N_13145,N_12139,N_12502);
or U13146 (N_13146,N_12117,N_12629);
nor U13147 (N_13147,N_12650,N_12335);
or U13148 (N_13148,N_12561,N_12258);
xor U13149 (N_13149,N_12131,N_12090);
and U13150 (N_13150,N_12649,N_12706);
and U13151 (N_13151,N_12668,N_12244);
and U13152 (N_13152,N_12142,N_12563);
nand U13153 (N_13153,N_12304,N_12406);
xnor U13154 (N_13154,N_12479,N_12631);
and U13155 (N_13155,N_12675,N_12328);
or U13156 (N_13156,N_12173,N_12580);
nor U13157 (N_13157,N_12554,N_12577);
nand U13158 (N_13158,N_12035,N_12655);
xor U13159 (N_13159,N_12006,N_12493);
and U13160 (N_13160,N_12119,N_12421);
or U13161 (N_13161,N_12316,N_12660);
or U13162 (N_13162,N_12632,N_12659);
or U13163 (N_13163,N_12323,N_12141);
nand U13164 (N_13164,N_12734,N_12389);
or U13165 (N_13165,N_12733,N_12227);
xor U13166 (N_13166,N_12273,N_12494);
or U13167 (N_13167,N_12480,N_12585);
and U13168 (N_13168,N_12655,N_12068);
nor U13169 (N_13169,N_12707,N_12156);
and U13170 (N_13170,N_12087,N_12568);
or U13171 (N_13171,N_12205,N_12050);
or U13172 (N_13172,N_12475,N_12365);
nor U13173 (N_13173,N_12490,N_12061);
and U13174 (N_13174,N_12598,N_12351);
nand U13175 (N_13175,N_12511,N_12255);
and U13176 (N_13176,N_12038,N_12161);
xnor U13177 (N_13177,N_12415,N_12689);
xnor U13178 (N_13178,N_12584,N_12716);
or U13179 (N_13179,N_12726,N_12403);
or U13180 (N_13180,N_12234,N_12368);
nand U13181 (N_13181,N_12205,N_12316);
xor U13182 (N_13182,N_12224,N_12030);
nand U13183 (N_13183,N_12342,N_12488);
or U13184 (N_13184,N_12105,N_12668);
nand U13185 (N_13185,N_12022,N_12728);
nor U13186 (N_13186,N_12005,N_12593);
and U13187 (N_13187,N_12225,N_12632);
nand U13188 (N_13188,N_12339,N_12504);
nor U13189 (N_13189,N_12717,N_12211);
nand U13190 (N_13190,N_12207,N_12708);
nand U13191 (N_13191,N_12059,N_12671);
nand U13192 (N_13192,N_12414,N_12070);
nor U13193 (N_13193,N_12742,N_12119);
and U13194 (N_13194,N_12405,N_12314);
or U13195 (N_13195,N_12468,N_12661);
nor U13196 (N_13196,N_12410,N_12700);
and U13197 (N_13197,N_12335,N_12089);
and U13198 (N_13198,N_12503,N_12122);
and U13199 (N_13199,N_12500,N_12725);
and U13200 (N_13200,N_12670,N_12217);
nand U13201 (N_13201,N_12222,N_12010);
nor U13202 (N_13202,N_12343,N_12656);
or U13203 (N_13203,N_12577,N_12239);
nand U13204 (N_13204,N_12313,N_12456);
xor U13205 (N_13205,N_12723,N_12253);
or U13206 (N_13206,N_12118,N_12651);
nand U13207 (N_13207,N_12507,N_12650);
nor U13208 (N_13208,N_12065,N_12530);
xor U13209 (N_13209,N_12440,N_12191);
nor U13210 (N_13210,N_12664,N_12500);
or U13211 (N_13211,N_12416,N_12662);
and U13212 (N_13212,N_12502,N_12664);
and U13213 (N_13213,N_12421,N_12162);
nor U13214 (N_13214,N_12347,N_12046);
or U13215 (N_13215,N_12351,N_12552);
nor U13216 (N_13216,N_12694,N_12243);
nor U13217 (N_13217,N_12595,N_12179);
and U13218 (N_13218,N_12584,N_12534);
nand U13219 (N_13219,N_12052,N_12391);
or U13220 (N_13220,N_12274,N_12197);
xnor U13221 (N_13221,N_12483,N_12643);
or U13222 (N_13222,N_12346,N_12617);
xnor U13223 (N_13223,N_12627,N_12060);
or U13224 (N_13224,N_12370,N_12640);
or U13225 (N_13225,N_12284,N_12475);
nand U13226 (N_13226,N_12023,N_12057);
nand U13227 (N_13227,N_12635,N_12267);
xnor U13228 (N_13228,N_12050,N_12431);
or U13229 (N_13229,N_12259,N_12282);
and U13230 (N_13230,N_12406,N_12626);
or U13231 (N_13231,N_12681,N_12467);
nand U13232 (N_13232,N_12355,N_12181);
nor U13233 (N_13233,N_12327,N_12053);
nor U13234 (N_13234,N_12210,N_12291);
xnor U13235 (N_13235,N_12726,N_12077);
nor U13236 (N_13236,N_12200,N_12526);
xnor U13237 (N_13237,N_12052,N_12266);
nand U13238 (N_13238,N_12504,N_12700);
and U13239 (N_13239,N_12074,N_12346);
nor U13240 (N_13240,N_12088,N_12241);
and U13241 (N_13241,N_12378,N_12082);
nor U13242 (N_13242,N_12546,N_12562);
xnor U13243 (N_13243,N_12464,N_12358);
and U13244 (N_13244,N_12632,N_12663);
xnor U13245 (N_13245,N_12436,N_12362);
xor U13246 (N_13246,N_12642,N_12566);
nand U13247 (N_13247,N_12257,N_12343);
and U13248 (N_13248,N_12164,N_12551);
and U13249 (N_13249,N_12596,N_12641);
or U13250 (N_13250,N_12513,N_12316);
nor U13251 (N_13251,N_12042,N_12350);
nor U13252 (N_13252,N_12720,N_12625);
or U13253 (N_13253,N_12320,N_12177);
and U13254 (N_13254,N_12483,N_12055);
or U13255 (N_13255,N_12176,N_12071);
xor U13256 (N_13256,N_12199,N_12661);
xnor U13257 (N_13257,N_12307,N_12250);
and U13258 (N_13258,N_12067,N_12392);
xor U13259 (N_13259,N_12516,N_12694);
nand U13260 (N_13260,N_12324,N_12711);
and U13261 (N_13261,N_12612,N_12691);
and U13262 (N_13262,N_12588,N_12655);
nor U13263 (N_13263,N_12737,N_12299);
nand U13264 (N_13264,N_12492,N_12452);
and U13265 (N_13265,N_12653,N_12089);
nand U13266 (N_13266,N_12394,N_12162);
nand U13267 (N_13267,N_12541,N_12249);
or U13268 (N_13268,N_12266,N_12337);
nor U13269 (N_13269,N_12184,N_12380);
or U13270 (N_13270,N_12151,N_12527);
or U13271 (N_13271,N_12681,N_12383);
or U13272 (N_13272,N_12610,N_12136);
nand U13273 (N_13273,N_12225,N_12137);
xnor U13274 (N_13274,N_12274,N_12524);
and U13275 (N_13275,N_12371,N_12130);
and U13276 (N_13276,N_12618,N_12471);
xnor U13277 (N_13277,N_12439,N_12502);
and U13278 (N_13278,N_12203,N_12227);
xor U13279 (N_13279,N_12638,N_12642);
xor U13280 (N_13280,N_12703,N_12171);
nand U13281 (N_13281,N_12729,N_12046);
xor U13282 (N_13282,N_12452,N_12009);
or U13283 (N_13283,N_12120,N_12294);
nand U13284 (N_13284,N_12420,N_12044);
nor U13285 (N_13285,N_12051,N_12357);
or U13286 (N_13286,N_12232,N_12437);
xnor U13287 (N_13287,N_12626,N_12366);
nor U13288 (N_13288,N_12597,N_12132);
nor U13289 (N_13289,N_12691,N_12469);
and U13290 (N_13290,N_12466,N_12043);
nand U13291 (N_13291,N_12454,N_12564);
and U13292 (N_13292,N_12507,N_12377);
nand U13293 (N_13293,N_12748,N_12357);
and U13294 (N_13294,N_12202,N_12429);
nand U13295 (N_13295,N_12011,N_12556);
nor U13296 (N_13296,N_12705,N_12159);
or U13297 (N_13297,N_12441,N_12198);
xor U13298 (N_13298,N_12716,N_12681);
xnor U13299 (N_13299,N_12428,N_12343);
or U13300 (N_13300,N_12487,N_12162);
nor U13301 (N_13301,N_12402,N_12292);
xor U13302 (N_13302,N_12492,N_12691);
and U13303 (N_13303,N_12407,N_12265);
and U13304 (N_13304,N_12654,N_12520);
or U13305 (N_13305,N_12590,N_12254);
and U13306 (N_13306,N_12238,N_12158);
nor U13307 (N_13307,N_12666,N_12084);
xor U13308 (N_13308,N_12391,N_12063);
xnor U13309 (N_13309,N_12651,N_12272);
and U13310 (N_13310,N_12516,N_12052);
and U13311 (N_13311,N_12049,N_12583);
and U13312 (N_13312,N_12212,N_12375);
nand U13313 (N_13313,N_12529,N_12582);
nor U13314 (N_13314,N_12469,N_12583);
and U13315 (N_13315,N_12628,N_12345);
xnor U13316 (N_13316,N_12433,N_12437);
nor U13317 (N_13317,N_12003,N_12157);
xor U13318 (N_13318,N_12153,N_12490);
nand U13319 (N_13319,N_12302,N_12127);
xnor U13320 (N_13320,N_12221,N_12155);
or U13321 (N_13321,N_12101,N_12005);
nand U13322 (N_13322,N_12041,N_12726);
nand U13323 (N_13323,N_12623,N_12661);
nand U13324 (N_13324,N_12723,N_12231);
nor U13325 (N_13325,N_12052,N_12176);
nor U13326 (N_13326,N_12264,N_12140);
nand U13327 (N_13327,N_12275,N_12507);
nor U13328 (N_13328,N_12015,N_12258);
and U13329 (N_13329,N_12618,N_12045);
nand U13330 (N_13330,N_12007,N_12741);
and U13331 (N_13331,N_12343,N_12189);
xor U13332 (N_13332,N_12502,N_12417);
nor U13333 (N_13333,N_12285,N_12256);
or U13334 (N_13334,N_12434,N_12059);
nor U13335 (N_13335,N_12298,N_12328);
and U13336 (N_13336,N_12547,N_12551);
nor U13337 (N_13337,N_12054,N_12341);
nor U13338 (N_13338,N_12108,N_12555);
or U13339 (N_13339,N_12247,N_12678);
nand U13340 (N_13340,N_12291,N_12592);
nor U13341 (N_13341,N_12572,N_12514);
nand U13342 (N_13342,N_12451,N_12565);
xor U13343 (N_13343,N_12474,N_12452);
and U13344 (N_13344,N_12424,N_12672);
and U13345 (N_13345,N_12646,N_12073);
nand U13346 (N_13346,N_12515,N_12065);
nor U13347 (N_13347,N_12077,N_12385);
or U13348 (N_13348,N_12541,N_12489);
nor U13349 (N_13349,N_12523,N_12396);
nand U13350 (N_13350,N_12309,N_12435);
nand U13351 (N_13351,N_12510,N_12115);
xor U13352 (N_13352,N_12717,N_12440);
nand U13353 (N_13353,N_12312,N_12010);
xor U13354 (N_13354,N_12327,N_12123);
xnor U13355 (N_13355,N_12620,N_12454);
nand U13356 (N_13356,N_12694,N_12311);
or U13357 (N_13357,N_12326,N_12030);
or U13358 (N_13358,N_12203,N_12142);
nor U13359 (N_13359,N_12662,N_12608);
nor U13360 (N_13360,N_12545,N_12219);
nor U13361 (N_13361,N_12696,N_12241);
and U13362 (N_13362,N_12214,N_12178);
and U13363 (N_13363,N_12710,N_12628);
nor U13364 (N_13364,N_12082,N_12572);
and U13365 (N_13365,N_12647,N_12388);
and U13366 (N_13366,N_12060,N_12016);
or U13367 (N_13367,N_12002,N_12221);
xnor U13368 (N_13368,N_12633,N_12248);
or U13369 (N_13369,N_12400,N_12669);
nand U13370 (N_13370,N_12082,N_12007);
nand U13371 (N_13371,N_12183,N_12295);
nor U13372 (N_13372,N_12385,N_12078);
nand U13373 (N_13373,N_12297,N_12519);
xnor U13374 (N_13374,N_12561,N_12309);
or U13375 (N_13375,N_12714,N_12272);
nor U13376 (N_13376,N_12167,N_12178);
or U13377 (N_13377,N_12018,N_12078);
xnor U13378 (N_13378,N_12330,N_12246);
or U13379 (N_13379,N_12158,N_12258);
or U13380 (N_13380,N_12268,N_12094);
nor U13381 (N_13381,N_12508,N_12259);
nand U13382 (N_13382,N_12016,N_12114);
or U13383 (N_13383,N_12217,N_12157);
nand U13384 (N_13384,N_12221,N_12266);
nor U13385 (N_13385,N_12073,N_12557);
and U13386 (N_13386,N_12013,N_12447);
xnor U13387 (N_13387,N_12238,N_12598);
nand U13388 (N_13388,N_12416,N_12299);
nand U13389 (N_13389,N_12509,N_12063);
xnor U13390 (N_13390,N_12525,N_12343);
nor U13391 (N_13391,N_12523,N_12550);
and U13392 (N_13392,N_12724,N_12298);
xor U13393 (N_13393,N_12653,N_12294);
and U13394 (N_13394,N_12097,N_12238);
xnor U13395 (N_13395,N_12582,N_12641);
and U13396 (N_13396,N_12449,N_12219);
nand U13397 (N_13397,N_12321,N_12293);
nor U13398 (N_13398,N_12618,N_12403);
nand U13399 (N_13399,N_12019,N_12233);
or U13400 (N_13400,N_12554,N_12519);
nor U13401 (N_13401,N_12058,N_12122);
or U13402 (N_13402,N_12365,N_12680);
nor U13403 (N_13403,N_12577,N_12094);
and U13404 (N_13404,N_12582,N_12630);
and U13405 (N_13405,N_12198,N_12458);
nor U13406 (N_13406,N_12475,N_12348);
nand U13407 (N_13407,N_12381,N_12354);
or U13408 (N_13408,N_12728,N_12440);
xor U13409 (N_13409,N_12311,N_12339);
and U13410 (N_13410,N_12641,N_12480);
nor U13411 (N_13411,N_12548,N_12528);
or U13412 (N_13412,N_12699,N_12546);
and U13413 (N_13413,N_12180,N_12736);
nor U13414 (N_13414,N_12168,N_12114);
or U13415 (N_13415,N_12637,N_12431);
nand U13416 (N_13416,N_12641,N_12278);
nor U13417 (N_13417,N_12725,N_12131);
nor U13418 (N_13418,N_12139,N_12287);
and U13419 (N_13419,N_12634,N_12457);
nand U13420 (N_13420,N_12214,N_12398);
xor U13421 (N_13421,N_12155,N_12269);
or U13422 (N_13422,N_12637,N_12661);
nor U13423 (N_13423,N_12152,N_12220);
nand U13424 (N_13424,N_12182,N_12080);
xnor U13425 (N_13425,N_12324,N_12114);
nand U13426 (N_13426,N_12549,N_12474);
xor U13427 (N_13427,N_12266,N_12681);
nand U13428 (N_13428,N_12128,N_12270);
xnor U13429 (N_13429,N_12071,N_12235);
nor U13430 (N_13430,N_12049,N_12693);
nand U13431 (N_13431,N_12527,N_12573);
or U13432 (N_13432,N_12360,N_12461);
xor U13433 (N_13433,N_12483,N_12695);
and U13434 (N_13434,N_12157,N_12222);
and U13435 (N_13435,N_12189,N_12176);
nor U13436 (N_13436,N_12532,N_12268);
and U13437 (N_13437,N_12597,N_12683);
or U13438 (N_13438,N_12499,N_12231);
or U13439 (N_13439,N_12570,N_12748);
and U13440 (N_13440,N_12565,N_12595);
or U13441 (N_13441,N_12496,N_12292);
and U13442 (N_13442,N_12409,N_12651);
xor U13443 (N_13443,N_12085,N_12196);
nor U13444 (N_13444,N_12067,N_12167);
nand U13445 (N_13445,N_12744,N_12052);
and U13446 (N_13446,N_12519,N_12441);
nand U13447 (N_13447,N_12595,N_12320);
or U13448 (N_13448,N_12115,N_12294);
nor U13449 (N_13449,N_12746,N_12153);
or U13450 (N_13450,N_12176,N_12087);
and U13451 (N_13451,N_12238,N_12472);
and U13452 (N_13452,N_12645,N_12230);
or U13453 (N_13453,N_12705,N_12593);
xnor U13454 (N_13454,N_12723,N_12187);
nor U13455 (N_13455,N_12572,N_12538);
nor U13456 (N_13456,N_12671,N_12282);
or U13457 (N_13457,N_12395,N_12483);
nand U13458 (N_13458,N_12229,N_12411);
and U13459 (N_13459,N_12416,N_12449);
nor U13460 (N_13460,N_12695,N_12697);
or U13461 (N_13461,N_12597,N_12581);
or U13462 (N_13462,N_12006,N_12465);
nor U13463 (N_13463,N_12252,N_12708);
or U13464 (N_13464,N_12669,N_12577);
xnor U13465 (N_13465,N_12018,N_12056);
xnor U13466 (N_13466,N_12712,N_12367);
or U13467 (N_13467,N_12226,N_12012);
or U13468 (N_13468,N_12485,N_12654);
or U13469 (N_13469,N_12722,N_12646);
nor U13470 (N_13470,N_12302,N_12662);
nor U13471 (N_13471,N_12624,N_12666);
nor U13472 (N_13472,N_12553,N_12546);
nand U13473 (N_13473,N_12446,N_12201);
nor U13474 (N_13474,N_12673,N_12108);
xor U13475 (N_13475,N_12694,N_12415);
nand U13476 (N_13476,N_12478,N_12419);
xor U13477 (N_13477,N_12541,N_12041);
nor U13478 (N_13478,N_12300,N_12466);
nor U13479 (N_13479,N_12463,N_12243);
and U13480 (N_13480,N_12630,N_12587);
or U13481 (N_13481,N_12375,N_12191);
or U13482 (N_13482,N_12742,N_12530);
or U13483 (N_13483,N_12244,N_12567);
xnor U13484 (N_13484,N_12645,N_12238);
and U13485 (N_13485,N_12405,N_12525);
and U13486 (N_13486,N_12148,N_12149);
nand U13487 (N_13487,N_12472,N_12230);
nand U13488 (N_13488,N_12443,N_12282);
and U13489 (N_13489,N_12398,N_12128);
and U13490 (N_13490,N_12262,N_12601);
nand U13491 (N_13491,N_12746,N_12242);
xnor U13492 (N_13492,N_12583,N_12333);
nand U13493 (N_13493,N_12069,N_12511);
nand U13494 (N_13494,N_12153,N_12024);
or U13495 (N_13495,N_12685,N_12485);
nor U13496 (N_13496,N_12153,N_12657);
xor U13497 (N_13497,N_12100,N_12184);
nand U13498 (N_13498,N_12454,N_12327);
nand U13499 (N_13499,N_12486,N_12653);
or U13500 (N_13500,N_13455,N_12771);
or U13501 (N_13501,N_12961,N_12833);
nor U13502 (N_13502,N_12899,N_13036);
or U13503 (N_13503,N_12984,N_13389);
nor U13504 (N_13504,N_13067,N_12819);
nand U13505 (N_13505,N_13025,N_13121);
xnor U13506 (N_13506,N_13008,N_13382);
xnor U13507 (N_13507,N_13256,N_13410);
xor U13508 (N_13508,N_12886,N_12891);
or U13509 (N_13509,N_13004,N_13139);
nor U13510 (N_13510,N_13064,N_13391);
and U13511 (N_13511,N_13229,N_13166);
or U13512 (N_13512,N_12755,N_12832);
and U13513 (N_13513,N_13110,N_12820);
and U13514 (N_13514,N_13078,N_13251);
xor U13515 (N_13515,N_13173,N_12841);
xor U13516 (N_13516,N_13109,N_12861);
and U13517 (N_13517,N_12962,N_13363);
nor U13518 (N_13518,N_13050,N_12940);
xnor U13519 (N_13519,N_13113,N_12999);
and U13520 (N_13520,N_12966,N_13326);
nor U13521 (N_13521,N_12969,N_12894);
or U13522 (N_13522,N_13108,N_13432);
nor U13523 (N_13523,N_13292,N_12917);
and U13524 (N_13524,N_13190,N_12920);
nand U13525 (N_13525,N_13453,N_13320);
or U13526 (N_13526,N_12773,N_13131);
xnor U13527 (N_13527,N_13269,N_12968);
xnor U13528 (N_13528,N_13007,N_13200);
and U13529 (N_13529,N_13300,N_13371);
nand U13530 (N_13530,N_13026,N_12928);
and U13531 (N_13531,N_13181,N_13101);
or U13532 (N_13532,N_12864,N_13234);
xor U13533 (N_13533,N_13017,N_13021);
or U13534 (N_13534,N_13446,N_12827);
nor U13535 (N_13535,N_12812,N_13277);
nor U13536 (N_13536,N_13381,N_12798);
or U13537 (N_13537,N_13442,N_12845);
or U13538 (N_13538,N_12925,N_13295);
or U13539 (N_13539,N_13048,N_13095);
xnor U13540 (N_13540,N_13129,N_13408);
nor U13541 (N_13541,N_13270,N_12912);
xnor U13542 (N_13542,N_13069,N_12880);
nand U13543 (N_13543,N_12837,N_13312);
or U13544 (N_13544,N_13288,N_13143);
or U13545 (N_13545,N_13049,N_12958);
xnor U13546 (N_13546,N_12835,N_13032);
and U13547 (N_13547,N_13000,N_13339);
or U13548 (N_13548,N_13237,N_13020);
nand U13549 (N_13549,N_13354,N_12865);
and U13550 (N_13550,N_13412,N_12764);
xor U13551 (N_13551,N_13448,N_13016);
and U13552 (N_13552,N_13289,N_12751);
nor U13553 (N_13553,N_13028,N_12997);
nand U13554 (N_13554,N_12873,N_13182);
and U13555 (N_13555,N_13411,N_12821);
and U13556 (N_13556,N_13247,N_12916);
or U13557 (N_13557,N_12898,N_13039);
or U13558 (N_13558,N_12776,N_13183);
nor U13559 (N_13559,N_13169,N_12998);
or U13560 (N_13560,N_12838,N_13188);
nand U13561 (N_13561,N_13255,N_13174);
nand U13562 (N_13562,N_13468,N_12807);
or U13563 (N_13563,N_13119,N_12879);
nand U13564 (N_13564,N_13340,N_13218);
nor U13565 (N_13565,N_13073,N_13350);
and U13566 (N_13566,N_13486,N_13490);
and U13567 (N_13567,N_13465,N_13332);
nand U13568 (N_13568,N_12889,N_12933);
and U13569 (N_13569,N_13060,N_13158);
or U13570 (N_13570,N_13435,N_13123);
or U13571 (N_13571,N_13226,N_13231);
nor U13572 (N_13572,N_12834,N_13195);
xnor U13573 (N_13573,N_12926,N_13212);
nor U13574 (N_13574,N_12923,N_13063);
and U13575 (N_13575,N_12825,N_13290);
nor U13576 (N_13576,N_13429,N_13407);
and U13577 (N_13577,N_12911,N_12974);
nor U13578 (N_13578,N_13058,N_12803);
xnor U13579 (N_13579,N_13168,N_13047);
and U13580 (N_13580,N_12823,N_13274);
xnor U13581 (N_13581,N_12766,N_12976);
nor U13582 (N_13582,N_13244,N_13437);
or U13583 (N_13583,N_13140,N_12818);
and U13584 (N_13584,N_13092,N_12982);
and U13585 (N_13585,N_12794,N_13003);
and U13586 (N_13586,N_12822,N_12765);
or U13587 (N_13587,N_12900,N_13287);
xor U13588 (N_13588,N_13071,N_12789);
or U13589 (N_13589,N_13464,N_12762);
nor U13590 (N_13590,N_12876,N_13471);
and U13591 (N_13591,N_13070,N_13431);
xnor U13592 (N_13592,N_12759,N_13379);
nor U13593 (N_13593,N_13308,N_12957);
nand U13594 (N_13594,N_13248,N_13100);
or U13595 (N_13595,N_12955,N_13498);
and U13596 (N_13596,N_12948,N_13461);
xor U13597 (N_13597,N_12813,N_13030);
nand U13598 (N_13598,N_13319,N_12839);
nand U13599 (N_13599,N_12842,N_12878);
nor U13600 (N_13600,N_13154,N_13337);
and U13601 (N_13601,N_13355,N_13359);
and U13602 (N_13602,N_13044,N_13238);
xor U13603 (N_13603,N_13357,N_13424);
and U13604 (N_13604,N_13336,N_12768);
xnor U13605 (N_13605,N_12913,N_13368);
nor U13606 (N_13606,N_13157,N_12932);
or U13607 (N_13607,N_13062,N_13367);
xor U13608 (N_13608,N_13488,N_12866);
xor U13609 (N_13609,N_13045,N_13115);
xor U13610 (N_13610,N_13040,N_12977);
or U13611 (N_13611,N_13055,N_12885);
or U13612 (N_13612,N_12824,N_13365);
or U13613 (N_13613,N_13019,N_12910);
and U13614 (N_13614,N_13481,N_13005);
nand U13615 (N_13615,N_13074,N_13191);
xor U13616 (N_13616,N_13315,N_13083);
and U13617 (N_13617,N_12863,N_13006);
nand U13618 (N_13618,N_12929,N_13388);
nand U13619 (N_13619,N_12817,N_13478);
or U13620 (N_13620,N_12901,N_12849);
nor U13621 (N_13621,N_13086,N_13459);
and U13622 (N_13622,N_12978,N_12882);
nor U13623 (N_13623,N_13399,N_12987);
xnor U13624 (N_13624,N_13227,N_12959);
nor U13625 (N_13625,N_13241,N_13002);
and U13626 (N_13626,N_12934,N_13102);
nor U13627 (N_13627,N_12874,N_13324);
nand U13628 (N_13628,N_13103,N_13395);
and U13629 (N_13629,N_12906,N_13059);
nor U13630 (N_13630,N_13066,N_13273);
nand U13631 (N_13631,N_12964,N_13243);
xor U13632 (N_13632,N_12951,N_13202);
xor U13633 (N_13633,N_13106,N_13076);
nor U13634 (N_13634,N_12903,N_13136);
xor U13635 (N_13635,N_13334,N_13392);
nor U13636 (N_13636,N_13088,N_12947);
nor U13637 (N_13637,N_13281,N_13299);
and U13638 (N_13638,N_13305,N_13322);
and U13639 (N_13639,N_12750,N_13348);
and U13640 (N_13640,N_13201,N_12809);
nand U13641 (N_13641,N_13239,N_12854);
and U13642 (N_13642,N_13477,N_13219);
nor U13643 (N_13643,N_13484,N_13138);
xor U13644 (N_13644,N_12868,N_13254);
xor U13645 (N_13645,N_13462,N_12888);
nor U13646 (N_13646,N_13483,N_12884);
xor U13647 (N_13647,N_12902,N_13268);
nand U13648 (N_13648,N_13165,N_13061);
nor U13649 (N_13649,N_12780,N_13469);
xnor U13650 (N_13650,N_13031,N_13333);
and U13651 (N_13651,N_13041,N_13375);
and U13652 (N_13652,N_12796,N_12972);
nor U13653 (N_13653,N_12938,N_13180);
or U13654 (N_13654,N_13027,N_13185);
nor U13655 (N_13655,N_13034,N_13015);
nand U13656 (N_13656,N_12829,N_13485);
nand U13657 (N_13657,N_12853,N_12857);
or U13658 (N_13658,N_13346,N_13010);
nand U13659 (N_13659,N_13151,N_12952);
nor U13660 (N_13660,N_12814,N_13208);
or U13661 (N_13661,N_13250,N_12760);
nand U13662 (N_13662,N_12956,N_13366);
and U13663 (N_13663,N_12935,N_12785);
xnor U13664 (N_13664,N_12790,N_12808);
or U13665 (N_13665,N_13114,N_13489);
or U13666 (N_13666,N_12752,N_13072);
xnor U13667 (N_13667,N_13042,N_13438);
or U13668 (N_13668,N_12883,N_13450);
and U13669 (N_13669,N_12828,N_13341);
xor U13670 (N_13670,N_13351,N_13282);
nor U13671 (N_13671,N_13285,N_13096);
and U13672 (N_13672,N_13403,N_12862);
or U13673 (N_13673,N_13497,N_13130);
and U13674 (N_13674,N_13492,N_13172);
xor U13675 (N_13675,N_13137,N_13321);
nor U13676 (N_13676,N_12769,N_12981);
or U13677 (N_13677,N_12836,N_13405);
and U13678 (N_13678,N_12783,N_12777);
xor U13679 (N_13679,N_13311,N_12770);
xor U13680 (N_13680,N_13146,N_12754);
nor U13681 (N_13681,N_13394,N_13402);
xor U13682 (N_13682,N_12846,N_12867);
and U13683 (N_13683,N_13085,N_12847);
xor U13684 (N_13684,N_12816,N_13451);
and U13685 (N_13685,N_13262,N_13235);
nor U13686 (N_13686,N_13033,N_12870);
nor U13687 (N_13687,N_13024,N_13360);
or U13688 (N_13688,N_12985,N_13470);
and U13689 (N_13689,N_12904,N_12996);
and U13690 (N_13690,N_13144,N_13342);
nor U13691 (N_13691,N_12782,N_12810);
xor U13692 (N_13692,N_13203,N_12896);
or U13693 (N_13693,N_12930,N_13252);
and U13694 (N_13694,N_12756,N_13362);
xor U13695 (N_13695,N_12919,N_13303);
and U13696 (N_13696,N_13406,N_13145);
or U13697 (N_13697,N_13038,N_13495);
nand U13698 (N_13698,N_12793,N_12800);
and U13699 (N_13699,N_13105,N_13463);
and U13700 (N_13700,N_13077,N_13344);
or U13701 (N_13701,N_13449,N_12897);
nor U13702 (N_13702,N_12826,N_12954);
xor U13703 (N_13703,N_13271,N_13263);
nor U13704 (N_13704,N_13224,N_13189);
xor U13705 (N_13705,N_13267,N_13482);
nand U13706 (N_13706,N_12772,N_13493);
or U13707 (N_13707,N_13018,N_12909);
or U13708 (N_13708,N_13206,N_12804);
and U13709 (N_13709,N_12843,N_13091);
or U13710 (N_13710,N_13349,N_12973);
or U13711 (N_13711,N_13439,N_13198);
nor U13712 (N_13712,N_13257,N_13358);
or U13713 (N_13713,N_13196,N_13009);
nand U13714 (N_13714,N_13253,N_13258);
nand U13715 (N_13715,N_13184,N_12830);
and U13716 (N_13716,N_13387,N_13283);
nor U13717 (N_13717,N_13499,N_12806);
and U13718 (N_13718,N_13428,N_12775);
nand U13719 (N_13719,N_13338,N_13318);
and U13720 (N_13720,N_13159,N_12767);
xnor U13721 (N_13721,N_13376,N_13310);
or U13722 (N_13722,N_13443,N_12960);
and U13723 (N_13723,N_13156,N_12946);
nand U13724 (N_13724,N_13436,N_12753);
nand U13725 (N_13725,N_13246,N_13452);
xor U13726 (N_13726,N_13401,N_13116);
or U13727 (N_13727,N_13053,N_13421);
xnor U13728 (N_13728,N_13249,N_13161);
nor U13729 (N_13729,N_12914,N_13433);
or U13730 (N_13730,N_12908,N_12949);
nand U13731 (N_13731,N_12792,N_12831);
xor U13732 (N_13732,N_13475,N_13147);
xnor U13733 (N_13733,N_12983,N_13314);
nor U13734 (N_13734,N_13491,N_13094);
and U13735 (N_13735,N_13479,N_13192);
and U13736 (N_13736,N_12915,N_13230);
nand U13737 (N_13737,N_13386,N_13309);
xor U13738 (N_13738,N_13217,N_13013);
nand U13739 (N_13739,N_13221,N_12855);
or U13740 (N_13740,N_13284,N_12774);
or U13741 (N_13741,N_13458,N_13107);
nor U13742 (N_13742,N_13361,N_13396);
and U13743 (N_13743,N_12986,N_13372);
nand U13744 (N_13744,N_13390,N_12895);
or U13745 (N_13745,N_12869,N_13068);
nand U13746 (N_13746,N_13193,N_13135);
nand U13747 (N_13747,N_13126,N_13054);
xor U13748 (N_13748,N_12758,N_13204);
xnor U13749 (N_13749,N_12788,N_13141);
and U13750 (N_13750,N_13306,N_13400);
nor U13751 (N_13751,N_13467,N_13232);
nor U13752 (N_13752,N_13177,N_13425);
nor U13753 (N_13753,N_12802,N_13325);
and U13754 (N_13754,N_13409,N_12995);
or U13755 (N_13755,N_13487,N_12943);
or U13756 (N_13756,N_13280,N_13447);
xor U13757 (N_13757,N_13261,N_12967);
nor U13758 (N_13758,N_13245,N_13082);
and U13759 (N_13759,N_13323,N_13132);
xor U13760 (N_13760,N_12988,N_13415);
nand U13761 (N_13761,N_12763,N_13427);
xor U13762 (N_13762,N_13046,N_13171);
nor U13763 (N_13763,N_13331,N_13293);
nand U13764 (N_13764,N_13111,N_13398);
or U13765 (N_13765,N_12850,N_12872);
nor U13766 (N_13766,N_13220,N_13117);
nor U13767 (N_13767,N_12787,N_13084);
or U13768 (N_13768,N_12941,N_13301);
nand U13769 (N_13769,N_12791,N_13385);
or U13770 (N_13770,N_13223,N_13369);
nor U13771 (N_13771,N_13298,N_13222);
or U13772 (N_13772,N_13089,N_12881);
xnor U13773 (N_13773,N_13418,N_13377);
xnor U13774 (N_13774,N_13148,N_13397);
and U13775 (N_13775,N_12887,N_13302);
xor U13776 (N_13776,N_13120,N_12795);
nor U13777 (N_13777,N_13454,N_12805);
or U13778 (N_13778,N_12875,N_12953);
or U13779 (N_13779,N_13474,N_13090);
and U13780 (N_13780,N_13207,N_13393);
or U13781 (N_13781,N_13374,N_13279);
or U13782 (N_13782,N_12924,N_12781);
nand U13783 (N_13783,N_13133,N_13476);
nand U13784 (N_13784,N_12945,N_13441);
or U13785 (N_13785,N_13012,N_13426);
and U13786 (N_13786,N_13264,N_13414);
or U13787 (N_13787,N_12859,N_13199);
and U13788 (N_13788,N_13416,N_13260);
xor U13789 (N_13789,N_13276,N_12936);
nor U13790 (N_13790,N_12778,N_13297);
and U13791 (N_13791,N_13329,N_13104);
nor U13792 (N_13792,N_13051,N_13215);
xor U13793 (N_13793,N_12971,N_12931);
and U13794 (N_13794,N_12950,N_13125);
or U13795 (N_13795,N_13317,N_13413);
nor U13796 (N_13796,N_12980,N_13343);
nand U13797 (N_13797,N_13286,N_13356);
nand U13798 (N_13798,N_12921,N_13175);
xnor U13799 (N_13799,N_13233,N_13347);
and U13800 (N_13800,N_13327,N_13434);
and U13801 (N_13801,N_13128,N_13170);
and U13802 (N_13802,N_13153,N_12840);
nand U13803 (N_13803,N_13473,N_13466);
nor U13804 (N_13804,N_13057,N_12815);
and U13805 (N_13805,N_12801,N_13328);
nor U13806 (N_13806,N_12922,N_12970);
nand U13807 (N_13807,N_12994,N_12877);
nand U13808 (N_13808,N_12892,N_13162);
and U13809 (N_13809,N_12848,N_13098);
nand U13810 (N_13810,N_12893,N_13014);
or U13811 (N_13811,N_13052,N_13149);
nand U13812 (N_13812,N_13186,N_13445);
or U13813 (N_13813,N_12890,N_13001);
xnor U13814 (N_13814,N_13080,N_12779);
nor U13815 (N_13815,N_13081,N_13210);
nand U13816 (N_13816,N_12989,N_13122);
xor U13817 (N_13817,N_12963,N_13240);
and U13818 (N_13818,N_12965,N_13278);
nor U13819 (N_13819,N_13440,N_13404);
nand U13820 (N_13820,N_13087,N_13093);
or U13821 (N_13821,N_12844,N_13029);
nor U13822 (N_13822,N_12852,N_13420);
or U13823 (N_13823,N_12993,N_13457);
or U13824 (N_13824,N_12907,N_13228);
and U13825 (N_13825,N_12905,N_13127);
nand U13826 (N_13826,N_13211,N_12797);
xnor U13827 (N_13827,N_13307,N_13197);
xnor U13828 (N_13828,N_13294,N_12937);
or U13829 (N_13829,N_13383,N_13496);
or U13830 (N_13830,N_13335,N_13205);
nor U13831 (N_13831,N_13417,N_12860);
nor U13832 (N_13832,N_12871,N_13056);
and U13833 (N_13833,N_12757,N_12944);
or U13834 (N_13834,N_13384,N_12927);
nor U13835 (N_13835,N_13176,N_13134);
xnor U13836 (N_13836,N_13035,N_13022);
or U13837 (N_13837,N_13352,N_12918);
or U13838 (N_13838,N_12811,N_13330);
nor U13839 (N_13839,N_13265,N_13313);
xnor U13840 (N_13840,N_13214,N_13216);
xor U13841 (N_13841,N_13296,N_12858);
and U13842 (N_13842,N_13378,N_13155);
nor U13843 (N_13843,N_13494,N_13075);
xnor U13844 (N_13844,N_13079,N_12856);
nor U13845 (N_13845,N_13179,N_13370);
or U13846 (N_13846,N_13011,N_12990);
nor U13847 (N_13847,N_13419,N_13023);
nor U13848 (N_13848,N_13380,N_13164);
or U13849 (N_13849,N_13422,N_13345);
nand U13850 (N_13850,N_13304,N_13194);
xnor U13851 (N_13851,N_13444,N_13213);
nor U13852 (N_13852,N_12979,N_12992);
xor U13853 (N_13853,N_13037,N_13097);
xnor U13854 (N_13854,N_13150,N_13043);
xnor U13855 (N_13855,N_13364,N_13236);
and U13856 (N_13856,N_13178,N_12942);
or U13857 (N_13857,N_13430,N_12851);
and U13858 (N_13858,N_13456,N_13272);
or U13859 (N_13859,N_13099,N_13266);
nand U13860 (N_13860,N_13187,N_12991);
and U13861 (N_13861,N_13472,N_13160);
or U13862 (N_13862,N_13242,N_13118);
nand U13863 (N_13863,N_13065,N_13112);
or U13864 (N_13864,N_13163,N_13460);
xor U13865 (N_13865,N_13142,N_13353);
and U13866 (N_13866,N_12799,N_13316);
nand U13867 (N_13867,N_13275,N_13225);
or U13868 (N_13868,N_12786,N_13373);
nor U13869 (N_13869,N_13167,N_13152);
nand U13870 (N_13870,N_13480,N_13423);
nand U13871 (N_13871,N_12939,N_13291);
or U13872 (N_13872,N_13259,N_12761);
nor U13873 (N_13873,N_13124,N_12975);
and U13874 (N_13874,N_13209,N_12784);
xor U13875 (N_13875,N_13490,N_13359);
xnor U13876 (N_13876,N_12827,N_13281);
or U13877 (N_13877,N_13051,N_13079);
or U13878 (N_13878,N_13085,N_12775);
and U13879 (N_13879,N_13409,N_13389);
and U13880 (N_13880,N_12965,N_13285);
and U13881 (N_13881,N_12957,N_13364);
xnor U13882 (N_13882,N_13069,N_13317);
nor U13883 (N_13883,N_12934,N_12847);
or U13884 (N_13884,N_13117,N_13142);
nand U13885 (N_13885,N_13322,N_12766);
xnor U13886 (N_13886,N_13071,N_13421);
or U13887 (N_13887,N_13476,N_13471);
xor U13888 (N_13888,N_13400,N_12835);
and U13889 (N_13889,N_12811,N_12830);
or U13890 (N_13890,N_13268,N_13484);
nand U13891 (N_13891,N_13379,N_13284);
nor U13892 (N_13892,N_13028,N_12800);
or U13893 (N_13893,N_13053,N_12790);
xnor U13894 (N_13894,N_12809,N_13097);
or U13895 (N_13895,N_13126,N_12969);
nor U13896 (N_13896,N_13393,N_12759);
xor U13897 (N_13897,N_13215,N_13081);
nor U13898 (N_13898,N_13314,N_13143);
or U13899 (N_13899,N_12892,N_13482);
xnor U13900 (N_13900,N_12897,N_12892);
xor U13901 (N_13901,N_12983,N_13361);
nand U13902 (N_13902,N_13317,N_12781);
and U13903 (N_13903,N_12815,N_12750);
nor U13904 (N_13904,N_13052,N_13224);
nand U13905 (N_13905,N_12831,N_12895);
nand U13906 (N_13906,N_12853,N_12898);
nor U13907 (N_13907,N_13346,N_12818);
nand U13908 (N_13908,N_13197,N_13424);
xor U13909 (N_13909,N_13439,N_13140);
and U13910 (N_13910,N_13067,N_13150);
xnor U13911 (N_13911,N_13002,N_13126);
nand U13912 (N_13912,N_12860,N_13358);
nand U13913 (N_13913,N_12891,N_12853);
nor U13914 (N_13914,N_12982,N_13451);
and U13915 (N_13915,N_13268,N_13137);
xor U13916 (N_13916,N_13369,N_13380);
and U13917 (N_13917,N_13266,N_13265);
nor U13918 (N_13918,N_13199,N_12910);
and U13919 (N_13919,N_13033,N_12807);
and U13920 (N_13920,N_12805,N_13396);
nor U13921 (N_13921,N_12914,N_13083);
and U13922 (N_13922,N_13427,N_13077);
and U13923 (N_13923,N_13377,N_13431);
or U13924 (N_13924,N_13302,N_12845);
nor U13925 (N_13925,N_12963,N_12928);
and U13926 (N_13926,N_12833,N_13102);
nand U13927 (N_13927,N_12910,N_12908);
and U13928 (N_13928,N_12935,N_13199);
or U13929 (N_13929,N_13401,N_13111);
xor U13930 (N_13930,N_13017,N_13435);
and U13931 (N_13931,N_13252,N_13334);
nand U13932 (N_13932,N_12932,N_13295);
nor U13933 (N_13933,N_12791,N_13186);
or U13934 (N_13934,N_13346,N_13466);
xnor U13935 (N_13935,N_13452,N_13090);
nand U13936 (N_13936,N_13016,N_12975);
nor U13937 (N_13937,N_12998,N_12782);
nand U13938 (N_13938,N_13373,N_13197);
and U13939 (N_13939,N_12915,N_12985);
and U13940 (N_13940,N_12893,N_13108);
nor U13941 (N_13941,N_12794,N_13296);
nor U13942 (N_13942,N_12876,N_12925);
xnor U13943 (N_13943,N_13258,N_12885);
or U13944 (N_13944,N_12979,N_13359);
and U13945 (N_13945,N_13371,N_13133);
xnor U13946 (N_13946,N_12950,N_13038);
xnor U13947 (N_13947,N_13380,N_12917);
and U13948 (N_13948,N_12891,N_13416);
xor U13949 (N_13949,N_13097,N_13479);
or U13950 (N_13950,N_13353,N_13413);
xor U13951 (N_13951,N_13084,N_13349);
and U13952 (N_13952,N_13466,N_13099);
or U13953 (N_13953,N_13029,N_12960);
or U13954 (N_13954,N_13025,N_13393);
and U13955 (N_13955,N_13401,N_12969);
or U13956 (N_13956,N_12927,N_12986);
and U13957 (N_13957,N_13335,N_13336);
or U13958 (N_13958,N_13254,N_12914);
nor U13959 (N_13959,N_12983,N_12766);
and U13960 (N_13960,N_12959,N_12926);
or U13961 (N_13961,N_13080,N_13452);
xor U13962 (N_13962,N_12805,N_13460);
nand U13963 (N_13963,N_13381,N_13253);
and U13964 (N_13964,N_13175,N_13337);
or U13965 (N_13965,N_13465,N_13011);
and U13966 (N_13966,N_13358,N_13246);
or U13967 (N_13967,N_13208,N_13243);
and U13968 (N_13968,N_13052,N_13384);
nand U13969 (N_13969,N_13162,N_12820);
nor U13970 (N_13970,N_13082,N_13319);
xnor U13971 (N_13971,N_12874,N_13227);
xor U13972 (N_13972,N_13443,N_12807);
and U13973 (N_13973,N_13143,N_13269);
xor U13974 (N_13974,N_12933,N_13470);
nand U13975 (N_13975,N_12837,N_13081);
nor U13976 (N_13976,N_13154,N_12824);
or U13977 (N_13977,N_12898,N_13079);
or U13978 (N_13978,N_13314,N_13147);
or U13979 (N_13979,N_13406,N_13260);
nor U13980 (N_13980,N_13491,N_13333);
nor U13981 (N_13981,N_12837,N_13278);
or U13982 (N_13982,N_13213,N_12912);
xor U13983 (N_13983,N_13132,N_13137);
nor U13984 (N_13984,N_13164,N_13151);
xnor U13985 (N_13985,N_12938,N_13205);
nand U13986 (N_13986,N_12907,N_12820);
xor U13987 (N_13987,N_13489,N_12763);
nor U13988 (N_13988,N_13495,N_13218);
and U13989 (N_13989,N_13343,N_13497);
or U13990 (N_13990,N_13118,N_13087);
and U13991 (N_13991,N_12835,N_13024);
or U13992 (N_13992,N_13104,N_12952);
nand U13993 (N_13993,N_13391,N_13494);
nand U13994 (N_13994,N_13425,N_12998);
nor U13995 (N_13995,N_13217,N_13283);
or U13996 (N_13996,N_13416,N_13234);
nor U13997 (N_13997,N_13431,N_12846);
nand U13998 (N_13998,N_13216,N_12847);
xnor U13999 (N_13999,N_13436,N_13279);
xnor U14000 (N_14000,N_12814,N_13100);
and U14001 (N_14001,N_13177,N_12799);
and U14002 (N_14002,N_12892,N_13077);
nor U14003 (N_14003,N_13192,N_13115);
and U14004 (N_14004,N_13226,N_12797);
or U14005 (N_14005,N_13336,N_12871);
nor U14006 (N_14006,N_12989,N_13060);
or U14007 (N_14007,N_12790,N_13326);
xor U14008 (N_14008,N_13362,N_13281);
or U14009 (N_14009,N_12944,N_13105);
nand U14010 (N_14010,N_12866,N_12907);
xor U14011 (N_14011,N_12994,N_12940);
and U14012 (N_14012,N_12876,N_13029);
xor U14013 (N_14013,N_13061,N_13413);
nor U14014 (N_14014,N_13215,N_13326);
nand U14015 (N_14015,N_13465,N_12894);
nand U14016 (N_14016,N_12863,N_13382);
and U14017 (N_14017,N_13387,N_13090);
nand U14018 (N_14018,N_13269,N_12972);
or U14019 (N_14019,N_13277,N_13391);
xnor U14020 (N_14020,N_12871,N_13495);
nand U14021 (N_14021,N_12790,N_13195);
xor U14022 (N_14022,N_13135,N_12950);
nor U14023 (N_14023,N_12835,N_13367);
nand U14024 (N_14024,N_13080,N_13005);
xor U14025 (N_14025,N_13393,N_13084);
nand U14026 (N_14026,N_12880,N_13162);
nor U14027 (N_14027,N_12928,N_12977);
and U14028 (N_14028,N_12973,N_12757);
nor U14029 (N_14029,N_12878,N_13408);
nand U14030 (N_14030,N_13198,N_13044);
and U14031 (N_14031,N_12929,N_12976);
or U14032 (N_14032,N_12818,N_13424);
nand U14033 (N_14033,N_13072,N_13134);
nor U14034 (N_14034,N_12879,N_13278);
nand U14035 (N_14035,N_13028,N_13137);
nor U14036 (N_14036,N_12779,N_13098);
nor U14037 (N_14037,N_13057,N_12989);
xor U14038 (N_14038,N_13112,N_13323);
nand U14039 (N_14039,N_13454,N_12829);
or U14040 (N_14040,N_13206,N_13148);
and U14041 (N_14041,N_13138,N_12796);
or U14042 (N_14042,N_13261,N_13098);
nor U14043 (N_14043,N_13443,N_13256);
or U14044 (N_14044,N_12750,N_12951);
nand U14045 (N_14045,N_13152,N_13275);
and U14046 (N_14046,N_13392,N_12858);
and U14047 (N_14047,N_13275,N_12907);
and U14048 (N_14048,N_12981,N_12841);
and U14049 (N_14049,N_13246,N_13216);
xor U14050 (N_14050,N_13347,N_12807);
nor U14051 (N_14051,N_12844,N_13233);
nor U14052 (N_14052,N_13215,N_13166);
and U14053 (N_14053,N_13075,N_12830);
and U14054 (N_14054,N_12779,N_13315);
nand U14055 (N_14055,N_13216,N_13037);
or U14056 (N_14056,N_12861,N_13430);
xor U14057 (N_14057,N_13064,N_13393);
or U14058 (N_14058,N_13434,N_13107);
nand U14059 (N_14059,N_13178,N_12986);
xor U14060 (N_14060,N_13467,N_12869);
nand U14061 (N_14061,N_12890,N_13249);
xor U14062 (N_14062,N_13010,N_13437);
nor U14063 (N_14063,N_13217,N_12799);
nand U14064 (N_14064,N_13446,N_12841);
and U14065 (N_14065,N_12784,N_13095);
xor U14066 (N_14066,N_13064,N_13244);
or U14067 (N_14067,N_13439,N_13152);
nor U14068 (N_14068,N_12900,N_13448);
and U14069 (N_14069,N_13463,N_13288);
nor U14070 (N_14070,N_12998,N_13375);
or U14071 (N_14071,N_13213,N_13336);
or U14072 (N_14072,N_13309,N_13165);
and U14073 (N_14073,N_13264,N_12962);
or U14074 (N_14074,N_12932,N_12802);
nor U14075 (N_14075,N_13214,N_12908);
and U14076 (N_14076,N_12813,N_13126);
nand U14077 (N_14077,N_13253,N_13061);
and U14078 (N_14078,N_13293,N_13268);
xor U14079 (N_14079,N_13459,N_12922);
nor U14080 (N_14080,N_13122,N_13093);
or U14081 (N_14081,N_13236,N_13381);
and U14082 (N_14082,N_13489,N_12804);
nor U14083 (N_14083,N_13145,N_13188);
and U14084 (N_14084,N_13487,N_13470);
xor U14085 (N_14085,N_13362,N_13117);
and U14086 (N_14086,N_13233,N_12998);
nand U14087 (N_14087,N_13209,N_13487);
nor U14088 (N_14088,N_13069,N_13036);
nand U14089 (N_14089,N_13015,N_13448);
and U14090 (N_14090,N_13106,N_12818);
and U14091 (N_14091,N_13333,N_12794);
nand U14092 (N_14092,N_12804,N_13297);
or U14093 (N_14093,N_13012,N_12812);
nand U14094 (N_14094,N_13057,N_13221);
and U14095 (N_14095,N_12970,N_13280);
xnor U14096 (N_14096,N_12810,N_13000);
or U14097 (N_14097,N_12790,N_13051);
and U14098 (N_14098,N_13055,N_13353);
and U14099 (N_14099,N_13372,N_13212);
nor U14100 (N_14100,N_13335,N_13333);
or U14101 (N_14101,N_12850,N_12968);
nor U14102 (N_14102,N_13180,N_13259);
nor U14103 (N_14103,N_13180,N_13170);
nor U14104 (N_14104,N_13229,N_13329);
or U14105 (N_14105,N_13275,N_12784);
or U14106 (N_14106,N_12836,N_12886);
nor U14107 (N_14107,N_12913,N_13348);
and U14108 (N_14108,N_13005,N_13172);
and U14109 (N_14109,N_13463,N_13026);
and U14110 (N_14110,N_12867,N_13154);
nand U14111 (N_14111,N_12762,N_13063);
nand U14112 (N_14112,N_13371,N_13157);
xor U14113 (N_14113,N_13258,N_13483);
xor U14114 (N_14114,N_12947,N_12769);
or U14115 (N_14115,N_12930,N_13023);
nor U14116 (N_14116,N_13109,N_13217);
nor U14117 (N_14117,N_13169,N_13042);
and U14118 (N_14118,N_13424,N_12993);
xnor U14119 (N_14119,N_13057,N_12806);
nor U14120 (N_14120,N_12850,N_13032);
xor U14121 (N_14121,N_12758,N_12974);
and U14122 (N_14122,N_12750,N_13316);
xnor U14123 (N_14123,N_13079,N_13184);
nand U14124 (N_14124,N_13157,N_12752);
nand U14125 (N_14125,N_13396,N_13375);
xor U14126 (N_14126,N_13388,N_12897);
or U14127 (N_14127,N_12796,N_13120);
and U14128 (N_14128,N_12810,N_12936);
nand U14129 (N_14129,N_13037,N_13322);
or U14130 (N_14130,N_13326,N_12938);
xnor U14131 (N_14131,N_13387,N_13405);
nand U14132 (N_14132,N_13120,N_13172);
nor U14133 (N_14133,N_12984,N_12774);
nand U14134 (N_14134,N_12764,N_12886);
and U14135 (N_14135,N_12750,N_12937);
nor U14136 (N_14136,N_13481,N_13459);
and U14137 (N_14137,N_13448,N_13091);
nor U14138 (N_14138,N_13008,N_13207);
xor U14139 (N_14139,N_12981,N_13390);
nand U14140 (N_14140,N_13433,N_12919);
nand U14141 (N_14141,N_13267,N_12843);
and U14142 (N_14142,N_13364,N_13102);
or U14143 (N_14143,N_13369,N_13289);
nand U14144 (N_14144,N_13242,N_13413);
or U14145 (N_14145,N_13369,N_13165);
nor U14146 (N_14146,N_12761,N_12808);
xnor U14147 (N_14147,N_13097,N_12964);
nand U14148 (N_14148,N_13025,N_12892);
and U14149 (N_14149,N_12921,N_13201);
or U14150 (N_14150,N_13067,N_13262);
nor U14151 (N_14151,N_12780,N_12901);
nand U14152 (N_14152,N_13091,N_12892);
and U14153 (N_14153,N_12973,N_13015);
nand U14154 (N_14154,N_13160,N_13042);
or U14155 (N_14155,N_13147,N_13295);
nand U14156 (N_14156,N_12856,N_13496);
and U14157 (N_14157,N_12991,N_12949);
and U14158 (N_14158,N_13019,N_13034);
nand U14159 (N_14159,N_13345,N_13418);
xor U14160 (N_14160,N_13480,N_13159);
xnor U14161 (N_14161,N_13483,N_12842);
nor U14162 (N_14162,N_12816,N_12823);
xnor U14163 (N_14163,N_13342,N_13023);
and U14164 (N_14164,N_12898,N_13385);
or U14165 (N_14165,N_12942,N_13438);
nand U14166 (N_14166,N_13400,N_13459);
and U14167 (N_14167,N_12790,N_13330);
or U14168 (N_14168,N_13311,N_13408);
nand U14169 (N_14169,N_13241,N_12804);
nor U14170 (N_14170,N_13329,N_12919);
nand U14171 (N_14171,N_13297,N_13094);
and U14172 (N_14172,N_13261,N_13143);
nand U14173 (N_14173,N_12997,N_13260);
nor U14174 (N_14174,N_12784,N_12998);
nor U14175 (N_14175,N_13469,N_13256);
xnor U14176 (N_14176,N_13286,N_13433);
and U14177 (N_14177,N_13489,N_12836);
nand U14178 (N_14178,N_13292,N_13207);
or U14179 (N_14179,N_12930,N_13092);
or U14180 (N_14180,N_13340,N_13184);
nand U14181 (N_14181,N_13492,N_13431);
nor U14182 (N_14182,N_13396,N_12929);
or U14183 (N_14183,N_13030,N_13448);
or U14184 (N_14184,N_12783,N_13245);
nand U14185 (N_14185,N_12867,N_13264);
or U14186 (N_14186,N_13147,N_13108);
nand U14187 (N_14187,N_13105,N_13070);
or U14188 (N_14188,N_13145,N_13286);
or U14189 (N_14189,N_12953,N_13030);
nor U14190 (N_14190,N_12764,N_12994);
nand U14191 (N_14191,N_13067,N_12750);
and U14192 (N_14192,N_12912,N_13225);
nand U14193 (N_14193,N_12975,N_13257);
nand U14194 (N_14194,N_13455,N_13076);
and U14195 (N_14195,N_13323,N_13347);
nand U14196 (N_14196,N_13053,N_13475);
or U14197 (N_14197,N_13316,N_13394);
and U14198 (N_14198,N_13136,N_12833);
nand U14199 (N_14199,N_13126,N_13105);
xor U14200 (N_14200,N_13383,N_13381);
xor U14201 (N_14201,N_13041,N_13497);
or U14202 (N_14202,N_12787,N_12805);
nand U14203 (N_14203,N_13123,N_13430);
and U14204 (N_14204,N_13376,N_12966);
nor U14205 (N_14205,N_12800,N_13075);
xnor U14206 (N_14206,N_12945,N_12981);
nor U14207 (N_14207,N_13153,N_13007);
or U14208 (N_14208,N_13336,N_12949);
and U14209 (N_14209,N_12832,N_13439);
and U14210 (N_14210,N_12972,N_12756);
nor U14211 (N_14211,N_13021,N_13401);
or U14212 (N_14212,N_13407,N_13496);
or U14213 (N_14213,N_12898,N_13377);
or U14214 (N_14214,N_13398,N_13284);
nor U14215 (N_14215,N_13431,N_12905);
nor U14216 (N_14216,N_12974,N_12919);
and U14217 (N_14217,N_13307,N_13441);
xnor U14218 (N_14218,N_13239,N_12853);
nand U14219 (N_14219,N_13056,N_13346);
xor U14220 (N_14220,N_12826,N_13497);
or U14221 (N_14221,N_12793,N_12753);
or U14222 (N_14222,N_12891,N_13308);
or U14223 (N_14223,N_12918,N_13310);
nand U14224 (N_14224,N_12987,N_12976);
or U14225 (N_14225,N_13364,N_13313);
nand U14226 (N_14226,N_12944,N_12807);
xnor U14227 (N_14227,N_13144,N_13311);
nand U14228 (N_14228,N_13449,N_13228);
or U14229 (N_14229,N_13263,N_12756);
xor U14230 (N_14230,N_12907,N_13117);
xnor U14231 (N_14231,N_13145,N_13425);
or U14232 (N_14232,N_13109,N_12775);
nand U14233 (N_14233,N_13340,N_12816);
nor U14234 (N_14234,N_12809,N_13195);
or U14235 (N_14235,N_13068,N_12875);
and U14236 (N_14236,N_13384,N_13150);
or U14237 (N_14237,N_12902,N_12777);
and U14238 (N_14238,N_13087,N_13302);
nand U14239 (N_14239,N_12886,N_13376);
xor U14240 (N_14240,N_13441,N_13444);
xnor U14241 (N_14241,N_12936,N_12803);
and U14242 (N_14242,N_13245,N_12817);
nor U14243 (N_14243,N_12844,N_12829);
and U14244 (N_14244,N_13453,N_12902);
nor U14245 (N_14245,N_13264,N_12777);
nor U14246 (N_14246,N_13397,N_13460);
and U14247 (N_14247,N_13442,N_12984);
or U14248 (N_14248,N_13215,N_13060);
and U14249 (N_14249,N_13366,N_12795);
xnor U14250 (N_14250,N_14161,N_13980);
nor U14251 (N_14251,N_13872,N_14249);
nor U14252 (N_14252,N_13763,N_14143);
nand U14253 (N_14253,N_14159,N_13533);
or U14254 (N_14254,N_13971,N_13664);
and U14255 (N_14255,N_14202,N_14215);
or U14256 (N_14256,N_13642,N_13524);
nand U14257 (N_14257,N_13956,N_13873);
or U14258 (N_14258,N_13929,N_13516);
nand U14259 (N_14259,N_13688,N_14188);
or U14260 (N_14260,N_13705,N_13736);
nand U14261 (N_14261,N_14244,N_14149);
nor U14262 (N_14262,N_14189,N_14076);
nand U14263 (N_14263,N_13969,N_13834);
xnor U14264 (N_14264,N_13689,N_13882);
and U14265 (N_14265,N_13948,N_13660);
xor U14266 (N_14266,N_13543,N_13846);
xnor U14267 (N_14267,N_13618,N_13845);
nor U14268 (N_14268,N_14198,N_14062);
xor U14269 (N_14269,N_13601,N_13706);
nor U14270 (N_14270,N_13778,N_13953);
nand U14271 (N_14271,N_13596,N_13805);
nor U14272 (N_14272,N_13627,N_14007);
nor U14273 (N_14273,N_13878,N_13780);
or U14274 (N_14274,N_14193,N_13728);
xor U14275 (N_14275,N_13727,N_14068);
or U14276 (N_14276,N_13506,N_13982);
xor U14277 (N_14277,N_13636,N_14024);
or U14278 (N_14278,N_13761,N_14028);
xnor U14279 (N_14279,N_14183,N_14191);
or U14280 (N_14280,N_14069,N_13707);
and U14281 (N_14281,N_13988,N_14242);
nor U14282 (N_14282,N_13735,N_13546);
or U14283 (N_14283,N_14199,N_13509);
xor U14284 (N_14284,N_13749,N_13928);
nand U14285 (N_14285,N_13906,N_13926);
or U14286 (N_14286,N_13607,N_14072);
nor U14287 (N_14287,N_14174,N_13766);
nand U14288 (N_14288,N_13807,N_13698);
and U14289 (N_14289,N_14040,N_14019);
nor U14290 (N_14290,N_14119,N_13526);
xnor U14291 (N_14291,N_13934,N_13922);
and U14292 (N_14292,N_13528,N_13508);
and U14293 (N_14293,N_13574,N_14032);
and U14294 (N_14294,N_13976,N_13904);
nor U14295 (N_14295,N_13853,N_14105);
or U14296 (N_14296,N_13573,N_13768);
nand U14297 (N_14297,N_13898,N_13530);
and U14298 (N_14298,N_13571,N_13876);
nand U14299 (N_14299,N_13624,N_14139);
and U14300 (N_14300,N_13639,N_13667);
and U14301 (N_14301,N_14134,N_13915);
and U14302 (N_14302,N_14085,N_14235);
or U14303 (N_14303,N_14186,N_14027);
or U14304 (N_14304,N_14065,N_13638);
or U14305 (N_14305,N_14165,N_13567);
nand U14306 (N_14306,N_13558,N_13927);
nor U14307 (N_14307,N_13994,N_13998);
nand U14308 (N_14308,N_13850,N_14131);
or U14309 (N_14309,N_13616,N_13540);
nand U14310 (N_14310,N_13593,N_13726);
nand U14311 (N_14311,N_14043,N_13937);
and U14312 (N_14312,N_13968,N_13762);
nor U14313 (N_14313,N_13751,N_13656);
and U14314 (N_14314,N_13787,N_13697);
xnor U14315 (N_14315,N_13868,N_13923);
and U14316 (N_14316,N_13914,N_14035);
xor U14317 (N_14317,N_13774,N_13966);
nor U14318 (N_14318,N_13580,N_13828);
nor U14319 (N_14319,N_14100,N_13967);
nand U14320 (N_14320,N_14126,N_14058);
nand U14321 (N_14321,N_14030,N_13676);
or U14322 (N_14322,N_13916,N_13894);
xnor U14323 (N_14323,N_14155,N_14000);
nor U14324 (N_14324,N_14104,N_13869);
nor U14325 (N_14325,N_14201,N_13946);
xor U14326 (N_14326,N_14051,N_14167);
xnor U14327 (N_14327,N_14010,N_14082);
nor U14328 (N_14328,N_13970,N_13619);
xnor U14329 (N_14329,N_13589,N_13913);
and U14330 (N_14330,N_13901,N_13510);
nor U14331 (N_14331,N_13678,N_13765);
nand U14332 (N_14332,N_13613,N_13769);
or U14333 (N_14333,N_14037,N_13957);
and U14334 (N_14334,N_13572,N_13786);
and U14335 (N_14335,N_14209,N_14148);
and U14336 (N_14336,N_13889,N_13659);
xor U14337 (N_14337,N_14020,N_13757);
nand U14338 (N_14338,N_13544,N_14166);
nand U14339 (N_14339,N_14208,N_13531);
nor U14340 (N_14340,N_13603,N_13663);
nand U14341 (N_14341,N_13704,N_13941);
or U14342 (N_14342,N_13611,N_14224);
or U14343 (N_14343,N_14049,N_14177);
xnor U14344 (N_14344,N_13724,N_14021);
nand U14345 (N_14345,N_13855,N_13770);
and U14346 (N_14346,N_14234,N_14197);
xnor U14347 (N_14347,N_14173,N_14237);
and U14348 (N_14348,N_13793,N_13692);
or U14349 (N_14349,N_13799,N_13826);
nand U14350 (N_14350,N_13819,N_13744);
xnor U14351 (N_14351,N_13553,N_13653);
and U14352 (N_14352,N_13715,N_14026);
nor U14353 (N_14353,N_14182,N_13909);
xor U14354 (N_14354,N_13892,N_14054);
or U14355 (N_14355,N_14239,N_14179);
nor U14356 (N_14356,N_14236,N_14133);
and U14357 (N_14357,N_13885,N_14107);
nor U14358 (N_14358,N_14081,N_14073);
nand U14359 (N_14359,N_13905,N_13746);
xnor U14360 (N_14360,N_13818,N_13903);
and U14361 (N_14361,N_13500,N_13979);
or U14362 (N_14362,N_13599,N_14246);
or U14363 (N_14363,N_13515,N_13794);
nand U14364 (N_14364,N_14078,N_13888);
and U14365 (N_14365,N_14226,N_13628);
or U14366 (N_14366,N_14011,N_13645);
nor U14367 (N_14367,N_13716,N_13925);
and U14368 (N_14368,N_13985,N_13932);
nor U14369 (N_14369,N_14125,N_13641);
and U14370 (N_14370,N_13841,N_13810);
or U14371 (N_14371,N_14036,N_13734);
and U14372 (N_14372,N_13512,N_13760);
nor U14373 (N_14373,N_13521,N_13759);
or U14374 (N_14374,N_14106,N_13576);
and U14375 (N_14375,N_14109,N_13874);
nor U14376 (N_14376,N_13983,N_13550);
or U14377 (N_14377,N_13962,N_14114);
or U14378 (N_14378,N_13804,N_14238);
or U14379 (N_14379,N_13963,N_13847);
nor U14380 (N_14380,N_13696,N_14146);
xor U14381 (N_14381,N_13854,N_13835);
and U14382 (N_14382,N_13960,N_13505);
nor U14383 (N_14383,N_13527,N_13857);
nand U14384 (N_14384,N_13560,N_13816);
nand U14385 (N_14385,N_14016,N_13917);
nand U14386 (N_14386,N_14214,N_13750);
or U14387 (N_14387,N_13949,N_13989);
nand U14388 (N_14388,N_14158,N_13814);
nor U14389 (N_14389,N_14211,N_14074);
nand U14390 (N_14390,N_14175,N_14206);
nor U14391 (N_14391,N_14045,N_14135);
nor U14392 (N_14392,N_13900,N_13785);
nand U14393 (N_14393,N_13635,N_14136);
nand U14394 (N_14394,N_14151,N_13538);
xor U14395 (N_14395,N_13710,N_14142);
nor U14396 (N_14396,N_13658,N_13891);
and U14397 (N_14397,N_13525,N_14110);
nand U14398 (N_14398,N_13858,N_13681);
nand U14399 (N_14399,N_13594,N_13670);
and U14400 (N_14400,N_14034,N_13859);
xor U14401 (N_14401,N_13518,N_13893);
xnor U14402 (N_14402,N_13532,N_13789);
nand U14403 (N_14403,N_14240,N_14123);
and U14404 (N_14404,N_14077,N_13732);
nand U14405 (N_14405,N_14241,N_13931);
and U14406 (N_14406,N_14042,N_13836);
nor U14407 (N_14407,N_13748,N_13779);
xnor U14408 (N_14408,N_13864,N_14171);
xnor U14409 (N_14409,N_13647,N_13803);
xor U14410 (N_14410,N_13943,N_13741);
and U14411 (N_14411,N_13517,N_14200);
xor U14412 (N_14412,N_13733,N_14092);
xnor U14413 (N_14413,N_13686,N_13790);
nand U14414 (N_14414,N_13502,N_13569);
nor U14415 (N_14415,N_13899,N_13783);
xor U14416 (N_14416,N_14229,N_13911);
xor U14417 (N_14417,N_13651,N_13671);
nor U14418 (N_14418,N_13504,N_14163);
and U14419 (N_14419,N_13827,N_13883);
and U14420 (N_14420,N_13597,N_13902);
nand U14421 (N_14421,N_14162,N_13791);
or U14422 (N_14422,N_13687,N_13661);
nand U14423 (N_14423,N_13880,N_14232);
nand U14424 (N_14424,N_13861,N_14031);
nand U14425 (N_14425,N_13867,N_14121);
and U14426 (N_14426,N_14095,N_13919);
nand U14427 (N_14427,N_14122,N_13609);
xor U14428 (N_14428,N_13501,N_13579);
or U14429 (N_14429,N_13650,N_14220);
xnor U14430 (N_14430,N_13514,N_13712);
nand U14431 (N_14431,N_13622,N_14061);
nor U14432 (N_14432,N_13737,N_14101);
and U14433 (N_14433,N_14212,N_13623);
nor U14434 (N_14434,N_14225,N_14086);
nor U14435 (N_14435,N_13592,N_14137);
xnor U14436 (N_14436,N_13672,N_13897);
and U14437 (N_14437,N_13837,N_14227);
nand U14438 (N_14438,N_13981,N_13764);
nand U14439 (N_14439,N_13947,N_13930);
or U14440 (N_14440,N_13582,N_13644);
nor U14441 (N_14441,N_13695,N_14052);
nor U14442 (N_14442,N_14132,N_13964);
or U14443 (N_14443,N_13577,N_14181);
nand U14444 (N_14444,N_13634,N_14172);
or U14445 (N_14445,N_13870,N_13871);
xnor U14446 (N_14446,N_14128,N_13993);
xor U14447 (N_14447,N_14084,N_13598);
nand U14448 (N_14448,N_14001,N_13554);
or U14449 (N_14449,N_13513,N_13851);
and U14450 (N_14450,N_14029,N_13811);
nand U14451 (N_14451,N_13722,N_13523);
xor U14452 (N_14452,N_14117,N_14176);
nand U14453 (N_14453,N_13895,N_13718);
nor U14454 (N_14454,N_13997,N_13723);
xor U14455 (N_14455,N_13954,N_14120);
or U14456 (N_14456,N_13731,N_14097);
nor U14457 (N_14457,N_13729,N_14102);
and U14458 (N_14458,N_13843,N_14184);
xor U14459 (N_14459,N_13797,N_13940);
or U14460 (N_14460,N_13529,N_14127);
nand U14461 (N_14461,N_13605,N_13669);
nor U14462 (N_14462,N_14196,N_13583);
or U14463 (N_14463,N_14023,N_14055);
or U14464 (N_14464,N_14017,N_13564);
xnor U14465 (N_14465,N_13784,N_14025);
or U14466 (N_14466,N_13974,N_13752);
nor U14467 (N_14467,N_14070,N_13632);
xor U14468 (N_14468,N_13747,N_13955);
and U14469 (N_14469,N_13829,N_14195);
xor U14470 (N_14470,N_13581,N_13996);
nand U14471 (N_14471,N_13758,N_14190);
xnor U14472 (N_14472,N_13615,N_13772);
xor U14473 (N_14473,N_13781,N_13547);
nor U14474 (N_14474,N_13792,N_13708);
xor U14475 (N_14475,N_13961,N_13555);
xnor U14476 (N_14476,N_14247,N_13944);
and U14477 (N_14477,N_14060,N_14009);
nor U14478 (N_14478,N_13920,N_14218);
xnor U14479 (N_14479,N_13652,N_13975);
and U14480 (N_14480,N_13884,N_14205);
and U14481 (N_14481,N_14228,N_14090);
nand U14482 (N_14482,N_13701,N_14003);
xnor U14483 (N_14483,N_13725,N_13959);
nor U14484 (N_14484,N_14170,N_13668);
and U14485 (N_14485,N_13511,N_13536);
and U14486 (N_14486,N_14187,N_13693);
xor U14487 (N_14487,N_14079,N_13566);
and U14488 (N_14488,N_13646,N_14147);
and U14489 (N_14489,N_13987,N_13684);
xor U14490 (N_14490,N_14013,N_14207);
nand U14491 (N_14491,N_13753,N_14156);
xnor U14492 (N_14492,N_13865,N_13977);
nand U14493 (N_14493,N_13631,N_13935);
or U14494 (N_14494,N_14064,N_13559);
or U14495 (N_14495,N_13548,N_13742);
and U14496 (N_14496,N_14071,N_14178);
and U14497 (N_14497,N_13682,N_13924);
xnor U14498 (N_14498,N_13626,N_14004);
or U14499 (N_14499,N_13965,N_13995);
nor U14500 (N_14500,N_13938,N_13815);
xnor U14501 (N_14501,N_13612,N_14152);
and U14502 (N_14502,N_13714,N_13796);
or U14503 (N_14503,N_14113,N_13739);
xnor U14504 (N_14504,N_14103,N_14075);
or U14505 (N_14505,N_14180,N_13685);
nand U14506 (N_14506,N_13606,N_13625);
and U14507 (N_14507,N_13823,N_13990);
and U14508 (N_14508,N_13557,N_13675);
nor U14509 (N_14509,N_13640,N_14231);
or U14510 (N_14510,N_13570,N_13662);
nor U14511 (N_14511,N_13575,N_13630);
or U14512 (N_14512,N_14185,N_14112);
nand U14513 (N_14513,N_13522,N_13838);
xor U14514 (N_14514,N_13694,N_13798);
or U14515 (N_14515,N_13812,N_14088);
nor U14516 (N_14516,N_13629,N_14005);
or U14517 (N_14517,N_14059,N_14008);
or U14518 (N_14518,N_13849,N_13621);
nor U14519 (N_14519,N_13825,N_13951);
nand U14520 (N_14520,N_13740,N_13999);
nand U14521 (N_14521,N_13713,N_13939);
or U14522 (N_14522,N_13881,N_13918);
xnor U14523 (N_14523,N_13795,N_13711);
nand U14524 (N_14524,N_13585,N_14083);
nand U14525 (N_14525,N_14015,N_14141);
and U14526 (N_14526,N_13950,N_14157);
nor U14527 (N_14527,N_13691,N_13912);
nand U14528 (N_14528,N_14216,N_13802);
xnor U14529 (N_14529,N_13756,N_14115);
xor U14530 (N_14530,N_14044,N_13649);
nor U14531 (N_14531,N_13972,N_13562);
xnor U14532 (N_14532,N_14038,N_13984);
nand U14533 (N_14533,N_13860,N_13866);
and U14534 (N_14534,N_13936,N_14098);
or U14535 (N_14535,N_13844,N_13657);
nand U14536 (N_14536,N_14046,N_14138);
nand U14537 (N_14537,N_13648,N_13842);
nand U14538 (N_14538,N_13771,N_14140);
xor U14539 (N_14539,N_13637,N_14160);
xnor U14540 (N_14540,N_13703,N_14111);
or U14541 (N_14541,N_13820,N_13863);
or U14542 (N_14542,N_13534,N_14014);
xor U14543 (N_14543,N_13767,N_13776);
nor U14544 (N_14544,N_13745,N_13610);
or U14545 (N_14545,N_13720,N_14144);
xor U14546 (N_14546,N_14217,N_14050);
xor U14547 (N_14547,N_13824,N_13680);
nand U14548 (N_14548,N_14248,N_13683);
xor U14549 (N_14549,N_13856,N_13709);
and U14550 (N_14550,N_13958,N_13578);
or U14551 (N_14551,N_14048,N_13832);
nand U14552 (N_14552,N_13717,N_14006);
xnor U14553 (N_14553,N_13921,N_13831);
or U14554 (N_14554,N_14099,N_13743);
nor U14555 (N_14555,N_14204,N_13690);
nand U14556 (N_14556,N_14153,N_14066);
or U14557 (N_14557,N_14057,N_14047);
xor U14558 (N_14558,N_13933,N_14033);
or U14559 (N_14559,N_13602,N_13537);
or U14560 (N_14560,N_13586,N_13945);
and U14561 (N_14561,N_13549,N_14067);
nor U14562 (N_14562,N_13520,N_14012);
and U14563 (N_14563,N_13801,N_13702);
nor U14564 (N_14564,N_13556,N_13721);
xor U14565 (N_14565,N_13822,N_13617);
and U14566 (N_14566,N_13782,N_13840);
or U14567 (N_14567,N_13839,N_13942);
and U14568 (N_14568,N_13614,N_13852);
xor U14569 (N_14569,N_13907,N_13677);
and U14570 (N_14570,N_13890,N_14118);
or U14571 (N_14571,N_14154,N_13788);
and U14572 (N_14572,N_13674,N_13620);
nor U14573 (N_14573,N_13565,N_13552);
and U14574 (N_14574,N_14223,N_13862);
nor U14575 (N_14575,N_13755,N_14219);
and U14576 (N_14576,N_13666,N_13535);
nor U14577 (N_14577,N_14129,N_14053);
and U14578 (N_14578,N_13886,N_13821);
or U14579 (N_14579,N_14039,N_14002);
xnor U14580 (N_14580,N_13875,N_13633);
nand U14581 (N_14581,N_14221,N_13809);
xor U14582 (N_14582,N_13973,N_13775);
and U14583 (N_14583,N_14108,N_14203);
nor U14584 (N_14584,N_13738,N_14093);
or U14585 (N_14585,N_13673,N_13503);
nor U14586 (N_14586,N_13910,N_13600);
or U14587 (N_14587,N_13654,N_14041);
nand U14588 (N_14588,N_14230,N_13679);
or U14589 (N_14589,N_13800,N_14145);
and U14590 (N_14590,N_14022,N_13991);
and U14591 (N_14591,N_13551,N_13877);
and U14592 (N_14592,N_13595,N_14096);
nor U14593 (N_14593,N_14124,N_14210);
nor U14594 (N_14594,N_13808,N_13908);
xnor U14595 (N_14595,N_13665,N_14194);
nand U14596 (N_14596,N_13700,N_13519);
or U14597 (N_14597,N_13590,N_13608);
and U14598 (N_14598,N_13773,N_14164);
nor U14599 (N_14599,N_13584,N_14245);
or U14600 (N_14600,N_13978,N_13541);
and U14601 (N_14601,N_14018,N_13699);
or U14602 (N_14602,N_13561,N_13539);
xnor U14603 (N_14603,N_13587,N_13887);
xor U14604 (N_14604,N_13655,N_13545);
nand U14605 (N_14605,N_13830,N_13542);
and U14606 (N_14606,N_13813,N_14130);
nor U14607 (N_14607,N_13604,N_13806);
and U14608 (N_14608,N_14150,N_14080);
nor U14609 (N_14609,N_14089,N_13568);
or U14610 (N_14610,N_13563,N_14213);
or U14611 (N_14611,N_13833,N_13777);
nand U14612 (N_14612,N_13588,N_13992);
xnor U14613 (N_14613,N_14063,N_14233);
xnor U14614 (N_14614,N_14222,N_14094);
or U14615 (N_14615,N_13817,N_13730);
nand U14616 (N_14616,N_14192,N_13986);
nor U14617 (N_14617,N_14168,N_13591);
nand U14618 (N_14618,N_14116,N_14056);
or U14619 (N_14619,N_13507,N_13643);
xor U14620 (N_14620,N_14087,N_14091);
nand U14621 (N_14621,N_14169,N_13719);
xnor U14622 (N_14622,N_13879,N_14243);
or U14623 (N_14623,N_13896,N_13952);
nand U14624 (N_14624,N_13754,N_13848);
nor U14625 (N_14625,N_14160,N_14023);
nand U14626 (N_14626,N_14139,N_14227);
and U14627 (N_14627,N_14121,N_13559);
nand U14628 (N_14628,N_14229,N_13940);
or U14629 (N_14629,N_13675,N_14055);
nor U14630 (N_14630,N_13568,N_13592);
and U14631 (N_14631,N_13736,N_14189);
or U14632 (N_14632,N_14162,N_13692);
nor U14633 (N_14633,N_13775,N_13946);
nand U14634 (N_14634,N_13995,N_14032);
nand U14635 (N_14635,N_13968,N_13887);
nand U14636 (N_14636,N_14009,N_13835);
nor U14637 (N_14637,N_14058,N_13942);
nor U14638 (N_14638,N_13799,N_13622);
nand U14639 (N_14639,N_14032,N_14027);
nor U14640 (N_14640,N_13646,N_13622);
xnor U14641 (N_14641,N_13625,N_13958);
and U14642 (N_14642,N_13788,N_13574);
xnor U14643 (N_14643,N_14157,N_14122);
and U14644 (N_14644,N_13822,N_13638);
nand U14645 (N_14645,N_13584,N_13697);
nand U14646 (N_14646,N_14239,N_13528);
nor U14647 (N_14647,N_13976,N_13644);
and U14648 (N_14648,N_13579,N_14192);
and U14649 (N_14649,N_13603,N_14068);
or U14650 (N_14650,N_14137,N_13631);
nand U14651 (N_14651,N_13715,N_13993);
xnor U14652 (N_14652,N_14069,N_13697);
nand U14653 (N_14653,N_13530,N_14161);
xnor U14654 (N_14654,N_13721,N_13952);
nor U14655 (N_14655,N_13737,N_14086);
or U14656 (N_14656,N_13556,N_14242);
or U14657 (N_14657,N_13730,N_13795);
nor U14658 (N_14658,N_13962,N_13981);
nand U14659 (N_14659,N_13980,N_13610);
and U14660 (N_14660,N_14136,N_14222);
nand U14661 (N_14661,N_13646,N_13806);
xnor U14662 (N_14662,N_14074,N_14025);
nand U14663 (N_14663,N_13794,N_13709);
nand U14664 (N_14664,N_13551,N_14228);
nor U14665 (N_14665,N_13601,N_13725);
xnor U14666 (N_14666,N_13922,N_14026);
or U14667 (N_14667,N_13657,N_13601);
xor U14668 (N_14668,N_14116,N_14126);
nand U14669 (N_14669,N_13677,N_13564);
xnor U14670 (N_14670,N_13935,N_14067);
xnor U14671 (N_14671,N_14214,N_14160);
nor U14672 (N_14672,N_13869,N_13777);
xnor U14673 (N_14673,N_13562,N_13786);
or U14674 (N_14674,N_13958,N_14232);
xor U14675 (N_14675,N_13560,N_13799);
nand U14676 (N_14676,N_13632,N_14156);
and U14677 (N_14677,N_13599,N_14190);
nor U14678 (N_14678,N_13568,N_13525);
nand U14679 (N_14679,N_13610,N_14148);
xor U14680 (N_14680,N_13761,N_14188);
nand U14681 (N_14681,N_14108,N_14189);
xnor U14682 (N_14682,N_14015,N_13536);
xor U14683 (N_14683,N_13997,N_13836);
or U14684 (N_14684,N_13964,N_13948);
and U14685 (N_14685,N_13534,N_14035);
xor U14686 (N_14686,N_13687,N_13691);
xor U14687 (N_14687,N_14075,N_13890);
or U14688 (N_14688,N_13650,N_14125);
nand U14689 (N_14689,N_14175,N_13669);
xor U14690 (N_14690,N_14223,N_14185);
nand U14691 (N_14691,N_13646,N_13574);
nor U14692 (N_14692,N_13661,N_13570);
nand U14693 (N_14693,N_13866,N_13848);
nand U14694 (N_14694,N_13542,N_14194);
nor U14695 (N_14695,N_13901,N_14066);
and U14696 (N_14696,N_13662,N_13879);
or U14697 (N_14697,N_13581,N_13979);
nor U14698 (N_14698,N_13802,N_13701);
nor U14699 (N_14699,N_13535,N_14143);
xnor U14700 (N_14700,N_14212,N_13604);
xor U14701 (N_14701,N_14209,N_13520);
xnor U14702 (N_14702,N_13754,N_13527);
or U14703 (N_14703,N_13901,N_13562);
xor U14704 (N_14704,N_13678,N_13944);
or U14705 (N_14705,N_14016,N_14021);
and U14706 (N_14706,N_14043,N_13700);
nor U14707 (N_14707,N_13680,N_13960);
xor U14708 (N_14708,N_14004,N_13961);
or U14709 (N_14709,N_14235,N_13597);
nand U14710 (N_14710,N_13803,N_14040);
nor U14711 (N_14711,N_13918,N_13836);
nand U14712 (N_14712,N_14010,N_13510);
and U14713 (N_14713,N_13685,N_13590);
nand U14714 (N_14714,N_14151,N_14227);
and U14715 (N_14715,N_14158,N_14053);
xnor U14716 (N_14716,N_13964,N_14120);
xor U14717 (N_14717,N_14021,N_14033);
xnor U14718 (N_14718,N_14224,N_13730);
or U14719 (N_14719,N_13718,N_13617);
or U14720 (N_14720,N_13581,N_14100);
and U14721 (N_14721,N_13578,N_14236);
or U14722 (N_14722,N_13891,N_13923);
or U14723 (N_14723,N_13686,N_13982);
xnor U14724 (N_14724,N_14032,N_14199);
or U14725 (N_14725,N_13981,N_13861);
and U14726 (N_14726,N_13844,N_14085);
xnor U14727 (N_14727,N_13694,N_14050);
and U14728 (N_14728,N_13561,N_13713);
xor U14729 (N_14729,N_14128,N_13986);
or U14730 (N_14730,N_13698,N_13845);
or U14731 (N_14731,N_14077,N_14122);
nand U14732 (N_14732,N_13644,N_14129);
or U14733 (N_14733,N_14074,N_14132);
nor U14734 (N_14734,N_13741,N_14249);
nand U14735 (N_14735,N_14171,N_13925);
nand U14736 (N_14736,N_13956,N_13613);
nor U14737 (N_14737,N_13541,N_14098);
and U14738 (N_14738,N_14216,N_13930);
nand U14739 (N_14739,N_13751,N_13577);
nor U14740 (N_14740,N_13850,N_14176);
nor U14741 (N_14741,N_14212,N_14023);
xor U14742 (N_14742,N_13529,N_14247);
and U14743 (N_14743,N_14182,N_13553);
or U14744 (N_14744,N_13862,N_14006);
and U14745 (N_14745,N_13574,N_13912);
and U14746 (N_14746,N_14087,N_14172);
and U14747 (N_14747,N_14191,N_14032);
or U14748 (N_14748,N_13872,N_13568);
nand U14749 (N_14749,N_13872,N_14004);
nor U14750 (N_14750,N_14051,N_13542);
and U14751 (N_14751,N_14177,N_13820);
nor U14752 (N_14752,N_13593,N_14081);
and U14753 (N_14753,N_14046,N_14095);
and U14754 (N_14754,N_13786,N_13861);
nor U14755 (N_14755,N_13866,N_13755);
xor U14756 (N_14756,N_13927,N_13911);
nand U14757 (N_14757,N_14150,N_13745);
or U14758 (N_14758,N_14060,N_13575);
xnor U14759 (N_14759,N_13899,N_13752);
or U14760 (N_14760,N_13691,N_14070);
or U14761 (N_14761,N_13783,N_14136);
nor U14762 (N_14762,N_14076,N_13640);
nand U14763 (N_14763,N_13939,N_14020);
nand U14764 (N_14764,N_14078,N_14204);
and U14765 (N_14765,N_13728,N_13796);
and U14766 (N_14766,N_13877,N_13801);
or U14767 (N_14767,N_14185,N_14102);
and U14768 (N_14768,N_13887,N_13910);
nand U14769 (N_14769,N_14078,N_14036);
or U14770 (N_14770,N_14051,N_13873);
or U14771 (N_14771,N_13786,N_13801);
nor U14772 (N_14772,N_13966,N_14180);
or U14773 (N_14773,N_14184,N_14186);
nor U14774 (N_14774,N_13851,N_13640);
nand U14775 (N_14775,N_13628,N_13817);
and U14776 (N_14776,N_13647,N_13509);
nor U14777 (N_14777,N_14234,N_13896);
xnor U14778 (N_14778,N_13569,N_13907);
nor U14779 (N_14779,N_14104,N_14190);
or U14780 (N_14780,N_13994,N_14047);
nand U14781 (N_14781,N_13790,N_13633);
or U14782 (N_14782,N_13694,N_13864);
nor U14783 (N_14783,N_13685,N_13696);
or U14784 (N_14784,N_13594,N_13687);
or U14785 (N_14785,N_14242,N_13726);
or U14786 (N_14786,N_14132,N_14138);
nor U14787 (N_14787,N_13955,N_13535);
nand U14788 (N_14788,N_13894,N_13600);
or U14789 (N_14789,N_13887,N_13944);
or U14790 (N_14790,N_13846,N_14211);
nor U14791 (N_14791,N_13770,N_13937);
xnor U14792 (N_14792,N_13734,N_13783);
xor U14793 (N_14793,N_13942,N_14092);
and U14794 (N_14794,N_14201,N_14217);
or U14795 (N_14795,N_13663,N_13926);
and U14796 (N_14796,N_14239,N_13719);
nor U14797 (N_14797,N_13601,N_13888);
xor U14798 (N_14798,N_13773,N_14045);
nand U14799 (N_14799,N_13861,N_13523);
nand U14800 (N_14800,N_14017,N_13573);
and U14801 (N_14801,N_14247,N_13804);
and U14802 (N_14802,N_14100,N_14149);
and U14803 (N_14803,N_13849,N_13692);
xnor U14804 (N_14804,N_14242,N_13532);
xnor U14805 (N_14805,N_14005,N_13773);
and U14806 (N_14806,N_13730,N_13527);
nor U14807 (N_14807,N_13563,N_14085);
or U14808 (N_14808,N_14035,N_14169);
nand U14809 (N_14809,N_13510,N_13656);
xnor U14810 (N_14810,N_14173,N_13753);
xor U14811 (N_14811,N_13796,N_13669);
and U14812 (N_14812,N_13983,N_13772);
nand U14813 (N_14813,N_14138,N_13799);
nor U14814 (N_14814,N_14016,N_13781);
or U14815 (N_14815,N_14097,N_14178);
xor U14816 (N_14816,N_14118,N_13569);
nor U14817 (N_14817,N_14185,N_13662);
nand U14818 (N_14818,N_14226,N_13846);
nor U14819 (N_14819,N_14042,N_13529);
xor U14820 (N_14820,N_14143,N_13520);
or U14821 (N_14821,N_14151,N_14074);
nor U14822 (N_14822,N_13510,N_14160);
nor U14823 (N_14823,N_14124,N_13992);
nand U14824 (N_14824,N_13586,N_13940);
and U14825 (N_14825,N_14002,N_13596);
and U14826 (N_14826,N_13831,N_13720);
or U14827 (N_14827,N_13701,N_14128);
nor U14828 (N_14828,N_13863,N_14073);
or U14829 (N_14829,N_13539,N_13715);
nand U14830 (N_14830,N_13657,N_14113);
or U14831 (N_14831,N_13523,N_13536);
nand U14832 (N_14832,N_13915,N_14056);
or U14833 (N_14833,N_13789,N_13730);
nor U14834 (N_14834,N_13638,N_13608);
or U14835 (N_14835,N_13608,N_13974);
xor U14836 (N_14836,N_13887,N_13613);
nor U14837 (N_14837,N_14198,N_14076);
xnor U14838 (N_14838,N_13764,N_13503);
and U14839 (N_14839,N_14213,N_14186);
or U14840 (N_14840,N_13826,N_13771);
or U14841 (N_14841,N_13932,N_13995);
nor U14842 (N_14842,N_13750,N_13890);
xnor U14843 (N_14843,N_14148,N_14197);
and U14844 (N_14844,N_14195,N_13861);
xor U14845 (N_14845,N_14245,N_13507);
or U14846 (N_14846,N_14059,N_14052);
nand U14847 (N_14847,N_13890,N_13507);
and U14848 (N_14848,N_13932,N_13528);
or U14849 (N_14849,N_13943,N_13865);
or U14850 (N_14850,N_14061,N_13599);
nor U14851 (N_14851,N_14121,N_13736);
nor U14852 (N_14852,N_13674,N_13997);
and U14853 (N_14853,N_14228,N_13803);
and U14854 (N_14854,N_14153,N_13802);
and U14855 (N_14855,N_13684,N_14129);
and U14856 (N_14856,N_13624,N_13590);
nand U14857 (N_14857,N_13658,N_13509);
xor U14858 (N_14858,N_14119,N_13999);
or U14859 (N_14859,N_13684,N_13763);
and U14860 (N_14860,N_14137,N_14226);
xor U14861 (N_14861,N_13700,N_13837);
or U14862 (N_14862,N_13738,N_13637);
nand U14863 (N_14863,N_13710,N_13507);
nor U14864 (N_14864,N_13637,N_13566);
or U14865 (N_14865,N_13659,N_14246);
xor U14866 (N_14866,N_14100,N_14160);
and U14867 (N_14867,N_14169,N_13607);
xnor U14868 (N_14868,N_14174,N_13829);
and U14869 (N_14869,N_13896,N_13518);
or U14870 (N_14870,N_14218,N_14118);
nor U14871 (N_14871,N_14099,N_14065);
xnor U14872 (N_14872,N_13784,N_13870);
and U14873 (N_14873,N_13845,N_13860);
nor U14874 (N_14874,N_13632,N_14207);
nor U14875 (N_14875,N_14035,N_13804);
nor U14876 (N_14876,N_13781,N_13640);
and U14877 (N_14877,N_14205,N_13523);
xnor U14878 (N_14878,N_13642,N_13514);
xnor U14879 (N_14879,N_14065,N_14186);
xnor U14880 (N_14880,N_13947,N_13854);
and U14881 (N_14881,N_13848,N_13789);
and U14882 (N_14882,N_13633,N_14094);
or U14883 (N_14883,N_13953,N_14013);
xnor U14884 (N_14884,N_13692,N_14090);
or U14885 (N_14885,N_13618,N_14037);
nor U14886 (N_14886,N_13747,N_14198);
and U14887 (N_14887,N_13698,N_13808);
or U14888 (N_14888,N_14239,N_13832);
and U14889 (N_14889,N_13930,N_14012);
xor U14890 (N_14890,N_14125,N_13960);
xor U14891 (N_14891,N_14218,N_14105);
nand U14892 (N_14892,N_13754,N_13692);
and U14893 (N_14893,N_14024,N_14030);
nand U14894 (N_14894,N_13973,N_13882);
and U14895 (N_14895,N_13720,N_14187);
nor U14896 (N_14896,N_13699,N_13564);
and U14897 (N_14897,N_13601,N_13726);
nand U14898 (N_14898,N_13595,N_14025);
nor U14899 (N_14899,N_13801,N_13594);
nor U14900 (N_14900,N_13952,N_13681);
nand U14901 (N_14901,N_13973,N_13996);
nor U14902 (N_14902,N_13653,N_14177);
and U14903 (N_14903,N_13630,N_14118);
or U14904 (N_14904,N_14034,N_13990);
and U14905 (N_14905,N_14029,N_14140);
xor U14906 (N_14906,N_13683,N_13607);
or U14907 (N_14907,N_14148,N_14046);
or U14908 (N_14908,N_13708,N_14163);
nand U14909 (N_14909,N_14220,N_13744);
nor U14910 (N_14910,N_13861,N_13746);
nor U14911 (N_14911,N_13894,N_14157);
nand U14912 (N_14912,N_13599,N_13777);
and U14913 (N_14913,N_14179,N_14096);
xor U14914 (N_14914,N_13744,N_13816);
nor U14915 (N_14915,N_13649,N_13565);
xor U14916 (N_14916,N_13562,N_13645);
or U14917 (N_14917,N_13613,N_13776);
nor U14918 (N_14918,N_13990,N_14044);
xnor U14919 (N_14919,N_13665,N_13924);
nor U14920 (N_14920,N_13914,N_13972);
and U14921 (N_14921,N_13786,N_13616);
or U14922 (N_14922,N_13778,N_13908);
and U14923 (N_14923,N_13766,N_13888);
or U14924 (N_14924,N_14051,N_14223);
or U14925 (N_14925,N_13529,N_14032);
or U14926 (N_14926,N_14211,N_13746);
nand U14927 (N_14927,N_13885,N_14032);
or U14928 (N_14928,N_14061,N_13767);
nand U14929 (N_14929,N_13691,N_13840);
or U14930 (N_14930,N_13897,N_13695);
nand U14931 (N_14931,N_13828,N_14121);
or U14932 (N_14932,N_13805,N_14191);
or U14933 (N_14933,N_13525,N_13610);
xor U14934 (N_14934,N_14204,N_14016);
nand U14935 (N_14935,N_13781,N_14190);
xnor U14936 (N_14936,N_13756,N_13673);
xnor U14937 (N_14937,N_14178,N_14199);
xnor U14938 (N_14938,N_13955,N_13789);
or U14939 (N_14939,N_13621,N_13625);
nor U14940 (N_14940,N_13983,N_13888);
nand U14941 (N_14941,N_13657,N_13896);
and U14942 (N_14942,N_13611,N_14059);
nand U14943 (N_14943,N_13572,N_13983);
nand U14944 (N_14944,N_13821,N_13631);
nor U14945 (N_14945,N_13837,N_13791);
nand U14946 (N_14946,N_13572,N_13621);
nand U14947 (N_14947,N_13739,N_13925);
and U14948 (N_14948,N_13839,N_14208);
and U14949 (N_14949,N_13939,N_13968);
or U14950 (N_14950,N_14170,N_13537);
and U14951 (N_14951,N_13616,N_13836);
nand U14952 (N_14952,N_13635,N_14017);
nor U14953 (N_14953,N_14170,N_13866);
and U14954 (N_14954,N_14043,N_14226);
or U14955 (N_14955,N_13874,N_13724);
nand U14956 (N_14956,N_13814,N_13590);
xnor U14957 (N_14957,N_13685,N_13781);
nand U14958 (N_14958,N_13864,N_13867);
or U14959 (N_14959,N_13891,N_14016);
nor U14960 (N_14960,N_13825,N_13545);
nand U14961 (N_14961,N_13965,N_14084);
and U14962 (N_14962,N_13745,N_13970);
xnor U14963 (N_14963,N_13659,N_13662);
and U14964 (N_14964,N_13574,N_14205);
nand U14965 (N_14965,N_13731,N_14173);
nand U14966 (N_14966,N_14015,N_13684);
and U14967 (N_14967,N_13820,N_13818);
and U14968 (N_14968,N_13690,N_13919);
or U14969 (N_14969,N_13781,N_13791);
nor U14970 (N_14970,N_13592,N_13574);
xnor U14971 (N_14971,N_13853,N_13929);
and U14972 (N_14972,N_13724,N_13630);
and U14973 (N_14973,N_14053,N_13799);
or U14974 (N_14974,N_13700,N_13713);
nand U14975 (N_14975,N_13681,N_13502);
xnor U14976 (N_14976,N_14162,N_14000);
xor U14977 (N_14977,N_13735,N_13527);
and U14978 (N_14978,N_13510,N_14100);
xnor U14979 (N_14979,N_13570,N_13540);
nor U14980 (N_14980,N_14058,N_13562);
xor U14981 (N_14981,N_14030,N_13700);
and U14982 (N_14982,N_13861,N_14081);
and U14983 (N_14983,N_14175,N_14197);
xor U14984 (N_14984,N_13543,N_14155);
and U14985 (N_14985,N_13747,N_14170);
or U14986 (N_14986,N_13527,N_14120);
or U14987 (N_14987,N_14213,N_13680);
or U14988 (N_14988,N_13651,N_13918);
or U14989 (N_14989,N_13585,N_13762);
nor U14990 (N_14990,N_14021,N_14065);
or U14991 (N_14991,N_13631,N_13998);
xnor U14992 (N_14992,N_14104,N_13725);
xnor U14993 (N_14993,N_13806,N_13523);
and U14994 (N_14994,N_13995,N_13540);
xor U14995 (N_14995,N_14047,N_13969);
and U14996 (N_14996,N_14146,N_14100);
or U14997 (N_14997,N_13876,N_14227);
nor U14998 (N_14998,N_13663,N_13526);
or U14999 (N_14999,N_14230,N_13692);
or UO_0 (O_0,N_14745,N_14705);
or UO_1 (O_1,N_14980,N_14550);
nand UO_2 (O_2,N_14585,N_14554);
or UO_3 (O_3,N_14326,N_14424);
or UO_4 (O_4,N_14532,N_14610);
or UO_5 (O_5,N_14770,N_14301);
nor UO_6 (O_6,N_14358,N_14310);
and UO_7 (O_7,N_14759,N_14841);
and UO_8 (O_8,N_14413,N_14653);
nand UO_9 (O_9,N_14958,N_14643);
nor UO_10 (O_10,N_14697,N_14575);
nand UO_11 (O_11,N_14817,N_14518);
or UO_12 (O_12,N_14461,N_14443);
nand UO_13 (O_13,N_14953,N_14494);
nand UO_14 (O_14,N_14276,N_14539);
nor UO_15 (O_15,N_14719,N_14456);
and UO_16 (O_16,N_14870,N_14606);
xnor UO_17 (O_17,N_14497,N_14440);
xnor UO_18 (O_18,N_14383,N_14996);
xor UO_19 (O_19,N_14305,N_14436);
nand UO_20 (O_20,N_14888,N_14347);
and UO_21 (O_21,N_14355,N_14264);
or UO_22 (O_22,N_14598,N_14277);
xor UO_23 (O_23,N_14956,N_14954);
or UO_24 (O_24,N_14914,N_14921);
nand UO_25 (O_25,N_14803,N_14471);
or UO_26 (O_26,N_14454,N_14685);
or UO_27 (O_27,N_14593,N_14570);
nand UO_28 (O_28,N_14331,N_14903);
nand UO_29 (O_29,N_14569,N_14478);
xor UO_30 (O_30,N_14474,N_14579);
nand UO_31 (O_31,N_14269,N_14935);
and UO_32 (O_32,N_14741,N_14822);
xnor UO_33 (O_33,N_14352,N_14736);
nand UO_34 (O_34,N_14687,N_14945);
and UO_35 (O_35,N_14732,N_14372);
and UO_36 (O_36,N_14889,N_14618);
or UO_37 (O_37,N_14540,N_14441);
and UO_38 (O_38,N_14800,N_14414);
nor UO_39 (O_39,N_14853,N_14769);
nand UO_40 (O_40,N_14711,N_14545);
and UO_41 (O_41,N_14313,N_14785);
and UO_42 (O_42,N_14616,N_14701);
and UO_43 (O_43,N_14819,N_14967);
nor UO_44 (O_44,N_14726,N_14951);
xnor UO_45 (O_45,N_14892,N_14434);
nor UO_46 (O_46,N_14648,N_14321);
nand UO_47 (O_47,N_14897,N_14345);
and UO_48 (O_48,N_14997,N_14353);
and UO_49 (O_49,N_14799,N_14564);
xnor UO_50 (O_50,N_14948,N_14354);
and UO_51 (O_51,N_14964,N_14915);
or UO_52 (O_52,N_14297,N_14872);
xor UO_53 (O_53,N_14343,N_14916);
or UO_54 (O_54,N_14809,N_14303);
xnor UO_55 (O_55,N_14480,N_14720);
nand UO_56 (O_56,N_14279,N_14565);
and UO_57 (O_57,N_14484,N_14315);
nor UO_58 (O_58,N_14563,N_14308);
nand UO_59 (O_59,N_14586,N_14983);
and UO_60 (O_60,N_14510,N_14882);
xnor UO_61 (O_61,N_14342,N_14725);
nor UO_62 (O_62,N_14943,N_14576);
nand UO_63 (O_63,N_14501,N_14735);
xnor UO_64 (O_64,N_14415,N_14560);
nand UO_65 (O_65,N_14363,N_14587);
or UO_66 (O_66,N_14574,N_14638);
nor UO_67 (O_67,N_14737,N_14455);
or UO_68 (O_68,N_14254,N_14934);
nor UO_69 (O_69,N_14581,N_14479);
xor UO_70 (O_70,N_14986,N_14549);
or UO_71 (O_71,N_14761,N_14831);
xor UO_72 (O_72,N_14529,N_14306);
or UO_73 (O_73,N_14790,N_14700);
or UO_74 (O_74,N_14784,N_14664);
and UO_75 (O_75,N_14294,N_14366);
nor UO_76 (O_76,N_14428,N_14546);
or UO_77 (O_77,N_14465,N_14665);
xor UO_78 (O_78,N_14668,N_14690);
nand UO_79 (O_79,N_14292,N_14272);
or UO_80 (O_80,N_14905,N_14670);
nor UO_81 (O_81,N_14318,N_14262);
and UO_82 (O_82,N_14582,N_14509);
xnor UO_83 (O_83,N_14349,N_14982);
xor UO_84 (O_84,N_14333,N_14757);
or UO_85 (O_85,N_14774,N_14512);
or UO_86 (O_86,N_14868,N_14388);
nand UO_87 (O_87,N_14857,N_14703);
or UO_88 (O_88,N_14884,N_14328);
or UO_89 (O_89,N_14802,N_14544);
nand UO_90 (O_90,N_14410,N_14991);
and UO_91 (O_91,N_14714,N_14708);
nor UO_92 (O_92,N_14312,N_14617);
or UO_93 (O_93,N_14583,N_14814);
or UO_94 (O_94,N_14823,N_14612);
nand UO_95 (O_95,N_14722,N_14608);
and UO_96 (O_96,N_14660,N_14758);
and UO_97 (O_97,N_14522,N_14707);
and UO_98 (O_98,N_14968,N_14693);
or UO_99 (O_99,N_14930,N_14886);
nand UO_100 (O_100,N_14675,N_14346);
nor UO_101 (O_101,N_14577,N_14869);
and UO_102 (O_102,N_14742,N_14439);
and UO_103 (O_103,N_14256,N_14846);
and UO_104 (O_104,N_14604,N_14922);
or UO_105 (O_105,N_14397,N_14694);
nand UO_106 (O_106,N_14752,N_14252);
or UO_107 (O_107,N_14537,N_14295);
nor UO_108 (O_108,N_14588,N_14712);
and UO_109 (O_109,N_14258,N_14810);
nand UO_110 (O_110,N_14289,N_14419);
xor UO_111 (O_111,N_14828,N_14282);
xor UO_112 (O_112,N_14332,N_14852);
nand UO_113 (O_113,N_14734,N_14449);
or UO_114 (O_114,N_14382,N_14526);
xnor UO_115 (O_115,N_14939,N_14808);
and UO_116 (O_116,N_14572,N_14796);
xor UO_117 (O_117,N_14629,N_14874);
xor UO_118 (O_118,N_14778,N_14950);
and UO_119 (O_119,N_14265,N_14816);
xor UO_120 (O_120,N_14314,N_14840);
nand UO_121 (O_121,N_14684,N_14866);
nor UO_122 (O_122,N_14843,N_14881);
and UO_123 (O_123,N_14408,N_14597);
nor UO_124 (O_124,N_14985,N_14592);
or UO_125 (O_125,N_14845,N_14891);
nor UO_126 (O_126,N_14847,N_14286);
and UO_127 (O_127,N_14678,N_14350);
xor UO_128 (O_128,N_14826,N_14482);
xor UO_129 (O_129,N_14601,N_14910);
nor UO_130 (O_130,N_14299,N_14362);
or UO_131 (O_131,N_14718,N_14250);
or UO_132 (O_132,N_14955,N_14596);
and UO_133 (O_133,N_14671,N_14261);
nand UO_134 (O_134,N_14864,N_14302);
nand UO_135 (O_135,N_14691,N_14406);
nand UO_136 (O_136,N_14786,N_14669);
or UO_137 (O_137,N_14534,N_14371);
xnor UO_138 (O_138,N_14942,N_14444);
and UO_139 (O_139,N_14491,N_14862);
and UO_140 (O_140,N_14263,N_14339);
nand UO_141 (O_141,N_14733,N_14538);
nor UO_142 (O_142,N_14599,N_14842);
nand UO_143 (O_143,N_14860,N_14435);
or UO_144 (O_144,N_14965,N_14492);
nor UO_145 (O_145,N_14777,N_14476);
nor UO_146 (O_146,N_14381,N_14337);
nor UO_147 (O_147,N_14856,N_14688);
nand UO_148 (O_148,N_14792,N_14837);
or UO_149 (O_149,N_14635,N_14767);
xnor UO_150 (O_150,N_14475,N_14839);
nand UO_151 (O_151,N_14977,N_14630);
nor UO_152 (O_152,N_14829,N_14788);
and UO_153 (O_153,N_14573,N_14438);
or UO_154 (O_154,N_14754,N_14404);
xnor UO_155 (O_155,N_14513,N_14765);
and UO_156 (O_156,N_14972,N_14365);
nand UO_157 (O_157,N_14644,N_14298);
nand UO_158 (O_158,N_14502,N_14871);
nand UO_159 (O_159,N_14291,N_14779);
xnor UO_160 (O_160,N_14485,N_14548);
nor UO_161 (O_161,N_14525,N_14724);
xor UO_162 (O_162,N_14713,N_14403);
nand UO_163 (O_163,N_14755,N_14268);
nor UO_164 (O_164,N_14698,N_14373);
and UO_165 (O_165,N_14894,N_14386);
and UO_166 (O_166,N_14390,N_14919);
and UO_167 (O_167,N_14925,N_14834);
or UO_168 (O_168,N_14949,N_14970);
and UO_169 (O_169,N_14278,N_14812);
or UO_170 (O_170,N_14394,N_14266);
xor UO_171 (O_171,N_14746,N_14999);
nor UO_172 (O_172,N_14821,N_14429);
or UO_173 (O_173,N_14917,N_14280);
and UO_174 (O_174,N_14775,N_14651);
xor UO_175 (O_175,N_14677,N_14738);
and UO_176 (O_176,N_14824,N_14959);
or UO_177 (O_177,N_14259,N_14895);
nor UO_178 (O_178,N_14338,N_14706);
nand UO_179 (O_179,N_14928,N_14483);
and UO_180 (O_180,N_14727,N_14561);
or UO_181 (O_181,N_14452,N_14811);
nand UO_182 (O_182,N_14666,N_14551);
or UO_183 (O_183,N_14993,N_14274);
nor UO_184 (O_184,N_14854,N_14595);
and UO_185 (O_185,N_14432,N_14876);
nand UO_186 (O_186,N_14877,N_14511);
xor UO_187 (O_187,N_14271,N_14374);
nand UO_188 (O_188,N_14680,N_14740);
xor UO_189 (O_189,N_14749,N_14607);
xnor UO_190 (O_190,N_14348,N_14764);
or UO_191 (O_191,N_14334,N_14887);
or UO_192 (O_192,N_14571,N_14743);
nand UO_193 (O_193,N_14251,N_14542);
xnor UO_194 (O_194,N_14378,N_14931);
nor UO_195 (O_195,N_14489,N_14637);
or UO_196 (O_196,N_14625,N_14364);
or UO_197 (O_197,N_14798,N_14920);
or UO_198 (O_198,N_14851,N_14420);
or UO_199 (O_199,N_14830,N_14589);
nand UO_200 (O_200,N_14393,N_14940);
nand UO_201 (O_201,N_14361,N_14640);
nand UO_202 (O_202,N_14418,N_14899);
nand UO_203 (O_203,N_14379,N_14901);
and UO_204 (O_204,N_14890,N_14402);
xor UO_205 (O_205,N_14833,N_14918);
nand UO_206 (O_206,N_14801,N_14609);
nor UO_207 (O_207,N_14753,N_14649);
or UO_208 (O_208,N_14260,N_14807);
or UO_209 (O_209,N_14676,N_14966);
and UO_210 (O_210,N_14605,N_14674);
xnor UO_211 (O_211,N_14624,N_14470);
xor UO_212 (O_212,N_14760,N_14642);
nor UO_213 (O_213,N_14813,N_14836);
nor UO_214 (O_214,N_14686,N_14656);
and UO_215 (O_215,N_14503,N_14750);
nand UO_216 (O_216,N_14530,N_14791);
nor UO_217 (O_217,N_14445,N_14827);
or UO_218 (O_218,N_14531,N_14360);
or UO_219 (O_219,N_14751,N_14661);
and UO_220 (O_220,N_14281,N_14825);
nand UO_221 (O_221,N_14789,N_14627);
xor UO_222 (O_222,N_14771,N_14621);
and UO_223 (O_223,N_14927,N_14508);
nor UO_224 (O_224,N_14387,N_14729);
nand UO_225 (O_225,N_14499,N_14613);
nor UO_226 (O_226,N_14620,N_14699);
nand UO_227 (O_227,N_14963,N_14359);
nand UO_228 (O_228,N_14384,N_14768);
nand UO_229 (O_229,N_14850,N_14893);
or UO_230 (O_230,N_14663,N_14351);
xor UO_231 (O_231,N_14543,N_14748);
nand UO_232 (O_232,N_14401,N_14391);
nand UO_233 (O_233,N_14655,N_14336);
nor UO_234 (O_234,N_14309,N_14427);
nand UO_235 (O_235,N_14527,N_14568);
and UO_236 (O_236,N_14944,N_14960);
or UO_237 (O_237,N_14591,N_14451);
or UO_238 (O_238,N_14523,N_14317);
nor UO_239 (O_239,N_14929,N_14679);
and UO_240 (O_240,N_14602,N_14794);
xor UO_241 (O_241,N_14990,N_14578);
and UO_242 (O_242,N_14488,N_14590);
nor UO_243 (O_243,N_14739,N_14462);
nor UO_244 (O_244,N_14773,N_14396);
nor UO_245 (O_245,N_14975,N_14562);
nand UO_246 (O_246,N_14498,N_14368);
nand UO_247 (O_247,N_14647,N_14936);
nor UO_248 (O_248,N_14976,N_14495);
nand UO_249 (O_249,N_14426,N_14457);
nand UO_250 (O_250,N_14692,N_14375);
xor UO_251 (O_251,N_14673,N_14453);
nand UO_252 (O_252,N_14340,N_14776);
xnor UO_253 (O_253,N_14873,N_14437);
xnor UO_254 (O_254,N_14904,N_14623);
xor UO_255 (O_255,N_14552,N_14952);
nand UO_256 (O_256,N_14710,N_14422);
and UO_257 (O_257,N_14516,N_14376);
or UO_258 (O_258,N_14399,N_14988);
and UO_259 (O_259,N_14311,N_14646);
nand UO_260 (O_260,N_14995,N_14329);
nor UO_261 (O_261,N_14433,N_14556);
nand UO_262 (O_262,N_14356,N_14447);
nand UO_263 (O_263,N_14766,N_14411);
xor UO_264 (O_264,N_14584,N_14377);
and UO_265 (O_265,N_14463,N_14580);
nand UO_266 (O_266,N_14622,N_14533);
nor UO_267 (O_267,N_14412,N_14500);
xnor UO_268 (O_268,N_14324,N_14709);
nand UO_269 (O_269,N_14815,N_14514);
nor UO_270 (O_270,N_14989,N_14744);
xor UO_271 (O_271,N_14645,N_14307);
or UO_272 (O_272,N_14658,N_14566);
xor UO_273 (O_273,N_14619,N_14818);
and UO_274 (O_274,N_14267,N_14902);
or UO_275 (O_275,N_14486,N_14937);
nand UO_276 (O_276,N_14721,N_14938);
xor UO_277 (O_277,N_14528,N_14287);
or UO_278 (O_278,N_14473,N_14797);
nand UO_279 (O_279,N_14878,N_14793);
nand UO_280 (O_280,N_14762,N_14763);
nor UO_281 (O_281,N_14536,N_14662);
xor UO_282 (O_282,N_14981,N_14723);
xor UO_283 (O_283,N_14505,N_14273);
nand UO_284 (O_284,N_14628,N_14861);
nand UO_285 (O_285,N_14865,N_14304);
nand UO_286 (O_286,N_14466,N_14639);
xnor UO_287 (O_287,N_14341,N_14855);
nand UO_288 (O_288,N_14290,N_14875);
xor UO_289 (O_289,N_14520,N_14787);
or UO_290 (O_290,N_14389,N_14316);
and UO_291 (O_291,N_14496,N_14689);
xnor UO_292 (O_292,N_14896,N_14553);
nand UO_293 (O_293,N_14780,N_14469);
nand UO_294 (O_294,N_14715,N_14781);
or UO_295 (O_295,N_14716,N_14631);
nand UO_296 (O_296,N_14367,N_14863);
nor UO_297 (O_297,N_14459,N_14650);
or UO_298 (O_298,N_14270,N_14987);
xnor UO_299 (O_299,N_14880,N_14879);
nand UO_300 (O_300,N_14913,N_14398);
xnor UO_301 (O_301,N_14322,N_14695);
or UO_302 (O_302,N_14933,N_14357);
nand UO_303 (O_303,N_14535,N_14425);
xnor UO_304 (O_304,N_14327,N_14641);
nor UO_305 (O_305,N_14506,N_14898);
nand UO_306 (O_306,N_14652,N_14407);
or UO_307 (O_307,N_14490,N_14672);
or UO_308 (O_308,N_14472,N_14795);
nor UO_309 (O_309,N_14524,N_14832);
nor UO_310 (O_310,N_14405,N_14519);
nand UO_311 (O_311,N_14731,N_14417);
nand UO_312 (O_312,N_14446,N_14567);
nand UO_313 (O_313,N_14541,N_14421);
and UO_314 (O_314,N_14883,N_14416);
xnor UO_315 (O_315,N_14848,N_14969);
nor UO_316 (O_316,N_14978,N_14460);
nand UO_317 (O_317,N_14450,N_14804);
or UO_318 (O_318,N_14932,N_14558);
or UO_319 (O_319,N_14369,N_14838);
nor UO_320 (O_320,N_14730,N_14431);
xnor UO_321 (O_321,N_14844,N_14820);
and UO_322 (O_322,N_14923,N_14335);
nand UO_323 (O_323,N_14626,N_14979);
nand UO_324 (O_324,N_14507,N_14395);
xnor UO_325 (O_325,N_14907,N_14559);
and UO_326 (O_326,N_14926,N_14900);
and UO_327 (O_327,N_14517,N_14783);
nand UO_328 (O_328,N_14634,N_14998);
or UO_329 (O_329,N_14611,N_14941);
nor UO_330 (O_330,N_14806,N_14555);
nor UO_331 (O_331,N_14380,N_14717);
or UO_332 (O_332,N_14255,N_14300);
or UO_333 (O_333,N_14320,N_14594);
and UO_334 (O_334,N_14957,N_14504);
xor UO_335 (O_335,N_14946,N_14323);
nand UO_336 (O_336,N_14992,N_14908);
or UO_337 (O_337,N_14994,N_14906);
nand UO_338 (O_338,N_14458,N_14962);
nor UO_339 (O_339,N_14947,N_14481);
nand UO_340 (O_340,N_14487,N_14867);
and UO_341 (O_341,N_14659,N_14961);
nand UO_342 (O_342,N_14515,N_14284);
and UO_343 (O_343,N_14728,N_14696);
and UO_344 (O_344,N_14330,N_14319);
and UO_345 (O_345,N_14468,N_14702);
xor UO_346 (O_346,N_14283,N_14615);
and UO_347 (O_347,N_14682,N_14911);
or UO_348 (O_348,N_14667,N_14614);
xor UO_349 (O_349,N_14325,N_14683);
and UO_350 (O_350,N_14971,N_14973);
nand UO_351 (O_351,N_14275,N_14557);
nor UO_352 (O_352,N_14885,N_14400);
or UO_353 (O_353,N_14296,N_14392);
or UO_354 (O_354,N_14849,N_14858);
nor UO_355 (O_355,N_14603,N_14805);
and UO_356 (O_356,N_14909,N_14442);
nor UO_357 (O_357,N_14756,N_14924);
and UO_358 (O_358,N_14772,N_14344);
nor UO_359 (O_359,N_14477,N_14423);
and UO_360 (O_360,N_14253,N_14385);
xor UO_361 (O_361,N_14547,N_14370);
and UO_362 (O_362,N_14912,N_14600);
nor UO_363 (O_363,N_14859,N_14521);
or UO_364 (O_364,N_14654,N_14633);
nand UO_365 (O_365,N_14493,N_14409);
xnor UO_366 (O_366,N_14464,N_14467);
xnor UO_367 (O_367,N_14782,N_14430);
nand UO_368 (O_368,N_14974,N_14285);
nand UO_369 (O_369,N_14747,N_14835);
xor UO_370 (O_370,N_14984,N_14293);
xnor UO_371 (O_371,N_14657,N_14632);
xnor UO_372 (O_372,N_14448,N_14288);
nor UO_373 (O_373,N_14704,N_14636);
or UO_374 (O_374,N_14257,N_14681);
and UO_375 (O_375,N_14714,N_14644);
or UO_376 (O_376,N_14919,N_14646);
xor UO_377 (O_377,N_14663,N_14756);
and UO_378 (O_378,N_14824,N_14616);
nand UO_379 (O_379,N_14730,N_14355);
xor UO_380 (O_380,N_14274,N_14338);
or UO_381 (O_381,N_14802,N_14647);
or UO_382 (O_382,N_14965,N_14711);
nand UO_383 (O_383,N_14304,N_14485);
or UO_384 (O_384,N_14969,N_14387);
nor UO_385 (O_385,N_14526,N_14421);
or UO_386 (O_386,N_14832,N_14393);
and UO_387 (O_387,N_14729,N_14814);
or UO_388 (O_388,N_14580,N_14471);
nor UO_389 (O_389,N_14669,N_14850);
and UO_390 (O_390,N_14907,N_14549);
or UO_391 (O_391,N_14908,N_14841);
nor UO_392 (O_392,N_14703,N_14659);
and UO_393 (O_393,N_14968,N_14780);
xnor UO_394 (O_394,N_14339,N_14360);
nand UO_395 (O_395,N_14518,N_14304);
or UO_396 (O_396,N_14926,N_14265);
xor UO_397 (O_397,N_14738,N_14303);
nand UO_398 (O_398,N_14573,N_14402);
nand UO_399 (O_399,N_14888,N_14671);
and UO_400 (O_400,N_14689,N_14870);
xnor UO_401 (O_401,N_14702,N_14823);
nand UO_402 (O_402,N_14767,N_14685);
or UO_403 (O_403,N_14692,N_14470);
and UO_404 (O_404,N_14682,N_14448);
and UO_405 (O_405,N_14423,N_14525);
and UO_406 (O_406,N_14769,N_14273);
nand UO_407 (O_407,N_14909,N_14984);
and UO_408 (O_408,N_14487,N_14937);
xnor UO_409 (O_409,N_14638,N_14536);
or UO_410 (O_410,N_14883,N_14894);
xnor UO_411 (O_411,N_14559,N_14767);
or UO_412 (O_412,N_14674,N_14829);
or UO_413 (O_413,N_14948,N_14699);
nor UO_414 (O_414,N_14442,N_14874);
xnor UO_415 (O_415,N_14629,N_14985);
nand UO_416 (O_416,N_14378,N_14707);
xor UO_417 (O_417,N_14864,N_14581);
nor UO_418 (O_418,N_14405,N_14279);
xor UO_419 (O_419,N_14412,N_14391);
and UO_420 (O_420,N_14391,N_14842);
nand UO_421 (O_421,N_14969,N_14376);
xor UO_422 (O_422,N_14601,N_14546);
or UO_423 (O_423,N_14833,N_14332);
nor UO_424 (O_424,N_14954,N_14424);
nor UO_425 (O_425,N_14303,N_14426);
and UO_426 (O_426,N_14477,N_14540);
or UO_427 (O_427,N_14362,N_14509);
or UO_428 (O_428,N_14448,N_14783);
nor UO_429 (O_429,N_14654,N_14291);
nand UO_430 (O_430,N_14436,N_14332);
and UO_431 (O_431,N_14493,N_14305);
nor UO_432 (O_432,N_14489,N_14761);
nor UO_433 (O_433,N_14455,N_14862);
or UO_434 (O_434,N_14595,N_14396);
and UO_435 (O_435,N_14831,N_14592);
nand UO_436 (O_436,N_14444,N_14551);
and UO_437 (O_437,N_14262,N_14332);
and UO_438 (O_438,N_14411,N_14960);
xor UO_439 (O_439,N_14653,N_14965);
xnor UO_440 (O_440,N_14368,N_14826);
or UO_441 (O_441,N_14798,N_14698);
and UO_442 (O_442,N_14658,N_14835);
or UO_443 (O_443,N_14379,N_14512);
nor UO_444 (O_444,N_14316,N_14551);
xnor UO_445 (O_445,N_14519,N_14782);
xnor UO_446 (O_446,N_14434,N_14831);
xnor UO_447 (O_447,N_14644,N_14938);
or UO_448 (O_448,N_14798,N_14470);
nand UO_449 (O_449,N_14630,N_14327);
nand UO_450 (O_450,N_14353,N_14443);
nand UO_451 (O_451,N_14332,N_14296);
and UO_452 (O_452,N_14320,N_14613);
xnor UO_453 (O_453,N_14589,N_14844);
nor UO_454 (O_454,N_14929,N_14433);
nand UO_455 (O_455,N_14616,N_14816);
xor UO_456 (O_456,N_14663,N_14593);
and UO_457 (O_457,N_14316,N_14289);
xnor UO_458 (O_458,N_14757,N_14882);
xor UO_459 (O_459,N_14726,N_14406);
nor UO_460 (O_460,N_14735,N_14524);
and UO_461 (O_461,N_14824,N_14841);
and UO_462 (O_462,N_14294,N_14695);
xnor UO_463 (O_463,N_14614,N_14333);
or UO_464 (O_464,N_14341,N_14340);
nand UO_465 (O_465,N_14296,N_14408);
and UO_466 (O_466,N_14402,N_14793);
nor UO_467 (O_467,N_14381,N_14826);
xnor UO_468 (O_468,N_14608,N_14463);
nor UO_469 (O_469,N_14574,N_14662);
nor UO_470 (O_470,N_14720,N_14857);
or UO_471 (O_471,N_14714,N_14476);
xnor UO_472 (O_472,N_14320,N_14989);
xnor UO_473 (O_473,N_14682,N_14561);
and UO_474 (O_474,N_14579,N_14567);
nor UO_475 (O_475,N_14391,N_14828);
nor UO_476 (O_476,N_14905,N_14970);
nor UO_477 (O_477,N_14419,N_14300);
or UO_478 (O_478,N_14585,N_14616);
xnor UO_479 (O_479,N_14285,N_14712);
nand UO_480 (O_480,N_14348,N_14531);
or UO_481 (O_481,N_14717,N_14284);
or UO_482 (O_482,N_14399,N_14867);
nand UO_483 (O_483,N_14457,N_14310);
nand UO_484 (O_484,N_14820,N_14869);
nand UO_485 (O_485,N_14644,N_14694);
and UO_486 (O_486,N_14830,N_14277);
nor UO_487 (O_487,N_14807,N_14263);
and UO_488 (O_488,N_14952,N_14894);
or UO_489 (O_489,N_14920,N_14695);
and UO_490 (O_490,N_14356,N_14484);
nor UO_491 (O_491,N_14280,N_14571);
nor UO_492 (O_492,N_14309,N_14492);
nor UO_493 (O_493,N_14828,N_14574);
xnor UO_494 (O_494,N_14445,N_14836);
or UO_495 (O_495,N_14854,N_14268);
nand UO_496 (O_496,N_14955,N_14571);
or UO_497 (O_497,N_14430,N_14976);
nand UO_498 (O_498,N_14624,N_14607);
nor UO_499 (O_499,N_14740,N_14947);
and UO_500 (O_500,N_14592,N_14425);
nand UO_501 (O_501,N_14868,N_14289);
xor UO_502 (O_502,N_14621,N_14572);
nand UO_503 (O_503,N_14581,N_14751);
xor UO_504 (O_504,N_14274,N_14788);
nand UO_505 (O_505,N_14340,N_14257);
and UO_506 (O_506,N_14801,N_14394);
nand UO_507 (O_507,N_14533,N_14445);
xor UO_508 (O_508,N_14784,N_14680);
nor UO_509 (O_509,N_14972,N_14763);
or UO_510 (O_510,N_14975,N_14854);
nand UO_511 (O_511,N_14521,N_14913);
nand UO_512 (O_512,N_14284,N_14854);
xor UO_513 (O_513,N_14978,N_14464);
or UO_514 (O_514,N_14650,N_14271);
nor UO_515 (O_515,N_14742,N_14749);
and UO_516 (O_516,N_14766,N_14611);
xor UO_517 (O_517,N_14569,N_14542);
and UO_518 (O_518,N_14469,N_14695);
and UO_519 (O_519,N_14818,N_14373);
and UO_520 (O_520,N_14979,N_14384);
and UO_521 (O_521,N_14617,N_14323);
or UO_522 (O_522,N_14868,N_14606);
or UO_523 (O_523,N_14357,N_14455);
or UO_524 (O_524,N_14630,N_14790);
xor UO_525 (O_525,N_14701,N_14493);
and UO_526 (O_526,N_14339,N_14757);
xnor UO_527 (O_527,N_14897,N_14552);
or UO_528 (O_528,N_14306,N_14722);
xor UO_529 (O_529,N_14847,N_14309);
nand UO_530 (O_530,N_14500,N_14858);
nor UO_531 (O_531,N_14383,N_14527);
nand UO_532 (O_532,N_14977,N_14345);
and UO_533 (O_533,N_14418,N_14384);
or UO_534 (O_534,N_14371,N_14946);
and UO_535 (O_535,N_14634,N_14483);
nand UO_536 (O_536,N_14933,N_14470);
or UO_537 (O_537,N_14306,N_14405);
or UO_538 (O_538,N_14262,N_14728);
and UO_539 (O_539,N_14644,N_14985);
xor UO_540 (O_540,N_14917,N_14674);
and UO_541 (O_541,N_14524,N_14806);
nand UO_542 (O_542,N_14777,N_14398);
nor UO_543 (O_543,N_14641,N_14493);
nor UO_544 (O_544,N_14596,N_14402);
nand UO_545 (O_545,N_14648,N_14534);
nor UO_546 (O_546,N_14722,N_14892);
xnor UO_547 (O_547,N_14338,N_14817);
nor UO_548 (O_548,N_14894,N_14595);
or UO_549 (O_549,N_14519,N_14789);
nor UO_550 (O_550,N_14834,N_14994);
xor UO_551 (O_551,N_14485,N_14600);
and UO_552 (O_552,N_14479,N_14992);
and UO_553 (O_553,N_14915,N_14731);
and UO_554 (O_554,N_14801,N_14305);
nor UO_555 (O_555,N_14913,N_14592);
nand UO_556 (O_556,N_14500,N_14607);
xnor UO_557 (O_557,N_14738,N_14445);
nor UO_558 (O_558,N_14975,N_14856);
nand UO_559 (O_559,N_14969,N_14633);
nor UO_560 (O_560,N_14576,N_14999);
xor UO_561 (O_561,N_14605,N_14509);
nor UO_562 (O_562,N_14628,N_14433);
xnor UO_563 (O_563,N_14943,N_14822);
nand UO_564 (O_564,N_14602,N_14603);
xor UO_565 (O_565,N_14511,N_14522);
xor UO_566 (O_566,N_14951,N_14389);
and UO_567 (O_567,N_14353,N_14807);
xnor UO_568 (O_568,N_14962,N_14271);
and UO_569 (O_569,N_14419,N_14318);
nand UO_570 (O_570,N_14817,N_14276);
xor UO_571 (O_571,N_14651,N_14539);
and UO_572 (O_572,N_14776,N_14570);
nand UO_573 (O_573,N_14312,N_14284);
nand UO_574 (O_574,N_14650,N_14942);
xor UO_575 (O_575,N_14594,N_14657);
nand UO_576 (O_576,N_14400,N_14735);
and UO_577 (O_577,N_14736,N_14575);
xor UO_578 (O_578,N_14752,N_14792);
xor UO_579 (O_579,N_14484,N_14393);
nand UO_580 (O_580,N_14608,N_14466);
and UO_581 (O_581,N_14652,N_14465);
or UO_582 (O_582,N_14602,N_14394);
nand UO_583 (O_583,N_14376,N_14297);
xnor UO_584 (O_584,N_14365,N_14861);
or UO_585 (O_585,N_14494,N_14510);
nor UO_586 (O_586,N_14372,N_14556);
and UO_587 (O_587,N_14933,N_14691);
or UO_588 (O_588,N_14981,N_14542);
nor UO_589 (O_589,N_14297,N_14580);
nand UO_590 (O_590,N_14659,N_14379);
and UO_591 (O_591,N_14798,N_14807);
xnor UO_592 (O_592,N_14662,N_14818);
xor UO_593 (O_593,N_14776,N_14437);
nand UO_594 (O_594,N_14994,N_14397);
or UO_595 (O_595,N_14719,N_14859);
xnor UO_596 (O_596,N_14259,N_14935);
xnor UO_597 (O_597,N_14740,N_14980);
and UO_598 (O_598,N_14851,N_14879);
xor UO_599 (O_599,N_14833,N_14368);
and UO_600 (O_600,N_14400,N_14310);
nor UO_601 (O_601,N_14606,N_14995);
nand UO_602 (O_602,N_14423,N_14534);
nand UO_603 (O_603,N_14875,N_14308);
and UO_604 (O_604,N_14620,N_14264);
xor UO_605 (O_605,N_14525,N_14790);
or UO_606 (O_606,N_14458,N_14517);
nand UO_607 (O_607,N_14675,N_14560);
and UO_608 (O_608,N_14679,N_14758);
xnor UO_609 (O_609,N_14274,N_14613);
xor UO_610 (O_610,N_14303,N_14322);
nand UO_611 (O_611,N_14543,N_14444);
or UO_612 (O_612,N_14895,N_14913);
nor UO_613 (O_613,N_14357,N_14803);
or UO_614 (O_614,N_14843,N_14402);
and UO_615 (O_615,N_14696,N_14378);
or UO_616 (O_616,N_14259,N_14947);
and UO_617 (O_617,N_14984,N_14881);
nor UO_618 (O_618,N_14649,N_14366);
and UO_619 (O_619,N_14518,N_14693);
xnor UO_620 (O_620,N_14529,N_14536);
nand UO_621 (O_621,N_14809,N_14507);
nand UO_622 (O_622,N_14734,N_14899);
nand UO_623 (O_623,N_14916,N_14744);
and UO_624 (O_624,N_14876,N_14900);
nor UO_625 (O_625,N_14692,N_14379);
nor UO_626 (O_626,N_14675,N_14460);
and UO_627 (O_627,N_14879,N_14836);
xnor UO_628 (O_628,N_14266,N_14319);
nand UO_629 (O_629,N_14724,N_14805);
or UO_630 (O_630,N_14301,N_14336);
and UO_631 (O_631,N_14318,N_14860);
and UO_632 (O_632,N_14418,N_14385);
and UO_633 (O_633,N_14985,N_14763);
nand UO_634 (O_634,N_14478,N_14528);
and UO_635 (O_635,N_14976,N_14687);
nor UO_636 (O_636,N_14849,N_14351);
xnor UO_637 (O_637,N_14642,N_14578);
and UO_638 (O_638,N_14845,N_14520);
xor UO_639 (O_639,N_14937,N_14766);
and UO_640 (O_640,N_14958,N_14689);
nand UO_641 (O_641,N_14906,N_14805);
or UO_642 (O_642,N_14793,N_14844);
nand UO_643 (O_643,N_14572,N_14775);
or UO_644 (O_644,N_14636,N_14346);
nand UO_645 (O_645,N_14819,N_14840);
or UO_646 (O_646,N_14836,N_14490);
nor UO_647 (O_647,N_14307,N_14814);
and UO_648 (O_648,N_14620,N_14443);
or UO_649 (O_649,N_14738,N_14741);
or UO_650 (O_650,N_14956,N_14813);
nand UO_651 (O_651,N_14509,N_14504);
nand UO_652 (O_652,N_14264,N_14962);
or UO_653 (O_653,N_14582,N_14532);
and UO_654 (O_654,N_14403,N_14959);
xnor UO_655 (O_655,N_14594,N_14345);
nor UO_656 (O_656,N_14356,N_14641);
xor UO_657 (O_657,N_14884,N_14786);
nor UO_658 (O_658,N_14365,N_14834);
nor UO_659 (O_659,N_14262,N_14322);
nand UO_660 (O_660,N_14840,N_14318);
xor UO_661 (O_661,N_14402,N_14597);
xor UO_662 (O_662,N_14587,N_14308);
or UO_663 (O_663,N_14696,N_14513);
nor UO_664 (O_664,N_14842,N_14420);
nor UO_665 (O_665,N_14978,N_14945);
xor UO_666 (O_666,N_14933,N_14701);
nand UO_667 (O_667,N_14566,N_14880);
nor UO_668 (O_668,N_14791,N_14607);
nand UO_669 (O_669,N_14836,N_14825);
nor UO_670 (O_670,N_14831,N_14709);
xor UO_671 (O_671,N_14883,N_14377);
xor UO_672 (O_672,N_14296,N_14453);
or UO_673 (O_673,N_14876,N_14448);
nor UO_674 (O_674,N_14699,N_14827);
nand UO_675 (O_675,N_14704,N_14811);
xor UO_676 (O_676,N_14399,N_14644);
nor UO_677 (O_677,N_14374,N_14913);
xor UO_678 (O_678,N_14373,N_14437);
or UO_679 (O_679,N_14471,N_14784);
and UO_680 (O_680,N_14724,N_14602);
xnor UO_681 (O_681,N_14651,N_14750);
nor UO_682 (O_682,N_14760,N_14978);
or UO_683 (O_683,N_14608,N_14513);
nand UO_684 (O_684,N_14479,N_14821);
or UO_685 (O_685,N_14763,N_14711);
nand UO_686 (O_686,N_14292,N_14596);
nand UO_687 (O_687,N_14746,N_14507);
nand UO_688 (O_688,N_14310,N_14996);
xnor UO_689 (O_689,N_14586,N_14685);
xnor UO_690 (O_690,N_14904,N_14940);
nor UO_691 (O_691,N_14522,N_14371);
or UO_692 (O_692,N_14834,N_14485);
nand UO_693 (O_693,N_14647,N_14287);
nand UO_694 (O_694,N_14454,N_14256);
nand UO_695 (O_695,N_14831,N_14841);
and UO_696 (O_696,N_14917,N_14435);
xnor UO_697 (O_697,N_14449,N_14709);
xor UO_698 (O_698,N_14284,N_14421);
and UO_699 (O_699,N_14476,N_14440);
and UO_700 (O_700,N_14539,N_14848);
nor UO_701 (O_701,N_14347,N_14544);
nor UO_702 (O_702,N_14359,N_14308);
nor UO_703 (O_703,N_14828,N_14830);
nand UO_704 (O_704,N_14762,N_14664);
and UO_705 (O_705,N_14797,N_14471);
nand UO_706 (O_706,N_14719,N_14494);
nand UO_707 (O_707,N_14279,N_14536);
nand UO_708 (O_708,N_14401,N_14858);
nor UO_709 (O_709,N_14698,N_14968);
nand UO_710 (O_710,N_14908,N_14767);
xor UO_711 (O_711,N_14514,N_14873);
nor UO_712 (O_712,N_14460,N_14618);
and UO_713 (O_713,N_14405,N_14533);
xnor UO_714 (O_714,N_14489,N_14314);
xor UO_715 (O_715,N_14302,N_14590);
xor UO_716 (O_716,N_14830,N_14302);
nor UO_717 (O_717,N_14932,N_14861);
nand UO_718 (O_718,N_14260,N_14409);
or UO_719 (O_719,N_14311,N_14294);
xor UO_720 (O_720,N_14581,N_14829);
nor UO_721 (O_721,N_14951,N_14353);
nand UO_722 (O_722,N_14997,N_14474);
nand UO_723 (O_723,N_14768,N_14774);
or UO_724 (O_724,N_14355,N_14764);
or UO_725 (O_725,N_14922,N_14672);
and UO_726 (O_726,N_14720,N_14880);
xor UO_727 (O_727,N_14718,N_14340);
and UO_728 (O_728,N_14803,N_14461);
or UO_729 (O_729,N_14791,N_14777);
xor UO_730 (O_730,N_14788,N_14584);
nand UO_731 (O_731,N_14842,N_14306);
xnor UO_732 (O_732,N_14508,N_14716);
and UO_733 (O_733,N_14783,N_14942);
and UO_734 (O_734,N_14636,N_14908);
nand UO_735 (O_735,N_14444,N_14768);
or UO_736 (O_736,N_14560,N_14544);
nor UO_737 (O_737,N_14967,N_14538);
nor UO_738 (O_738,N_14544,N_14798);
nor UO_739 (O_739,N_14611,N_14585);
or UO_740 (O_740,N_14553,N_14546);
or UO_741 (O_741,N_14821,N_14265);
xnor UO_742 (O_742,N_14939,N_14436);
and UO_743 (O_743,N_14415,N_14987);
nand UO_744 (O_744,N_14925,N_14844);
and UO_745 (O_745,N_14972,N_14920);
or UO_746 (O_746,N_14267,N_14453);
xnor UO_747 (O_747,N_14336,N_14529);
and UO_748 (O_748,N_14612,N_14743);
and UO_749 (O_749,N_14585,N_14704);
nor UO_750 (O_750,N_14496,N_14628);
nand UO_751 (O_751,N_14279,N_14635);
xor UO_752 (O_752,N_14590,N_14760);
or UO_753 (O_753,N_14627,N_14413);
and UO_754 (O_754,N_14336,N_14857);
and UO_755 (O_755,N_14562,N_14460);
nor UO_756 (O_756,N_14651,N_14598);
or UO_757 (O_757,N_14456,N_14967);
and UO_758 (O_758,N_14395,N_14893);
xor UO_759 (O_759,N_14771,N_14413);
and UO_760 (O_760,N_14615,N_14679);
and UO_761 (O_761,N_14996,N_14986);
or UO_762 (O_762,N_14885,N_14602);
xnor UO_763 (O_763,N_14460,N_14919);
xor UO_764 (O_764,N_14302,N_14711);
xnor UO_765 (O_765,N_14546,N_14587);
nand UO_766 (O_766,N_14604,N_14592);
nand UO_767 (O_767,N_14589,N_14809);
and UO_768 (O_768,N_14740,N_14787);
xnor UO_769 (O_769,N_14369,N_14695);
xnor UO_770 (O_770,N_14952,N_14704);
nand UO_771 (O_771,N_14300,N_14992);
xnor UO_772 (O_772,N_14680,N_14777);
nor UO_773 (O_773,N_14324,N_14968);
and UO_774 (O_774,N_14879,N_14661);
and UO_775 (O_775,N_14884,N_14514);
nand UO_776 (O_776,N_14942,N_14575);
nand UO_777 (O_777,N_14555,N_14472);
and UO_778 (O_778,N_14309,N_14491);
xor UO_779 (O_779,N_14941,N_14392);
xnor UO_780 (O_780,N_14842,N_14645);
nor UO_781 (O_781,N_14778,N_14568);
xnor UO_782 (O_782,N_14887,N_14337);
xor UO_783 (O_783,N_14897,N_14577);
nor UO_784 (O_784,N_14658,N_14928);
nand UO_785 (O_785,N_14805,N_14502);
nor UO_786 (O_786,N_14990,N_14449);
nand UO_787 (O_787,N_14693,N_14740);
xor UO_788 (O_788,N_14328,N_14695);
nor UO_789 (O_789,N_14860,N_14412);
nand UO_790 (O_790,N_14726,N_14285);
nand UO_791 (O_791,N_14523,N_14521);
nand UO_792 (O_792,N_14433,N_14753);
or UO_793 (O_793,N_14529,N_14831);
and UO_794 (O_794,N_14425,N_14494);
or UO_795 (O_795,N_14772,N_14518);
or UO_796 (O_796,N_14739,N_14652);
or UO_797 (O_797,N_14476,N_14578);
nand UO_798 (O_798,N_14749,N_14280);
xor UO_799 (O_799,N_14560,N_14484);
and UO_800 (O_800,N_14552,N_14568);
nor UO_801 (O_801,N_14725,N_14314);
or UO_802 (O_802,N_14351,N_14746);
nand UO_803 (O_803,N_14924,N_14431);
and UO_804 (O_804,N_14287,N_14466);
nand UO_805 (O_805,N_14310,N_14903);
nand UO_806 (O_806,N_14999,N_14597);
or UO_807 (O_807,N_14542,N_14764);
xnor UO_808 (O_808,N_14888,N_14336);
nor UO_809 (O_809,N_14929,N_14980);
and UO_810 (O_810,N_14978,N_14624);
nor UO_811 (O_811,N_14405,N_14696);
xor UO_812 (O_812,N_14685,N_14286);
nor UO_813 (O_813,N_14576,N_14658);
and UO_814 (O_814,N_14998,N_14938);
xor UO_815 (O_815,N_14864,N_14435);
xnor UO_816 (O_816,N_14872,N_14376);
xnor UO_817 (O_817,N_14599,N_14674);
and UO_818 (O_818,N_14659,N_14602);
nand UO_819 (O_819,N_14643,N_14327);
and UO_820 (O_820,N_14432,N_14785);
nor UO_821 (O_821,N_14628,N_14303);
and UO_822 (O_822,N_14794,N_14287);
nor UO_823 (O_823,N_14316,N_14524);
nor UO_824 (O_824,N_14334,N_14896);
or UO_825 (O_825,N_14461,N_14366);
and UO_826 (O_826,N_14538,N_14276);
xnor UO_827 (O_827,N_14948,N_14947);
nor UO_828 (O_828,N_14889,N_14497);
and UO_829 (O_829,N_14700,N_14804);
and UO_830 (O_830,N_14640,N_14810);
xnor UO_831 (O_831,N_14842,N_14547);
xor UO_832 (O_832,N_14669,N_14428);
nand UO_833 (O_833,N_14360,N_14839);
xnor UO_834 (O_834,N_14697,N_14728);
nor UO_835 (O_835,N_14914,N_14626);
or UO_836 (O_836,N_14822,N_14545);
and UO_837 (O_837,N_14812,N_14393);
xnor UO_838 (O_838,N_14657,N_14967);
or UO_839 (O_839,N_14322,N_14337);
xor UO_840 (O_840,N_14285,N_14869);
nor UO_841 (O_841,N_14344,N_14539);
nand UO_842 (O_842,N_14806,N_14553);
xor UO_843 (O_843,N_14817,N_14955);
xnor UO_844 (O_844,N_14264,N_14425);
nor UO_845 (O_845,N_14675,N_14605);
or UO_846 (O_846,N_14909,N_14608);
xor UO_847 (O_847,N_14574,N_14458);
and UO_848 (O_848,N_14292,N_14812);
nand UO_849 (O_849,N_14336,N_14852);
and UO_850 (O_850,N_14267,N_14789);
or UO_851 (O_851,N_14924,N_14501);
or UO_852 (O_852,N_14335,N_14269);
nor UO_853 (O_853,N_14839,N_14439);
or UO_854 (O_854,N_14965,N_14531);
nor UO_855 (O_855,N_14491,N_14303);
or UO_856 (O_856,N_14275,N_14464);
and UO_857 (O_857,N_14268,N_14711);
xor UO_858 (O_858,N_14757,N_14818);
nand UO_859 (O_859,N_14486,N_14423);
xor UO_860 (O_860,N_14445,N_14398);
nand UO_861 (O_861,N_14502,N_14488);
xor UO_862 (O_862,N_14969,N_14550);
nand UO_863 (O_863,N_14971,N_14807);
nor UO_864 (O_864,N_14423,N_14939);
nor UO_865 (O_865,N_14839,N_14520);
nand UO_866 (O_866,N_14288,N_14364);
nor UO_867 (O_867,N_14935,N_14812);
or UO_868 (O_868,N_14524,N_14679);
and UO_869 (O_869,N_14336,N_14303);
nand UO_870 (O_870,N_14543,N_14754);
xnor UO_871 (O_871,N_14508,N_14403);
and UO_872 (O_872,N_14732,N_14398);
nand UO_873 (O_873,N_14505,N_14518);
and UO_874 (O_874,N_14802,N_14516);
nand UO_875 (O_875,N_14692,N_14689);
xor UO_876 (O_876,N_14432,N_14964);
or UO_877 (O_877,N_14546,N_14500);
xor UO_878 (O_878,N_14715,N_14643);
nand UO_879 (O_879,N_14456,N_14615);
or UO_880 (O_880,N_14990,N_14697);
xor UO_881 (O_881,N_14312,N_14415);
or UO_882 (O_882,N_14728,N_14516);
or UO_883 (O_883,N_14944,N_14288);
nand UO_884 (O_884,N_14554,N_14749);
nand UO_885 (O_885,N_14926,N_14605);
and UO_886 (O_886,N_14684,N_14736);
nor UO_887 (O_887,N_14892,N_14874);
nand UO_888 (O_888,N_14998,N_14582);
nand UO_889 (O_889,N_14632,N_14706);
nand UO_890 (O_890,N_14397,N_14507);
and UO_891 (O_891,N_14938,N_14976);
or UO_892 (O_892,N_14881,N_14594);
and UO_893 (O_893,N_14978,N_14885);
and UO_894 (O_894,N_14377,N_14262);
nand UO_895 (O_895,N_14800,N_14290);
nand UO_896 (O_896,N_14751,N_14494);
and UO_897 (O_897,N_14791,N_14626);
or UO_898 (O_898,N_14429,N_14727);
xor UO_899 (O_899,N_14707,N_14412);
or UO_900 (O_900,N_14514,N_14918);
and UO_901 (O_901,N_14765,N_14799);
and UO_902 (O_902,N_14508,N_14818);
xnor UO_903 (O_903,N_14498,N_14441);
nand UO_904 (O_904,N_14601,N_14611);
nor UO_905 (O_905,N_14334,N_14700);
nor UO_906 (O_906,N_14312,N_14814);
nor UO_907 (O_907,N_14455,N_14968);
and UO_908 (O_908,N_14607,N_14439);
and UO_909 (O_909,N_14730,N_14328);
nand UO_910 (O_910,N_14286,N_14464);
or UO_911 (O_911,N_14885,N_14664);
nand UO_912 (O_912,N_14802,N_14541);
nor UO_913 (O_913,N_14840,N_14399);
nand UO_914 (O_914,N_14973,N_14653);
or UO_915 (O_915,N_14726,N_14402);
nor UO_916 (O_916,N_14720,N_14614);
and UO_917 (O_917,N_14851,N_14687);
nor UO_918 (O_918,N_14375,N_14992);
or UO_919 (O_919,N_14461,N_14616);
xnor UO_920 (O_920,N_14578,N_14513);
xnor UO_921 (O_921,N_14316,N_14983);
nor UO_922 (O_922,N_14785,N_14740);
and UO_923 (O_923,N_14992,N_14897);
and UO_924 (O_924,N_14258,N_14923);
nor UO_925 (O_925,N_14836,N_14351);
nand UO_926 (O_926,N_14876,N_14743);
nand UO_927 (O_927,N_14794,N_14647);
or UO_928 (O_928,N_14729,N_14582);
nor UO_929 (O_929,N_14295,N_14734);
or UO_930 (O_930,N_14463,N_14645);
or UO_931 (O_931,N_14582,N_14466);
nor UO_932 (O_932,N_14582,N_14458);
or UO_933 (O_933,N_14640,N_14410);
or UO_934 (O_934,N_14948,N_14703);
and UO_935 (O_935,N_14716,N_14340);
or UO_936 (O_936,N_14341,N_14749);
nor UO_937 (O_937,N_14262,N_14343);
nand UO_938 (O_938,N_14768,N_14736);
or UO_939 (O_939,N_14566,N_14408);
xor UO_940 (O_940,N_14706,N_14447);
xnor UO_941 (O_941,N_14683,N_14727);
nand UO_942 (O_942,N_14772,N_14962);
nand UO_943 (O_943,N_14628,N_14921);
or UO_944 (O_944,N_14476,N_14989);
nand UO_945 (O_945,N_14607,N_14376);
or UO_946 (O_946,N_14921,N_14770);
xor UO_947 (O_947,N_14693,N_14895);
xor UO_948 (O_948,N_14681,N_14902);
nand UO_949 (O_949,N_14464,N_14705);
or UO_950 (O_950,N_14802,N_14349);
nor UO_951 (O_951,N_14865,N_14296);
nand UO_952 (O_952,N_14698,N_14853);
nand UO_953 (O_953,N_14729,N_14861);
nor UO_954 (O_954,N_14353,N_14453);
and UO_955 (O_955,N_14722,N_14386);
xnor UO_956 (O_956,N_14781,N_14800);
nand UO_957 (O_957,N_14909,N_14310);
xor UO_958 (O_958,N_14791,N_14397);
nand UO_959 (O_959,N_14290,N_14656);
nor UO_960 (O_960,N_14252,N_14546);
or UO_961 (O_961,N_14945,N_14531);
nand UO_962 (O_962,N_14636,N_14318);
nor UO_963 (O_963,N_14751,N_14708);
and UO_964 (O_964,N_14802,N_14703);
and UO_965 (O_965,N_14387,N_14957);
or UO_966 (O_966,N_14299,N_14614);
nand UO_967 (O_967,N_14884,N_14430);
nor UO_968 (O_968,N_14952,N_14812);
nor UO_969 (O_969,N_14591,N_14364);
nand UO_970 (O_970,N_14830,N_14292);
nor UO_971 (O_971,N_14601,N_14301);
nand UO_972 (O_972,N_14485,N_14473);
xor UO_973 (O_973,N_14889,N_14698);
nor UO_974 (O_974,N_14830,N_14427);
xnor UO_975 (O_975,N_14878,N_14343);
or UO_976 (O_976,N_14445,N_14773);
xor UO_977 (O_977,N_14830,N_14780);
or UO_978 (O_978,N_14598,N_14618);
nor UO_979 (O_979,N_14541,N_14656);
xnor UO_980 (O_980,N_14740,N_14429);
nor UO_981 (O_981,N_14697,N_14479);
nor UO_982 (O_982,N_14894,N_14562);
xnor UO_983 (O_983,N_14729,N_14970);
and UO_984 (O_984,N_14551,N_14933);
xor UO_985 (O_985,N_14378,N_14758);
and UO_986 (O_986,N_14359,N_14894);
nor UO_987 (O_987,N_14432,N_14333);
or UO_988 (O_988,N_14407,N_14689);
nand UO_989 (O_989,N_14366,N_14993);
and UO_990 (O_990,N_14780,N_14726);
xnor UO_991 (O_991,N_14717,N_14900);
nand UO_992 (O_992,N_14978,N_14593);
nor UO_993 (O_993,N_14462,N_14945);
nand UO_994 (O_994,N_14974,N_14262);
xor UO_995 (O_995,N_14859,N_14915);
or UO_996 (O_996,N_14863,N_14429);
or UO_997 (O_997,N_14891,N_14987);
nor UO_998 (O_998,N_14932,N_14752);
and UO_999 (O_999,N_14325,N_14565);
and UO_1000 (O_1000,N_14474,N_14297);
xor UO_1001 (O_1001,N_14381,N_14770);
nor UO_1002 (O_1002,N_14466,N_14621);
and UO_1003 (O_1003,N_14904,N_14838);
xor UO_1004 (O_1004,N_14848,N_14692);
and UO_1005 (O_1005,N_14381,N_14408);
nor UO_1006 (O_1006,N_14398,N_14340);
and UO_1007 (O_1007,N_14493,N_14479);
nand UO_1008 (O_1008,N_14981,N_14351);
and UO_1009 (O_1009,N_14573,N_14743);
nor UO_1010 (O_1010,N_14387,N_14891);
or UO_1011 (O_1011,N_14522,N_14830);
xnor UO_1012 (O_1012,N_14653,N_14359);
and UO_1013 (O_1013,N_14484,N_14405);
and UO_1014 (O_1014,N_14417,N_14519);
nor UO_1015 (O_1015,N_14348,N_14511);
nor UO_1016 (O_1016,N_14731,N_14406);
or UO_1017 (O_1017,N_14882,N_14459);
nand UO_1018 (O_1018,N_14707,N_14589);
and UO_1019 (O_1019,N_14692,N_14404);
or UO_1020 (O_1020,N_14850,N_14463);
and UO_1021 (O_1021,N_14440,N_14984);
xnor UO_1022 (O_1022,N_14636,N_14711);
nand UO_1023 (O_1023,N_14291,N_14681);
nor UO_1024 (O_1024,N_14957,N_14578);
or UO_1025 (O_1025,N_14432,N_14745);
nand UO_1026 (O_1026,N_14436,N_14550);
nor UO_1027 (O_1027,N_14601,N_14694);
nand UO_1028 (O_1028,N_14381,N_14457);
and UO_1029 (O_1029,N_14553,N_14703);
and UO_1030 (O_1030,N_14942,N_14587);
nand UO_1031 (O_1031,N_14668,N_14266);
and UO_1032 (O_1032,N_14922,N_14795);
nand UO_1033 (O_1033,N_14689,N_14603);
or UO_1034 (O_1034,N_14704,N_14336);
or UO_1035 (O_1035,N_14847,N_14585);
xor UO_1036 (O_1036,N_14333,N_14635);
nor UO_1037 (O_1037,N_14864,N_14268);
nor UO_1038 (O_1038,N_14298,N_14537);
nand UO_1039 (O_1039,N_14722,N_14322);
nand UO_1040 (O_1040,N_14821,N_14837);
nand UO_1041 (O_1041,N_14808,N_14784);
xor UO_1042 (O_1042,N_14501,N_14319);
xor UO_1043 (O_1043,N_14409,N_14676);
nand UO_1044 (O_1044,N_14585,N_14530);
xor UO_1045 (O_1045,N_14648,N_14780);
nand UO_1046 (O_1046,N_14513,N_14667);
xor UO_1047 (O_1047,N_14506,N_14876);
or UO_1048 (O_1048,N_14875,N_14637);
nor UO_1049 (O_1049,N_14948,N_14923);
and UO_1050 (O_1050,N_14993,N_14672);
nor UO_1051 (O_1051,N_14730,N_14402);
xnor UO_1052 (O_1052,N_14564,N_14855);
and UO_1053 (O_1053,N_14488,N_14783);
xnor UO_1054 (O_1054,N_14612,N_14362);
nor UO_1055 (O_1055,N_14398,N_14266);
nand UO_1056 (O_1056,N_14288,N_14927);
nor UO_1057 (O_1057,N_14658,N_14644);
and UO_1058 (O_1058,N_14640,N_14903);
nor UO_1059 (O_1059,N_14967,N_14688);
xor UO_1060 (O_1060,N_14588,N_14674);
or UO_1061 (O_1061,N_14452,N_14344);
nand UO_1062 (O_1062,N_14717,N_14957);
nand UO_1063 (O_1063,N_14513,N_14687);
xor UO_1064 (O_1064,N_14480,N_14513);
nor UO_1065 (O_1065,N_14621,N_14858);
and UO_1066 (O_1066,N_14417,N_14363);
and UO_1067 (O_1067,N_14761,N_14958);
and UO_1068 (O_1068,N_14328,N_14896);
xor UO_1069 (O_1069,N_14569,N_14898);
nand UO_1070 (O_1070,N_14422,N_14512);
nand UO_1071 (O_1071,N_14302,N_14641);
nand UO_1072 (O_1072,N_14312,N_14584);
or UO_1073 (O_1073,N_14834,N_14773);
and UO_1074 (O_1074,N_14916,N_14675);
or UO_1075 (O_1075,N_14778,N_14453);
and UO_1076 (O_1076,N_14862,N_14305);
xnor UO_1077 (O_1077,N_14764,N_14735);
or UO_1078 (O_1078,N_14395,N_14441);
or UO_1079 (O_1079,N_14530,N_14435);
or UO_1080 (O_1080,N_14558,N_14942);
nor UO_1081 (O_1081,N_14888,N_14424);
and UO_1082 (O_1082,N_14892,N_14519);
and UO_1083 (O_1083,N_14954,N_14776);
nor UO_1084 (O_1084,N_14535,N_14685);
and UO_1085 (O_1085,N_14377,N_14773);
and UO_1086 (O_1086,N_14275,N_14425);
nand UO_1087 (O_1087,N_14537,N_14959);
or UO_1088 (O_1088,N_14570,N_14715);
nor UO_1089 (O_1089,N_14774,N_14722);
and UO_1090 (O_1090,N_14259,N_14432);
or UO_1091 (O_1091,N_14650,N_14889);
or UO_1092 (O_1092,N_14504,N_14822);
nand UO_1093 (O_1093,N_14370,N_14463);
nand UO_1094 (O_1094,N_14292,N_14532);
or UO_1095 (O_1095,N_14892,N_14699);
nand UO_1096 (O_1096,N_14337,N_14656);
and UO_1097 (O_1097,N_14407,N_14388);
nor UO_1098 (O_1098,N_14489,N_14575);
or UO_1099 (O_1099,N_14544,N_14713);
nand UO_1100 (O_1100,N_14963,N_14484);
nand UO_1101 (O_1101,N_14975,N_14936);
and UO_1102 (O_1102,N_14327,N_14372);
nor UO_1103 (O_1103,N_14359,N_14526);
nand UO_1104 (O_1104,N_14924,N_14673);
xnor UO_1105 (O_1105,N_14479,N_14662);
nor UO_1106 (O_1106,N_14527,N_14406);
and UO_1107 (O_1107,N_14829,N_14960);
or UO_1108 (O_1108,N_14971,N_14372);
xnor UO_1109 (O_1109,N_14643,N_14400);
nand UO_1110 (O_1110,N_14380,N_14852);
or UO_1111 (O_1111,N_14948,N_14538);
nor UO_1112 (O_1112,N_14962,N_14822);
nor UO_1113 (O_1113,N_14728,N_14805);
and UO_1114 (O_1114,N_14300,N_14780);
and UO_1115 (O_1115,N_14932,N_14605);
xnor UO_1116 (O_1116,N_14331,N_14936);
nor UO_1117 (O_1117,N_14417,N_14735);
and UO_1118 (O_1118,N_14891,N_14977);
and UO_1119 (O_1119,N_14257,N_14488);
xnor UO_1120 (O_1120,N_14345,N_14670);
xnor UO_1121 (O_1121,N_14970,N_14451);
nand UO_1122 (O_1122,N_14816,N_14257);
or UO_1123 (O_1123,N_14977,N_14652);
nor UO_1124 (O_1124,N_14447,N_14479);
and UO_1125 (O_1125,N_14861,N_14303);
nand UO_1126 (O_1126,N_14415,N_14944);
nand UO_1127 (O_1127,N_14323,N_14343);
or UO_1128 (O_1128,N_14673,N_14689);
nand UO_1129 (O_1129,N_14925,N_14351);
xor UO_1130 (O_1130,N_14256,N_14871);
nand UO_1131 (O_1131,N_14664,N_14505);
nor UO_1132 (O_1132,N_14659,N_14308);
nor UO_1133 (O_1133,N_14757,N_14470);
xor UO_1134 (O_1134,N_14949,N_14526);
or UO_1135 (O_1135,N_14855,N_14474);
and UO_1136 (O_1136,N_14391,N_14608);
nor UO_1137 (O_1137,N_14652,N_14778);
and UO_1138 (O_1138,N_14709,N_14936);
nor UO_1139 (O_1139,N_14700,N_14529);
nand UO_1140 (O_1140,N_14848,N_14255);
or UO_1141 (O_1141,N_14431,N_14256);
nor UO_1142 (O_1142,N_14794,N_14984);
or UO_1143 (O_1143,N_14446,N_14926);
and UO_1144 (O_1144,N_14962,N_14294);
nor UO_1145 (O_1145,N_14775,N_14934);
nor UO_1146 (O_1146,N_14430,N_14898);
nor UO_1147 (O_1147,N_14983,N_14805);
and UO_1148 (O_1148,N_14734,N_14723);
nor UO_1149 (O_1149,N_14422,N_14973);
or UO_1150 (O_1150,N_14473,N_14496);
or UO_1151 (O_1151,N_14539,N_14434);
and UO_1152 (O_1152,N_14497,N_14980);
nor UO_1153 (O_1153,N_14258,N_14489);
or UO_1154 (O_1154,N_14627,N_14970);
nor UO_1155 (O_1155,N_14486,N_14411);
nor UO_1156 (O_1156,N_14329,N_14616);
and UO_1157 (O_1157,N_14822,N_14606);
and UO_1158 (O_1158,N_14498,N_14581);
and UO_1159 (O_1159,N_14501,N_14855);
or UO_1160 (O_1160,N_14572,N_14934);
or UO_1161 (O_1161,N_14398,N_14493);
or UO_1162 (O_1162,N_14965,N_14395);
and UO_1163 (O_1163,N_14633,N_14761);
nor UO_1164 (O_1164,N_14778,N_14807);
nand UO_1165 (O_1165,N_14971,N_14643);
nand UO_1166 (O_1166,N_14468,N_14916);
nand UO_1167 (O_1167,N_14582,N_14584);
nor UO_1168 (O_1168,N_14690,N_14933);
nor UO_1169 (O_1169,N_14466,N_14595);
nand UO_1170 (O_1170,N_14498,N_14437);
or UO_1171 (O_1171,N_14259,N_14567);
xnor UO_1172 (O_1172,N_14848,N_14603);
or UO_1173 (O_1173,N_14882,N_14749);
or UO_1174 (O_1174,N_14851,N_14540);
xnor UO_1175 (O_1175,N_14284,N_14640);
and UO_1176 (O_1176,N_14324,N_14393);
nand UO_1177 (O_1177,N_14993,N_14783);
nor UO_1178 (O_1178,N_14973,N_14735);
nand UO_1179 (O_1179,N_14309,N_14962);
or UO_1180 (O_1180,N_14419,N_14498);
xor UO_1181 (O_1181,N_14905,N_14574);
nor UO_1182 (O_1182,N_14545,N_14809);
and UO_1183 (O_1183,N_14848,N_14353);
xnor UO_1184 (O_1184,N_14297,N_14637);
nor UO_1185 (O_1185,N_14870,N_14977);
or UO_1186 (O_1186,N_14444,N_14471);
xnor UO_1187 (O_1187,N_14432,N_14421);
nor UO_1188 (O_1188,N_14925,N_14412);
or UO_1189 (O_1189,N_14297,N_14536);
nand UO_1190 (O_1190,N_14469,N_14373);
and UO_1191 (O_1191,N_14488,N_14412);
and UO_1192 (O_1192,N_14499,N_14974);
and UO_1193 (O_1193,N_14813,N_14529);
nand UO_1194 (O_1194,N_14808,N_14629);
nand UO_1195 (O_1195,N_14660,N_14391);
nand UO_1196 (O_1196,N_14651,N_14777);
nor UO_1197 (O_1197,N_14440,N_14971);
nand UO_1198 (O_1198,N_14804,N_14478);
or UO_1199 (O_1199,N_14751,N_14636);
nand UO_1200 (O_1200,N_14862,N_14594);
and UO_1201 (O_1201,N_14612,N_14519);
nor UO_1202 (O_1202,N_14682,N_14303);
nand UO_1203 (O_1203,N_14503,N_14775);
or UO_1204 (O_1204,N_14279,N_14281);
or UO_1205 (O_1205,N_14410,N_14726);
or UO_1206 (O_1206,N_14313,N_14792);
and UO_1207 (O_1207,N_14944,N_14356);
nor UO_1208 (O_1208,N_14671,N_14621);
or UO_1209 (O_1209,N_14364,N_14878);
nor UO_1210 (O_1210,N_14815,N_14968);
nor UO_1211 (O_1211,N_14660,N_14566);
nor UO_1212 (O_1212,N_14465,N_14899);
nand UO_1213 (O_1213,N_14497,N_14928);
and UO_1214 (O_1214,N_14656,N_14698);
or UO_1215 (O_1215,N_14969,N_14290);
or UO_1216 (O_1216,N_14414,N_14300);
or UO_1217 (O_1217,N_14441,N_14562);
and UO_1218 (O_1218,N_14821,N_14503);
nor UO_1219 (O_1219,N_14840,N_14664);
xor UO_1220 (O_1220,N_14712,N_14830);
xnor UO_1221 (O_1221,N_14386,N_14697);
and UO_1222 (O_1222,N_14289,N_14932);
nor UO_1223 (O_1223,N_14402,N_14965);
nor UO_1224 (O_1224,N_14666,N_14636);
and UO_1225 (O_1225,N_14558,N_14656);
nand UO_1226 (O_1226,N_14835,N_14570);
xnor UO_1227 (O_1227,N_14793,N_14444);
or UO_1228 (O_1228,N_14690,N_14418);
or UO_1229 (O_1229,N_14840,N_14410);
nand UO_1230 (O_1230,N_14397,N_14686);
xor UO_1231 (O_1231,N_14434,N_14381);
xor UO_1232 (O_1232,N_14985,N_14732);
or UO_1233 (O_1233,N_14807,N_14374);
nand UO_1234 (O_1234,N_14765,N_14553);
nand UO_1235 (O_1235,N_14990,N_14395);
and UO_1236 (O_1236,N_14540,N_14818);
nor UO_1237 (O_1237,N_14575,N_14791);
nor UO_1238 (O_1238,N_14791,N_14595);
and UO_1239 (O_1239,N_14953,N_14689);
nand UO_1240 (O_1240,N_14484,N_14499);
nand UO_1241 (O_1241,N_14413,N_14286);
nand UO_1242 (O_1242,N_14692,N_14490);
xnor UO_1243 (O_1243,N_14461,N_14663);
nor UO_1244 (O_1244,N_14506,N_14972);
nand UO_1245 (O_1245,N_14711,N_14338);
and UO_1246 (O_1246,N_14976,N_14326);
nand UO_1247 (O_1247,N_14871,N_14569);
nor UO_1248 (O_1248,N_14324,N_14525);
nand UO_1249 (O_1249,N_14668,N_14827);
nor UO_1250 (O_1250,N_14471,N_14737);
nand UO_1251 (O_1251,N_14749,N_14697);
nor UO_1252 (O_1252,N_14544,N_14382);
or UO_1253 (O_1253,N_14481,N_14655);
xor UO_1254 (O_1254,N_14533,N_14856);
or UO_1255 (O_1255,N_14278,N_14349);
nor UO_1256 (O_1256,N_14278,N_14928);
xor UO_1257 (O_1257,N_14367,N_14812);
or UO_1258 (O_1258,N_14836,N_14976);
xor UO_1259 (O_1259,N_14567,N_14559);
nand UO_1260 (O_1260,N_14765,N_14940);
nor UO_1261 (O_1261,N_14451,N_14878);
nand UO_1262 (O_1262,N_14264,N_14991);
xor UO_1263 (O_1263,N_14693,N_14945);
nand UO_1264 (O_1264,N_14519,N_14264);
nor UO_1265 (O_1265,N_14920,N_14507);
or UO_1266 (O_1266,N_14900,N_14283);
xor UO_1267 (O_1267,N_14466,N_14340);
and UO_1268 (O_1268,N_14587,N_14903);
and UO_1269 (O_1269,N_14835,N_14699);
nand UO_1270 (O_1270,N_14728,N_14792);
or UO_1271 (O_1271,N_14514,N_14577);
nand UO_1272 (O_1272,N_14402,N_14409);
xnor UO_1273 (O_1273,N_14262,N_14406);
or UO_1274 (O_1274,N_14623,N_14665);
xnor UO_1275 (O_1275,N_14714,N_14640);
nor UO_1276 (O_1276,N_14372,N_14478);
or UO_1277 (O_1277,N_14384,N_14645);
nor UO_1278 (O_1278,N_14655,N_14896);
nor UO_1279 (O_1279,N_14939,N_14435);
and UO_1280 (O_1280,N_14265,N_14373);
nand UO_1281 (O_1281,N_14957,N_14255);
nand UO_1282 (O_1282,N_14577,N_14513);
xor UO_1283 (O_1283,N_14840,N_14298);
and UO_1284 (O_1284,N_14699,N_14984);
nor UO_1285 (O_1285,N_14836,N_14404);
nand UO_1286 (O_1286,N_14370,N_14552);
nand UO_1287 (O_1287,N_14712,N_14538);
nand UO_1288 (O_1288,N_14884,N_14400);
and UO_1289 (O_1289,N_14433,N_14545);
nor UO_1290 (O_1290,N_14858,N_14672);
or UO_1291 (O_1291,N_14446,N_14646);
or UO_1292 (O_1292,N_14620,N_14887);
nand UO_1293 (O_1293,N_14323,N_14955);
and UO_1294 (O_1294,N_14531,N_14336);
nor UO_1295 (O_1295,N_14868,N_14520);
or UO_1296 (O_1296,N_14762,N_14736);
xnor UO_1297 (O_1297,N_14776,N_14733);
xnor UO_1298 (O_1298,N_14327,N_14515);
xor UO_1299 (O_1299,N_14362,N_14906);
and UO_1300 (O_1300,N_14580,N_14304);
nor UO_1301 (O_1301,N_14262,N_14327);
nand UO_1302 (O_1302,N_14939,N_14634);
or UO_1303 (O_1303,N_14848,N_14322);
xor UO_1304 (O_1304,N_14532,N_14770);
or UO_1305 (O_1305,N_14262,N_14555);
or UO_1306 (O_1306,N_14711,N_14461);
or UO_1307 (O_1307,N_14306,N_14967);
nand UO_1308 (O_1308,N_14348,N_14855);
nor UO_1309 (O_1309,N_14923,N_14811);
or UO_1310 (O_1310,N_14308,N_14600);
or UO_1311 (O_1311,N_14358,N_14782);
nor UO_1312 (O_1312,N_14567,N_14645);
nand UO_1313 (O_1313,N_14649,N_14574);
nor UO_1314 (O_1314,N_14787,N_14623);
nor UO_1315 (O_1315,N_14835,N_14394);
and UO_1316 (O_1316,N_14793,N_14308);
or UO_1317 (O_1317,N_14774,N_14370);
and UO_1318 (O_1318,N_14403,N_14720);
or UO_1319 (O_1319,N_14712,N_14320);
xnor UO_1320 (O_1320,N_14669,N_14333);
nor UO_1321 (O_1321,N_14434,N_14811);
or UO_1322 (O_1322,N_14366,N_14409);
nand UO_1323 (O_1323,N_14949,N_14747);
xnor UO_1324 (O_1324,N_14873,N_14552);
nand UO_1325 (O_1325,N_14915,N_14918);
nand UO_1326 (O_1326,N_14911,N_14663);
or UO_1327 (O_1327,N_14918,N_14720);
nand UO_1328 (O_1328,N_14536,N_14466);
nand UO_1329 (O_1329,N_14987,N_14257);
nor UO_1330 (O_1330,N_14500,N_14599);
and UO_1331 (O_1331,N_14566,N_14416);
nand UO_1332 (O_1332,N_14825,N_14464);
nand UO_1333 (O_1333,N_14730,N_14656);
xnor UO_1334 (O_1334,N_14868,N_14477);
nand UO_1335 (O_1335,N_14582,N_14764);
nand UO_1336 (O_1336,N_14633,N_14417);
and UO_1337 (O_1337,N_14676,N_14360);
nand UO_1338 (O_1338,N_14281,N_14999);
nor UO_1339 (O_1339,N_14259,N_14281);
nor UO_1340 (O_1340,N_14402,N_14749);
nand UO_1341 (O_1341,N_14314,N_14920);
nor UO_1342 (O_1342,N_14273,N_14835);
nand UO_1343 (O_1343,N_14678,N_14904);
nor UO_1344 (O_1344,N_14459,N_14756);
and UO_1345 (O_1345,N_14540,N_14726);
and UO_1346 (O_1346,N_14375,N_14920);
xnor UO_1347 (O_1347,N_14655,N_14703);
nor UO_1348 (O_1348,N_14444,N_14965);
and UO_1349 (O_1349,N_14554,N_14259);
and UO_1350 (O_1350,N_14829,N_14359);
xnor UO_1351 (O_1351,N_14719,N_14306);
xnor UO_1352 (O_1352,N_14566,N_14858);
xnor UO_1353 (O_1353,N_14597,N_14691);
nor UO_1354 (O_1354,N_14696,N_14923);
nand UO_1355 (O_1355,N_14611,N_14490);
nor UO_1356 (O_1356,N_14469,N_14996);
or UO_1357 (O_1357,N_14624,N_14882);
and UO_1358 (O_1358,N_14890,N_14578);
nand UO_1359 (O_1359,N_14406,N_14342);
nor UO_1360 (O_1360,N_14936,N_14429);
nand UO_1361 (O_1361,N_14866,N_14757);
xor UO_1362 (O_1362,N_14369,N_14697);
nand UO_1363 (O_1363,N_14422,N_14825);
or UO_1364 (O_1364,N_14941,N_14887);
and UO_1365 (O_1365,N_14584,N_14387);
or UO_1366 (O_1366,N_14266,N_14329);
or UO_1367 (O_1367,N_14607,N_14256);
nand UO_1368 (O_1368,N_14772,N_14847);
xor UO_1369 (O_1369,N_14569,N_14695);
xnor UO_1370 (O_1370,N_14769,N_14669);
nand UO_1371 (O_1371,N_14412,N_14312);
nor UO_1372 (O_1372,N_14770,N_14738);
and UO_1373 (O_1373,N_14922,N_14525);
or UO_1374 (O_1374,N_14306,N_14810);
nor UO_1375 (O_1375,N_14569,N_14750);
nand UO_1376 (O_1376,N_14819,N_14677);
xor UO_1377 (O_1377,N_14821,N_14832);
and UO_1378 (O_1378,N_14928,N_14816);
nor UO_1379 (O_1379,N_14395,N_14758);
nor UO_1380 (O_1380,N_14397,N_14876);
or UO_1381 (O_1381,N_14581,N_14686);
nand UO_1382 (O_1382,N_14364,N_14700);
xnor UO_1383 (O_1383,N_14892,N_14474);
nor UO_1384 (O_1384,N_14823,N_14615);
nor UO_1385 (O_1385,N_14715,N_14795);
and UO_1386 (O_1386,N_14508,N_14266);
xor UO_1387 (O_1387,N_14784,N_14842);
xnor UO_1388 (O_1388,N_14984,N_14375);
xnor UO_1389 (O_1389,N_14415,N_14359);
and UO_1390 (O_1390,N_14907,N_14714);
or UO_1391 (O_1391,N_14846,N_14748);
and UO_1392 (O_1392,N_14743,N_14390);
nand UO_1393 (O_1393,N_14858,N_14300);
and UO_1394 (O_1394,N_14479,N_14272);
and UO_1395 (O_1395,N_14721,N_14536);
nand UO_1396 (O_1396,N_14883,N_14553);
and UO_1397 (O_1397,N_14586,N_14485);
or UO_1398 (O_1398,N_14775,N_14839);
and UO_1399 (O_1399,N_14303,N_14584);
xor UO_1400 (O_1400,N_14588,N_14444);
nand UO_1401 (O_1401,N_14519,N_14631);
xnor UO_1402 (O_1402,N_14287,N_14323);
nor UO_1403 (O_1403,N_14339,N_14399);
and UO_1404 (O_1404,N_14594,N_14693);
xnor UO_1405 (O_1405,N_14352,N_14762);
or UO_1406 (O_1406,N_14813,N_14636);
nor UO_1407 (O_1407,N_14744,N_14895);
or UO_1408 (O_1408,N_14837,N_14665);
xor UO_1409 (O_1409,N_14639,N_14877);
xnor UO_1410 (O_1410,N_14411,N_14365);
nor UO_1411 (O_1411,N_14804,N_14323);
xnor UO_1412 (O_1412,N_14844,N_14717);
nor UO_1413 (O_1413,N_14494,N_14639);
or UO_1414 (O_1414,N_14277,N_14843);
nand UO_1415 (O_1415,N_14491,N_14353);
or UO_1416 (O_1416,N_14971,N_14476);
or UO_1417 (O_1417,N_14563,N_14499);
or UO_1418 (O_1418,N_14722,N_14725);
nand UO_1419 (O_1419,N_14742,N_14988);
and UO_1420 (O_1420,N_14665,N_14922);
xor UO_1421 (O_1421,N_14974,N_14629);
or UO_1422 (O_1422,N_14865,N_14656);
xor UO_1423 (O_1423,N_14889,N_14839);
nand UO_1424 (O_1424,N_14505,N_14339);
nand UO_1425 (O_1425,N_14876,N_14391);
xor UO_1426 (O_1426,N_14750,N_14453);
and UO_1427 (O_1427,N_14478,N_14585);
xor UO_1428 (O_1428,N_14639,N_14633);
and UO_1429 (O_1429,N_14311,N_14555);
and UO_1430 (O_1430,N_14965,N_14280);
and UO_1431 (O_1431,N_14616,N_14645);
or UO_1432 (O_1432,N_14832,N_14332);
nand UO_1433 (O_1433,N_14762,N_14435);
nand UO_1434 (O_1434,N_14678,N_14773);
and UO_1435 (O_1435,N_14398,N_14462);
nor UO_1436 (O_1436,N_14604,N_14895);
nand UO_1437 (O_1437,N_14485,N_14495);
or UO_1438 (O_1438,N_14607,N_14445);
and UO_1439 (O_1439,N_14469,N_14403);
xnor UO_1440 (O_1440,N_14711,N_14542);
xnor UO_1441 (O_1441,N_14919,N_14790);
or UO_1442 (O_1442,N_14433,N_14446);
and UO_1443 (O_1443,N_14255,N_14622);
or UO_1444 (O_1444,N_14700,N_14994);
nand UO_1445 (O_1445,N_14534,N_14517);
and UO_1446 (O_1446,N_14864,N_14651);
or UO_1447 (O_1447,N_14558,N_14317);
nand UO_1448 (O_1448,N_14497,N_14328);
and UO_1449 (O_1449,N_14320,N_14466);
nand UO_1450 (O_1450,N_14597,N_14927);
nor UO_1451 (O_1451,N_14750,N_14848);
or UO_1452 (O_1452,N_14674,N_14611);
or UO_1453 (O_1453,N_14934,N_14443);
nand UO_1454 (O_1454,N_14610,N_14656);
and UO_1455 (O_1455,N_14608,N_14530);
nor UO_1456 (O_1456,N_14376,N_14686);
or UO_1457 (O_1457,N_14522,N_14458);
or UO_1458 (O_1458,N_14928,N_14965);
xor UO_1459 (O_1459,N_14416,N_14279);
and UO_1460 (O_1460,N_14907,N_14340);
nand UO_1461 (O_1461,N_14258,N_14781);
nand UO_1462 (O_1462,N_14983,N_14579);
nor UO_1463 (O_1463,N_14775,N_14360);
xor UO_1464 (O_1464,N_14915,N_14441);
and UO_1465 (O_1465,N_14724,N_14336);
xor UO_1466 (O_1466,N_14778,N_14748);
nand UO_1467 (O_1467,N_14280,N_14643);
nand UO_1468 (O_1468,N_14763,N_14664);
nand UO_1469 (O_1469,N_14747,N_14744);
or UO_1470 (O_1470,N_14623,N_14688);
nor UO_1471 (O_1471,N_14256,N_14657);
and UO_1472 (O_1472,N_14959,N_14751);
nand UO_1473 (O_1473,N_14681,N_14817);
nor UO_1474 (O_1474,N_14893,N_14450);
xnor UO_1475 (O_1475,N_14365,N_14927);
xor UO_1476 (O_1476,N_14323,N_14854);
or UO_1477 (O_1477,N_14816,N_14824);
nor UO_1478 (O_1478,N_14781,N_14544);
nand UO_1479 (O_1479,N_14335,N_14659);
or UO_1480 (O_1480,N_14396,N_14884);
or UO_1481 (O_1481,N_14255,N_14751);
nor UO_1482 (O_1482,N_14546,N_14289);
or UO_1483 (O_1483,N_14301,N_14934);
xnor UO_1484 (O_1484,N_14649,N_14991);
nor UO_1485 (O_1485,N_14912,N_14416);
nand UO_1486 (O_1486,N_14804,N_14940);
or UO_1487 (O_1487,N_14558,N_14613);
or UO_1488 (O_1488,N_14475,N_14325);
or UO_1489 (O_1489,N_14756,N_14722);
xor UO_1490 (O_1490,N_14643,N_14370);
or UO_1491 (O_1491,N_14558,N_14653);
nand UO_1492 (O_1492,N_14445,N_14524);
or UO_1493 (O_1493,N_14891,N_14269);
nand UO_1494 (O_1494,N_14649,N_14757);
nor UO_1495 (O_1495,N_14766,N_14719);
nor UO_1496 (O_1496,N_14926,N_14898);
or UO_1497 (O_1497,N_14447,N_14690);
or UO_1498 (O_1498,N_14929,N_14498);
nand UO_1499 (O_1499,N_14313,N_14632);
nor UO_1500 (O_1500,N_14367,N_14370);
nand UO_1501 (O_1501,N_14500,N_14832);
xor UO_1502 (O_1502,N_14534,N_14385);
nor UO_1503 (O_1503,N_14573,N_14708);
nand UO_1504 (O_1504,N_14772,N_14343);
and UO_1505 (O_1505,N_14288,N_14918);
nor UO_1506 (O_1506,N_14997,N_14437);
nand UO_1507 (O_1507,N_14987,N_14748);
and UO_1508 (O_1508,N_14258,N_14972);
xor UO_1509 (O_1509,N_14803,N_14387);
nor UO_1510 (O_1510,N_14789,N_14864);
or UO_1511 (O_1511,N_14606,N_14520);
nand UO_1512 (O_1512,N_14716,N_14613);
nand UO_1513 (O_1513,N_14676,N_14326);
nor UO_1514 (O_1514,N_14350,N_14752);
xnor UO_1515 (O_1515,N_14678,N_14317);
and UO_1516 (O_1516,N_14392,N_14787);
and UO_1517 (O_1517,N_14274,N_14634);
xnor UO_1518 (O_1518,N_14352,N_14787);
or UO_1519 (O_1519,N_14354,N_14845);
nor UO_1520 (O_1520,N_14628,N_14983);
nor UO_1521 (O_1521,N_14820,N_14902);
and UO_1522 (O_1522,N_14895,N_14937);
nor UO_1523 (O_1523,N_14625,N_14574);
and UO_1524 (O_1524,N_14407,N_14729);
and UO_1525 (O_1525,N_14543,N_14831);
and UO_1526 (O_1526,N_14910,N_14426);
nand UO_1527 (O_1527,N_14574,N_14587);
and UO_1528 (O_1528,N_14475,N_14738);
and UO_1529 (O_1529,N_14567,N_14719);
nor UO_1530 (O_1530,N_14732,N_14754);
xnor UO_1531 (O_1531,N_14320,N_14773);
or UO_1532 (O_1532,N_14572,N_14402);
nand UO_1533 (O_1533,N_14786,N_14412);
or UO_1534 (O_1534,N_14970,N_14250);
xnor UO_1535 (O_1535,N_14724,N_14512);
nand UO_1536 (O_1536,N_14516,N_14420);
xor UO_1537 (O_1537,N_14322,N_14769);
or UO_1538 (O_1538,N_14568,N_14289);
xor UO_1539 (O_1539,N_14922,N_14927);
nand UO_1540 (O_1540,N_14594,N_14447);
nor UO_1541 (O_1541,N_14771,N_14430);
or UO_1542 (O_1542,N_14949,N_14415);
and UO_1543 (O_1543,N_14421,N_14644);
nand UO_1544 (O_1544,N_14382,N_14377);
or UO_1545 (O_1545,N_14612,N_14583);
nor UO_1546 (O_1546,N_14964,N_14312);
nor UO_1547 (O_1547,N_14806,N_14986);
nand UO_1548 (O_1548,N_14583,N_14682);
nor UO_1549 (O_1549,N_14795,N_14860);
or UO_1550 (O_1550,N_14883,N_14588);
nand UO_1551 (O_1551,N_14576,N_14698);
nand UO_1552 (O_1552,N_14935,N_14775);
nand UO_1553 (O_1553,N_14579,N_14425);
or UO_1554 (O_1554,N_14892,N_14929);
and UO_1555 (O_1555,N_14830,N_14581);
nor UO_1556 (O_1556,N_14533,N_14960);
nor UO_1557 (O_1557,N_14602,N_14317);
xnor UO_1558 (O_1558,N_14816,N_14775);
xnor UO_1559 (O_1559,N_14999,N_14655);
nor UO_1560 (O_1560,N_14899,N_14597);
or UO_1561 (O_1561,N_14784,N_14361);
xnor UO_1562 (O_1562,N_14474,N_14798);
nand UO_1563 (O_1563,N_14463,N_14541);
xor UO_1564 (O_1564,N_14913,N_14327);
xnor UO_1565 (O_1565,N_14890,N_14511);
nor UO_1566 (O_1566,N_14449,N_14646);
nand UO_1567 (O_1567,N_14321,N_14657);
xor UO_1568 (O_1568,N_14597,N_14872);
nand UO_1569 (O_1569,N_14596,N_14903);
and UO_1570 (O_1570,N_14507,N_14637);
or UO_1571 (O_1571,N_14514,N_14659);
and UO_1572 (O_1572,N_14628,N_14535);
nand UO_1573 (O_1573,N_14443,N_14326);
or UO_1574 (O_1574,N_14781,N_14402);
nand UO_1575 (O_1575,N_14624,N_14657);
nor UO_1576 (O_1576,N_14353,N_14611);
xnor UO_1577 (O_1577,N_14757,N_14608);
nand UO_1578 (O_1578,N_14603,N_14786);
nand UO_1579 (O_1579,N_14360,N_14583);
nor UO_1580 (O_1580,N_14491,N_14439);
nand UO_1581 (O_1581,N_14273,N_14964);
nand UO_1582 (O_1582,N_14674,N_14818);
xor UO_1583 (O_1583,N_14719,N_14356);
nand UO_1584 (O_1584,N_14267,N_14370);
and UO_1585 (O_1585,N_14615,N_14828);
nor UO_1586 (O_1586,N_14504,N_14384);
and UO_1587 (O_1587,N_14801,N_14293);
and UO_1588 (O_1588,N_14436,N_14442);
nand UO_1589 (O_1589,N_14838,N_14266);
or UO_1590 (O_1590,N_14701,N_14677);
nor UO_1591 (O_1591,N_14331,N_14948);
nor UO_1592 (O_1592,N_14791,N_14582);
xnor UO_1593 (O_1593,N_14629,N_14799);
and UO_1594 (O_1594,N_14536,N_14272);
xor UO_1595 (O_1595,N_14465,N_14511);
and UO_1596 (O_1596,N_14250,N_14829);
nand UO_1597 (O_1597,N_14869,N_14317);
nand UO_1598 (O_1598,N_14328,N_14648);
and UO_1599 (O_1599,N_14620,N_14945);
and UO_1600 (O_1600,N_14392,N_14415);
nor UO_1601 (O_1601,N_14572,N_14665);
and UO_1602 (O_1602,N_14951,N_14428);
nor UO_1603 (O_1603,N_14455,N_14379);
and UO_1604 (O_1604,N_14372,N_14563);
and UO_1605 (O_1605,N_14570,N_14845);
or UO_1606 (O_1606,N_14436,N_14517);
nor UO_1607 (O_1607,N_14435,N_14652);
nor UO_1608 (O_1608,N_14358,N_14368);
or UO_1609 (O_1609,N_14695,N_14376);
nor UO_1610 (O_1610,N_14682,N_14469);
or UO_1611 (O_1611,N_14562,N_14654);
or UO_1612 (O_1612,N_14359,N_14719);
nor UO_1613 (O_1613,N_14719,N_14360);
nand UO_1614 (O_1614,N_14609,N_14347);
or UO_1615 (O_1615,N_14505,N_14562);
or UO_1616 (O_1616,N_14375,N_14842);
nor UO_1617 (O_1617,N_14855,N_14527);
xnor UO_1618 (O_1618,N_14561,N_14419);
or UO_1619 (O_1619,N_14920,N_14876);
xnor UO_1620 (O_1620,N_14916,N_14752);
xor UO_1621 (O_1621,N_14352,N_14312);
and UO_1622 (O_1622,N_14788,N_14901);
or UO_1623 (O_1623,N_14927,N_14252);
nor UO_1624 (O_1624,N_14589,N_14686);
and UO_1625 (O_1625,N_14624,N_14277);
and UO_1626 (O_1626,N_14273,N_14699);
xor UO_1627 (O_1627,N_14697,N_14512);
nor UO_1628 (O_1628,N_14382,N_14393);
nor UO_1629 (O_1629,N_14490,N_14972);
and UO_1630 (O_1630,N_14581,N_14945);
and UO_1631 (O_1631,N_14518,N_14700);
and UO_1632 (O_1632,N_14356,N_14824);
xor UO_1633 (O_1633,N_14461,N_14453);
nand UO_1634 (O_1634,N_14282,N_14362);
nor UO_1635 (O_1635,N_14991,N_14805);
or UO_1636 (O_1636,N_14561,N_14827);
nor UO_1637 (O_1637,N_14825,N_14973);
nand UO_1638 (O_1638,N_14769,N_14417);
or UO_1639 (O_1639,N_14317,N_14699);
xnor UO_1640 (O_1640,N_14873,N_14351);
and UO_1641 (O_1641,N_14948,N_14790);
xor UO_1642 (O_1642,N_14440,N_14528);
or UO_1643 (O_1643,N_14933,N_14360);
or UO_1644 (O_1644,N_14732,N_14725);
or UO_1645 (O_1645,N_14914,N_14576);
xor UO_1646 (O_1646,N_14468,N_14424);
and UO_1647 (O_1647,N_14927,N_14701);
nand UO_1648 (O_1648,N_14470,N_14976);
nor UO_1649 (O_1649,N_14822,N_14506);
nor UO_1650 (O_1650,N_14609,N_14342);
nand UO_1651 (O_1651,N_14617,N_14640);
nor UO_1652 (O_1652,N_14720,N_14703);
and UO_1653 (O_1653,N_14746,N_14811);
nand UO_1654 (O_1654,N_14260,N_14655);
nand UO_1655 (O_1655,N_14652,N_14625);
and UO_1656 (O_1656,N_14572,N_14580);
or UO_1657 (O_1657,N_14875,N_14816);
nand UO_1658 (O_1658,N_14696,N_14703);
nand UO_1659 (O_1659,N_14752,N_14665);
nor UO_1660 (O_1660,N_14939,N_14626);
xor UO_1661 (O_1661,N_14596,N_14939);
xnor UO_1662 (O_1662,N_14375,N_14533);
and UO_1663 (O_1663,N_14928,N_14277);
nand UO_1664 (O_1664,N_14874,N_14711);
or UO_1665 (O_1665,N_14473,N_14380);
nand UO_1666 (O_1666,N_14874,N_14501);
or UO_1667 (O_1667,N_14731,N_14961);
nand UO_1668 (O_1668,N_14262,N_14931);
or UO_1669 (O_1669,N_14848,N_14321);
nor UO_1670 (O_1670,N_14255,N_14899);
xnor UO_1671 (O_1671,N_14337,N_14595);
and UO_1672 (O_1672,N_14397,N_14646);
and UO_1673 (O_1673,N_14820,N_14492);
nand UO_1674 (O_1674,N_14481,N_14338);
nor UO_1675 (O_1675,N_14718,N_14818);
xor UO_1676 (O_1676,N_14642,N_14550);
and UO_1677 (O_1677,N_14647,N_14684);
xor UO_1678 (O_1678,N_14611,N_14847);
nand UO_1679 (O_1679,N_14270,N_14925);
xnor UO_1680 (O_1680,N_14951,N_14378);
xnor UO_1681 (O_1681,N_14503,N_14954);
nor UO_1682 (O_1682,N_14964,N_14826);
nand UO_1683 (O_1683,N_14356,N_14561);
and UO_1684 (O_1684,N_14624,N_14777);
xor UO_1685 (O_1685,N_14988,N_14269);
xnor UO_1686 (O_1686,N_14536,N_14503);
nand UO_1687 (O_1687,N_14680,N_14888);
xnor UO_1688 (O_1688,N_14771,N_14799);
nand UO_1689 (O_1689,N_14393,N_14641);
and UO_1690 (O_1690,N_14986,N_14959);
or UO_1691 (O_1691,N_14450,N_14264);
or UO_1692 (O_1692,N_14363,N_14430);
and UO_1693 (O_1693,N_14879,N_14809);
xor UO_1694 (O_1694,N_14256,N_14437);
nand UO_1695 (O_1695,N_14992,N_14503);
nand UO_1696 (O_1696,N_14700,N_14360);
xor UO_1697 (O_1697,N_14858,N_14998);
nand UO_1698 (O_1698,N_14283,N_14870);
or UO_1699 (O_1699,N_14997,N_14436);
xor UO_1700 (O_1700,N_14703,N_14477);
nor UO_1701 (O_1701,N_14953,N_14816);
xor UO_1702 (O_1702,N_14505,N_14391);
and UO_1703 (O_1703,N_14889,N_14944);
and UO_1704 (O_1704,N_14813,N_14970);
nor UO_1705 (O_1705,N_14703,N_14851);
nor UO_1706 (O_1706,N_14720,N_14944);
xnor UO_1707 (O_1707,N_14998,N_14909);
and UO_1708 (O_1708,N_14822,N_14800);
or UO_1709 (O_1709,N_14300,N_14957);
nand UO_1710 (O_1710,N_14730,N_14542);
or UO_1711 (O_1711,N_14659,N_14674);
nor UO_1712 (O_1712,N_14816,N_14628);
xnor UO_1713 (O_1713,N_14777,N_14311);
nand UO_1714 (O_1714,N_14446,N_14352);
nand UO_1715 (O_1715,N_14501,N_14254);
nor UO_1716 (O_1716,N_14315,N_14570);
nor UO_1717 (O_1717,N_14831,N_14828);
xnor UO_1718 (O_1718,N_14613,N_14755);
nand UO_1719 (O_1719,N_14382,N_14734);
xor UO_1720 (O_1720,N_14578,N_14719);
xnor UO_1721 (O_1721,N_14468,N_14330);
or UO_1722 (O_1722,N_14999,N_14925);
nand UO_1723 (O_1723,N_14335,N_14389);
and UO_1724 (O_1724,N_14891,N_14979);
nand UO_1725 (O_1725,N_14291,N_14567);
xor UO_1726 (O_1726,N_14743,N_14498);
nor UO_1727 (O_1727,N_14957,N_14283);
and UO_1728 (O_1728,N_14799,N_14388);
xor UO_1729 (O_1729,N_14759,N_14659);
or UO_1730 (O_1730,N_14845,N_14978);
nand UO_1731 (O_1731,N_14837,N_14881);
nand UO_1732 (O_1732,N_14921,N_14507);
and UO_1733 (O_1733,N_14255,N_14282);
nor UO_1734 (O_1734,N_14803,N_14919);
nand UO_1735 (O_1735,N_14726,N_14893);
nand UO_1736 (O_1736,N_14734,N_14606);
nor UO_1737 (O_1737,N_14278,N_14473);
and UO_1738 (O_1738,N_14262,N_14748);
xnor UO_1739 (O_1739,N_14964,N_14329);
or UO_1740 (O_1740,N_14761,N_14708);
nand UO_1741 (O_1741,N_14960,N_14468);
nor UO_1742 (O_1742,N_14573,N_14560);
or UO_1743 (O_1743,N_14840,N_14648);
and UO_1744 (O_1744,N_14763,N_14734);
or UO_1745 (O_1745,N_14723,N_14905);
nor UO_1746 (O_1746,N_14299,N_14897);
nor UO_1747 (O_1747,N_14866,N_14577);
and UO_1748 (O_1748,N_14281,N_14355);
or UO_1749 (O_1749,N_14336,N_14600);
nand UO_1750 (O_1750,N_14346,N_14377);
xor UO_1751 (O_1751,N_14875,N_14550);
and UO_1752 (O_1752,N_14500,N_14475);
and UO_1753 (O_1753,N_14544,N_14699);
nand UO_1754 (O_1754,N_14781,N_14370);
or UO_1755 (O_1755,N_14748,N_14459);
and UO_1756 (O_1756,N_14972,N_14529);
xor UO_1757 (O_1757,N_14305,N_14650);
nor UO_1758 (O_1758,N_14909,N_14758);
or UO_1759 (O_1759,N_14804,N_14972);
or UO_1760 (O_1760,N_14315,N_14646);
and UO_1761 (O_1761,N_14529,N_14592);
nand UO_1762 (O_1762,N_14362,N_14829);
and UO_1763 (O_1763,N_14479,N_14515);
nand UO_1764 (O_1764,N_14355,N_14713);
and UO_1765 (O_1765,N_14497,N_14872);
and UO_1766 (O_1766,N_14399,N_14735);
or UO_1767 (O_1767,N_14435,N_14904);
and UO_1768 (O_1768,N_14367,N_14510);
or UO_1769 (O_1769,N_14481,N_14518);
nor UO_1770 (O_1770,N_14458,N_14630);
and UO_1771 (O_1771,N_14325,N_14720);
or UO_1772 (O_1772,N_14815,N_14766);
or UO_1773 (O_1773,N_14863,N_14857);
nand UO_1774 (O_1774,N_14392,N_14535);
and UO_1775 (O_1775,N_14897,N_14620);
nor UO_1776 (O_1776,N_14687,N_14962);
or UO_1777 (O_1777,N_14428,N_14837);
xnor UO_1778 (O_1778,N_14614,N_14391);
nand UO_1779 (O_1779,N_14897,N_14704);
nand UO_1780 (O_1780,N_14426,N_14771);
xnor UO_1781 (O_1781,N_14635,N_14270);
nor UO_1782 (O_1782,N_14860,N_14567);
and UO_1783 (O_1783,N_14842,N_14379);
nand UO_1784 (O_1784,N_14800,N_14559);
or UO_1785 (O_1785,N_14542,N_14297);
nand UO_1786 (O_1786,N_14525,N_14569);
or UO_1787 (O_1787,N_14568,N_14926);
and UO_1788 (O_1788,N_14597,N_14803);
nand UO_1789 (O_1789,N_14606,N_14923);
xor UO_1790 (O_1790,N_14453,N_14664);
or UO_1791 (O_1791,N_14347,N_14770);
xor UO_1792 (O_1792,N_14812,N_14681);
nand UO_1793 (O_1793,N_14806,N_14565);
xnor UO_1794 (O_1794,N_14949,N_14429);
or UO_1795 (O_1795,N_14945,N_14952);
or UO_1796 (O_1796,N_14648,N_14344);
and UO_1797 (O_1797,N_14666,N_14680);
xnor UO_1798 (O_1798,N_14438,N_14702);
and UO_1799 (O_1799,N_14574,N_14718);
and UO_1800 (O_1800,N_14998,N_14398);
xnor UO_1801 (O_1801,N_14299,N_14978);
nand UO_1802 (O_1802,N_14945,N_14723);
nor UO_1803 (O_1803,N_14464,N_14991);
xnor UO_1804 (O_1804,N_14276,N_14593);
and UO_1805 (O_1805,N_14905,N_14679);
or UO_1806 (O_1806,N_14277,N_14474);
nand UO_1807 (O_1807,N_14828,N_14628);
and UO_1808 (O_1808,N_14373,N_14289);
nor UO_1809 (O_1809,N_14885,N_14512);
nand UO_1810 (O_1810,N_14614,N_14469);
xor UO_1811 (O_1811,N_14863,N_14865);
or UO_1812 (O_1812,N_14293,N_14978);
and UO_1813 (O_1813,N_14543,N_14664);
nand UO_1814 (O_1814,N_14623,N_14919);
or UO_1815 (O_1815,N_14430,N_14767);
or UO_1816 (O_1816,N_14540,N_14567);
nor UO_1817 (O_1817,N_14635,N_14443);
xnor UO_1818 (O_1818,N_14307,N_14809);
and UO_1819 (O_1819,N_14943,N_14873);
and UO_1820 (O_1820,N_14715,N_14635);
or UO_1821 (O_1821,N_14845,N_14402);
nand UO_1822 (O_1822,N_14804,N_14644);
nor UO_1823 (O_1823,N_14582,N_14833);
nand UO_1824 (O_1824,N_14442,N_14539);
xor UO_1825 (O_1825,N_14464,N_14446);
nand UO_1826 (O_1826,N_14329,N_14999);
xnor UO_1827 (O_1827,N_14808,N_14252);
and UO_1828 (O_1828,N_14966,N_14959);
xor UO_1829 (O_1829,N_14378,N_14366);
nand UO_1830 (O_1830,N_14664,N_14269);
xor UO_1831 (O_1831,N_14468,N_14739);
xnor UO_1832 (O_1832,N_14681,N_14328);
nor UO_1833 (O_1833,N_14660,N_14943);
xor UO_1834 (O_1834,N_14899,N_14442);
nor UO_1835 (O_1835,N_14769,N_14353);
nor UO_1836 (O_1836,N_14980,N_14930);
and UO_1837 (O_1837,N_14257,N_14986);
nor UO_1838 (O_1838,N_14495,N_14617);
nand UO_1839 (O_1839,N_14592,N_14565);
nor UO_1840 (O_1840,N_14803,N_14666);
or UO_1841 (O_1841,N_14759,N_14615);
or UO_1842 (O_1842,N_14372,N_14466);
and UO_1843 (O_1843,N_14261,N_14392);
nand UO_1844 (O_1844,N_14696,N_14840);
nand UO_1845 (O_1845,N_14331,N_14841);
nand UO_1846 (O_1846,N_14948,N_14788);
nor UO_1847 (O_1847,N_14641,N_14528);
nor UO_1848 (O_1848,N_14765,N_14454);
xor UO_1849 (O_1849,N_14655,N_14916);
xor UO_1850 (O_1850,N_14965,N_14832);
xor UO_1851 (O_1851,N_14662,N_14514);
nor UO_1852 (O_1852,N_14347,N_14504);
nor UO_1853 (O_1853,N_14686,N_14569);
nor UO_1854 (O_1854,N_14949,N_14627);
nand UO_1855 (O_1855,N_14610,N_14576);
nand UO_1856 (O_1856,N_14469,N_14741);
or UO_1857 (O_1857,N_14702,N_14758);
nor UO_1858 (O_1858,N_14372,N_14780);
nand UO_1859 (O_1859,N_14332,N_14616);
and UO_1860 (O_1860,N_14487,N_14703);
xnor UO_1861 (O_1861,N_14800,N_14788);
or UO_1862 (O_1862,N_14470,N_14416);
xor UO_1863 (O_1863,N_14394,N_14643);
nand UO_1864 (O_1864,N_14563,N_14322);
nand UO_1865 (O_1865,N_14644,N_14483);
nand UO_1866 (O_1866,N_14338,N_14253);
nand UO_1867 (O_1867,N_14280,N_14424);
or UO_1868 (O_1868,N_14680,N_14412);
or UO_1869 (O_1869,N_14677,N_14260);
and UO_1870 (O_1870,N_14837,N_14435);
nand UO_1871 (O_1871,N_14679,N_14727);
nor UO_1872 (O_1872,N_14538,N_14554);
nand UO_1873 (O_1873,N_14919,N_14273);
or UO_1874 (O_1874,N_14322,N_14451);
xnor UO_1875 (O_1875,N_14601,N_14273);
or UO_1876 (O_1876,N_14530,N_14973);
xnor UO_1877 (O_1877,N_14280,N_14604);
nor UO_1878 (O_1878,N_14387,N_14502);
nand UO_1879 (O_1879,N_14500,N_14724);
nor UO_1880 (O_1880,N_14395,N_14469);
nor UO_1881 (O_1881,N_14782,N_14806);
and UO_1882 (O_1882,N_14522,N_14273);
or UO_1883 (O_1883,N_14572,N_14748);
nand UO_1884 (O_1884,N_14871,N_14942);
nor UO_1885 (O_1885,N_14951,N_14775);
nor UO_1886 (O_1886,N_14554,N_14666);
and UO_1887 (O_1887,N_14295,N_14670);
and UO_1888 (O_1888,N_14391,N_14913);
or UO_1889 (O_1889,N_14994,N_14330);
or UO_1890 (O_1890,N_14544,N_14327);
xor UO_1891 (O_1891,N_14381,N_14259);
or UO_1892 (O_1892,N_14723,N_14395);
or UO_1893 (O_1893,N_14754,N_14579);
nor UO_1894 (O_1894,N_14964,N_14401);
and UO_1895 (O_1895,N_14788,N_14728);
and UO_1896 (O_1896,N_14716,N_14450);
and UO_1897 (O_1897,N_14304,N_14998);
xor UO_1898 (O_1898,N_14951,N_14364);
or UO_1899 (O_1899,N_14982,N_14808);
or UO_1900 (O_1900,N_14283,N_14319);
and UO_1901 (O_1901,N_14467,N_14361);
and UO_1902 (O_1902,N_14956,N_14286);
nand UO_1903 (O_1903,N_14456,N_14827);
nor UO_1904 (O_1904,N_14830,N_14993);
or UO_1905 (O_1905,N_14608,N_14408);
and UO_1906 (O_1906,N_14419,N_14596);
or UO_1907 (O_1907,N_14836,N_14273);
nand UO_1908 (O_1908,N_14691,N_14615);
and UO_1909 (O_1909,N_14483,N_14784);
nand UO_1910 (O_1910,N_14632,N_14469);
nor UO_1911 (O_1911,N_14867,N_14559);
nand UO_1912 (O_1912,N_14403,N_14632);
xnor UO_1913 (O_1913,N_14991,N_14986);
nor UO_1914 (O_1914,N_14763,N_14520);
nand UO_1915 (O_1915,N_14431,N_14941);
and UO_1916 (O_1916,N_14653,N_14282);
and UO_1917 (O_1917,N_14333,N_14692);
nand UO_1918 (O_1918,N_14936,N_14281);
and UO_1919 (O_1919,N_14793,N_14690);
xnor UO_1920 (O_1920,N_14258,N_14597);
xnor UO_1921 (O_1921,N_14635,N_14834);
nor UO_1922 (O_1922,N_14607,N_14811);
or UO_1923 (O_1923,N_14703,N_14261);
xnor UO_1924 (O_1924,N_14950,N_14695);
or UO_1925 (O_1925,N_14511,N_14612);
nand UO_1926 (O_1926,N_14413,N_14341);
or UO_1927 (O_1927,N_14930,N_14385);
nand UO_1928 (O_1928,N_14423,N_14587);
and UO_1929 (O_1929,N_14576,N_14260);
nand UO_1930 (O_1930,N_14588,N_14909);
nand UO_1931 (O_1931,N_14474,N_14682);
and UO_1932 (O_1932,N_14558,N_14587);
nand UO_1933 (O_1933,N_14625,N_14296);
and UO_1934 (O_1934,N_14678,N_14533);
or UO_1935 (O_1935,N_14743,N_14745);
xor UO_1936 (O_1936,N_14504,N_14260);
and UO_1937 (O_1937,N_14608,N_14847);
xor UO_1938 (O_1938,N_14470,N_14912);
nor UO_1939 (O_1939,N_14765,N_14525);
xor UO_1940 (O_1940,N_14997,N_14761);
xor UO_1941 (O_1941,N_14299,N_14667);
xnor UO_1942 (O_1942,N_14255,N_14893);
and UO_1943 (O_1943,N_14586,N_14696);
and UO_1944 (O_1944,N_14436,N_14425);
and UO_1945 (O_1945,N_14900,N_14707);
xor UO_1946 (O_1946,N_14444,N_14737);
and UO_1947 (O_1947,N_14675,N_14917);
and UO_1948 (O_1948,N_14308,N_14503);
or UO_1949 (O_1949,N_14309,N_14511);
and UO_1950 (O_1950,N_14587,N_14957);
nor UO_1951 (O_1951,N_14858,N_14888);
and UO_1952 (O_1952,N_14420,N_14961);
or UO_1953 (O_1953,N_14565,N_14509);
nand UO_1954 (O_1954,N_14919,N_14452);
or UO_1955 (O_1955,N_14896,N_14589);
and UO_1956 (O_1956,N_14923,N_14910);
nand UO_1957 (O_1957,N_14494,N_14787);
nor UO_1958 (O_1958,N_14659,N_14554);
nor UO_1959 (O_1959,N_14256,N_14592);
or UO_1960 (O_1960,N_14756,N_14793);
xnor UO_1961 (O_1961,N_14975,N_14974);
and UO_1962 (O_1962,N_14734,N_14794);
xnor UO_1963 (O_1963,N_14518,N_14767);
and UO_1964 (O_1964,N_14913,N_14307);
xnor UO_1965 (O_1965,N_14600,N_14797);
xor UO_1966 (O_1966,N_14695,N_14775);
nand UO_1967 (O_1967,N_14331,N_14284);
nor UO_1968 (O_1968,N_14368,N_14987);
or UO_1969 (O_1969,N_14484,N_14927);
or UO_1970 (O_1970,N_14289,N_14747);
nand UO_1971 (O_1971,N_14515,N_14986);
or UO_1972 (O_1972,N_14365,N_14307);
nand UO_1973 (O_1973,N_14291,N_14640);
nand UO_1974 (O_1974,N_14426,N_14787);
nand UO_1975 (O_1975,N_14659,N_14594);
xor UO_1976 (O_1976,N_14251,N_14914);
or UO_1977 (O_1977,N_14894,N_14913);
nor UO_1978 (O_1978,N_14911,N_14797);
or UO_1979 (O_1979,N_14346,N_14693);
and UO_1980 (O_1980,N_14970,N_14982);
nor UO_1981 (O_1981,N_14610,N_14946);
and UO_1982 (O_1982,N_14342,N_14534);
xor UO_1983 (O_1983,N_14535,N_14979);
nor UO_1984 (O_1984,N_14739,N_14697);
or UO_1985 (O_1985,N_14876,N_14739);
or UO_1986 (O_1986,N_14617,N_14813);
and UO_1987 (O_1987,N_14315,N_14590);
or UO_1988 (O_1988,N_14548,N_14911);
nand UO_1989 (O_1989,N_14397,N_14982);
nand UO_1990 (O_1990,N_14278,N_14570);
nand UO_1991 (O_1991,N_14668,N_14711);
nor UO_1992 (O_1992,N_14857,N_14762);
nor UO_1993 (O_1993,N_14976,N_14635);
nor UO_1994 (O_1994,N_14528,N_14628);
and UO_1995 (O_1995,N_14583,N_14868);
nor UO_1996 (O_1996,N_14911,N_14618);
and UO_1997 (O_1997,N_14839,N_14448);
xnor UO_1998 (O_1998,N_14745,N_14333);
nor UO_1999 (O_1999,N_14472,N_14900);
endmodule