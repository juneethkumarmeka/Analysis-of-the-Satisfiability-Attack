module basic_500_3000_500_5_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_115,In_91);
nand U1 (N_1,In_74,In_46);
nor U2 (N_2,In_223,In_194);
or U3 (N_3,In_459,In_295);
nor U4 (N_4,In_259,In_362);
xor U5 (N_5,In_449,In_275);
nor U6 (N_6,In_492,In_483);
nor U7 (N_7,In_11,In_25);
nor U8 (N_8,In_388,In_28);
nor U9 (N_9,In_370,In_340);
or U10 (N_10,In_256,In_88);
or U11 (N_11,In_489,In_135);
nand U12 (N_12,In_393,In_382);
nor U13 (N_13,In_157,In_389);
nand U14 (N_14,In_493,In_298);
or U15 (N_15,In_161,In_238);
and U16 (N_16,In_211,In_243);
nor U17 (N_17,In_54,In_479);
and U18 (N_18,In_332,In_284);
nand U19 (N_19,In_212,In_222);
nor U20 (N_20,In_187,In_499);
nand U21 (N_21,In_267,In_113);
or U22 (N_22,In_443,In_354);
or U23 (N_23,In_90,In_159);
nand U24 (N_24,In_346,In_55);
nand U25 (N_25,In_283,In_162);
xor U26 (N_26,In_359,In_109);
and U27 (N_27,In_118,In_53);
or U28 (N_28,In_77,In_40);
and U29 (N_29,In_179,In_271);
nor U30 (N_30,In_35,In_152);
nor U31 (N_31,In_117,In_232);
and U32 (N_32,In_425,In_444);
or U33 (N_33,In_254,In_0);
nand U34 (N_34,In_186,In_349);
nand U35 (N_35,In_430,In_305);
nor U36 (N_36,In_96,In_148);
or U37 (N_37,In_233,In_155);
nand U38 (N_38,In_182,In_355);
and U39 (N_39,In_178,In_381);
and U40 (N_40,In_323,In_468);
or U41 (N_41,In_282,In_228);
nor U42 (N_42,In_438,In_239);
xor U43 (N_43,In_318,In_201);
and U44 (N_44,In_312,In_268);
nand U45 (N_45,In_94,In_79);
and U46 (N_46,In_445,In_313);
nand U47 (N_47,In_151,In_81);
or U48 (N_48,In_202,In_5);
and U49 (N_49,In_276,In_361);
and U50 (N_50,In_423,In_487);
or U51 (N_51,In_221,In_420);
nor U52 (N_52,In_21,In_171);
nor U53 (N_53,In_336,In_266);
nand U54 (N_54,In_291,In_408);
nor U55 (N_55,In_101,In_396);
xor U56 (N_56,In_435,In_30);
or U57 (N_57,In_341,In_22);
and U58 (N_58,In_378,In_10);
and U59 (N_59,In_24,In_39);
nand U60 (N_60,In_188,In_411);
and U61 (N_61,In_472,In_263);
or U62 (N_62,In_484,In_87);
or U63 (N_63,In_288,In_33);
and U64 (N_64,In_17,In_92);
or U65 (N_65,In_415,In_216);
or U66 (N_66,In_432,In_251);
nor U67 (N_67,In_153,In_235);
or U68 (N_68,In_156,In_429);
nand U69 (N_69,In_246,In_36);
xor U70 (N_70,In_441,In_392);
or U71 (N_71,In_121,In_304);
and U72 (N_72,In_12,In_130);
xnor U73 (N_73,In_486,In_352);
nor U74 (N_74,In_71,In_245);
xnor U75 (N_75,In_103,In_20);
and U76 (N_76,In_37,In_398);
or U77 (N_77,In_350,In_19);
nor U78 (N_78,In_287,In_66);
or U79 (N_79,In_200,In_124);
nor U80 (N_80,In_248,In_437);
nor U81 (N_81,In_448,In_427);
and U82 (N_82,In_440,In_456);
and U83 (N_83,In_100,In_401);
and U84 (N_84,In_102,In_250);
or U85 (N_85,In_62,In_466);
xor U86 (N_86,In_139,In_150);
and U87 (N_87,In_405,In_72);
and U88 (N_88,In_460,In_457);
nand U89 (N_89,In_439,In_49);
or U90 (N_90,In_442,In_120);
or U91 (N_91,In_368,In_369);
and U92 (N_92,In_281,In_183);
xor U93 (N_93,In_122,In_253);
and U94 (N_94,In_390,In_67);
nand U95 (N_95,In_126,In_98);
nor U96 (N_96,In_70,In_6);
and U97 (N_97,In_86,In_197);
and U98 (N_98,In_321,In_106);
or U99 (N_99,In_317,In_131);
xnor U100 (N_100,In_63,In_351);
or U101 (N_101,In_365,In_99);
and U102 (N_102,In_230,In_480);
nand U103 (N_103,In_301,In_132);
nand U104 (N_104,In_7,In_3);
or U105 (N_105,In_44,In_315);
nor U106 (N_106,In_15,In_112);
nor U107 (N_107,In_454,In_82);
or U108 (N_108,In_60,In_488);
nor U109 (N_109,In_470,In_136);
nor U110 (N_110,In_145,In_164);
xnor U111 (N_111,In_335,In_142);
and U112 (N_112,In_129,In_261);
nand U113 (N_113,In_342,In_47);
nand U114 (N_114,In_134,In_83);
nand U115 (N_115,In_296,In_140);
or U116 (N_116,In_462,In_363);
nor U117 (N_117,In_203,In_147);
and U118 (N_118,In_114,In_289);
nand U119 (N_119,In_292,In_307);
nor U120 (N_120,In_137,In_476);
nand U121 (N_121,In_8,In_177);
or U122 (N_122,In_310,In_377);
nand U123 (N_123,In_34,In_208);
or U124 (N_124,In_417,In_174);
nand U125 (N_125,In_185,In_302);
or U126 (N_126,In_229,In_219);
nor U127 (N_127,In_144,In_399);
and U128 (N_128,In_224,In_421);
and U129 (N_129,In_226,In_13);
nor U130 (N_130,In_311,In_277);
nor U131 (N_131,In_149,In_84);
nand U132 (N_132,In_218,In_234);
nor U133 (N_133,In_196,In_204);
and U134 (N_134,In_165,In_241);
or U135 (N_135,In_426,In_104);
nor U136 (N_136,In_303,In_56);
and U137 (N_137,In_29,In_394);
nand U138 (N_138,In_257,In_357);
and U139 (N_139,In_481,In_400);
xor U140 (N_140,In_331,In_14);
and U141 (N_141,In_364,In_308);
or U142 (N_142,In_416,In_294);
xor U143 (N_143,In_265,In_347);
nand U144 (N_144,In_309,In_469);
xnor U145 (N_145,In_57,In_41);
or U146 (N_146,In_58,In_299);
nor U147 (N_147,In_372,In_371);
or U148 (N_148,In_85,In_451);
nor U149 (N_149,In_403,In_45);
xnor U150 (N_150,In_333,In_89);
nor U151 (N_151,In_498,In_475);
and U152 (N_152,In_409,In_367);
nand U153 (N_153,In_97,In_477);
nand U154 (N_154,In_279,In_119);
xnor U155 (N_155,In_192,In_463);
nand U156 (N_156,In_206,In_376);
nand U157 (N_157,In_193,In_348);
and U158 (N_158,In_184,In_328);
xnor U159 (N_159,In_80,In_1);
and U160 (N_160,In_455,In_384);
and U161 (N_161,In_31,In_76);
or U162 (N_162,In_320,In_181);
or U163 (N_163,In_107,In_494);
nor U164 (N_164,In_464,In_434);
xor U165 (N_165,In_240,In_32);
xnor U166 (N_166,In_141,In_418);
or U167 (N_167,In_339,In_2);
and U168 (N_168,In_190,In_269);
xnor U169 (N_169,In_436,In_446);
and U170 (N_170,In_412,In_64);
or U171 (N_171,In_326,In_458);
nand U172 (N_172,In_258,In_207);
or U173 (N_173,In_387,In_293);
and U174 (N_174,In_297,In_123);
nor U175 (N_175,In_18,In_375);
or U176 (N_176,In_490,In_48);
and U177 (N_177,In_314,In_272);
nand U178 (N_178,In_158,In_474);
xor U179 (N_179,In_497,In_495);
nand U180 (N_180,In_236,In_419);
and U181 (N_181,In_461,In_59);
xnor U182 (N_182,In_385,In_38);
or U183 (N_183,In_225,In_338);
nor U184 (N_184,In_356,In_395);
or U185 (N_185,In_379,In_199);
and U186 (N_186,In_397,In_337);
nor U187 (N_187,In_127,In_478);
or U188 (N_188,In_273,In_146);
nor U189 (N_189,In_386,In_324);
nand U190 (N_190,In_231,In_260);
nand U191 (N_191,In_374,In_249);
nor U192 (N_192,In_402,In_4);
xnor U193 (N_193,In_110,In_215);
or U194 (N_194,In_26,In_467);
or U195 (N_195,In_280,In_93);
xor U196 (N_196,In_78,In_69);
xor U197 (N_197,In_343,In_143);
nor U198 (N_198,In_61,In_496);
nand U199 (N_199,In_111,In_406);
or U200 (N_200,In_452,In_205);
xor U201 (N_201,In_264,In_168);
and U202 (N_202,In_220,In_50);
nand U203 (N_203,In_353,In_471);
or U204 (N_204,In_431,In_176);
or U205 (N_205,In_278,In_209);
xor U206 (N_206,In_65,In_175);
and U207 (N_207,In_485,In_491);
or U208 (N_208,In_105,In_16);
nand U209 (N_209,In_422,In_198);
or U210 (N_210,In_173,In_237);
or U211 (N_211,In_217,In_9);
nor U212 (N_212,In_270,In_383);
xor U213 (N_213,In_255,In_380);
nor U214 (N_214,In_330,In_154);
or U215 (N_215,In_213,In_170);
and U216 (N_216,In_160,In_95);
xnor U217 (N_217,In_358,In_482);
and U218 (N_218,In_108,In_242);
nand U219 (N_219,In_172,In_290);
and U220 (N_220,In_163,In_465);
nand U221 (N_221,In_391,In_75);
or U222 (N_222,In_138,In_428);
xnor U223 (N_223,In_128,In_407);
or U224 (N_224,In_210,In_68);
nand U225 (N_225,In_334,In_306);
nor U226 (N_226,In_125,In_191);
nor U227 (N_227,In_42,In_189);
nor U228 (N_228,In_116,In_169);
and U229 (N_229,In_360,In_447);
nor U230 (N_230,In_453,In_319);
xor U231 (N_231,In_366,In_450);
and U232 (N_232,In_286,In_413);
and U233 (N_233,In_27,In_166);
or U234 (N_234,In_227,In_316);
nand U235 (N_235,In_327,In_133);
and U236 (N_236,In_180,In_274);
nand U237 (N_237,In_404,In_410);
nor U238 (N_238,In_322,In_325);
nor U239 (N_239,In_195,In_247);
nor U240 (N_240,In_345,In_167);
and U241 (N_241,In_43,In_344);
nand U242 (N_242,In_262,In_424);
or U243 (N_243,In_52,In_23);
nand U244 (N_244,In_73,In_244);
and U245 (N_245,In_414,In_252);
or U246 (N_246,In_214,In_51);
and U247 (N_247,In_373,In_285);
nor U248 (N_248,In_329,In_473);
xor U249 (N_249,In_433,In_300);
and U250 (N_250,In_189,In_239);
nor U251 (N_251,In_155,In_356);
or U252 (N_252,In_383,In_279);
nor U253 (N_253,In_320,In_147);
nand U254 (N_254,In_60,In_245);
nor U255 (N_255,In_494,In_164);
nand U256 (N_256,In_163,In_15);
nand U257 (N_257,In_50,In_329);
and U258 (N_258,In_114,In_275);
nor U259 (N_259,In_253,In_218);
nor U260 (N_260,In_289,In_30);
and U261 (N_261,In_245,In_413);
or U262 (N_262,In_325,In_283);
and U263 (N_263,In_183,In_163);
and U264 (N_264,In_267,In_418);
nor U265 (N_265,In_451,In_100);
nand U266 (N_266,In_448,In_19);
or U267 (N_267,In_79,In_380);
nand U268 (N_268,In_301,In_313);
or U269 (N_269,In_95,In_19);
xor U270 (N_270,In_280,In_15);
xnor U271 (N_271,In_133,In_124);
nand U272 (N_272,In_436,In_399);
or U273 (N_273,In_217,In_86);
nor U274 (N_274,In_335,In_195);
and U275 (N_275,In_114,In_38);
nand U276 (N_276,In_232,In_336);
and U277 (N_277,In_298,In_331);
and U278 (N_278,In_435,In_317);
nor U279 (N_279,In_381,In_292);
nor U280 (N_280,In_477,In_124);
and U281 (N_281,In_411,In_161);
or U282 (N_282,In_433,In_313);
nand U283 (N_283,In_283,In_437);
or U284 (N_284,In_364,In_170);
xor U285 (N_285,In_292,In_302);
nand U286 (N_286,In_497,In_291);
or U287 (N_287,In_459,In_209);
xor U288 (N_288,In_150,In_301);
and U289 (N_289,In_211,In_328);
or U290 (N_290,In_294,In_133);
xnor U291 (N_291,In_5,In_369);
xnor U292 (N_292,In_456,In_66);
and U293 (N_293,In_244,In_66);
or U294 (N_294,In_456,In_275);
or U295 (N_295,In_181,In_65);
nand U296 (N_296,In_321,In_275);
nor U297 (N_297,In_364,In_47);
nor U298 (N_298,In_162,In_312);
nor U299 (N_299,In_221,In_479);
or U300 (N_300,In_464,In_23);
nand U301 (N_301,In_485,In_142);
or U302 (N_302,In_45,In_102);
nand U303 (N_303,In_67,In_298);
nor U304 (N_304,In_395,In_2);
nor U305 (N_305,In_56,In_205);
and U306 (N_306,In_459,In_187);
and U307 (N_307,In_219,In_8);
xor U308 (N_308,In_253,In_181);
nor U309 (N_309,In_367,In_65);
and U310 (N_310,In_406,In_81);
or U311 (N_311,In_469,In_128);
nor U312 (N_312,In_1,In_478);
nor U313 (N_313,In_353,In_454);
or U314 (N_314,In_247,In_99);
nand U315 (N_315,In_104,In_23);
or U316 (N_316,In_243,In_43);
and U317 (N_317,In_495,In_15);
or U318 (N_318,In_14,In_74);
nand U319 (N_319,In_175,In_341);
or U320 (N_320,In_122,In_39);
or U321 (N_321,In_0,In_59);
nor U322 (N_322,In_31,In_412);
or U323 (N_323,In_259,In_481);
and U324 (N_324,In_211,In_147);
nand U325 (N_325,In_203,In_56);
nor U326 (N_326,In_456,In_234);
nor U327 (N_327,In_393,In_292);
or U328 (N_328,In_205,In_336);
xor U329 (N_329,In_496,In_481);
nor U330 (N_330,In_207,In_105);
nand U331 (N_331,In_201,In_161);
nand U332 (N_332,In_380,In_403);
nand U333 (N_333,In_374,In_497);
and U334 (N_334,In_111,In_110);
and U335 (N_335,In_214,In_410);
nand U336 (N_336,In_139,In_272);
or U337 (N_337,In_6,In_361);
nand U338 (N_338,In_377,In_348);
xor U339 (N_339,In_487,In_404);
nand U340 (N_340,In_98,In_191);
or U341 (N_341,In_404,In_74);
and U342 (N_342,In_321,In_308);
nor U343 (N_343,In_379,In_39);
or U344 (N_344,In_255,In_332);
and U345 (N_345,In_84,In_431);
or U346 (N_346,In_1,In_146);
or U347 (N_347,In_61,In_63);
nand U348 (N_348,In_430,In_132);
or U349 (N_349,In_2,In_204);
or U350 (N_350,In_267,In_30);
nor U351 (N_351,In_159,In_167);
or U352 (N_352,In_495,In_486);
nand U353 (N_353,In_102,In_273);
nand U354 (N_354,In_152,In_20);
nor U355 (N_355,In_152,In_108);
nand U356 (N_356,In_325,In_28);
nor U357 (N_357,In_471,In_129);
or U358 (N_358,In_264,In_99);
nand U359 (N_359,In_85,In_12);
nand U360 (N_360,In_118,In_393);
nor U361 (N_361,In_223,In_417);
nor U362 (N_362,In_30,In_64);
nor U363 (N_363,In_232,In_267);
nand U364 (N_364,In_397,In_498);
or U365 (N_365,In_185,In_41);
xnor U366 (N_366,In_88,In_276);
or U367 (N_367,In_348,In_184);
nor U368 (N_368,In_66,In_260);
or U369 (N_369,In_55,In_44);
or U370 (N_370,In_395,In_450);
and U371 (N_371,In_377,In_109);
nand U372 (N_372,In_169,In_317);
nor U373 (N_373,In_19,In_17);
nor U374 (N_374,In_24,In_239);
or U375 (N_375,In_67,In_36);
nand U376 (N_376,In_270,In_135);
or U377 (N_377,In_451,In_326);
nand U378 (N_378,In_391,In_15);
nand U379 (N_379,In_407,In_146);
and U380 (N_380,In_446,In_282);
nand U381 (N_381,In_439,In_184);
nand U382 (N_382,In_366,In_13);
xor U383 (N_383,In_345,In_242);
and U384 (N_384,In_9,In_66);
xor U385 (N_385,In_332,In_45);
or U386 (N_386,In_440,In_143);
nand U387 (N_387,In_287,In_375);
or U388 (N_388,In_447,In_1);
nand U389 (N_389,In_383,In_231);
and U390 (N_390,In_410,In_473);
or U391 (N_391,In_262,In_120);
nand U392 (N_392,In_405,In_343);
nand U393 (N_393,In_474,In_380);
or U394 (N_394,In_128,In_19);
or U395 (N_395,In_380,In_383);
and U396 (N_396,In_255,In_51);
nor U397 (N_397,In_262,In_188);
xnor U398 (N_398,In_22,In_338);
or U399 (N_399,In_55,In_239);
or U400 (N_400,In_269,In_168);
or U401 (N_401,In_370,In_133);
nand U402 (N_402,In_177,In_98);
xnor U403 (N_403,In_352,In_198);
or U404 (N_404,In_351,In_381);
nand U405 (N_405,In_351,In_48);
and U406 (N_406,In_216,In_68);
and U407 (N_407,In_6,In_489);
or U408 (N_408,In_87,In_451);
xnor U409 (N_409,In_497,In_165);
and U410 (N_410,In_322,In_167);
nand U411 (N_411,In_231,In_62);
nor U412 (N_412,In_94,In_370);
nor U413 (N_413,In_60,In_153);
nor U414 (N_414,In_233,In_98);
nor U415 (N_415,In_202,In_341);
nand U416 (N_416,In_53,In_156);
nor U417 (N_417,In_141,In_327);
nor U418 (N_418,In_469,In_362);
or U419 (N_419,In_87,In_353);
and U420 (N_420,In_94,In_83);
or U421 (N_421,In_411,In_244);
nand U422 (N_422,In_307,In_370);
nand U423 (N_423,In_147,In_110);
nand U424 (N_424,In_354,In_225);
nor U425 (N_425,In_228,In_258);
nor U426 (N_426,In_246,In_482);
and U427 (N_427,In_45,In_85);
and U428 (N_428,In_78,In_152);
or U429 (N_429,In_106,In_365);
and U430 (N_430,In_405,In_313);
xor U431 (N_431,In_380,In_210);
and U432 (N_432,In_250,In_345);
or U433 (N_433,In_226,In_260);
nand U434 (N_434,In_22,In_163);
or U435 (N_435,In_228,In_303);
and U436 (N_436,In_220,In_62);
or U437 (N_437,In_122,In_109);
and U438 (N_438,In_196,In_77);
and U439 (N_439,In_81,In_138);
or U440 (N_440,In_424,In_397);
nand U441 (N_441,In_405,In_23);
nand U442 (N_442,In_89,In_415);
nand U443 (N_443,In_433,In_268);
nand U444 (N_444,In_42,In_494);
nor U445 (N_445,In_498,In_424);
nand U446 (N_446,In_366,In_118);
nand U447 (N_447,In_496,In_448);
nand U448 (N_448,In_289,In_470);
or U449 (N_449,In_373,In_415);
or U450 (N_450,In_34,In_352);
or U451 (N_451,In_269,In_33);
or U452 (N_452,In_424,In_43);
nor U453 (N_453,In_421,In_371);
xor U454 (N_454,In_240,In_219);
and U455 (N_455,In_157,In_188);
nor U456 (N_456,In_121,In_109);
or U457 (N_457,In_158,In_219);
and U458 (N_458,In_495,In_163);
and U459 (N_459,In_212,In_56);
xor U460 (N_460,In_196,In_280);
nand U461 (N_461,In_450,In_67);
nand U462 (N_462,In_338,In_315);
and U463 (N_463,In_50,In_298);
xor U464 (N_464,In_177,In_93);
xor U465 (N_465,In_65,In_66);
or U466 (N_466,In_23,In_303);
nand U467 (N_467,In_498,In_77);
and U468 (N_468,In_336,In_364);
nand U469 (N_469,In_161,In_266);
or U470 (N_470,In_318,In_235);
nand U471 (N_471,In_52,In_375);
nor U472 (N_472,In_261,In_331);
xor U473 (N_473,In_279,In_396);
and U474 (N_474,In_197,In_85);
or U475 (N_475,In_244,In_347);
nor U476 (N_476,In_23,In_407);
xor U477 (N_477,In_429,In_61);
and U478 (N_478,In_177,In_304);
and U479 (N_479,In_462,In_359);
or U480 (N_480,In_144,In_320);
nand U481 (N_481,In_50,In_386);
and U482 (N_482,In_342,In_257);
nor U483 (N_483,In_270,In_96);
and U484 (N_484,In_118,In_91);
nor U485 (N_485,In_42,In_401);
or U486 (N_486,In_286,In_365);
nor U487 (N_487,In_422,In_256);
xnor U488 (N_488,In_101,In_172);
or U489 (N_489,In_469,In_45);
nand U490 (N_490,In_58,In_205);
and U491 (N_491,In_369,In_358);
nor U492 (N_492,In_16,In_143);
nand U493 (N_493,In_239,In_331);
and U494 (N_494,In_127,In_235);
or U495 (N_495,In_163,In_301);
and U496 (N_496,In_176,In_131);
and U497 (N_497,In_92,In_178);
and U498 (N_498,In_193,In_270);
and U499 (N_499,In_61,In_262);
or U500 (N_500,In_48,In_234);
and U501 (N_501,In_408,In_27);
xor U502 (N_502,In_319,In_354);
nand U503 (N_503,In_456,In_171);
nand U504 (N_504,In_35,In_270);
nand U505 (N_505,In_396,In_413);
xor U506 (N_506,In_82,In_375);
nor U507 (N_507,In_95,In_459);
nor U508 (N_508,In_423,In_167);
nor U509 (N_509,In_17,In_221);
nor U510 (N_510,In_98,In_74);
and U511 (N_511,In_363,In_352);
or U512 (N_512,In_1,In_12);
or U513 (N_513,In_462,In_110);
and U514 (N_514,In_335,In_419);
nor U515 (N_515,In_274,In_204);
or U516 (N_516,In_82,In_11);
nor U517 (N_517,In_362,In_24);
nor U518 (N_518,In_213,In_446);
and U519 (N_519,In_479,In_310);
and U520 (N_520,In_65,In_112);
and U521 (N_521,In_359,In_80);
and U522 (N_522,In_357,In_37);
or U523 (N_523,In_195,In_14);
nor U524 (N_524,In_331,In_400);
nor U525 (N_525,In_460,In_455);
or U526 (N_526,In_228,In_439);
nor U527 (N_527,In_280,In_68);
or U528 (N_528,In_117,In_406);
or U529 (N_529,In_491,In_386);
nor U530 (N_530,In_157,In_371);
and U531 (N_531,In_317,In_11);
nor U532 (N_532,In_101,In_240);
and U533 (N_533,In_283,In_402);
xnor U534 (N_534,In_231,In_222);
xnor U535 (N_535,In_366,In_38);
nand U536 (N_536,In_469,In_228);
nand U537 (N_537,In_499,In_384);
xor U538 (N_538,In_24,In_249);
or U539 (N_539,In_139,In_65);
or U540 (N_540,In_192,In_319);
or U541 (N_541,In_304,In_9);
xor U542 (N_542,In_423,In_25);
nor U543 (N_543,In_444,In_147);
nor U544 (N_544,In_145,In_291);
nor U545 (N_545,In_370,In_195);
nand U546 (N_546,In_325,In_372);
or U547 (N_547,In_162,In_288);
nand U548 (N_548,In_172,In_202);
nor U549 (N_549,In_69,In_227);
nor U550 (N_550,In_355,In_296);
nor U551 (N_551,In_350,In_50);
nand U552 (N_552,In_203,In_331);
nand U553 (N_553,In_404,In_378);
and U554 (N_554,In_374,In_281);
and U555 (N_555,In_46,In_497);
nand U556 (N_556,In_19,In_60);
and U557 (N_557,In_219,In_345);
nor U558 (N_558,In_419,In_358);
and U559 (N_559,In_436,In_310);
and U560 (N_560,In_410,In_439);
and U561 (N_561,In_142,In_256);
xor U562 (N_562,In_52,In_134);
xnor U563 (N_563,In_199,In_476);
nor U564 (N_564,In_256,In_276);
nand U565 (N_565,In_158,In_3);
nor U566 (N_566,In_139,In_375);
nor U567 (N_567,In_227,In_238);
nand U568 (N_568,In_62,In_82);
and U569 (N_569,In_258,In_94);
nor U570 (N_570,In_337,In_353);
nand U571 (N_571,In_404,In_63);
and U572 (N_572,In_447,In_426);
and U573 (N_573,In_403,In_226);
and U574 (N_574,In_364,In_435);
nor U575 (N_575,In_365,In_71);
nor U576 (N_576,In_212,In_452);
nor U577 (N_577,In_252,In_272);
and U578 (N_578,In_266,In_4);
xnor U579 (N_579,In_395,In_100);
and U580 (N_580,In_226,In_195);
nand U581 (N_581,In_192,In_254);
or U582 (N_582,In_176,In_114);
or U583 (N_583,In_68,In_368);
nor U584 (N_584,In_126,In_6);
and U585 (N_585,In_231,In_332);
and U586 (N_586,In_226,In_259);
and U587 (N_587,In_251,In_219);
xor U588 (N_588,In_431,In_236);
xnor U589 (N_589,In_42,In_294);
nand U590 (N_590,In_288,In_431);
nand U591 (N_591,In_240,In_96);
and U592 (N_592,In_44,In_325);
or U593 (N_593,In_340,In_430);
nand U594 (N_594,In_184,In_370);
xor U595 (N_595,In_233,In_292);
nand U596 (N_596,In_457,In_325);
and U597 (N_597,In_265,In_259);
nor U598 (N_598,In_205,In_137);
or U599 (N_599,In_208,In_422);
nor U600 (N_600,N_151,N_114);
nand U601 (N_601,N_106,N_162);
nor U602 (N_602,N_298,N_459);
or U603 (N_603,N_243,N_235);
or U604 (N_604,N_398,N_122);
and U605 (N_605,N_217,N_263);
nor U606 (N_606,N_95,N_268);
nand U607 (N_607,N_517,N_148);
nand U608 (N_608,N_455,N_374);
nor U609 (N_609,N_325,N_200);
nor U610 (N_610,N_257,N_593);
nor U611 (N_611,N_242,N_313);
or U612 (N_612,N_103,N_135);
nor U613 (N_613,N_205,N_211);
and U614 (N_614,N_157,N_288);
or U615 (N_615,N_564,N_232);
or U616 (N_616,N_396,N_83);
nand U617 (N_617,N_289,N_482);
or U618 (N_618,N_477,N_33);
and U619 (N_619,N_516,N_264);
and U620 (N_620,N_328,N_9);
nand U621 (N_621,N_269,N_230);
nand U622 (N_622,N_185,N_565);
nor U623 (N_623,N_542,N_177);
xor U624 (N_624,N_154,N_433);
and U625 (N_625,N_493,N_387);
or U626 (N_626,N_373,N_457);
nand U627 (N_627,N_45,N_484);
or U628 (N_628,N_201,N_342);
nor U629 (N_629,N_81,N_173);
nand U630 (N_630,N_300,N_402);
nand U631 (N_631,N_52,N_98);
and U632 (N_632,N_391,N_485);
xor U633 (N_633,N_146,N_204);
nand U634 (N_634,N_527,N_577);
and U635 (N_635,N_216,N_592);
or U636 (N_636,N_164,N_237);
nand U637 (N_637,N_296,N_567);
nand U638 (N_638,N_41,N_510);
or U639 (N_639,N_348,N_572);
or U640 (N_640,N_29,N_432);
or U641 (N_641,N_584,N_134);
and U642 (N_642,N_74,N_30);
or U643 (N_643,N_421,N_440);
nand U644 (N_644,N_299,N_419);
nor U645 (N_645,N_522,N_405);
or U646 (N_646,N_339,N_65);
or U647 (N_647,N_520,N_557);
nor U648 (N_648,N_105,N_236);
nor U649 (N_649,N_426,N_350);
or U650 (N_650,N_110,N_182);
nor U651 (N_651,N_305,N_72);
nor U652 (N_652,N_153,N_219);
xor U653 (N_653,N_505,N_344);
nor U654 (N_654,N_561,N_128);
nand U655 (N_655,N_218,N_524);
nand U656 (N_656,N_434,N_131);
or U657 (N_657,N_360,N_14);
xor U658 (N_658,N_191,N_293);
nor U659 (N_659,N_221,N_258);
and U660 (N_660,N_531,N_539);
xnor U661 (N_661,N_479,N_279);
nor U662 (N_662,N_453,N_247);
xor U663 (N_663,N_447,N_1);
or U664 (N_664,N_306,N_111);
nor U665 (N_665,N_294,N_165);
nand U666 (N_666,N_196,N_591);
and U667 (N_667,N_48,N_290);
nor U668 (N_668,N_498,N_424);
nand U669 (N_669,N_580,N_598);
nand U670 (N_670,N_140,N_476);
nor U671 (N_671,N_275,N_280);
and U672 (N_672,N_368,N_112);
or U673 (N_673,N_208,N_176);
and U674 (N_674,N_12,N_530);
nor U675 (N_675,N_443,N_521);
or U676 (N_676,N_563,N_227);
nor U677 (N_677,N_251,N_502);
nand U678 (N_678,N_423,N_207);
and U679 (N_679,N_382,N_108);
and U680 (N_680,N_213,N_341);
or U681 (N_681,N_101,N_538);
nor U682 (N_682,N_533,N_2);
or U683 (N_683,N_158,N_399);
and U684 (N_684,N_214,N_241);
or U685 (N_685,N_333,N_470);
or U686 (N_686,N_511,N_137);
and U687 (N_687,N_49,N_354);
nand U688 (N_688,N_377,N_425);
nor U689 (N_689,N_535,N_195);
or U690 (N_690,N_392,N_460);
xnor U691 (N_691,N_389,N_24);
or U692 (N_692,N_576,N_599);
or U693 (N_693,N_570,N_64);
or U694 (N_694,N_141,N_249);
nor U695 (N_695,N_94,N_320);
nand U696 (N_696,N_19,N_166);
nor U697 (N_697,N_85,N_515);
and U698 (N_698,N_430,N_347);
and U699 (N_699,N_272,N_507);
nor U700 (N_700,N_285,N_70);
and U701 (N_701,N_465,N_406);
and U702 (N_702,N_458,N_509);
or U703 (N_703,N_337,N_283);
or U704 (N_704,N_566,N_228);
xnor U705 (N_705,N_132,N_192);
nor U706 (N_706,N_34,N_159);
and U707 (N_707,N_316,N_332);
or U708 (N_708,N_252,N_15);
or U709 (N_709,N_60,N_536);
and U710 (N_710,N_256,N_528);
and U711 (N_711,N_17,N_439);
and U712 (N_712,N_359,N_197);
nor U713 (N_713,N_203,N_513);
or U714 (N_714,N_560,N_278);
nor U715 (N_715,N_273,N_326);
nand U716 (N_716,N_54,N_68);
nor U717 (N_717,N_362,N_178);
and U718 (N_718,N_353,N_260);
or U719 (N_719,N_469,N_35);
nand U720 (N_720,N_427,N_78);
and U721 (N_721,N_22,N_156);
nor U722 (N_722,N_59,N_555);
xor U723 (N_723,N_590,N_315);
or U724 (N_724,N_335,N_152);
nor U725 (N_725,N_518,N_297);
nand U726 (N_726,N_578,N_548);
nand U727 (N_727,N_194,N_163);
nor U728 (N_728,N_383,N_361);
and U729 (N_729,N_544,N_464);
or U730 (N_730,N_394,N_384);
and U731 (N_731,N_117,N_345);
nand U732 (N_732,N_307,N_80);
or U733 (N_733,N_473,N_220);
nor U734 (N_734,N_231,N_11);
nor U735 (N_735,N_107,N_483);
xnor U736 (N_736,N_526,N_579);
nor U737 (N_737,N_545,N_596);
nor U738 (N_738,N_364,N_202);
and U739 (N_739,N_26,N_181);
nand U740 (N_740,N_376,N_388);
or U741 (N_741,N_16,N_130);
or U742 (N_742,N_451,N_149);
and U743 (N_743,N_93,N_274);
and U744 (N_744,N_73,N_317);
nor U745 (N_745,N_336,N_188);
or U746 (N_746,N_481,N_450);
and U747 (N_747,N_547,N_248);
and U748 (N_748,N_575,N_301);
nand U749 (N_749,N_120,N_343);
nor U750 (N_750,N_222,N_329);
nor U751 (N_751,N_187,N_304);
nor U752 (N_752,N_338,N_3);
or U753 (N_753,N_327,N_552);
or U754 (N_754,N_551,N_210);
and U755 (N_755,N_125,N_184);
xor U756 (N_756,N_136,N_346);
and U757 (N_757,N_116,N_77);
nand U758 (N_758,N_127,N_379);
nand U759 (N_759,N_109,N_415);
and U760 (N_760,N_523,N_238);
xnor U761 (N_761,N_67,N_287);
xor U762 (N_762,N_139,N_369);
or U763 (N_763,N_586,N_322);
and U764 (N_764,N_129,N_261);
nor U765 (N_765,N_411,N_244);
and U766 (N_766,N_161,N_47);
and U767 (N_767,N_553,N_413);
nor U768 (N_768,N_250,N_71);
nor U769 (N_769,N_6,N_365);
nand U770 (N_770,N_58,N_417);
nor U771 (N_771,N_574,N_319);
or U772 (N_772,N_10,N_492);
nand U773 (N_773,N_0,N_223);
nand U774 (N_774,N_89,N_349);
and U775 (N_775,N_282,N_234);
nor U776 (N_776,N_486,N_104);
xor U777 (N_777,N_529,N_437);
and U778 (N_778,N_587,N_597);
or U779 (N_779,N_50,N_167);
or U780 (N_780,N_562,N_489);
or U781 (N_781,N_314,N_96);
xor U782 (N_782,N_594,N_534);
nor U783 (N_783,N_255,N_265);
nand U784 (N_784,N_412,N_401);
nor U785 (N_785,N_118,N_262);
nand U786 (N_786,N_546,N_514);
nand U787 (N_787,N_142,N_418);
or U788 (N_788,N_206,N_56);
nor U789 (N_789,N_340,N_53);
or U790 (N_790,N_504,N_147);
and U791 (N_791,N_454,N_429);
nor U792 (N_792,N_400,N_324);
and U793 (N_793,N_267,N_284);
and U794 (N_794,N_276,N_386);
nand U795 (N_795,N_583,N_259);
xor U796 (N_796,N_186,N_441);
and U797 (N_797,N_121,N_155);
nand U798 (N_798,N_436,N_435);
and U799 (N_799,N_233,N_519);
nor U800 (N_800,N_445,N_23);
nor U801 (N_801,N_31,N_372);
xor U802 (N_802,N_295,N_496);
nand U803 (N_803,N_75,N_225);
xor U804 (N_804,N_254,N_308);
nand U805 (N_805,N_99,N_82);
xnor U806 (N_806,N_356,N_449);
and U807 (N_807,N_488,N_487);
nand U808 (N_808,N_174,N_366);
and U809 (N_809,N_568,N_160);
xnor U810 (N_810,N_506,N_588);
nand U811 (N_811,N_199,N_76);
nand U812 (N_812,N_46,N_8);
or U813 (N_813,N_277,N_390);
xnor U814 (N_814,N_585,N_172);
nand U815 (N_815,N_138,N_13);
nand U816 (N_816,N_7,N_474);
or U817 (N_817,N_318,N_170);
and U818 (N_818,N_475,N_471);
and U819 (N_819,N_97,N_495);
and U820 (N_820,N_480,N_28);
or U821 (N_821,N_503,N_51);
or U822 (N_822,N_303,N_358);
or U823 (N_823,N_79,N_370);
xnor U824 (N_824,N_271,N_478);
nor U825 (N_825,N_462,N_44);
or U826 (N_826,N_215,N_532);
nand U827 (N_827,N_330,N_168);
nand U828 (N_828,N_537,N_549);
nand U829 (N_829,N_589,N_119);
nand U830 (N_830,N_87,N_126);
nor U831 (N_831,N_43,N_407);
nand U832 (N_832,N_352,N_42);
or U833 (N_833,N_569,N_408);
or U834 (N_834,N_190,N_183);
nor U835 (N_835,N_57,N_169);
and U836 (N_836,N_92,N_66);
and U837 (N_837,N_312,N_84);
nand U838 (N_838,N_150,N_371);
and U839 (N_839,N_375,N_380);
nor U840 (N_840,N_212,N_448);
and U841 (N_841,N_102,N_438);
or U842 (N_842,N_461,N_355);
nor U843 (N_843,N_209,N_452);
or U844 (N_844,N_229,N_189);
xor U845 (N_845,N_309,N_403);
nand U846 (N_846,N_573,N_541);
or U847 (N_847,N_500,N_409);
nor U848 (N_848,N_18,N_144);
and U849 (N_849,N_311,N_497);
nor U850 (N_850,N_404,N_422);
and U851 (N_851,N_175,N_397);
and U852 (N_852,N_351,N_323);
nor U853 (N_853,N_385,N_357);
or U854 (N_854,N_395,N_554);
nor U855 (N_855,N_63,N_499);
and U856 (N_856,N_331,N_226);
or U857 (N_857,N_334,N_270);
nand U858 (N_858,N_456,N_39);
and U859 (N_859,N_310,N_302);
nand U860 (N_860,N_179,N_363);
or U861 (N_861,N_21,N_291);
nand U862 (N_862,N_25,N_467);
and U863 (N_863,N_145,N_556);
and U864 (N_864,N_428,N_253);
and U865 (N_865,N_180,N_468);
nand U866 (N_866,N_133,N_525);
and U867 (N_867,N_442,N_286);
nand U868 (N_868,N_466,N_198);
nand U869 (N_869,N_420,N_36);
or U870 (N_870,N_86,N_540);
nor U871 (N_871,N_27,N_37);
nand U872 (N_872,N_410,N_490);
nand U873 (N_873,N_113,N_472);
or U874 (N_874,N_32,N_62);
xor U875 (N_875,N_463,N_431);
and U876 (N_876,N_61,N_543);
nand U877 (N_877,N_266,N_91);
nor U878 (N_878,N_100,N_40);
nor U879 (N_879,N_444,N_582);
nand U880 (N_880,N_367,N_381);
and U881 (N_881,N_124,N_4);
and U882 (N_882,N_321,N_246);
and U883 (N_883,N_88,N_20);
nand U884 (N_884,N_494,N_512);
and U885 (N_885,N_5,N_115);
or U886 (N_886,N_55,N_171);
or U887 (N_887,N_571,N_123);
or U888 (N_888,N_90,N_581);
nand U889 (N_889,N_245,N_393);
or U890 (N_890,N_143,N_193);
or U891 (N_891,N_550,N_239);
xor U892 (N_892,N_416,N_491);
and U893 (N_893,N_446,N_559);
nand U894 (N_894,N_224,N_414);
nand U895 (N_895,N_558,N_378);
nand U896 (N_896,N_292,N_501);
and U897 (N_897,N_595,N_508);
nand U898 (N_898,N_281,N_38);
or U899 (N_899,N_240,N_69);
nand U900 (N_900,N_383,N_227);
and U901 (N_901,N_230,N_263);
nand U902 (N_902,N_15,N_55);
nand U903 (N_903,N_116,N_51);
nand U904 (N_904,N_270,N_178);
and U905 (N_905,N_368,N_569);
or U906 (N_906,N_576,N_60);
and U907 (N_907,N_253,N_520);
xnor U908 (N_908,N_146,N_513);
nand U909 (N_909,N_135,N_555);
nor U910 (N_910,N_464,N_493);
nand U911 (N_911,N_519,N_158);
nand U912 (N_912,N_405,N_534);
and U913 (N_913,N_80,N_593);
nor U914 (N_914,N_542,N_313);
nand U915 (N_915,N_287,N_260);
nor U916 (N_916,N_532,N_205);
and U917 (N_917,N_136,N_120);
nor U918 (N_918,N_382,N_376);
or U919 (N_919,N_101,N_574);
nand U920 (N_920,N_106,N_212);
and U921 (N_921,N_277,N_312);
and U922 (N_922,N_103,N_268);
and U923 (N_923,N_341,N_553);
nor U924 (N_924,N_216,N_384);
and U925 (N_925,N_23,N_124);
or U926 (N_926,N_326,N_426);
nor U927 (N_927,N_484,N_430);
xnor U928 (N_928,N_125,N_278);
nor U929 (N_929,N_352,N_573);
nor U930 (N_930,N_186,N_535);
and U931 (N_931,N_219,N_283);
nand U932 (N_932,N_300,N_379);
xnor U933 (N_933,N_551,N_381);
nor U934 (N_934,N_83,N_528);
nor U935 (N_935,N_378,N_176);
or U936 (N_936,N_71,N_468);
or U937 (N_937,N_455,N_464);
xnor U938 (N_938,N_286,N_91);
nand U939 (N_939,N_495,N_492);
or U940 (N_940,N_304,N_170);
or U941 (N_941,N_250,N_104);
or U942 (N_942,N_32,N_40);
and U943 (N_943,N_32,N_17);
and U944 (N_944,N_29,N_273);
and U945 (N_945,N_59,N_182);
nor U946 (N_946,N_111,N_37);
and U947 (N_947,N_525,N_500);
xor U948 (N_948,N_379,N_283);
nand U949 (N_949,N_260,N_17);
or U950 (N_950,N_413,N_308);
xnor U951 (N_951,N_193,N_73);
nand U952 (N_952,N_295,N_242);
nor U953 (N_953,N_13,N_126);
nor U954 (N_954,N_142,N_237);
or U955 (N_955,N_508,N_368);
and U956 (N_956,N_210,N_10);
nor U957 (N_957,N_204,N_45);
nor U958 (N_958,N_347,N_173);
xor U959 (N_959,N_523,N_166);
or U960 (N_960,N_419,N_51);
xnor U961 (N_961,N_349,N_305);
or U962 (N_962,N_494,N_161);
or U963 (N_963,N_257,N_173);
nor U964 (N_964,N_243,N_578);
nor U965 (N_965,N_91,N_122);
and U966 (N_966,N_133,N_562);
and U967 (N_967,N_114,N_476);
or U968 (N_968,N_274,N_468);
or U969 (N_969,N_175,N_52);
or U970 (N_970,N_492,N_568);
nand U971 (N_971,N_91,N_22);
or U972 (N_972,N_74,N_519);
or U973 (N_973,N_66,N_444);
and U974 (N_974,N_218,N_574);
and U975 (N_975,N_351,N_466);
nor U976 (N_976,N_195,N_527);
xor U977 (N_977,N_507,N_572);
xnor U978 (N_978,N_283,N_385);
nor U979 (N_979,N_263,N_380);
nand U980 (N_980,N_327,N_65);
nand U981 (N_981,N_327,N_505);
and U982 (N_982,N_567,N_505);
or U983 (N_983,N_49,N_524);
nand U984 (N_984,N_53,N_469);
nor U985 (N_985,N_329,N_479);
and U986 (N_986,N_302,N_546);
and U987 (N_987,N_597,N_321);
or U988 (N_988,N_498,N_99);
xnor U989 (N_989,N_466,N_480);
nand U990 (N_990,N_95,N_354);
or U991 (N_991,N_555,N_353);
and U992 (N_992,N_346,N_145);
or U993 (N_993,N_34,N_366);
and U994 (N_994,N_459,N_66);
and U995 (N_995,N_247,N_541);
nand U996 (N_996,N_566,N_378);
xnor U997 (N_997,N_329,N_233);
nor U998 (N_998,N_473,N_274);
nand U999 (N_999,N_174,N_415);
nand U1000 (N_1000,N_409,N_475);
and U1001 (N_1001,N_579,N_544);
and U1002 (N_1002,N_358,N_427);
nand U1003 (N_1003,N_527,N_413);
nor U1004 (N_1004,N_198,N_471);
nor U1005 (N_1005,N_424,N_410);
and U1006 (N_1006,N_430,N_181);
or U1007 (N_1007,N_580,N_303);
nor U1008 (N_1008,N_179,N_337);
nor U1009 (N_1009,N_277,N_335);
or U1010 (N_1010,N_472,N_178);
nand U1011 (N_1011,N_591,N_491);
nor U1012 (N_1012,N_545,N_252);
or U1013 (N_1013,N_319,N_488);
nand U1014 (N_1014,N_5,N_518);
or U1015 (N_1015,N_268,N_373);
xor U1016 (N_1016,N_367,N_189);
and U1017 (N_1017,N_149,N_503);
and U1018 (N_1018,N_110,N_502);
xor U1019 (N_1019,N_53,N_536);
nand U1020 (N_1020,N_122,N_28);
nand U1021 (N_1021,N_249,N_422);
nand U1022 (N_1022,N_542,N_400);
nor U1023 (N_1023,N_566,N_192);
and U1024 (N_1024,N_233,N_380);
and U1025 (N_1025,N_532,N_318);
or U1026 (N_1026,N_145,N_150);
and U1027 (N_1027,N_236,N_422);
xor U1028 (N_1028,N_305,N_403);
nor U1029 (N_1029,N_281,N_15);
or U1030 (N_1030,N_361,N_327);
or U1031 (N_1031,N_515,N_595);
nand U1032 (N_1032,N_201,N_46);
nand U1033 (N_1033,N_250,N_41);
nor U1034 (N_1034,N_214,N_146);
or U1035 (N_1035,N_319,N_228);
or U1036 (N_1036,N_291,N_23);
and U1037 (N_1037,N_586,N_223);
nor U1038 (N_1038,N_332,N_157);
nor U1039 (N_1039,N_247,N_543);
nand U1040 (N_1040,N_47,N_401);
nor U1041 (N_1041,N_543,N_331);
nand U1042 (N_1042,N_87,N_439);
and U1043 (N_1043,N_270,N_97);
or U1044 (N_1044,N_461,N_104);
nand U1045 (N_1045,N_161,N_170);
nor U1046 (N_1046,N_51,N_177);
and U1047 (N_1047,N_158,N_163);
and U1048 (N_1048,N_222,N_181);
xnor U1049 (N_1049,N_446,N_526);
or U1050 (N_1050,N_221,N_189);
nand U1051 (N_1051,N_55,N_96);
nor U1052 (N_1052,N_270,N_424);
or U1053 (N_1053,N_373,N_596);
or U1054 (N_1054,N_212,N_55);
and U1055 (N_1055,N_556,N_513);
and U1056 (N_1056,N_400,N_80);
nor U1057 (N_1057,N_40,N_69);
and U1058 (N_1058,N_339,N_237);
nor U1059 (N_1059,N_434,N_51);
or U1060 (N_1060,N_240,N_450);
nand U1061 (N_1061,N_465,N_281);
or U1062 (N_1062,N_258,N_129);
nand U1063 (N_1063,N_524,N_253);
nand U1064 (N_1064,N_458,N_155);
nand U1065 (N_1065,N_445,N_595);
or U1066 (N_1066,N_137,N_588);
or U1067 (N_1067,N_157,N_305);
or U1068 (N_1068,N_474,N_280);
nor U1069 (N_1069,N_197,N_98);
xor U1070 (N_1070,N_507,N_508);
or U1071 (N_1071,N_155,N_380);
nor U1072 (N_1072,N_64,N_593);
nand U1073 (N_1073,N_42,N_427);
or U1074 (N_1074,N_152,N_496);
and U1075 (N_1075,N_49,N_449);
or U1076 (N_1076,N_89,N_104);
nand U1077 (N_1077,N_316,N_596);
and U1078 (N_1078,N_197,N_150);
nor U1079 (N_1079,N_486,N_246);
nor U1080 (N_1080,N_423,N_275);
or U1081 (N_1081,N_33,N_18);
nand U1082 (N_1082,N_168,N_498);
or U1083 (N_1083,N_25,N_408);
and U1084 (N_1084,N_469,N_277);
nor U1085 (N_1085,N_546,N_99);
nor U1086 (N_1086,N_542,N_419);
nor U1087 (N_1087,N_62,N_522);
and U1088 (N_1088,N_266,N_416);
and U1089 (N_1089,N_13,N_228);
and U1090 (N_1090,N_246,N_420);
or U1091 (N_1091,N_343,N_366);
and U1092 (N_1092,N_446,N_81);
xnor U1093 (N_1093,N_109,N_71);
nand U1094 (N_1094,N_538,N_394);
or U1095 (N_1095,N_578,N_577);
xor U1096 (N_1096,N_466,N_380);
nand U1097 (N_1097,N_429,N_108);
or U1098 (N_1098,N_121,N_124);
and U1099 (N_1099,N_10,N_259);
nor U1100 (N_1100,N_37,N_238);
and U1101 (N_1101,N_539,N_21);
nor U1102 (N_1102,N_498,N_417);
nor U1103 (N_1103,N_539,N_204);
nor U1104 (N_1104,N_507,N_267);
nor U1105 (N_1105,N_66,N_230);
xnor U1106 (N_1106,N_490,N_223);
nand U1107 (N_1107,N_497,N_419);
xor U1108 (N_1108,N_220,N_423);
xnor U1109 (N_1109,N_185,N_544);
nor U1110 (N_1110,N_246,N_482);
and U1111 (N_1111,N_355,N_295);
or U1112 (N_1112,N_284,N_446);
and U1113 (N_1113,N_244,N_546);
nand U1114 (N_1114,N_84,N_280);
nor U1115 (N_1115,N_419,N_326);
nand U1116 (N_1116,N_407,N_251);
or U1117 (N_1117,N_589,N_167);
nand U1118 (N_1118,N_431,N_357);
nand U1119 (N_1119,N_97,N_67);
and U1120 (N_1120,N_495,N_153);
nor U1121 (N_1121,N_255,N_474);
nand U1122 (N_1122,N_403,N_535);
nor U1123 (N_1123,N_573,N_370);
and U1124 (N_1124,N_551,N_368);
and U1125 (N_1125,N_191,N_397);
nand U1126 (N_1126,N_346,N_447);
and U1127 (N_1127,N_10,N_414);
nor U1128 (N_1128,N_44,N_318);
nor U1129 (N_1129,N_302,N_461);
and U1130 (N_1130,N_416,N_43);
or U1131 (N_1131,N_412,N_107);
or U1132 (N_1132,N_101,N_265);
xnor U1133 (N_1133,N_226,N_18);
xor U1134 (N_1134,N_145,N_137);
and U1135 (N_1135,N_449,N_482);
nor U1136 (N_1136,N_486,N_474);
nand U1137 (N_1137,N_386,N_122);
nor U1138 (N_1138,N_519,N_599);
or U1139 (N_1139,N_71,N_34);
nor U1140 (N_1140,N_364,N_328);
or U1141 (N_1141,N_56,N_327);
nor U1142 (N_1142,N_302,N_466);
and U1143 (N_1143,N_191,N_380);
and U1144 (N_1144,N_19,N_40);
or U1145 (N_1145,N_418,N_185);
and U1146 (N_1146,N_269,N_313);
nor U1147 (N_1147,N_521,N_598);
or U1148 (N_1148,N_565,N_412);
or U1149 (N_1149,N_463,N_171);
and U1150 (N_1150,N_49,N_220);
and U1151 (N_1151,N_266,N_517);
nand U1152 (N_1152,N_345,N_562);
xor U1153 (N_1153,N_0,N_329);
xor U1154 (N_1154,N_248,N_44);
or U1155 (N_1155,N_220,N_357);
and U1156 (N_1156,N_322,N_346);
or U1157 (N_1157,N_490,N_101);
and U1158 (N_1158,N_100,N_250);
or U1159 (N_1159,N_460,N_581);
nand U1160 (N_1160,N_440,N_164);
nand U1161 (N_1161,N_286,N_387);
nand U1162 (N_1162,N_84,N_463);
or U1163 (N_1163,N_266,N_120);
or U1164 (N_1164,N_358,N_514);
or U1165 (N_1165,N_406,N_326);
and U1166 (N_1166,N_50,N_542);
nand U1167 (N_1167,N_97,N_368);
nand U1168 (N_1168,N_316,N_537);
and U1169 (N_1169,N_575,N_130);
and U1170 (N_1170,N_169,N_466);
or U1171 (N_1171,N_297,N_355);
xnor U1172 (N_1172,N_84,N_150);
nand U1173 (N_1173,N_286,N_476);
nor U1174 (N_1174,N_51,N_267);
and U1175 (N_1175,N_543,N_339);
and U1176 (N_1176,N_63,N_89);
nand U1177 (N_1177,N_150,N_298);
or U1178 (N_1178,N_150,N_310);
and U1179 (N_1179,N_8,N_545);
nor U1180 (N_1180,N_436,N_92);
nand U1181 (N_1181,N_478,N_197);
nor U1182 (N_1182,N_541,N_403);
nor U1183 (N_1183,N_516,N_160);
nor U1184 (N_1184,N_524,N_12);
nor U1185 (N_1185,N_356,N_112);
or U1186 (N_1186,N_286,N_253);
or U1187 (N_1187,N_474,N_319);
or U1188 (N_1188,N_579,N_35);
or U1189 (N_1189,N_222,N_308);
xor U1190 (N_1190,N_450,N_409);
and U1191 (N_1191,N_383,N_36);
and U1192 (N_1192,N_311,N_264);
nand U1193 (N_1193,N_247,N_473);
nand U1194 (N_1194,N_181,N_575);
or U1195 (N_1195,N_45,N_285);
or U1196 (N_1196,N_41,N_280);
nor U1197 (N_1197,N_133,N_541);
nor U1198 (N_1198,N_254,N_280);
nand U1199 (N_1199,N_56,N_168);
or U1200 (N_1200,N_1129,N_1151);
xnor U1201 (N_1201,N_1011,N_986);
nand U1202 (N_1202,N_613,N_841);
nand U1203 (N_1203,N_719,N_1157);
and U1204 (N_1204,N_1020,N_1114);
nand U1205 (N_1205,N_1058,N_786);
or U1206 (N_1206,N_631,N_1182);
and U1207 (N_1207,N_881,N_1130);
nor U1208 (N_1208,N_853,N_602);
and U1209 (N_1209,N_980,N_996);
and U1210 (N_1210,N_1110,N_1031);
or U1211 (N_1211,N_933,N_1173);
or U1212 (N_1212,N_718,N_643);
xnor U1213 (N_1213,N_805,N_738);
and U1214 (N_1214,N_971,N_1100);
or U1215 (N_1215,N_769,N_647);
and U1216 (N_1216,N_761,N_1174);
nor U1217 (N_1217,N_651,N_867);
or U1218 (N_1218,N_1112,N_1023);
or U1219 (N_1219,N_720,N_1098);
nor U1220 (N_1220,N_1022,N_886);
and U1221 (N_1221,N_840,N_808);
or U1222 (N_1222,N_1097,N_1106);
or U1223 (N_1223,N_1179,N_776);
and U1224 (N_1224,N_1070,N_1059);
and U1225 (N_1225,N_952,N_1089);
nand U1226 (N_1226,N_844,N_1145);
or U1227 (N_1227,N_610,N_794);
nor U1228 (N_1228,N_1030,N_764);
xnor U1229 (N_1229,N_1121,N_953);
nor U1230 (N_1230,N_984,N_681);
nand U1231 (N_1231,N_949,N_977);
or U1232 (N_1232,N_685,N_692);
xnor U1233 (N_1233,N_729,N_1139);
and U1234 (N_1234,N_1156,N_1144);
xor U1235 (N_1235,N_889,N_833);
nand U1236 (N_1236,N_1021,N_660);
or U1237 (N_1237,N_967,N_749);
or U1238 (N_1238,N_698,N_675);
or U1239 (N_1239,N_939,N_988);
nand U1240 (N_1240,N_696,N_1077);
nand U1241 (N_1241,N_1005,N_1009);
nor U1242 (N_1242,N_883,N_708);
nor U1243 (N_1243,N_1010,N_960);
or U1244 (N_1244,N_969,N_891);
or U1245 (N_1245,N_796,N_1135);
or U1246 (N_1246,N_918,N_1045);
and U1247 (N_1247,N_1085,N_614);
nor U1248 (N_1248,N_983,N_911);
or U1249 (N_1249,N_603,N_703);
and U1250 (N_1250,N_740,N_1159);
nand U1251 (N_1251,N_783,N_722);
and U1252 (N_1252,N_1087,N_807);
and U1253 (N_1253,N_734,N_1169);
and U1254 (N_1254,N_965,N_1187);
xnor U1255 (N_1255,N_1136,N_732);
nand U1256 (N_1256,N_816,N_1060);
nand U1257 (N_1257,N_970,N_682);
nor U1258 (N_1258,N_612,N_780);
or U1259 (N_1259,N_680,N_1111);
nand U1260 (N_1260,N_1091,N_1033);
nand U1261 (N_1261,N_1126,N_672);
or U1262 (N_1262,N_1189,N_802);
nand U1263 (N_1263,N_752,N_845);
or U1264 (N_1264,N_858,N_1071);
nor U1265 (N_1265,N_778,N_901);
nor U1266 (N_1266,N_1083,N_1047);
xnor U1267 (N_1267,N_1184,N_875);
or U1268 (N_1268,N_850,N_893);
and U1269 (N_1269,N_1119,N_1188);
or U1270 (N_1270,N_723,N_1143);
or U1271 (N_1271,N_750,N_691);
or U1272 (N_1272,N_644,N_617);
nor U1273 (N_1273,N_1049,N_630);
or U1274 (N_1274,N_982,N_627);
and U1275 (N_1275,N_846,N_639);
and U1276 (N_1276,N_1192,N_871);
xor U1277 (N_1277,N_1109,N_1040);
or U1278 (N_1278,N_999,N_632);
or U1279 (N_1279,N_1102,N_768);
and U1280 (N_1280,N_607,N_882);
or U1281 (N_1281,N_677,N_834);
nor U1282 (N_1282,N_1123,N_950);
nor U1283 (N_1283,N_1046,N_623);
nand U1284 (N_1284,N_878,N_756);
or U1285 (N_1285,N_709,N_766);
or U1286 (N_1286,N_605,N_945);
or U1287 (N_1287,N_1177,N_1050);
or U1288 (N_1288,N_1062,N_803);
nand U1289 (N_1289,N_1054,N_1073);
nand U1290 (N_1290,N_784,N_1028);
xnor U1291 (N_1291,N_827,N_633);
or U1292 (N_1292,N_801,N_777);
nand U1293 (N_1293,N_648,N_782);
and U1294 (N_1294,N_812,N_1007);
and U1295 (N_1295,N_962,N_940);
and U1296 (N_1296,N_820,N_1137);
and U1297 (N_1297,N_809,N_645);
and U1298 (N_1298,N_892,N_767);
nand U1299 (N_1299,N_929,N_819);
nor U1300 (N_1300,N_913,N_1080);
xor U1301 (N_1301,N_1079,N_731);
and U1302 (N_1302,N_890,N_1132);
xnor U1303 (N_1303,N_1168,N_813);
and U1304 (N_1304,N_877,N_1194);
or U1305 (N_1305,N_669,N_1148);
nand U1306 (N_1306,N_944,N_1064);
and U1307 (N_1307,N_955,N_1035);
and U1308 (N_1308,N_751,N_688);
or U1309 (N_1309,N_1092,N_1014);
nor U1310 (N_1310,N_1025,N_862);
nand U1311 (N_1311,N_626,N_637);
nand U1312 (N_1312,N_695,N_1118);
nor U1313 (N_1313,N_973,N_715);
or U1314 (N_1314,N_1082,N_914);
nand U1315 (N_1315,N_611,N_1038);
and U1316 (N_1316,N_941,N_868);
and U1317 (N_1317,N_924,N_628);
and U1318 (N_1318,N_759,N_1138);
or U1319 (N_1319,N_1176,N_652);
nor U1320 (N_1320,N_624,N_699);
or U1321 (N_1321,N_717,N_800);
and U1322 (N_1322,N_1147,N_727);
or U1323 (N_1323,N_873,N_900);
nor U1324 (N_1324,N_774,N_753);
and U1325 (N_1325,N_859,N_615);
nor U1326 (N_1326,N_1048,N_728);
and U1327 (N_1327,N_1003,N_1150);
nand U1328 (N_1328,N_638,N_765);
xor U1329 (N_1329,N_981,N_993);
xnor U1330 (N_1330,N_673,N_1072);
or U1331 (N_1331,N_898,N_1044);
and U1332 (N_1332,N_710,N_895);
xnor U1333 (N_1333,N_1037,N_1018);
and U1334 (N_1334,N_1076,N_619);
nand U1335 (N_1335,N_974,N_915);
xor U1336 (N_1336,N_1052,N_604);
nor U1337 (N_1337,N_1093,N_991);
nand U1338 (N_1338,N_625,N_842);
and U1339 (N_1339,N_757,N_706);
nand U1340 (N_1340,N_856,N_985);
nor U1341 (N_1341,N_847,N_702);
nor U1342 (N_1342,N_671,N_748);
nand U1343 (N_1343,N_676,N_1081);
or U1344 (N_1344,N_831,N_864);
and U1345 (N_1345,N_1034,N_811);
or U1346 (N_1346,N_855,N_919);
nor U1347 (N_1347,N_1131,N_649);
xor U1348 (N_1348,N_1190,N_742);
xnor U1349 (N_1349,N_655,N_1001);
nand U1350 (N_1350,N_1012,N_640);
nor U1351 (N_1351,N_1108,N_1133);
or U1352 (N_1352,N_658,N_926);
xor U1353 (N_1353,N_665,N_931);
nand U1354 (N_1354,N_679,N_656);
and U1355 (N_1355,N_1006,N_1004);
nand U1356 (N_1356,N_650,N_747);
xor U1357 (N_1357,N_785,N_951);
xnor U1358 (N_1358,N_843,N_832);
nor U1359 (N_1359,N_1122,N_927);
and U1360 (N_1360,N_733,N_791);
and U1361 (N_1361,N_606,N_908);
nand U1362 (N_1362,N_1146,N_1162);
xor U1363 (N_1363,N_998,N_775);
or U1364 (N_1364,N_1128,N_1027);
or U1365 (N_1365,N_662,N_959);
or U1366 (N_1366,N_642,N_818);
xnor U1367 (N_1367,N_888,N_787);
or U1368 (N_1368,N_1165,N_792);
nor U1369 (N_1369,N_1068,N_760);
nand U1370 (N_1370,N_629,N_957);
nand U1371 (N_1371,N_1199,N_724);
and U1372 (N_1372,N_1026,N_1008);
nand U1373 (N_1373,N_1096,N_608);
nand U1374 (N_1374,N_746,N_1164);
and U1375 (N_1375,N_664,N_961);
nand U1376 (N_1376,N_975,N_925);
and U1377 (N_1377,N_795,N_948);
nand U1378 (N_1378,N_1013,N_1183);
nand U1379 (N_1379,N_869,N_601);
or U1380 (N_1380,N_815,N_958);
nand U1381 (N_1381,N_989,N_1103);
and U1382 (N_1382,N_799,N_1029);
xnor U1383 (N_1383,N_726,N_872);
or U1384 (N_1384,N_1115,N_997);
and U1385 (N_1385,N_1041,N_880);
or U1386 (N_1386,N_1043,N_700);
nor U1387 (N_1387,N_1036,N_1061);
nor U1388 (N_1388,N_1066,N_1032);
or U1389 (N_1389,N_790,N_852);
and U1390 (N_1390,N_865,N_670);
and U1391 (N_1391,N_1154,N_826);
xor U1392 (N_1392,N_896,N_705);
nor U1393 (N_1393,N_741,N_1000);
nor U1394 (N_1394,N_635,N_641);
nand U1395 (N_1395,N_1180,N_636);
nor U1396 (N_1396,N_861,N_1153);
or U1397 (N_1397,N_909,N_894);
xor U1398 (N_1398,N_755,N_912);
nand U1399 (N_1399,N_674,N_866);
and U1400 (N_1400,N_904,N_1116);
or U1401 (N_1401,N_1024,N_838);
and U1402 (N_1402,N_793,N_810);
nor U1403 (N_1403,N_646,N_1160);
nand U1404 (N_1404,N_713,N_976);
nand U1405 (N_1405,N_657,N_972);
nand U1406 (N_1406,N_1069,N_716);
or U1407 (N_1407,N_707,N_762);
or U1408 (N_1408,N_1063,N_902);
xor U1409 (N_1409,N_1057,N_835);
nand U1410 (N_1410,N_622,N_744);
or U1411 (N_1411,N_863,N_1056);
nor U1412 (N_1412,N_1163,N_916);
nor U1413 (N_1413,N_876,N_689);
and U1414 (N_1414,N_1055,N_1053);
nand U1415 (N_1415,N_666,N_1172);
nor U1416 (N_1416,N_823,N_600);
or U1417 (N_1417,N_1042,N_1161);
and U1418 (N_1418,N_798,N_987);
and U1419 (N_1419,N_1084,N_770);
nor U1420 (N_1420,N_854,N_874);
nor U1421 (N_1421,N_1170,N_1075);
nand U1422 (N_1422,N_887,N_737);
nor U1423 (N_1423,N_1166,N_721);
and U1424 (N_1424,N_966,N_788);
or U1425 (N_1425,N_697,N_839);
and U1426 (N_1426,N_1140,N_947);
and U1427 (N_1427,N_824,N_936);
and U1428 (N_1428,N_1065,N_781);
nor U1429 (N_1429,N_797,N_735);
and U1430 (N_1430,N_621,N_828);
nand U1431 (N_1431,N_905,N_990);
or U1432 (N_1432,N_1178,N_897);
nand U1433 (N_1433,N_921,N_995);
nand U1434 (N_1434,N_903,N_694);
nand U1435 (N_1435,N_964,N_712);
xor U1436 (N_1436,N_686,N_693);
xnor U1437 (N_1437,N_857,N_884);
or U1438 (N_1438,N_1094,N_779);
xnor U1439 (N_1439,N_1155,N_968);
or U1440 (N_1440,N_725,N_938);
and U1441 (N_1441,N_1107,N_930);
nor U1442 (N_1442,N_634,N_879);
xor U1443 (N_1443,N_711,N_917);
xnor U1444 (N_1444,N_817,N_848);
and U1445 (N_1445,N_849,N_932);
and U1446 (N_1446,N_979,N_992);
nor U1447 (N_1447,N_653,N_899);
and U1448 (N_1448,N_773,N_1142);
nor U1449 (N_1449,N_1167,N_736);
nor U1450 (N_1450,N_1193,N_1195);
nand U1451 (N_1451,N_829,N_616);
nor U1452 (N_1452,N_1120,N_923);
nand U1453 (N_1453,N_825,N_870);
xnor U1454 (N_1454,N_851,N_609);
and U1455 (N_1455,N_1186,N_763);
nand U1456 (N_1456,N_1019,N_739);
or U1457 (N_1457,N_618,N_684);
and U1458 (N_1458,N_1152,N_822);
nand U1459 (N_1459,N_1197,N_1051);
and U1460 (N_1460,N_1141,N_1002);
nand U1461 (N_1461,N_928,N_804);
nor U1462 (N_1462,N_920,N_754);
nor U1463 (N_1463,N_814,N_663);
nand U1464 (N_1464,N_830,N_678);
and U1465 (N_1465,N_683,N_789);
nand U1466 (N_1466,N_1127,N_1088);
or U1467 (N_1467,N_1074,N_687);
and U1468 (N_1468,N_758,N_885);
nand U1469 (N_1469,N_1117,N_836);
nand U1470 (N_1470,N_743,N_1125);
nor U1471 (N_1471,N_1134,N_946);
or U1472 (N_1472,N_1090,N_690);
and U1473 (N_1473,N_1086,N_667);
nor U1474 (N_1474,N_837,N_907);
and U1475 (N_1475,N_745,N_860);
and U1476 (N_1476,N_1104,N_730);
nand U1477 (N_1477,N_1175,N_954);
xnor U1478 (N_1478,N_910,N_1171);
nor U1479 (N_1479,N_1017,N_934);
nor U1480 (N_1480,N_956,N_1113);
and U1481 (N_1481,N_1039,N_963);
and U1482 (N_1482,N_772,N_668);
or U1483 (N_1483,N_937,N_661);
xnor U1484 (N_1484,N_1124,N_922);
nand U1485 (N_1485,N_1101,N_943);
nand U1486 (N_1486,N_1185,N_1015);
nand U1487 (N_1487,N_821,N_1158);
nor U1488 (N_1488,N_1191,N_806);
xnor U1489 (N_1489,N_714,N_771);
nand U1490 (N_1490,N_654,N_620);
nand U1491 (N_1491,N_701,N_935);
nor U1492 (N_1492,N_1196,N_1181);
and U1493 (N_1493,N_704,N_906);
nor U1494 (N_1494,N_1105,N_942);
or U1495 (N_1495,N_659,N_1078);
and U1496 (N_1496,N_1016,N_1198);
and U1497 (N_1497,N_978,N_1095);
nor U1498 (N_1498,N_1149,N_1067);
nand U1499 (N_1499,N_1099,N_994);
and U1500 (N_1500,N_791,N_1008);
or U1501 (N_1501,N_1127,N_892);
nand U1502 (N_1502,N_794,N_940);
nand U1503 (N_1503,N_998,N_710);
and U1504 (N_1504,N_812,N_1167);
nand U1505 (N_1505,N_1049,N_1187);
or U1506 (N_1506,N_713,N_966);
or U1507 (N_1507,N_843,N_679);
or U1508 (N_1508,N_658,N_736);
xnor U1509 (N_1509,N_1067,N_884);
and U1510 (N_1510,N_1043,N_605);
and U1511 (N_1511,N_1107,N_1183);
nand U1512 (N_1512,N_999,N_869);
xor U1513 (N_1513,N_874,N_1004);
nand U1514 (N_1514,N_965,N_850);
or U1515 (N_1515,N_619,N_982);
or U1516 (N_1516,N_948,N_632);
and U1517 (N_1517,N_748,N_921);
or U1518 (N_1518,N_886,N_781);
nand U1519 (N_1519,N_830,N_877);
and U1520 (N_1520,N_1078,N_830);
xnor U1521 (N_1521,N_689,N_635);
xor U1522 (N_1522,N_1036,N_618);
nor U1523 (N_1523,N_764,N_907);
or U1524 (N_1524,N_717,N_1090);
or U1525 (N_1525,N_1184,N_1029);
nand U1526 (N_1526,N_1092,N_877);
or U1527 (N_1527,N_1099,N_658);
and U1528 (N_1528,N_907,N_676);
or U1529 (N_1529,N_894,N_968);
nand U1530 (N_1530,N_787,N_768);
nor U1531 (N_1531,N_1011,N_701);
nor U1532 (N_1532,N_1088,N_615);
and U1533 (N_1533,N_911,N_619);
or U1534 (N_1534,N_807,N_1000);
or U1535 (N_1535,N_658,N_681);
nor U1536 (N_1536,N_902,N_857);
nor U1537 (N_1537,N_757,N_1057);
and U1538 (N_1538,N_941,N_724);
and U1539 (N_1539,N_830,N_1127);
and U1540 (N_1540,N_1195,N_1098);
and U1541 (N_1541,N_605,N_713);
and U1542 (N_1542,N_843,N_1004);
xnor U1543 (N_1543,N_960,N_772);
and U1544 (N_1544,N_1143,N_1158);
and U1545 (N_1545,N_1069,N_651);
and U1546 (N_1546,N_693,N_890);
nor U1547 (N_1547,N_1077,N_643);
nor U1548 (N_1548,N_779,N_880);
or U1549 (N_1549,N_954,N_618);
nor U1550 (N_1550,N_1075,N_1155);
or U1551 (N_1551,N_1026,N_966);
nor U1552 (N_1552,N_953,N_740);
nor U1553 (N_1553,N_1088,N_812);
xor U1554 (N_1554,N_771,N_802);
nor U1555 (N_1555,N_630,N_743);
and U1556 (N_1556,N_1124,N_870);
or U1557 (N_1557,N_1071,N_961);
xnor U1558 (N_1558,N_1017,N_790);
nor U1559 (N_1559,N_1117,N_950);
xnor U1560 (N_1560,N_1151,N_1062);
and U1561 (N_1561,N_1015,N_899);
nand U1562 (N_1562,N_1112,N_839);
nor U1563 (N_1563,N_1146,N_976);
or U1564 (N_1564,N_661,N_894);
or U1565 (N_1565,N_1040,N_1191);
nor U1566 (N_1566,N_964,N_967);
nand U1567 (N_1567,N_1083,N_911);
xor U1568 (N_1568,N_831,N_1008);
nand U1569 (N_1569,N_727,N_1020);
nand U1570 (N_1570,N_799,N_712);
or U1571 (N_1571,N_1021,N_1109);
nor U1572 (N_1572,N_939,N_934);
xnor U1573 (N_1573,N_727,N_709);
nand U1574 (N_1574,N_1141,N_911);
nand U1575 (N_1575,N_895,N_947);
and U1576 (N_1576,N_682,N_858);
nand U1577 (N_1577,N_825,N_1033);
nor U1578 (N_1578,N_1115,N_1090);
and U1579 (N_1579,N_646,N_711);
and U1580 (N_1580,N_1184,N_819);
xor U1581 (N_1581,N_1119,N_626);
nand U1582 (N_1582,N_1072,N_806);
or U1583 (N_1583,N_773,N_1023);
nand U1584 (N_1584,N_770,N_675);
or U1585 (N_1585,N_1132,N_1026);
or U1586 (N_1586,N_1199,N_1022);
and U1587 (N_1587,N_619,N_1021);
nor U1588 (N_1588,N_707,N_970);
nand U1589 (N_1589,N_749,N_1030);
nand U1590 (N_1590,N_1147,N_929);
nand U1591 (N_1591,N_737,N_701);
and U1592 (N_1592,N_970,N_619);
or U1593 (N_1593,N_620,N_779);
or U1594 (N_1594,N_1123,N_905);
nor U1595 (N_1595,N_1047,N_683);
nor U1596 (N_1596,N_810,N_783);
and U1597 (N_1597,N_828,N_1069);
or U1598 (N_1598,N_722,N_962);
or U1599 (N_1599,N_954,N_926);
or U1600 (N_1600,N_1172,N_1190);
xor U1601 (N_1601,N_711,N_730);
nor U1602 (N_1602,N_1153,N_958);
and U1603 (N_1603,N_645,N_882);
nand U1604 (N_1604,N_655,N_1114);
nor U1605 (N_1605,N_1010,N_1014);
or U1606 (N_1606,N_711,N_733);
or U1607 (N_1607,N_855,N_1024);
or U1608 (N_1608,N_665,N_1193);
nand U1609 (N_1609,N_1041,N_601);
and U1610 (N_1610,N_643,N_722);
nor U1611 (N_1611,N_701,N_1175);
nor U1612 (N_1612,N_801,N_722);
nand U1613 (N_1613,N_1164,N_1075);
xor U1614 (N_1614,N_1116,N_1106);
nand U1615 (N_1615,N_786,N_931);
nor U1616 (N_1616,N_1121,N_657);
and U1617 (N_1617,N_714,N_992);
or U1618 (N_1618,N_1138,N_1047);
nor U1619 (N_1619,N_947,N_1133);
nand U1620 (N_1620,N_1031,N_1153);
and U1621 (N_1621,N_607,N_822);
nor U1622 (N_1622,N_815,N_709);
nand U1623 (N_1623,N_603,N_881);
xor U1624 (N_1624,N_1189,N_671);
nor U1625 (N_1625,N_871,N_781);
or U1626 (N_1626,N_699,N_828);
nor U1627 (N_1627,N_904,N_637);
nor U1628 (N_1628,N_1099,N_670);
nor U1629 (N_1629,N_796,N_896);
or U1630 (N_1630,N_880,N_675);
xnor U1631 (N_1631,N_643,N_864);
or U1632 (N_1632,N_1143,N_639);
or U1633 (N_1633,N_626,N_1189);
nand U1634 (N_1634,N_1001,N_1010);
or U1635 (N_1635,N_612,N_1199);
nand U1636 (N_1636,N_931,N_1082);
nor U1637 (N_1637,N_1059,N_902);
nand U1638 (N_1638,N_964,N_1152);
or U1639 (N_1639,N_740,N_1181);
nor U1640 (N_1640,N_913,N_734);
and U1641 (N_1641,N_633,N_1092);
and U1642 (N_1642,N_1162,N_1184);
and U1643 (N_1643,N_717,N_868);
nand U1644 (N_1644,N_776,N_719);
nand U1645 (N_1645,N_601,N_954);
nand U1646 (N_1646,N_873,N_644);
nor U1647 (N_1647,N_733,N_1108);
or U1648 (N_1648,N_1075,N_1147);
or U1649 (N_1649,N_667,N_911);
nand U1650 (N_1650,N_930,N_901);
and U1651 (N_1651,N_835,N_1181);
nor U1652 (N_1652,N_904,N_649);
and U1653 (N_1653,N_1183,N_953);
or U1654 (N_1654,N_1092,N_824);
nor U1655 (N_1655,N_869,N_792);
nand U1656 (N_1656,N_1095,N_734);
or U1657 (N_1657,N_908,N_706);
nand U1658 (N_1658,N_1078,N_1022);
and U1659 (N_1659,N_621,N_835);
or U1660 (N_1660,N_1139,N_1151);
xor U1661 (N_1661,N_1090,N_1076);
nand U1662 (N_1662,N_1182,N_1195);
nand U1663 (N_1663,N_767,N_949);
xor U1664 (N_1664,N_882,N_821);
and U1665 (N_1665,N_1025,N_1109);
and U1666 (N_1666,N_637,N_1135);
xor U1667 (N_1667,N_937,N_654);
xor U1668 (N_1668,N_1108,N_881);
nor U1669 (N_1669,N_1070,N_1028);
or U1670 (N_1670,N_984,N_955);
and U1671 (N_1671,N_909,N_1119);
xnor U1672 (N_1672,N_1097,N_936);
nand U1673 (N_1673,N_1163,N_1113);
or U1674 (N_1674,N_857,N_1099);
nand U1675 (N_1675,N_815,N_1002);
and U1676 (N_1676,N_1157,N_815);
and U1677 (N_1677,N_733,N_692);
xor U1678 (N_1678,N_1162,N_605);
xnor U1679 (N_1679,N_677,N_660);
nand U1680 (N_1680,N_792,N_864);
and U1681 (N_1681,N_904,N_901);
or U1682 (N_1682,N_1118,N_693);
or U1683 (N_1683,N_614,N_954);
or U1684 (N_1684,N_671,N_931);
and U1685 (N_1685,N_1082,N_682);
and U1686 (N_1686,N_668,N_797);
xor U1687 (N_1687,N_686,N_973);
xnor U1688 (N_1688,N_1020,N_603);
nor U1689 (N_1689,N_834,N_704);
and U1690 (N_1690,N_1133,N_767);
xor U1691 (N_1691,N_648,N_1134);
or U1692 (N_1692,N_1015,N_956);
or U1693 (N_1693,N_605,N_823);
nand U1694 (N_1694,N_1049,N_1065);
and U1695 (N_1695,N_1092,N_855);
and U1696 (N_1696,N_930,N_1164);
nor U1697 (N_1697,N_905,N_770);
nor U1698 (N_1698,N_1077,N_918);
and U1699 (N_1699,N_918,N_718);
nor U1700 (N_1700,N_816,N_778);
nand U1701 (N_1701,N_1118,N_838);
nand U1702 (N_1702,N_653,N_720);
xnor U1703 (N_1703,N_1095,N_731);
or U1704 (N_1704,N_721,N_730);
nand U1705 (N_1705,N_884,N_737);
nor U1706 (N_1706,N_740,N_639);
or U1707 (N_1707,N_859,N_630);
and U1708 (N_1708,N_1143,N_925);
or U1709 (N_1709,N_634,N_927);
nor U1710 (N_1710,N_963,N_769);
xor U1711 (N_1711,N_1081,N_637);
nor U1712 (N_1712,N_795,N_1089);
nand U1713 (N_1713,N_716,N_630);
and U1714 (N_1714,N_1163,N_714);
and U1715 (N_1715,N_700,N_739);
or U1716 (N_1716,N_718,N_789);
and U1717 (N_1717,N_639,N_980);
or U1718 (N_1718,N_1013,N_625);
nand U1719 (N_1719,N_799,N_1139);
or U1720 (N_1720,N_1051,N_716);
nand U1721 (N_1721,N_735,N_907);
xor U1722 (N_1722,N_976,N_1162);
nor U1723 (N_1723,N_955,N_977);
or U1724 (N_1724,N_980,N_921);
and U1725 (N_1725,N_906,N_773);
or U1726 (N_1726,N_726,N_690);
and U1727 (N_1727,N_1180,N_1083);
or U1728 (N_1728,N_608,N_868);
and U1729 (N_1729,N_1105,N_1030);
nor U1730 (N_1730,N_731,N_1071);
and U1731 (N_1731,N_1081,N_1182);
xnor U1732 (N_1732,N_1125,N_777);
xnor U1733 (N_1733,N_937,N_986);
and U1734 (N_1734,N_656,N_690);
nand U1735 (N_1735,N_741,N_1158);
and U1736 (N_1736,N_771,N_998);
nand U1737 (N_1737,N_1063,N_608);
nor U1738 (N_1738,N_692,N_705);
and U1739 (N_1739,N_719,N_936);
and U1740 (N_1740,N_653,N_1012);
or U1741 (N_1741,N_945,N_795);
nor U1742 (N_1742,N_754,N_768);
or U1743 (N_1743,N_858,N_704);
xor U1744 (N_1744,N_989,N_896);
nor U1745 (N_1745,N_720,N_854);
nand U1746 (N_1746,N_1007,N_807);
nor U1747 (N_1747,N_1042,N_798);
or U1748 (N_1748,N_855,N_902);
and U1749 (N_1749,N_741,N_970);
nor U1750 (N_1750,N_651,N_816);
nor U1751 (N_1751,N_966,N_1020);
or U1752 (N_1752,N_1009,N_1099);
or U1753 (N_1753,N_827,N_935);
nor U1754 (N_1754,N_1141,N_841);
nand U1755 (N_1755,N_637,N_608);
or U1756 (N_1756,N_1119,N_930);
or U1757 (N_1757,N_650,N_1154);
xor U1758 (N_1758,N_958,N_651);
or U1759 (N_1759,N_738,N_830);
nor U1760 (N_1760,N_1181,N_1175);
or U1761 (N_1761,N_730,N_906);
or U1762 (N_1762,N_949,N_1063);
nor U1763 (N_1763,N_678,N_831);
or U1764 (N_1764,N_1172,N_675);
and U1765 (N_1765,N_850,N_742);
nor U1766 (N_1766,N_691,N_673);
or U1767 (N_1767,N_823,N_1179);
and U1768 (N_1768,N_936,N_841);
and U1769 (N_1769,N_1061,N_1129);
nor U1770 (N_1770,N_939,N_682);
and U1771 (N_1771,N_700,N_924);
nand U1772 (N_1772,N_914,N_1153);
nand U1773 (N_1773,N_877,N_644);
and U1774 (N_1774,N_1099,N_981);
or U1775 (N_1775,N_1034,N_654);
xor U1776 (N_1776,N_757,N_809);
nor U1777 (N_1777,N_984,N_1038);
and U1778 (N_1778,N_743,N_948);
and U1779 (N_1779,N_1162,N_690);
nor U1780 (N_1780,N_968,N_1189);
and U1781 (N_1781,N_1187,N_1029);
nand U1782 (N_1782,N_883,N_746);
nor U1783 (N_1783,N_609,N_762);
nand U1784 (N_1784,N_1072,N_982);
nor U1785 (N_1785,N_672,N_868);
nor U1786 (N_1786,N_935,N_784);
or U1787 (N_1787,N_1120,N_749);
or U1788 (N_1788,N_604,N_946);
and U1789 (N_1789,N_676,N_944);
nand U1790 (N_1790,N_1054,N_898);
nand U1791 (N_1791,N_1142,N_715);
and U1792 (N_1792,N_904,N_600);
or U1793 (N_1793,N_734,N_707);
and U1794 (N_1794,N_980,N_969);
nand U1795 (N_1795,N_728,N_1136);
and U1796 (N_1796,N_630,N_604);
nand U1797 (N_1797,N_1138,N_1148);
and U1798 (N_1798,N_892,N_810);
or U1799 (N_1799,N_783,N_1141);
and U1800 (N_1800,N_1344,N_1652);
or U1801 (N_1801,N_1567,N_1633);
and U1802 (N_1802,N_1675,N_1636);
xor U1803 (N_1803,N_1651,N_1484);
nand U1804 (N_1804,N_1530,N_1708);
and U1805 (N_1805,N_1786,N_1538);
and U1806 (N_1806,N_1333,N_1524);
and U1807 (N_1807,N_1368,N_1635);
and U1808 (N_1808,N_1458,N_1730);
nand U1809 (N_1809,N_1658,N_1372);
nor U1810 (N_1810,N_1650,N_1439);
or U1811 (N_1811,N_1315,N_1792);
nand U1812 (N_1812,N_1715,N_1479);
or U1813 (N_1813,N_1420,N_1232);
nor U1814 (N_1814,N_1396,N_1326);
nand U1815 (N_1815,N_1417,N_1663);
and U1816 (N_1816,N_1343,N_1548);
or U1817 (N_1817,N_1696,N_1661);
and U1818 (N_1818,N_1625,N_1339);
or U1819 (N_1819,N_1248,N_1491);
and U1820 (N_1820,N_1265,N_1593);
nand U1821 (N_1821,N_1296,N_1698);
nor U1822 (N_1822,N_1258,N_1649);
or U1823 (N_1823,N_1209,N_1744);
nand U1824 (N_1824,N_1240,N_1674);
and U1825 (N_1825,N_1781,N_1342);
or U1826 (N_1826,N_1543,N_1203);
and U1827 (N_1827,N_1383,N_1345);
nor U1828 (N_1828,N_1415,N_1582);
xnor U1829 (N_1829,N_1462,N_1602);
nand U1830 (N_1830,N_1388,N_1551);
or U1831 (N_1831,N_1359,N_1676);
nand U1832 (N_1832,N_1532,N_1742);
nor U1833 (N_1833,N_1774,N_1419);
nand U1834 (N_1834,N_1711,N_1644);
and U1835 (N_1835,N_1773,N_1719);
xor U1836 (N_1836,N_1374,N_1743);
or U1837 (N_1837,N_1778,N_1793);
nor U1838 (N_1838,N_1717,N_1303);
nand U1839 (N_1839,N_1401,N_1499);
nor U1840 (N_1840,N_1686,N_1590);
nor U1841 (N_1841,N_1723,N_1520);
xor U1842 (N_1842,N_1346,N_1560);
nand U1843 (N_1843,N_1596,N_1377);
and U1844 (N_1844,N_1550,N_1795);
nand U1845 (N_1845,N_1615,N_1647);
nand U1846 (N_1846,N_1208,N_1277);
xnor U1847 (N_1847,N_1279,N_1679);
or U1848 (N_1848,N_1256,N_1755);
and U1849 (N_1849,N_1317,N_1463);
nor U1850 (N_1850,N_1225,N_1340);
or U1851 (N_1851,N_1496,N_1216);
nor U1852 (N_1852,N_1525,N_1271);
or U1853 (N_1853,N_1607,N_1581);
and U1854 (N_1854,N_1580,N_1294);
nor U1855 (N_1855,N_1475,N_1626);
nor U1856 (N_1856,N_1378,N_1290);
and U1857 (N_1857,N_1362,N_1796);
or U1858 (N_1858,N_1302,N_1666);
nor U1859 (N_1859,N_1270,N_1735);
nor U1860 (N_1860,N_1628,N_1734);
xnor U1861 (N_1861,N_1230,N_1571);
nor U1862 (N_1862,N_1461,N_1214);
or U1863 (N_1863,N_1695,N_1613);
xnor U1864 (N_1864,N_1512,N_1598);
nor U1865 (N_1865,N_1211,N_1490);
nand U1866 (N_1866,N_1467,N_1752);
nor U1867 (N_1867,N_1609,N_1349);
nand U1868 (N_1868,N_1448,N_1684);
nor U1869 (N_1869,N_1367,N_1753);
nor U1870 (N_1870,N_1737,N_1478);
nor U1871 (N_1871,N_1263,N_1437);
or U1872 (N_1872,N_1562,N_1575);
and U1873 (N_1873,N_1757,N_1706);
or U1874 (N_1874,N_1207,N_1329);
and U1875 (N_1875,N_1432,N_1382);
nor U1876 (N_1876,N_1487,N_1255);
nand U1877 (N_1877,N_1336,N_1619);
nor U1878 (N_1878,N_1281,N_1239);
nand U1879 (N_1879,N_1614,N_1794);
nand U1880 (N_1880,N_1561,N_1295);
xnor U1881 (N_1881,N_1447,N_1264);
nor U1882 (N_1882,N_1418,N_1699);
nor U1883 (N_1883,N_1276,N_1384);
nand U1884 (N_1884,N_1784,N_1435);
nand U1885 (N_1885,N_1732,N_1429);
xor U1886 (N_1886,N_1622,N_1300);
nor U1887 (N_1887,N_1768,N_1506);
or U1888 (N_1888,N_1334,N_1728);
nor U1889 (N_1889,N_1783,N_1411);
or U1890 (N_1890,N_1714,N_1772);
and U1891 (N_1891,N_1597,N_1299);
nand U1892 (N_1892,N_1514,N_1246);
or U1893 (N_1893,N_1451,N_1671);
nor U1894 (N_1894,N_1552,N_1251);
and U1895 (N_1895,N_1243,N_1495);
nand U1896 (N_1896,N_1456,N_1351);
or U1897 (N_1897,N_1599,N_1505);
or U1898 (N_1898,N_1481,N_1528);
nand U1899 (N_1899,N_1617,N_1703);
nor U1900 (N_1900,N_1309,N_1438);
and U1901 (N_1901,N_1564,N_1779);
or U1902 (N_1902,N_1399,N_1412);
nand U1903 (N_1903,N_1523,N_1535);
or U1904 (N_1904,N_1387,N_1219);
nor U1905 (N_1905,N_1709,N_1400);
nand U1906 (N_1906,N_1369,N_1526);
and U1907 (N_1907,N_1254,N_1366);
xor U1908 (N_1908,N_1665,N_1540);
nand U1909 (N_1909,N_1226,N_1641);
nand U1910 (N_1910,N_1568,N_1591);
nor U1911 (N_1911,N_1325,N_1252);
nor U1912 (N_1912,N_1788,N_1515);
xnor U1913 (N_1913,N_1569,N_1237);
or U1914 (N_1914,N_1238,N_1537);
and U1915 (N_1915,N_1414,N_1332);
nand U1916 (N_1916,N_1354,N_1430);
nor U1917 (N_1917,N_1606,N_1397);
nor U1918 (N_1918,N_1427,N_1498);
or U1919 (N_1919,N_1555,N_1511);
nor U1920 (N_1920,N_1316,N_1223);
and U1921 (N_1921,N_1749,N_1260);
or U1922 (N_1922,N_1282,N_1765);
nand U1923 (N_1923,N_1693,N_1747);
nand U1924 (N_1924,N_1492,N_1426);
and U1925 (N_1925,N_1690,N_1454);
nand U1926 (N_1926,N_1659,N_1452);
and U1927 (N_1927,N_1241,N_1639);
nor U1928 (N_1928,N_1646,N_1390);
nor U1929 (N_1929,N_1436,N_1470);
nor U1930 (N_1930,N_1578,N_1485);
xnor U1931 (N_1931,N_1403,N_1740);
nand U1932 (N_1932,N_1306,N_1688);
and U1933 (N_1933,N_1691,N_1465);
or U1934 (N_1934,N_1477,N_1245);
nand U1935 (N_1935,N_1363,N_1664);
and U1936 (N_1936,N_1267,N_1750);
xor U1937 (N_1937,N_1413,N_1404);
or U1938 (N_1938,N_1656,N_1364);
or U1939 (N_1939,N_1601,N_1761);
nand U1940 (N_1940,N_1236,N_1573);
and U1941 (N_1941,N_1228,N_1433);
nand U1942 (N_1942,N_1331,N_1247);
nand U1943 (N_1943,N_1657,N_1507);
nand U1944 (N_1944,N_1450,N_1341);
nor U1945 (N_1945,N_1431,N_1324);
nor U1946 (N_1946,N_1545,N_1457);
and U1947 (N_1947,N_1678,N_1231);
or U1948 (N_1948,N_1780,N_1321);
nor U1949 (N_1949,N_1565,N_1623);
or U1950 (N_1950,N_1503,N_1553);
nor U1951 (N_1951,N_1529,N_1518);
or U1952 (N_1952,N_1718,N_1350);
or U1953 (N_1953,N_1308,N_1705);
xor U1954 (N_1954,N_1358,N_1204);
nand U1955 (N_1955,N_1253,N_1672);
nand U1956 (N_1956,N_1497,N_1767);
nand U1957 (N_1957,N_1513,N_1392);
or U1958 (N_1958,N_1476,N_1455);
nand U1959 (N_1959,N_1365,N_1287);
and U1960 (N_1960,N_1785,N_1704);
xnor U1961 (N_1961,N_1517,N_1293);
nor U1962 (N_1962,N_1616,N_1588);
nor U1963 (N_1963,N_1787,N_1782);
nand U1964 (N_1964,N_1681,N_1791);
or U1965 (N_1965,N_1662,N_1729);
nor U1966 (N_1966,N_1673,N_1554);
xor U1967 (N_1967,N_1637,N_1508);
and U1968 (N_1968,N_1670,N_1353);
nand U1969 (N_1969,N_1655,N_1471);
or U1970 (N_1970,N_1756,N_1269);
or U1971 (N_1971,N_1422,N_1604);
xor U1972 (N_1972,N_1483,N_1280);
and U1973 (N_1973,N_1371,N_1776);
or U1974 (N_1974,N_1583,N_1612);
nor U1975 (N_1975,N_1579,N_1224);
and U1976 (N_1976,N_1539,N_1777);
nand U1977 (N_1977,N_1234,N_1534);
or U1978 (N_1978,N_1307,N_1489);
nand U1979 (N_1979,N_1373,N_1504);
or U1980 (N_1980,N_1473,N_1592);
nand U1981 (N_1981,N_1653,N_1298);
xor U1982 (N_1982,N_1421,N_1542);
and U1983 (N_1983,N_1394,N_1682);
nand U1984 (N_1984,N_1493,N_1213);
nor U1985 (N_1985,N_1547,N_1640);
xnor U1986 (N_1986,N_1683,N_1510);
or U1987 (N_1987,N_1305,N_1328);
nand U1988 (N_1988,N_1301,N_1707);
or U1989 (N_1989,N_1629,N_1393);
nor U1990 (N_1990,N_1449,N_1304);
and U1991 (N_1991,N_1770,N_1235);
nor U1992 (N_1992,N_1720,N_1611);
or U1993 (N_1993,N_1405,N_1731);
nand U1994 (N_1994,N_1559,N_1408);
or U1995 (N_1995,N_1288,N_1566);
and U1996 (N_1996,N_1721,N_1763);
nor U1997 (N_1997,N_1710,N_1500);
and U1998 (N_1998,N_1310,N_1775);
and U1999 (N_1999,N_1425,N_1466);
nand U2000 (N_2000,N_1533,N_1380);
nor U2001 (N_2001,N_1585,N_1220);
or U2002 (N_2002,N_1416,N_1689);
or U2003 (N_2003,N_1259,N_1677);
and U2004 (N_2004,N_1445,N_1262);
nand U2005 (N_2005,N_1712,N_1621);
nand U2006 (N_2006,N_1292,N_1480);
nor U2007 (N_2007,N_1268,N_1557);
nand U2008 (N_2008,N_1217,N_1318);
xor U2009 (N_2009,N_1212,N_1798);
nand U2010 (N_2010,N_1522,N_1297);
nand U2011 (N_2011,N_1702,N_1386);
nor U2012 (N_2012,N_1531,N_1521);
nor U2013 (N_2013,N_1771,N_1726);
nand U2014 (N_2014,N_1697,N_1229);
or U2015 (N_2015,N_1274,N_1584);
nor U2016 (N_2016,N_1409,N_1746);
and U2017 (N_2017,N_1634,N_1642);
nor U2018 (N_2018,N_1284,N_1440);
or U2019 (N_2019,N_1638,N_1685);
nor U2020 (N_2020,N_1700,N_1724);
or U2021 (N_2021,N_1605,N_1618);
or U2022 (N_2022,N_1407,N_1441);
and U2023 (N_2023,N_1218,N_1244);
nand U2024 (N_2024,N_1736,N_1687);
xor U2025 (N_2025,N_1563,N_1327);
nor U2026 (N_2026,N_1630,N_1586);
and U2027 (N_2027,N_1589,N_1221);
nand U2028 (N_2028,N_1311,N_1745);
nor U2029 (N_2029,N_1716,N_1337);
or U2030 (N_2030,N_1398,N_1319);
or U2031 (N_2031,N_1249,N_1527);
nor U2032 (N_2032,N_1357,N_1556);
nor U2033 (N_2033,N_1453,N_1754);
xor U2034 (N_2034,N_1261,N_1648);
nand U2035 (N_2035,N_1289,N_1395);
nand U2036 (N_2036,N_1572,N_1667);
nand U2037 (N_2037,N_1516,N_1587);
and U2038 (N_2038,N_1222,N_1206);
nand U2039 (N_2039,N_1541,N_1227);
or U2040 (N_2040,N_1335,N_1286);
and U2041 (N_2041,N_1257,N_1424);
or U2042 (N_2042,N_1410,N_1608);
and U2043 (N_2043,N_1722,N_1469);
xor U2044 (N_2044,N_1789,N_1460);
or U2045 (N_2045,N_1370,N_1645);
nand U2046 (N_2046,N_1660,N_1624);
nand U2047 (N_2047,N_1355,N_1741);
or U2048 (N_2048,N_1570,N_1643);
nor U2049 (N_2049,N_1330,N_1549);
nor U2050 (N_2050,N_1283,N_1313);
and U2051 (N_2051,N_1797,N_1320);
nor U2052 (N_2052,N_1733,N_1338);
or U2053 (N_2053,N_1273,N_1620);
nand U2054 (N_2054,N_1764,N_1694);
or U2055 (N_2055,N_1356,N_1278);
xnor U2056 (N_2056,N_1758,N_1576);
or U2057 (N_2057,N_1352,N_1502);
and U2058 (N_2058,N_1443,N_1361);
nor U2059 (N_2059,N_1202,N_1762);
and U2060 (N_2060,N_1200,N_1360);
and U2061 (N_2061,N_1347,N_1323);
and U2062 (N_2062,N_1205,N_1442);
or U2063 (N_2063,N_1428,N_1468);
nand U2064 (N_2064,N_1434,N_1546);
and U2065 (N_2065,N_1536,N_1266);
xor U2066 (N_2066,N_1769,N_1668);
and U2067 (N_2067,N_1486,N_1391);
or U2068 (N_2068,N_1760,N_1375);
or U2069 (N_2069,N_1314,N_1488);
xnor U2070 (N_2070,N_1631,N_1603);
or U2071 (N_2071,N_1713,N_1739);
and U2072 (N_2072,N_1242,N_1444);
or U2073 (N_2073,N_1632,N_1381);
or U2074 (N_2074,N_1669,N_1385);
nor U2075 (N_2075,N_1285,N_1759);
or U2076 (N_2076,N_1348,N_1680);
and U2077 (N_2077,N_1692,N_1406);
or U2078 (N_2078,N_1766,N_1446);
xnor U2079 (N_2079,N_1610,N_1389);
or U2080 (N_2080,N_1701,N_1727);
nand U2081 (N_2081,N_1574,N_1312);
nand U2082 (N_2082,N_1799,N_1402);
and U2083 (N_2083,N_1544,N_1233);
nor U2084 (N_2084,N_1250,N_1751);
or U2085 (N_2085,N_1494,N_1210);
nand U2086 (N_2086,N_1654,N_1595);
and U2087 (N_2087,N_1215,N_1577);
nor U2088 (N_2088,N_1738,N_1790);
nand U2089 (N_2089,N_1459,N_1275);
xor U2090 (N_2090,N_1201,N_1472);
nand U2091 (N_2091,N_1725,N_1474);
and U2092 (N_2092,N_1509,N_1627);
and U2093 (N_2093,N_1322,N_1482);
or U2094 (N_2094,N_1501,N_1748);
or U2095 (N_2095,N_1379,N_1519);
or U2096 (N_2096,N_1423,N_1558);
and U2097 (N_2097,N_1291,N_1600);
and U2098 (N_2098,N_1376,N_1594);
nand U2099 (N_2099,N_1464,N_1272);
nor U2100 (N_2100,N_1392,N_1584);
nor U2101 (N_2101,N_1540,N_1300);
nor U2102 (N_2102,N_1220,N_1344);
nor U2103 (N_2103,N_1424,N_1742);
or U2104 (N_2104,N_1419,N_1400);
nand U2105 (N_2105,N_1696,N_1329);
nand U2106 (N_2106,N_1638,N_1750);
nor U2107 (N_2107,N_1466,N_1730);
and U2108 (N_2108,N_1413,N_1716);
or U2109 (N_2109,N_1211,N_1501);
nand U2110 (N_2110,N_1518,N_1536);
nor U2111 (N_2111,N_1490,N_1336);
or U2112 (N_2112,N_1766,N_1252);
or U2113 (N_2113,N_1643,N_1595);
and U2114 (N_2114,N_1242,N_1520);
or U2115 (N_2115,N_1414,N_1520);
nor U2116 (N_2116,N_1363,N_1542);
or U2117 (N_2117,N_1445,N_1649);
nand U2118 (N_2118,N_1232,N_1500);
and U2119 (N_2119,N_1658,N_1524);
nand U2120 (N_2120,N_1257,N_1403);
nor U2121 (N_2121,N_1312,N_1706);
or U2122 (N_2122,N_1338,N_1656);
nor U2123 (N_2123,N_1549,N_1687);
nor U2124 (N_2124,N_1204,N_1752);
and U2125 (N_2125,N_1244,N_1670);
nand U2126 (N_2126,N_1728,N_1515);
or U2127 (N_2127,N_1272,N_1604);
or U2128 (N_2128,N_1636,N_1611);
nand U2129 (N_2129,N_1407,N_1360);
xnor U2130 (N_2130,N_1658,N_1311);
nor U2131 (N_2131,N_1659,N_1493);
and U2132 (N_2132,N_1644,N_1393);
xor U2133 (N_2133,N_1215,N_1570);
and U2134 (N_2134,N_1742,N_1766);
nor U2135 (N_2135,N_1596,N_1710);
and U2136 (N_2136,N_1666,N_1428);
nand U2137 (N_2137,N_1491,N_1744);
or U2138 (N_2138,N_1544,N_1258);
or U2139 (N_2139,N_1647,N_1219);
nand U2140 (N_2140,N_1620,N_1309);
nand U2141 (N_2141,N_1285,N_1760);
nor U2142 (N_2142,N_1566,N_1791);
nand U2143 (N_2143,N_1262,N_1411);
nand U2144 (N_2144,N_1453,N_1796);
or U2145 (N_2145,N_1383,N_1609);
nor U2146 (N_2146,N_1448,N_1248);
nand U2147 (N_2147,N_1254,N_1495);
nand U2148 (N_2148,N_1637,N_1264);
xor U2149 (N_2149,N_1621,N_1383);
or U2150 (N_2150,N_1736,N_1599);
nand U2151 (N_2151,N_1337,N_1433);
or U2152 (N_2152,N_1790,N_1443);
nand U2153 (N_2153,N_1219,N_1371);
and U2154 (N_2154,N_1666,N_1782);
xnor U2155 (N_2155,N_1385,N_1630);
nor U2156 (N_2156,N_1535,N_1348);
or U2157 (N_2157,N_1293,N_1429);
or U2158 (N_2158,N_1288,N_1603);
nor U2159 (N_2159,N_1255,N_1784);
nor U2160 (N_2160,N_1345,N_1514);
and U2161 (N_2161,N_1510,N_1549);
xnor U2162 (N_2162,N_1717,N_1759);
xor U2163 (N_2163,N_1638,N_1445);
xnor U2164 (N_2164,N_1443,N_1235);
nor U2165 (N_2165,N_1263,N_1322);
nand U2166 (N_2166,N_1650,N_1699);
nor U2167 (N_2167,N_1771,N_1743);
xnor U2168 (N_2168,N_1517,N_1505);
or U2169 (N_2169,N_1214,N_1749);
xnor U2170 (N_2170,N_1438,N_1421);
xnor U2171 (N_2171,N_1658,N_1704);
nor U2172 (N_2172,N_1351,N_1309);
xnor U2173 (N_2173,N_1578,N_1603);
and U2174 (N_2174,N_1344,N_1704);
xor U2175 (N_2175,N_1308,N_1620);
xnor U2176 (N_2176,N_1703,N_1489);
nor U2177 (N_2177,N_1603,N_1760);
nor U2178 (N_2178,N_1789,N_1681);
nand U2179 (N_2179,N_1644,N_1654);
or U2180 (N_2180,N_1496,N_1702);
nand U2181 (N_2181,N_1356,N_1778);
nand U2182 (N_2182,N_1778,N_1332);
or U2183 (N_2183,N_1381,N_1747);
nor U2184 (N_2184,N_1442,N_1351);
nand U2185 (N_2185,N_1629,N_1703);
or U2186 (N_2186,N_1244,N_1601);
xor U2187 (N_2187,N_1639,N_1632);
nand U2188 (N_2188,N_1471,N_1794);
and U2189 (N_2189,N_1671,N_1655);
nor U2190 (N_2190,N_1511,N_1391);
or U2191 (N_2191,N_1411,N_1672);
nand U2192 (N_2192,N_1748,N_1600);
and U2193 (N_2193,N_1755,N_1746);
nand U2194 (N_2194,N_1744,N_1691);
nor U2195 (N_2195,N_1760,N_1766);
or U2196 (N_2196,N_1222,N_1413);
nand U2197 (N_2197,N_1712,N_1614);
nand U2198 (N_2198,N_1710,N_1227);
and U2199 (N_2199,N_1471,N_1208);
nor U2200 (N_2200,N_1243,N_1721);
nand U2201 (N_2201,N_1644,N_1763);
nor U2202 (N_2202,N_1274,N_1529);
xnor U2203 (N_2203,N_1441,N_1242);
nand U2204 (N_2204,N_1429,N_1694);
nand U2205 (N_2205,N_1577,N_1370);
and U2206 (N_2206,N_1512,N_1504);
nand U2207 (N_2207,N_1499,N_1395);
nand U2208 (N_2208,N_1503,N_1311);
nand U2209 (N_2209,N_1235,N_1568);
nand U2210 (N_2210,N_1665,N_1489);
or U2211 (N_2211,N_1639,N_1515);
nor U2212 (N_2212,N_1364,N_1347);
or U2213 (N_2213,N_1569,N_1246);
nor U2214 (N_2214,N_1206,N_1649);
xnor U2215 (N_2215,N_1256,N_1430);
nand U2216 (N_2216,N_1204,N_1551);
nor U2217 (N_2217,N_1358,N_1380);
or U2218 (N_2218,N_1713,N_1222);
or U2219 (N_2219,N_1714,N_1556);
nor U2220 (N_2220,N_1684,N_1306);
nor U2221 (N_2221,N_1734,N_1422);
or U2222 (N_2222,N_1617,N_1397);
and U2223 (N_2223,N_1282,N_1684);
nor U2224 (N_2224,N_1218,N_1491);
and U2225 (N_2225,N_1244,N_1498);
nor U2226 (N_2226,N_1386,N_1345);
nor U2227 (N_2227,N_1734,N_1611);
or U2228 (N_2228,N_1526,N_1613);
and U2229 (N_2229,N_1506,N_1254);
nor U2230 (N_2230,N_1762,N_1747);
and U2231 (N_2231,N_1442,N_1629);
nand U2232 (N_2232,N_1506,N_1539);
and U2233 (N_2233,N_1772,N_1203);
or U2234 (N_2234,N_1675,N_1444);
and U2235 (N_2235,N_1254,N_1343);
nor U2236 (N_2236,N_1420,N_1272);
nor U2237 (N_2237,N_1696,N_1674);
nand U2238 (N_2238,N_1680,N_1760);
nor U2239 (N_2239,N_1645,N_1733);
nor U2240 (N_2240,N_1548,N_1485);
and U2241 (N_2241,N_1696,N_1398);
nor U2242 (N_2242,N_1242,N_1383);
nand U2243 (N_2243,N_1458,N_1255);
and U2244 (N_2244,N_1551,N_1696);
nand U2245 (N_2245,N_1359,N_1701);
nor U2246 (N_2246,N_1590,N_1672);
nand U2247 (N_2247,N_1342,N_1392);
nand U2248 (N_2248,N_1619,N_1785);
or U2249 (N_2249,N_1468,N_1496);
nor U2250 (N_2250,N_1772,N_1561);
and U2251 (N_2251,N_1532,N_1343);
nand U2252 (N_2252,N_1433,N_1781);
or U2253 (N_2253,N_1508,N_1391);
or U2254 (N_2254,N_1453,N_1287);
or U2255 (N_2255,N_1319,N_1425);
nor U2256 (N_2256,N_1472,N_1438);
nand U2257 (N_2257,N_1347,N_1661);
and U2258 (N_2258,N_1757,N_1334);
or U2259 (N_2259,N_1298,N_1668);
and U2260 (N_2260,N_1244,N_1772);
nor U2261 (N_2261,N_1584,N_1435);
xnor U2262 (N_2262,N_1468,N_1545);
or U2263 (N_2263,N_1622,N_1795);
and U2264 (N_2264,N_1288,N_1627);
or U2265 (N_2265,N_1517,N_1538);
or U2266 (N_2266,N_1200,N_1704);
and U2267 (N_2267,N_1306,N_1434);
nor U2268 (N_2268,N_1649,N_1237);
xnor U2269 (N_2269,N_1708,N_1360);
and U2270 (N_2270,N_1433,N_1233);
nand U2271 (N_2271,N_1420,N_1221);
and U2272 (N_2272,N_1335,N_1795);
nand U2273 (N_2273,N_1246,N_1306);
and U2274 (N_2274,N_1778,N_1211);
and U2275 (N_2275,N_1360,N_1493);
nand U2276 (N_2276,N_1792,N_1321);
nor U2277 (N_2277,N_1584,N_1744);
nand U2278 (N_2278,N_1610,N_1672);
nand U2279 (N_2279,N_1759,N_1732);
nand U2280 (N_2280,N_1322,N_1574);
and U2281 (N_2281,N_1675,N_1388);
nand U2282 (N_2282,N_1774,N_1275);
and U2283 (N_2283,N_1708,N_1788);
and U2284 (N_2284,N_1595,N_1205);
nor U2285 (N_2285,N_1242,N_1542);
or U2286 (N_2286,N_1400,N_1463);
nand U2287 (N_2287,N_1607,N_1390);
xnor U2288 (N_2288,N_1215,N_1478);
nor U2289 (N_2289,N_1449,N_1240);
and U2290 (N_2290,N_1337,N_1422);
xor U2291 (N_2291,N_1214,N_1327);
and U2292 (N_2292,N_1561,N_1760);
and U2293 (N_2293,N_1299,N_1783);
or U2294 (N_2294,N_1644,N_1392);
and U2295 (N_2295,N_1744,N_1253);
or U2296 (N_2296,N_1406,N_1267);
and U2297 (N_2297,N_1521,N_1384);
or U2298 (N_2298,N_1787,N_1426);
and U2299 (N_2299,N_1292,N_1266);
or U2300 (N_2300,N_1483,N_1399);
nor U2301 (N_2301,N_1723,N_1569);
and U2302 (N_2302,N_1620,N_1312);
or U2303 (N_2303,N_1268,N_1676);
and U2304 (N_2304,N_1356,N_1302);
or U2305 (N_2305,N_1477,N_1465);
nor U2306 (N_2306,N_1442,N_1681);
nor U2307 (N_2307,N_1267,N_1335);
and U2308 (N_2308,N_1375,N_1555);
nor U2309 (N_2309,N_1278,N_1339);
and U2310 (N_2310,N_1263,N_1323);
nor U2311 (N_2311,N_1218,N_1646);
nor U2312 (N_2312,N_1559,N_1447);
and U2313 (N_2313,N_1461,N_1475);
and U2314 (N_2314,N_1302,N_1393);
and U2315 (N_2315,N_1786,N_1203);
nand U2316 (N_2316,N_1329,N_1374);
or U2317 (N_2317,N_1544,N_1469);
nor U2318 (N_2318,N_1568,N_1375);
nand U2319 (N_2319,N_1429,N_1403);
xnor U2320 (N_2320,N_1495,N_1701);
and U2321 (N_2321,N_1743,N_1276);
and U2322 (N_2322,N_1496,N_1443);
or U2323 (N_2323,N_1503,N_1430);
or U2324 (N_2324,N_1442,N_1262);
nor U2325 (N_2325,N_1684,N_1315);
and U2326 (N_2326,N_1254,N_1431);
xnor U2327 (N_2327,N_1464,N_1551);
nor U2328 (N_2328,N_1268,N_1263);
or U2329 (N_2329,N_1314,N_1268);
or U2330 (N_2330,N_1427,N_1337);
and U2331 (N_2331,N_1492,N_1291);
nor U2332 (N_2332,N_1735,N_1798);
nor U2333 (N_2333,N_1654,N_1347);
nand U2334 (N_2334,N_1449,N_1506);
xor U2335 (N_2335,N_1203,N_1408);
nor U2336 (N_2336,N_1355,N_1599);
nor U2337 (N_2337,N_1273,N_1603);
nand U2338 (N_2338,N_1370,N_1656);
nand U2339 (N_2339,N_1425,N_1678);
and U2340 (N_2340,N_1640,N_1797);
and U2341 (N_2341,N_1572,N_1285);
xor U2342 (N_2342,N_1288,N_1610);
and U2343 (N_2343,N_1600,N_1608);
nor U2344 (N_2344,N_1616,N_1200);
and U2345 (N_2345,N_1372,N_1226);
or U2346 (N_2346,N_1284,N_1736);
and U2347 (N_2347,N_1507,N_1278);
nand U2348 (N_2348,N_1533,N_1564);
nor U2349 (N_2349,N_1351,N_1207);
and U2350 (N_2350,N_1208,N_1275);
or U2351 (N_2351,N_1673,N_1222);
nand U2352 (N_2352,N_1643,N_1781);
nand U2353 (N_2353,N_1209,N_1598);
nor U2354 (N_2354,N_1541,N_1537);
nand U2355 (N_2355,N_1571,N_1746);
nor U2356 (N_2356,N_1727,N_1548);
nor U2357 (N_2357,N_1292,N_1401);
or U2358 (N_2358,N_1268,N_1742);
nand U2359 (N_2359,N_1345,N_1461);
nor U2360 (N_2360,N_1662,N_1273);
or U2361 (N_2361,N_1577,N_1794);
or U2362 (N_2362,N_1770,N_1501);
nand U2363 (N_2363,N_1410,N_1470);
nor U2364 (N_2364,N_1607,N_1582);
xor U2365 (N_2365,N_1428,N_1489);
and U2366 (N_2366,N_1215,N_1243);
or U2367 (N_2367,N_1271,N_1297);
nor U2368 (N_2368,N_1287,N_1326);
nand U2369 (N_2369,N_1408,N_1334);
and U2370 (N_2370,N_1281,N_1746);
nor U2371 (N_2371,N_1393,N_1247);
or U2372 (N_2372,N_1321,N_1790);
xor U2373 (N_2373,N_1749,N_1494);
nand U2374 (N_2374,N_1748,N_1799);
nand U2375 (N_2375,N_1792,N_1723);
nor U2376 (N_2376,N_1482,N_1556);
nor U2377 (N_2377,N_1778,N_1545);
and U2378 (N_2378,N_1705,N_1689);
nor U2379 (N_2379,N_1521,N_1427);
and U2380 (N_2380,N_1391,N_1626);
and U2381 (N_2381,N_1483,N_1595);
or U2382 (N_2382,N_1374,N_1259);
nand U2383 (N_2383,N_1273,N_1319);
or U2384 (N_2384,N_1373,N_1258);
nand U2385 (N_2385,N_1460,N_1321);
and U2386 (N_2386,N_1581,N_1299);
or U2387 (N_2387,N_1577,N_1686);
xor U2388 (N_2388,N_1326,N_1377);
nor U2389 (N_2389,N_1244,N_1574);
and U2390 (N_2390,N_1794,N_1524);
nand U2391 (N_2391,N_1749,N_1500);
nor U2392 (N_2392,N_1671,N_1206);
and U2393 (N_2393,N_1232,N_1516);
or U2394 (N_2394,N_1362,N_1604);
nand U2395 (N_2395,N_1498,N_1280);
and U2396 (N_2396,N_1244,N_1552);
nor U2397 (N_2397,N_1393,N_1201);
or U2398 (N_2398,N_1426,N_1453);
xor U2399 (N_2399,N_1725,N_1795);
or U2400 (N_2400,N_1883,N_1965);
and U2401 (N_2401,N_2392,N_2062);
nand U2402 (N_2402,N_2336,N_1888);
or U2403 (N_2403,N_2399,N_2226);
and U2404 (N_2404,N_1946,N_1818);
nor U2405 (N_2405,N_2203,N_1939);
nor U2406 (N_2406,N_2111,N_2260);
nand U2407 (N_2407,N_2097,N_2123);
nor U2408 (N_2408,N_2258,N_2051);
or U2409 (N_2409,N_1897,N_2214);
and U2410 (N_2410,N_2301,N_2177);
or U2411 (N_2411,N_1985,N_1806);
and U2412 (N_2412,N_1983,N_2371);
nor U2413 (N_2413,N_2311,N_2199);
and U2414 (N_2414,N_2144,N_2181);
or U2415 (N_2415,N_2276,N_2208);
nand U2416 (N_2416,N_2356,N_2113);
nand U2417 (N_2417,N_2143,N_2202);
and U2418 (N_2418,N_1866,N_2188);
nor U2419 (N_2419,N_2344,N_1921);
and U2420 (N_2420,N_2076,N_2159);
or U2421 (N_2421,N_2384,N_1846);
nor U2422 (N_2422,N_2207,N_1932);
nand U2423 (N_2423,N_2006,N_1831);
nand U2424 (N_2424,N_2066,N_1892);
nand U2425 (N_2425,N_2286,N_2186);
xor U2426 (N_2426,N_2105,N_2281);
nor U2427 (N_2427,N_2334,N_1978);
and U2428 (N_2428,N_2237,N_1802);
nor U2429 (N_2429,N_2102,N_2138);
xor U2430 (N_2430,N_1886,N_1904);
nor U2431 (N_2431,N_2329,N_2124);
xor U2432 (N_2432,N_2103,N_1996);
or U2433 (N_2433,N_1926,N_2373);
nand U2434 (N_2434,N_2232,N_1875);
and U2435 (N_2435,N_2331,N_2023);
nor U2436 (N_2436,N_2034,N_2026);
xor U2437 (N_2437,N_1857,N_2121);
and U2438 (N_2438,N_2139,N_2067);
nand U2439 (N_2439,N_2055,N_2095);
and U2440 (N_2440,N_1872,N_2291);
or U2441 (N_2441,N_1879,N_2312);
or U2442 (N_2442,N_2154,N_2212);
nand U2443 (N_2443,N_2283,N_1943);
or U2444 (N_2444,N_2321,N_2092);
nor U2445 (N_2445,N_1936,N_2394);
or U2446 (N_2446,N_1925,N_2059);
and U2447 (N_2447,N_2350,N_1972);
or U2448 (N_2448,N_1917,N_1870);
or U2449 (N_2449,N_1922,N_2275);
and U2450 (N_2450,N_2145,N_2249);
and U2451 (N_2451,N_1986,N_2183);
and U2452 (N_2452,N_1848,N_2146);
and U2453 (N_2453,N_2036,N_2018);
nor U2454 (N_2454,N_1938,N_1861);
and U2455 (N_2455,N_1902,N_1898);
nand U2456 (N_2456,N_1804,N_1919);
nand U2457 (N_2457,N_1858,N_2106);
nor U2458 (N_2458,N_2250,N_2206);
nor U2459 (N_2459,N_1997,N_2288);
and U2460 (N_2460,N_2169,N_2358);
nand U2461 (N_2461,N_2068,N_2315);
or U2462 (N_2462,N_1825,N_2219);
or U2463 (N_2463,N_2090,N_2192);
or U2464 (N_2464,N_2369,N_2011);
nand U2465 (N_2465,N_2343,N_1918);
or U2466 (N_2466,N_2112,N_1871);
or U2467 (N_2467,N_2222,N_1891);
and U2468 (N_2468,N_1819,N_2171);
nand U2469 (N_2469,N_1821,N_2099);
nand U2470 (N_2470,N_2221,N_2104);
and U2471 (N_2471,N_2077,N_2367);
or U2472 (N_2472,N_2255,N_2048);
and U2473 (N_2473,N_2108,N_2082);
and U2474 (N_2474,N_2056,N_2125);
xor U2475 (N_2475,N_2282,N_1882);
nand U2476 (N_2476,N_2253,N_2040);
and U2477 (N_2477,N_2119,N_1878);
or U2478 (N_2478,N_2323,N_2267);
or U2479 (N_2479,N_2337,N_2107);
nor U2480 (N_2480,N_2053,N_2341);
nor U2481 (N_2481,N_2047,N_1828);
nor U2482 (N_2482,N_2028,N_2225);
and U2483 (N_2483,N_1993,N_2012);
nand U2484 (N_2484,N_1877,N_2167);
and U2485 (N_2485,N_1853,N_2080);
nor U2486 (N_2486,N_1907,N_2101);
and U2487 (N_2487,N_1906,N_1817);
nor U2488 (N_2488,N_2294,N_2382);
and U2489 (N_2489,N_1952,N_2269);
nor U2490 (N_2490,N_1976,N_2293);
nand U2491 (N_2491,N_2128,N_1987);
and U2492 (N_2492,N_2148,N_2360);
nand U2493 (N_2493,N_2016,N_2365);
nand U2494 (N_2494,N_2284,N_2228);
and U2495 (N_2495,N_1933,N_2393);
nand U2496 (N_2496,N_2085,N_1984);
or U2497 (N_2497,N_2227,N_1865);
or U2498 (N_2498,N_2003,N_2020);
nand U2499 (N_2499,N_2240,N_2239);
nand U2500 (N_2500,N_2335,N_2060);
nand U2501 (N_2501,N_2300,N_1931);
or U2502 (N_2502,N_1900,N_2378);
nand U2503 (N_2503,N_2210,N_1814);
xor U2504 (N_2504,N_1957,N_2326);
nand U2505 (N_2505,N_1830,N_2141);
nor U2506 (N_2506,N_1839,N_2245);
and U2507 (N_2507,N_1851,N_2093);
nand U2508 (N_2508,N_2271,N_2140);
and U2509 (N_2509,N_2084,N_2218);
nand U2510 (N_2510,N_1948,N_2109);
and U2511 (N_2511,N_2024,N_2162);
and U2512 (N_2512,N_2175,N_2096);
nand U2513 (N_2513,N_2390,N_1927);
or U2514 (N_2514,N_1940,N_2303);
and U2515 (N_2515,N_2120,N_2320);
xnor U2516 (N_2516,N_2070,N_2174);
nand U2517 (N_2517,N_2327,N_2285);
or U2518 (N_2518,N_1915,N_1805);
nor U2519 (N_2519,N_2074,N_2347);
xnor U2520 (N_2520,N_1994,N_2165);
and U2521 (N_2521,N_1955,N_2355);
or U2522 (N_2522,N_2304,N_1868);
nor U2523 (N_2523,N_1855,N_1937);
nor U2524 (N_2524,N_1971,N_2058);
and U2525 (N_2525,N_2163,N_2265);
nor U2526 (N_2526,N_2223,N_2340);
nand U2527 (N_2527,N_2397,N_1808);
xor U2528 (N_2528,N_2242,N_2098);
and U2529 (N_2529,N_1956,N_1944);
nand U2530 (N_2530,N_2262,N_1884);
nor U2531 (N_2531,N_2130,N_2037);
xnor U2532 (N_2532,N_2000,N_1977);
nand U2533 (N_2533,N_2254,N_2158);
nand U2534 (N_2534,N_2061,N_1823);
or U2535 (N_2535,N_2362,N_1842);
or U2536 (N_2536,N_2180,N_2266);
and U2537 (N_2537,N_2117,N_2160);
or U2538 (N_2538,N_2178,N_2135);
nand U2539 (N_2539,N_2359,N_1905);
or U2540 (N_2540,N_2087,N_1838);
nand U2541 (N_2541,N_2019,N_2234);
nor U2542 (N_2542,N_1881,N_2328);
and U2543 (N_2543,N_1887,N_1923);
or U2544 (N_2544,N_2136,N_1850);
nor U2545 (N_2545,N_1859,N_2306);
or U2546 (N_2546,N_2314,N_1809);
and U2547 (N_2547,N_2134,N_2372);
nor U2548 (N_2548,N_2263,N_2187);
nand U2549 (N_2549,N_2235,N_1928);
and U2550 (N_2550,N_2147,N_2049);
or U2551 (N_2551,N_2078,N_2391);
nor U2552 (N_2552,N_1960,N_1822);
or U2553 (N_2553,N_2027,N_2010);
xor U2554 (N_2554,N_2172,N_1934);
and U2555 (N_2555,N_1832,N_1880);
nor U2556 (N_2556,N_1949,N_2065);
and U2557 (N_2557,N_2116,N_1967);
nand U2558 (N_2558,N_2357,N_1980);
nand U2559 (N_2559,N_1899,N_2377);
and U2560 (N_2560,N_2149,N_2013);
and U2561 (N_2561,N_2368,N_2088);
or U2562 (N_2562,N_2273,N_2386);
nor U2563 (N_2563,N_2342,N_1837);
xnor U2564 (N_2564,N_2002,N_1836);
or U2565 (N_2565,N_1969,N_2057);
nor U2566 (N_2566,N_1950,N_2071);
nand U2567 (N_2567,N_1910,N_2161);
nor U2568 (N_2568,N_2277,N_2316);
xnor U2569 (N_2569,N_2079,N_1992);
nand U2570 (N_2570,N_2339,N_2094);
or U2571 (N_2571,N_1889,N_2072);
nand U2572 (N_2572,N_1862,N_1867);
xor U2573 (N_2573,N_2122,N_1930);
and U2574 (N_2574,N_2319,N_1901);
nand U2575 (N_2575,N_1841,N_2173);
xnor U2576 (N_2576,N_2398,N_2025);
and U2577 (N_2577,N_2164,N_2153);
xor U2578 (N_2578,N_1869,N_1954);
nor U2579 (N_2579,N_1909,N_1893);
xnor U2580 (N_2580,N_2274,N_2252);
or U2581 (N_2581,N_2083,N_2166);
or U2582 (N_2582,N_2388,N_1833);
nand U2583 (N_2583,N_1966,N_2195);
and U2584 (N_2584,N_2395,N_2015);
or U2585 (N_2585,N_2209,N_2259);
nor U2586 (N_2586,N_1968,N_2270);
or U2587 (N_2587,N_2264,N_1981);
nand U2588 (N_2588,N_2333,N_2224);
xnor U2589 (N_2589,N_1801,N_1942);
or U2590 (N_2590,N_2137,N_2182);
nor U2591 (N_2591,N_2292,N_1912);
nor U2592 (N_2592,N_2200,N_1908);
nor U2593 (N_2593,N_2132,N_2041);
and U2594 (N_2594,N_2313,N_2380);
nor U2595 (N_2595,N_2290,N_2115);
and U2596 (N_2596,N_1803,N_2194);
or U2597 (N_2597,N_1963,N_2152);
xor U2598 (N_2598,N_2004,N_2091);
nand U2599 (N_2599,N_2353,N_2133);
xnor U2600 (N_2600,N_2230,N_2370);
nor U2601 (N_2601,N_2309,N_1824);
nand U2602 (N_2602,N_2296,N_1820);
nand U2603 (N_2603,N_1953,N_2032);
nand U2604 (N_2604,N_1945,N_2381);
or U2605 (N_2605,N_2150,N_1876);
nand U2606 (N_2606,N_2063,N_1826);
and U2607 (N_2607,N_2349,N_2042);
and U2608 (N_2608,N_2366,N_1852);
nor U2609 (N_2609,N_2376,N_2008);
nor U2610 (N_2610,N_1811,N_2351);
nor U2611 (N_2611,N_2151,N_2324);
nor U2612 (N_2612,N_2215,N_2089);
xor U2613 (N_2613,N_2383,N_2044);
and U2614 (N_2614,N_2193,N_1844);
nand U2615 (N_2615,N_2029,N_2389);
nand U2616 (N_2616,N_1964,N_2318);
nand U2617 (N_2617,N_2075,N_1947);
nand U2618 (N_2618,N_2216,N_2142);
or U2619 (N_2619,N_2302,N_2014);
xnor U2620 (N_2620,N_2069,N_2211);
or U2621 (N_2621,N_2196,N_1863);
and U2622 (N_2622,N_2190,N_2217);
and U2623 (N_2623,N_2043,N_1815);
xnor U2624 (N_2624,N_1991,N_2305);
nor U2625 (N_2625,N_2131,N_2021);
xnor U2626 (N_2626,N_1975,N_1911);
and U2627 (N_2627,N_2031,N_1913);
and U2628 (N_2628,N_1916,N_1988);
nand U2629 (N_2629,N_2272,N_2241);
nand U2630 (N_2630,N_1834,N_2033);
or U2631 (N_2631,N_2379,N_2114);
nand U2632 (N_2632,N_2039,N_2050);
xor U2633 (N_2633,N_2198,N_1990);
nand U2634 (N_2634,N_1827,N_2385);
nor U2635 (N_2635,N_1995,N_1941);
nand U2636 (N_2636,N_2201,N_2155);
or U2637 (N_2637,N_1847,N_1962);
nand U2638 (N_2638,N_2354,N_1895);
or U2639 (N_2639,N_2236,N_2278);
and U2640 (N_2640,N_1959,N_2268);
nor U2641 (N_2641,N_2352,N_1813);
nand U2642 (N_2642,N_1840,N_2127);
nand U2643 (N_2643,N_2157,N_2297);
or U2644 (N_2644,N_2345,N_2213);
xor U2645 (N_2645,N_1989,N_2396);
nand U2646 (N_2646,N_2364,N_2257);
or U2647 (N_2647,N_2387,N_2322);
nand U2648 (N_2648,N_1845,N_2045);
nand U2649 (N_2649,N_2247,N_2289);
xnor U2650 (N_2650,N_2035,N_2298);
or U2651 (N_2651,N_2046,N_1903);
and U2652 (N_2652,N_2204,N_1961);
nand U2653 (N_2653,N_1974,N_1951);
nand U2654 (N_2654,N_2007,N_2005);
and U2655 (N_2655,N_2038,N_1920);
and U2656 (N_2656,N_2110,N_1999);
nor U2657 (N_2657,N_1843,N_2001);
nor U2658 (N_2658,N_2361,N_1810);
and U2659 (N_2659,N_1812,N_2244);
and U2660 (N_2660,N_1973,N_2179);
and U2661 (N_2661,N_1800,N_2299);
and U2662 (N_2662,N_2052,N_2022);
nand U2663 (N_2663,N_2220,N_2086);
nand U2664 (N_2664,N_1896,N_1929);
or U2665 (N_2665,N_1982,N_2184);
and U2666 (N_2666,N_2374,N_2229);
and U2667 (N_2667,N_2176,N_2348);
or U2668 (N_2668,N_1849,N_2317);
or U2669 (N_2669,N_1914,N_1890);
and U2670 (N_2670,N_2081,N_2129);
nand U2671 (N_2671,N_2310,N_1807);
xor U2672 (N_2672,N_2248,N_2295);
and U2673 (N_2673,N_2233,N_2073);
or U2674 (N_2674,N_2168,N_1856);
nand U2675 (N_2675,N_2243,N_1958);
xor U2676 (N_2676,N_1829,N_2308);
or U2677 (N_2677,N_2375,N_2261);
or U2678 (N_2678,N_1935,N_2256);
or U2679 (N_2679,N_1816,N_2307);
nand U2680 (N_2680,N_2170,N_1998);
nor U2681 (N_2681,N_2126,N_2238);
and U2682 (N_2682,N_1970,N_2346);
and U2683 (N_2683,N_2251,N_1885);
nor U2684 (N_2684,N_2280,N_2231);
nor U2685 (N_2685,N_2017,N_1979);
nand U2686 (N_2686,N_1860,N_2205);
or U2687 (N_2687,N_2332,N_2118);
nand U2688 (N_2688,N_2054,N_1873);
and U2689 (N_2689,N_2246,N_1924);
and U2690 (N_2690,N_2191,N_1874);
nand U2691 (N_2691,N_2279,N_2325);
and U2692 (N_2692,N_2100,N_2185);
or U2693 (N_2693,N_2287,N_1894);
nand U2694 (N_2694,N_2338,N_2189);
and U2695 (N_2695,N_2363,N_2197);
and U2696 (N_2696,N_2156,N_2009);
nor U2697 (N_2697,N_2330,N_1835);
xor U2698 (N_2698,N_1864,N_2030);
nand U2699 (N_2699,N_1854,N_2064);
xor U2700 (N_2700,N_1932,N_2358);
and U2701 (N_2701,N_2213,N_1809);
or U2702 (N_2702,N_1810,N_2092);
xnor U2703 (N_2703,N_2066,N_2350);
and U2704 (N_2704,N_2316,N_1996);
nand U2705 (N_2705,N_2016,N_2304);
xor U2706 (N_2706,N_1952,N_1853);
nor U2707 (N_2707,N_2284,N_2357);
or U2708 (N_2708,N_2058,N_2133);
nor U2709 (N_2709,N_1999,N_2241);
or U2710 (N_2710,N_2077,N_1973);
or U2711 (N_2711,N_1853,N_2196);
and U2712 (N_2712,N_2049,N_2129);
and U2713 (N_2713,N_2381,N_1958);
or U2714 (N_2714,N_1972,N_2045);
nand U2715 (N_2715,N_1838,N_1993);
and U2716 (N_2716,N_1950,N_1865);
nor U2717 (N_2717,N_2047,N_2226);
or U2718 (N_2718,N_2057,N_2159);
xor U2719 (N_2719,N_2019,N_1932);
and U2720 (N_2720,N_1870,N_1952);
xor U2721 (N_2721,N_2243,N_1834);
or U2722 (N_2722,N_2377,N_1810);
nand U2723 (N_2723,N_1811,N_1941);
or U2724 (N_2724,N_2310,N_2162);
nor U2725 (N_2725,N_2388,N_2175);
nand U2726 (N_2726,N_2209,N_1828);
or U2727 (N_2727,N_2004,N_1895);
nand U2728 (N_2728,N_1930,N_1829);
nor U2729 (N_2729,N_2090,N_2300);
nand U2730 (N_2730,N_2261,N_2226);
and U2731 (N_2731,N_2246,N_2319);
nand U2732 (N_2732,N_2021,N_1898);
nand U2733 (N_2733,N_1903,N_2172);
nor U2734 (N_2734,N_2102,N_2352);
nand U2735 (N_2735,N_2370,N_1844);
nand U2736 (N_2736,N_2194,N_2003);
or U2737 (N_2737,N_2280,N_2105);
nand U2738 (N_2738,N_2000,N_2167);
or U2739 (N_2739,N_2086,N_2029);
and U2740 (N_2740,N_2271,N_1922);
or U2741 (N_2741,N_2333,N_1880);
nand U2742 (N_2742,N_2198,N_1858);
nor U2743 (N_2743,N_2179,N_1823);
nand U2744 (N_2744,N_2378,N_2168);
xor U2745 (N_2745,N_1826,N_2235);
and U2746 (N_2746,N_1893,N_1911);
nand U2747 (N_2747,N_2329,N_2064);
nor U2748 (N_2748,N_2069,N_2071);
nor U2749 (N_2749,N_1822,N_2393);
nor U2750 (N_2750,N_2254,N_2042);
nor U2751 (N_2751,N_2192,N_2010);
and U2752 (N_2752,N_1852,N_2015);
and U2753 (N_2753,N_2370,N_2383);
and U2754 (N_2754,N_2313,N_1973);
and U2755 (N_2755,N_2378,N_1803);
and U2756 (N_2756,N_2279,N_1925);
or U2757 (N_2757,N_2249,N_2281);
nand U2758 (N_2758,N_2190,N_1940);
nand U2759 (N_2759,N_1961,N_1904);
nor U2760 (N_2760,N_2324,N_2145);
xor U2761 (N_2761,N_2191,N_1898);
and U2762 (N_2762,N_2191,N_1982);
nor U2763 (N_2763,N_2030,N_2200);
and U2764 (N_2764,N_2261,N_1987);
xor U2765 (N_2765,N_1915,N_2188);
nor U2766 (N_2766,N_1976,N_2281);
or U2767 (N_2767,N_2116,N_2361);
or U2768 (N_2768,N_2395,N_1938);
and U2769 (N_2769,N_2389,N_2252);
nand U2770 (N_2770,N_2363,N_2389);
or U2771 (N_2771,N_1966,N_2247);
and U2772 (N_2772,N_1824,N_2228);
or U2773 (N_2773,N_1892,N_2286);
nor U2774 (N_2774,N_1951,N_2133);
or U2775 (N_2775,N_2018,N_1934);
or U2776 (N_2776,N_1892,N_2382);
nor U2777 (N_2777,N_2083,N_1853);
nor U2778 (N_2778,N_2045,N_1985);
and U2779 (N_2779,N_2140,N_2305);
and U2780 (N_2780,N_1815,N_1985);
nor U2781 (N_2781,N_2375,N_2364);
xnor U2782 (N_2782,N_1933,N_2009);
and U2783 (N_2783,N_2238,N_2197);
and U2784 (N_2784,N_1803,N_2244);
and U2785 (N_2785,N_2107,N_2256);
nor U2786 (N_2786,N_1890,N_2073);
nand U2787 (N_2787,N_1965,N_1874);
and U2788 (N_2788,N_1908,N_2287);
or U2789 (N_2789,N_1997,N_1947);
nand U2790 (N_2790,N_1814,N_2176);
and U2791 (N_2791,N_1914,N_2219);
and U2792 (N_2792,N_1979,N_2113);
nor U2793 (N_2793,N_2109,N_2336);
nand U2794 (N_2794,N_1929,N_1832);
and U2795 (N_2795,N_2100,N_2068);
or U2796 (N_2796,N_1950,N_2298);
nand U2797 (N_2797,N_2243,N_2265);
xnor U2798 (N_2798,N_2019,N_2070);
and U2799 (N_2799,N_2036,N_2191);
nor U2800 (N_2800,N_2137,N_1874);
nand U2801 (N_2801,N_1899,N_2079);
nand U2802 (N_2802,N_2012,N_1961);
and U2803 (N_2803,N_2334,N_2140);
and U2804 (N_2804,N_2067,N_1835);
or U2805 (N_2805,N_1834,N_1950);
and U2806 (N_2806,N_1972,N_1853);
nand U2807 (N_2807,N_2375,N_2329);
nand U2808 (N_2808,N_1819,N_2242);
xor U2809 (N_2809,N_1929,N_1918);
and U2810 (N_2810,N_1909,N_2017);
or U2811 (N_2811,N_2006,N_2163);
xor U2812 (N_2812,N_1823,N_2092);
nand U2813 (N_2813,N_2391,N_2298);
and U2814 (N_2814,N_1889,N_2129);
nand U2815 (N_2815,N_2122,N_2025);
or U2816 (N_2816,N_2358,N_2387);
nor U2817 (N_2817,N_2095,N_1891);
nor U2818 (N_2818,N_2074,N_2190);
and U2819 (N_2819,N_1805,N_2141);
or U2820 (N_2820,N_1846,N_2312);
or U2821 (N_2821,N_1850,N_2285);
nor U2822 (N_2822,N_2198,N_2184);
xnor U2823 (N_2823,N_1941,N_2364);
or U2824 (N_2824,N_2019,N_2328);
and U2825 (N_2825,N_2309,N_1838);
or U2826 (N_2826,N_2015,N_2235);
nor U2827 (N_2827,N_2065,N_2348);
or U2828 (N_2828,N_1819,N_2262);
nand U2829 (N_2829,N_2120,N_2002);
or U2830 (N_2830,N_2095,N_2212);
nand U2831 (N_2831,N_1809,N_2009);
nand U2832 (N_2832,N_1951,N_2251);
or U2833 (N_2833,N_1911,N_2141);
nor U2834 (N_2834,N_1891,N_2226);
and U2835 (N_2835,N_2398,N_2172);
nand U2836 (N_2836,N_2292,N_2092);
and U2837 (N_2837,N_2249,N_2282);
or U2838 (N_2838,N_2209,N_2261);
and U2839 (N_2839,N_2080,N_1911);
and U2840 (N_2840,N_1908,N_1832);
or U2841 (N_2841,N_1830,N_1872);
nor U2842 (N_2842,N_2062,N_2368);
nand U2843 (N_2843,N_2012,N_2179);
nor U2844 (N_2844,N_2364,N_1833);
or U2845 (N_2845,N_1886,N_2100);
and U2846 (N_2846,N_2308,N_2162);
nand U2847 (N_2847,N_2324,N_2353);
nor U2848 (N_2848,N_2363,N_2214);
and U2849 (N_2849,N_2358,N_2017);
and U2850 (N_2850,N_2301,N_1907);
or U2851 (N_2851,N_1942,N_1842);
and U2852 (N_2852,N_1998,N_2291);
and U2853 (N_2853,N_2094,N_2124);
or U2854 (N_2854,N_2063,N_2242);
xnor U2855 (N_2855,N_1806,N_2213);
or U2856 (N_2856,N_1952,N_1961);
or U2857 (N_2857,N_2180,N_1919);
nor U2858 (N_2858,N_1961,N_2365);
nor U2859 (N_2859,N_1926,N_2304);
or U2860 (N_2860,N_1948,N_2013);
xnor U2861 (N_2861,N_2033,N_2181);
and U2862 (N_2862,N_2263,N_2260);
or U2863 (N_2863,N_2210,N_1889);
xnor U2864 (N_2864,N_2359,N_2278);
nand U2865 (N_2865,N_2361,N_1927);
nor U2866 (N_2866,N_1942,N_2126);
xnor U2867 (N_2867,N_2209,N_2057);
or U2868 (N_2868,N_2005,N_2025);
or U2869 (N_2869,N_1977,N_2302);
nor U2870 (N_2870,N_2057,N_2365);
xor U2871 (N_2871,N_2131,N_2112);
nor U2872 (N_2872,N_2195,N_2391);
or U2873 (N_2873,N_1920,N_1880);
or U2874 (N_2874,N_2298,N_2079);
nor U2875 (N_2875,N_1835,N_1860);
xnor U2876 (N_2876,N_2287,N_2154);
nand U2877 (N_2877,N_2066,N_1856);
or U2878 (N_2878,N_1837,N_2120);
or U2879 (N_2879,N_1988,N_1907);
xor U2880 (N_2880,N_1997,N_2305);
nor U2881 (N_2881,N_1887,N_2193);
or U2882 (N_2882,N_1931,N_2008);
nand U2883 (N_2883,N_2166,N_1984);
and U2884 (N_2884,N_2396,N_2175);
or U2885 (N_2885,N_2029,N_2334);
nor U2886 (N_2886,N_2368,N_1937);
xnor U2887 (N_2887,N_2244,N_2186);
nor U2888 (N_2888,N_2055,N_1923);
and U2889 (N_2889,N_2015,N_2089);
xor U2890 (N_2890,N_1985,N_2068);
nor U2891 (N_2891,N_2396,N_1913);
or U2892 (N_2892,N_1840,N_2224);
xnor U2893 (N_2893,N_2015,N_1927);
or U2894 (N_2894,N_2069,N_2258);
or U2895 (N_2895,N_2176,N_1924);
or U2896 (N_2896,N_2149,N_2084);
and U2897 (N_2897,N_2254,N_1910);
nand U2898 (N_2898,N_2277,N_2364);
nand U2899 (N_2899,N_2002,N_2208);
nand U2900 (N_2900,N_1804,N_2199);
or U2901 (N_2901,N_2289,N_2223);
xnor U2902 (N_2902,N_1848,N_2025);
or U2903 (N_2903,N_2121,N_2172);
nand U2904 (N_2904,N_2033,N_2327);
or U2905 (N_2905,N_1861,N_2233);
or U2906 (N_2906,N_1937,N_2366);
and U2907 (N_2907,N_2142,N_2003);
and U2908 (N_2908,N_2168,N_2132);
or U2909 (N_2909,N_2226,N_2062);
xnor U2910 (N_2910,N_1861,N_2220);
nor U2911 (N_2911,N_1849,N_2392);
nand U2912 (N_2912,N_2336,N_1989);
and U2913 (N_2913,N_2397,N_2224);
nor U2914 (N_2914,N_2229,N_1842);
and U2915 (N_2915,N_2026,N_1842);
or U2916 (N_2916,N_1951,N_2232);
and U2917 (N_2917,N_2045,N_2113);
and U2918 (N_2918,N_2352,N_2190);
nor U2919 (N_2919,N_1905,N_1955);
and U2920 (N_2920,N_1996,N_2389);
and U2921 (N_2921,N_1920,N_1854);
and U2922 (N_2922,N_1902,N_1803);
nor U2923 (N_2923,N_1964,N_1963);
and U2924 (N_2924,N_1846,N_2115);
nor U2925 (N_2925,N_1812,N_2140);
nand U2926 (N_2926,N_1859,N_2148);
and U2927 (N_2927,N_2237,N_1967);
and U2928 (N_2928,N_1907,N_2222);
nor U2929 (N_2929,N_1918,N_1893);
nand U2930 (N_2930,N_1953,N_2222);
and U2931 (N_2931,N_2069,N_2123);
xor U2932 (N_2932,N_2300,N_2154);
and U2933 (N_2933,N_2206,N_2254);
and U2934 (N_2934,N_2327,N_1998);
nand U2935 (N_2935,N_1844,N_2081);
and U2936 (N_2936,N_2069,N_2197);
xnor U2937 (N_2937,N_1840,N_2035);
or U2938 (N_2938,N_2242,N_1836);
or U2939 (N_2939,N_2288,N_2061);
and U2940 (N_2940,N_2244,N_1950);
and U2941 (N_2941,N_1849,N_2125);
and U2942 (N_2942,N_1800,N_2089);
and U2943 (N_2943,N_1899,N_2082);
xor U2944 (N_2944,N_2363,N_2380);
nand U2945 (N_2945,N_2240,N_2023);
nor U2946 (N_2946,N_2151,N_2268);
or U2947 (N_2947,N_2270,N_2052);
nand U2948 (N_2948,N_2263,N_1955);
nor U2949 (N_2949,N_1835,N_2042);
and U2950 (N_2950,N_2005,N_1907);
nor U2951 (N_2951,N_2207,N_2312);
nand U2952 (N_2952,N_2196,N_1937);
nand U2953 (N_2953,N_2121,N_2091);
nand U2954 (N_2954,N_2092,N_2080);
and U2955 (N_2955,N_2127,N_2274);
or U2956 (N_2956,N_2318,N_2182);
nor U2957 (N_2957,N_2243,N_1809);
and U2958 (N_2958,N_2293,N_2217);
and U2959 (N_2959,N_2109,N_1926);
and U2960 (N_2960,N_1812,N_2208);
nand U2961 (N_2961,N_2174,N_2014);
nand U2962 (N_2962,N_1915,N_1853);
and U2963 (N_2963,N_2287,N_2216);
nand U2964 (N_2964,N_1872,N_2087);
nand U2965 (N_2965,N_2064,N_1982);
or U2966 (N_2966,N_2202,N_2359);
nor U2967 (N_2967,N_2280,N_2390);
or U2968 (N_2968,N_2083,N_1803);
or U2969 (N_2969,N_2081,N_2383);
xnor U2970 (N_2970,N_2015,N_2142);
nand U2971 (N_2971,N_2257,N_1860);
nand U2972 (N_2972,N_1910,N_1963);
nor U2973 (N_2973,N_2061,N_1932);
nand U2974 (N_2974,N_1801,N_2391);
xor U2975 (N_2975,N_2008,N_2011);
and U2976 (N_2976,N_2044,N_1918);
and U2977 (N_2977,N_2096,N_2035);
nand U2978 (N_2978,N_2217,N_2390);
and U2979 (N_2979,N_1983,N_2257);
or U2980 (N_2980,N_1999,N_2136);
nand U2981 (N_2981,N_1925,N_2361);
nor U2982 (N_2982,N_2331,N_2231);
nor U2983 (N_2983,N_1931,N_2270);
and U2984 (N_2984,N_1934,N_1860);
or U2985 (N_2985,N_2291,N_2033);
and U2986 (N_2986,N_2169,N_2248);
xnor U2987 (N_2987,N_2190,N_2030);
nand U2988 (N_2988,N_1967,N_2273);
nor U2989 (N_2989,N_2081,N_2255);
and U2990 (N_2990,N_2198,N_2162);
or U2991 (N_2991,N_1898,N_2324);
or U2992 (N_2992,N_2152,N_2339);
xnor U2993 (N_2993,N_2177,N_1922);
and U2994 (N_2994,N_2322,N_2159);
nand U2995 (N_2995,N_1951,N_1901);
xnor U2996 (N_2996,N_2207,N_2075);
or U2997 (N_2997,N_2193,N_1966);
nand U2998 (N_2998,N_2189,N_2150);
nor U2999 (N_2999,N_2339,N_2266);
nor UO_0 (O_0,N_2554,N_2827);
xnor UO_1 (O_1,N_2676,N_2994);
nor UO_2 (O_2,N_2490,N_2691);
or UO_3 (O_3,N_2956,N_2749);
or UO_4 (O_4,N_2760,N_2534);
or UO_5 (O_5,N_2654,N_2848);
or UO_6 (O_6,N_2682,N_2674);
or UO_7 (O_7,N_2401,N_2973);
or UO_8 (O_8,N_2750,N_2969);
nor UO_9 (O_9,N_2511,N_2884);
or UO_10 (O_10,N_2709,N_2469);
nor UO_11 (O_11,N_2810,N_2872);
xor UO_12 (O_12,N_2700,N_2640);
or UO_13 (O_13,N_2793,N_2896);
nor UO_14 (O_14,N_2651,N_2916);
nand UO_15 (O_15,N_2587,N_2719);
or UO_16 (O_16,N_2831,N_2561);
nand UO_17 (O_17,N_2404,N_2656);
nand UO_18 (O_18,N_2608,N_2781);
xnor UO_19 (O_19,N_2443,N_2703);
or UO_20 (O_20,N_2935,N_2641);
nand UO_21 (O_21,N_2958,N_2509);
or UO_22 (O_22,N_2748,N_2697);
nor UO_23 (O_23,N_2966,N_2786);
nor UO_24 (O_24,N_2811,N_2938);
nand UO_25 (O_25,N_2742,N_2413);
nand UO_26 (O_26,N_2594,N_2568);
and UO_27 (O_27,N_2504,N_2463);
nand UO_28 (O_28,N_2814,N_2546);
nor UO_29 (O_29,N_2930,N_2495);
nor UO_30 (O_30,N_2454,N_2537);
nand UO_31 (O_31,N_2763,N_2430);
nand UO_32 (O_32,N_2970,N_2677);
nand UO_33 (O_33,N_2954,N_2602);
and UO_34 (O_34,N_2738,N_2788);
nor UO_35 (O_35,N_2552,N_2411);
nand UO_36 (O_36,N_2603,N_2455);
nand UO_37 (O_37,N_2532,N_2550);
or UO_38 (O_38,N_2467,N_2657);
nor UO_39 (O_39,N_2575,N_2542);
or UO_40 (O_40,N_2426,N_2687);
nor UO_41 (O_41,N_2547,N_2835);
nand UO_42 (O_42,N_2451,N_2672);
xor UO_43 (O_43,N_2637,N_2799);
xor UO_44 (O_44,N_2609,N_2984);
nand UO_45 (O_45,N_2869,N_2435);
xor UO_46 (O_46,N_2658,N_2620);
and UO_47 (O_47,N_2744,N_2596);
nor UO_48 (O_48,N_2864,N_2861);
nor UO_49 (O_49,N_2647,N_2929);
and UO_50 (O_50,N_2502,N_2485);
nand UO_51 (O_51,N_2478,N_2421);
and UO_52 (O_52,N_2758,N_2695);
and UO_53 (O_53,N_2424,N_2645);
and UO_54 (O_54,N_2418,N_2733);
nor UO_55 (O_55,N_2627,N_2937);
nor UO_56 (O_56,N_2458,N_2735);
or UO_57 (O_57,N_2655,N_2952);
nor UO_58 (O_58,N_2518,N_2834);
or UO_59 (O_59,N_2795,N_2907);
nand UO_60 (O_60,N_2803,N_2425);
nor UO_61 (O_61,N_2584,N_2601);
and UO_62 (O_62,N_2633,N_2809);
or UO_63 (O_63,N_2711,N_2959);
and UO_64 (O_64,N_2893,N_2898);
or UO_65 (O_65,N_2871,N_2901);
nor UO_66 (O_66,N_2447,N_2612);
nor UO_67 (O_67,N_2648,N_2948);
or UO_68 (O_68,N_2432,N_2897);
or UO_69 (O_69,N_2420,N_2885);
or UO_70 (O_70,N_2888,N_2974);
or UO_71 (O_71,N_2611,N_2494);
nand UO_72 (O_72,N_2780,N_2972);
nand UO_73 (O_73,N_2999,N_2510);
nor UO_74 (O_74,N_2556,N_2644);
xor UO_75 (O_75,N_2823,N_2774);
nor UO_76 (O_76,N_2820,N_2626);
nor UO_77 (O_77,N_2488,N_2940);
and UO_78 (O_78,N_2993,N_2673);
nor UO_79 (O_79,N_2762,N_2965);
nor UO_80 (O_80,N_2448,N_2837);
and UO_81 (O_81,N_2798,N_2816);
and UO_82 (O_82,N_2649,N_2472);
nor UO_83 (O_83,N_2881,N_2863);
nand UO_84 (O_84,N_2931,N_2479);
nor UO_85 (O_85,N_2493,N_2899);
xor UO_86 (O_86,N_2544,N_2942);
or UO_87 (O_87,N_2543,N_2595);
or UO_88 (O_88,N_2977,N_2830);
xnor UO_89 (O_89,N_2530,N_2932);
or UO_90 (O_90,N_2489,N_2553);
or UO_91 (O_91,N_2414,N_2782);
nand UO_92 (O_92,N_2927,N_2650);
nand UO_93 (O_93,N_2908,N_2766);
xnor UO_94 (O_94,N_2819,N_2875);
nor UO_95 (O_95,N_2551,N_2500);
nand UO_96 (O_96,N_2470,N_2773);
nand UO_97 (O_97,N_2909,N_2890);
nand UO_98 (O_98,N_2739,N_2736);
nand UO_99 (O_99,N_2685,N_2610);
and UO_100 (O_100,N_2843,N_2902);
nand UO_101 (O_101,N_2690,N_2868);
and UO_102 (O_102,N_2765,N_2725);
or UO_103 (O_103,N_2545,N_2905);
nor UO_104 (O_104,N_2410,N_2794);
nand UO_105 (O_105,N_2617,N_2491);
nand UO_106 (O_106,N_2813,N_2987);
and UO_107 (O_107,N_2417,N_2593);
or UO_108 (O_108,N_2581,N_2950);
nor UO_109 (O_109,N_2403,N_2779);
nor UO_110 (O_110,N_2806,N_2515);
nor UO_111 (O_111,N_2720,N_2566);
and UO_112 (O_112,N_2548,N_2800);
and UO_113 (O_113,N_2946,N_2713);
or UO_114 (O_114,N_2579,N_2990);
and UO_115 (O_115,N_2538,N_2856);
and UO_116 (O_116,N_2712,N_2892);
nor UO_117 (O_117,N_2777,N_2785);
or UO_118 (O_118,N_2808,N_2850);
or UO_119 (O_119,N_2746,N_2475);
or UO_120 (O_120,N_2797,N_2628);
nand UO_121 (O_121,N_2625,N_2876);
and UO_122 (O_122,N_2877,N_2768);
nor UO_123 (O_123,N_2464,N_2846);
nand UO_124 (O_124,N_2433,N_2833);
xnor UO_125 (O_125,N_2462,N_2913);
nor UO_126 (O_126,N_2858,N_2844);
nand UO_127 (O_127,N_2659,N_2729);
nor UO_128 (O_128,N_2558,N_2460);
or UO_129 (O_129,N_2436,N_2906);
or UO_130 (O_130,N_2636,N_2666);
and UO_131 (O_131,N_2634,N_2517);
nand UO_132 (O_132,N_2971,N_2943);
nand UO_133 (O_133,N_2870,N_2439);
and UO_134 (O_134,N_2632,N_2698);
nor UO_135 (O_135,N_2562,N_2734);
and UO_136 (O_136,N_2635,N_2847);
nor UO_137 (O_137,N_2519,N_2526);
or UO_138 (O_138,N_2496,N_2702);
nand UO_139 (O_139,N_2638,N_2409);
and UO_140 (O_140,N_2976,N_2671);
and UO_141 (O_141,N_2730,N_2539);
nor UO_142 (O_142,N_2880,N_2535);
or UO_143 (O_143,N_2928,N_2576);
nor UO_144 (O_144,N_2559,N_2582);
or UO_145 (O_145,N_2665,N_2752);
nor UO_146 (O_146,N_2474,N_2572);
xor UO_147 (O_147,N_2944,N_2874);
and UO_148 (O_148,N_2726,N_2705);
or UO_149 (O_149,N_2771,N_2402);
nor UO_150 (O_150,N_2699,N_2440);
nand UO_151 (O_151,N_2731,N_2481);
nor UO_152 (O_152,N_2669,N_2453);
or UO_153 (O_153,N_2564,N_2829);
or UO_154 (O_154,N_2505,N_2585);
nor UO_155 (O_155,N_2714,N_2933);
nor UO_156 (O_156,N_2855,N_2516);
nand UO_157 (O_157,N_2471,N_2533);
or UO_158 (O_158,N_2925,N_2804);
and UO_159 (O_159,N_2577,N_2434);
and UO_160 (O_160,N_2939,N_2678);
nor UO_161 (O_161,N_2988,N_2801);
nor UO_162 (O_162,N_2921,N_2821);
nand UO_163 (O_163,N_2936,N_2701);
nor UO_164 (O_164,N_2422,N_2822);
or UO_165 (O_165,N_2688,N_2560);
nand UO_166 (O_166,N_2461,N_2442);
and UO_167 (O_167,N_2614,N_2631);
or UO_168 (O_168,N_2525,N_2465);
nor UO_169 (O_169,N_2476,N_2900);
nor UO_170 (O_170,N_2477,N_2981);
and UO_171 (O_171,N_2660,N_2784);
nor UO_172 (O_172,N_2783,N_2613);
and UO_173 (O_173,N_2588,N_2737);
and UO_174 (O_174,N_2865,N_2512);
or UO_175 (O_175,N_2605,N_2415);
and UO_176 (O_176,N_2549,N_2486);
or UO_177 (O_177,N_2643,N_2416);
or UO_178 (O_178,N_2718,N_2567);
xnor UO_179 (O_179,N_2859,N_2668);
and UO_180 (O_180,N_2772,N_2692);
and UO_181 (O_181,N_2842,N_2923);
or UO_182 (O_182,N_2751,N_2497);
and UO_183 (O_183,N_2642,N_2445);
nand UO_184 (O_184,N_2825,N_2894);
nor UO_185 (O_185,N_2991,N_2732);
or UO_186 (O_186,N_2604,N_2446);
or UO_187 (O_187,N_2599,N_2652);
nor UO_188 (O_188,N_2926,N_2583);
and UO_189 (O_189,N_2524,N_2840);
nand UO_190 (O_190,N_2589,N_2428);
or UO_191 (O_191,N_2503,N_2407);
and UO_192 (O_192,N_2607,N_2911);
and UO_193 (O_193,N_2873,N_2618);
or UO_194 (O_194,N_2429,N_2487);
nor UO_195 (O_195,N_2978,N_2694);
nor UO_196 (O_196,N_2621,N_2606);
and UO_197 (O_197,N_2807,N_2639);
nand UO_198 (O_198,N_2903,N_2895);
or UO_199 (O_199,N_2918,N_2826);
and UO_200 (O_200,N_2802,N_2484);
xnor UO_201 (O_201,N_2506,N_2574);
nor UO_202 (O_202,N_2696,N_2889);
nand UO_203 (O_203,N_2787,N_2419);
or UO_204 (O_204,N_2757,N_2841);
and UO_205 (O_205,N_2679,N_2400);
xnor UO_206 (O_206,N_2444,N_2716);
or UO_207 (O_207,N_2832,N_2767);
and UO_208 (O_208,N_2629,N_2653);
nor UO_209 (O_209,N_2680,N_2924);
nor UO_210 (O_210,N_2790,N_2466);
nor UO_211 (O_211,N_2597,N_2828);
or UO_212 (O_212,N_2957,N_2619);
or UO_213 (O_213,N_2449,N_2514);
nand UO_214 (O_214,N_2857,N_2437);
and UO_215 (O_215,N_2707,N_2507);
and UO_216 (O_216,N_2945,N_2427);
nor UO_217 (O_217,N_2778,N_2891);
or UO_218 (O_218,N_2681,N_2616);
xor UO_219 (O_219,N_2912,N_2759);
nand UO_220 (O_220,N_2845,N_2473);
or UO_221 (O_221,N_2986,N_2522);
or UO_222 (O_222,N_2975,N_2934);
or UO_223 (O_223,N_2789,N_2520);
or UO_224 (O_224,N_2684,N_2852);
xor UO_225 (O_225,N_2964,N_2527);
nand UO_226 (O_226,N_2992,N_2776);
nand UO_227 (O_227,N_2963,N_2910);
xor UO_228 (O_228,N_2743,N_2882);
nor UO_229 (O_229,N_2412,N_2883);
and UO_230 (O_230,N_2715,N_2770);
or UO_231 (O_231,N_2862,N_2623);
nor UO_232 (O_232,N_2866,N_2630);
nand UO_233 (O_233,N_2995,N_2513);
or UO_234 (O_234,N_2967,N_2755);
nand UO_235 (O_235,N_2683,N_2792);
or UO_236 (O_236,N_2423,N_2663);
or UO_237 (O_237,N_2849,N_2498);
and UO_238 (O_238,N_2624,N_2569);
and UO_239 (O_239,N_2838,N_2570);
nor UO_240 (O_240,N_2989,N_2754);
nand UO_241 (O_241,N_2915,N_2886);
and UO_242 (O_242,N_2727,N_2615);
or UO_243 (O_243,N_2578,N_2483);
and UO_244 (O_244,N_2710,N_2997);
nand UO_245 (O_245,N_2879,N_2557);
nor UO_246 (O_246,N_2480,N_2686);
nand UO_247 (O_247,N_2555,N_2867);
and UO_248 (O_248,N_2741,N_2482);
xor UO_249 (O_249,N_2662,N_2468);
nand UO_250 (O_250,N_2675,N_2824);
nand UO_251 (O_251,N_2791,N_2457);
xnor UO_252 (O_252,N_2728,N_2756);
nor UO_253 (O_253,N_2531,N_2528);
or UO_254 (O_254,N_2878,N_2590);
nor UO_255 (O_255,N_2796,N_2573);
nand UO_256 (O_256,N_2920,N_2953);
and UO_257 (O_257,N_2704,N_2775);
nand UO_258 (O_258,N_2961,N_2769);
or UO_259 (O_259,N_2405,N_2523);
or UO_260 (O_260,N_2586,N_2996);
or UO_261 (O_261,N_2723,N_2854);
nand UO_262 (O_262,N_2919,N_2955);
and UO_263 (O_263,N_2408,N_2968);
nand UO_264 (O_264,N_2456,N_2706);
or UO_265 (O_265,N_2521,N_2851);
xnor UO_266 (O_266,N_2904,N_2722);
or UO_267 (O_267,N_2985,N_2951);
nor UO_268 (O_268,N_2661,N_2565);
and UO_269 (O_269,N_2646,N_2753);
and UO_270 (O_270,N_2812,N_2563);
nor UO_271 (O_271,N_2805,N_2914);
and UO_272 (O_272,N_2492,N_2693);
nor UO_273 (O_273,N_2431,N_2917);
and UO_274 (O_274,N_2721,N_2960);
nor UO_275 (O_275,N_2580,N_2600);
and UO_276 (O_276,N_2571,N_2839);
and UO_277 (O_277,N_2450,N_2541);
or UO_278 (O_278,N_2745,N_2860);
nand UO_279 (O_279,N_2717,N_2536);
nor UO_280 (O_280,N_2592,N_2962);
nand UO_281 (O_281,N_2540,N_2747);
and UO_282 (O_282,N_2836,N_2501);
or UO_283 (O_283,N_2817,N_2815);
and UO_284 (O_284,N_2983,N_2664);
and UO_285 (O_285,N_2441,N_2949);
nand UO_286 (O_286,N_2922,N_2947);
nand UO_287 (O_287,N_2508,N_2761);
or UO_288 (O_288,N_2853,N_2529);
and UO_289 (O_289,N_2708,N_2406);
and UO_290 (O_290,N_2689,N_2764);
and UO_291 (O_291,N_2818,N_2941);
and UO_292 (O_292,N_2598,N_2740);
and UO_293 (O_293,N_2459,N_2622);
xnor UO_294 (O_294,N_2499,N_2982);
nor UO_295 (O_295,N_2724,N_2979);
nor UO_296 (O_296,N_2998,N_2438);
xnor UO_297 (O_297,N_2452,N_2887);
or UO_298 (O_298,N_2667,N_2670);
nor UO_299 (O_299,N_2591,N_2980);
nand UO_300 (O_300,N_2971,N_2691);
or UO_301 (O_301,N_2599,N_2966);
or UO_302 (O_302,N_2473,N_2905);
xnor UO_303 (O_303,N_2966,N_2784);
and UO_304 (O_304,N_2810,N_2710);
or UO_305 (O_305,N_2995,N_2675);
or UO_306 (O_306,N_2490,N_2826);
nand UO_307 (O_307,N_2424,N_2553);
nor UO_308 (O_308,N_2595,N_2520);
nand UO_309 (O_309,N_2490,N_2999);
and UO_310 (O_310,N_2790,N_2941);
nor UO_311 (O_311,N_2803,N_2740);
or UO_312 (O_312,N_2826,N_2467);
xor UO_313 (O_313,N_2556,N_2617);
nor UO_314 (O_314,N_2721,N_2805);
nor UO_315 (O_315,N_2906,N_2713);
or UO_316 (O_316,N_2847,N_2631);
or UO_317 (O_317,N_2767,N_2797);
nor UO_318 (O_318,N_2856,N_2631);
nand UO_319 (O_319,N_2920,N_2649);
nor UO_320 (O_320,N_2924,N_2782);
nor UO_321 (O_321,N_2799,N_2615);
and UO_322 (O_322,N_2744,N_2767);
or UO_323 (O_323,N_2557,N_2977);
nand UO_324 (O_324,N_2651,N_2940);
nand UO_325 (O_325,N_2785,N_2790);
and UO_326 (O_326,N_2419,N_2464);
and UO_327 (O_327,N_2918,N_2784);
xnor UO_328 (O_328,N_2987,N_2870);
or UO_329 (O_329,N_2658,N_2576);
or UO_330 (O_330,N_2812,N_2757);
nand UO_331 (O_331,N_2465,N_2607);
or UO_332 (O_332,N_2950,N_2873);
xnor UO_333 (O_333,N_2944,N_2533);
nand UO_334 (O_334,N_2438,N_2792);
nand UO_335 (O_335,N_2501,N_2977);
xor UO_336 (O_336,N_2654,N_2800);
nor UO_337 (O_337,N_2749,N_2935);
or UO_338 (O_338,N_2703,N_2807);
or UO_339 (O_339,N_2708,N_2938);
or UO_340 (O_340,N_2577,N_2918);
or UO_341 (O_341,N_2474,N_2984);
nand UO_342 (O_342,N_2484,N_2700);
or UO_343 (O_343,N_2471,N_2832);
nand UO_344 (O_344,N_2781,N_2984);
nor UO_345 (O_345,N_2440,N_2612);
and UO_346 (O_346,N_2643,N_2743);
and UO_347 (O_347,N_2873,N_2766);
or UO_348 (O_348,N_2778,N_2931);
xnor UO_349 (O_349,N_2752,N_2834);
xnor UO_350 (O_350,N_2822,N_2525);
nand UO_351 (O_351,N_2543,N_2949);
nor UO_352 (O_352,N_2984,N_2581);
nand UO_353 (O_353,N_2907,N_2869);
or UO_354 (O_354,N_2905,N_2980);
and UO_355 (O_355,N_2609,N_2574);
and UO_356 (O_356,N_2817,N_2967);
or UO_357 (O_357,N_2501,N_2443);
or UO_358 (O_358,N_2963,N_2969);
nand UO_359 (O_359,N_2608,N_2864);
nand UO_360 (O_360,N_2505,N_2588);
or UO_361 (O_361,N_2766,N_2797);
nor UO_362 (O_362,N_2703,N_2821);
nor UO_363 (O_363,N_2405,N_2563);
xnor UO_364 (O_364,N_2512,N_2893);
nand UO_365 (O_365,N_2762,N_2684);
and UO_366 (O_366,N_2563,N_2986);
xor UO_367 (O_367,N_2678,N_2473);
nand UO_368 (O_368,N_2569,N_2938);
nand UO_369 (O_369,N_2787,N_2576);
nand UO_370 (O_370,N_2608,N_2889);
or UO_371 (O_371,N_2792,N_2670);
or UO_372 (O_372,N_2469,N_2796);
or UO_373 (O_373,N_2578,N_2627);
and UO_374 (O_374,N_2506,N_2561);
nand UO_375 (O_375,N_2466,N_2783);
or UO_376 (O_376,N_2536,N_2501);
nand UO_377 (O_377,N_2579,N_2552);
xnor UO_378 (O_378,N_2637,N_2920);
or UO_379 (O_379,N_2402,N_2731);
xnor UO_380 (O_380,N_2999,N_2876);
nor UO_381 (O_381,N_2454,N_2696);
or UO_382 (O_382,N_2832,N_2535);
or UO_383 (O_383,N_2848,N_2990);
nor UO_384 (O_384,N_2420,N_2409);
and UO_385 (O_385,N_2646,N_2610);
nand UO_386 (O_386,N_2743,N_2695);
nor UO_387 (O_387,N_2442,N_2922);
nor UO_388 (O_388,N_2885,N_2510);
and UO_389 (O_389,N_2911,N_2771);
and UO_390 (O_390,N_2826,N_2564);
and UO_391 (O_391,N_2996,N_2955);
or UO_392 (O_392,N_2494,N_2988);
nand UO_393 (O_393,N_2423,N_2415);
and UO_394 (O_394,N_2465,N_2796);
nor UO_395 (O_395,N_2726,N_2648);
nor UO_396 (O_396,N_2910,N_2873);
nand UO_397 (O_397,N_2859,N_2755);
nand UO_398 (O_398,N_2428,N_2585);
nor UO_399 (O_399,N_2869,N_2839);
xnor UO_400 (O_400,N_2711,N_2471);
nor UO_401 (O_401,N_2471,N_2503);
xnor UO_402 (O_402,N_2940,N_2910);
nor UO_403 (O_403,N_2455,N_2987);
nor UO_404 (O_404,N_2721,N_2817);
nor UO_405 (O_405,N_2974,N_2574);
or UO_406 (O_406,N_2679,N_2593);
nor UO_407 (O_407,N_2552,N_2692);
xnor UO_408 (O_408,N_2735,N_2723);
and UO_409 (O_409,N_2462,N_2513);
nand UO_410 (O_410,N_2472,N_2929);
xor UO_411 (O_411,N_2963,N_2973);
and UO_412 (O_412,N_2699,N_2580);
and UO_413 (O_413,N_2545,N_2403);
nor UO_414 (O_414,N_2554,N_2810);
and UO_415 (O_415,N_2572,N_2555);
nand UO_416 (O_416,N_2926,N_2952);
or UO_417 (O_417,N_2489,N_2782);
nor UO_418 (O_418,N_2501,N_2682);
or UO_419 (O_419,N_2680,N_2934);
nor UO_420 (O_420,N_2971,N_2829);
and UO_421 (O_421,N_2923,N_2461);
or UO_422 (O_422,N_2830,N_2786);
or UO_423 (O_423,N_2783,N_2843);
and UO_424 (O_424,N_2555,N_2793);
or UO_425 (O_425,N_2839,N_2622);
and UO_426 (O_426,N_2965,N_2719);
or UO_427 (O_427,N_2787,N_2454);
nand UO_428 (O_428,N_2410,N_2574);
nor UO_429 (O_429,N_2955,N_2734);
nor UO_430 (O_430,N_2668,N_2734);
or UO_431 (O_431,N_2570,N_2869);
nand UO_432 (O_432,N_2668,N_2611);
nor UO_433 (O_433,N_2988,N_2549);
or UO_434 (O_434,N_2735,N_2831);
or UO_435 (O_435,N_2639,N_2426);
or UO_436 (O_436,N_2819,N_2987);
xnor UO_437 (O_437,N_2914,N_2869);
nor UO_438 (O_438,N_2963,N_2991);
xor UO_439 (O_439,N_2797,N_2989);
xor UO_440 (O_440,N_2520,N_2824);
xnor UO_441 (O_441,N_2551,N_2567);
nor UO_442 (O_442,N_2622,N_2868);
or UO_443 (O_443,N_2759,N_2677);
nand UO_444 (O_444,N_2907,N_2586);
and UO_445 (O_445,N_2815,N_2515);
nor UO_446 (O_446,N_2623,N_2915);
nand UO_447 (O_447,N_2925,N_2969);
nand UO_448 (O_448,N_2750,N_2793);
and UO_449 (O_449,N_2553,N_2504);
nor UO_450 (O_450,N_2793,N_2538);
and UO_451 (O_451,N_2614,N_2906);
nand UO_452 (O_452,N_2957,N_2772);
nand UO_453 (O_453,N_2875,N_2954);
or UO_454 (O_454,N_2861,N_2902);
or UO_455 (O_455,N_2562,N_2666);
nand UO_456 (O_456,N_2954,N_2787);
nor UO_457 (O_457,N_2408,N_2912);
and UO_458 (O_458,N_2459,N_2669);
nand UO_459 (O_459,N_2447,N_2893);
and UO_460 (O_460,N_2968,N_2489);
or UO_461 (O_461,N_2773,N_2493);
nor UO_462 (O_462,N_2553,N_2636);
nand UO_463 (O_463,N_2869,N_2806);
nor UO_464 (O_464,N_2406,N_2911);
and UO_465 (O_465,N_2779,N_2722);
or UO_466 (O_466,N_2973,N_2421);
nand UO_467 (O_467,N_2823,N_2879);
nor UO_468 (O_468,N_2882,N_2533);
and UO_469 (O_469,N_2931,N_2932);
and UO_470 (O_470,N_2610,N_2535);
nand UO_471 (O_471,N_2863,N_2448);
or UO_472 (O_472,N_2807,N_2618);
nor UO_473 (O_473,N_2405,N_2740);
nor UO_474 (O_474,N_2738,N_2915);
nand UO_475 (O_475,N_2542,N_2482);
nor UO_476 (O_476,N_2475,N_2405);
nand UO_477 (O_477,N_2488,N_2712);
or UO_478 (O_478,N_2696,N_2679);
nand UO_479 (O_479,N_2809,N_2564);
and UO_480 (O_480,N_2457,N_2746);
xnor UO_481 (O_481,N_2654,N_2726);
or UO_482 (O_482,N_2837,N_2455);
nor UO_483 (O_483,N_2477,N_2478);
and UO_484 (O_484,N_2434,N_2745);
or UO_485 (O_485,N_2737,N_2591);
xor UO_486 (O_486,N_2570,N_2606);
nor UO_487 (O_487,N_2808,N_2804);
and UO_488 (O_488,N_2740,N_2678);
nand UO_489 (O_489,N_2925,N_2927);
nor UO_490 (O_490,N_2943,N_2582);
and UO_491 (O_491,N_2692,N_2865);
nand UO_492 (O_492,N_2809,N_2630);
xnor UO_493 (O_493,N_2973,N_2890);
and UO_494 (O_494,N_2464,N_2762);
nor UO_495 (O_495,N_2690,N_2911);
nor UO_496 (O_496,N_2511,N_2433);
and UO_497 (O_497,N_2610,N_2575);
or UO_498 (O_498,N_2494,N_2713);
nand UO_499 (O_499,N_2706,N_2972);
endmodule