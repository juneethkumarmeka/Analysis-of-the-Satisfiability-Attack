module basic_500_3000_500_60_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_303,In_435);
or U1 (N_1,In_344,In_149);
and U2 (N_2,In_23,In_385);
nand U3 (N_3,In_295,In_419);
or U4 (N_4,In_146,In_114);
nand U5 (N_5,In_299,In_498);
nor U6 (N_6,In_212,In_313);
nand U7 (N_7,In_264,In_266);
and U8 (N_8,In_221,In_242);
or U9 (N_9,In_357,In_274);
nor U10 (N_10,In_230,In_423);
or U11 (N_11,In_410,In_120);
nand U12 (N_12,In_27,In_191);
nor U13 (N_13,In_144,In_99);
nand U14 (N_14,In_178,In_20);
nand U15 (N_15,In_224,In_424);
and U16 (N_16,In_436,In_170);
or U17 (N_17,In_129,In_259);
nand U18 (N_18,In_91,In_452);
and U19 (N_19,In_281,In_46);
and U20 (N_20,In_422,In_387);
nand U21 (N_21,In_258,In_217);
nor U22 (N_22,In_347,In_163);
or U23 (N_23,In_416,In_108);
or U24 (N_24,In_225,In_94);
xor U25 (N_25,In_199,In_67);
or U26 (N_26,In_362,In_493);
nor U27 (N_27,In_378,In_147);
and U28 (N_28,In_336,In_138);
nor U29 (N_29,In_280,In_492);
and U30 (N_30,In_255,In_375);
or U31 (N_31,In_234,In_126);
and U32 (N_32,In_162,In_449);
nor U33 (N_33,In_480,In_263);
or U34 (N_34,In_155,In_366);
xnor U35 (N_35,In_222,In_239);
and U36 (N_36,In_157,In_428);
or U37 (N_37,In_211,In_327);
or U38 (N_38,In_245,In_437);
nand U39 (N_39,In_92,In_297);
or U40 (N_40,In_17,In_343);
nand U41 (N_41,In_409,In_18);
and U42 (N_42,In_55,In_139);
nand U43 (N_43,In_88,In_481);
and U44 (N_44,In_68,In_451);
nand U45 (N_45,In_30,In_250);
nand U46 (N_46,In_175,In_107);
or U47 (N_47,In_220,In_432);
nor U48 (N_48,In_499,In_391);
nor U49 (N_49,In_190,In_286);
nor U50 (N_50,In_329,In_197);
and U51 (N_51,In_478,In_156);
nand U52 (N_52,In_397,In_322);
nand U53 (N_53,In_270,In_124);
or U54 (N_54,In_355,N_5);
nor U55 (N_55,In_66,In_81);
and U56 (N_56,In_62,In_232);
or U57 (N_57,N_49,In_41);
nand U58 (N_58,In_458,In_292);
nor U59 (N_59,In_354,In_373);
nand U60 (N_60,In_381,In_341);
nor U61 (N_61,In_213,In_383);
and U62 (N_62,In_348,N_3);
or U63 (N_63,In_202,In_179);
nor U64 (N_64,In_145,In_188);
nor U65 (N_65,In_434,In_330);
nand U66 (N_66,In_164,In_122);
nor U67 (N_67,In_102,In_168);
and U68 (N_68,In_491,In_421);
nand U69 (N_69,In_128,In_87);
nor U70 (N_70,In_117,N_39);
or U71 (N_71,N_41,In_85);
and U72 (N_72,In_314,In_9);
and U73 (N_73,In_448,In_417);
nand U74 (N_74,In_334,In_187);
or U75 (N_75,In_365,In_60);
or U76 (N_76,In_185,In_171);
and U77 (N_77,In_294,In_352);
nor U78 (N_78,In_69,In_45);
and U79 (N_79,In_226,In_489);
nor U80 (N_80,In_33,In_119);
and U81 (N_81,In_214,In_218);
or U82 (N_82,In_2,In_390);
nand U83 (N_83,In_254,In_184);
nor U84 (N_84,In_4,In_453);
nor U85 (N_85,N_15,In_261);
and U86 (N_86,In_360,In_291);
xnor U87 (N_87,In_488,In_337);
and U88 (N_88,In_172,In_283);
and U89 (N_89,In_29,In_364);
nor U90 (N_90,In_43,In_363);
or U91 (N_91,In_472,N_24);
nor U92 (N_92,In_31,In_111);
xor U93 (N_93,In_65,In_406);
nor U94 (N_94,In_186,In_192);
xor U95 (N_95,In_229,In_160);
nor U96 (N_96,In_350,In_228);
and U97 (N_97,In_326,In_466);
nor U98 (N_98,In_77,In_426);
and U99 (N_99,In_133,In_316);
or U100 (N_100,N_77,N_44);
or U101 (N_101,N_95,In_444);
nand U102 (N_102,In_7,In_84);
nor U103 (N_103,In_93,In_310);
or U104 (N_104,In_482,In_265);
and U105 (N_105,In_32,In_318);
nor U106 (N_106,In_39,In_16);
and U107 (N_107,N_21,N_75);
or U108 (N_108,In_96,N_94);
or U109 (N_109,In_408,In_253);
nor U110 (N_110,In_269,In_47);
or U111 (N_111,N_14,In_433);
and U112 (N_112,In_233,In_332);
and U113 (N_113,In_331,In_44);
and U114 (N_114,In_300,In_462);
nor U115 (N_115,In_181,In_14);
nor U116 (N_116,N_88,In_219);
nor U117 (N_117,In_112,N_60);
nand U118 (N_118,In_298,N_51);
nor U119 (N_119,In_97,In_396);
and U120 (N_120,In_34,N_22);
and U121 (N_121,N_33,In_1);
nor U122 (N_122,In_374,In_143);
nor U123 (N_123,In_152,In_306);
or U124 (N_124,In_57,In_401);
or U125 (N_125,In_389,In_319);
and U126 (N_126,N_48,N_54);
nand U127 (N_127,In_438,In_210);
or U128 (N_128,In_456,In_338);
nand U129 (N_129,N_9,N_43);
and U130 (N_130,In_174,In_372);
xnor U131 (N_131,In_321,In_340);
nand U132 (N_132,In_324,In_285);
nor U133 (N_133,In_59,N_7);
nand U134 (N_134,N_74,In_35);
nand U135 (N_135,In_400,N_46);
or U136 (N_136,In_257,In_247);
or U137 (N_137,In_86,In_246);
nand U138 (N_138,N_89,In_182);
nand U139 (N_139,In_459,N_73);
and U140 (N_140,In_414,In_19);
nand U141 (N_141,In_279,In_477);
or U142 (N_142,In_442,In_72);
nor U143 (N_143,N_11,In_439);
nor U144 (N_144,In_369,In_209);
nand U145 (N_145,In_325,In_474);
nor U146 (N_146,In_0,In_305);
nor U147 (N_147,N_28,In_398);
nor U148 (N_148,In_130,In_113);
or U149 (N_149,N_42,In_388);
and U150 (N_150,N_56,N_32);
or U151 (N_151,In_6,N_4);
nor U152 (N_152,In_427,N_31);
and U153 (N_153,N_66,In_167);
nor U154 (N_154,In_312,In_443);
and U155 (N_155,In_148,N_124);
and U156 (N_156,N_53,N_90);
and U157 (N_157,N_142,In_301);
or U158 (N_158,In_345,In_116);
or U159 (N_159,N_81,In_193);
and U160 (N_160,In_278,In_356);
nor U161 (N_161,In_158,In_431);
or U162 (N_162,N_133,N_109);
nor U163 (N_163,N_85,In_37);
nand U164 (N_164,In_260,N_122);
and U165 (N_165,In_207,In_403);
nor U166 (N_166,In_275,In_430);
or U167 (N_167,In_342,In_73);
and U168 (N_168,In_105,N_16);
nor U169 (N_169,N_13,In_351);
nand U170 (N_170,In_25,In_415);
nor U171 (N_171,In_201,In_249);
nor U172 (N_172,In_244,N_68);
nor U173 (N_173,In_71,N_40);
nand U174 (N_174,In_315,In_287);
and U175 (N_175,In_317,In_471);
and U176 (N_176,N_107,N_72);
or U177 (N_177,In_237,In_289);
or U178 (N_178,In_495,N_116);
and U179 (N_179,In_36,In_479);
or U180 (N_180,N_62,N_135);
nand U181 (N_181,In_311,In_455);
nand U182 (N_182,In_240,In_150);
nand U183 (N_183,N_104,In_216);
or U184 (N_184,In_349,N_121);
and U185 (N_185,In_418,In_272);
nor U186 (N_186,In_26,N_82);
or U187 (N_187,In_70,N_125);
nand U188 (N_188,In_40,In_204);
nor U189 (N_189,In_195,N_141);
nor U190 (N_190,In_79,N_36);
nor U191 (N_191,N_118,In_487);
nand U192 (N_192,N_110,N_128);
and U193 (N_193,In_49,In_282);
nand U194 (N_194,N_8,In_243);
nor U195 (N_195,In_177,N_138);
nor U196 (N_196,N_97,N_80);
nor U197 (N_197,In_132,In_441);
and U198 (N_198,In_486,In_323);
or U199 (N_199,N_145,In_166);
nand U200 (N_200,N_103,N_57);
and U201 (N_201,N_158,In_159);
nor U202 (N_202,In_328,N_139);
and U203 (N_203,In_238,In_196);
and U204 (N_204,N_137,N_86);
nor U205 (N_205,N_112,In_288);
nor U206 (N_206,N_63,In_11);
nor U207 (N_207,In_395,In_53);
and U208 (N_208,N_114,In_123);
xor U209 (N_209,N_161,In_52);
nand U210 (N_210,In_135,N_98);
nand U211 (N_211,N_69,N_19);
or U212 (N_212,N_65,N_61);
nand U213 (N_213,In_5,In_429);
or U214 (N_214,N_195,N_123);
nor U215 (N_215,N_134,N_76);
nand U216 (N_216,N_34,N_197);
nand U217 (N_217,In_110,In_180);
nand U218 (N_218,In_63,N_192);
and U219 (N_219,N_152,In_484);
or U220 (N_220,In_194,In_256);
or U221 (N_221,N_83,N_185);
nor U222 (N_222,N_164,In_154);
nor U223 (N_223,In_8,In_464);
and U224 (N_224,N_119,In_42);
nand U225 (N_225,N_59,N_143);
or U226 (N_226,N_25,In_377);
nor U227 (N_227,In_267,N_55);
and U228 (N_228,In_203,In_339);
nor U229 (N_229,N_27,N_10);
xnor U230 (N_230,In_425,N_193);
and U231 (N_231,In_125,N_126);
nand U232 (N_232,N_157,In_273);
and U233 (N_233,In_165,In_22);
or U234 (N_234,N_198,In_335);
and U235 (N_235,In_473,N_160);
nor U236 (N_236,N_189,N_102);
nand U237 (N_237,In_227,In_76);
or U238 (N_238,In_208,In_371);
nand U239 (N_239,N_18,In_284);
nor U240 (N_240,N_99,N_93);
and U241 (N_241,In_21,In_136);
nand U242 (N_242,In_460,In_15);
nor U243 (N_243,In_64,In_56);
nor U244 (N_244,In_386,N_180);
and U245 (N_245,In_320,N_131);
nand U246 (N_246,In_54,In_333);
nor U247 (N_247,In_346,In_109);
nor U248 (N_248,N_174,In_361);
nor U249 (N_249,In_142,N_58);
nand U250 (N_250,In_153,N_222);
nand U251 (N_251,N_196,In_137);
and U252 (N_252,In_307,In_12);
or U253 (N_253,In_141,In_470);
nor U254 (N_254,In_309,In_497);
nor U255 (N_255,N_239,In_118);
or U256 (N_256,In_413,N_0);
nor U257 (N_257,N_212,In_370);
nor U258 (N_258,N_163,In_98);
and U259 (N_259,In_74,N_204);
nand U260 (N_260,N_190,In_83);
or U261 (N_261,In_205,In_293);
or U262 (N_262,In_106,N_183);
or U263 (N_263,N_223,In_476);
nor U264 (N_264,N_227,In_151);
or U265 (N_265,N_2,N_225);
nand U266 (N_266,N_153,N_35);
and U267 (N_267,N_181,N_228);
or U268 (N_268,In_475,In_95);
or U269 (N_269,N_247,N_168);
nor U270 (N_270,N_167,N_246);
nor U271 (N_271,In_103,In_276);
nor U272 (N_272,N_232,N_224);
or U273 (N_273,N_177,N_87);
and U274 (N_274,N_146,N_249);
or U275 (N_275,N_84,In_277);
or U276 (N_276,N_26,N_182);
and U277 (N_277,N_67,N_231);
nor U278 (N_278,N_179,In_48);
nand U279 (N_279,N_6,In_50);
nand U280 (N_280,In_367,In_446);
nand U281 (N_281,N_23,N_241);
nand U282 (N_282,N_113,In_236);
nand U283 (N_283,In_420,In_394);
nor U284 (N_284,In_121,In_393);
nor U285 (N_285,N_100,In_235);
nor U286 (N_286,N_150,In_304);
nand U287 (N_287,In_379,In_176);
nand U288 (N_288,N_170,In_490);
nor U289 (N_289,In_252,N_71);
nand U290 (N_290,In_271,N_237);
or U291 (N_291,N_218,In_463);
xnor U292 (N_292,N_208,In_198);
nor U293 (N_293,In_101,N_199);
nor U294 (N_294,N_203,In_461);
or U295 (N_295,In_100,N_171);
or U296 (N_296,In_469,N_120);
nand U297 (N_297,N_205,N_155);
and U298 (N_298,In_468,In_173);
nor U299 (N_299,N_129,In_61);
nand U300 (N_300,In_104,N_215);
nor U301 (N_301,N_288,N_37);
or U302 (N_302,N_281,N_149);
or U303 (N_303,N_295,N_176);
or U304 (N_304,In_28,N_202);
nand U305 (N_305,N_240,N_299);
and U306 (N_306,In_440,N_30);
nand U307 (N_307,N_220,In_496);
or U308 (N_308,N_130,N_284);
nor U309 (N_309,N_173,N_186);
nand U310 (N_310,In_404,N_271);
and U311 (N_311,In_302,N_217);
nand U312 (N_312,N_259,N_156);
nor U313 (N_313,In_206,N_206);
nand U314 (N_314,In_231,In_445);
or U315 (N_315,N_233,N_254);
nor U316 (N_316,N_159,In_13);
xor U317 (N_317,N_132,In_411);
or U318 (N_318,N_266,N_296);
nor U319 (N_319,In_454,N_96);
nor U320 (N_320,N_144,N_274);
or U321 (N_321,N_243,N_229);
or U322 (N_322,In_447,N_270);
or U323 (N_323,N_207,N_263);
and U324 (N_324,N_108,N_275);
or U325 (N_325,In_78,In_75);
nand U326 (N_326,N_166,N_209);
or U327 (N_327,In_353,N_50);
nor U328 (N_328,In_358,In_382);
or U329 (N_329,N_261,N_175);
nor U330 (N_330,N_105,N_169);
or U331 (N_331,In_376,N_238);
nor U332 (N_332,N_127,N_47);
nand U333 (N_333,In_89,N_283);
or U334 (N_334,In_115,N_214);
and U335 (N_335,N_267,N_286);
nand U336 (N_336,N_244,N_255);
and U337 (N_337,N_101,N_252);
nand U338 (N_338,N_273,N_1);
nor U339 (N_339,N_264,N_234);
or U340 (N_340,N_194,N_178);
nor U341 (N_341,In_457,N_70);
nand U342 (N_342,In_380,N_64);
and U343 (N_343,In_223,In_467);
xnor U344 (N_344,N_235,N_290);
or U345 (N_345,In_465,N_148);
or U346 (N_346,N_52,In_368);
and U347 (N_347,N_293,N_91);
or U348 (N_348,In_392,N_269);
nand U349 (N_349,In_134,In_24);
nor U350 (N_350,N_311,N_282);
or U351 (N_351,N_337,N_294);
nand U352 (N_352,N_279,In_131);
nand U353 (N_353,N_260,N_184);
or U354 (N_354,N_313,N_219);
or U355 (N_355,N_291,N_257);
or U356 (N_356,N_278,N_314);
nor U357 (N_357,In_268,N_298);
and U358 (N_358,N_346,N_265);
and U359 (N_359,N_251,N_276);
nor U360 (N_360,In_90,In_200);
or U361 (N_361,N_304,N_335);
and U362 (N_362,N_322,N_210);
and U363 (N_363,N_336,In_359);
nand U364 (N_364,In_215,N_285);
nand U365 (N_365,N_330,N_200);
nor U366 (N_366,N_253,N_349);
or U367 (N_367,N_318,N_277);
or U368 (N_368,N_309,N_348);
nor U369 (N_369,N_29,In_485);
and U370 (N_370,N_301,In_251);
or U371 (N_371,N_341,In_161);
or U372 (N_372,In_127,N_17);
or U373 (N_373,N_310,In_80);
nor U374 (N_374,N_316,N_20);
and U375 (N_375,N_312,N_165);
or U376 (N_376,N_306,N_319);
nor U377 (N_377,N_45,In_450);
or U378 (N_378,In_308,N_211);
or U379 (N_379,In_248,N_287);
and U380 (N_380,N_188,N_324);
and U381 (N_381,N_332,In_296);
nor U382 (N_382,N_320,N_216);
nor U383 (N_383,N_106,N_262);
and U384 (N_384,N_292,In_407);
and U385 (N_385,In_405,N_162);
xnor U386 (N_386,N_230,In_412);
or U387 (N_387,N_115,N_226);
or U388 (N_388,In_51,N_321);
nand U389 (N_389,N_315,In_58);
nor U390 (N_390,N_331,N_289);
and U391 (N_391,N_272,In_494);
or U392 (N_392,N_302,N_111);
nand U393 (N_393,N_329,N_256);
xor U394 (N_394,N_305,In_3);
or U395 (N_395,N_151,N_258);
nand U396 (N_396,N_140,In_262);
and U397 (N_397,In_290,N_79);
xnor U398 (N_398,N_268,N_136);
nand U399 (N_399,N_334,N_191);
nor U400 (N_400,N_317,N_303);
or U401 (N_401,N_366,N_359);
and U402 (N_402,N_375,N_343);
nand U403 (N_403,In_241,N_371);
or U404 (N_404,In_183,In_384);
nand U405 (N_405,N_382,N_387);
nand U406 (N_406,N_397,N_38);
nand U407 (N_407,N_388,N_297);
or U408 (N_408,N_364,N_344);
and U409 (N_409,N_376,N_78);
or U410 (N_410,N_147,N_392);
and U411 (N_411,N_354,N_326);
or U412 (N_412,N_245,N_377);
or U413 (N_413,N_356,N_342);
and U414 (N_414,N_352,N_340);
or U415 (N_415,N_386,N_391);
or U416 (N_416,N_351,N_333);
or U417 (N_417,N_399,N_307);
or U418 (N_418,In_483,N_373);
xor U419 (N_419,N_221,N_201);
nor U420 (N_420,N_362,In_399);
and U421 (N_421,N_347,N_381);
or U422 (N_422,N_353,N_361);
nand U423 (N_423,N_365,N_280);
or U424 (N_424,N_389,N_350);
or U425 (N_425,N_242,N_250);
or U426 (N_426,In_10,N_172);
or U427 (N_427,In_38,N_372);
or U428 (N_428,In_82,N_396);
nor U429 (N_429,N_355,N_248);
nor U430 (N_430,In_402,N_394);
nand U431 (N_431,N_367,N_360);
or U432 (N_432,N_393,N_325);
and U433 (N_433,N_383,N_374);
nand U434 (N_434,N_380,N_368);
nand U435 (N_435,N_187,N_154);
nand U436 (N_436,In_189,N_379);
or U437 (N_437,N_398,N_370);
nand U438 (N_438,N_338,N_328);
nand U439 (N_439,N_390,N_369);
nor U440 (N_440,N_300,N_117);
nand U441 (N_441,N_385,In_169);
nand U442 (N_442,N_345,N_358);
and U443 (N_443,N_308,N_378);
nand U444 (N_444,N_323,In_140);
xnor U445 (N_445,N_339,N_363);
and U446 (N_446,N_92,N_384);
nand U447 (N_447,N_236,N_213);
nor U448 (N_448,N_12,N_395);
nor U449 (N_449,N_327,N_357);
or U450 (N_450,N_402,N_404);
nor U451 (N_451,N_434,N_448);
and U452 (N_452,N_414,N_410);
nand U453 (N_453,N_431,N_418);
or U454 (N_454,N_407,N_433);
and U455 (N_455,N_420,N_437);
and U456 (N_456,N_416,N_417);
or U457 (N_457,N_409,N_425);
xor U458 (N_458,N_444,N_447);
nor U459 (N_459,N_415,N_406);
nor U460 (N_460,N_441,N_401);
nand U461 (N_461,N_408,N_400);
nor U462 (N_462,N_411,N_429);
and U463 (N_463,N_412,N_419);
and U464 (N_464,N_439,N_422);
xnor U465 (N_465,N_449,N_424);
or U466 (N_466,N_427,N_446);
nor U467 (N_467,N_440,N_435);
nand U468 (N_468,N_423,N_413);
and U469 (N_469,N_426,N_445);
or U470 (N_470,N_405,N_438);
or U471 (N_471,N_421,N_432);
nor U472 (N_472,N_436,N_403);
nor U473 (N_473,N_430,N_428);
and U474 (N_474,N_443,N_442);
nor U475 (N_475,N_425,N_405);
xnor U476 (N_476,N_413,N_441);
nor U477 (N_477,N_422,N_403);
and U478 (N_478,N_449,N_437);
nand U479 (N_479,N_449,N_439);
nor U480 (N_480,N_437,N_426);
or U481 (N_481,N_441,N_423);
and U482 (N_482,N_412,N_401);
nand U483 (N_483,N_428,N_434);
nor U484 (N_484,N_421,N_449);
nand U485 (N_485,N_445,N_407);
or U486 (N_486,N_417,N_423);
nor U487 (N_487,N_422,N_438);
or U488 (N_488,N_445,N_441);
nand U489 (N_489,N_403,N_430);
nor U490 (N_490,N_416,N_424);
or U491 (N_491,N_424,N_440);
nand U492 (N_492,N_410,N_433);
nor U493 (N_493,N_422,N_401);
and U494 (N_494,N_421,N_414);
nor U495 (N_495,N_414,N_439);
and U496 (N_496,N_415,N_423);
and U497 (N_497,N_412,N_443);
nor U498 (N_498,N_405,N_423);
and U499 (N_499,N_408,N_445);
nand U500 (N_500,N_463,N_478);
or U501 (N_501,N_481,N_457);
and U502 (N_502,N_454,N_458);
or U503 (N_503,N_470,N_482);
or U504 (N_504,N_467,N_484);
or U505 (N_505,N_479,N_462);
nand U506 (N_506,N_495,N_489);
nand U507 (N_507,N_475,N_491);
and U508 (N_508,N_474,N_476);
or U509 (N_509,N_468,N_455);
and U510 (N_510,N_477,N_493);
and U511 (N_511,N_486,N_473);
nand U512 (N_512,N_451,N_472);
and U513 (N_513,N_460,N_487);
nor U514 (N_514,N_485,N_459);
nor U515 (N_515,N_497,N_456);
nand U516 (N_516,N_480,N_488);
or U517 (N_517,N_452,N_496);
and U518 (N_518,N_492,N_469);
nor U519 (N_519,N_466,N_499);
nand U520 (N_520,N_465,N_471);
and U521 (N_521,N_464,N_450);
and U522 (N_522,N_453,N_490);
nor U523 (N_523,N_498,N_494);
nand U524 (N_524,N_461,N_483);
xor U525 (N_525,N_476,N_462);
nor U526 (N_526,N_486,N_488);
nand U527 (N_527,N_482,N_453);
nor U528 (N_528,N_478,N_489);
nand U529 (N_529,N_459,N_467);
or U530 (N_530,N_484,N_496);
and U531 (N_531,N_496,N_469);
and U532 (N_532,N_453,N_493);
or U533 (N_533,N_485,N_470);
or U534 (N_534,N_493,N_459);
nor U535 (N_535,N_484,N_488);
or U536 (N_536,N_467,N_479);
xnor U537 (N_537,N_454,N_488);
or U538 (N_538,N_471,N_455);
and U539 (N_539,N_470,N_451);
and U540 (N_540,N_482,N_465);
nor U541 (N_541,N_499,N_452);
nand U542 (N_542,N_480,N_486);
nand U543 (N_543,N_475,N_472);
or U544 (N_544,N_498,N_464);
or U545 (N_545,N_494,N_453);
or U546 (N_546,N_477,N_482);
nor U547 (N_547,N_498,N_469);
or U548 (N_548,N_484,N_465);
nand U549 (N_549,N_493,N_486);
and U550 (N_550,N_548,N_528);
or U551 (N_551,N_527,N_511);
and U552 (N_552,N_508,N_506);
nor U553 (N_553,N_513,N_536);
nor U554 (N_554,N_517,N_500);
nor U555 (N_555,N_544,N_505);
nor U556 (N_556,N_525,N_510);
and U557 (N_557,N_507,N_530);
nand U558 (N_558,N_526,N_509);
or U559 (N_559,N_533,N_539);
nand U560 (N_560,N_545,N_504);
nor U561 (N_561,N_520,N_515);
or U562 (N_562,N_516,N_524);
and U563 (N_563,N_532,N_521);
nand U564 (N_564,N_537,N_535);
nand U565 (N_565,N_512,N_549);
nor U566 (N_566,N_531,N_541);
or U567 (N_567,N_514,N_501);
nor U568 (N_568,N_543,N_519);
nor U569 (N_569,N_540,N_534);
or U570 (N_570,N_523,N_546);
xnor U571 (N_571,N_503,N_529);
and U572 (N_572,N_547,N_522);
or U573 (N_573,N_542,N_502);
nand U574 (N_574,N_538,N_518);
or U575 (N_575,N_521,N_503);
or U576 (N_576,N_543,N_527);
and U577 (N_577,N_537,N_541);
or U578 (N_578,N_502,N_513);
nand U579 (N_579,N_516,N_514);
and U580 (N_580,N_503,N_538);
nand U581 (N_581,N_537,N_544);
nor U582 (N_582,N_524,N_519);
nand U583 (N_583,N_544,N_511);
nor U584 (N_584,N_519,N_517);
or U585 (N_585,N_522,N_518);
and U586 (N_586,N_526,N_511);
and U587 (N_587,N_521,N_502);
and U588 (N_588,N_527,N_517);
and U589 (N_589,N_531,N_527);
or U590 (N_590,N_548,N_525);
nor U591 (N_591,N_536,N_516);
nand U592 (N_592,N_546,N_547);
or U593 (N_593,N_546,N_505);
nor U594 (N_594,N_514,N_528);
nor U595 (N_595,N_524,N_530);
xor U596 (N_596,N_540,N_505);
or U597 (N_597,N_513,N_518);
or U598 (N_598,N_545,N_518);
nor U599 (N_599,N_538,N_542);
or U600 (N_600,N_560,N_593);
or U601 (N_601,N_585,N_568);
and U602 (N_602,N_599,N_550);
nor U603 (N_603,N_582,N_595);
nand U604 (N_604,N_556,N_597);
or U605 (N_605,N_579,N_590);
and U606 (N_606,N_566,N_563);
nand U607 (N_607,N_583,N_555);
or U608 (N_608,N_558,N_596);
or U609 (N_609,N_564,N_571);
nand U610 (N_610,N_591,N_576);
nand U611 (N_611,N_572,N_554);
nor U612 (N_612,N_562,N_559);
or U613 (N_613,N_580,N_589);
and U614 (N_614,N_594,N_569);
nand U615 (N_615,N_553,N_598);
nor U616 (N_616,N_561,N_567);
nand U617 (N_617,N_557,N_584);
nand U618 (N_618,N_592,N_565);
nand U619 (N_619,N_577,N_574);
xor U620 (N_620,N_588,N_575);
or U621 (N_621,N_552,N_587);
nand U622 (N_622,N_573,N_586);
and U623 (N_623,N_551,N_581);
nor U624 (N_624,N_570,N_578);
xnor U625 (N_625,N_591,N_594);
and U626 (N_626,N_571,N_552);
nand U627 (N_627,N_583,N_572);
or U628 (N_628,N_553,N_563);
nor U629 (N_629,N_589,N_597);
and U630 (N_630,N_577,N_580);
or U631 (N_631,N_567,N_575);
or U632 (N_632,N_553,N_590);
or U633 (N_633,N_569,N_574);
or U634 (N_634,N_562,N_594);
nor U635 (N_635,N_550,N_584);
or U636 (N_636,N_582,N_590);
and U637 (N_637,N_589,N_583);
and U638 (N_638,N_594,N_578);
and U639 (N_639,N_592,N_560);
and U640 (N_640,N_564,N_551);
and U641 (N_641,N_597,N_585);
nand U642 (N_642,N_559,N_557);
or U643 (N_643,N_559,N_582);
nand U644 (N_644,N_552,N_560);
and U645 (N_645,N_578,N_572);
nor U646 (N_646,N_560,N_582);
or U647 (N_647,N_595,N_583);
and U648 (N_648,N_586,N_563);
nand U649 (N_649,N_570,N_583);
and U650 (N_650,N_624,N_608);
nor U651 (N_651,N_631,N_609);
nand U652 (N_652,N_628,N_612);
nand U653 (N_653,N_630,N_643);
nand U654 (N_654,N_638,N_620);
nand U655 (N_655,N_648,N_633);
nand U656 (N_656,N_636,N_635);
nor U657 (N_657,N_647,N_621);
and U658 (N_658,N_607,N_637);
nor U659 (N_659,N_601,N_611);
nand U660 (N_660,N_629,N_649);
and U661 (N_661,N_602,N_640);
nor U662 (N_662,N_626,N_622);
xnor U663 (N_663,N_603,N_639);
or U664 (N_664,N_615,N_619);
nor U665 (N_665,N_605,N_645);
nand U666 (N_666,N_600,N_604);
or U667 (N_667,N_623,N_614);
or U668 (N_668,N_610,N_642);
nor U669 (N_669,N_646,N_625);
nand U670 (N_670,N_641,N_617);
or U671 (N_671,N_632,N_634);
nand U672 (N_672,N_644,N_616);
or U673 (N_673,N_606,N_618);
xor U674 (N_674,N_627,N_613);
and U675 (N_675,N_605,N_614);
or U676 (N_676,N_617,N_645);
or U677 (N_677,N_608,N_636);
nand U678 (N_678,N_610,N_635);
and U679 (N_679,N_619,N_610);
or U680 (N_680,N_630,N_642);
xor U681 (N_681,N_638,N_603);
nand U682 (N_682,N_640,N_611);
nor U683 (N_683,N_638,N_615);
or U684 (N_684,N_606,N_633);
nand U685 (N_685,N_613,N_646);
nand U686 (N_686,N_619,N_629);
or U687 (N_687,N_605,N_611);
and U688 (N_688,N_619,N_641);
and U689 (N_689,N_609,N_623);
or U690 (N_690,N_621,N_603);
or U691 (N_691,N_609,N_639);
or U692 (N_692,N_629,N_602);
nor U693 (N_693,N_639,N_630);
or U694 (N_694,N_640,N_639);
nor U695 (N_695,N_625,N_641);
nor U696 (N_696,N_626,N_604);
or U697 (N_697,N_616,N_632);
and U698 (N_698,N_619,N_627);
nand U699 (N_699,N_600,N_628);
nand U700 (N_700,N_691,N_668);
and U701 (N_701,N_669,N_686);
nand U702 (N_702,N_697,N_687);
and U703 (N_703,N_694,N_681);
xor U704 (N_704,N_665,N_675);
nor U705 (N_705,N_690,N_655);
or U706 (N_706,N_678,N_696);
and U707 (N_707,N_679,N_663);
nand U708 (N_708,N_698,N_667);
and U709 (N_709,N_673,N_692);
nand U710 (N_710,N_670,N_695);
and U711 (N_711,N_688,N_666);
and U712 (N_712,N_661,N_659);
and U713 (N_713,N_653,N_676);
nor U714 (N_714,N_664,N_652);
nand U715 (N_715,N_650,N_651);
nand U716 (N_716,N_671,N_657);
or U717 (N_717,N_699,N_672);
nand U718 (N_718,N_654,N_684);
nor U719 (N_719,N_662,N_660);
nor U720 (N_720,N_674,N_682);
nand U721 (N_721,N_677,N_685);
or U722 (N_722,N_683,N_656);
and U723 (N_723,N_689,N_693);
or U724 (N_724,N_680,N_658);
or U725 (N_725,N_699,N_697);
nand U726 (N_726,N_658,N_651);
and U727 (N_727,N_680,N_668);
and U728 (N_728,N_662,N_691);
and U729 (N_729,N_675,N_668);
and U730 (N_730,N_698,N_684);
or U731 (N_731,N_683,N_687);
nor U732 (N_732,N_660,N_690);
and U733 (N_733,N_666,N_684);
nand U734 (N_734,N_651,N_669);
xor U735 (N_735,N_661,N_663);
nand U736 (N_736,N_656,N_663);
and U737 (N_737,N_662,N_680);
nor U738 (N_738,N_687,N_690);
or U739 (N_739,N_666,N_677);
xor U740 (N_740,N_664,N_655);
nand U741 (N_741,N_698,N_694);
nand U742 (N_742,N_664,N_653);
or U743 (N_743,N_678,N_654);
nand U744 (N_744,N_663,N_698);
nor U745 (N_745,N_658,N_682);
nand U746 (N_746,N_699,N_681);
nand U747 (N_747,N_690,N_669);
and U748 (N_748,N_673,N_650);
nor U749 (N_749,N_667,N_662);
xor U750 (N_750,N_717,N_702);
nand U751 (N_751,N_705,N_748);
nor U752 (N_752,N_725,N_703);
nor U753 (N_753,N_704,N_746);
nor U754 (N_754,N_700,N_714);
nor U755 (N_755,N_706,N_718);
nand U756 (N_756,N_745,N_708);
xnor U757 (N_757,N_738,N_724);
or U758 (N_758,N_735,N_716);
nand U759 (N_759,N_744,N_723);
nor U760 (N_760,N_721,N_719);
or U761 (N_761,N_720,N_726);
or U762 (N_762,N_734,N_712);
or U763 (N_763,N_741,N_747);
nand U764 (N_764,N_736,N_707);
nand U765 (N_765,N_713,N_740);
nand U766 (N_766,N_711,N_742);
nand U767 (N_767,N_739,N_737);
or U768 (N_768,N_715,N_722);
or U769 (N_769,N_709,N_730);
or U770 (N_770,N_749,N_743);
nand U771 (N_771,N_728,N_731);
nand U772 (N_772,N_710,N_732);
or U773 (N_773,N_729,N_727);
and U774 (N_774,N_701,N_733);
or U775 (N_775,N_725,N_734);
and U776 (N_776,N_732,N_748);
xnor U777 (N_777,N_701,N_732);
xnor U778 (N_778,N_743,N_704);
nor U779 (N_779,N_705,N_725);
and U780 (N_780,N_719,N_739);
or U781 (N_781,N_748,N_746);
nand U782 (N_782,N_700,N_718);
and U783 (N_783,N_715,N_706);
and U784 (N_784,N_704,N_701);
nand U785 (N_785,N_718,N_736);
and U786 (N_786,N_714,N_711);
nand U787 (N_787,N_721,N_744);
nand U788 (N_788,N_716,N_741);
and U789 (N_789,N_703,N_721);
and U790 (N_790,N_705,N_747);
nand U791 (N_791,N_734,N_726);
nand U792 (N_792,N_706,N_741);
or U793 (N_793,N_705,N_744);
nand U794 (N_794,N_705,N_732);
and U795 (N_795,N_732,N_736);
and U796 (N_796,N_743,N_718);
nor U797 (N_797,N_737,N_701);
nand U798 (N_798,N_749,N_732);
and U799 (N_799,N_730,N_749);
and U800 (N_800,N_772,N_780);
nand U801 (N_801,N_768,N_794);
or U802 (N_802,N_793,N_761);
and U803 (N_803,N_777,N_786);
and U804 (N_804,N_764,N_762);
or U805 (N_805,N_756,N_751);
and U806 (N_806,N_785,N_757);
nor U807 (N_807,N_787,N_760);
nand U808 (N_808,N_784,N_753);
nor U809 (N_809,N_765,N_798);
nand U810 (N_810,N_755,N_797);
nand U811 (N_811,N_795,N_782);
and U812 (N_812,N_783,N_767);
or U813 (N_813,N_769,N_776);
nand U814 (N_814,N_779,N_788);
and U815 (N_815,N_774,N_778);
and U816 (N_816,N_799,N_752);
nor U817 (N_817,N_781,N_750);
or U818 (N_818,N_790,N_796);
or U819 (N_819,N_754,N_766);
nor U820 (N_820,N_791,N_775);
and U821 (N_821,N_763,N_789);
or U822 (N_822,N_773,N_759);
and U823 (N_823,N_758,N_770);
or U824 (N_824,N_771,N_792);
or U825 (N_825,N_782,N_765);
nand U826 (N_826,N_750,N_779);
nor U827 (N_827,N_797,N_774);
nor U828 (N_828,N_766,N_750);
nand U829 (N_829,N_783,N_797);
or U830 (N_830,N_760,N_796);
and U831 (N_831,N_788,N_796);
nor U832 (N_832,N_776,N_779);
or U833 (N_833,N_774,N_757);
and U834 (N_834,N_774,N_764);
and U835 (N_835,N_799,N_754);
nor U836 (N_836,N_784,N_762);
nand U837 (N_837,N_788,N_769);
nand U838 (N_838,N_766,N_782);
or U839 (N_839,N_786,N_752);
nor U840 (N_840,N_797,N_765);
or U841 (N_841,N_763,N_770);
nand U842 (N_842,N_786,N_762);
nand U843 (N_843,N_796,N_770);
nand U844 (N_844,N_784,N_787);
nand U845 (N_845,N_778,N_793);
and U846 (N_846,N_780,N_777);
or U847 (N_847,N_751,N_755);
nand U848 (N_848,N_776,N_772);
and U849 (N_849,N_793,N_786);
nand U850 (N_850,N_809,N_847);
nand U851 (N_851,N_839,N_848);
and U852 (N_852,N_800,N_819);
nand U853 (N_853,N_849,N_842);
or U854 (N_854,N_834,N_820);
and U855 (N_855,N_845,N_822);
or U856 (N_856,N_827,N_818);
nor U857 (N_857,N_836,N_808);
nor U858 (N_858,N_830,N_841);
nand U859 (N_859,N_831,N_815);
or U860 (N_860,N_814,N_817);
nor U861 (N_861,N_825,N_838);
nor U862 (N_862,N_835,N_810);
or U863 (N_863,N_816,N_844);
and U864 (N_864,N_846,N_811);
and U865 (N_865,N_806,N_843);
xor U866 (N_866,N_803,N_801);
nor U867 (N_867,N_832,N_833);
and U868 (N_868,N_807,N_813);
nand U869 (N_869,N_823,N_812);
nand U870 (N_870,N_840,N_804);
or U871 (N_871,N_828,N_826);
or U872 (N_872,N_805,N_821);
and U873 (N_873,N_802,N_829);
nand U874 (N_874,N_837,N_824);
or U875 (N_875,N_812,N_844);
and U876 (N_876,N_814,N_822);
and U877 (N_877,N_847,N_837);
nand U878 (N_878,N_845,N_842);
or U879 (N_879,N_832,N_811);
nand U880 (N_880,N_820,N_821);
nor U881 (N_881,N_847,N_824);
and U882 (N_882,N_809,N_813);
nor U883 (N_883,N_808,N_812);
and U884 (N_884,N_824,N_846);
and U885 (N_885,N_808,N_831);
nor U886 (N_886,N_808,N_804);
or U887 (N_887,N_839,N_835);
and U888 (N_888,N_803,N_822);
nor U889 (N_889,N_800,N_816);
or U890 (N_890,N_803,N_812);
or U891 (N_891,N_845,N_808);
and U892 (N_892,N_830,N_828);
xnor U893 (N_893,N_832,N_809);
or U894 (N_894,N_829,N_807);
and U895 (N_895,N_828,N_823);
and U896 (N_896,N_813,N_825);
nand U897 (N_897,N_846,N_847);
or U898 (N_898,N_800,N_820);
nor U899 (N_899,N_804,N_806);
nor U900 (N_900,N_855,N_898);
and U901 (N_901,N_892,N_899);
nand U902 (N_902,N_859,N_886);
and U903 (N_903,N_863,N_878);
nor U904 (N_904,N_853,N_869);
and U905 (N_905,N_852,N_856);
nand U906 (N_906,N_873,N_887);
nand U907 (N_907,N_880,N_860);
or U908 (N_908,N_866,N_888);
or U909 (N_909,N_868,N_861);
nor U910 (N_910,N_851,N_854);
nand U911 (N_911,N_872,N_876);
and U912 (N_912,N_858,N_881);
and U913 (N_913,N_875,N_865);
and U914 (N_914,N_889,N_882);
and U915 (N_915,N_896,N_897);
nor U916 (N_916,N_870,N_864);
nand U917 (N_917,N_884,N_890);
or U918 (N_918,N_893,N_895);
and U919 (N_919,N_877,N_885);
nand U920 (N_920,N_891,N_871);
or U921 (N_921,N_857,N_850);
or U922 (N_922,N_883,N_867);
nor U923 (N_923,N_894,N_862);
or U924 (N_924,N_874,N_879);
nor U925 (N_925,N_861,N_885);
nand U926 (N_926,N_897,N_852);
or U927 (N_927,N_851,N_877);
and U928 (N_928,N_873,N_875);
nor U929 (N_929,N_872,N_888);
nand U930 (N_930,N_878,N_875);
nor U931 (N_931,N_878,N_862);
nand U932 (N_932,N_872,N_899);
or U933 (N_933,N_868,N_854);
or U934 (N_934,N_857,N_858);
or U935 (N_935,N_873,N_898);
or U936 (N_936,N_882,N_892);
nand U937 (N_937,N_894,N_869);
nand U938 (N_938,N_881,N_861);
and U939 (N_939,N_852,N_860);
or U940 (N_940,N_881,N_862);
or U941 (N_941,N_880,N_868);
nand U942 (N_942,N_861,N_894);
and U943 (N_943,N_887,N_882);
or U944 (N_944,N_851,N_852);
xnor U945 (N_945,N_862,N_865);
and U946 (N_946,N_854,N_858);
or U947 (N_947,N_882,N_878);
or U948 (N_948,N_887,N_856);
and U949 (N_949,N_870,N_898);
and U950 (N_950,N_918,N_924);
nand U951 (N_951,N_923,N_936);
nand U952 (N_952,N_937,N_926);
nand U953 (N_953,N_909,N_935);
or U954 (N_954,N_944,N_932);
or U955 (N_955,N_921,N_906);
nor U956 (N_956,N_920,N_943);
nor U957 (N_957,N_945,N_940);
nand U958 (N_958,N_904,N_910);
or U959 (N_959,N_946,N_930);
nand U960 (N_960,N_917,N_933);
nand U961 (N_961,N_927,N_922);
or U962 (N_962,N_905,N_902);
or U963 (N_963,N_939,N_925);
xnor U964 (N_964,N_915,N_914);
and U965 (N_965,N_942,N_901);
nand U966 (N_966,N_907,N_931);
nor U967 (N_967,N_900,N_947);
nand U968 (N_968,N_908,N_912);
or U969 (N_969,N_911,N_928);
nand U970 (N_970,N_941,N_903);
nand U971 (N_971,N_934,N_949);
or U972 (N_972,N_919,N_948);
and U973 (N_973,N_916,N_938);
nand U974 (N_974,N_913,N_929);
and U975 (N_975,N_905,N_940);
nor U976 (N_976,N_935,N_920);
and U977 (N_977,N_909,N_937);
and U978 (N_978,N_932,N_934);
nand U979 (N_979,N_904,N_900);
or U980 (N_980,N_901,N_909);
and U981 (N_981,N_929,N_928);
and U982 (N_982,N_911,N_915);
or U983 (N_983,N_910,N_949);
nor U984 (N_984,N_939,N_915);
nand U985 (N_985,N_945,N_944);
or U986 (N_986,N_934,N_902);
or U987 (N_987,N_904,N_925);
nor U988 (N_988,N_919,N_946);
nor U989 (N_989,N_941,N_931);
nand U990 (N_990,N_941,N_909);
nand U991 (N_991,N_904,N_926);
nor U992 (N_992,N_922,N_925);
and U993 (N_993,N_904,N_923);
nand U994 (N_994,N_925,N_921);
nor U995 (N_995,N_937,N_943);
and U996 (N_996,N_922,N_932);
nor U997 (N_997,N_932,N_939);
or U998 (N_998,N_942,N_923);
nand U999 (N_999,N_939,N_922);
nand U1000 (N_1000,N_998,N_951);
nor U1001 (N_1001,N_993,N_968);
or U1002 (N_1002,N_984,N_985);
or U1003 (N_1003,N_953,N_988);
nand U1004 (N_1004,N_960,N_973);
nand U1005 (N_1005,N_977,N_969);
and U1006 (N_1006,N_978,N_964);
nor U1007 (N_1007,N_972,N_963);
nand U1008 (N_1008,N_979,N_958);
and U1009 (N_1009,N_991,N_996);
nor U1010 (N_1010,N_961,N_954);
or U1011 (N_1011,N_982,N_970);
and U1012 (N_1012,N_976,N_959);
nand U1013 (N_1013,N_955,N_965);
or U1014 (N_1014,N_986,N_950);
nand U1015 (N_1015,N_987,N_952);
and U1016 (N_1016,N_994,N_956);
and U1017 (N_1017,N_997,N_971);
nor U1018 (N_1018,N_995,N_974);
nor U1019 (N_1019,N_980,N_967);
nand U1020 (N_1020,N_975,N_981);
nand U1021 (N_1021,N_992,N_990);
or U1022 (N_1022,N_999,N_966);
nand U1023 (N_1023,N_957,N_989);
nand U1024 (N_1024,N_983,N_962);
nor U1025 (N_1025,N_953,N_960);
nand U1026 (N_1026,N_976,N_993);
nand U1027 (N_1027,N_958,N_967);
nor U1028 (N_1028,N_990,N_971);
and U1029 (N_1029,N_967,N_965);
or U1030 (N_1030,N_967,N_963);
nand U1031 (N_1031,N_972,N_970);
and U1032 (N_1032,N_973,N_955);
and U1033 (N_1033,N_972,N_953);
and U1034 (N_1034,N_980,N_994);
nand U1035 (N_1035,N_985,N_967);
nand U1036 (N_1036,N_974,N_975);
and U1037 (N_1037,N_965,N_986);
nand U1038 (N_1038,N_955,N_988);
and U1039 (N_1039,N_982,N_965);
xor U1040 (N_1040,N_956,N_971);
or U1041 (N_1041,N_994,N_985);
and U1042 (N_1042,N_955,N_983);
nor U1043 (N_1043,N_998,N_956);
nand U1044 (N_1044,N_983,N_956);
nand U1045 (N_1045,N_972,N_995);
or U1046 (N_1046,N_973,N_954);
nor U1047 (N_1047,N_975,N_990);
and U1048 (N_1048,N_995,N_984);
xnor U1049 (N_1049,N_975,N_976);
and U1050 (N_1050,N_1045,N_1049);
or U1051 (N_1051,N_1047,N_1038);
nand U1052 (N_1052,N_1010,N_1015);
nand U1053 (N_1053,N_1003,N_1013);
and U1054 (N_1054,N_1020,N_1005);
nand U1055 (N_1055,N_1034,N_1024);
or U1056 (N_1056,N_1048,N_1025);
or U1057 (N_1057,N_1000,N_1028);
or U1058 (N_1058,N_1008,N_1011);
nand U1059 (N_1059,N_1041,N_1042);
and U1060 (N_1060,N_1031,N_1018);
xor U1061 (N_1061,N_1004,N_1002);
nor U1062 (N_1062,N_1026,N_1029);
and U1063 (N_1063,N_1033,N_1044);
or U1064 (N_1064,N_1046,N_1007);
or U1065 (N_1065,N_1030,N_1021);
nand U1066 (N_1066,N_1036,N_1017);
nand U1067 (N_1067,N_1016,N_1039);
nand U1068 (N_1068,N_1014,N_1040);
and U1069 (N_1069,N_1022,N_1032);
nand U1070 (N_1070,N_1035,N_1037);
and U1071 (N_1071,N_1006,N_1009);
and U1072 (N_1072,N_1001,N_1023);
nor U1073 (N_1073,N_1043,N_1012);
xnor U1074 (N_1074,N_1019,N_1027);
nand U1075 (N_1075,N_1009,N_1004);
nor U1076 (N_1076,N_1002,N_1014);
nand U1077 (N_1077,N_1000,N_1039);
nand U1078 (N_1078,N_1027,N_1013);
nor U1079 (N_1079,N_1027,N_1029);
and U1080 (N_1080,N_1020,N_1025);
nor U1081 (N_1081,N_1041,N_1021);
and U1082 (N_1082,N_1000,N_1008);
nand U1083 (N_1083,N_1000,N_1013);
nor U1084 (N_1084,N_1027,N_1015);
nand U1085 (N_1085,N_1040,N_1011);
and U1086 (N_1086,N_1016,N_1023);
nand U1087 (N_1087,N_1028,N_1036);
or U1088 (N_1088,N_1026,N_1007);
or U1089 (N_1089,N_1038,N_1029);
nand U1090 (N_1090,N_1049,N_1007);
nand U1091 (N_1091,N_1039,N_1010);
and U1092 (N_1092,N_1011,N_1019);
nor U1093 (N_1093,N_1005,N_1016);
and U1094 (N_1094,N_1045,N_1003);
nor U1095 (N_1095,N_1038,N_1009);
nand U1096 (N_1096,N_1028,N_1033);
or U1097 (N_1097,N_1030,N_1008);
nor U1098 (N_1098,N_1040,N_1010);
nor U1099 (N_1099,N_1027,N_1039);
and U1100 (N_1100,N_1057,N_1076);
xnor U1101 (N_1101,N_1094,N_1078);
nor U1102 (N_1102,N_1059,N_1081);
or U1103 (N_1103,N_1065,N_1071);
nand U1104 (N_1104,N_1069,N_1098);
nand U1105 (N_1105,N_1056,N_1090);
and U1106 (N_1106,N_1054,N_1064);
nor U1107 (N_1107,N_1063,N_1084);
nand U1108 (N_1108,N_1088,N_1066);
nand U1109 (N_1109,N_1095,N_1072);
nor U1110 (N_1110,N_1080,N_1061);
nand U1111 (N_1111,N_1091,N_1050);
and U1112 (N_1112,N_1058,N_1079);
nand U1113 (N_1113,N_1097,N_1052);
and U1114 (N_1114,N_1082,N_1087);
nor U1115 (N_1115,N_1075,N_1089);
nand U1116 (N_1116,N_1051,N_1085);
nor U1117 (N_1117,N_1073,N_1062);
or U1118 (N_1118,N_1083,N_1053);
nor U1119 (N_1119,N_1092,N_1086);
and U1120 (N_1120,N_1060,N_1096);
or U1121 (N_1121,N_1068,N_1074);
or U1122 (N_1122,N_1077,N_1070);
nor U1123 (N_1123,N_1067,N_1099);
nor U1124 (N_1124,N_1055,N_1093);
and U1125 (N_1125,N_1085,N_1090);
and U1126 (N_1126,N_1089,N_1097);
and U1127 (N_1127,N_1059,N_1051);
nor U1128 (N_1128,N_1055,N_1053);
and U1129 (N_1129,N_1099,N_1052);
or U1130 (N_1130,N_1088,N_1070);
nand U1131 (N_1131,N_1053,N_1092);
and U1132 (N_1132,N_1084,N_1071);
or U1133 (N_1133,N_1074,N_1097);
and U1134 (N_1134,N_1067,N_1081);
nand U1135 (N_1135,N_1070,N_1093);
and U1136 (N_1136,N_1086,N_1076);
and U1137 (N_1137,N_1059,N_1072);
nand U1138 (N_1138,N_1086,N_1066);
and U1139 (N_1139,N_1083,N_1078);
nand U1140 (N_1140,N_1080,N_1062);
nand U1141 (N_1141,N_1092,N_1055);
and U1142 (N_1142,N_1061,N_1075);
and U1143 (N_1143,N_1061,N_1071);
and U1144 (N_1144,N_1052,N_1066);
nor U1145 (N_1145,N_1063,N_1075);
xor U1146 (N_1146,N_1064,N_1097);
nor U1147 (N_1147,N_1090,N_1092);
and U1148 (N_1148,N_1065,N_1093);
nor U1149 (N_1149,N_1056,N_1050);
or U1150 (N_1150,N_1131,N_1126);
nor U1151 (N_1151,N_1110,N_1108);
nand U1152 (N_1152,N_1112,N_1133);
and U1153 (N_1153,N_1134,N_1109);
or U1154 (N_1154,N_1149,N_1123);
and U1155 (N_1155,N_1107,N_1114);
or U1156 (N_1156,N_1143,N_1145);
xnor U1157 (N_1157,N_1144,N_1146);
or U1158 (N_1158,N_1142,N_1136);
nor U1159 (N_1159,N_1111,N_1132);
nand U1160 (N_1160,N_1104,N_1115);
nand U1161 (N_1161,N_1140,N_1137);
nor U1162 (N_1162,N_1120,N_1113);
or U1163 (N_1163,N_1117,N_1130);
and U1164 (N_1164,N_1102,N_1122);
and U1165 (N_1165,N_1128,N_1100);
and U1166 (N_1166,N_1135,N_1147);
nand U1167 (N_1167,N_1139,N_1129);
nor U1168 (N_1168,N_1124,N_1125);
nor U1169 (N_1169,N_1106,N_1105);
nor U1170 (N_1170,N_1103,N_1141);
nor U1171 (N_1171,N_1127,N_1119);
or U1172 (N_1172,N_1121,N_1148);
and U1173 (N_1173,N_1138,N_1101);
xnor U1174 (N_1174,N_1118,N_1116);
nor U1175 (N_1175,N_1106,N_1102);
and U1176 (N_1176,N_1149,N_1112);
or U1177 (N_1177,N_1142,N_1146);
nand U1178 (N_1178,N_1119,N_1131);
or U1179 (N_1179,N_1100,N_1141);
nor U1180 (N_1180,N_1108,N_1128);
or U1181 (N_1181,N_1130,N_1113);
nor U1182 (N_1182,N_1145,N_1140);
or U1183 (N_1183,N_1120,N_1122);
or U1184 (N_1184,N_1147,N_1134);
or U1185 (N_1185,N_1140,N_1104);
or U1186 (N_1186,N_1114,N_1149);
nand U1187 (N_1187,N_1105,N_1131);
nand U1188 (N_1188,N_1145,N_1133);
or U1189 (N_1189,N_1135,N_1115);
and U1190 (N_1190,N_1136,N_1103);
xnor U1191 (N_1191,N_1116,N_1140);
and U1192 (N_1192,N_1106,N_1149);
or U1193 (N_1193,N_1127,N_1111);
nor U1194 (N_1194,N_1124,N_1120);
xor U1195 (N_1195,N_1108,N_1119);
and U1196 (N_1196,N_1130,N_1109);
or U1197 (N_1197,N_1125,N_1115);
nand U1198 (N_1198,N_1132,N_1141);
nand U1199 (N_1199,N_1130,N_1133);
nand U1200 (N_1200,N_1168,N_1178);
nor U1201 (N_1201,N_1182,N_1199);
and U1202 (N_1202,N_1188,N_1158);
nor U1203 (N_1203,N_1154,N_1192);
nor U1204 (N_1204,N_1163,N_1151);
nor U1205 (N_1205,N_1194,N_1167);
nand U1206 (N_1206,N_1150,N_1197);
nor U1207 (N_1207,N_1170,N_1185);
nand U1208 (N_1208,N_1156,N_1175);
nand U1209 (N_1209,N_1161,N_1196);
or U1210 (N_1210,N_1172,N_1162);
nor U1211 (N_1211,N_1160,N_1166);
and U1212 (N_1212,N_1183,N_1184);
or U1213 (N_1213,N_1193,N_1187);
nand U1214 (N_1214,N_1198,N_1171);
nand U1215 (N_1215,N_1165,N_1180);
and U1216 (N_1216,N_1179,N_1186);
nor U1217 (N_1217,N_1177,N_1152);
and U1218 (N_1218,N_1176,N_1169);
or U1219 (N_1219,N_1164,N_1157);
and U1220 (N_1220,N_1190,N_1195);
and U1221 (N_1221,N_1173,N_1181);
and U1222 (N_1222,N_1159,N_1155);
nor U1223 (N_1223,N_1174,N_1189);
or U1224 (N_1224,N_1153,N_1191);
nand U1225 (N_1225,N_1181,N_1152);
nand U1226 (N_1226,N_1191,N_1174);
nor U1227 (N_1227,N_1191,N_1184);
and U1228 (N_1228,N_1168,N_1150);
nor U1229 (N_1229,N_1188,N_1195);
nor U1230 (N_1230,N_1162,N_1180);
nor U1231 (N_1231,N_1169,N_1190);
nand U1232 (N_1232,N_1156,N_1150);
and U1233 (N_1233,N_1186,N_1188);
or U1234 (N_1234,N_1198,N_1194);
and U1235 (N_1235,N_1151,N_1157);
or U1236 (N_1236,N_1197,N_1158);
and U1237 (N_1237,N_1166,N_1159);
nor U1238 (N_1238,N_1183,N_1164);
and U1239 (N_1239,N_1150,N_1160);
or U1240 (N_1240,N_1168,N_1188);
nand U1241 (N_1241,N_1153,N_1163);
or U1242 (N_1242,N_1176,N_1180);
or U1243 (N_1243,N_1154,N_1185);
nor U1244 (N_1244,N_1177,N_1170);
nand U1245 (N_1245,N_1173,N_1179);
or U1246 (N_1246,N_1198,N_1152);
or U1247 (N_1247,N_1196,N_1160);
or U1248 (N_1248,N_1195,N_1182);
and U1249 (N_1249,N_1199,N_1193);
or U1250 (N_1250,N_1227,N_1240);
and U1251 (N_1251,N_1214,N_1246);
nor U1252 (N_1252,N_1249,N_1202);
nor U1253 (N_1253,N_1216,N_1237);
nand U1254 (N_1254,N_1205,N_1220);
and U1255 (N_1255,N_1211,N_1239);
nand U1256 (N_1256,N_1203,N_1244);
or U1257 (N_1257,N_1221,N_1248);
or U1258 (N_1258,N_1218,N_1247);
nor U1259 (N_1259,N_1228,N_1231);
and U1260 (N_1260,N_1245,N_1201);
and U1261 (N_1261,N_1215,N_1209);
xnor U1262 (N_1262,N_1235,N_1229);
nor U1263 (N_1263,N_1226,N_1213);
nor U1264 (N_1264,N_1241,N_1222);
and U1265 (N_1265,N_1206,N_1208);
and U1266 (N_1266,N_1242,N_1234);
nor U1267 (N_1267,N_1232,N_1219);
or U1268 (N_1268,N_1210,N_1223);
and U1269 (N_1269,N_1212,N_1238);
nand U1270 (N_1270,N_1200,N_1225);
xnor U1271 (N_1271,N_1243,N_1207);
xnor U1272 (N_1272,N_1204,N_1224);
xnor U1273 (N_1273,N_1236,N_1233);
nand U1274 (N_1274,N_1217,N_1230);
nor U1275 (N_1275,N_1248,N_1214);
or U1276 (N_1276,N_1209,N_1230);
or U1277 (N_1277,N_1217,N_1214);
or U1278 (N_1278,N_1201,N_1246);
and U1279 (N_1279,N_1246,N_1217);
and U1280 (N_1280,N_1239,N_1220);
and U1281 (N_1281,N_1247,N_1235);
or U1282 (N_1282,N_1246,N_1234);
and U1283 (N_1283,N_1247,N_1217);
and U1284 (N_1284,N_1242,N_1231);
nand U1285 (N_1285,N_1206,N_1244);
nor U1286 (N_1286,N_1212,N_1216);
or U1287 (N_1287,N_1206,N_1212);
nor U1288 (N_1288,N_1228,N_1212);
or U1289 (N_1289,N_1205,N_1239);
or U1290 (N_1290,N_1205,N_1216);
or U1291 (N_1291,N_1207,N_1244);
or U1292 (N_1292,N_1239,N_1237);
or U1293 (N_1293,N_1238,N_1235);
nand U1294 (N_1294,N_1212,N_1223);
and U1295 (N_1295,N_1208,N_1249);
or U1296 (N_1296,N_1243,N_1241);
nand U1297 (N_1297,N_1218,N_1225);
and U1298 (N_1298,N_1222,N_1234);
or U1299 (N_1299,N_1246,N_1236);
nand U1300 (N_1300,N_1299,N_1287);
or U1301 (N_1301,N_1283,N_1297);
or U1302 (N_1302,N_1296,N_1258);
and U1303 (N_1303,N_1268,N_1280);
or U1304 (N_1304,N_1264,N_1262);
or U1305 (N_1305,N_1266,N_1298);
nor U1306 (N_1306,N_1255,N_1277);
or U1307 (N_1307,N_1286,N_1291);
nand U1308 (N_1308,N_1257,N_1260);
and U1309 (N_1309,N_1256,N_1275);
nor U1310 (N_1310,N_1253,N_1274);
and U1311 (N_1311,N_1278,N_1289);
nand U1312 (N_1312,N_1279,N_1261);
and U1313 (N_1313,N_1270,N_1290);
nand U1314 (N_1314,N_1265,N_1259);
nand U1315 (N_1315,N_1267,N_1285);
or U1316 (N_1316,N_1284,N_1295);
nor U1317 (N_1317,N_1282,N_1263);
nor U1318 (N_1318,N_1292,N_1254);
or U1319 (N_1319,N_1288,N_1252);
nor U1320 (N_1320,N_1271,N_1251);
nor U1321 (N_1321,N_1250,N_1272);
nand U1322 (N_1322,N_1293,N_1294);
nor U1323 (N_1323,N_1281,N_1273);
nor U1324 (N_1324,N_1276,N_1269);
or U1325 (N_1325,N_1290,N_1257);
nand U1326 (N_1326,N_1269,N_1277);
or U1327 (N_1327,N_1267,N_1263);
nor U1328 (N_1328,N_1286,N_1265);
or U1329 (N_1329,N_1257,N_1268);
nor U1330 (N_1330,N_1252,N_1261);
or U1331 (N_1331,N_1297,N_1299);
nand U1332 (N_1332,N_1289,N_1294);
nor U1333 (N_1333,N_1299,N_1255);
or U1334 (N_1334,N_1265,N_1283);
nand U1335 (N_1335,N_1267,N_1282);
or U1336 (N_1336,N_1291,N_1267);
or U1337 (N_1337,N_1260,N_1253);
and U1338 (N_1338,N_1270,N_1295);
xnor U1339 (N_1339,N_1289,N_1292);
and U1340 (N_1340,N_1250,N_1270);
nor U1341 (N_1341,N_1278,N_1294);
or U1342 (N_1342,N_1291,N_1274);
or U1343 (N_1343,N_1254,N_1279);
nor U1344 (N_1344,N_1265,N_1298);
or U1345 (N_1345,N_1257,N_1288);
and U1346 (N_1346,N_1298,N_1294);
nor U1347 (N_1347,N_1264,N_1289);
nor U1348 (N_1348,N_1258,N_1282);
and U1349 (N_1349,N_1257,N_1280);
nor U1350 (N_1350,N_1340,N_1316);
nor U1351 (N_1351,N_1321,N_1348);
nand U1352 (N_1352,N_1317,N_1333);
nand U1353 (N_1353,N_1300,N_1318);
and U1354 (N_1354,N_1322,N_1309);
nor U1355 (N_1355,N_1311,N_1331);
or U1356 (N_1356,N_1338,N_1302);
nand U1357 (N_1357,N_1330,N_1327);
or U1358 (N_1358,N_1347,N_1306);
nor U1359 (N_1359,N_1319,N_1332);
or U1360 (N_1360,N_1341,N_1308);
xor U1361 (N_1361,N_1314,N_1305);
or U1362 (N_1362,N_1349,N_1342);
nand U1363 (N_1363,N_1339,N_1323);
nor U1364 (N_1364,N_1310,N_1325);
and U1365 (N_1365,N_1343,N_1326);
nand U1366 (N_1366,N_1303,N_1315);
nand U1367 (N_1367,N_1344,N_1346);
or U1368 (N_1368,N_1329,N_1313);
and U1369 (N_1369,N_1304,N_1334);
nand U1370 (N_1370,N_1307,N_1335);
nand U1371 (N_1371,N_1320,N_1301);
nand U1372 (N_1372,N_1312,N_1337);
nand U1373 (N_1373,N_1336,N_1328);
or U1374 (N_1374,N_1345,N_1324);
nor U1375 (N_1375,N_1308,N_1333);
or U1376 (N_1376,N_1310,N_1339);
nor U1377 (N_1377,N_1330,N_1333);
or U1378 (N_1378,N_1340,N_1301);
and U1379 (N_1379,N_1348,N_1337);
or U1380 (N_1380,N_1322,N_1316);
nand U1381 (N_1381,N_1321,N_1329);
xnor U1382 (N_1382,N_1316,N_1332);
and U1383 (N_1383,N_1339,N_1305);
nand U1384 (N_1384,N_1320,N_1330);
nor U1385 (N_1385,N_1310,N_1306);
nor U1386 (N_1386,N_1321,N_1346);
nand U1387 (N_1387,N_1315,N_1332);
nor U1388 (N_1388,N_1300,N_1314);
or U1389 (N_1389,N_1315,N_1314);
nor U1390 (N_1390,N_1328,N_1325);
and U1391 (N_1391,N_1329,N_1326);
and U1392 (N_1392,N_1316,N_1345);
and U1393 (N_1393,N_1321,N_1338);
nor U1394 (N_1394,N_1310,N_1341);
nand U1395 (N_1395,N_1329,N_1345);
xnor U1396 (N_1396,N_1328,N_1305);
nor U1397 (N_1397,N_1317,N_1306);
nor U1398 (N_1398,N_1338,N_1311);
and U1399 (N_1399,N_1315,N_1307);
nand U1400 (N_1400,N_1366,N_1396);
nor U1401 (N_1401,N_1391,N_1377);
nor U1402 (N_1402,N_1373,N_1370);
nor U1403 (N_1403,N_1382,N_1362);
or U1404 (N_1404,N_1381,N_1379);
nand U1405 (N_1405,N_1374,N_1357);
nor U1406 (N_1406,N_1376,N_1375);
nand U1407 (N_1407,N_1361,N_1371);
nand U1408 (N_1408,N_1378,N_1397);
or U1409 (N_1409,N_1390,N_1392);
nand U1410 (N_1410,N_1383,N_1354);
nand U1411 (N_1411,N_1358,N_1364);
nand U1412 (N_1412,N_1360,N_1352);
or U1413 (N_1413,N_1398,N_1387);
and U1414 (N_1414,N_1367,N_1359);
and U1415 (N_1415,N_1368,N_1372);
nand U1416 (N_1416,N_1394,N_1399);
or U1417 (N_1417,N_1395,N_1386);
or U1418 (N_1418,N_1353,N_1356);
and U1419 (N_1419,N_1384,N_1355);
nor U1420 (N_1420,N_1380,N_1393);
and U1421 (N_1421,N_1369,N_1388);
nor U1422 (N_1422,N_1385,N_1365);
xor U1423 (N_1423,N_1363,N_1351);
and U1424 (N_1424,N_1389,N_1350);
and U1425 (N_1425,N_1369,N_1385);
nand U1426 (N_1426,N_1379,N_1359);
xor U1427 (N_1427,N_1357,N_1376);
nor U1428 (N_1428,N_1363,N_1399);
and U1429 (N_1429,N_1352,N_1392);
and U1430 (N_1430,N_1390,N_1360);
nor U1431 (N_1431,N_1383,N_1370);
and U1432 (N_1432,N_1397,N_1355);
and U1433 (N_1433,N_1386,N_1385);
nand U1434 (N_1434,N_1375,N_1390);
nand U1435 (N_1435,N_1356,N_1387);
nor U1436 (N_1436,N_1359,N_1372);
or U1437 (N_1437,N_1377,N_1350);
or U1438 (N_1438,N_1398,N_1357);
and U1439 (N_1439,N_1377,N_1378);
nor U1440 (N_1440,N_1363,N_1396);
and U1441 (N_1441,N_1355,N_1370);
and U1442 (N_1442,N_1364,N_1388);
nor U1443 (N_1443,N_1394,N_1358);
nand U1444 (N_1444,N_1373,N_1387);
or U1445 (N_1445,N_1379,N_1367);
nor U1446 (N_1446,N_1381,N_1387);
nand U1447 (N_1447,N_1350,N_1362);
xnor U1448 (N_1448,N_1358,N_1360);
nor U1449 (N_1449,N_1372,N_1392);
and U1450 (N_1450,N_1414,N_1430);
nor U1451 (N_1451,N_1441,N_1406);
nand U1452 (N_1452,N_1424,N_1427);
and U1453 (N_1453,N_1405,N_1433);
nand U1454 (N_1454,N_1407,N_1431);
and U1455 (N_1455,N_1448,N_1416);
or U1456 (N_1456,N_1408,N_1437);
nand U1457 (N_1457,N_1403,N_1421);
and U1458 (N_1458,N_1428,N_1402);
or U1459 (N_1459,N_1404,N_1435);
or U1460 (N_1460,N_1419,N_1432);
nand U1461 (N_1461,N_1415,N_1445);
nand U1462 (N_1462,N_1438,N_1411);
nand U1463 (N_1463,N_1426,N_1440);
nand U1464 (N_1464,N_1422,N_1423);
or U1465 (N_1465,N_1417,N_1444);
or U1466 (N_1466,N_1434,N_1429);
nor U1467 (N_1467,N_1409,N_1425);
and U1468 (N_1468,N_1418,N_1420);
and U1469 (N_1469,N_1412,N_1443);
nand U1470 (N_1470,N_1410,N_1439);
and U1471 (N_1471,N_1446,N_1447);
nor U1472 (N_1472,N_1400,N_1401);
xnor U1473 (N_1473,N_1442,N_1413);
and U1474 (N_1474,N_1449,N_1436);
and U1475 (N_1475,N_1410,N_1427);
nor U1476 (N_1476,N_1420,N_1413);
nand U1477 (N_1477,N_1408,N_1431);
nand U1478 (N_1478,N_1423,N_1442);
nand U1479 (N_1479,N_1410,N_1430);
or U1480 (N_1480,N_1443,N_1438);
or U1481 (N_1481,N_1408,N_1429);
nor U1482 (N_1482,N_1413,N_1402);
nand U1483 (N_1483,N_1432,N_1425);
or U1484 (N_1484,N_1430,N_1404);
or U1485 (N_1485,N_1404,N_1440);
nand U1486 (N_1486,N_1439,N_1415);
nor U1487 (N_1487,N_1445,N_1430);
or U1488 (N_1488,N_1434,N_1409);
and U1489 (N_1489,N_1428,N_1407);
xnor U1490 (N_1490,N_1411,N_1407);
nor U1491 (N_1491,N_1431,N_1400);
or U1492 (N_1492,N_1416,N_1444);
nor U1493 (N_1493,N_1448,N_1433);
or U1494 (N_1494,N_1420,N_1419);
nor U1495 (N_1495,N_1426,N_1439);
nor U1496 (N_1496,N_1439,N_1427);
or U1497 (N_1497,N_1404,N_1448);
or U1498 (N_1498,N_1436,N_1405);
or U1499 (N_1499,N_1418,N_1426);
and U1500 (N_1500,N_1484,N_1491);
nor U1501 (N_1501,N_1494,N_1489);
nor U1502 (N_1502,N_1480,N_1476);
and U1503 (N_1503,N_1497,N_1467);
or U1504 (N_1504,N_1487,N_1473);
nor U1505 (N_1505,N_1479,N_1459);
and U1506 (N_1506,N_1455,N_1460);
or U1507 (N_1507,N_1498,N_1495);
nand U1508 (N_1508,N_1469,N_1493);
and U1509 (N_1509,N_1463,N_1451);
nor U1510 (N_1510,N_1456,N_1453);
nand U1511 (N_1511,N_1477,N_1496);
or U1512 (N_1512,N_1466,N_1450);
and U1513 (N_1513,N_1472,N_1499);
and U1514 (N_1514,N_1468,N_1486);
or U1515 (N_1515,N_1488,N_1452);
nor U1516 (N_1516,N_1481,N_1464);
and U1517 (N_1517,N_1485,N_1458);
xor U1518 (N_1518,N_1492,N_1471);
nand U1519 (N_1519,N_1482,N_1461);
and U1520 (N_1520,N_1490,N_1454);
xnor U1521 (N_1521,N_1457,N_1483);
nor U1522 (N_1522,N_1478,N_1470);
nand U1523 (N_1523,N_1474,N_1462);
and U1524 (N_1524,N_1475,N_1465);
or U1525 (N_1525,N_1469,N_1453);
nor U1526 (N_1526,N_1481,N_1462);
or U1527 (N_1527,N_1452,N_1461);
and U1528 (N_1528,N_1498,N_1499);
and U1529 (N_1529,N_1461,N_1468);
nor U1530 (N_1530,N_1469,N_1454);
and U1531 (N_1531,N_1458,N_1467);
xor U1532 (N_1532,N_1488,N_1468);
nor U1533 (N_1533,N_1480,N_1451);
and U1534 (N_1534,N_1471,N_1472);
nand U1535 (N_1535,N_1482,N_1451);
and U1536 (N_1536,N_1478,N_1492);
nand U1537 (N_1537,N_1459,N_1457);
or U1538 (N_1538,N_1478,N_1467);
nor U1539 (N_1539,N_1458,N_1495);
or U1540 (N_1540,N_1468,N_1459);
nand U1541 (N_1541,N_1492,N_1470);
or U1542 (N_1542,N_1452,N_1489);
nand U1543 (N_1543,N_1454,N_1458);
nor U1544 (N_1544,N_1481,N_1468);
and U1545 (N_1545,N_1480,N_1477);
nand U1546 (N_1546,N_1490,N_1471);
nor U1547 (N_1547,N_1480,N_1492);
nand U1548 (N_1548,N_1475,N_1481);
nand U1549 (N_1549,N_1450,N_1457);
and U1550 (N_1550,N_1535,N_1514);
nand U1551 (N_1551,N_1504,N_1538);
xor U1552 (N_1552,N_1505,N_1544);
nor U1553 (N_1553,N_1500,N_1518);
and U1554 (N_1554,N_1512,N_1531);
nor U1555 (N_1555,N_1524,N_1547);
nor U1556 (N_1556,N_1533,N_1517);
nor U1557 (N_1557,N_1549,N_1502);
nand U1558 (N_1558,N_1523,N_1507);
or U1559 (N_1559,N_1537,N_1540);
nand U1560 (N_1560,N_1521,N_1542);
nor U1561 (N_1561,N_1525,N_1516);
and U1562 (N_1562,N_1541,N_1513);
and U1563 (N_1563,N_1508,N_1539);
nand U1564 (N_1564,N_1527,N_1506);
nor U1565 (N_1565,N_1520,N_1510);
or U1566 (N_1566,N_1530,N_1548);
nand U1567 (N_1567,N_1515,N_1528);
nor U1568 (N_1568,N_1503,N_1526);
and U1569 (N_1569,N_1501,N_1511);
nand U1570 (N_1570,N_1545,N_1509);
nor U1571 (N_1571,N_1529,N_1534);
nor U1572 (N_1572,N_1532,N_1536);
and U1573 (N_1573,N_1519,N_1522);
nor U1574 (N_1574,N_1546,N_1543);
or U1575 (N_1575,N_1514,N_1523);
nor U1576 (N_1576,N_1532,N_1534);
nor U1577 (N_1577,N_1520,N_1540);
or U1578 (N_1578,N_1519,N_1512);
nor U1579 (N_1579,N_1526,N_1548);
or U1580 (N_1580,N_1516,N_1522);
nand U1581 (N_1581,N_1523,N_1545);
nor U1582 (N_1582,N_1514,N_1538);
nor U1583 (N_1583,N_1526,N_1527);
and U1584 (N_1584,N_1529,N_1533);
or U1585 (N_1585,N_1517,N_1549);
nand U1586 (N_1586,N_1508,N_1520);
nand U1587 (N_1587,N_1542,N_1531);
nor U1588 (N_1588,N_1511,N_1509);
or U1589 (N_1589,N_1507,N_1547);
and U1590 (N_1590,N_1514,N_1525);
or U1591 (N_1591,N_1545,N_1526);
nor U1592 (N_1592,N_1535,N_1545);
nand U1593 (N_1593,N_1503,N_1536);
and U1594 (N_1594,N_1523,N_1536);
and U1595 (N_1595,N_1511,N_1549);
or U1596 (N_1596,N_1517,N_1516);
or U1597 (N_1597,N_1534,N_1524);
nand U1598 (N_1598,N_1549,N_1548);
or U1599 (N_1599,N_1548,N_1534);
or U1600 (N_1600,N_1588,N_1563);
or U1601 (N_1601,N_1593,N_1559);
nor U1602 (N_1602,N_1576,N_1571);
or U1603 (N_1603,N_1598,N_1567);
and U1604 (N_1604,N_1592,N_1555);
nor U1605 (N_1605,N_1586,N_1565);
nand U1606 (N_1606,N_1552,N_1580);
and U1607 (N_1607,N_1597,N_1574);
nand U1608 (N_1608,N_1550,N_1568);
nand U1609 (N_1609,N_1595,N_1590);
nand U1610 (N_1610,N_1573,N_1553);
nor U1611 (N_1611,N_1554,N_1551);
or U1612 (N_1612,N_1584,N_1564);
or U1613 (N_1613,N_1577,N_1589);
nand U1614 (N_1614,N_1582,N_1578);
nand U1615 (N_1615,N_1587,N_1591);
nor U1616 (N_1616,N_1599,N_1566);
nor U1617 (N_1617,N_1575,N_1560);
nand U1618 (N_1618,N_1557,N_1583);
and U1619 (N_1619,N_1570,N_1596);
nor U1620 (N_1620,N_1558,N_1569);
nand U1621 (N_1621,N_1572,N_1581);
or U1622 (N_1622,N_1556,N_1585);
nand U1623 (N_1623,N_1561,N_1579);
or U1624 (N_1624,N_1562,N_1594);
or U1625 (N_1625,N_1599,N_1581);
and U1626 (N_1626,N_1582,N_1584);
nand U1627 (N_1627,N_1577,N_1554);
nor U1628 (N_1628,N_1574,N_1599);
nor U1629 (N_1629,N_1576,N_1570);
and U1630 (N_1630,N_1569,N_1594);
and U1631 (N_1631,N_1571,N_1567);
xnor U1632 (N_1632,N_1599,N_1563);
or U1633 (N_1633,N_1597,N_1598);
nor U1634 (N_1634,N_1578,N_1594);
and U1635 (N_1635,N_1572,N_1560);
nor U1636 (N_1636,N_1585,N_1557);
and U1637 (N_1637,N_1567,N_1580);
nand U1638 (N_1638,N_1577,N_1558);
and U1639 (N_1639,N_1589,N_1571);
nor U1640 (N_1640,N_1586,N_1558);
and U1641 (N_1641,N_1571,N_1588);
nand U1642 (N_1642,N_1582,N_1596);
nand U1643 (N_1643,N_1568,N_1561);
nand U1644 (N_1644,N_1576,N_1567);
or U1645 (N_1645,N_1582,N_1560);
nand U1646 (N_1646,N_1553,N_1586);
nand U1647 (N_1647,N_1551,N_1581);
and U1648 (N_1648,N_1594,N_1579);
nand U1649 (N_1649,N_1560,N_1598);
nor U1650 (N_1650,N_1610,N_1642);
and U1651 (N_1651,N_1626,N_1649);
nor U1652 (N_1652,N_1623,N_1627);
and U1653 (N_1653,N_1632,N_1645);
or U1654 (N_1654,N_1612,N_1637);
or U1655 (N_1655,N_1647,N_1630);
or U1656 (N_1656,N_1639,N_1611);
nor U1657 (N_1657,N_1600,N_1604);
nand U1658 (N_1658,N_1614,N_1608);
nor U1659 (N_1659,N_1644,N_1603);
nor U1660 (N_1660,N_1617,N_1635);
or U1661 (N_1661,N_1615,N_1640);
and U1662 (N_1662,N_1634,N_1621);
or U1663 (N_1663,N_1613,N_1633);
or U1664 (N_1664,N_1636,N_1619);
nor U1665 (N_1665,N_1628,N_1646);
nor U1666 (N_1666,N_1618,N_1631);
nor U1667 (N_1667,N_1605,N_1643);
or U1668 (N_1668,N_1641,N_1602);
nand U1669 (N_1669,N_1620,N_1622);
nor U1670 (N_1670,N_1625,N_1624);
and U1671 (N_1671,N_1607,N_1648);
nand U1672 (N_1672,N_1638,N_1609);
and U1673 (N_1673,N_1601,N_1629);
or U1674 (N_1674,N_1616,N_1606);
or U1675 (N_1675,N_1605,N_1613);
or U1676 (N_1676,N_1615,N_1606);
nand U1677 (N_1677,N_1614,N_1617);
nand U1678 (N_1678,N_1641,N_1633);
and U1679 (N_1679,N_1622,N_1602);
nand U1680 (N_1680,N_1646,N_1601);
or U1681 (N_1681,N_1616,N_1636);
nand U1682 (N_1682,N_1625,N_1622);
and U1683 (N_1683,N_1631,N_1607);
and U1684 (N_1684,N_1610,N_1633);
nor U1685 (N_1685,N_1617,N_1638);
nand U1686 (N_1686,N_1636,N_1621);
xnor U1687 (N_1687,N_1622,N_1636);
and U1688 (N_1688,N_1645,N_1631);
nand U1689 (N_1689,N_1624,N_1636);
and U1690 (N_1690,N_1641,N_1607);
nor U1691 (N_1691,N_1649,N_1615);
and U1692 (N_1692,N_1618,N_1625);
nor U1693 (N_1693,N_1604,N_1630);
or U1694 (N_1694,N_1610,N_1635);
nand U1695 (N_1695,N_1647,N_1629);
and U1696 (N_1696,N_1605,N_1610);
and U1697 (N_1697,N_1621,N_1615);
nand U1698 (N_1698,N_1635,N_1643);
nor U1699 (N_1699,N_1620,N_1621);
and U1700 (N_1700,N_1688,N_1670);
or U1701 (N_1701,N_1653,N_1669);
or U1702 (N_1702,N_1687,N_1682);
and U1703 (N_1703,N_1660,N_1659);
or U1704 (N_1704,N_1698,N_1677);
nor U1705 (N_1705,N_1685,N_1690);
and U1706 (N_1706,N_1662,N_1697);
and U1707 (N_1707,N_1696,N_1651);
nand U1708 (N_1708,N_1652,N_1694);
and U1709 (N_1709,N_1668,N_1691);
or U1710 (N_1710,N_1664,N_1657);
nand U1711 (N_1711,N_1695,N_1656);
or U1712 (N_1712,N_1684,N_1675);
or U1713 (N_1713,N_1676,N_1678);
or U1714 (N_1714,N_1661,N_1672);
or U1715 (N_1715,N_1681,N_1689);
nor U1716 (N_1716,N_1654,N_1692);
or U1717 (N_1717,N_1686,N_1683);
nand U1718 (N_1718,N_1667,N_1674);
and U1719 (N_1719,N_1663,N_1680);
and U1720 (N_1720,N_1671,N_1666);
nor U1721 (N_1721,N_1673,N_1699);
and U1722 (N_1722,N_1693,N_1658);
nor U1723 (N_1723,N_1655,N_1665);
or U1724 (N_1724,N_1679,N_1650);
or U1725 (N_1725,N_1679,N_1689);
nand U1726 (N_1726,N_1681,N_1664);
nor U1727 (N_1727,N_1670,N_1663);
and U1728 (N_1728,N_1678,N_1688);
nor U1729 (N_1729,N_1681,N_1650);
nand U1730 (N_1730,N_1688,N_1686);
or U1731 (N_1731,N_1685,N_1683);
or U1732 (N_1732,N_1692,N_1699);
and U1733 (N_1733,N_1676,N_1686);
or U1734 (N_1734,N_1660,N_1674);
or U1735 (N_1735,N_1671,N_1688);
or U1736 (N_1736,N_1668,N_1689);
nor U1737 (N_1737,N_1665,N_1672);
and U1738 (N_1738,N_1651,N_1654);
or U1739 (N_1739,N_1679,N_1662);
nor U1740 (N_1740,N_1659,N_1675);
nand U1741 (N_1741,N_1655,N_1697);
nand U1742 (N_1742,N_1683,N_1665);
nand U1743 (N_1743,N_1664,N_1694);
and U1744 (N_1744,N_1666,N_1697);
nor U1745 (N_1745,N_1662,N_1685);
nor U1746 (N_1746,N_1652,N_1699);
nand U1747 (N_1747,N_1678,N_1670);
nor U1748 (N_1748,N_1698,N_1682);
and U1749 (N_1749,N_1675,N_1697);
nand U1750 (N_1750,N_1702,N_1736);
or U1751 (N_1751,N_1734,N_1717);
or U1752 (N_1752,N_1741,N_1723);
nor U1753 (N_1753,N_1744,N_1746);
nand U1754 (N_1754,N_1711,N_1743);
nor U1755 (N_1755,N_1716,N_1708);
nor U1756 (N_1756,N_1721,N_1701);
nand U1757 (N_1757,N_1738,N_1724);
nor U1758 (N_1758,N_1709,N_1729);
xor U1759 (N_1759,N_1727,N_1722);
and U1760 (N_1760,N_1732,N_1719);
nor U1761 (N_1761,N_1715,N_1706);
and U1762 (N_1762,N_1712,N_1713);
and U1763 (N_1763,N_1730,N_1704);
or U1764 (N_1764,N_1707,N_1705);
or U1765 (N_1765,N_1720,N_1735);
and U1766 (N_1766,N_1740,N_1748);
nor U1767 (N_1767,N_1731,N_1726);
xor U1768 (N_1768,N_1737,N_1733);
or U1769 (N_1769,N_1728,N_1700);
nor U1770 (N_1770,N_1703,N_1725);
nand U1771 (N_1771,N_1747,N_1714);
or U1772 (N_1772,N_1749,N_1745);
and U1773 (N_1773,N_1710,N_1739);
nand U1774 (N_1774,N_1742,N_1718);
and U1775 (N_1775,N_1747,N_1718);
or U1776 (N_1776,N_1724,N_1726);
nor U1777 (N_1777,N_1712,N_1740);
or U1778 (N_1778,N_1733,N_1716);
nor U1779 (N_1779,N_1741,N_1731);
and U1780 (N_1780,N_1734,N_1706);
nand U1781 (N_1781,N_1724,N_1721);
nor U1782 (N_1782,N_1707,N_1732);
nand U1783 (N_1783,N_1715,N_1703);
nor U1784 (N_1784,N_1732,N_1703);
and U1785 (N_1785,N_1724,N_1737);
and U1786 (N_1786,N_1730,N_1745);
or U1787 (N_1787,N_1709,N_1701);
or U1788 (N_1788,N_1713,N_1721);
or U1789 (N_1789,N_1709,N_1730);
and U1790 (N_1790,N_1748,N_1736);
nor U1791 (N_1791,N_1726,N_1714);
nand U1792 (N_1792,N_1714,N_1748);
or U1793 (N_1793,N_1722,N_1737);
nor U1794 (N_1794,N_1747,N_1721);
nand U1795 (N_1795,N_1731,N_1718);
or U1796 (N_1796,N_1749,N_1726);
or U1797 (N_1797,N_1726,N_1700);
and U1798 (N_1798,N_1710,N_1735);
and U1799 (N_1799,N_1716,N_1700);
nand U1800 (N_1800,N_1795,N_1754);
nor U1801 (N_1801,N_1784,N_1772);
nand U1802 (N_1802,N_1798,N_1780);
nand U1803 (N_1803,N_1771,N_1777);
nand U1804 (N_1804,N_1773,N_1765);
or U1805 (N_1805,N_1786,N_1787);
and U1806 (N_1806,N_1750,N_1751);
and U1807 (N_1807,N_1791,N_1783);
nor U1808 (N_1808,N_1752,N_1790);
nand U1809 (N_1809,N_1767,N_1796);
nand U1810 (N_1810,N_1760,N_1768);
xnor U1811 (N_1811,N_1758,N_1782);
nor U1812 (N_1812,N_1757,N_1774);
or U1813 (N_1813,N_1759,N_1761);
or U1814 (N_1814,N_1770,N_1799);
nand U1815 (N_1815,N_1769,N_1781);
and U1816 (N_1816,N_1766,N_1789);
or U1817 (N_1817,N_1755,N_1763);
nor U1818 (N_1818,N_1794,N_1778);
nand U1819 (N_1819,N_1779,N_1785);
nor U1820 (N_1820,N_1793,N_1788);
and U1821 (N_1821,N_1753,N_1797);
nor U1822 (N_1822,N_1775,N_1792);
and U1823 (N_1823,N_1756,N_1764);
or U1824 (N_1824,N_1762,N_1776);
and U1825 (N_1825,N_1772,N_1769);
nor U1826 (N_1826,N_1793,N_1758);
nand U1827 (N_1827,N_1782,N_1779);
or U1828 (N_1828,N_1785,N_1784);
and U1829 (N_1829,N_1781,N_1773);
nor U1830 (N_1830,N_1792,N_1759);
nor U1831 (N_1831,N_1789,N_1773);
and U1832 (N_1832,N_1772,N_1763);
or U1833 (N_1833,N_1777,N_1766);
nor U1834 (N_1834,N_1774,N_1764);
and U1835 (N_1835,N_1771,N_1788);
nor U1836 (N_1836,N_1798,N_1750);
or U1837 (N_1837,N_1754,N_1772);
nor U1838 (N_1838,N_1786,N_1788);
and U1839 (N_1839,N_1763,N_1790);
nor U1840 (N_1840,N_1782,N_1756);
and U1841 (N_1841,N_1755,N_1779);
nand U1842 (N_1842,N_1764,N_1767);
or U1843 (N_1843,N_1797,N_1768);
nand U1844 (N_1844,N_1789,N_1772);
nor U1845 (N_1845,N_1774,N_1795);
or U1846 (N_1846,N_1759,N_1775);
nor U1847 (N_1847,N_1778,N_1758);
xor U1848 (N_1848,N_1799,N_1775);
nor U1849 (N_1849,N_1758,N_1769);
or U1850 (N_1850,N_1811,N_1843);
and U1851 (N_1851,N_1815,N_1831);
or U1852 (N_1852,N_1824,N_1803);
or U1853 (N_1853,N_1846,N_1804);
nor U1854 (N_1854,N_1822,N_1819);
and U1855 (N_1855,N_1835,N_1836);
and U1856 (N_1856,N_1844,N_1818);
and U1857 (N_1857,N_1809,N_1801);
nand U1858 (N_1858,N_1800,N_1848);
nand U1859 (N_1859,N_1821,N_1838);
nor U1860 (N_1860,N_1814,N_1830);
or U1861 (N_1861,N_1847,N_1841);
nand U1862 (N_1862,N_1837,N_1825);
and U1863 (N_1863,N_1807,N_1802);
or U1864 (N_1864,N_1828,N_1805);
and U1865 (N_1865,N_1823,N_1845);
nor U1866 (N_1866,N_1832,N_1834);
nor U1867 (N_1867,N_1816,N_1810);
nor U1868 (N_1868,N_1840,N_1813);
or U1869 (N_1869,N_1842,N_1808);
nor U1870 (N_1870,N_1833,N_1849);
and U1871 (N_1871,N_1817,N_1820);
or U1872 (N_1872,N_1839,N_1827);
xor U1873 (N_1873,N_1812,N_1826);
nand U1874 (N_1874,N_1806,N_1829);
or U1875 (N_1875,N_1831,N_1847);
and U1876 (N_1876,N_1845,N_1825);
and U1877 (N_1877,N_1835,N_1802);
nand U1878 (N_1878,N_1834,N_1845);
or U1879 (N_1879,N_1830,N_1822);
nor U1880 (N_1880,N_1828,N_1804);
nor U1881 (N_1881,N_1819,N_1833);
or U1882 (N_1882,N_1824,N_1845);
or U1883 (N_1883,N_1813,N_1804);
or U1884 (N_1884,N_1800,N_1802);
or U1885 (N_1885,N_1830,N_1828);
nand U1886 (N_1886,N_1819,N_1810);
and U1887 (N_1887,N_1828,N_1801);
nand U1888 (N_1888,N_1848,N_1810);
nor U1889 (N_1889,N_1847,N_1835);
nor U1890 (N_1890,N_1822,N_1838);
nand U1891 (N_1891,N_1804,N_1840);
or U1892 (N_1892,N_1841,N_1843);
nand U1893 (N_1893,N_1805,N_1841);
nand U1894 (N_1894,N_1820,N_1831);
nor U1895 (N_1895,N_1800,N_1843);
or U1896 (N_1896,N_1843,N_1848);
nand U1897 (N_1897,N_1823,N_1849);
or U1898 (N_1898,N_1836,N_1807);
nor U1899 (N_1899,N_1811,N_1845);
nand U1900 (N_1900,N_1851,N_1858);
and U1901 (N_1901,N_1880,N_1887);
or U1902 (N_1902,N_1895,N_1892);
and U1903 (N_1903,N_1871,N_1896);
nand U1904 (N_1904,N_1877,N_1864);
nor U1905 (N_1905,N_1894,N_1898);
nand U1906 (N_1906,N_1859,N_1852);
xnor U1907 (N_1907,N_1897,N_1854);
and U1908 (N_1908,N_1891,N_1850);
nor U1909 (N_1909,N_1868,N_1899);
and U1910 (N_1910,N_1869,N_1893);
or U1911 (N_1911,N_1870,N_1855);
nor U1912 (N_1912,N_1884,N_1881);
or U1913 (N_1913,N_1867,N_1890);
or U1914 (N_1914,N_1865,N_1873);
nand U1915 (N_1915,N_1874,N_1885);
nor U1916 (N_1916,N_1882,N_1876);
and U1917 (N_1917,N_1857,N_1860);
nor U1918 (N_1918,N_1862,N_1872);
nand U1919 (N_1919,N_1853,N_1863);
or U1920 (N_1920,N_1875,N_1861);
or U1921 (N_1921,N_1856,N_1888);
nand U1922 (N_1922,N_1883,N_1879);
or U1923 (N_1923,N_1889,N_1878);
nand U1924 (N_1924,N_1886,N_1866);
and U1925 (N_1925,N_1882,N_1865);
and U1926 (N_1926,N_1874,N_1865);
nor U1927 (N_1927,N_1869,N_1851);
nand U1928 (N_1928,N_1854,N_1899);
nand U1929 (N_1929,N_1899,N_1874);
nand U1930 (N_1930,N_1888,N_1861);
nand U1931 (N_1931,N_1869,N_1855);
nand U1932 (N_1932,N_1885,N_1872);
nor U1933 (N_1933,N_1859,N_1865);
nor U1934 (N_1934,N_1869,N_1897);
and U1935 (N_1935,N_1854,N_1893);
or U1936 (N_1936,N_1863,N_1888);
and U1937 (N_1937,N_1867,N_1897);
and U1938 (N_1938,N_1893,N_1894);
nor U1939 (N_1939,N_1874,N_1877);
nor U1940 (N_1940,N_1864,N_1865);
or U1941 (N_1941,N_1888,N_1879);
nor U1942 (N_1942,N_1872,N_1891);
and U1943 (N_1943,N_1868,N_1857);
nand U1944 (N_1944,N_1899,N_1869);
nand U1945 (N_1945,N_1887,N_1891);
nand U1946 (N_1946,N_1875,N_1897);
nand U1947 (N_1947,N_1881,N_1852);
or U1948 (N_1948,N_1892,N_1874);
or U1949 (N_1949,N_1889,N_1893);
nor U1950 (N_1950,N_1937,N_1936);
nor U1951 (N_1951,N_1923,N_1922);
or U1952 (N_1952,N_1900,N_1946);
and U1953 (N_1953,N_1916,N_1917);
xnor U1954 (N_1954,N_1935,N_1941);
nor U1955 (N_1955,N_1929,N_1939);
nand U1956 (N_1956,N_1931,N_1943);
nor U1957 (N_1957,N_1924,N_1927);
and U1958 (N_1958,N_1921,N_1918);
or U1959 (N_1959,N_1940,N_1906);
and U1960 (N_1960,N_1912,N_1904);
and U1961 (N_1961,N_1908,N_1911);
or U1962 (N_1962,N_1933,N_1910);
or U1963 (N_1963,N_1945,N_1914);
nor U1964 (N_1964,N_1930,N_1925);
and U1965 (N_1965,N_1944,N_1919);
nor U1966 (N_1966,N_1915,N_1902);
and U1967 (N_1967,N_1942,N_1938);
nand U1968 (N_1968,N_1949,N_1901);
nand U1969 (N_1969,N_1909,N_1932);
nor U1970 (N_1970,N_1948,N_1934);
or U1971 (N_1971,N_1905,N_1913);
or U1972 (N_1972,N_1926,N_1928);
nor U1973 (N_1973,N_1920,N_1907);
nand U1974 (N_1974,N_1903,N_1947);
or U1975 (N_1975,N_1946,N_1932);
and U1976 (N_1976,N_1935,N_1923);
nor U1977 (N_1977,N_1940,N_1924);
and U1978 (N_1978,N_1931,N_1904);
nand U1979 (N_1979,N_1946,N_1935);
nor U1980 (N_1980,N_1906,N_1948);
and U1981 (N_1981,N_1931,N_1900);
and U1982 (N_1982,N_1924,N_1935);
xnor U1983 (N_1983,N_1926,N_1915);
or U1984 (N_1984,N_1904,N_1913);
or U1985 (N_1985,N_1939,N_1927);
and U1986 (N_1986,N_1918,N_1929);
nor U1987 (N_1987,N_1901,N_1902);
or U1988 (N_1988,N_1935,N_1907);
nand U1989 (N_1989,N_1943,N_1936);
nand U1990 (N_1990,N_1901,N_1914);
nor U1991 (N_1991,N_1911,N_1904);
and U1992 (N_1992,N_1933,N_1924);
and U1993 (N_1993,N_1920,N_1914);
and U1994 (N_1994,N_1940,N_1901);
or U1995 (N_1995,N_1932,N_1931);
and U1996 (N_1996,N_1947,N_1927);
or U1997 (N_1997,N_1914,N_1919);
nand U1998 (N_1998,N_1910,N_1904);
nand U1999 (N_1999,N_1921,N_1947);
nor U2000 (N_2000,N_1980,N_1954);
nor U2001 (N_2001,N_1966,N_1970);
nor U2002 (N_2002,N_1995,N_1975);
and U2003 (N_2003,N_1968,N_1961);
nand U2004 (N_2004,N_1988,N_1973);
or U2005 (N_2005,N_1981,N_1994);
nand U2006 (N_2006,N_1967,N_1987);
nor U2007 (N_2007,N_1974,N_1989);
or U2008 (N_2008,N_1985,N_1993);
nand U2009 (N_2009,N_1957,N_1956);
or U2010 (N_2010,N_1963,N_1986);
or U2011 (N_2011,N_1983,N_1984);
or U2012 (N_2012,N_1960,N_1982);
nand U2013 (N_2013,N_1951,N_1992);
nand U2014 (N_2014,N_1964,N_1969);
and U2015 (N_2015,N_1996,N_1971);
or U2016 (N_2016,N_1962,N_1991);
nand U2017 (N_2017,N_1979,N_1955);
nand U2018 (N_2018,N_1958,N_1965);
nor U2019 (N_2019,N_1976,N_1950);
or U2020 (N_2020,N_1999,N_1998);
nor U2021 (N_2021,N_1952,N_1978);
nand U2022 (N_2022,N_1977,N_1990);
nand U2023 (N_2023,N_1953,N_1972);
or U2024 (N_2024,N_1959,N_1997);
and U2025 (N_2025,N_1966,N_1998);
nand U2026 (N_2026,N_1950,N_1956);
and U2027 (N_2027,N_1985,N_1957);
and U2028 (N_2028,N_1967,N_1960);
nor U2029 (N_2029,N_1999,N_1996);
nand U2030 (N_2030,N_1960,N_1971);
or U2031 (N_2031,N_1972,N_1995);
or U2032 (N_2032,N_1952,N_1987);
nor U2033 (N_2033,N_1978,N_1977);
nor U2034 (N_2034,N_1960,N_1968);
nand U2035 (N_2035,N_1988,N_1985);
nor U2036 (N_2036,N_1995,N_1989);
or U2037 (N_2037,N_1996,N_1979);
nand U2038 (N_2038,N_1987,N_1984);
xnor U2039 (N_2039,N_1989,N_1969);
or U2040 (N_2040,N_1990,N_1956);
or U2041 (N_2041,N_1970,N_1996);
nand U2042 (N_2042,N_1955,N_1969);
and U2043 (N_2043,N_1980,N_1973);
nor U2044 (N_2044,N_1964,N_1963);
nor U2045 (N_2045,N_1961,N_1977);
and U2046 (N_2046,N_1995,N_1964);
and U2047 (N_2047,N_1962,N_1971);
nor U2048 (N_2048,N_1999,N_1953);
and U2049 (N_2049,N_1999,N_1989);
and U2050 (N_2050,N_2049,N_2048);
and U2051 (N_2051,N_2012,N_2033);
nor U2052 (N_2052,N_2015,N_2034);
nor U2053 (N_2053,N_2017,N_2025);
xnor U2054 (N_2054,N_2032,N_2020);
or U2055 (N_2055,N_2029,N_2008);
nand U2056 (N_2056,N_2001,N_2042);
and U2057 (N_2057,N_2023,N_2036);
or U2058 (N_2058,N_2045,N_2005);
nand U2059 (N_2059,N_2041,N_2006);
nand U2060 (N_2060,N_2022,N_2046);
nor U2061 (N_2061,N_2030,N_2013);
nor U2062 (N_2062,N_2039,N_2002);
or U2063 (N_2063,N_2026,N_2004);
nand U2064 (N_2064,N_2037,N_2031);
nand U2065 (N_2065,N_2021,N_2000);
and U2066 (N_2066,N_2040,N_2038);
or U2067 (N_2067,N_2014,N_2024);
nor U2068 (N_2068,N_2019,N_2010);
xor U2069 (N_2069,N_2043,N_2016);
or U2070 (N_2070,N_2028,N_2044);
or U2071 (N_2071,N_2047,N_2018);
or U2072 (N_2072,N_2011,N_2003);
nor U2073 (N_2073,N_2027,N_2035);
and U2074 (N_2074,N_2009,N_2007);
nand U2075 (N_2075,N_2032,N_2040);
nor U2076 (N_2076,N_2001,N_2004);
nor U2077 (N_2077,N_2010,N_2004);
or U2078 (N_2078,N_2030,N_2027);
and U2079 (N_2079,N_2009,N_2016);
and U2080 (N_2080,N_2002,N_2003);
nor U2081 (N_2081,N_2027,N_2007);
and U2082 (N_2082,N_2026,N_2010);
xor U2083 (N_2083,N_2035,N_2002);
or U2084 (N_2084,N_2009,N_2048);
nor U2085 (N_2085,N_2037,N_2025);
and U2086 (N_2086,N_2034,N_2021);
or U2087 (N_2087,N_2015,N_2025);
and U2088 (N_2088,N_2023,N_2024);
nor U2089 (N_2089,N_2013,N_2022);
or U2090 (N_2090,N_2039,N_2007);
nand U2091 (N_2091,N_2038,N_2024);
nand U2092 (N_2092,N_2000,N_2032);
nand U2093 (N_2093,N_2015,N_2023);
and U2094 (N_2094,N_2006,N_2049);
and U2095 (N_2095,N_2036,N_2049);
nor U2096 (N_2096,N_2016,N_2049);
or U2097 (N_2097,N_2041,N_2028);
and U2098 (N_2098,N_2011,N_2004);
nor U2099 (N_2099,N_2039,N_2013);
nand U2100 (N_2100,N_2070,N_2053);
nand U2101 (N_2101,N_2052,N_2073);
or U2102 (N_2102,N_2090,N_2074);
nor U2103 (N_2103,N_2050,N_2089);
nor U2104 (N_2104,N_2086,N_2096);
nor U2105 (N_2105,N_2092,N_2064);
nand U2106 (N_2106,N_2098,N_2083);
or U2107 (N_2107,N_2060,N_2059);
nand U2108 (N_2108,N_2063,N_2061);
and U2109 (N_2109,N_2065,N_2077);
nand U2110 (N_2110,N_2091,N_2068);
nand U2111 (N_2111,N_2056,N_2082);
and U2112 (N_2112,N_2067,N_2093);
nor U2113 (N_2113,N_2079,N_2076);
nand U2114 (N_2114,N_2075,N_2084);
xor U2115 (N_2115,N_2080,N_2087);
nand U2116 (N_2116,N_2078,N_2055);
nor U2117 (N_2117,N_2057,N_2054);
nor U2118 (N_2118,N_2097,N_2072);
nor U2119 (N_2119,N_2081,N_2069);
or U2120 (N_2120,N_2085,N_2066);
and U2121 (N_2121,N_2051,N_2088);
or U2122 (N_2122,N_2062,N_2099);
and U2123 (N_2123,N_2095,N_2058);
nand U2124 (N_2124,N_2071,N_2094);
nand U2125 (N_2125,N_2086,N_2067);
or U2126 (N_2126,N_2074,N_2097);
and U2127 (N_2127,N_2051,N_2073);
nor U2128 (N_2128,N_2070,N_2062);
xnor U2129 (N_2129,N_2054,N_2070);
or U2130 (N_2130,N_2072,N_2090);
nand U2131 (N_2131,N_2078,N_2083);
nor U2132 (N_2132,N_2066,N_2090);
and U2133 (N_2133,N_2060,N_2056);
or U2134 (N_2134,N_2093,N_2082);
or U2135 (N_2135,N_2062,N_2057);
nand U2136 (N_2136,N_2094,N_2096);
nand U2137 (N_2137,N_2079,N_2066);
or U2138 (N_2138,N_2081,N_2051);
and U2139 (N_2139,N_2092,N_2051);
nand U2140 (N_2140,N_2053,N_2097);
nor U2141 (N_2141,N_2068,N_2087);
or U2142 (N_2142,N_2091,N_2077);
nand U2143 (N_2143,N_2087,N_2093);
nor U2144 (N_2144,N_2053,N_2079);
or U2145 (N_2145,N_2054,N_2074);
xnor U2146 (N_2146,N_2062,N_2068);
or U2147 (N_2147,N_2085,N_2054);
or U2148 (N_2148,N_2055,N_2058);
and U2149 (N_2149,N_2076,N_2087);
or U2150 (N_2150,N_2128,N_2137);
and U2151 (N_2151,N_2132,N_2130);
nand U2152 (N_2152,N_2126,N_2142);
and U2153 (N_2153,N_2122,N_2139);
nor U2154 (N_2154,N_2104,N_2127);
or U2155 (N_2155,N_2120,N_2110);
nor U2156 (N_2156,N_2108,N_2109);
nor U2157 (N_2157,N_2145,N_2105);
nand U2158 (N_2158,N_2134,N_2144);
and U2159 (N_2159,N_2101,N_2138);
and U2160 (N_2160,N_2102,N_2100);
and U2161 (N_2161,N_2131,N_2124);
nor U2162 (N_2162,N_2123,N_2113);
nand U2163 (N_2163,N_2121,N_2103);
nor U2164 (N_2164,N_2129,N_2136);
nor U2165 (N_2165,N_2146,N_2125);
and U2166 (N_2166,N_2117,N_2141);
and U2167 (N_2167,N_2148,N_2111);
nand U2168 (N_2168,N_2119,N_2106);
nor U2169 (N_2169,N_2149,N_2114);
and U2170 (N_2170,N_2133,N_2118);
or U2171 (N_2171,N_2140,N_2107);
nand U2172 (N_2172,N_2116,N_2115);
or U2173 (N_2173,N_2135,N_2147);
nand U2174 (N_2174,N_2112,N_2143);
nor U2175 (N_2175,N_2110,N_2144);
nand U2176 (N_2176,N_2104,N_2103);
or U2177 (N_2177,N_2149,N_2146);
nand U2178 (N_2178,N_2144,N_2124);
nor U2179 (N_2179,N_2109,N_2146);
or U2180 (N_2180,N_2115,N_2143);
xor U2181 (N_2181,N_2143,N_2106);
or U2182 (N_2182,N_2117,N_2112);
nand U2183 (N_2183,N_2107,N_2118);
and U2184 (N_2184,N_2138,N_2111);
and U2185 (N_2185,N_2142,N_2123);
nor U2186 (N_2186,N_2146,N_2124);
nor U2187 (N_2187,N_2143,N_2124);
nor U2188 (N_2188,N_2139,N_2127);
nand U2189 (N_2189,N_2102,N_2143);
or U2190 (N_2190,N_2129,N_2139);
nand U2191 (N_2191,N_2125,N_2137);
nor U2192 (N_2192,N_2115,N_2108);
nor U2193 (N_2193,N_2106,N_2141);
and U2194 (N_2194,N_2110,N_2114);
and U2195 (N_2195,N_2140,N_2145);
or U2196 (N_2196,N_2149,N_2130);
nor U2197 (N_2197,N_2113,N_2145);
nor U2198 (N_2198,N_2131,N_2144);
nand U2199 (N_2199,N_2125,N_2105);
nor U2200 (N_2200,N_2153,N_2198);
nor U2201 (N_2201,N_2187,N_2186);
nor U2202 (N_2202,N_2164,N_2199);
nor U2203 (N_2203,N_2154,N_2179);
or U2204 (N_2204,N_2152,N_2174);
and U2205 (N_2205,N_2150,N_2160);
nand U2206 (N_2206,N_2196,N_2151);
nand U2207 (N_2207,N_2189,N_2184);
and U2208 (N_2208,N_2180,N_2163);
or U2209 (N_2209,N_2156,N_2157);
nand U2210 (N_2210,N_2168,N_2190);
and U2211 (N_2211,N_2194,N_2195);
nor U2212 (N_2212,N_2191,N_2181);
and U2213 (N_2213,N_2188,N_2175);
nor U2214 (N_2214,N_2170,N_2193);
nand U2215 (N_2215,N_2171,N_2172);
nor U2216 (N_2216,N_2173,N_2176);
and U2217 (N_2217,N_2159,N_2178);
or U2218 (N_2218,N_2161,N_2165);
nor U2219 (N_2219,N_2169,N_2183);
nand U2220 (N_2220,N_2155,N_2192);
nand U2221 (N_2221,N_2167,N_2158);
and U2222 (N_2222,N_2182,N_2185);
nor U2223 (N_2223,N_2162,N_2197);
and U2224 (N_2224,N_2166,N_2177);
or U2225 (N_2225,N_2179,N_2172);
nand U2226 (N_2226,N_2193,N_2177);
nor U2227 (N_2227,N_2159,N_2172);
and U2228 (N_2228,N_2153,N_2188);
nand U2229 (N_2229,N_2178,N_2164);
nand U2230 (N_2230,N_2167,N_2155);
and U2231 (N_2231,N_2198,N_2162);
nor U2232 (N_2232,N_2161,N_2196);
nand U2233 (N_2233,N_2161,N_2178);
or U2234 (N_2234,N_2168,N_2157);
nand U2235 (N_2235,N_2170,N_2190);
and U2236 (N_2236,N_2188,N_2156);
or U2237 (N_2237,N_2152,N_2171);
and U2238 (N_2238,N_2198,N_2194);
or U2239 (N_2239,N_2151,N_2154);
nor U2240 (N_2240,N_2184,N_2175);
nand U2241 (N_2241,N_2161,N_2170);
or U2242 (N_2242,N_2198,N_2151);
nor U2243 (N_2243,N_2192,N_2165);
and U2244 (N_2244,N_2176,N_2151);
nor U2245 (N_2245,N_2157,N_2195);
or U2246 (N_2246,N_2186,N_2199);
and U2247 (N_2247,N_2161,N_2174);
and U2248 (N_2248,N_2162,N_2173);
or U2249 (N_2249,N_2194,N_2185);
or U2250 (N_2250,N_2201,N_2231);
nor U2251 (N_2251,N_2205,N_2210);
or U2252 (N_2252,N_2226,N_2232);
nor U2253 (N_2253,N_2247,N_2238);
nor U2254 (N_2254,N_2204,N_2218);
and U2255 (N_2255,N_2223,N_2220);
and U2256 (N_2256,N_2230,N_2240);
or U2257 (N_2257,N_2228,N_2207);
and U2258 (N_2258,N_2221,N_2234);
nor U2259 (N_2259,N_2224,N_2244);
and U2260 (N_2260,N_2245,N_2206);
nand U2261 (N_2261,N_2242,N_2248);
or U2262 (N_2262,N_2249,N_2214);
nor U2263 (N_2263,N_2200,N_2222);
or U2264 (N_2264,N_2203,N_2217);
or U2265 (N_2265,N_2202,N_2227);
and U2266 (N_2266,N_2219,N_2239);
nor U2267 (N_2267,N_2225,N_2213);
or U2268 (N_2268,N_2212,N_2243);
nand U2269 (N_2269,N_2211,N_2246);
nand U2270 (N_2270,N_2208,N_2216);
nand U2271 (N_2271,N_2236,N_2235);
or U2272 (N_2272,N_2209,N_2233);
nor U2273 (N_2273,N_2241,N_2237);
xor U2274 (N_2274,N_2229,N_2215);
and U2275 (N_2275,N_2202,N_2245);
nand U2276 (N_2276,N_2217,N_2238);
nand U2277 (N_2277,N_2231,N_2237);
nand U2278 (N_2278,N_2203,N_2220);
nor U2279 (N_2279,N_2244,N_2248);
nor U2280 (N_2280,N_2210,N_2219);
and U2281 (N_2281,N_2228,N_2246);
or U2282 (N_2282,N_2239,N_2204);
nor U2283 (N_2283,N_2234,N_2207);
nor U2284 (N_2284,N_2235,N_2230);
nand U2285 (N_2285,N_2241,N_2232);
or U2286 (N_2286,N_2225,N_2228);
nor U2287 (N_2287,N_2234,N_2239);
nand U2288 (N_2288,N_2247,N_2241);
nand U2289 (N_2289,N_2207,N_2233);
nor U2290 (N_2290,N_2226,N_2209);
and U2291 (N_2291,N_2248,N_2246);
nor U2292 (N_2292,N_2238,N_2222);
nand U2293 (N_2293,N_2218,N_2217);
or U2294 (N_2294,N_2205,N_2222);
and U2295 (N_2295,N_2246,N_2218);
nand U2296 (N_2296,N_2246,N_2216);
nand U2297 (N_2297,N_2240,N_2200);
or U2298 (N_2298,N_2227,N_2218);
or U2299 (N_2299,N_2207,N_2201);
nor U2300 (N_2300,N_2287,N_2266);
nand U2301 (N_2301,N_2285,N_2286);
nand U2302 (N_2302,N_2282,N_2281);
or U2303 (N_2303,N_2297,N_2261);
nand U2304 (N_2304,N_2255,N_2295);
nand U2305 (N_2305,N_2283,N_2260);
or U2306 (N_2306,N_2262,N_2263);
nand U2307 (N_2307,N_2269,N_2253);
nor U2308 (N_2308,N_2256,N_2268);
and U2309 (N_2309,N_2277,N_2280);
nand U2310 (N_2310,N_2290,N_2288);
nand U2311 (N_2311,N_2267,N_2276);
and U2312 (N_2312,N_2271,N_2272);
or U2313 (N_2313,N_2252,N_2293);
nand U2314 (N_2314,N_2291,N_2257);
nand U2315 (N_2315,N_2251,N_2265);
nor U2316 (N_2316,N_2298,N_2289);
or U2317 (N_2317,N_2264,N_2273);
nor U2318 (N_2318,N_2274,N_2284);
or U2319 (N_2319,N_2254,N_2278);
nand U2320 (N_2320,N_2292,N_2299);
nor U2321 (N_2321,N_2258,N_2270);
nor U2322 (N_2322,N_2259,N_2275);
xor U2323 (N_2323,N_2250,N_2296);
nand U2324 (N_2324,N_2279,N_2294);
nor U2325 (N_2325,N_2295,N_2286);
and U2326 (N_2326,N_2256,N_2261);
nand U2327 (N_2327,N_2292,N_2262);
and U2328 (N_2328,N_2253,N_2251);
and U2329 (N_2329,N_2272,N_2286);
and U2330 (N_2330,N_2289,N_2252);
nand U2331 (N_2331,N_2270,N_2295);
and U2332 (N_2332,N_2275,N_2268);
nor U2333 (N_2333,N_2276,N_2263);
nand U2334 (N_2334,N_2267,N_2281);
and U2335 (N_2335,N_2297,N_2252);
and U2336 (N_2336,N_2259,N_2263);
nor U2337 (N_2337,N_2284,N_2297);
nor U2338 (N_2338,N_2263,N_2291);
nand U2339 (N_2339,N_2298,N_2285);
or U2340 (N_2340,N_2277,N_2275);
and U2341 (N_2341,N_2289,N_2257);
and U2342 (N_2342,N_2292,N_2259);
nor U2343 (N_2343,N_2297,N_2294);
xor U2344 (N_2344,N_2288,N_2284);
and U2345 (N_2345,N_2259,N_2284);
or U2346 (N_2346,N_2291,N_2269);
nor U2347 (N_2347,N_2282,N_2298);
nand U2348 (N_2348,N_2284,N_2260);
nand U2349 (N_2349,N_2276,N_2255);
or U2350 (N_2350,N_2344,N_2325);
or U2351 (N_2351,N_2346,N_2320);
nor U2352 (N_2352,N_2300,N_2335);
and U2353 (N_2353,N_2333,N_2309);
and U2354 (N_2354,N_2310,N_2305);
nand U2355 (N_2355,N_2339,N_2308);
xnor U2356 (N_2356,N_2304,N_2317);
nor U2357 (N_2357,N_2312,N_2340);
nor U2358 (N_2358,N_2348,N_2319);
and U2359 (N_2359,N_2311,N_2323);
and U2360 (N_2360,N_2338,N_2330);
or U2361 (N_2361,N_2327,N_2318);
nor U2362 (N_2362,N_2343,N_2345);
nor U2363 (N_2363,N_2336,N_2332);
nand U2364 (N_2364,N_2307,N_2331);
and U2365 (N_2365,N_2303,N_2316);
nor U2366 (N_2366,N_2334,N_2302);
or U2367 (N_2367,N_2321,N_2313);
and U2368 (N_2368,N_2328,N_2349);
or U2369 (N_2369,N_2306,N_2324);
nor U2370 (N_2370,N_2314,N_2329);
and U2371 (N_2371,N_2341,N_2301);
or U2372 (N_2372,N_2326,N_2315);
and U2373 (N_2373,N_2322,N_2347);
nor U2374 (N_2374,N_2342,N_2337);
and U2375 (N_2375,N_2328,N_2346);
or U2376 (N_2376,N_2324,N_2345);
nand U2377 (N_2377,N_2308,N_2310);
or U2378 (N_2378,N_2312,N_2313);
nand U2379 (N_2379,N_2347,N_2340);
and U2380 (N_2380,N_2331,N_2311);
nor U2381 (N_2381,N_2319,N_2337);
nand U2382 (N_2382,N_2342,N_2339);
or U2383 (N_2383,N_2337,N_2335);
nor U2384 (N_2384,N_2341,N_2335);
nand U2385 (N_2385,N_2309,N_2307);
or U2386 (N_2386,N_2338,N_2333);
and U2387 (N_2387,N_2333,N_2317);
nand U2388 (N_2388,N_2309,N_2322);
nor U2389 (N_2389,N_2349,N_2314);
nor U2390 (N_2390,N_2322,N_2307);
nand U2391 (N_2391,N_2307,N_2339);
or U2392 (N_2392,N_2307,N_2315);
nand U2393 (N_2393,N_2334,N_2339);
nand U2394 (N_2394,N_2321,N_2326);
or U2395 (N_2395,N_2338,N_2305);
nor U2396 (N_2396,N_2330,N_2318);
or U2397 (N_2397,N_2332,N_2305);
nor U2398 (N_2398,N_2302,N_2305);
or U2399 (N_2399,N_2315,N_2300);
nand U2400 (N_2400,N_2382,N_2364);
or U2401 (N_2401,N_2390,N_2368);
and U2402 (N_2402,N_2356,N_2393);
xnor U2403 (N_2403,N_2354,N_2383);
and U2404 (N_2404,N_2358,N_2353);
nor U2405 (N_2405,N_2360,N_2372);
or U2406 (N_2406,N_2381,N_2395);
and U2407 (N_2407,N_2369,N_2376);
nand U2408 (N_2408,N_2367,N_2365);
nor U2409 (N_2409,N_2361,N_2380);
or U2410 (N_2410,N_2392,N_2384);
nand U2411 (N_2411,N_2394,N_2386);
or U2412 (N_2412,N_2397,N_2375);
and U2413 (N_2413,N_2378,N_2389);
xor U2414 (N_2414,N_2396,N_2391);
or U2415 (N_2415,N_2350,N_2370);
or U2416 (N_2416,N_2377,N_2398);
nor U2417 (N_2417,N_2399,N_2355);
or U2418 (N_2418,N_2359,N_2357);
or U2419 (N_2419,N_2352,N_2388);
or U2420 (N_2420,N_2385,N_2363);
nor U2421 (N_2421,N_2373,N_2371);
nor U2422 (N_2422,N_2366,N_2362);
or U2423 (N_2423,N_2374,N_2379);
nand U2424 (N_2424,N_2351,N_2387);
nand U2425 (N_2425,N_2380,N_2399);
nor U2426 (N_2426,N_2373,N_2395);
nand U2427 (N_2427,N_2350,N_2376);
or U2428 (N_2428,N_2359,N_2371);
nor U2429 (N_2429,N_2396,N_2376);
nand U2430 (N_2430,N_2399,N_2381);
or U2431 (N_2431,N_2385,N_2374);
nand U2432 (N_2432,N_2396,N_2353);
nand U2433 (N_2433,N_2395,N_2363);
nor U2434 (N_2434,N_2394,N_2397);
nand U2435 (N_2435,N_2368,N_2367);
nor U2436 (N_2436,N_2394,N_2371);
nand U2437 (N_2437,N_2365,N_2357);
and U2438 (N_2438,N_2374,N_2390);
nand U2439 (N_2439,N_2371,N_2372);
and U2440 (N_2440,N_2355,N_2394);
or U2441 (N_2441,N_2387,N_2366);
nor U2442 (N_2442,N_2356,N_2365);
or U2443 (N_2443,N_2394,N_2380);
nor U2444 (N_2444,N_2350,N_2375);
and U2445 (N_2445,N_2380,N_2381);
and U2446 (N_2446,N_2358,N_2371);
or U2447 (N_2447,N_2395,N_2353);
nor U2448 (N_2448,N_2375,N_2383);
nand U2449 (N_2449,N_2352,N_2353);
nand U2450 (N_2450,N_2422,N_2408);
and U2451 (N_2451,N_2441,N_2417);
nand U2452 (N_2452,N_2400,N_2433);
or U2453 (N_2453,N_2410,N_2424);
and U2454 (N_2454,N_2445,N_2446);
and U2455 (N_2455,N_2429,N_2412);
and U2456 (N_2456,N_2418,N_2448);
and U2457 (N_2457,N_2423,N_2416);
nor U2458 (N_2458,N_2413,N_2406);
and U2459 (N_2459,N_2442,N_2440);
and U2460 (N_2460,N_2405,N_2425);
and U2461 (N_2461,N_2407,N_2403);
nand U2462 (N_2462,N_2427,N_2404);
nand U2463 (N_2463,N_2438,N_2447);
and U2464 (N_2464,N_2434,N_2437);
nor U2465 (N_2465,N_2402,N_2430);
and U2466 (N_2466,N_2401,N_2414);
or U2467 (N_2467,N_2415,N_2421);
nor U2468 (N_2468,N_2449,N_2439);
nand U2469 (N_2469,N_2426,N_2435);
xor U2470 (N_2470,N_2443,N_2431);
nor U2471 (N_2471,N_2419,N_2444);
or U2472 (N_2472,N_2420,N_2432);
nand U2473 (N_2473,N_2436,N_2409);
and U2474 (N_2474,N_2411,N_2428);
nand U2475 (N_2475,N_2447,N_2422);
or U2476 (N_2476,N_2417,N_2430);
and U2477 (N_2477,N_2401,N_2413);
and U2478 (N_2478,N_2447,N_2409);
or U2479 (N_2479,N_2444,N_2447);
or U2480 (N_2480,N_2432,N_2417);
or U2481 (N_2481,N_2422,N_2433);
and U2482 (N_2482,N_2444,N_2435);
nand U2483 (N_2483,N_2423,N_2441);
nor U2484 (N_2484,N_2441,N_2433);
nor U2485 (N_2485,N_2446,N_2436);
or U2486 (N_2486,N_2424,N_2407);
or U2487 (N_2487,N_2410,N_2430);
xor U2488 (N_2488,N_2404,N_2419);
and U2489 (N_2489,N_2414,N_2448);
nor U2490 (N_2490,N_2436,N_2434);
nand U2491 (N_2491,N_2444,N_2413);
or U2492 (N_2492,N_2422,N_2434);
nand U2493 (N_2493,N_2440,N_2427);
nand U2494 (N_2494,N_2433,N_2415);
or U2495 (N_2495,N_2415,N_2441);
and U2496 (N_2496,N_2426,N_2449);
nor U2497 (N_2497,N_2424,N_2409);
and U2498 (N_2498,N_2428,N_2425);
or U2499 (N_2499,N_2438,N_2412);
xor U2500 (N_2500,N_2466,N_2498);
nand U2501 (N_2501,N_2472,N_2461);
nor U2502 (N_2502,N_2473,N_2471);
nand U2503 (N_2503,N_2487,N_2483);
nand U2504 (N_2504,N_2459,N_2492);
nand U2505 (N_2505,N_2494,N_2495);
nand U2506 (N_2506,N_2490,N_2460);
or U2507 (N_2507,N_2479,N_2480);
nand U2508 (N_2508,N_2465,N_2488);
and U2509 (N_2509,N_2453,N_2481);
nand U2510 (N_2510,N_2474,N_2462);
nand U2511 (N_2511,N_2486,N_2477);
and U2512 (N_2512,N_2470,N_2496);
nor U2513 (N_2513,N_2491,N_2458);
or U2514 (N_2514,N_2478,N_2463);
and U2515 (N_2515,N_2468,N_2476);
or U2516 (N_2516,N_2469,N_2454);
and U2517 (N_2517,N_2497,N_2464);
nand U2518 (N_2518,N_2456,N_2489);
nor U2519 (N_2519,N_2467,N_2499);
nand U2520 (N_2520,N_2484,N_2457);
and U2521 (N_2521,N_2455,N_2493);
xor U2522 (N_2522,N_2452,N_2485);
or U2523 (N_2523,N_2450,N_2482);
or U2524 (N_2524,N_2475,N_2451);
or U2525 (N_2525,N_2452,N_2494);
and U2526 (N_2526,N_2484,N_2456);
nand U2527 (N_2527,N_2495,N_2488);
or U2528 (N_2528,N_2455,N_2474);
or U2529 (N_2529,N_2466,N_2456);
or U2530 (N_2530,N_2475,N_2472);
or U2531 (N_2531,N_2481,N_2499);
or U2532 (N_2532,N_2489,N_2491);
and U2533 (N_2533,N_2489,N_2494);
or U2534 (N_2534,N_2452,N_2476);
and U2535 (N_2535,N_2464,N_2463);
or U2536 (N_2536,N_2466,N_2486);
or U2537 (N_2537,N_2461,N_2477);
or U2538 (N_2538,N_2458,N_2475);
nand U2539 (N_2539,N_2491,N_2493);
and U2540 (N_2540,N_2455,N_2452);
or U2541 (N_2541,N_2458,N_2463);
nand U2542 (N_2542,N_2469,N_2470);
xnor U2543 (N_2543,N_2460,N_2469);
and U2544 (N_2544,N_2466,N_2459);
or U2545 (N_2545,N_2451,N_2480);
nor U2546 (N_2546,N_2479,N_2492);
nor U2547 (N_2547,N_2488,N_2486);
nand U2548 (N_2548,N_2496,N_2478);
and U2549 (N_2549,N_2468,N_2451);
or U2550 (N_2550,N_2511,N_2522);
and U2551 (N_2551,N_2527,N_2514);
nor U2552 (N_2552,N_2540,N_2521);
and U2553 (N_2553,N_2518,N_2523);
and U2554 (N_2554,N_2535,N_2547);
or U2555 (N_2555,N_2543,N_2529);
or U2556 (N_2556,N_2525,N_2526);
nand U2557 (N_2557,N_2509,N_2504);
nor U2558 (N_2558,N_2542,N_2545);
and U2559 (N_2559,N_2531,N_2532);
nand U2560 (N_2560,N_2506,N_2541);
nand U2561 (N_2561,N_2537,N_2517);
or U2562 (N_2562,N_2546,N_2502);
nor U2563 (N_2563,N_2500,N_2510);
nand U2564 (N_2564,N_2508,N_2536);
or U2565 (N_2565,N_2524,N_2505);
and U2566 (N_2566,N_2548,N_2533);
xor U2567 (N_2567,N_2539,N_2530);
and U2568 (N_2568,N_2528,N_2512);
nor U2569 (N_2569,N_2538,N_2544);
or U2570 (N_2570,N_2534,N_2515);
nor U2571 (N_2571,N_2520,N_2513);
nand U2572 (N_2572,N_2516,N_2507);
nor U2573 (N_2573,N_2501,N_2503);
nand U2574 (N_2574,N_2549,N_2519);
nor U2575 (N_2575,N_2528,N_2503);
nand U2576 (N_2576,N_2509,N_2513);
and U2577 (N_2577,N_2541,N_2522);
nand U2578 (N_2578,N_2527,N_2510);
and U2579 (N_2579,N_2519,N_2509);
nand U2580 (N_2580,N_2502,N_2520);
nor U2581 (N_2581,N_2531,N_2543);
nor U2582 (N_2582,N_2507,N_2520);
and U2583 (N_2583,N_2523,N_2522);
nand U2584 (N_2584,N_2547,N_2507);
xnor U2585 (N_2585,N_2505,N_2521);
or U2586 (N_2586,N_2536,N_2507);
nor U2587 (N_2587,N_2540,N_2507);
and U2588 (N_2588,N_2549,N_2532);
and U2589 (N_2589,N_2520,N_2534);
and U2590 (N_2590,N_2513,N_2524);
nor U2591 (N_2591,N_2518,N_2527);
nand U2592 (N_2592,N_2549,N_2536);
or U2593 (N_2593,N_2505,N_2529);
or U2594 (N_2594,N_2526,N_2548);
nor U2595 (N_2595,N_2524,N_2523);
nand U2596 (N_2596,N_2513,N_2516);
or U2597 (N_2597,N_2522,N_2535);
or U2598 (N_2598,N_2516,N_2521);
nor U2599 (N_2599,N_2549,N_2516);
or U2600 (N_2600,N_2569,N_2592);
and U2601 (N_2601,N_2561,N_2572);
or U2602 (N_2602,N_2593,N_2553);
or U2603 (N_2603,N_2590,N_2564);
and U2604 (N_2604,N_2579,N_2556);
xnor U2605 (N_2605,N_2557,N_2588);
nand U2606 (N_2606,N_2570,N_2552);
nor U2607 (N_2607,N_2574,N_2575);
nand U2608 (N_2608,N_2566,N_2550);
or U2609 (N_2609,N_2578,N_2597);
and U2610 (N_2610,N_2551,N_2596);
nand U2611 (N_2611,N_2586,N_2563);
or U2612 (N_2612,N_2585,N_2595);
and U2613 (N_2613,N_2587,N_2599);
nand U2614 (N_2614,N_2571,N_2568);
nand U2615 (N_2615,N_2573,N_2594);
nand U2616 (N_2616,N_2555,N_2567);
and U2617 (N_2617,N_2560,N_2580);
nand U2618 (N_2618,N_2558,N_2584);
and U2619 (N_2619,N_2562,N_2559);
nor U2620 (N_2620,N_2581,N_2591);
nand U2621 (N_2621,N_2582,N_2589);
nand U2622 (N_2622,N_2598,N_2554);
nand U2623 (N_2623,N_2565,N_2576);
or U2624 (N_2624,N_2577,N_2583);
nand U2625 (N_2625,N_2568,N_2577);
nand U2626 (N_2626,N_2580,N_2581);
or U2627 (N_2627,N_2592,N_2551);
nor U2628 (N_2628,N_2584,N_2559);
and U2629 (N_2629,N_2579,N_2561);
nor U2630 (N_2630,N_2596,N_2583);
or U2631 (N_2631,N_2580,N_2554);
and U2632 (N_2632,N_2554,N_2596);
nor U2633 (N_2633,N_2551,N_2574);
or U2634 (N_2634,N_2585,N_2581);
xor U2635 (N_2635,N_2594,N_2563);
and U2636 (N_2636,N_2594,N_2568);
nand U2637 (N_2637,N_2588,N_2560);
and U2638 (N_2638,N_2558,N_2588);
or U2639 (N_2639,N_2574,N_2555);
and U2640 (N_2640,N_2580,N_2599);
or U2641 (N_2641,N_2568,N_2574);
or U2642 (N_2642,N_2587,N_2589);
nor U2643 (N_2643,N_2576,N_2585);
and U2644 (N_2644,N_2560,N_2581);
nor U2645 (N_2645,N_2571,N_2585);
and U2646 (N_2646,N_2556,N_2582);
and U2647 (N_2647,N_2571,N_2575);
nor U2648 (N_2648,N_2579,N_2593);
or U2649 (N_2649,N_2550,N_2597);
nand U2650 (N_2650,N_2638,N_2611);
nand U2651 (N_2651,N_2630,N_2604);
xnor U2652 (N_2652,N_2614,N_2618);
or U2653 (N_2653,N_2602,N_2648);
or U2654 (N_2654,N_2616,N_2649);
nor U2655 (N_2655,N_2647,N_2627);
or U2656 (N_2656,N_2606,N_2629);
or U2657 (N_2657,N_2615,N_2642);
and U2658 (N_2658,N_2644,N_2619);
nand U2659 (N_2659,N_2622,N_2605);
nand U2660 (N_2660,N_2628,N_2645);
nor U2661 (N_2661,N_2610,N_2613);
nand U2662 (N_2662,N_2612,N_2631);
nor U2663 (N_2663,N_2624,N_2633);
or U2664 (N_2664,N_2639,N_2617);
nand U2665 (N_2665,N_2621,N_2646);
nor U2666 (N_2666,N_2632,N_2636);
nand U2667 (N_2667,N_2609,N_2635);
nand U2668 (N_2668,N_2623,N_2626);
nand U2669 (N_2669,N_2640,N_2608);
and U2670 (N_2670,N_2625,N_2603);
and U2671 (N_2671,N_2620,N_2600);
and U2672 (N_2672,N_2607,N_2637);
and U2673 (N_2673,N_2643,N_2641);
nand U2674 (N_2674,N_2634,N_2601);
or U2675 (N_2675,N_2623,N_2611);
or U2676 (N_2676,N_2612,N_2611);
and U2677 (N_2677,N_2637,N_2613);
nand U2678 (N_2678,N_2636,N_2635);
or U2679 (N_2679,N_2637,N_2642);
or U2680 (N_2680,N_2604,N_2603);
and U2681 (N_2681,N_2626,N_2607);
nor U2682 (N_2682,N_2645,N_2600);
nor U2683 (N_2683,N_2628,N_2615);
nor U2684 (N_2684,N_2633,N_2635);
nand U2685 (N_2685,N_2612,N_2632);
nor U2686 (N_2686,N_2622,N_2637);
or U2687 (N_2687,N_2641,N_2614);
nor U2688 (N_2688,N_2626,N_2619);
nand U2689 (N_2689,N_2643,N_2631);
or U2690 (N_2690,N_2621,N_2619);
and U2691 (N_2691,N_2620,N_2630);
or U2692 (N_2692,N_2634,N_2614);
nand U2693 (N_2693,N_2623,N_2639);
nand U2694 (N_2694,N_2604,N_2627);
nand U2695 (N_2695,N_2640,N_2625);
nand U2696 (N_2696,N_2622,N_2601);
and U2697 (N_2697,N_2644,N_2623);
xnor U2698 (N_2698,N_2611,N_2643);
or U2699 (N_2699,N_2618,N_2624);
nand U2700 (N_2700,N_2689,N_2678);
or U2701 (N_2701,N_2659,N_2680);
and U2702 (N_2702,N_2679,N_2676);
and U2703 (N_2703,N_2681,N_2699);
nand U2704 (N_2704,N_2661,N_2654);
and U2705 (N_2705,N_2677,N_2682);
nand U2706 (N_2706,N_2669,N_2657);
or U2707 (N_2707,N_2686,N_2663);
nand U2708 (N_2708,N_2653,N_2696);
nand U2709 (N_2709,N_2660,N_2674);
or U2710 (N_2710,N_2662,N_2668);
nand U2711 (N_2711,N_2675,N_2697);
nand U2712 (N_2712,N_2673,N_2664);
nand U2713 (N_2713,N_2684,N_2693);
nand U2714 (N_2714,N_2687,N_2698);
nor U2715 (N_2715,N_2650,N_2658);
or U2716 (N_2716,N_2670,N_2672);
or U2717 (N_2717,N_2655,N_2665);
nand U2718 (N_2718,N_2671,N_2691);
nor U2719 (N_2719,N_2690,N_2694);
nor U2720 (N_2720,N_2656,N_2666);
or U2721 (N_2721,N_2695,N_2651);
or U2722 (N_2722,N_2683,N_2692);
nor U2723 (N_2723,N_2652,N_2667);
nor U2724 (N_2724,N_2688,N_2685);
or U2725 (N_2725,N_2653,N_2694);
nand U2726 (N_2726,N_2652,N_2671);
nand U2727 (N_2727,N_2681,N_2658);
or U2728 (N_2728,N_2651,N_2672);
nand U2729 (N_2729,N_2683,N_2688);
and U2730 (N_2730,N_2657,N_2688);
and U2731 (N_2731,N_2691,N_2682);
or U2732 (N_2732,N_2669,N_2688);
nand U2733 (N_2733,N_2674,N_2692);
nor U2734 (N_2734,N_2661,N_2663);
or U2735 (N_2735,N_2667,N_2658);
nor U2736 (N_2736,N_2650,N_2661);
nand U2737 (N_2737,N_2677,N_2691);
or U2738 (N_2738,N_2652,N_2656);
nor U2739 (N_2739,N_2661,N_2668);
or U2740 (N_2740,N_2656,N_2657);
nor U2741 (N_2741,N_2690,N_2673);
or U2742 (N_2742,N_2691,N_2659);
and U2743 (N_2743,N_2655,N_2689);
nor U2744 (N_2744,N_2681,N_2675);
nor U2745 (N_2745,N_2682,N_2689);
or U2746 (N_2746,N_2676,N_2684);
or U2747 (N_2747,N_2676,N_2696);
and U2748 (N_2748,N_2674,N_2683);
and U2749 (N_2749,N_2670,N_2659);
or U2750 (N_2750,N_2723,N_2739);
nand U2751 (N_2751,N_2706,N_2724);
or U2752 (N_2752,N_2741,N_2701);
or U2753 (N_2753,N_2743,N_2744);
nor U2754 (N_2754,N_2709,N_2703);
or U2755 (N_2755,N_2748,N_2712);
nor U2756 (N_2756,N_2715,N_2738);
nand U2757 (N_2757,N_2730,N_2726);
nor U2758 (N_2758,N_2725,N_2708);
nor U2759 (N_2759,N_2721,N_2731);
nand U2760 (N_2760,N_2710,N_2702);
nand U2761 (N_2761,N_2713,N_2736);
or U2762 (N_2762,N_2742,N_2727);
nand U2763 (N_2763,N_2737,N_2745);
and U2764 (N_2764,N_2749,N_2720);
or U2765 (N_2765,N_2734,N_2704);
nand U2766 (N_2766,N_2728,N_2732);
and U2767 (N_2767,N_2729,N_2700);
and U2768 (N_2768,N_2714,N_2717);
nand U2769 (N_2769,N_2707,N_2705);
nand U2770 (N_2770,N_2746,N_2722);
and U2771 (N_2771,N_2735,N_2711);
nand U2772 (N_2772,N_2718,N_2747);
nor U2773 (N_2773,N_2719,N_2733);
nor U2774 (N_2774,N_2740,N_2716);
nor U2775 (N_2775,N_2736,N_2708);
or U2776 (N_2776,N_2719,N_2744);
nor U2777 (N_2777,N_2708,N_2740);
or U2778 (N_2778,N_2740,N_2710);
nand U2779 (N_2779,N_2725,N_2735);
or U2780 (N_2780,N_2730,N_2706);
nand U2781 (N_2781,N_2721,N_2718);
nand U2782 (N_2782,N_2713,N_2745);
nand U2783 (N_2783,N_2705,N_2721);
nor U2784 (N_2784,N_2705,N_2749);
and U2785 (N_2785,N_2748,N_2716);
nor U2786 (N_2786,N_2716,N_2714);
nand U2787 (N_2787,N_2747,N_2729);
nor U2788 (N_2788,N_2703,N_2721);
nand U2789 (N_2789,N_2727,N_2714);
or U2790 (N_2790,N_2737,N_2701);
or U2791 (N_2791,N_2712,N_2709);
nor U2792 (N_2792,N_2748,N_2729);
and U2793 (N_2793,N_2749,N_2728);
or U2794 (N_2794,N_2724,N_2738);
or U2795 (N_2795,N_2733,N_2738);
and U2796 (N_2796,N_2748,N_2705);
and U2797 (N_2797,N_2718,N_2734);
nand U2798 (N_2798,N_2749,N_2702);
or U2799 (N_2799,N_2724,N_2735);
nor U2800 (N_2800,N_2766,N_2762);
or U2801 (N_2801,N_2780,N_2788);
or U2802 (N_2802,N_2774,N_2775);
or U2803 (N_2803,N_2760,N_2795);
and U2804 (N_2804,N_2776,N_2756);
or U2805 (N_2805,N_2781,N_2798);
nand U2806 (N_2806,N_2772,N_2789);
or U2807 (N_2807,N_2761,N_2791);
or U2808 (N_2808,N_2771,N_2770);
and U2809 (N_2809,N_2773,N_2790);
or U2810 (N_2810,N_2784,N_2782);
and U2811 (N_2811,N_2786,N_2765);
xor U2812 (N_2812,N_2750,N_2757);
nor U2813 (N_2813,N_2796,N_2752);
and U2814 (N_2814,N_2783,N_2769);
nand U2815 (N_2815,N_2755,N_2753);
nor U2816 (N_2816,N_2767,N_2797);
nor U2817 (N_2817,N_2793,N_2792);
xnor U2818 (N_2818,N_2785,N_2787);
nand U2819 (N_2819,N_2759,N_2764);
and U2820 (N_2820,N_2777,N_2754);
or U2821 (N_2821,N_2751,N_2768);
and U2822 (N_2822,N_2779,N_2794);
and U2823 (N_2823,N_2799,N_2758);
nand U2824 (N_2824,N_2778,N_2763);
nor U2825 (N_2825,N_2769,N_2763);
and U2826 (N_2826,N_2766,N_2778);
nand U2827 (N_2827,N_2761,N_2768);
nand U2828 (N_2828,N_2767,N_2776);
nand U2829 (N_2829,N_2781,N_2771);
or U2830 (N_2830,N_2793,N_2774);
nor U2831 (N_2831,N_2780,N_2771);
nand U2832 (N_2832,N_2767,N_2758);
and U2833 (N_2833,N_2780,N_2753);
nor U2834 (N_2834,N_2759,N_2783);
nor U2835 (N_2835,N_2778,N_2761);
and U2836 (N_2836,N_2758,N_2790);
and U2837 (N_2837,N_2768,N_2753);
or U2838 (N_2838,N_2796,N_2769);
nor U2839 (N_2839,N_2780,N_2765);
nand U2840 (N_2840,N_2789,N_2752);
nor U2841 (N_2841,N_2798,N_2757);
or U2842 (N_2842,N_2794,N_2793);
nand U2843 (N_2843,N_2768,N_2788);
nand U2844 (N_2844,N_2769,N_2798);
and U2845 (N_2845,N_2783,N_2786);
or U2846 (N_2846,N_2792,N_2755);
nand U2847 (N_2847,N_2755,N_2777);
nand U2848 (N_2848,N_2770,N_2772);
nand U2849 (N_2849,N_2791,N_2763);
and U2850 (N_2850,N_2805,N_2821);
and U2851 (N_2851,N_2815,N_2814);
or U2852 (N_2852,N_2838,N_2845);
nand U2853 (N_2853,N_2802,N_2808);
nand U2854 (N_2854,N_2836,N_2810);
and U2855 (N_2855,N_2834,N_2848);
nor U2856 (N_2856,N_2811,N_2846);
and U2857 (N_2857,N_2804,N_2822);
nor U2858 (N_2858,N_2803,N_2849);
or U2859 (N_2859,N_2823,N_2807);
and U2860 (N_2860,N_2817,N_2813);
or U2861 (N_2861,N_2841,N_2833);
nand U2862 (N_2862,N_2827,N_2809);
nor U2863 (N_2863,N_2844,N_2840);
nand U2864 (N_2864,N_2835,N_2832);
nand U2865 (N_2865,N_2825,N_2816);
nor U2866 (N_2866,N_2837,N_2812);
nor U2867 (N_2867,N_2847,N_2819);
and U2868 (N_2868,N_2831,N_2826);
nor U2869 (N_2869,N_2824,N_2820);
or U2870 (N_2870,N_2842,N_2843);
xnor U2871 (N_2871,N_2801,N_2818);
nand U2872 (N_2872,N_2828,N_2806);
and U2873 (N_2873,N_2830,N_2829);
nor U2874 (N_2874,N_2839,N_2800);
and U2875 (N_2875,N_2842,N_2829);
or U2876 (N_2876,N_2837,N_2845);
or U2877 (N_2877,N_2807,N_2811);
or U2878 (N_2878,N_2831,N_2807);
or U2879 (N_2879,N_2831,N_2840);
or U2880 (N_2880,N_2847,N_2811);
nor U2881 (N_2881,N_2821,N_2810);
nor U2882 (N_2882,N_2834,N_2846);
and U2883 (N_2883,N_2820,N_2830);
and U2884 (N_2884,N_2806,N_2829);
or U2885 (N_2885,N_2811,N_2827);
nor U2886 (N_2886,N_2803,N_2836);
or U2887 (N_2887,N_2849,N_2824);
or U2888 (N_2888,N_2834,N_2828);
xor U2889 (N_2889,N_2843,N_2804);
or U2890 (N_2890,N_2826,N_2846);
or U2891 (N_2891,N_2809,N_2843);
and U2892 (N_2892,N_2812,N_2825);
nand U2893 (N_2893,N_2806,N_2800);
xnor U2894 (N_2894,N_2827,N_2830);
xnor U2895 (N_2895,N_2809,N_2841);
nand U2896 (N_2896,N_2814,N_2809);
nand U2897 (N_2897,N_2810,N_2841);
nand U2898 (N_2898,N_2805,N_2810);
or U2899 (N_2899,N_2813,N_2811);
or U2900 (N_2900,N_2879,N_2884);
and U2901 (N_2901,N_2883,N_2889);
and U2902 (N_2902,N_2861,N_2874);
nand U2903 (N_2903,N_2851,N_2856);
nor U2904 (N_2904,N_2887,N_2872);
nand U2905 (N_2905,N_2896,N_2885);
and U2906 (N_2906,N_2870,N_2873);
nand U2907 (N_2907,N_2881,N_2871);
nand U2908 (N_2908,N_2897,N_2868);
nand U2909 (N_2909,N_2880,N_2888);
nor U2910 (N_2910,N_2855,N_2899);
or U2911 (N_2911,N_2886,N_2863);
nand U2912 (N_2912,N_2866,N_2898);
nor U2913 (N_2913,N_2894,N_2893);
nand U2914 (N_2914,N_2858,N_2865);
and U2915 (N_2915,N_2895,N_2867);
or U2916 (N_2916,N_2852,N_2882);
nor U2917 (N_2917,N_2878,N_2854);
nand U2918 (N_2918,N_2869,N_2860);
xnor U2919 (N_2919,N_2857,N_2892);
nor U2920 (N_2920,N_2891,N_2850);
or U2921 (N_2921,N_2890,N_2876);
nor U2922 (N_2922,N_2864,N_2859);
or U2923 (N_2923,N_2875,N_2862);
nor U2924 (N_2924,N_2877,N_2853);
or U2925 (N_2925,N_2864,N_2853);
or U2926 (N_2926,N_2896,N_2863);
nand U2927 (N_2927,N_2892,N_2854);
or U2928 (N_2928,N_2858,N_2854);
nor U2929 (N_2929,N_2884,N_2882);
or U2930 (N_2930,N_2887,N_2875);
or U2931 (N_2931,N_2884,N_2861);
nor U2932 (N_2932,N_2888,N_2877);
nor U2933 (N_2933,N_2860,N_2886);
and U2934 (N_2934,N_2883,N_2891);
xor U2935 (N_2935,N_2889,N_2862);
and U2936 (N_2936,N_2876,N_2873);
and U2937 (N_2937,N_2871,N_2878);
nor U2938 (N_2938,N_2898,N_2860);
nand U2939 (N_2939,N_2887,N_2879);
xor U2940 (N_2940,N_2898,N_2870);
nand U2941 (N_2941,N_2869,N_2850);
nand U2942 (N_2942,N_2865,N_2883);
and U2943 (N_2943,N_2877,N_2894);
xor U2944 (N_2944,N_2880,N_2859);
nand U2945 (N_2945,N_2865,N_2895);
or U2946 (N_2946,N_2879,N_2855);
nand U2947 (N_2947,N_2858,N_2851);
nor U2948 (N_2948,N_2893,N_2879);
and U2949 (N_2949,N_2878,N_2870);
and U2950 (N_2950,N_2938,N_2911);
or U2951 (N_2951,N_2905,N_2947);
or U2952 (N_2952,N_2913,N_2918);
nor U2953 (N_2953,N_2904,N_2940);
nand U2954 (N_2954,N_2931,N_2903);
nor U2955 (N_2955,N_2917,N_2927);
nand U2956 (N_2956,N_2926,N_2937);
xnor U2957 (N_2957,N_2934,N_2902);
nand U2958 (N_2958,N_2909,N_2949);
and U2959 (N_2959,N_2936,N_2906);
nand U2960 (N_2960,N_2943,N_2942);
or U2961 (N_2961,N_2908,N_2919);
and U2962 (N_2962,N_2916,N_2932);
and U2963 (N_2963,N_2925,N_2921);
nor U2964 (N_2964,N_2920,N_2933);
nand U2965 (N_2965,N_2941,N_2900);
nor U2966 (N_2966,N_2946,N_2923);
nand U2967 (N_2967,N_2929,N_2901);
and U2968 (N_2968,N_2945,N_2922);
nand U2969 (N_2969,N_2910,N_2930);
nor U2970 (N_2970,N_2928,N_2935);
nand U2971 (N_2971,N_2924,N_2944);
nand U2972 (N_2972,N_2915,N_2948);
nor U2973 (N_2973,N_2912,N_2939);
or U2974 (N_2974,N_2907,N_2914);
nor U2975 (N_2975,N_2920,N_2932);
nand U2976 (N_2976,N_2920,N_2946);
nor U2977 (N_2977,N_2945,N_2949);
nand U2978 (N_2978,N_2921,N_2902);
and U2979 (N_2979,N_2919,N_2924);
nand U2980 (N_2980,N_2905,N_2919);
nand U2981 (N_2981,N_2943,N_2918);
and U2982 (N_2982,N_2933,N_2949);
or U2983 (N_2983,N_2912,N_2946);
nand U2984 (N_2984,N_2945,N_2948);
nor U2985 (N_2985,N_2936,N_2924);
xor U2986 (N_2986,N_2944,N_2904);
nand U2987 (N_2987,N_2905,N_2949);
nand U2988 (N_2988,N_2920,N_2934);
nor U2989 (N_2989,N_2937,N_2944);
and U2990 (N_2990,N_2932,N_2902);
nand U2991 (N_2991,N_2920,N_2913);
or U2992 (N_2992,N_2945,N_2947);
nor U2993 (N_2993,N_2940,N_2921);
nand U2994 (N_2994,N_2912,N_2928);
and U2995 (N_2995,N_2915,N_2949);
nor U2996 (N_2996,N_2917,N_2915);
or U2997 (N_2997,N_2938,N_2933);
nor U2998 (N_2998,N_2904,N_2902);
nand U2999 (N_2999,N_2905,N_2912);
nor UO_0 (O_0,N_2996,N_2970);
xnor UO_1 (O_1,N_2987,N_2990);
nor UO_2 (O_2,N_2989,N_2961);
or UO_3 (O_3,N_2980,N_2995);
and UO_4 (O_4,N_2953,N_2975);
nand UO_5 (O_5,N_2967,N_2963);
and UO_6 (O_6,N_2977,N_2992);
nand UO_7 (O_7,N_2973,N_2968);
nand UO_8 (O_8,N_2982,N_2960);
nand UO_9 (O_9,N_2957,N_2969);
nor UO_10 (O_10,N_2986,N_2962);
or UO_11 (O_11,N_2978,N_2979);
or UO_12 (O_12,N_2966,N_2972);
and UO_13 (O_13,N_2991,N_2954);
or UO_14 (O_14,N_2955,N_2964);
or UO_15 (O_15,N_2993,N_2965);
nand UO_16 (O_16,N_2999,N_2981);
and UO_17 (O_17,N_2983,N_2997);
and UO_18 (O_18,N_2952,N_2951);
and UO_19 (O_19,N_2984,N_2958);
and UO_20 (O_20,N_2994,N_2956);
and UO_21 (O_21,N_2998,N_2976);
xor UO_22 (O_22,N_2959,N_2985);
nand UO_23 (O_23,N_2974,N_2950);
nor UO_24 (O_24,N_2988,N_2971);
nor UO_25 (O_25,N_2988,N_2953);
nor UO_26 (O_26,N_2997,N_2994);
nor UO_27 (O_27,N_2981,N_2966);
and UO_28 (O_28,N_2986,N_2957);
nand UO_29 (O_29,N_2981,N_2970);
or UO_30 (O_30,N_2950,N_2962);
nand UO_31 (O_31,N_2964,N_2954);
or UO_32 (O_32,N_2993,N_2983);
nor UO_33 (O_33,N_2964,N_2992);
and UO_34 (O_34,N_2984,N_2987);
nor UO_35 (O_35,N_2976,N_2956);
nor UO_36 (O_36,N_2986,N_2987);
nand UO_37 (O_37,N_2950,N_2984);
xnor UO_38 (O_38,N_2968,N_2976);
xnor UO_39 (O_39,N_2985,N_2960);
and UO_40 (O_40,N_2994,N_2999);
and UO_41 (O_41,N_2967,N_2974);
or UO_42 (O_42,N_2970,N_2957);
nor UO_43 (O_43,N_2983,N_2964);
nand UO_44 (O_44,N_2957,N_2971);
and UO_45 (O_45,N_2998,N_2951);
or UO_46 (O_46,N_2967,N_2997);
and UO_47 (O_47,N_2954,N_2980);
nand UO_48 (O_48,N_2953,N_2991);
nand UO_49 (O_49,N_2953,N_2999);
or UO_50 (O_50,N_2964,N_2993);
or UO_51 (O_51,N_2983,N_2960);
and UO_52 (O_52,N_2984,N_2971);
nor UO_53 (O_53,N_2979,N_2971);
nand UO_54 (O_54,N_2986,N_2966);
and UO_55 (O_55,N_2989,N_2974);
nand UO_56 (O_56,N_2979,N_2969);
or UO_57 (O_57,N_2974,N_2992);
nand UO_58 (O_58,N_2989,N_2994);
and UO_59 (O_59,N_2969,N_2999);
or UO_60 (O_60,N_2982,N_2970);
or UO_61 (O_61,N_2997,N_2992);
nand UO_62 (O_62,N_2952,N_2990);
and UO_63 (O_63,N_2999,N_2973);
and UO_64 (O_64,N_2972,N_2987);
nand UO_65 (O_65,N_2973,N_2978);
or UO_66 (O_66,N_2951,N_2969);
or UO_67 (O_67,N_2982,N_2983);
or UO_68 (O_68,N_2996,N_2973);
or UO_69 (O_69,N_2973,N_2951);
and UO_70 (O_70,N_2957,N_2989);
nor UO_71 (O_71,N_2956,N_2993);
or UO_72 (O_72,N_2970,N_2955);
nand UO_73 (O_73,N_2972,N_2992);
nor UO_74 (O_74,N_2975,N_2980);
nand UO_75 (O_75,N_2964,N_2995);
or UO_76 (O_76,N_2971,N_2990);
nand UO_77 (O_77,N_2982,N_2998);
nor UO_78 (O_78,N_2976,N_2975);
or UO_79 (O_79,N_2994,N_2968);
nand UO_80 (O_80,N_2954,N_2966);
and UO_81 (O_81,N_2981,N_2964);
and UO_82 (O_82,N_2994,N_2950);
and UO_83 (O_83,N_2988,N_2959);
nor UO_84 (O_84,N_2974,N_2976);
nand UO_85 (O_85,N_2970,N_2989);
and UO_86 (O_86,N_2963,N_2990);
or UO_87 (O_87,N_2990,N_2989);
and UO_88 (O_88,N_2950,N_2973);
or UO_89 (O_89,N_2997,N_2987);
nand UO_90 (O_90,N_2990,N_2972);
and UO_91 (O_91,N_2990,N_2974);
or UO_92 (O_92,N_2959,N_2993);
nor UO_93 (O_93,N_2957,N_2975);
and UO_94 (O_94,N_2950,N_2963);
nor UO_95 (O_95,N_2977,N_2975);
and UO_96 (O_96,N_2979,N_2957);
nor UO_97 (O_97,N_2999,N_2979);
and UO_98 (O_98,N_2977,N_2962);
nor UO_99 (O_99,N_2964,N_2972);
nand UO_100 (O_100,N_2957,N_2966);
nor UO_101 (O_101,N_2955,N_2967);
and UO_102 (O_102,N_2983,N_2985);
nand UO_103 (O_103,N_2990,N_2977);
nor UO_104 (O_104,N_2973,N_2991);
and UO_105 (O_105,N_2984,N_2983);
nand UO_106 (O_106,N_2957,N_2964);
nand UO_107 (O_107,N_2991,N_2965);
and UO_108 (O_108,N_2967,N_2999);
or UO_109 (O_109,N_2952,N_2986);
nor UO_110 (O_110,N_2965,N_2961);
or UO_111 (O_111,N_2967,N_2994);
nor UO_112 (O_112,N_2976,N_2971);
and UO_113 (O_113,N_2954,N_2975);
or UO_114 (O_114,N_2982,N_2987);
and UO_115 (O_115,N_2961,N_2990);
and UO_116 (O_116,N_2955,N_2957);
nand UO_117 (O_117,N_2953,N_2961);
nor UO_118 (O_118,N_2969,N_2997);
nor UO_119 (O_119,N_2993,N_2950);
or UO_120 (O_120,N_2988,N_2963);
or UO_121 (O_121,N_2958,N_2950);
or UO_122 (O_122,N_2982,N_2986);
nand UO_123 (O_123,N_2956,N_2974);
and UO_124 (O_124,N_2995,N_2984);
or UO_125 (O_125,N_2968,N_2983);
nor UO_126 (O_126,N_2961,N_2972);
nor UO_127 (O_127,N_2992,N_2961);
and UO_128 (O_128,N_2997,N_2962);
and UO_129 (O_129,N_2951,N_2971);
nand UO_130 (O_130,N_2966,N_2984);
xnor UO_131 (O_131,N_2968,N_2986);
nand UO_132 (O_132,N_2958,N_2957);
and UO_133 (O_133,N_2959,N_2994);
nor UO_134 (O_134,N_2970,N_2950);
or UO_135 (O_135,N_2986,N_2974);
xor UO_136 (O_136,N_2958,N_2966);
nand UO_137 (O_137,N_2963,N_2972);
nand UO_138 (O_138,N_2981,N_2951);
or UO_139 (O_139,N_2966,N_2977);
nand UO_140 (O_140,N_2980,N_2983);
nor UO_141 (O_141,N_2990,N_2975);
nand UO_142 (O_142,N_2978,N_2990);
nor UO_143 (O_143,N_2994,N_2965);
and UO_144 (O_144,N_2958,N_2963);
and UO_145 (O_145,N_2993,N_2979);
and UO_146 (O_146,N_2956,N_2979);
nor UO_147 (O_147,N_2966,N_2988);
nand UO_148 (O_148,N_2969,N_2985);
or UO_149 (O_149,N_2951,N_2950);
or UO_150 (O_150,N_2995,N_2965);
nand UO_151 (O_151,N_2985,N_2972);
or UO_152 (O_152,N_2969,N_2970);
nor UO_153 (O_153,N_2953,N_2964);
nand UO_154 (O_154,N_2954,N_2985);
or UO_155 (O_155,N_2963,N_2979);
and UO_156 (O_156,N_2960,N_2993);
and UO_157 (O_157,N_2985,N_2978);
nor UO_158 (O_158,N_2981,N_2958);
or UO_159 (O_159,N_2999,N_2954);
or UO_160 (O_160,N_2973,N_2993);
nand UO_161 (O_161,N_2954,N_2988);
and UO_162 (O_162,N_2999,N_2992);
and UO_163 (O_163,N_2998,N_2987);
nor UO_164 (O_164,N_2961,N_2956);
or UO_165 (O_165,N_2971,N_2962);
nand UO_166 (O_166,N_2960,N_2965);
or UO_167 (O_167,N_2958,N_2968);
and UO_168 (O_168,N_2997,N_2973);
nand UO_169 (O_169,N_2973,N_2953);
or UO_170 (O_170,N_2950,N_2985);
nor UO_171 (O_171,N_2980,N_2968);
nand UO_172 (O_172,N_2981,N_2954);
or UO_173 (O_173,N_2967,N_2984);
nand UO_174 (O_174,N_2958,N_2952);
or UO_175 (O_175,N_2983,N_2998);
and UO_176 (O_176,N_2952,N_2992);
or UO_177 (O_177,N_2998,N_2977);
and UO_178 (O_178,N_2951,N_2978);
and UO_179 (O_179,N_2983,N_2999);
nand UO_180 (O_180,N_2994,N_2953);
nor UO_181 (O_181,N_2953,N_2968);
nor UO_182 (O_182,N_2990,N_2969);
and UO_183 (O_183,N_2983,N_2965);
or UO_184 (O_184,N_2950,N_2981);
xor UO_185 (O_185,N_2958,N_2971);
or UO_186 (O_186,N_2997,N_2968);
and UO_187 (O_187,N_2993,N_2995);
nand UO_188 (O_188,N_2986,N_2979);
nand UO_189 (O_189,N_2966,N_2976);
and UO_190 (O_190,N_2991,N_2989);
nor UO_191 (O_191,N_2988,N_2980);
nand UO_192 (O_192,N_2952,N_2968);
nor UO_193 (O_193,N_2997,N_2990);
and UO_194 (O_194,N_2950,N_2980);
and UO_195 (O_195,N_2983,N_2995);
nor UO_196 (O_196,N_2967,N_2979);
nor UO_197 (O_197,N_2958,N_2979);
nor UO_198 (O_198,N_2960,N_2956);
nand UO_199 (O_199,N_2959,N_2996);
and UO_200 (O_200,N_2957,N_2990);
and UO_201 (O_201,N_2986,N_2969);
and UO_202 (O_202,N_2953,N_2990);
or UO_203 (O_203,N_2987,N_2989);
nor UO_204 (O_204,N_2968,N_2950);
or UO_205 (O_205,N_2962,N_2954);
and UO_206 (O_206,N_2953,N_2987);
nor UO_207 (O_207,N_2963,N_2968);
or UO_208 (O_208,N_2951,N_2987);
nor UO_209 (O_209,N_2986,N_2983);
nor UO_210 (O_210,N_2999,N_2989);
nand UO_211 (O_211,N_2952,N_2993);
nand UO_212 (O_212,N_2976,N_2959);
and UO_213 (O_213,N_2956,N_2982);
nor UO_214 (O_214,N_2953,N_2986);
and UO_215 (O_215,N_2961,N_2950);
nand UO_216 (O_216,N_2956,N_2990);
or UO_217 (O_217,N_2971,N_2977);
nand UO_218 (O_218,N_2971,N_2972);
nor UO_219 (O_219,N_2976,N_2991);
xnor UO_220 (O_220,N_2958,N_2989);
nand UO_221 (O_221,N_2960,N_2991);
nor UO_222 (O_222,N_2999,N_2978);
nor UO_223 (O_223,N_2983,N_2978);
nor UO_224 (O_224,N_2958,N_2973);
nor UO_225 (O_225,N_2988,N_2997);
nand UO_226 (O_226,N_2960,N_2999);
nor UO_227 (O_227,N_2976,N_2989);
nand UO_228 (O_228,N_2992,N_2958);
xor UO_229 (O_229,N_2996,N_2954);
nor UO_230 (O_230,N_2984,N_2973);
nand UO_231 (O_231,N_2955,N_2980);
nand UO_232 (O_232,N_2957,N_2973);
and UO_233 (O_233,N_2995,N_2961);
and UO_234 (O_234,N_2965,N_2985);
or UO_235 (O_235,N_2974,N_2994);
nand UO_236 (O_236,N_2989,N_2979);
or UO_237 (O_237,N_2962,N_2996);
and UO_238 (O_238,N_2951,N_2989);
and UO_239 (O_239,N_2973,N_2987);
or UO_240 (O_240,N_2974,N_2964);
nor UO_241 (O_241,N_2956,N_2973);
and UO_242 (O_242,N_2953,N_2972);
and UO_243 (O_243,N_2961,N_2960);
and UO_244 (O_244,N_2967,N_2989);
or UO_245 (O_245,N_2990,N_2954);
nand UO_246 (O_246,N_2993,N_2996);
nor UO_247 (O_247,N_2982,N_2952);
and UO_248 (O_248,N_2967,N_2980);
nand UO_249 (O_249,N_2986,N_2965);
or UO_250 (O_250,N_2970,N_2994);
nand UO_251 (O_251,N_2995,N_2955);
nor UO_252 (O_252,N_2992,N_2962);
and UO_253 (O_253,N_2960,N_2974);
nor UO_254 (O_254,N_2976,N_2962);
nor UO_255 (O_255,N_2993,N_2992);
or UO_256 (O_256,N_2989,N_2954);
or UO_257 (O_257,N_2997,N_2980);
or UO_258 (O_258,N_2955,N_2992);
or UO_259 (O_259,N_2964,N_2996);
nand UO_260 (O_260,N_2961,N_2993);
or UO_261 (O_261,N_2995,N_2981);
or UO_262 (O_262,N_2956,N_2983);
nand UO_263 (O_263,N_2995,N_2971);
nor UO_264 (O_264,N_2967,N_2993);
or UO_265 (O_265,N_2997,N_2999);
xnor UO_266 (O_266,N_2989,N_2975);
or UO_267 (O_267,N_2958,N_2982);
or UO_268 (O_268,N_2971,N_2975);
nor UO_269 (O_269,N_2996,N_2998);
nand UO_270 (O_270,N_2977,N_2964);
or UO_271 (O_271,N_2979,N_2997);
nor UO_272 (O_272,N_2959,N_2980);
nand UO_273 (O_273,N_2980,N_2970);
and UO_274 (O_274,N_2959,N_2951);
nand UO_275 (O_275,N_2971,N_2974);
nand UO_276 (O_276,N_2984,N_2990);
nor UO_277 (O_277,N_2954,N_2950);
and UO_278 (O_278,N_2982,N_2991);
and UO_279 (O_279,N_2967,N_2962);
nor UO_280 (O_280,N_2968,N_2977);
nand UO_281 (O_281,N_2988,N_2978);
and UO_282 (O_282,N_2957,N_2954);
xnor UO_283 (O_283,N_2993,N_2953);
and UO_284 (O_284,N_2982,N_2996);
and UO_285 (O_285,N_2951,N_2985);
and UO_286 (O_286,N_2964,N_2990);
nor UO_287 (O_287,N_2984,N_2975);
nor UO_288 (O_288,N_2951,N_2977);
nor UO_289 (O_289,N_2986,N_2998);
nor UO_290 (O_290,N_2964,N_2994);
nor UO_291 (O_291,N_2988,N_2987);
nor UO_292 (O_292,N_2970,N_2958);
nand UO_293 (O_293,N_2981,N_2979);
xor UO_294 (O_294,N_2969,N_2976);
and UO_295 (O_295,N_2958,N_2964);
nand UO_296 (O_296,N_2965,N_2992);
xnor UO_297 (O_297,N_2993,N_2970);
or UO_298 (O_298,N_2965,N_2973);
nor UO_299 (O_299,N_2966,N_2951);
and UO_300 (O_300,N_2971,N_2993);
and UO_301 (O_301,N_2999,N_2985);
nor UO_302 (O_302,N_2991,N_2950);
nand UO_303 (O_303,N_2984,N_2980);
nor UO_304 (O_304,N_2964,N_2960);
nand UO_305 (O_305,N_2998,N_2954);
or UO_306 (O_306,N_2988,N_2970);
and UO_307 (O_307,N_2983,N_2972);
nand UO_308 (O_308,N_2954,N_2958);
nand UO_309 (O_309,N_2983,N_2951);
nor UO_310 (O_310,N_2983,N_2958);
nand UO_311 (O_311,N_2955,N_2971);
and UO_312 (O_312,N_2968,N_2991);
nor UO_313 (O_313,N_2965,N_2987);
nor UO_314 (O_314,N_2960,N_2989);
or UO_315 (O_315,N_2994,N_2987);
nand UO_316 (O_316,N_2988,N_2990);
and UO_317 (O_317,N_2967,N_2977);
and UO_318 (O_318,N_2981,N_2992);
and UO_319 (O_319,N_2976,N_2963);
and UO_320 (O_320,N_2981,N_2953);
or UO_321 (O_321,N_2994,N_2972);
xor UO_322 (O_322,N_2981,N_2977);
and UO_323 (O_323,N_2988,N_2972);
or UO_324 (O_324,N_2957,N_2963);
nand UO_325 (O_325,N_2972,N_2958);
and UO_326 (O_326,N_2986,N_2992);
nor UO_327 (O_327,N_2988,N_2952);
or UO_328 (O_328,N_2979,N_2994);
and UO_329 (O_329,N_2985,N_2995);
nor UO_330 (O_330,N_2976,N_2961);
nand UO_331 (O_331,N_2967,N_2995);
or UO_332 (O_332,N_2959,N_2961);
nand UO_333 (O_333,N_2984,N_2955);
and UO_334 (O_334,N_2958,N_2959);
nor UO_335 (O_335,N_2966,N_2973);
nand UO_336 (O_336,N_2950,N_2999);
and UO_337 (O_337,N_2975,N_2960);
nand UO_338 (O_338,N_2982,N_2985);
and UO_339 (O_339,N_2999,N_2971);
and UO_340 (O_340,N_2953,N_2956);
nand UO_341 (O_341,N_2966,N_2990);
nor UO_342 (O_342,N_2968,N_2993);
nor UO_343 (O_343,N_2970,N_2960);
or UO_344 (O_344,N_2969,N_2981);
nand UO_345 (O_345,N_2956,N_2996);
and UO_346 (O_346,N_2968,N_2966);
nor UO_347 (O_347,N_2997,N_2986);
nand UO_348 (O_348,N_2951,N_2954);
nor UO_349 (O_349,N_2968,N_2955);
and UO_350 (O_350,N_2968,N_2992);
and UO_351 (O_351,N_2960,N_2954);
nor UO_352 (O_352,N_2952,N_2964);
nor UO_353 (O_353,N_2970,N_2974);
nand UO_354 (O_354,N_2976,N_2983);
and UO_355 (O_355,N_2975,N_2956);
nor UO_356 (O_356,N_2997,N_2952);
and UO_357 (O_357,N_2977,N_2953);
or UO_358 (O_358,N_2998,N_2961);
nand UO_359 (O_359,N_2951,N_2994);
or UO_360 (O_360,N_2968,N_2995);
or UO_361 (O_361,N_2959,N_2990);
nor UO_362 (O_362,N_2955,N_2958);
nand UO_363 (O_363,N_2958,N_2991);
nand UO_364 (O_364,N_2979,N_2982);
nand UO_365 (O_365,N_2986,N_2960);
nand UO_366 (O_366,N_2956,N_2999);
nor UO_367 (O_367,N_2999,N_2955);
or UO_368 (O_368,N_2969,N_2950);
nand UO_369 (O_369,N_2979,N_2972);
xor UO_370 (O_370,N_2967,N_2953);
nor UO_371 (O_371,N_2996,N_2967);
and UO_372 (O_372,N_2978,N_2991);
and UO_373 (O_373,N_2953,N_2959);
nor UO_374 (O_374,N_2991,N_2967);
and UO_375 (O_375,N_2983,N_2981);
nor UO_376 (O_376,N_2970,N_2985);
nand UO_377 (O_377,N_2968,N_2972);
and UO_378 (O_378,N_2971,N_2980);
and UO_379 (O_379,N_2975,N_2988);
nor UO_380 (O_380,N_2951,N_2992);
nor UO_381 (O_381,N_2973,N_2961);
nand UO_382 (O_382,N_2990,N_2992);
nor UO_383 (O_383,N_2998,N_2973);
or UO_384 (O_384,N_2985,N_2957);
or UO_385 (O_385,N_2969,N_2961);
nand UO_386 (O_386,N_2979,N_2959);
and UO_387 (O_387,N_2967,N_2951);
or UO_388 (O_388,N_2958,N_2987);
or UO_389 (O_389,N_2967,N_2987);
and UO_390 (O_390,N_2966,N_2967);
and UO_391 (O_391,N_2964,N_2979);
and UO_392 (O_392,N_2976,N_2980);
and UO_393 (O_393,N_2953,N_2989);
nand UO_394 (O_394,N_2998,N_2978);
and UO_395 (O_395,N_2985,N_2964);
or UO_396 (O_396,N_2953,N_2992);
or UO_397 (O_397,N_2981,N_2956);
or UO_398 (O_398,N_2961,N_2997);
and UO_399 (O_399,N_2989,N_2950);
and UO_400 (O_400,N_2992,N_2989);
or UO_401 (O_401,N_2953,N_2963);
or UO_402 (O_402,N_2970,N_2997);
and UO_403 (O_403,N_2992,N_2988);
and UO_404 (O_404,N_2978,N_2982);
nor UO_405 (O_405,N_2978,N_2960);
nand UO_406 (O_406,N_2974,N_2977);
nand UO_407 (O_407,N_2970,N_2998);
or UO_408 (O_408,N_2982,N_2995);
nor UO_409 (O_409,N_2964,N_2989);
xor UO_410 (O_410,N_2953,N_2985);
nor UO_411 (O_411,N_2969,N_2977);
and UO_412 (O_412,N_2958,N_2988);
or UO_413 (O_413,N_2951,N_2958);
and UO_414 (O_414,N_2963,N_2951);
nor UO_415 (O_415,N_2956,N_2965);
or UO_416 (O_416,N_2966,N_2994);
or UO_417 (O_417,N_2973,N_2980);
nor UO_418 (O_418,N_2995,N_2979);
and UO_419 (O_419,N_2978,N_2955);
or UO_420 (O_420,N_2965,N_2980);
or UO_421 (O_421,N_2987,N_2960);
nor UO_422 (O_422,N_2991,N_2955);
nand UO_423 (O_423,N_2957,N_2993);
and UO_424 (O_424,N_2990,N_2950);
and UO_425 (O_425,N_2973,N_2992);
nor UO_426 (O_426,N_2986,N_2988);
and UO_427 (O_427,N_2979,N_2973);
or UO_428 (O_428,N_2999,N_2965);
and UO_429 (O_429,N_2985,N_2981);
nor UO_430 (O_430,N_2952,N_2950);
and UO_431 (O_431,N_2957,N_2961);
and UO_432 (O_432,N_2992,N_2976);
and UO_433 (O_433,N_2951,N_2997);
nand UO_434 (O_434,N_2995,N_2956);
or UO_435 (O_435,N_2959,N_2966);
and UO_436 (O_436,N_2990,N_2980);
or UO_437 (O_437,N_2967,N_2969);
nor UO_438 (O_438,N_2956,N_2985);
or UO_439 (O_439,N_2968,N_2999);
nand UO_440 (O_440,N_2976,N_2965);
nor UO_441 (O_441,N_2962,N_2984);
nand UO_442 (O_442,N_2991,N_2951);
and UO_443 (O_443,N_2985,N_2961);
or UO_444 (O_444,N_2979,N_2966);
or UO_445 (O_445,N_2971,N_2997);
xor UO_446 (O_446,N_2987,N_2950);
and UO_447 (O_447,N_2954,N_2986);
and UO_448 (O_448,N_2982,N_2954);
or UO_449 (O_449,N_2959,N_2997);
and UO_450 (O_450,N_2975,N_2983);
or UO_451 (O_451,N_2981,N_2987);
or UO_452 (O_452,N_2998,N_2990);
or UO_453 (O_453,N_2994,N_2977);
nand UO_454 (O_454,N_2970,N_2963);
and UO_455 (O_455,N_2964,N_2998);
or UO_456 (O_456,N_2981,N_2978);
nor UO_457 (O_457,N_2972,N_2954);
xnor UO_458 (O_458,N_2957,N_2999);
xor UO_459 (O_459,N_2967,N_2959);
or UO_460 (O_460,N_2984,N_2978);
nand UO_461 (O_461,N_2959,N_2971);
nor UO_462 (O_462,N_2974,N_2959);
or UO_463 (O_463,N_2989,N_2978);
or UO_464 (O_464,N_2986,N_2975);
and UO_465 (O_465,N_2970,N_2973);
nor UO_466 (O_466,N_2957,N_2962);
and UO_467 (O_467,N_2981,N_2974);
or UO_468 (O_468,N_2983,N_2990);
nand UO_469 (O_469,N_2988,N_2951);
and UO_470 (O_470,N_2960,N_2994);
nor UO_471 (O_471,N_2965,N_2988);
nor UO_472 (O_472,N_2980,N_2991);
nor UO_473 (O_473,N_2968,N_2990);
nand UO_474 (O_474,N_2984,N_2961);
nand UO_475 (O_475,N_2991,N_2969);
and UO_476 (O_476,N_2974,N_2988);
nor UO_477 (O_477,N_2997,N_2989);
and UO_478 (O_478,N_2993,N_2981);
and UO_479 (O_479,N_2953,N_2983);
and UO_480 (O_480,N_2953,N_2998);
nor UO_481 (O_481,N_2983,N_2977);
and UO_482 (O_482,N_2995,N_2973);
or UO_483 (O_483,N_2970,N_2967);
nor UO_484 (O_484,N_2984,N_2969);
or UO_485 (O_485,N_2963,N_2980);
nand UO_486 (O_486,N_2969,N_2958);
nor UO_487 (O_487,N_2989,N_2982);
and UO_488 (O_488,N_2998,N_2994);
nor UO_489 (O_489,N_2957,N_2974);
and UO_490 (O_490,N_2991,N_2959);
nor UO_491 (O_491,N_2996,N_2963);
or UO_492 (O_492,N_2973,N_2964);
and UO_493 (O_493,N_2953,N_2969);
and UO_494 (O_494,N_2981,N_2955);
nor UO_495 (O_495,N_2995,N_2986);
or UO_496 (O_496,N_2966,N_2974);
and UO_497 (O_497,N_2955,N_2954);
or UO_498 (O_498,N_2994,N_2978);
or UO_499 (O_499,N_2972,N_2974);
endmodule