module basic_500_3000_500_3_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_80,In_70);
and U1 (N_1,In_287,In_175);
and U2 (N_2,In_190,In_346);
nand U3 (N_3,In_363,In_253);
or U4 (N_4,In_197,In_294);
or U5 (N_5,In_440,In_411);
nand U6 (N_6,In_238,In_121);
nand U7 (N_7,In_176,In_482);
xor U8 (N_8,In_257,In_173);
or U9 (N_9,In_282,In_304);
xnor U10 (N_10,In_14,In_200);
or U11 (N_11,In_340,In_165);
nand U12 (N_12,In_481,In_405);
and U13 (N_13,In_447,In_279);
and U14 (N_14,In_320,In_296);
nand U15 (N_15,In_149,In_353);
xnor U16 (N_16,In_209,In_168);
and U17 (N_17,In_196,In_21);
nor U18 (N_18,In_409,In_63);
and U19 (N_19,In_206,In_295);
nor U20 (N_20,In_124,In_475);
and U21 (N_21,In_116,In_383);
or U22 (N_22,In_221,In_241);
or U23 (N_23,In_78,In_369);
or U24 (N_24,In_130,In_162);
nand U25 (N_25,In_289,In_329);
and U26 (N_26,In_177,In_372);
or U27 (N_27,In_260,In_429);
or U28 (N_28,In_64,In_258);
nor U29 (N_29,In_91,In_399);
and U30 (N_30,In_113,In_108);
and U31 (N_31,In_179,In_127);
and U32 (N_32,In_486,In_152);
nand U33 (N_33,In_213,In_438);
nand U34 (N_34,In_48,In_254);
nor U35 (N_35,In_459,In_73);
and U36 (N_36,In_55,In_1);
and U37 (N_37,In_193,In_249);
and U38 (N_38,In_366,In_473);
nand U39 (N_39,In_499,In_211);
xnor U40 (N_40,In_231,In_111);
and U41 (N_41,In_334,In_265);
nor U42 (N_42,In_240,In_34);
and U43 (N_43,In_266,In_134);
xor U44 (N_44,In_164,In_288);
or U45 (N_45,In_463,In_129);
nor U46 (N_46,In_110,In_285);
nand U47 (N_47,In_36,In_6);
or U48 (N_48,In_376,In_275);
nand U49 (N_49,In_7,In_77);
nand U50 (N_50,In_368,In_344);
and U51 (N_51,In_442,In_458);
and U52 (N_52,In_432,In_226);
nor U53 (N_53,In_484,In_439);
or U54 (N_54,In_72,In_410);
nand U55 (N_55,In_428,In_83);
nor U56 (N_56,In_443,In_256);
or U57 (N_57,In_359,In_341);
nor U58 (N_58,In_131,In_43);
or U59 (N_59,In_89,In_232);
nand U60 (N_60,In_23,In_395);
nand U61 (N_61,In_315,In_454);
and U62 (N_62,In_74,In_180);
nand U63 (N_63,In_337,In_332);
or U64 (N_64,In_472,In_184);
nor U65 (N_65,In_158,In_269);
nand U66 (N_66,In_106,In_93);
nand U67 (N_67,In_479,In_5);
nor U68 (N_68,In_434,In_189);
or U69 (N_69,In_140,In_328);
nor U70 (N_70,In_161,In_65);
or U71 (N_71,In_272,In_319);
nor U72 (N_72,In_485,In_22);
nand U73 (N_73,In_316,In_147);
or U74 (N_74,In_468,In_351);
or U75 (N_75,In_114,In_495);
nand U76 (N_76,In_321,In_387);
or U77 (N_77,In_248,In_471);
nand U78 (N_78,In_59,In_457);
nor U79 (N_79,In_26,In_31);
nor U80 (N_80,In_138,In_339);
and U81 (N_81,In_284,In_452);
or U82 (N_82,In_393,In_18);
and U83 (N_83,In_342,In_28);
nor U84 (N_84,In_268,In_33);
nor U85 (N_85,In_390,In_40);
nand U86 (N_86,In_470,In_414);
nor U87 (N_87,In_400,In_107);
nand U88 (N_88,In_16,In_476);
nand U89 (N_89,In_293,In_263);
and U90 (N_90,In_49,In_132);
nor U91 (N_91,In_174,In_223);
nand U92 (N_92,In_195,In_437);
nor U93 (N_93,In_301,In_178);
nor U94 (N_94,In_318,In_183);
nand U95 (N_95,In_228,In_385);
or U96 (N_96,In_51,In_493);
or U97 (N_97,In_283,In_92);
nor U98 (N_98,In_84,In_311);
and U99 (N_99,In_386,In_455);
or U100 (N_100,In_436,In_102);
nand U101 (N_101,In_126,In_456);
and U102 (N_102,In_298,In_233);
nor U103 (N_103,In_487,In_291);
nor U104 (N_104,In_103,In_322);
or U105 (N_105,In_188,In_67);
xnor U106 (N_106,In_276,In_66);
or U107 (N_107,In_413,In_199);
nor U108 (N_108,In_474,In_202);
and U109 (N_109,In_317,In_261);
nor U110 (N_110,In_203,In_309);
nor U111 (N_111,In_378,In_365);
nand U112 (N_112,In_3,In_109);
nand U113 (N_113,In_392,In_303);
or U114 (N_114,In_186,In_97);
xor U115 (N_115,In_2,In_277);
nor U116 (N_116,In_379,In_490);
xor U117 (N_117,In_305,In_45);
nor U118 (N_118,In_345,In_251);
nor U119 (N_119,In_388,In_4);
or U120 (N_120,In_208,In_201);
nand U121 (N_121,In_204,In_156);
nor U122 (N_122,In_128,In_46);
or U123 (N_123,In_497,In_99);
nor U124 (N_124,In_194,In_56);
and U125 (N_125,In_370,In_151);
nand U126 (N_126,In_354,In_42);
nor U127 (N_127,In_219,In_225);
or U128 (N_128,In_270,In_467);
or U129 (N_129,In_403,In_54);
nand U130 (N_130,In_215,In_492);
nand U131 (N_131,In_469,In_465);
and U132 (N_132,In_153,In_397);
nor U133 (N_133,In_53,In_19);
or U134 (N_134,In_185,In_35);
nor U135 (N_135,In_182,In_71);
or U136 (N_136,In_216,In_299);
nand U137 (N_137,In_314,In_466);
nand U138 (N_138,In_212,In_445);
nor U139 (N_139,In_488,In_462);
xnor U140 (N_140,In_133,In_308);
and U141 (N_141,In_252,In_426);
nand U142 (N_142,In_352,In_460);
nand U143 (N_143,In_112,In_86);
nand U144 (N_144,In_20,In_355);
nand U145 (N_145,In_449,In_313);
or U146 (N_146,In_243,In_494);
nand U147 (N_147,In_123,In_154);
and U148 (N_148,In_356,In_47);
nand U149 (N_149,In_214,In_453);
nand U150 (N_150,In_229,In_273);
nor U151 (N_151,In_491,In_159);
nor U152 (N_152,In_430,In_331);
and U153 (N_153,In_100,In_198);
nand U154 (N_154,In_171,In_38);
or U155 (N_155,In_274,In_167);
nand U156 (N_156,In_404,In_62);
or U157 (N_157,In_82,In_419);
nor U158 (N_158,In_325,In_30);
or U159 (N_159,In_478,In_420);
nand U160 (N_160,In_135,In_323);
xnor U161 (N_161,In_187,In_330);
nor U162 (N_162,In_95,In_297);
nand U163 (N_163,In_68,In_278);
and U164 (N_164,In_17,In_75);
nand U165 (N_165,In_343,In_286);
nand U166 (N_166,In_144,In_160);
or U167 (N_167,In_12,In_448);
nor U168 (N_168,In_224,In_181);
nor U169 (N_169,In_217,In_431);
and U170 (N_170,In_119,In_60);
or U171 (N_171,In_267,In_362);
and U172 (N_172,In_326,In_358);
nand U173 (N_173,In_408,In_192);
or U174 (N_174,In_451,In_24);
or U175 (N_175,In_25,In_307);
nand U176 (N_176,In_324,In_242);
nand U177 (N_177,In_424,In_489);
nand U178 (N_178,In_496,In_139);
nor U179 (N_179,In_327,In_338);
nor U180 (N_180,In_402,In_247);
xnor U181 (N_181,In_239,In_381);
or U182 (N_182,In_44,In_371);
and U183 (N_183,In_446,In_235);
nor U184 (N_184,In_172,In_333);
and U185 (N_185,In_88,In_349);
or U186 (N_186,In_382,In_39);
nor U187 (N_187,In_394,In_373);
nor U188 (N_188,In_58,In_170);
and U189 (N_189,In_104,In_364);
nand U190 (N_190,In_375,In_94);
xnor U191 (N_191,In_335,In_136);
or U192 (N_192,In_57,In_234);
and U193 (N_193,In_336,In_205);
or U194 (N_194,In_464,In_96);
or U195 (N_195,In_27,In_191);
or U196 (N_196,In_236,In_143);
and U197 (N_197,In_246,In_8);
nor U198 (N_198,In_396,In_118);
nand U199 (N_199,In_264,In_169);
nand U200 (N_200,In_347,In_271);
nor U201 (N_201,In_415,In_407);
or U202 (N_202,In_98,In_227);
nand U203 (N_203,In_122,In_444);
xnor U204 (N_204,In_81,In_441);
and U205 (N_205,In_141,In_117);
and U206 (N_206,In_69,In_9);
and U207 (N_207,In_61,In_230);
nor U208 (N_208,In_401,In_142);
or U209 (N_209,In_11,In_237);
nor U210 (N_210,In_306,In_163);
nand U211 (N_211,In_425,In_427);
nand U212 (N_212,In_145,In_435);
nand U213 (N_213,In_374,In_87);
and U214 (N_214,In_10,In_433);
nor U215 (N_215,In_312,In_417);
nor U216 (N_216,In_137,In_115);
and U217 (N_217,In_377,In_421);
or U218 (N_218,In_245,In_480);
nand U219 (N_219,In_155,In_281);
or U220 (N_220,In_357,In_348);
xnor U221 (N_221,In_222,In_244);
nand U222 (N_222,In_148,In_412);
nand U223 (N_223,In_37,In_422);
or U224 (N_224,In_477,In_210);
and U225 (N_225,In_90,In_15);
nor U226 (N_226,In_13,In_461);
nor U227 (N_227,In_384,In_101);
or U228 (N_228,In_259,In_76);
nor U229 (N_229,In_406,In_41);
nand U230 (N_230,In_280,In_255);
nor U231 (N_231,In_146,In_218);
and U232 (N_232,In_157,In_150);
and U233 (N_233,In_483,In_310);
or U234 (N_234,In_32,In_50);
or U235 (N_235,In_262,In_166);
xnor U236 (N_236,In_498,In_416);
and U237 (N_237,In_220,In_250);
and U238 (N_238,In_418,In_450);
or U239 (N_239,In_389,In_0);
xnor U240 (N_240,In_120,In_290);
or U241 (N_241,In_380,In_105);
and U242 (N_242,In_29,In_207);
nor U243 (N_243,In_360,In_300);
and U244 (N_244,In_361,In_350);
and U245 (N_245,In_302,In_79);
and U246 (N_246,In_391,In_423);
nor U247 (N_247,In_398,In_85);
nor U248 (N_248,In_292,In_52);
or U249 (N_249,In_125,In_367);
or U250 (N_250,In_255,In_444);
and U251 (N_251,In_169,In_86);
or U252 (N_252,In_207,In_292);
and U253 (N_253,In_303,In_132);
and U254 (N_254,In_355,In_293);
nor U255 (N_255,In_156,In_75);
and U256 (N_256,In_499,In_411);
nand U257 (N_257,In_224,In_431);
and U258 (N_258,In_348,In_21);
and U259 (N_259,In_48,In_359);
nand U260 (N_260,In_28,In_349);
nor U261 (N_261,In_4,In_293);
and U262 (N_262,In_268,In_116);
or U263 (N_263,In_230,In_222);
or U264 (N_264,In_240,In_451);
nor U265 (N_265,In_460,In_188);
xor U266 (N_266,In_412,In_384);
nand U267 (N_267,In_45,In_259);
nand U268 (N_268,In_10,In_459);
and U269 (N_269,In_149,In_250);
nand U270 (N_270,In_298,In_19);
or U271 (N_271,In_411,In_227);
nor U272 (N_272,In_379,In_212);
or U273 (N_273,In_329,In_387);
nor U274 (N_274,In_201,In_37);
and U275 (N_275,In_467,In_214);
and U276 (N_276,In_430,In_232);
and U277 (N_277,In_411,In_207);
or U278 (N_278,In_270,In_210);
and U279 (N_279,In_422,In_473);
nand U280 (N_280,In_450,In_82);
and U281 (N_281,In_314,In_309);
or U282 (N_282,In_239,In_333);
and U283 (N_283,In_424,In_47);
and U284 (N_284,In_370,In_158);
or U285 (N_285,In_320,In_482);
xnor U286 (N_286,In_499,In_8);
nand U287 (N_287,In_443,In_248);
or U288 (N_288,In_198,In_306);
nor U289 (N_289,In_350,In_419);
nor U290 (N_290,In_281,In_498);
nand U291 (N_291,In_342,In_488);
nand U292 (N_292,In_483,In_169);
nor U293 (N_293,In_435,In_420);
nor U294 (N_294,In_328,In_439);
nor U295 (N_295,In_430,In_7);
and U296 (N_296,In_71,In_233);
or U297 (N_297,In_265,In_80);
and U298 (N_298,In_348,In_87);
nor U299 (N_299,In_119,In_231);
nor U300 (N_300,In_49,In_27);
and U301 (N_301,In_58,In_46);
and U302 (N_302,In_33,In_59);
nand U303 (N_303,In_273,In_243);
nor U304 (N_304,In_273,In_362);
xnor U305 (N_305,In_474,In_265);
nor U306 (N_306,In_26,In_45);
nor U307 (N_307,In_263,In_37);
or U308 (N_308,In_230,In_196);
and U309 (N_309,In_367,In_261);
or U310 (N_310,In_186,In_420);
nor U311 (N_311,In_485,In_168);
and U312 (N_312,In_352,In_463);
nand U313 (N_313,In_192,In_236);
or U314 (N_314,In_352,In_161);
nor U315 (N_315,In_3,In_57);
nand U316 (N_316,In_199,In_228);
nor U317 (N_317,In_43,In_357);
nor U318 (N_318,In_258,In_484);
or U319 (N_319,In_44,In_411);
and U320 (N_320,In_85,In_408);
nor U321 (N_321,In_116,In_460);
nand U322 (N_322,In_496,In_467);
nand U323 (N_323,In_496,In_222);
or U324 (N_324,In_410,In_386);
and U325 (N_325,In_468,In_8);
and U326 (N_326,In_198,In_94);
and U327 (N_327,In_236,In_303);
and U328 (N_328,In_307,In_78);
and U329 (N_329,In_199,In_109);
nand U330 (N_330,In_457,In_466);
nand U331 (N_331,In_45,In_10);
nand U332 (N_332,In_477,In_241);
and U333 (N_333,In_357,In_367);
nor U334 (N_334,In_383,In_482);
nand U335 (N_335,In_56,In_434);
and U336 (N_336,In_95,In_383);
or U337 (N_337,In_171,In_429);
nand U338 (N_338,In_53,In_430);
or U339 (N_339,In_190,In_462);
and U340 (N_340,In_485,In_214);
nor U341 (N_341,In_3,In_172);
and U342 (N_342,In_61,In_314);
nand U343 (N_343,In_138,In_403);
nor U344 (N_344,In_99,In_234);
nor U345 (N_345,In_375,In_371);
nor U346 (N_346,In_475,In_201);
or U347 (N_347,In_440,In_183);
nor U348 (N_348,In_311,In_361);
xor U349 (N_349,In_234,In_414);
or U350 (N_350,In_424,In_7);
nor U351 (N_351,In_372,In_456);
nor U352 (N_352,In_317,In_155);
or U353 (N_353,In_59,In_166);
nor U354 (N_354,In_421,In_149);
nand U355 (N_355,In_191,In_391);
nor U356 (N_356,In_206,In_224);
nor U357 (N_357,In_282,In_110);
nand U358 (N_358,In_21,In_340);
nand U359 (N_359,In_223,In_320);
or U360 (N_360,In_226,In_197);
nor U361 (N_361,In_86,In_471);
nand U362 (N_362,In_415,In_205);
nand U363 (N_363,In_314,In_289);
nor U364 (N_364,In_455,In_65);
nor U365 (N_365,In_263,In_438);
and U366 (N_366,In_306,In_190);
or U367 (N_367,In_474,In_238);
nand U368 (N_368,In_395,In_192);
and U369 (N_369,In_255,In_323);
or U370 (N_370,In_187,In_199);
xnor U371 (N_371,In_307,In_17);
or U372 (N_372,In_470,In_197);
and U373 (N_373,In_83,In_367);
and U374 (N_374,In_195,In_160);
nor U375 (N_375,In_126,In_365);
and U376 (N_376,In_377,In_175);
or U377 (N_377,In_479,In_107);
nand U378 (N_378,In_268,In_75);
or U379 (N_379,In_310,In_449);
and U380 (N_380,In_288,In_135);
nor U381 (N_381,In_317,In_215);
nand U382 (N_382,In_164,In_413);
or U383 (N_383,In_176,In_278);
nand U384 (N_384,In_82,In_115);
or U385 (N_385,In_102,In_176);
or U386 (N_386,In_369,In_432);
nand U387 (N_387,In_395,In_455);
and U388 (N_388,In_325,In_370);
and U389 (N_389,In_346,In_138);
and U390 (N_390,In_237,In_454);
or U391 (N_391,In_208,In_248);
nor U392 (N_392,In_165,In_413);
and U393 (N_393,In_268,In_185);
and U394 (N_394,In_170,In_408);
and U395 (N_395,In_52,In_189);
nand U396 (N_396,In_281,In_24);
xor U397 (N_397,In_456,In_163);
or U398 (N_398,In_239,In_235);
and U399 (N_399,In_298,In_293);
nor U400 (N_400,In_385,In_170);
and U401 (N_401,In_301,In_203);
nand U402 (N_402,In_254,In_141);
nand U403 (N_403,In_446,In_488);
and U404 (N_404,In_50,In_73);
and U405 (N_405,In_112,In_187);
or U406 (N_406,In_84,In_6);
nand U407 (N_407,In_337,In_3);
or U408 (N_408,In_129,In_280);
nand U409 (N_409,In_304,In_94);
xnor U410 (N_410,In_345,In_162);
nor U411 (N_411,In_371,In_323);
and U412 (N_412,In_282,In_325);
or U413 (N_413,In_68,In_10);
nand U414 (N_414,In_235,In_2);
nand U415 (N_415,In_112,In_134);
nand U416 (N_416,In_360,In_40);
nor U417 (N_417,In_288,In_368);
nand U418 (N_418,In_457,In_284);
nor U419 (N_419,In_300,In_286);
and U420 (N_420,In_397,In_76);
or U421 (N_421,In_262,In_388);
nand U422 (N_422,In_136,In_304);
and U423 (N_423,In_305,In_108);
nand U424 (N_424,In_250,In_359);
or U425 (N_425,In_24,In_184);
nand U426 (N_426,In_268,In_66);
nor U427 (N_427,In_30,In_314);
nor U428 (N_428,In_419,In_365);
or U429 (N_429,In_4,In_188);
xnor U430 (N_430,In_351,In_262);
nor U431 (N_431,In_25,In_165);
nand U432 (N_432,In_101,In_4);
and U433 (N_433,In_348,In_471);
and U434 (N_434,In_101,In_20);
and U435 (N_435,In_256,In_183);
and U436 (N_436,In_119,In_386);
nor U437 (N_437,In_499,In_30);
nand U438 (N_438,In_164,In_16);
nor U439 (N_439,In_390,In_258);
nor U440 (N_440,In_257,In_379);
nand U441 (N_441,In_167,In_241);
or U442 (N_442,In_321,In_391);
or U443 (N_443,In_22,In_46);
nand U444 (N_444,In_73,In_416);
xnor U445 (N_445,In_414,In_358);
nand U446 (N_446,In_216,In_400);
or U447 (N_447,In_42,In_331);
and U448 (N_448,In_188,In_53);
and U449 (N_449,In_254,In_68);
and U450 (N_450,In_214,In_25);
xnor U451 (N_451,In_128,In_423);
nor U452 (N_452,In_15,In_496);
and U453 (N_453,In_269,In_415);
nor U454 (N_454,In_155,In_80);
nand U455 (N_455,In_445,In_194);
or U456 (N_456,In_188,In_404);
and U457 (N_457,In_190,In_376);
xor U458 (N_458,In_142,In_291);
and U459 (N_459,In_186,In_172);
or U460 (N_460,In_143,In_202);
nor U461 (N_461,In_474,In_258);
nand U462 (N_462,In_462,In_330);
or U463 (N_463,In_48,In_377);
and U464 (N_464,In_337,In_5);
nor U465 (N_465,In_303,In_17);
or U466 (N_466,In_446,In_24);
and U467 (N_467,In_381,In_26);
or U468 (N_468,In_141,In_382);
or U469 (N_469,In_141,In_355);
or U470 (N_470,In_453,In_86);
nand U471 (N_471,In_7,In_28);
or U472 (N_472,In_308,In_89);
and U473 (N_473,In_392,In_432);
and U474 (N_474,In_422,In_482);
or U475 (N_475,In_217,In_399);
or U476 (N_476,In_277,In_115);
xor U477 (N_477,In_276,In_30);
and U478 (N_478,In_62,In_36);
or U479 (N_479,In_413,In_433);
or U480 (N_480,In_247,In_362);
and U481 (N_481,In_308,In_188);
nor U482 (N_482,In_312,In_457);
or U483 (N_483,In_225,In_67);
and U484 (N_484,In_314,In_71);
and U485 (N_485,In_310,In_443);
nor U486 (N_486,In_183,In_418);
nand U487 (N_487,In_177,In_347);
nor U488 (N_488,In_257,In_86);
and U489 (N_489,In_424,In_316);
nand U490 (N_490,In_375,In_157);
or U491 (N_491,In_140,In_485);
and U492 (N_492,In_364,In_168);
nor U493 (N_493,In_145,In_164);
nor U494 (N_494,In_140,In_305);
and U495 (N_495,In_462,In_31);
nor U496 (N_496,In_286,In_5);
and U497 (N_497,In_490,In_239);
nand U498 (N_498,In_96,In_116);
and U499 (N_499,In_390,In_379);
or U500 (N_500,In_474,In_150);
nand U501 (N_501,In_400,In_1);
and U502 (N_502,In_346,In_358);
nand U503 (N_503,In_349,In_297);
nor U504 (N_504,In_349,In_416);
nor U505 (N_505,In_288,In_58);
nor U506 (N_506,In_336,In_320);
nor U507 (N_507,In_280,In_95);
nor U508 (N_508,In_104,In_18);
and U509 (N_509,In_357,In_199);
or U510 (N_510,In_341,In_74);
and U511 (N_511,In_136,In_131);
nand U512 (N_512,In_376,In_280);
nand U513 (N_513,In_85,In_336);
and U514 (N_514,In_224,In_69);
or U515 (N_515,In_413,In_283);
nand U516 (N_516,In_420,In_20);
xor U517 (N_517,In_172,In_96);
or U518 (N_518,In_415,In_486);
and U519 (N_519,In_25,In_450);
nand U520 (N_520,In_293,In_100);
nor U521 (N_521,In_308,In_403);
nand U522 (N_522,In_83,In_217);
nand U523 (N_523,In_200,In_58);
xor U524 (N_524,In_66,In_107);
or U525 (N_525,In_463,In_431);
nand U526 (N_526,In_78,In_384);
and U527 (N_527,In_39,In_113);
and U528 (N_528,In_479,In_208);
nand U529 (N_529,In_58,In_151);
and U530 (N_530,In_40,In_186);
and U531 (N_531,In_6,In_451);
nor U532 (N_532,In_34,In_432);
and U533 (N_533,In_439,In_290);
nand U534 (N_534,In_320,In_433);
and U535 (N_535,In_215,In_302);
and U536 (N_536,In_310,In_441);
and U537 (N_537,In_58,In_488);
or U538 (N_538,In_356,In_204);
nor U539 (N_539,In_392,In_270);
or U540 (N_540,In_95,In_374);
nand U541 (N_541,In_437,In_347);
and U542 (N_542,In_236,In_57);
and U543 (N_543,In_85,In_88);
nor U544 (N_544,In_180,In_233);
and U545 (N_545,In_409,In_452);
or U546 (N_546,In_259,In_233);
xor U547 (N_547,In_230,In_130);
nor U548 (N_548,In_347,In_230);
or U549 (N_549,In_232,In_225);
or U550 (N_550,In_158,In_224);
xnor U551 (N_551,In_215,In_252);
or U552 (N_552,In_68,In_366);
nor U553 (N_553,In_449,In_169);
and U554 (N_554,In_198,In_488);
nand U555 (N_555,In_300,In_232);
nor U556 (N_556,In_87,In_186);
nor U557 (N_557,In_449,In_299);
nor U558 (N_558,In_400,In_356);
xor U559 (N_559,In_90,In_258);
nand U560 (N_560,In_16,In_236);
xor U561 (N_561,In_469,In_131);
nor U562 (N_562,In_225,In_436);
or U563 (N_563,In_128,In_175);
and U564 (N_564,In_279,In_413);
nor U565 (N_565,In_174,In_9);
or U566 (N_566,In_82,In_471);
nand U567 (N_567,In_222,In_475);
nor U568 (N_568,In_415,In_216);
and U569 (N_569,In_269,In_414);
nand U570 (N_570,In_282,In_224);
or U571 (N_571,In_403,In_258);
nor U572 (N_572,In_379,In_231);
and U573 (N_573,In_165,In_57);
nor U574 (N_574,In_157,In_396);
or U575 (N_575,In_367,In_26);
nand U576 (N_576,In_253,In_400);
or U577 (N_577,In_249,In_33);
and U578 (N_578,In_10,In_114);
or U579 (N_579,In_186,In_353);
nor U580 (N_580,In_297,In_9);
nor U581 (N_581,In_435,In_84);
nand U582 (N_582,In_246,In_316);
or U583 (N_583,In_46,In_288);
or U584 (N_584,In_0,In_120);
nor U585 (N_585,In_461,In_399);
or U586 (N_586,In_84,In_319);
nand U587 (N_587,In_309,In_81);
nor U588 (N_588,In_476,In_497);
nor U589 (N_589,In_373,In_337);
or U590 (N_590,In_377,In_111);
and U591 (N_591,In_363,In_103);
nor U592 (N_592,In_217,In_33);
nand U593 (N_593,In_163,In_406);
or U594 (N_594,In_316,In_387);
nor U595 (N_595,In_427,In_193);
nand U596 (N_596,In_239,In_67);
or U597 (N_597,In_158,In_239);
nor U598 (N_598,In_41,In_415);
xor U599 (N_599,In_412,In_332);
and U600 (N_600,In_247,In_71);
and U601 (N_601,In_312,In_177);
and U602 (N_602,In_446,In_463);
and U603 (N_603,In_115,In_103);
nand U604 (N_604,In_404,In_121);
nor U605 (N_605,In_221,In_313);
xnor U606 (N_606,In_381,In_122);
nand U607 (N_607,In_147,In_340);
nor U608 (N_608,In_140,In_227);
nor U609 (N_609,In_379,In_314);
nand U610 (N_610,In_439,In_298);
nor U611 (N_611,In_459,In_88);
or U612 (N_612,In_371,In_450);
nor U613 (N_613,In_80,In_493);
nand U614 (N_614,In_109,In_414);
and U615 (N_615,In_475,In_372);
nor U616 (N_616,In_403,In_76);
or U617 (N_617,In_35,In_344);
and U618 (N_618,In_495,In_202);
nand U619 (N_619,In_438,In_400);
nand U620 (N_620,In_197,In_123);
nand U621 (N_621,In_48,In_38);
nand U622 (N_622,In_80,In_342);
nand U623 (N_623,In_228,In_274);
nand U624 (N_624,In_394,In_248);
or U625 (N_625,In_492,In_140);
and U626 (N_626,In_496,In_192);
nor U627 (N_627,In_84,In_122);
or U628 (N_628,In_30,In_41);
and U629 (N_629,In_105,In_415);
nor U630 (N_630,In_263,In_300);
nor U631 (N_631,In_222,In_149);
or U632 (N_632,In_228,In_202);
and U633 (N_633,In_463,In_232);
nand U634 (N_634,In_259,In_280);
or U635 (N_635,In_274,In_356);
or U636 (N_636,In_15,In_467);
nand U637 (N_637,In_323,In_421);
or U638 (N_638,In_344,In_496);
nor U639 (N_639,In_257,In_448);
and U640 (N_640,In_232,In_302);
and U641 (N_641,In_121,In_479);
nor U642 (N_642,In_436,In_65);
nand U643 (N_643,In_277,In_471);
nand U644 (N_644,In_351,In_71);
or U645 (N_645,In_138,In_411);
nand U646 (N_646,In_69,In_21);
and U647 (N_647,In_147,In_26);
nor U648 (N_648,In_280,In_422);
and U649 (N_649,In_278,In_101);
and U650 (N_650,In_178,In_403);
and U651 (N_651,In_253,In_202);
or U652 (N_652,In_100,In_474);
and U653 (N_653,In_230,In_159);
and U654 (N_654,In_419,In_152);
nor U655 (N_655,In_184,In_336);
or U656 (N_656,In_231,In_9);
and U657 (N_657,In_357,In_302);
and U658 (N_658,In_170,In_139);
nor U659 (N_659,In_45,In_289);
nor U660 (N_660,In_98,In_401);
and U661 (N_661,In_463,In_269);
nand U662 (N_662,In_135,In_428);
nand U663 (N_663,In_421,In_281);
or U664 (N_664,In_194,In_474);
and U665 (N_665,In_231,In_140);
nand U666 (N_666,In_130,In_219);
xor U667 (N_667,In_296,In_167);
or U668 (N_668,In_204,In_488);
and U669 (N_669,In_22,In_459);
or U670 (N_670,In_325,In_111);
and U671 (N_671,In_244,In_187);
nand U672 (N_672,In_346,In_191);
nor U673 (N_673,In_448,In_273);
nor U674 (N_674,In_191,In_230);
nor U675 (N_675,In_266,In_421);
or U676 (N_676,In_66,In_366);
and U677 (N_677,In_46,In_164);
or U678 (N_678,In_191,In_30);
nor U679 (N_679,In_109,In_334);
nand U680 (N_680,In_154,In_343);
and U681 (N_681,In_425,In_434);
nor U682 (N_682,In_347,In_267);
nand U683 (N_683,In_115,In_79);
or U684 (N_684,In_153,In_402);
and U685 (N_685,In_276,In_117);
or U686 (N_686,In_332,In_114);
nand U687 (N_687,In_293,In_50);
nor U688 (N_688,In_225,In_371);
and U689 (N_689,In_50,In_490);
and U690 (N_690,In_58,In_233);
or U691 (N_691,In_337,In_433);
nor U692 (N_692,In_486,In_142);
nand U693 (N_693,In_308,In_118);
or U694 (N_694,In_338,In_400);
and U695 (N_695,In_376,In_413);
and U696 (N_696,In_484,In_217);
nor U697 (N_697,In_426,In_438);
nor U698 (N_698,In_82,In_447);
and U699 (N_699,In_240,In_337);
nand U700 (N_700,In_448,In_178);
nor U701 (N_701,In_340,In_142);
or U702 (N_702,In_105,In_442);
and U703 (N_703,In_161,In_226);
nand U704 (N_704,In_398,In_182);
and U705 (N_705,In_64,In_127);
or U706 (N_706,In_11,In_226);
or U707 (N_707,In_73,In_151);
or U708 (N_708,In_390,In_371);
nor U709 (N_709,In_459,In_402);
and U710 (N_710,In_2,In_449);
and U711 (N_711,In_123,In_252);
nand U712 (N_712,In_419,In_119);
nor U713 (N_713,In_281,In_359);
nor U714 (N_714,In_380,In_310);
or U715 (N_715,In_384,In_107);
and U716 (N_716,In_455,In_272);
or U717 (N_717,In_438,In_169);
nand U718 (N_718,In_463,In_265);
nand U719 (N_719,In_378,In_489);
nor U720 (N_720,In_94,In_173);
or U721 (N_721,In_46,In_205);
nand U722 (N_722,In_328,In_136);
nor U723 (N_723,In_346,In_40);
and U724 (N_724,In_417,In_316);
nor U725 (N_725,In_333,In_45);
nor U726 (N_726,In_47,In_414);
and U727 (N_727,In_92,In_471);
nor U728 (N_728,In_8,In_314);
nor U729 (N_729,In_292,In_224);
or U730 (N_730,In_38,In_147);
nor U731 (N_731,In_202,In_22);
nor U732 (N_732,In_80,In_344);
or U733 (N_733,In_123,In_305);
xnor U734 (N_734,In_65,In_165);
nand U735 (N_735,In_240,In_238);
or U736 (N_736,In_461,In_176);
and U737 (N_737,In_355,In_216);
or U738 (N_738,In_191,In_14);
or U739 (N_739,In_19,In_191);
nor U740 (N_740,In_366,In_116);
or U741 (N_741,In_408,In_421);
nor U742 (N_742,In_440,In_344);
and U743 (N_743,In_427,In_203);
and U744 (N_744,In_385,In_80);
and U745 (N_745,In_471,In_481);
or U746 (N_746,In_34,In_341);
or U747 (N_747,In_86,In_94);
nand U748 (N_748,In_93,In_68);
and U749 (N_749,In_205,In_381);
or U750 (N_750,In_456,In_487);
nand U751 (N_751,In_195,In_453);
nor U752 (N_752,In_257,In_457);
and U753 (N_753,In_304,In_495);
and U754 (N_754,In_75,In_166);
nor U755 (N_755,In_435,In_328);
and U756 (N_756,In_39,In_470);
or U757 (N_757,In_393,In_28);
nand U758 (N_758,In_270,In_225);
and U759 (N_759,In_493,In_445);
nor U760 (N_760,In_30,In_181);
nor U761 (N_761,In_188,In_153);
or U762 (N_762,In_126,In_275);
xor U763 (N_763,In_360,In_27);
or U764 (N_764,In_240,In_5);
nand U765 (N_765,In_486,In_422);
or U766 (N_766,In_52,In_493);
nand U767 (N_767,In_460,In_227);
or U768 (N_768,In_438,In_159);
nand U769 (N_769,In_246,In_377);
and U770 (N_770,In_307,In_309);
nand U771 (N_771,In_320,In_168);
and U772 (N_772,In_329,In_285);
nand U773 (N_773,In_24,In_308);
nand U774 (N_774,In_190,In_309);
nor U775 (N_775,In_489,In_436);
nand U776 (N_776,In_444,In_15);
or U777 (N_777,In_339,In_325);
and U778 (N_778,In_278,In_107);
or U779 (N_779,In_69,In_295);
or U780 (N_780,In_24,In_450);
or U781 (N_781,In_368,In_45);
nor U782 (N_782,In_224,In_372);
nor U783 (N_783,In_371,In_43);
or U784 (N_784,In_349,In_121);
and U785 (N_785,In_84,In_82);
nand U786 (N_786,In_5,In_338);
nand U787 (N_787,In_342,In_296);
nor U788 (N_788,In_115,In_285);
nand U789 (N_789,In_460,In_118);
nand U790 (N_790,In_65,In_153);
nor U791 (N_791,In_45,In_100);
nor U792 (N_792,In_75,In_70);
or U793 (N_793,In_300,In_214);
nand U794 (N_794,In_106,In_172);
or U795 (N_795,In_147,In_368);
nor U796 (N_796,In_296,In_349);
or U797 (N_797,In_386,In_445);
and U798 (N_798,In_493,In_300);
nand U799 (N_799,In_29,In_85);
nor U800 (N_800,In_313,In_54);
nand U801 (N_801,In_183,In_357);
nand U802 (N_802,In_326,In_111);
nor U803 (N_803,In_484,In_487);
nor U804 (N_804,In_405,In_298);
nor U805 (N_805,In_87,In_158);
and U806 (N_806,In_278,In_416);
and U807 (N_807,In_318,In_35);
or U808 (N_808,In_397,In_314);
nand U809 (N_809,In_386,In_446);
nor U810 (N_810,In_393,In_488);
or U811 (N_811,In_440,In_425);
nor U812 (N_812,In_462,In_316);
nor U813 (N_813,In_293,In_231);
or U814 (N_814,In_34,In_465);
and U815 (N_815,In_30,In_35);
nand U816 (N_816,In_411,In_40);
or U817 (N_817,In_106,In_397);
or U818 (N_818,In_280,In_50);
nand U819 (N_819,In_33,In_383);
nand U820 (N_820,In_225,In_406);
xor U821 (N_821,In_301,In_253);
or U822 (N_822,In_466,In_323);
nor U823 (N_823,In_204,In_406);
xor U824 (N_824,In_19,In_206);
nand U825 (N_825,In_351,In_406);
nor U826 (N_826,In_388,In_34);
nand U827 (N_827,In_383,In_344);
nand U828 (N_828,In_46,In_43);
or U829 (N_829,In_166,In_105);
or U830 (N_830,In_472,In_161);
nor U831 (N_831,In_481,In_93);
nor U832 (N_832,In_313,In_201);
nor U833 (N_833,In_376,In_225);
and U834 (N_834,In_29,In_275);
or U835 (N_835,In_75,In_150);
or U836 (N_836,In_253,In_308);
nand U837 (N_837,In_367,In_258);
and U838 (N_838,In_36,In_20);
and U839 (N_839,In_310,In_66);
nor U840 (N_840,In_216,In_499);
nor U841 (N_841,In_495,In_282);
nand U842 (N_842,In_153,In_190);
nand U843 (N_843,In_426,In_351);
or U844 (N_844,In_23,In_452);
and U845 (N_845,In_262,In_304);
nand U846 (N_846,In_426,In_198);
nor U847 (N_847,In_340,In_179);
nor U848 (N_848,In_39,In_198);
nor U849 (N_849,In_335,In_243);
nor U850 (N_850,In_79,In_100);
and U851 (N_851,In_42,In_475);
or U852 (N_852,In_289,In_469);
and U853 (N_853,In_474,In_250);
nand U854 (N_854,In_287,In_310);
nor U855 (N_855,In_299,In_424);
or U856 (N_856,In_481,In_213);
and U857 (N_857,In_225,In_148);
nor U858 (N_858,In_348,In_157);
and U859 (N_859,In_132,In_241);
nand U860 (N_860,In_267,In_130);
nand U861 (N_861,In_451,In_130);
or U862 (N_862,In_53,In_492);
xnor U863 (N_863,In_164,In_174);
and U864 (N_864,In_21,In_306);
and U865 (N_865,In_450,In_32);
or U866 (N_866,In_475,In_394);
nor U867 (N_867,In_300,In_246);
nor U868 (N_868,In_451,In_344);
nand U869 (N_869,In_237,In_105);
and U870 (N_870,In_468,In_179);
nor U871 (N_871,In_388,In_218);
nor U872 (N_872,In_143,In_144);
nor U873 (N_873,In_320,In_99);
xor U874 (N_874,In_372,In_490);
nor U875 (N_875,In_368,In_133);
and U876 (N_876,In_282,In_35);
and U877 (N_877,In_262,In_372);
nand U878 (N_878,In_445,In_354);
and U879 (N_879,In_28,In_113);
nand U880 (N_880,In_224,In_75);
or U881 (N_881,In_492,In_224);
nand U882 (N_882,In_300,In_55);
and U883 (N_883,In_149,In_206);
nor U884 (N_884,In_111,In_160);
or U885 (N_885,In_305,In_121);
nor U886 (N_886,In_118,In_409);
nand U887 (N_887,In_82,In_186);
nor U888 (N_888,In_287,In_383);
nand U889 (N_889,In_216,In_141);
or U890 (N_890,In_260,In_155);
nand U891 (N_891,In_113,In_269);
nand U892 (N_892,In_296,In_139);
or U893 (N_893,In_348,In_143);
and U894 (N_894,In_317,In_179);
nand U895 (N_895,In_88,In_182);
or U896 (N_896,In_426,In_2);
or U897 (N_897,In_366,In_321);
or U898 (N_898,In_421,In_32);
and U899 (N_899,In_438,In_268);
and U900 (N_900,In_195,In_471);
or U901 (N_901,In_282,In_146);
nand U902 (N_902,In_205,In_147);
and U903 (N_903,In_353,In_466);
and U904 (N_904,In_7,In_332);
nor U905 (N_905,In_119,In_380);
nand U906 (N_906,In_83,In_498);
nand U907 (N_907,In_118,In_394);
and U908 (N_908,In_78,In_408);
nor U909 (N_909,In_51,In_450);
and U910 (N_910,In_3,In_314);
and U911 (N_911,In_475,In_85);
nand U912 (N_912,In_472,In_64);
nand U913 (N_913,In_317,In_446);
nand U914 (N_914,In_475,In_410);
nor U915 (N_915,In_261,In_33);
or U916 (N_916,In_78,In_51);
nor U917 (N_917,In_255,In_57);
nor U918 (N_918,In_426,In_291);
or U919 (N_919,In_257,In_73);
or U920 (N_920,In_302,In_382);
or U921 (N_921,In_191,In_325);
and U922 (N_922,In_423,In_351);
and U923 (N_923,In_0,In_234);
and U924 (N_924,In_418,In_270);
nor U925 (N_925,In_169,In_154);
and U926 (N_926,In_353,In_339);
nor U927 (N_927,In_256,In_130);
and U928 (N_928,In_64,In_302);
or U929 (N_929,In_37,In_10);
or U930 (N_930,In_26,In_189);
nor U931 (N_931,In_366,In_268);
nor U932 (N_932,In_210,In_7);
and U933 (N_933,In_432,In_81);
nand U934 (N_934,In_354,In_209);
nor U935 (N_935,In_242,In_398);
nor U936 (N_936,In_91,In_122);
and U937 (N_937,In_498,In_153);
or U938 (N_938,In_63,In_463);
nand U939 (N_939,In_137,In_63);
or U940 (N_940,In_27,In_120);
and U941 (N_941,In_148,In_198);
or U942 (N_942,In_392,In_23);
or U943 (N_943,In_72,In_360);
nand U944 (N_944,In_87,In_104);
nand U945 (N_945,In_436,In_496);
and U946 (N_946,In_475,In_99);
or U947 (N_947,In_17,In_162);
nor U948 (N_948,In_430,In_174);
nor U949 (N_949,In_31,In_260);
nand U950 (N_950,In_221,In_365);
or U951 (N_951,In_344,In_164);
or U952 (N_952,In_136,In_13);
nand U953 (N_953,In_55,In_438);
and U954 (N_954,In_185,In_254);
xor U955 (N_955,In_31,In_333);
nor U956 (N_956,In_168,In_378);
nor U957 (N_957,In_360,In_144);
nor U958 (N_958,In_418,In_20);
nor U959 (N_959,In_138,In_74);
nor U960 (N_960,In_110,In_73);
and U961 (N_961,In_37,In_239);
or U962 (N_962,In_390,In_391);
nor U963 (N_963,In_434,In_17);
and U964 (N_964,In_322,In_308);
nor U965 (N_965,In_454,In_251);
nor U966 (N_966,In_345,In_306);
or U967 (N_967,In_60,In_281);
and U968 (N_968,In_7,In_367);
nand U969 (N_969,In_464,In_383);
nor U970 (N_970,In_231,In_134);
or U971 (N_971,In_314,In_136);
nor U972 (N_972,In_33,In_262);
or U973 (N_973,In_94,In_395);
nand U974 (N_974,In_285,In_219);
nand U975 (N_975,In_356,In_459);
and U976 (N_976,In_421,In_140);
or U977 (N_977,In_386,In_208);
nor U978 (N_978,In_174,In_19);
nand U979 (N_979,In_123,In_147);
nand U980 (N_980,In_66,In_274);
nor U981 (N_981,In_368,In_295);
xnor U982 (N_982,In_108,In_229);
nand U983 (N_983,In_182,In_307);
nand U984 (N_984,In_477,In_423);
nor U985 (N_985,In_94,In_472);
nor U986 (N_986,In_323,In_234);
or U987 (N_987,In_397,In_498);
and U988 (N_988,In_328,In_343);
nor U989 (N_989,In_129,In_479);
nand U990 (N_990,In_459,In_235);
xnor U991 (N_991,In_360,In_165);
nand U992 (N_992,In_305,In_189);
nand U993 (N_993,In_224,In_28);
nor U994 (N_994,In_186,In_383);
nor U995 (N_995,In_383,In_293);
nor U996 (N_996,In_488,In_249);
or U997 (N_997,In_62,In_445);
and U998 (N_998,In_155,In_82);
nor U999 (N_999,In_5,In_87);
and U1000 (N_1000,N_896,N_341);
and U1001 (N_1001,N_451,N_796);
or U1002 (N_1002,N_408,N_363);
xor U1003 (N_1003,N_786,N_19);
and U1004 (N_1004,N_249,N_885);
nor U1005 (N_1005,N_120,N_939);
or U1006 (N_1006,N_756,N_614);
and U1007 (N_1007,N_958,N_811);
and U1008 (N_1008,N_287,N_452);
and U1009 (N_1009,N_41,N_83);
and U1010 (N_1010,N_340,N_847);
nand U1011 (N_1011,N_623,N_213);
nand U1012 (N_1012,N_160,N_976);
xor U1013 (N_1013,N_822,N_436);
and U1014 (N_1014,N_33,N_357);
or U1015 (N_1015,N_409,N_520);
nand U1016 (N_1016,N_485,N_379);
or U1017 (N_1017,N_434,N_498);
and U1018 (N_1018,N_543,N_996);
xnor U1019 (N_1019,N_572,N_376);
nor U1020 (N_1020,N_37,N_992);
or U1021 (N_1021,N_365,N_948);
nand U1022 (N_1022,N_153,N_978);
nor U1023 (N_1023,N_273,N_626);
nor U1024 (N_1024,N_772,N_562);
nand U1025 (N_1025,N_182,N_905);
nand U1026 (N_1026,N_960,N_611);
or U1027 (N_1027,N_283,N_269);
nor U1028 (N_1028,N_123,N_410);
and U1029 (N_1029,N_58,N_570);
nor U1030 (N_1030,N_121,N_829);
nand U1031 (N_1031,N_834,N_916);
or U1032 (N_1032,N_350,N_494);
or U1033 (N_1033,N_354,N_762);
nand U1034 (N_1034,N_573,N_659);
and U1035 (N_1035,N_823,N_802);
nand U1036 (N_1036,N_858,N_922);
and U1037 (N_1037,N_103,N_920);
nor U1038 (N_1038,N_335,N_705);
nand U1039 (N_1039,N_233,N_857);
and U1040 (N_1040,N_583,N_691);
and U1041 (N_1041,N_398,N_527);
nor U1042 (N_1042,N_404,N_985);
or U1043 (N_1043,N_633,N_296);
nor U1044 (N_1044,N_568,N_293);
nand U1045 (N_1045,N_889,N_78);
and U1046 (N_1046,N_251,N_743);
or U1047 (N_1047,N_432,N_699);
xor U1048 (N_1048,N_940,N_644);
or U1049 (N_1049,N_735,N_918);
or U1050 (N_1050,N_443,N_62);
or U1051 (N_1051,N_446,N_926);
xor U1052 (N_1052,N_591,N_94);
or U1053 (N_1053,N_17,N_702);
and U1054 (N_1054,N_390,N_427);
or U1055 (N_1055,N_238,N_177);
nand U1056 (N_1056,N_197,N_710);
and U1057 (N_1057,N_317,N_368);
nand U1058 (N_1058,N_412,N_848);
or U1059 (N_1059,N_216,N_165);
and U1060 (N_1060,N_284,N_453);
nand U1061 (N_1061,N_618,N_79);
and U1062 (N_1062,N_619,N_264);
nand U1063 (N_1063,N_206,N_741);
nor U1064 (N_1064,N_47,N_88);
nand U1065 (N_1065,N_183,N_538);
nand U1066 (N_1066,N_243,N_556);
or U1067 (N_1067,N_674,N_860);
nor U1068 (N_1068,N_508,N_178);
nor U1069 (N_1069,N_715,N_113);
or U1070 (N_1070,N_731,N_465);
nand U1071 (N_1071,N_523,N_652);
nor U1072 (N_1072,N_106,N_956);
and U1073 (N_1073,N_791,N_513);
and U1074 (N_1074,N_827,N_999);
or U1075 (N_1075,N_764,N_28);
and U1076 (N_1076,N_587,N_330);
and U1077 (N_1077,N_227,N_535);
nand U1078 (N_1078,N_895,N_125);
nor U1079 (N_1079,N_819,N_342);
or U1080 (N_1080,N_696,N_625);
nor U1081 (N_1081,N_692,N_919);
and U1082 (N_1082,N_53,N_278);
and U1083 (N_1083,N_729,N_768);
and U1084 (N_1084,N_788,N_309);
nor U1085 (N_1085,N_405,N_704);
and U1086 (N_1086,N_9,N_884);
nand U1087 (N_1087,N_70,N_50);
or U1088 (N_1088,N_253,N_109);
nor U1089 (N_1089,N_850,N_226);
and U1090 (N_1090,N_344,N_987);
and U1091 (N_1091,N_105,N_218);
nand U1092 (N_1092,N_291,N_675);
and U1093 (N_1093,N_923,N_721);
or U1094 (N_1094,N_224,N_98);
or U1095 (N_1095,N_991,N_172);
and U1096 (N_1096,N_369,N_701);
nor U1097 (N_1097,N_30,N_541);
and U1098 (N_1098,N_616,N_897);
and U1099 (N_1099,N_399,N_727);
and U1100 (N_1100,N_942,N_998);
nor U1101 (N_1101,N_136,N_841);
and U1102 (N_1102,N_14,N_1);
and U1103 (N_1103,N_154,N_602);
or U1104 (N_1104,N_447,N_688);
nor U1105 (N_1105,N_258,N_846);
nor U1106 (N_1106,N_458,N_752);
nand U1107 (N_1107,N_893,N_630);
nand U1108 (N_1108,N_983,N_343);
nand U1109 (N_1109,N_129,N_910);
xnor U1110 (N_1110,N_724,N_657);
and U1111 (N_1111,N_124,N_256);
nor U1112 (N_1112,N_210,N_911);
and U1113 (N_1113,N_502,N_909);
or U1114 (N_1114,N_146,N_522);
nor U1115 (N_1115,N_953,N_687);
nor U1116 (N_1116,N_779,N_391);
nand U1117 (N_1117,N_155,N_989);
nand U1118 (N_1118,N_660,N_252);
and U1119 (N_1119,N_478,N_604);
or U1120 (N_1120,N_322,N_977);
or U1121 (N_1121,N_7,N_144);
or U1122 (N_1122,N_951,N_706);
nand U1123 (N_1123,N_529,N_496);
and U1124 (N_1124,N_755,N_548);
nor U1125 (N_1125,N_904,N_712);
and U1126 (N_1126,N_181,N_26);
nand U1127 (N_1127,N_874,N_605);
or U1128 (N_1128,N_305,N_800);
or U1129 (N_1129,N_0,N_45);
nand U1130 (N_1130,N_912,N_537);
or U1131 (N_1131,N_212,N_609);
or U1132 (N_1132,N_272,N_471);
or U1133 (N_1133,N_838,N_812);
nor U1134 (N_1134,N_198,N_737);
nor U1135 (N_1135,N_662,N_482);
nand U1136 (N_1136,N_351,N_333);
nand U1137 (N_1137,N_43,N_607);
or U1138 (N_1138,N_697,N_163);
and U1139 (N_1139,N_174,N_646);
nand U1140 (N_1140,N_949,N_323);
and U1141 (N_1141,N_65,N_444);
and U1142 (N_1142,N_792,N_509);
nand U1143 (N_1143,N_334,N_59);
nor U1144 (N_1144,N_894,N_759);
or U1145 (N_1145,N_859,N_931);
nor U1146 (N_1146,N_68,N_12);
and U1147 (N_1147,N_598,N_813);
and U1148 (N_1148,N_733,N_554);
and U1149 (N_1149,N_306,N_466);
and U1150 (N_1150,N_862,N_944);
nand U1151 (N_1151,N_864,N_339);
nor U1152 (N_1152,N_997,N_489);
and U1153 (N_1153,N_901,N_261);
and U1154 (N_1154,N_698,N_595);
and U1155 (N_1155,N_571,N_373);
and U1156 (N_1156,N_769,N_519);
nand U1157 (N_1157,N_915,N_319);
nor U1158 (N_1158,N_487,N_21);
nand U1159 (N_1159,N_279,N_990);
nand U1160 (N_1160,N_345,N_640);
nand U1161 (N_1161,N_484,N_938);
nand U1162 (N_1162,N_639,N_358);
nand U1163 (N_1163,N_966,N_219);
nor U1164 (N_1164,N_429,N_797);
and U1165 (N_1165,N_99,N_980);
and U1166 (N_1166,N_863,N_963);
or U1167 (N_1167,N_230,N_873);
or U1168 (N_1168,N_336,N_782);
nor U1169 (N_1169,N_31,N_158);
nor U1170 (N_1170,N_528,N_374);
nand U1171 (N_1171,N_961,N_540);
or U1172 (N_1172,N_580,N_442);
nand U1173 (N_1173,N_95,N_524);
nand U1174 (N_1174,N_673,N_265);
nor U1175 (N_1175,N_728,N_689);
nand U1176 (N_1176,N_377,N_669);
or U1177 (N_1177,N_209,N_254);
or U1178 (N_1178,N_842,N_423);
nor U1179 (N_1179,N_267,N_375);
and U1180 (N_1180,N_97,N_833);
nand U1181 (N_1181,N_744,N_981);
or U1182 (N_1182,N_10,N_214);
nor U1183 (N_1183,N_876,N_947);
nand U1184 (N_1184,N_512,N_780);
nor U1185 (N_1185,N_266,N_352);
nand U1186 (N_1186,N_292,N_488);
nor U1187 (N_1187,N_536,N_116);
nor U1188 (N_1188,N_921,N_854);
and U1189 (N_1189,N_865,N_395);
nand U1190 (N_1190,N_244,N_887);
and U1191 (N_1191,N_257,N_828);
nor U1192 (N_1192,N_285,N_681);
nand U1193 (N_1193,N_325,N_679);
nand U1194 (N_1194,N_167,N_126);
nand U1195 (N_1195,N_462,N_475);
nand U1196 (N_1196,N_808,N_208);
and U1197 (N_1197,N_449,N_288);
or U1198 (N_1198,N_734,N_582);
nand U1199 (N_1199,N_470,N_783);
nand U1200 (N_1200,N_241,N_972);
or U1201 (N_1201,N_653,N_937);
or U1202 (N_1202,N_145,N_445);
nor U1203 (N_1203,N_326,N_695);
nand U1204 (N_1204,N_713,N_191);
and U1205 (N_1205,N_479,N_52);
nor U1206 (N_1206,N_871,N_955);
and U1207 (N_1207,N_119,N_468);
nand U1208 (N_1208,N_166,N_816);
xnor U1209 (N_1209,N_366,N_970);
nand U1210 (N_1210,N_815,N_51);
and U1211 (N_1211,N_263,N_579);
and U1212 (N_1212,N_425,N_312);
nand U1213 (N_1213,N_81,N_565);
nor U1214 (N_1214,N_157,N_730);
and U1215 (N_1215,N_401,N_459);
and U1216 (N_1216,N_234,N_597);
or U1217 (N_1217,N_853,N_231);
nor U1218 (N_1218,N_670,N_275);
nor U1219 (N_1219,N_754,N_624);
nor U1220 (N_1220,N_592,N_647);
nor U1221 (N_1221,N_421,N_34);
and U1222 (N_1222,N_933,N_852);
nor U1223 (N_1223,N_469,N_386);
xor U1224 (N_1224,N_349,N_331);
and U1225 (N_1225,N_974,N_413);
nor U1226 (N_1226,N_986,N_515);
and U1227 (N_1227,N_294,N_236);
nand U1228 (N_1228,N_223,N_318);
or U1229 (N_1229,N_232,N_781);
and U1230 (N_1230,N_141,N_184);
or U1231 (N_1231,N_650,N_969);
nand U1232 (N_1232,N_690,N_44);
nand U1233 (N_1233,N_464,N_72);
nand U1234 (N_1234,N_907,N_608);
nor U1235 (N_1235,N_932,N_682);
and U1236 (N_1236,N_329,N_839);
nand U1237 (N_1237,N_775,N_222);
xnor U1238 (N_1238,N_709,N_821);
nand U1239 (N_1239,N_483,N_844);
nand U1240 (N_1240,N_631,N_656);
or U1241 (N_1241,N_620,N_883);
and U1242 (N_1242,N_908,N_108);
nor U1243 (N_1243,N_102,N_557);
or U1244 (N_1244,N_586,N_900);
or U1245 (N_1245,N_988,N_217);
and U1246 (N_1246,N_42,N_648);
or U1247 (N_1247,N_360,N_770);
nor U1248 (N_1248,N_76,N_80);
nand U1249 (N_1249,N_490,N_359);
or U1250 (N_1250,N_622,N_501);
nor U1251 (N_1251,N_307,N_192);
nand U1252 (N_1252,N_927,N_680);
nor U1253 (N_1253,N_477,N_248);
nor U1254 (N_1254,N_530,N_170);
nand U1255 (N_1255,N_240,N_371);
or U1256 (N_1256,N_411,N_651);
and U1257 (N_1257,N_869,N_215);
nor U1258 (N_1258,N_649,N_380);
or U1259 (N_1259,N_262,N_585);
nand U1260 (N_1260,N_247,N_671);
nor U1261 (N_1261,N_100,N_3);
or U1262 (N_1262,N_532,N_793);
nor U1263 (N_1263,N_118,N_694);
or U1264 (N_1264,N_658,N_531);
nor U1265 (N_1265,N_313,N_542);
or U1266 (N_1266,N_593,N_962);
or U1267 (N_1267,N_629,N_25);
nor U1268 (N_1268,N_845,N_250);
or U1269 (N_1269,N_387,N_771);
nor U1270 (N_1270,N_736,N_643);
or U1271 (N_1271,N_934,N_511);
nor U1272 (N_1272,N_686,N_474);
nor U1273 (N_1273,N_190,N_569);
nor U1274 (N_1274,N_514,N_40);
nand U1275 (N_1275,N_891,N_824);
xor U1276 (N_1276,N_161,N_946);
nand U1277 (N_1277,N_603,N_115);
or U1278 (N_1278,N_159,N_807);
or U1279 (N_1279,N_994,N_820);
nor U1280 (N_1280,N_187,N_110);
or U1281 (N_1281,N_799,N_700);
and U1282 (N_1282,N_11,N_112);
or U1283 (N_1283,N_935,N_422);
and U1284 (N_1284,N_601,N_903);
or U1285 (N_1285,N_551,N_617);
and U1286 (N_1286,N_282,N_750);
and U1287 (N_1287,N_8,N_148);
and U1288 (N_1288,N_460,N_5);
nand U1289 (N_1289,N_665,N_971);
nand U1290 (N_1290,N_281,N_301);
nor U1291 (N_1291,N_36,N_787);
nand U1292 (N_1292,N_24,N_73);
xor U1293 (N_1293,N_117,N_928);
nand U1294 (N_1294,N_594,N_806);
nand U1295 (N_1295,N_534,N_777);
and U1296 (N_1296,N_549,N_48);
or U1297 (N_1297,N_703,N_982);
or U1298 (N_1298,N_394,N_924);
nor U1299 (N_1299,N_661,N_726);
nor U1300 (N_1300,N_725,N_418);
or U1301 (N_1301,N_801,N_984);
nor U1302 (N_1302,N_431,N_199);
or U1303 (N_1303,N_577,N_152);
nand U1304 (N_1304,N_714,N_382);
and U1305 (N_1305,N_185,N_389);
nand U1306 (N_1306,N_965,N_563);
nand U1307 (N_1307,N_882,N_438);
and U1308 (N_1308,N_104,N_454);
or U1309 (N_1309,N_615,N_426);
nand U1310 (N_1310,N_967,N_773);
or U1311 (N_1311,N_881,N_836);
nor U1312 (N_1312,N_518,N_547);
nor U1313 (N_1313,N_663,N_60);
nor U1314 (N_1314,N_684,N_950);
or U1315 (N_1315,N_397,N_610);
and U1316 (N_1316,N_455,N_450);
and U1317 (N_1317,N_314,N_361);
or U1318 (N_1318,N_378,N_324);
and U1319 (N_1319,N_428,N_525);
and U1320 (N_1320,N_290,N_38);
nor U1321 (N_1321,N_180,N_90);
nand U1322 (N_1322,N_91,N_875);
and U1323 (N_1323,N_107,N_738);
nand U1324 (N_1324,N_481,N_716);
nand U1325 (N_1325,N_74,N_763);
nor U1326 (N_1326,N_861,N_825);
or U1327 (N_1327,N_635,N_131);
nor U1328 (N_1328,N_85,N_127);
xnor U1329 (N_1329,N_642,N_645);
nor U1330 (N_1330,N_552,N_718);
and U1331 (N_1331,N_930,N_173);
or U1332 (N_1332,N_228,N_114);
or U1333 (N_1333,N_299,N_414);
nor U1334 (N_1334,N_396,N_606);
or U1335 (N_1335,N_507,N_851);
nand U1336 (N_1336,N_201,N_321);
nor U1337 (N_1337,N_566,N_533);
nand U1338 (N_1338,N_320,N_590);
or U1339 (N_1339,N_872,N_56);
or U1340 (N_1340,N_840,N_943);
and U1341 (N_1341,N_751,N_311);
and U1342 (N_1342,N_186,N_628);
nand U1343 (N_1343,N_84,N_356);
nand U1344 (N_1344,N_289,N_150);
xnor U1345 (N_1345,N_843,N_456);
nor U1346 (N_1346,N_308,N_355);
nand U1347 (N_1347,N_463,N_567);
or U1348 (N_1348,N_722,N_588);
and U1349 (N_1349,N_143,N_13);
nand U1350 (N_1350,N_137,N_448);
xor U1351 (N_1351,N_15,N_316);
and U1352 (N_1352,N_435,N_268);
or U1353 (N_1353,N_561,N_613);
nand U1354 (N_1354,N_385,N_504);
nand U1355 (N_1355,N_211,N_742);
nand U1356 (N_1356,N_559,N_746);
or U1357 (N_1357,N_558,N_147);
or U1358 (N_1358,N_372,N_749);
and U1359 (N_1359,N_599,N_202);
or U1360 (N_1360,N_151,N_849);
nor U1361 (N_1361,N_899,N_20);
or U1362 (N_1362,N_139,N_433);
and U1363 (N_1363,N_457,N_200);
or U1364 (N_1364,N_664,N_245);
and U1365 (N_1365,N_495,N_473);
or U1366 (N_1366,N_886,N_560);
and U1367 (N_1367,N_975,N_169);
and U1368 (N_1368,N_817,N_437);
xor U1369 (N_1369,N_176,N_286);
and U1370 (N_1370,N_16,N_879);
nand U1371 (N_1371,N_388,N_4);
or U1372 (N_1372,N_235,N_776);
nor U1373 (N_1373,N_546,N_93);
xnor U1374 (N_1374,N_346,N_795);
or U1375 (N_1375,N_87,N_207);
nand U1376 (N_1376,N_758,N_668);
nor U1377 (N_1377,N_757,N_441);
nor U1378 (N_1378,N_499,N_555);
nand U1379 (N_1379,N_370,N_406);
or U1380 (N_1380,N_632,N_877);
nand U1381 (N_1381,N_790,N_765);
nor U1382 (N_1382,N_255,N_364);
and U1383 (N_1383,N_837,N_677);
and U1384 (N_1384,N_753,N_303);
or U1385 (N_1385,N_868,N_280);
nand U1386 (N_1386,N_637,N_747);
nor U1387 (N_1387,N_809,N_138);
nor U1388 (N_1388,N_492,N_954);
nor U1389 (N_1389,N_578,N_274);
nand U1390 (N_1390,N_237,N_835);
nand U1391 (N_1391,N_493,N_510);
xor U1392 (N_1392,N_784,N_353);
or U1393 (N_1393,N_740,N_23);
nand U1394 (N_1394,N_64,N_526);
and U1395 (N_1395,N_29,N_589);
xnor U1396 (N_1396,N_888,N_300);
nand U1397 (N_1397,N_805,N_539);
or U1398 (N_1398,N_168,N_732);
and U1399 (N_1399,N_205,N_766);
nor U1400 (N_1400,N_576,N_506);
nor U1401 (N_1401,N_979,N_189);
nor U1402 (N_1402,N_194,N_424);
nor U1403 (N_1403,N_134,N_128);
or U1404 (N_1404,N_774,N_898);
and U1405 (N_1405,N_277,N_870);
nor U1406 (N_1406,N_27,N_720);
nor U1407 (N_1407,N_71,N_270);
or U1408 (N_1408,N_612,N_193);
or U1409 (N_1409,N_392,N_310);
nor U1410 (N_1410,N_203,N_672);
nand U1411 (N_1411,N_407,N_332);
xor U1412 (N_1412,N_596,N_830);
nand U1413 (N_1413,N_63,N_239);
and U1414 (N_1414,N_867,N_667);
nand U1415 (N_1415,N_57,N_86);
and U1416 (N_1416,N_92,N_229);
and U1417 (N_1417,N_132,N_6);
or U1418 (N_1418,N_337,N_271);
or U1419 (N_1419,N_140,N_260);
nor U1420 (N_1420,N_32,N_500);
or U1421 (N_1421,N_798,N_505);
or U1422 (N_1422,N_69,N_717);
or U1423 (N_1423,N_521,N_347);
and U1424 (N_1424,N_130,N_472);
nor U1425 (N_1425,N_964,N_723);
and U1426 (N_1426,N_384,N_925);
nor U1427 (N_1427,N_929,N_348);
or U1428 (N_1428,N_693,N_878);
or U1429 (N_1429,N_297,N_259);
nand U1430 (N_1430,N_367,N_96);
xor U1431 (N_1431,N_403,N_634);
or U1432 (N_1432,N_242,N_66);
nor U1433 (N_1433,N_917,N_993);
and U1434 (N_1434,N_304,N_890);
and U1435 (N_1435,N_328,N_295);
nor U1436 (N_1436,N_803,N_420);
or U1437 (N_1437,N_122,N_164);
or U1438 (N_1438,N_902,N_461);
or U1439 (N_1439,N_503,N_35);
nor U1440 (N_1440,N_204,N_171);
nor U1441 (N_1441,N_913,N_149);
nand U1442 (N_1442,N_685,N_544);
nand U1443 (N_1443,N_61,N_162);
or U1444 (N_1444,N_195,N_627);
and U1445 (N_1445,N_952,N_683);
or U1446 (N_1446,N_18,N_545);
xnor U1447 (N_1447,N_584,N_402);
nor U1448 (N_1448,N_440,N_789);
nand U1449 (N_1449,N_550,N_761);
nor U1450 (N_1450,N_636,N_142);
nor U1451 (N_1451,N_973,N_748);
or U1452 (N_1452,N_221,N_739);
nor U1453 (N_1453,N_175,N_400);
or U1454 (N_1454,N_39,N_2);
or U1455 (N_1455,N_855,N_711);
nor U1456 (N_1456,N_276,N_600);
and U1457 (N_1457,N_415,N_760);
nand U1458 (N_1458,N_196,N_621);
nor U1459 (N_1459,N_968,N_517);
nor U1460 (N_1460,N_22,N_491);
nor U1461 (N_1461,N_46,N_77);
xor U1462 (N_1462,N_936,N_467);
or U1463 (N_1463,N_880,N_641);
xnor U1464 (N_1464,N_298,N_831);
nand U1465 (N_1465,N_804,N_581);
nand U1466 (N_1466,N_381,N_707);
or U1467 (N_1467,N_654,N_914);
or U1468 (N_1468,N_135,N_101);
nand U1469 (N_1469,N_678,N_564);
nor U1470 (N_1470,N_826,N_708);
nand U1471 (N_1471,N_832,N_785);
and U1472 (N_1472,N_778,N_89);
nand U1473 (N_1473,N_866,N_516);
and U1474 (N_1474,N_676,N_745);
nand U1475 (N_1475,N_818,N_486);
nand U1476 (N_1476,N_338,N_55);
nand U1477 (N_1477,N_416,N_49);
and U1478 (N_1478,N_75,N_439);
and U1479 (N_1479,N_246,N_941);
nor U1480 (N_1480,N_67,N_553);
nor U1481 (N_1481,N_133,N_430);
nor U1482 (N_1482,N_959,N_655);
nor U1483 (N_1483,N_957,N_574);
and U1484 (N_1484,N_767,N_54);
or U1485 (N_1485,N_480,N_666);
and U1486 (N_1486,N_945,N_156);
and U1487 (N_1487,N_220,N_327);
nor U1488 (N_1488,N_856,N_188);
nor U1489 (N_1489,N_497,N_719);
nor U1490 (N_1490,N_892,N_315);
xor U1491 (N_1491,N_810,N_393);
and U1492 (N_1492,N_302,N_906);
or U1493 (N_1493,N_476,N_995);
and U1494 (N_1494,N_225,N_82);
nor U1495 (N_1495,N_794,N_362);
nand U1496 (N_1496,N_179,N_111);
nor U1497 (N_1497,N_383,N_638);
or U1498 (N_1498,N_417,N_419);
or U1499 (N_1499,N_814,N_575);
or U1500 (N_1500,N_883,N_444);
nand U1501 (N_1501,N_430,N_424);
nor U1502 (N_1502,N_630,N_922);
nor U1503 (N_1503,N_634,N_843);
nand U1504 (N_1504,N_231,N_460);
nor U1505 (N_1505,N_913,N_476);
nand U1506 (N_1506,N_955,N_130);
xnor U1507 (N_1507,N_333,N_923);
or U1508 (N_1508,N_676,N_888);
and U1509 (N_1509,N_796,N_350);
and U1510 (N_1510,N_327,N_345);
and U1511 (N_1511,N_656,N_98);
nor U1512 (N_1512,N_97,N_449);
and U1513 (N_1513,N_330,N_947);
or U1514 (N_1514,N_32,N_309);
nor U1515 (N_1515,N_438,N_335);
nor U1516 (N_1516,N_266,N_90);
nand U1517 (N_1517,N_204,N_163);
nor U1518 (N_1518,N_154,N_706);
and U1519 (N_1519,N_105,N_440);
nand U1520 (N_1520,N_705,N_140);
nand U1521 (N_1521,N_642,N_724);
and U1522 (N_1522,N_444,N_531);
nand U1523 (N_1523,N_538,N_918);
nand U1524 (N_1524,N_386,N_280);
nor U1525 (N_1525,N_709,N_574);
nor U1526 (N_1526,N_185,N_595);
nand U1527 (N_1527,N_826,N_530);
and U1528 (N_1528,N_367,N_642);
xnor U1529 (N_1529,N_787,N_635);
and U1530 (N_1530,N_183,N_137);
nor U1531 (N_1531,N_190,N_525);
nor U1532 (N_1532,N_395,N_711);
or U1533 (N_1533,N_619,N_723);
nand U1534 (N_1534,N_437,N_94);
nor U1535 (N_1535,N_606,N_633);
and U1536 (N_1536,N_981,N_314);
nor U1537 (N_1537,N_578,N_808);
and U1538 (N_1538,N_16,N_747);
nand U1539 (N_1539,N_295,N_541);
xnor U1540 (N_1540,N_742,N_180);
or U1541 (N_1541,N_769,N_848);
nor U1542 (N_1542,N_631,N_161);
or U1543 (N_1543,N_990,N_78);
nor U1544 (N_1544,N_888,N_590);
or U1545 (N_1545,N_314,N_265);
or U1546 (N_1546,N_128,N_757);
or U1547 (N_1547,N_963,N_765);
nand U1548 (N_1548,N_373,N_190);
nand U1549 (N_1549,N_166,N_139);
and U1550 (N_1550,N_331,N_100);
or U1551 (N_1551,N_115,N_236);
nor U1552 (N_1552,N_594,N_207);
or U1553 (N_1553,N_487,N_500);
and U1554 (N_1554,N_322,N_243);
and U1555 (N_1555,N_817,N_579);
or U1556 (N_1556,N_231,N_141);
or U1557 (N_1557,N_940,N_62);
nor U1558 (N_1558,N_688,N_363);
nor U1559 (N_1559,N_9,N_325);
nor U1560 (N_1560,N_710,N_625);
or U1561 (N_1561,N_398,N_699);
nand U1562 (N_1562,N_369,N_898);
nand U1563 (N_1563,N_519,N_912);
nand U1564 (N_1564,N_220,N_443);
and U1565 (N_1565,N_137,N_389);
and U1566 (N_1566,N_930,N_931);
or U1567 (N_1567,N_691,N_786);
and U1568 (N_1568,N_734,N_43);
nand U1569 (N_1569,N_259,N_798);
and U1570 (N_1570,N_372,N_98);
or U1571 (N_1571,N_316,N_664);
or U1572 (N_1572,N_594,N_479);
nand U1573 (N_1573,N_12,N_73);
and U1574 (N_1574,N_764,N_68);
xnor U1575 (N_1575,N_991,N_443);
and U1576 (N_1576,N_864,N_486);
nor U1577 (N_1577,N_347,N_451);
and U1578 (N_1578,N_380,N_206);
nor U1579 (N_1579,N_480,N_359);
or U1580 (N_1580,N_662,N_373);
nand U1581 (N_1581,N_68,N_415);
and U1582 (N_1582,N_788,N_209);
nand U1583 (N_1583,N_774,N_67);
and U1584 (N_1584,N_325,N_426);
nand U1585 (N_1585,N_516,N_468);
or U1586 (N_1586,N_624,N_880);
or U1587 (N_1587,N_214,N_747);
and U1588 (N_1588,N_998,N_425);
and U1589 (N_1589,N_923,N_360);
and U1590 (N_1590,N_152,N_830);
and U1591 (N_1591,N_9,N_871);
nand U1592 (N_1592,N_337,N_101);
and U1593 (N_1593,N_272,N_433);
nand U1594 (N_1594,N_767,N_444);
or U1595 (N_1595,N_278,N_617);
nand U1596 (N_1596,N_597,N_376);
nand U1597 (N_1597,N_398,N_430);
and U1598 (N_1598,N_588,N_522);
nand U1599 (N_1599,N_778,N_186);
nand U1600 (N_1600,N_996,N_948);
nand U1601 (N_1601,N_302,N_951);
nand U1602 (N_1602,N_630,N_933);
and U1603 (N_1603,N_354,N_82);
nor U1604 (N_1604,N_64,N_740);
nor U1605 (N_1605,N_816,N_4);
nand U1606 (N_1606,N_606,N_533);
or U1607 (N_1607,N_261,N_250);
or U1608 (N_1608,N_527,N_209);
or U1609 (N_1609,N_632,N_847);
and U1610 (N_1610,N_397,N_899);
or U1611 (N_1611,N_603,N_225);
nand U1612 (N_1612,N_978,N_424);
nor U1613 (N_1613,N_465,N_723);
and U1614 (N_1614,N_679,N_563);
or U1615 (N_1615,N_680,N_286);
or U1616 (N_1616,N_717,N_914);
nand U1617 (N_1617,N_0,N_135);
or U1618 (N_1618,N_845,N_412);
nand U1619 (N_1619,N_753,N_920);
and U1620 (N_1620,N_323,N_544);
nor U1621 (N_1621,N_643,N_481);
nor U1622 (N_1622,N_969,N_928);
nand U1623 (N_1623,N_170,N_754);
nand U1624 (N_1624,N_727,N_486);
or U1625 (N_1625,N_270,N_503);
or U1626 (N_1626,N_400,N_549);
nor U1627 (N_1627,N_637,N_912);
nor U1628 (N_1628,N_876,N_964);
or U1629 (N_1629,N_131,N_517);
nand U1630 (N_1630,N_78,N_853);
and U1631 (N_1631,N_846,N_406);
and U1632 (N_1632,N_135,N_275);
nand U1633 (N_1633,N_125,N_487);
and U1634 (N_1634,N_336,N_855);
nor U1635 (N_1635,N_598,N_906);
nand U1636 (N_1636,N_9,N_393);
or U1637 (N_1637,N_942,N_554);
or U1638 (N_1638,N_944,N_48);
and U1639 (N_1639,N_752,N_321);
or U1640 (N_1640,N_476,N_761);
nand U1641 (N_1641,N_434,N_290);
nand U1642 (N_1642,N_208,N_845);
nor U1643 (N_1643,N_96,N_282);
or U1644 (N_1644,N_627,N_33);
or U1645 (N_1645,N_963,N_290);
nor U1646 (N_1646,N_658,N_651);
and U1647 (N_1647,N_737,N_972);
or U1648 (N_1648,N_387,N_689);
nor U1649 (N_1649,N_189,N_799);
nor U1650 (N_1650,N_455,N_983);
nor U1651 (N_1651,N_497,N_75);
or U1652 (N_1652,N_543,N_288);
nand U1653 (N_1653,N_48,N_156);
nor U1654 (N_1654,N_738,N_675);
and U1655 (N_1655,N_631,N_854);
nor U1656 (N_1656,N_512,N_697);
and U1657 (N_1657,N_707,N_760);
or U1658 (N_1658,N_210,N_251);
nand U1659 (N_1659,N_618,N_608);
or U1660 (N_1660,N_389,N_974);
xor U1661 (N_1661,N_278,N_204);
nor U1662 (N_1662,N_404,N_447);
or U1663 (N_1663,N_465,N_868);
nand U1664 (N_1664,N_638,N_946);
nand U1665 (N_1665,N_0,N_548);
or U1666 (N_1666,N_344,N_995);
and U1667 (N_1667,N_267,N_134);
and U1668 (N_1668,N_178,N_108);
xnor U1669 (N_1669,N_866,N_179);
nor U1670 (N_1670,N_33,N_206);
nor U1671 (N_1671,N_335,N_449);
nand U1672 (N_1672,N_299,N_335);
nand U1673 (N_1673,N_128,N_18);
xor U1674 (N_1674,N_250,N_608);
nand U1675 (N_1675,N_626,N_797);
nand U1676 (N_1676,N_737,N_538);
nand U1677 (N_1677,N_136,N_101);
and U1678 (N_1678,N_949,N_733);
nor U1679 (N_1679,N_584,N_301);
and U1680 (N_1680,N_534,N_328);
nor U1681 (N_1681,N_178,N_430);
and U1682 (N_1682,N_786,N_764);
and U1683 (N_1683,N_855,N_752);
or U1684 (N_1684,N_749,N_330);
nand U1685 (N_1685,N_26,N_868);
nand U1686 (N_1686,N_4,N_5);
or U1687 (N_1687,N_635,N_461);
nand U1688 (N_1688,N_77,N_398);
nand U1689 (N_1689,N_996,N_726);
nand U1690 (N_1690,N_936,N_19);
and U1691 (N_1691,N_815,N_248);
nand U1692 (N_1692,N_642,N_228);
nand U1693 (N_1693,N_925,N_934);
nor U1694 (N_1694,N_596,N_760);
nor U1695 (N_1695,N_974,N_725);
nor U1696 (N_1696,N_16,N_827);
nand U1697 (N_1697,N_485,N_919);
xor U1698 (N_1698,N_831,N_350);
nor U1699 (N_1699,N_319,N_745);
nor U1700 (N_1700,N_32,N_958);
nor U1701 (N_1701,N_495,N_319);
xnor U1702 (N_1702,N_760,N_19);
nand U1703 (N_1703,N_829,N_790);
and U1704 (N_1704,N_433,N_553);
nor U1705 (N_1705,N_324,N_546);
or U1706 (N_1706,N_635,N_566);
xnor U1707 (N_1707,N_21,N_294);
and U1708 (N_1708,N_905,N_300);
nand U1709 (N_1709,N_784,N_633);
or U1710 (N_1710,N_35,N_398);
or U1711 (N_1711,N_503,N_128);
or U1712 (N_1712,N_941,N_732);
or U1713 (N_1713,N_427,N_876);
or U1714 (N_1714,N_103,N_185);
or U1715 (N_1715,N_296,N_961);
and U1716 (N_1716,N_284,N_447);
or U1717 (N_1717,N_774,N_433);
nand U1718 (N_1718,N_858,N_900);
and U1719 (N_1719,N_877,N_508);
nand U1720 (N_1720,N_133,N_502);
nor U1721 (N_1721,N_220,N_473);
nand U1722 (N_1722,N_24,N_887);
nand U1723 (N_1723,N_41,N_370);
nor U1724 (N_1724,N_519,N_285);
and U1725 (N_1725,N_701,N_360);
and U1726 (N_1726,N_89,N_357);
and U1727 (N_1727,N_570,N_984);
or U1728 (N_1728,N_912,N_826);
nand U1729 (N_1729,N_679,N_183);
or U1730 (N_1730,N_91,N_659);
xnor U1731 (N_1731,N_19,N_733);
or U1732 (N_1732,N_769,N_853);
nor U1733 (N_1733,N_831,N_961);
or U1734 (N_1734,N_483,N_428);
nor U1735 (N_1735,N_826,N_993);
nand U1736 (N_1736,N_76,N_83);
or U1737 (N_1737,N_626,N_590);
or U1738 (N_1738,N_307,N_696);
and U1739 (N_1739,N_280,N_168);
nand U1740 (N_1740,N_440,N_269);
and U1741 (N_1741,N_508,N_810);
or U1742 (N_1742,N_574,N_328);
nor U1743 (N_1743,N_378,N_155);
and U1744 (N_1744,N_411,N_607);
and U1745 (N_1745,N_915,N_808);
and U1746 (N_1746,N_996,N_616);
nand U1747 (N_1747,N_674,N_510);
and U1748 (N_1748,N_811,N_11);
or U1749 (N_1749,N_38,N_604);
nand U1750 (N_1750,N_249,N_872);
and U1751 (N_1751,N_588,N_347);
or U1752 (N_1752,N_791,N_575);
or U1753 (N_1753,N_201,N_796);
or U1754 (N_1754,N_509,N_209);
and U1755 (N_1755,N_540,N_386);
or U1756 (N_1756,N_312,N_449);
and U1757 (N_1757,N_576,N_465);
nand U1758 (N_1758,N_542,N_695);
nand U1759 (N_1759,N_729,N_120);
nand U1760 (N_1760,N_963,N_165);
xor U1761 (N_1761,N_373,N_342);
nor U1762 (N_1762,N_825,N_731);
nor U1763 (N_1763,N_686,N_662);
and U1764 (N_1764,N_982,N_741);
nand U1765 (N_1765,N_150,N_661);
nand U1766 (N_1766,N_856,N_515);
nand U1767 (N_1767,N_468,N_505);
and U1768 (N_1768,N_862,N_688);
nand U1769 (N_1769,N_940,N_594);
or U1770 (N_1770,N_639,N_628);
or U1771 (N_1771,N_402,N_575);
or U1772 (N_1772,N_458,N_150);
nor U1773 (N_1773,N_523,N_164);
and U1774 (N_1774,N_568,N_753);
or U1775 (N_1775,N_763,N_544);
nand U1776 (N_1776,N_490,N_615);
or U1777 (N_1777,N_699,N_487);
or U1778 (N_1778,N_324,N_8);
and U1779 (N_1779,N_932,N_793);
and U1780 (N_1780,N_171,N_127);
or U1781 (N_1781,N_676,N_559);
nor U1782 (N_1782,N_987,N_369);
and U1783 (N_1783,N_452,N_246);
nor U1784 (N_1784,N_621,N_847);
nor U1785 (N_1785,N_530,N_620);
xnor U1786 (N_1786,N_739,N_780);
and U1787 (N_1787,N_918,N_594);
and U1788 (N_1788,N_415,N_101);
nand U1789 (N_1789,N_425,N_207);
and U1790 (N_1790,N_121,N_549);
nor U1791 (N_1791,N_560,N_140);
and U1792 (N_1792,N_813,N_359);
xor U1793 (N_1793,N_376,N_981);
nand U1794 (N_1794,N_748,N_366);
or U1795 (N_1795,N_115,N_69);
or U1796 (N_1796,N_581,N_913);
nor U1797 (N_1797,N_140,N_982);
nor U1798 (N_1798,N_932,N_421);
nand U1799 (N_1799,N_538,N_966);
nand U1800 (N_1800,N_582,N_437);
and U1801 (N_1801,N_483,N_733);
or U1802 (N_1802,N_206,N_706);
or U1803 (N_1803,N_504,N_891);
or U1804 (N_1804,N_660,N_300);
and U1805 (N_1805,N_57,N_114);
nor U1806 (N_1806,N_847,N_534);
and U1807 (N_1807,N_713,N_750);
and U1808 (N_1808,N_998,N_224);
nor U1809 (N_1809,N_163,N_461);
or U1810 (N_1810,N_696,N_102);
nor U1811 (N_1811,N_380,N_304);
or U1812 (N_1812,N_386,N_153);
or U1813 (N_1813,N_205,N_955);
nand U1814 (N_1814,N_402,N_629);
nor U1815 (N_1815,N_633,N_219);
nor U1816 (N_1816,N_440,N_10);
nand U1817 (N_1817,N_914,N_204);
or U1818 (N_1818,N_165,N_848);
nor U1819 (N_1819,N_875,N_19);
or U1820 (N_1820,N_369,N_707);
nand U1821 (N_1821,N_622,N_779);
and U1822 (N_1822,N_954,N_808);
or U1823 (N_1823,N_719,N_430);
or U1824 (N_1824,N_509,N_775);
or U1825 (N_1825,N_802,N_250);
nand U1826 (N_1826,N_132,N_759);
nand U1827 (N_1827,N_691,N_505);
nand U1828 (N_1828,N_290,N_128);
nand U1829 (N_1829,N_170,N_549);
and U1830 (N_1830,N_56,N_969);
nand U1831 (N_1831,N_991,N_688);
nand U1832 (N_1832,N_674,N_293);
nand U1833 (N_1833,N_854,N_806);
or U1834 (N_1834,N_962,N_537);
and U1835 (N_1835,N_496,N_872);
and U1836 (N_1836,N_139,N_406);
nor U1837 (N_1837,N_638,N_360);
and U1838 (N_1838,N_480,N_540);
and U1839 (N_1839,N_919,N_443);
and U1840 (N_1840,N_486,N_940);
and U1841 (N_1841,N_327,N_88);
nor U1842 (N_1842,N_640,N_903);
and U1843 (N_1843,N_903,N_305);
nor U1844 (N_1844,N_132,N_847);
nand U1845 (N_1845,N_110,N_643);
or U1846 (N_1846,N_220,N_10);
nor U1847 (N_1847,N_147,N_970);
or U1848 (N_1848,N_888,N_650);
and U1849 (N_1849,N_370,N_929);
and U1850 (N_1850,N_60,N_736);
nor U1851 (N_1851,N_949,N_191);
nand U1852 (N_1852,N_382,N_428);
nor U1853 (N_1853,N_881,N_550);
or U1854 (N_1854,N_204,N_207);
and U1855 (N_1855,N_17,N_384);
nand U1856 (N_1856,N_632,N_892);
nor U1857 (N_1857,N_265,N_753);
or U1858 (N_1858,N_894,N_939);
nor U1859 (N_1859,N_389,N_412);
xor U1860 (N_1860,N_706,N_303);
nor U1861 (N_1861,N_61,N_641);
nor U1862 (N_1862,N_972,N_184);
nand U1863 (N_1863,N_0,N_232);
and U1864 (N_1864,N_765,N_96);
nand U1865 (N_1865,N_178,N_964);
nand U1866 (N_1866,N_246,N_336);
nor U1867 (N_1867,N_239,N_667);
nand U1868 (N_1868,N_367,N_296);
nor U1869 (N_1869,N_55,N_3);
nor U1870 (N_1870,N_980,N_2);
and U1871 (N_1871,N_729,N_232);
nor U1872 (N_1872,N_237,N_771);
or U1873 (N_1873,N_198,N_695);
and U1874 (N_1874,N_169,N_953);
and U1875 (N_1875,N_576,N_877);
nor U1876 (N_1876,N_340,N_699);
nor U1877 (N_1877,N_268,N_833);
xor U1878 (N_1878,N_833,N_365);
and U1879 (N_1879,N_327,N_724);
and U1880 (N_1880,N_849,N_407);
nor U1881 (N_1881,N_497,N_306);
nand U1882 (N_1882,N_461,N_927);
or U1883 (N_1883,N_661,N_487);
nand U1884 (N_1884,N_988,N_334);
nor U1885 (N_1885,N_362,N_525);
and U1886 (N_1886,N_156,N_799);
or U1887 (N_1887,N_851,N_469);
xnor U1888 (N_1888,N_867,N_502);
nor U1889 (N_1889,N_678,N_411);
nor U1890 (N_1890,N_200,N_109);
and U1891 (N_1891,N_940,N_493);
and U1892 (N_1892,N_378,N_322);
and U1893 (N_1893,N_960,N_341);
and U1894 (N_1894,N_578,N_621);
or U1895 (N_1895,N_768,N_586);
nand U1896 (N_1896,N_618,N_936);
or U1897 (N_1897,N_802,N_514);
nand U1898 (N_1898,N_747,N_967);
nor U1899 (N_1899,N_341,N_256);
nand U1900 (N_1900,N_860,N_522);
nand U1901 (N_1901,N_126,N_516);
or U1902 (N_1902,N_619,N_790);
and U1903 (N_1903,N_746,N_476);
nor U1904 (N_1904,N_605,N_455);
nor U1905 (N_1905,N_351,N_22);
or U1906 (N_1906,N_972,N_271);
and U1907 (N_1907,N_377,N_416);
and U1908 (N_1908,N_941,N_793);
nor U1909 (N_1909,N_552,N_55);
nand U1910 (N_1910,N_763,N_586);
nand U1911 (N_1911,N_202,N_633);
or U1912 (N_1912,N_544,N_320);
nor U1913 (N_1913,N_868,N_439);
nor U1914 (N_1914,N_717,N_949);
and U1915 (N_1915,N_921,N_693);
nand U1916 (N_1916,N_210,N_734);
nand U1917 (N_1917,N_301,N_532);
or U1918 (N_1918,N_549,N_248);
nor U1919 (N_1919,N_245,N_949);
and U1920 (N_1920,N_609,N_915);
or U1921 (N_1921,N_639,N_528);
nor U1922 (N_1922,N_165,N_664);
nor U1923 (N_1923,N_572,N_6);
and U1924 (N_1924,N_502,N_680);
nand U1925 (N_1925,N_890,N_163);
and U1926 (N_1926,N_519,N_517);
and U1927 (N_1927,N_121,N_295);
nand U1928 (N_1928,N_772,N_775);
and U1929 (N_1929,N_573,N_384);
nand U1930 (N_1930,N_2,N_49);
or U1931 (N_1931,N_569,N_363);
and U1932 (N_1932,N_169,N_618);
and U1933 (N_1933,N_228,N_636);
nor U1934 (N_1934,N_905,N_231);
or U1935 (N_1935,N_40,N_5);
nand U1936 (N_1936,N_195,N_441);
nor U1937 (N_1937,N_126,N_72);
nor U1938 (N_1938,N_671,N_821);
or U1939 (N_1939,N_217,N_337);
or U1940 (N_1940,N_476,N_604);
or U1941 (N_1941,N_354,N_844);
nor U1942 (N_1942,N_24,N_329);
and U1943 (N_1943,N_291,N_173);
and U1944 (N_1944,N_780,N_249);
nor U1945 (N_1945,N_395,N_559);
nor U1946 (N_1946,N_448,N_541);
and U1947 (N_1947,N_938,N_431);
or U1948 (N_1948,N_765,N_654);
nor U1949 (N_1949,N_849,N_209);
nor U1950 (N_1950,N_440,N_458);
and U1951 (N_1951,N_787,N_11);
nor U1952 (N_1952,N_717,N_120);
nor U1953 (N_1953,N_612,N_638);
or U1954 (N_1954,N_395,N_787);
xnor U1955 (N_1955,N_43,N_264);
or U1956 (N_1956,N_343,N_552);
and U1957 (N_1957,N_621,N_167);
nand U1958 (N_1958,N_471,N_740);
nor U1959 (N_1959,N_326,N_501);
and U1960 (N_1960,N_712,N_162);
or U1961 (N_1961,N_492,N_723);
and U1962 (N_1962,N_94,N_727);
nand U1963 (N_1963,N_361,N_271);
or U1964 (N_1964,N_665,N_546);
or U1965 (N_1965,N_989,N_740);
or U1966 (N_1966,N_645,N_149);
nand U1967 (N_1967,N_742,N_855);
or U1968 (N_1968,N_769,N_247);
and U1969 (N_1969,N_567,N_496);
nor U1970 (N_1970,N_819,N_869);
nand U1971 (N_1971,N_624,N_456);
or U1972 (N_1972,N_125,N_373);
or U1973 (N_1973,N_179,N_677);
nand U1974 (N_1974,N_102,N_983);
nand U1975 (N_1975,N_552,N_600);
nand U1976 (N_1976,N_136,N_911);
nand U1977 (N_1977,N_462,N_594);
and U1978 (N_1978,N_145,N_297);
nor U1979 (N_1979,N_148,N_984);
or U1980 (N_1980,N_775,N_140);
or U1981 (N_1981,N_632,N_229);
or U1982 (N_1982,N_537,N_853);
or U1983 (N_1983,N_243,N_870);
nand U1984 (N_1984,N_34,N_983);
and U1985 (N_1985,N_924,N_80);
or U1986 (N_1986,N_681,N_16);
and U1987 (N_1987,N_86,N_162);
nor U1988 (N_1988,N_549,N_467);
and U1989 (N_1989,N_887,N_136);
xnor U1990 (N_1990,N_833,N_436);
or U1991 (N_1991,N_310,N_572);
nor U1992 (N_1992,N_867,N_827);
or U1993 (N_1993,N_431,N_151);
and U1994 (N_1994,N_627,N_92);
nor U1995 (N_1995,N_990,N_629);
or U1996 (N_1996,N_338,N_382);
and U1997 (N_1997,N_189,N_221);
nand U1998 (N_1998,N_238,N_922);
xnor U1999 (N_1999,N_361,N_986);
or U2000 (N_2000,N_1044,N_1053);
nor U2001 (N_2001,N_1819,N_1351);
or U2002 (N_2002,N_1847,N_1519);
and U2003 (N_2003,N_1197,N_1945);
and U2004 (N_2004,N_1024,N_1952);
or U2005 (N_2005,N_1811,N_1542);
and U2006 (N_2006,N_1290,N_1975);
or U2007 (N_2007,N_1579,N_1101);
nand U2008 (N_2008,N_1832,N_1442);
nor U2009 (N_2009,N_1453,N_1813);
nand U2010 (N_2010,N_1469,N_1795);
nand U2011 (N_2011,N_1349,N_1054);
and U2012 (N_2012,N_1876,N_1550);
or U2013 (N_2013,N_1438,N_1693);
nand U2014 (N_2014,N_1355,N_1367);
and U2015 (N_2015,N_1696,N_1708);
nor U2016 (N_2016,N_1884,N_1854);
or U2017 (N_2017,N_1386,N_1165);
nor U2018 (N_2018,N_1085,N_1371);
nor U2019 (N_2019,N_1892,N_1436);
nand U2020 (N_2020,N_1041,N_1889);
nor U2021 (N_2021,N_1651,N_1875);
and U2022 (N_2022,N_1957,N_1014);
or U2023 (N_2023,N_1548,N_1790);
xor U2024 (N_2024,N_1152,N_1269);
and U2025 (N_2025,N_1078,N_1585);
or U2026 (N_2026,N_1877,N_1200);
xnor U2027 (N_2027,N_1936,N_1241);
or U2028 (N_2028,N_1799,N_1091);
nand U2029 (N_2029,N_1973,N_1926);
and U2030 (N_2030,N_1285,N_1620);
nor U2031 (N_2031,N_1317,N_1781);
and U2032 (N_2032,N_1681,N_1201);
nor U2033 (N_2033,N_1263,N_1286);
nor U2034 (N_2034,N_1313,N_1746);
nand U2035 (N_2035,N_1028,N_1772);
and U2036 (N_2036,N_1996,N_1223);
xnor U2037 (N_2037,N_1977,N_1938);
and U2038 (N_2038,N_1480,N_1293);
nand U2039 (N_2039,N_1418,N_1424);
nand U2040 (N_2040,N_1803,N_1896);
and U2041 (N_2041,N_1870,N_1100);
and U2042 (N_2042,N_1029,N_1363);
nor U2043 (N_2043,N_1630,N_1648);
or U2044 (N_2044,N_1900,N_1590);
nand U2045 (N_2045,N_1478,N_1955);
or U2046 (N_2046,N_1009,N_1599);
nor U2047 (N_2047,N_1514,N_1976);
or U2048 (N_2048,N_1206,N_1256);
or U2049 (N_2049,N_1879,N_1511);
nand U2050 (N_2050,N_1466,N_1495);
and U2051 (N_2051,N_1916,N_1516);
and U2052 (N_2052,N_1503,N_1737);
nand U2053 (N_2053,N_1616,N_1930);
or U2054 (N_2054,N_1061,N_1712);
or U2055 (N_2055,N_1667,N_1445);
or U2056 (N_2056,N_1229,N_1523);
or U2057 (N_2057,N_1709,N_1244);
nor U2058 (N_2058,N_1485,N_1190);
or U2059 (N_2059,N_1069,N_1914);
nor U2060 (N_2060,N_1164,N_1988);
nor U2061 (N_2061,N_1807,N_1346);
and U2062 (N_2062,N_1268,N_1979);
nor U2063 (N_2063,N_1678,N_1082);
or U2064 (N_2064,N_1287,N_1486);
nand U2065 (N_2065,N_1419,N_1370);
or U2066 (N_2066,N_1236,N_1142);
xnor U2067 (N_2067,N_1198,N_1739);
or U2068 (N_2068,N_1228,N_1350);
nand U2069 (N_2069,N_1182,N_1220);
nand U2070 (N_2070,N_1076,N_1692);
nor U2071 (N_2071,N_1276,N_1720);
or U2072 (N_2072,N_1840,N_1661);
nand U2073 (N_2073,N_1233,N_1272);
and U2074 (N_2074,N_1831,N_1821);
or U2075 (N_2075,N_1217,N_1767);
nand U2076 (N_2076,N_1589,N_1862);
nor U2077 (N_2077,N_1907,N_1302);
nand U2078 (N_2078,N_1534,N_1656);
or U2079 (N_2079,N_1572,N_1869);
or U2080 (N_2080,N_1400,N_1646);
or U2081 (N_2081,N_1898,N_1038);
nand U2082 (N_2082,N_1570,N_1391);
nand U2083 (N_2083,N_1291,N_1405);
and U2084 (N_2084,N_1759,N_1617);
nand U2085 (N_2085,N_1963,N_1348);
and U2086 (N_2086,N_1281,N_1953);
nor U2087 (N_2087,N_1191,N_1556);
nand U2088 (N_2088,N_1360,N_1911);
and U2089 (N_2089,N_1120,N_1275);
or U2090 (N_2090,N_1064,N_1533);
nor U2091 (N_2091,N_1965,N_1747);
and U2092 (N_2092,N_1266,N_1726);
nand U2093 (N_2093,N_1116,N_1499);
or U2094 (N_2094,N_1912,N_1107);
and U2095 (N_2095,N_1493,N_1718);
nor U2096 (N_2096,N_1174,N_1562);
or U2097 (N_2097,N_1384,N_1219);
nand U2098 (N_2098,N_1112,N_1364);
or U2099 (N_2099,N_1212,N_1096);
nor U2100 (N_2100,N_1644,N_1810);
nand U2101 (N_2101,N_1950,N_1307);
or U2102 (N_2102,N_1624,N_1818);
or U2103 (N_2103,N_1923,N_1723);
nand U2104 (N_2104,N_1378,N_1939);
nand U2105 (N_2105,N_1434,N_1049);
nor U2106 (N_2106,N_1595,N_1763);
nor U2107 (N_2107,N_1968,N_1243);
nor U2108 (N_2108,N_1123,N_1702);
nor U2109 (N_2109,N_1608,N_1603);
and U2110 (N_2110,N_1460,N_1619);
nor U2111 (N_2111,N_1093,N_1150);
nor U2112 (N_2112,N_1403,N_1482);
nand U2113 (N_2113,N_1629,N_1551);
nand U2114 (N_2114,N_1594,N_1379);
or U2115 (N_2115,N_1398,N_1213);
nand U2116 (N_2116,N_1373,N_1188);
nor U2117 (N_2117,N_1043,N_1050);
or U2118 (N_2118,N_1447,N_1259);
nand U2119 (N_2119,N_1549,N_1894);
and U2120 (N_2120,N_1372,N_1784);
nand U2121 (N_2121,N_1856,N_1427);
nor U2122 (N_2122,N_1331,N_1871);
or U2123 (N_2123,N_1679,N_1669);
nor U2124 (N_2124,N_1114,N_1411);
xnor U2125 (N_2125,N_1488,N_1714);
and U2126 (N_2126,N_1311,N_1361);
and U2127 (N_2127,N_1340,N_1157);
xor U2128 (N_2128,N_1992,N_1828);
nand U2129 (N_2129,N_1280,N_1689);
nor U2130 (N_2130,N_1566,N_1358);
nand U2131 (N_2131,N_1423,N_1796);
nor U2132 (N_2132,N_1476,N_1637);
and U2133 (N_2133,N_1947,N_1305);
nand U2134 (N_2134,N_1541,N_1262);
or U2135 (N_2135,N_1985,N_1329);
xor U2136 (N_2136,N_1751,N_1867);
or U2137 (N_2137,N_1731,N_1187);
or U2138 (N_2138,N_1033,N_1180);
or U2139 (N_2139,N_1225,N_1941);
nand U2140 (N_2140,N_1322,N_1850);
nand U2141 (N_2141,N_1757,N_1470);
nand U2142 (N_2142,N_1376,N_1897);
and U2143 (N_2143,N_1066,N_1336);
nand U2144 (N_2144,N_1235,N_1011);
nor U2145 (N_2145,N_1834,N_1073);
nor U2146 (N_2146,N_1843,N_1088);
and U2147 (N_2147,N_1068,N_1464);
nand U2148 (N_2148,N_1168,N_1848);
and U2149 (N_2149,N_1902,N_1994);
nor U2150 (N_2150,N_1906,N_1508);
nand U2151 (N_2151,N_1859,N_1804);
nor U2152 (N_2152,N_1226,N_1688);
nor U2153 (N_2153,N_1318,N_1042);
nor U2154 (N_2154,N_1701,N_1295);
nor U2155 (N_2155,N_1177,N_1413);
nand U2156 (N_2156,N_1397,N_1539);
nand U2157 (N_2157,N_1904,N_1131);
and U2158 (N_2158,N_1124,N_1761);
nor U2159 (N_2159,N_1115,N_1341);
xnor U2160 (N_2160,N_1421,N_1760);
and U2161 (N_2161,N_1145,N_1734);
nand U2162 (N_2162,N_1582,N_1929);
nand U2163 (N_2163,N_1059,N_1525);
nand U2164 (N_2164,N_1086,N_1789);
and U2165 (N_2165,N_1048,N_1578);
and U2166 (N_2166,N_1778,N_1303);
nand U2167 (N_2167,N_1113,N_1817);
nor U2168 (N_2168,N_1196,N_1412);
or U2169 (N_2169,N_1079,N_1020);
nor U2170 (N_2170,N_1330,N_1097);
or U2171 (N_2171,N_1672,N_1785);
nand U2172 (N_2172,N_1487,N_1347);
and U2173 (N_2173,N_1312,N_1040);
or U2174 (N_2174,N_1333,N_1597);
or U2175 (N_2175,N_1838,N_1451);
nand U2176 (N_2176,N_1288,N_1027);
and U2177 (N_2177,N_1431,N_1273);
or U2178 (N_2178,N_1687,N_1260);
or U2179 (N_2179,N_1770,N_1366);
nor U2180 (N_2180,N_1297,N_1683);
nor U2181 (N_2181,N_1880,N_1969);
nand U2182 (N_2182,N_1354,N_1051);
nand U2183 (N_2183,N_1045,N_1492);
nand U2184 (N_2184,N_1638,N_1342);
nor U2185 (N_2185,N_1335,N_1927);
and U2186 (N_2186,N_1866,N_1375);
or U2187 (N_2187,N_1163,N_1674);
or U2188 (N_2188,N_1888,N_1522);
nand U2189 (N_2189,N_1855,N_1169);
nand U2190 (N_2190,N_1515,N_1798);
and U2191 (N_2191,N_1561,N_1357);
nor U2192 (N_2192,N_1238,N_1662);
and U2193 (N_2193,N_1129,N_1874);
nor U2194 (N_2194,N_1951,N_1270);
or U2195 (N_2195,N_1388,N_1218);
nand U2196 (N_2196,N_1294,N_1756);
xor U2197 (N_2197,N_1109,N_1748);
or U2198 (N_2198,N_1429,N_1265);
or U2199 (N_2199,N_1711,N_1094);
nand U2200 (N_2200,N_1455,N_1472);
nor U2201 (N_2201,N_1998,N_1016);
and U2202 (N_2202,N_1698,N_1389);
or U2203 (N_2203,N_1791,N_1545);
or U2204 (N_2204,N_1160,N_1697);
nor U2205 (N_2205,N_1841,N_1186);
nor U2206 (N_2206,N_1940,N_1546);
nor U2207 (N_2207,N_1510,N_1520);
or U2208 (N_2208,N_1873,N_1517);
nand U2209 (N_2209,N_1989,N_1035);
nor U2210 (N_2210,N_1494,N_1891);
or U2211 (N_2211,N_1993,N_1530);
nor U2212 (N_2212,N_1845,N_1685);
or U2213 (N_2213,N_1479,N_1394);
and U2214 (N_2214,N_1032,N_1345);
nor U2215 (N_2215,N_1860,N_1105);
nor U2216 (N_2216,N_1553,N_1618);
xnor U2217 (N_2217,N_1733,N_1820);
nand U2218 (N_2218,N_1296,N_1467);
nor U2219 (N_2219,N_1416,N_1095);
and U2220 (N_2220,N_1671,N_1443);
nor U2221 (N_2221,N_1623,N_1893);
nand U2222 (N_2222,N_1576,N_1208);
nand U2223 (N_2223,N_1261,N_1143);
nor U2224 (N_2224,N_1613,N_1161);
nand U2225 (N_2225,N_1321,N_1753);
nand U2226 (N_2226,N_1970,N_1128);
nor U2227 (N_2227,N_1924,N_1966);
or U2228 (N_2228,N_1183,N_1450);
and U2229 (N_2229,N_1359,N_1205);
nand U2230 (N_2230,N_1537,N_1111);
and U2231 (N_2231,N_1980,N_1657);
or U2232 (N_2232,N_1284,N_1247);
and U2233 (N_2233,N_1012,N_1991);
or U2234 (N_2234,N_1019,N_1749);
nor U2235 (N_2235,N_1021,N_1231);
or U2236 (N_2236,N_1323,N_1319);
xnor U2237 (N_2237,N_1155,N_1300);
nand U2238 (N_2238,N_1432,N_1385);
or U2239 (N_2239,N_1636,N_1690);
nor U2240 (N_2240,N_1609,N_1540);
or U2241 (N_2241,N_1090,N_1159);
or U2242 (N_2242,N_1649,N_1563);
nor U2243 (N_2243,N_1583,N_1117);
and U2244 (N_2244,N_1465,N_1369);
nor U2245 (N_2245,N_1250,N_1844);
nor U2246 (N_2246,N_1527,N_1395);
and U2247 (N_2247,N_1812,N_1267);
and U2248 (N_2248,N_1141,N_1658);
nand U2249 (N_2249,N_1308,N_1829);
xor U2250 (N_2250,N_1230,N_1179);
and U2251 (N_2251,N_1954,N_1199);
nor U2252 (N_2252,N_1249,N_1022);
nand U2253 (N_2253,N_1640,N_1399);
nand U2254 (N_2254,N_1611,N_1903);
nor U2255 (N_2255,N_1981,N_1668);
or U2256 (N_2256,N_1846,N_1127);
or U2257 (N_2257,N_1878,N_1513);
nor U2258 (N_2258,N_1118,N_1136);
and U2259 (N_2259,N_1962,N_1343);
nand U2260 (N_2260,N_1007,N_1569);
and U2261 (N_2261,N_1070,N_1207);
nor U2262 (N_2262,N_1650,N_1984);
nor U2263 (N_2263,N_1735,N_1065);
and U2264 (N_2264,N_1299,N_1908);
nor U2265 (N_2265,N_1864,N_1851);
nand U2266 (N_2266,N_1139,N_1377);
or U2267 (N_2267,N_1729,N_1380);
and U2268 (N_2268,N_1417,N_1706);
and U2269 (N_2269,N_1861,N_1822);
nor U2270 (N_2270,N_1383,N_1986);
or U2271 (N_2271,N_1928,N_1289);
or U2272 (N_2272,N_1933,N_1457);
nor U2273 (N_2273,N_1581,N_1214);
nand U2274 (N_2274,N_1635,N_1797);
and U2275 (N_2275,N_1224,N_1507);
nand U2276 (N_2276,N_1532,N_1448);
nor U2277 (N_2277,N_1942,N_1881);
nand U2278 (N_2278,N_1744,N_1792);
or U2279 (N_2279,N_1003,N_1353);
and U2280 (N_2280,N_1304,N_1919);
and U2281 (N_2281,N_1765,N_1144);
and U2282 (N_2282,N_1676,N_1309);
nand U2283 (N_2283,N_1222,N_1175);
and U2284 (N_2284,N_1645,N_1641);
nand U2285 (N_2285,N_1211,N_1584);
and U2286 (N_2286,N_1374,N_1245);
nor U2287 (N_2287,N_1614,N_1036);
and U2288 (N_2288,N_1758,N_1039);
and U2289 (N_2289,N_1588,N_1788);
or U2290 (N_2290,N_1102,N_1937);
nor U2291 (N_2291,N_1728,N_1406);
nand U2292 (N_2292,N_1741,N_1327);
nor U2293 (N_2293,N_1458,N_1382);
or U2294 (N_2294,N_1554,N_1543);
or U2295 (N_2295,N_1501,N_1456);
nor U2296 (N_2296,N_1010,N_1253);
xor U2297 (N_2297,N_1310,N_1762);
nor U2298 (N_2298,N_1887,N_1730);
or U2299 (N_2299,N_1184,N_1913);
nor U2300 (N_2300,N_1257,N_1018);
nor U2301 (N_2301,N_1509,N_1362);
nand U2302 (N_2302,N_1625,N_1555);
nor U2303 (N_2303,N_1704,N_1682);
nand U2304 (N_2304,N_1401,N_1857);
and U2305 (N_2305,N_1826,N_1771);
and U2306 (N_2306,N_1852,N_1837);
nor U2307 (N_2307,N_1793,N_1497);
or U2308 (N_2308,N_1099,N_1428);
nor U2309 (N_2309,N_1529,N_1080);
nor U2310 (N_2310,N_1081,N_1684);
or U2311 (N_2311,N_1596,N_1440);
nor U2312 (N_2312,N_1498,N_1356);
or U2313 (N_2313,N_1865,N_1982);
and U2314 (N_2314,N_1381,N_1087);
nand U2315 (N_2315,N_1568,N_1409);
and U2316 (N_2316,N_1621,N_1337);
nand U2317 (N_2317,N_1622,N_1430);
nand U2318 (N_2318,N_1320,N_1063);
or U2319 (N_2319,N_1536,N_1738);
or U2320 (N_2320,N_1189,N_1769);
nor U2321 (N_2321,N_1387,N_1017);
nand U2322 (N_2322,N_1591,N_1153);
or U2323 (N_2323,N_1454,N_1315);
nand U2324 (N_2324,N_1239,N_1971);
and U2325 (N_2325,N_1232,N_1632);
nor U2326 (N_2326,N_1119,N_1806);
nor U2327 (N_2327,N_1604,N_1481);
xor U2328 (N_2328,N_1148,N_1987);
nor U2329 (N_2329,N_1005,N_1802);
or U2330 (N_2330,N_1248,N_1132);
or U2331 (N_2331,N_1056,N_1827);
and U2332 (N_2332,N_1732,N_1058);
and U2333 (N_2333,N_1452,N_1166);
and U2334 (N_2334,N_1221,N_1176);
and U2335 (N_2335,N_1960,N_1414);
and U2336 (N_2336,N_1754,N_1607);
and U2337 (N_2337,N_1544,N_1890);
or U2338 (N_2338,N_1072,N_1755);
and U2339 (N_2339,N_1743,N_1531);
nand U2340 (N_2340,N_1439,N_1670);
nand U2341 (N_2341,N_1634,N_1943);
or U2342 (N_2342,N_1567,N_1408);
and U2343 (N_2343,N_1060,N_1872);
and U2344 (N_2344,N_1722,N_1396);
nor U2345 (N_2345,N_1326,N_1959);
and U2346 (N_2346,N_1067,N_1736);
nor U2347 (N_2347,N_1106,N_1823);
nand U2348 (N_2348,N_1203,N_1643);
or U2349 (N_2349,N_1918,N_1046);
and U2350 (N_2350,N_1612,N_1512);
or U2351 (N_2351,N_1133,N_1103);
or U2352 (N_2352,N_1282,N_1279);
and U2353 (N_2353,N_1449,N_1610);
or U2354 (N_2354,N_1901,N_1783);
nand U2355 (N_2355,N_1571,N_1505);
and U2356 (N_2356,N_1237,N_1437);
and U2357 (N_2357,N_1057,N_1149);
and U2358 (N_2358,N_1766,N_1008);
and U2359 (N_2359,N_1151,N_1167);
or U2360 (N_2360,N_1292,N_1627);
nor U2361 (N_2361,N_1606,N_1215);
and U2362 (N_2362,N_1277,N_1715);
and U2363 (N_2363,N_1653,N_1666);
nor U2364 (N_2364,N_1518,N_1463);
or U2365 (N_2365,N_1258,N_1949);
and U2366 (N_2366,N_1328,N_1673);
nor U2367 (N_2367,N_1209,N_1780);
and U2368 (N_2368,N_1332,N_1338);
nand U2369 (N_2369,N_1535,N_1974);
nand U2370 (N_2370,N_1573,N_1392);
nor U2371 (N_2371,N_1752,N_1863);
nor U2372 (N_2372,N_1283,N_1999);
nor U2373 (N_2373,N_1252,N_1528);
nand U2374 (N_2374,N_1716,N_1314);
or U2375 (N_2375,N_1663,N_1216);
nor U2376 (N_2376,N_1794,N_1402);
and U2377 (N_2377,N_1393,N_1601);
or U2378 (N_2378,N_1154,N_1325);
nor U2379 (N_2379,N_1602,N_1047);
nor U2380 (N_2380,N_1835,N_1271);
xor U2381 (N_2381,N_1204,N_1628);
xor U2382 (N_2382,N_1475,N_1306);
nand U2383 (N_2383,N_1909,N_1946);
nor U2384 (N_2384,N_1705,N_1592);
or U2385 (N_2385,N_1435,N_1776);
nand U2386 (N_2386,N_1193,N_1564);
or U2387 (N_2387,N_1703,N_1574);
and U2388 (N_2388,N_1830,N_1686);
xor U2389 (N_2389,N_1001,N_1839);
xor U2390 (N_2390,N_1768,N_1426);
nor U2391 (N_2391,N_1425,N_1185);
or U2392 (N_2392,N_1713,N_1967);
nand U2393 (N_2393,N_1171,N_1922);
xor U2394 (N_2394,N_1660,N_1978);
or U2395 (N_2395,N_1246,N_1410);
xnor U2396 (N_2396,N_1883,N_1137);
and U2397 (N_2397,N_1110,N_1098);
or U2398 (N_2398,N_1547,N_1719);
or U2399 (N_2399,N_1725,N_1422);
nor U2400 (N_2400,N_1652,N_1254);
nand U2401 (N_2401,N_1777,N_1524);
and U2402 (N_2402,N_1972,N_1773);
or U2403 (N_2403,N_1474,N_1062);
nor U2404 (N_2404,N_1092,N_1633);
or U2405 (N_2405,N_1575,N_1800);
and U2406 (N_2406,N_1932,N_1782);
or U2407 (N_2407,N_1600,N_1586);
and U2408 (N_2408,N_1565,N_1274);
nor U2409 (N_2409,N_1655,N_1334);
or U2410 (N_2410,N_1147,N_1352);
and U2411 (N_2411,N_1202,N_1931);
or U2412 (N_2412,N_1675,N_1108);
nand U2413 (N_2413,N_1013,N_1496);
and U2414 (N_2414,N_1026,N_1251);
nand U2415 (N_2415,N_1146,N_1779);
nand U2416 (N_2416,N_1178,N_1194);
or U2417 (N_2417,N_1724,N_1015);
nor U2418 (N_2418,N_1695,N_1825);
nand U2419 (N_2419,N_1764,N_1717);
nand U2420 (N_2420,N_1002,N_1089);
nor U2421 (N_2421,N_1631,N_1126);
nand U2422 (N_2422,N_1173,N_1407);
or U2423 (N_2423,N_1506,N_1156);
and U2424 (N_2424,N_1526,N_1234);
nand U2425 (N_2425,N_1801,N_1990);
nor U2426 (N_2426,N_1462,N_1000);
or U2427 (N_2427,N_1071,N_1468);
or U2428 (N_2428,N_1833,N_1004);
nand U2429 (N_2429,N_1025,N_1915);
and U2430 (N_2430,N_1473,N_1593);
or U2431 (N_2431,N_1654,N_1886);
or U2432 (N_2432,N_1134,N_1740);
nand U2433 (N_2433,N_1344,N_1598);
nand U2434 (N_2434,N_1444,N_1895);
nand U2435 (N_2435,N_1404,N_1842);
nor U2436 (N_2436,N_1917,N_1420);
nand U2437 (N_2437,N_1677,N_1944);
nor U2438 (N_2438,N_1242,N_1301);
and U2439 (N_2439,N_1983,N_1459);
nand U2440 (N_2440,N_1727,N_1006);
and U2441 (N_2441,N_1521,N_1316);
and U2442 (N_2442,N_1882,N_1483);
nor U2443 (N_2443,N_1775,N_1034);
nor U2444 (N_2444,N_1680,N_1477);
nand U2445 (N_2445,N_1615,N_1805);
and U2446 (N_2446,N_1023,N_1181);
or U2447 (N_2447,N_1138,N_1490);
nor U2448 (N_2448,N_1084,N_1786);
or U2449 (N_2449,N_1665,N_1433);
nor U2450 (N_2450,N_1774,N_1956);
nand U2451 (N_2451,N_1030,N_1552);
and U2452 (N_2452,N_1560,N_1824);
and U2453 (N_2453,N_1083,N_1809);
xnor U2454 (N_2454,N_1500,N_1037);
nor U2455 (N_2455,N_1122,N_1172);
and U2456 (N_2456,N_1885,N_1240);
nand U2457 (N_2457,N_1707,N_1816);
and U2458 (N_2458,N_1577,N_1721);
nor U2459 (N_2459,N_1557,N_1808);
xor U2460 (N_2460,N_1920,N_1659);
nor U2461 (N_2461,N_1958,N_1639);
nand U2462 (N_2462,N_1647,N_1836);
and U2463 (N_2463,N_1699,N_1750);
nor U2464 (N_2464,N_1264,N_1491);
and U2465 (N_2465,N_1121,N_1997);
and U2466 (N_2466,N_1052,N_1964);
nand U2467 (N_2467,N_1471,N_1125);
nor U2468 (N_2468,N_1899,N_1948);
nand U2469 (N_2469,N_1853,N_1642);
or U2470 (N_2470,N_1787,N_1195);
and U2471 (N_2471,N_1961,N_1227);
nand U2472 (N_2472,N_1055,N_1580);
nand U2473 (N_2473,N_1849,N_1691);
and U2474 (N_2474,N_1130,N_1192);
or U2475 (N_2475,N_1504,N_1605);
xor U2476 (N_2476,N_1745,N_1365);
and U2477 (N_2477,N_1031,N_1868);
and U2478 (N_2478,N_1905,N_1104);
or U2479 (N_2479,N_1484,N_1158);
or U2480 (N_2480,N_1415,N_1935);
nand U2481 (N_2481,N_1489,N_1910);
nand U2482 (N_2482,N_1502,N_1814);
or U2483 (N_2483,N_1559,N_1278);
nand U2484 (N_2484,N_1934,N_1446);
nor U2485 (N_2485,N_1339,N_1441);
or U2486 (N_2486,N_1710,N_1075);
nand U2487 (N_2487,N_1694,N_1390);
nand U2488 (N_2488,N_1815,N_1538);
or U2489 (N_2489,N_1324,N_1558);
and U2490 (N_2490,N_1162,N_1074);
and U2491 (N_2491,N_1858,N_1298);
nand U2492 (N_2492,N_1135,N_1664);
xor U2493 (N_2493,N_1626,N_1587);
nor U2494 (N_2494,N_1170,N_1700);
and U2495 (N_2495,N_1077,N_1140);
nor U2496 (N_2496,N_1921,N_1368);
and U2497 (N_2497,N_1210,N_1461);
or U2498 (N_2498,N_1925,N_1255);
nand U2499 (N_2499,N_1995,N_1742);
nor U2500 (N_2500,N_1516,N_1654);
nor U2501 (N_2501,N_1596,N_1760);
and U2502 (N_2502,N_1252,N_1189);
nor U2503 (N_2503,N_1670,N_1196);
nor U2504 (N_2504,N_1939,N_1202);
and U2505 (N_2505,N_1951,N_1506);
nand U2506 (N_2506,N_1552,N_1682);
nand U2507 (N_2507,N_1032,N_1064);
or U2508 (N_2508,N_1611,N_1403);
xnor U2509 (N_2509,N_1334,N_1177);
nor U2510 (N_2510,N_1422,N_1373);
nand U2511 (N_2511,N_1621,N_1081);
or U2512 (N_2512,N_1559,N_1730);
nor U2513 (N_2513,N_1687,N_1085);
nand U2514 (N_2514,N_1383,N_1901);
and U2515 (N_2515,N_1035,N_1176);
nor U2516 (N_2516,N_1699,N_1157);
nor U2517 (N_2517,N_1432,N_1506);
and U2518 (N_2518,N_1437,N_1957);
or U2519 (N_2519,N_1544,N_1918);
nand U2520 (N_2520,N_1862,N_1702);
nand U2521 (N_2521,N_1408,N_1086);
nor U2522 (N_2522,N_1575,N_1932);
nand U2523 (N_2523,N_1155,N_1951);
xnor U2524 (N_2524,N_1398,N_1396);
and U2525 (N_2525,N_1597,N_1830);
or U2526 (N_2526,N_1453,N_1328);
nand U2527 (N_2527,N_1970,N_1674);
or U2528 (N_2528,N_1981,N_1952);
and U2529 (N_2529,N_1711,N_1349);
nand U2530 (N_2530,N_1348,N_1109);
or U2531 (N_2531,N_1513,N_1642);
nand U2532 (N_2532,N_1936,N_1415);
nand U2533 (N_2533,N_1395,N_1386);
nand U2534 (N_2534,N_1498,N_1749);
or U2535 (N_2535,N_1835,N_1453);
nor U2536 (N_2536,N_1403,N_1318);
nand U2537 (N_2537,N_1787,N_1544);
xor U2538 (N_2538,N_1863,N_1468);
and U2539 (N_2539,N_1317,N_1868);
and U2540 (N_2540,N_1762,N_1236);
nor U2541 (N_2541,N_1437,N_1879);
nor U2542 (N_2542,N_1442,N_1522);
or U2543 (N_2543,N_1550,N_1699);
nand U2544 (N_2544,N_1006,N_1045);
and U2545 (N_2545,N_1479,N_1095);
and U2546 (N_2546,N_1331,N_1312);
and U2547 (N_2547,N_1139,N_1218);
and U2548 (N_2548,N_1504,N_1165);
nor U2549 (N_2549,N_1647,N_1337);
or U2550 (N_2550,N_1640,N_1240);
nand U2551 (N_2551,N_1616,N_1767);
nor U2552 (N_2552,N_1430,N_1649);
nor U2553 (N_2553,N_1726,N_1627);
nor U2554 (N_2554,N_1345,N_1670);
nor U2555 (N_2555,N_1154,N_1228);
and U2556 (N_2556,N_1991,N_1242);
or U2557 (N_2557,N_1148,N_1656);
nand U2558 (N_2558,N_1140,N_1129);
or U2559 (N_2559,N_1296,N_1006);
nand U2560 (N_2560,N_1694,N_1238);
and U2561 (N_2561,N_1850,N_1278);
xor U2562 (N_2562,N_1216,N_1548);
nand U2563 (N_2563,N_1236,N_1761);
or U2564 (N_2564,N_1672,N_1293);
and U2565 (N_2565,N_1730,N_1357);
nor U2566 (N_2566,N_1697,N_1342);
nand U2567 (N_2567,N_1750,N_1093);
or U2568 (N_2568,N_1584,N_1153);
or U2569 (N_2569,N_1010,N_1797);
nand U2570 (N_2570,N_1653,N_1671);
nor U2571 (N_2571,N_1677,N_1402);
nor U2572 (N_2572,N_1621,N_1393);
and U2573 (N_2573,N_1711,N_1787);
nand U2574 (N_2574,N_1161,N_1770);
or U2575 (N_2575,N_1858,N_1382);
nand U2576 (N_2576,N_1567,N_1613);
or U2577 (N_2577,N_1062,N_1470);
or U2578 (N_2578,N_1402,N_1072);
nor U2579 (N_2579,N_1172,N_1475);
or U2580 (N_2580,N_1704,N_1300);
nor U2581 (N_2581,N_1792,N_1716);
and U2582 (N_2582,N_1751,N_1645);
and U2583 (N_2583,N_1819,N_1795);
nand U2584 (N_2584,N_1839,N_1069);
or U2585 (N_2585,N_1552,N_1813);
nand U2586 (N_2586,N_1229,N_1830);
and U2587 (N_2587,N_1676,N_1031);
or U2588 (N_2588,N_1423,N_1814);
and U2589 (N_2589,N_1752,N_1882);
nor U2590 (N_2590,N_1346,N_1695);
and U2591 (N_2591,N_1335,N_1433);
nand U2592 (N_2592,N_1613,N_1976);
xnor U2593 (N_2593,N_1563,N_1307);
and U2594 (N_2594,N_1675,N_1608);
or U2595 (N_2595,N_1474,N_1190);
or U2596 (N_2596,N_1652,N_1870);
and U2597 (N_2597,N_1655,N_1603);
nor U2598 (N_2598,N_1704,N_1224);
or U2599 (N_2599,N_1087,N_1721);
nand U2600 (N_2600,N_1369,N_1297);
or U2601 (N_2601,N_1205,N_1168);
nand U2602 (N_2602,N_1674,N_1015);
nor U2603 (N_2603,N_1570,N_1432);
nor U2604 (N_2604,N_1228,N_1616);
nor U2605 (N_2605,N_1089,N_1324);
nor U2606 (N_2606,N_1050,N_1123);
nand U2607 (N_2607,N_1546,N_1733);
and U2608 (N_2608,N_1146,N_1693);
nor U2609 (N_2609,N_1953,N_1904);
or U2610 (N_2610,N_1827,N_1161);
or U2611 (N_2611,N_1773,N_1829);
nand U2612 (N_2612,N_1146,N_1900);
nand U2613 (N_2613,N_1049,N_1107);
xor U2614 (N_2614,N_1421,N_1379);
or U2615 (N_2615,N_1983,N_1614);
nand U2616 (N_2616,N_1023,N_1736);
nor U2617 (N_2617,N_1634,N_1152);
nand U2618 (N_2618,N_1275,N_1301);
and U2619 (N_2619,N_1403,N_1526);
nor U2620 (N_2620,N_1937,N_1882);
and U2621 (N_2621,N_1734,N_1032);
nor U2622 (N_2622,N_1193,N_1254);
nand U2623 (N_2623,N_1890,N_1163);
nand U2624 (N_2624,N_1313,N_1591);
nor U2625 (N_2625,N_1020,N_1866);
and U2626 (N_2626,N_1599,N_1696);
nand U2627 (N_2627,N_1355,N_1929);
and U2628 (N_2628,N_1429,N_1235);
nor U2629 (N_2629,N_1297,N_1329);
nor U2630 (N_2630,N_1648,N_1191);
nand U2631 (N_2631,N_1517,N_1939);
nand U2632 (N_2632,N_1574,N_1952);
and U2633 (N_2633,N_1521,N_1929);
xor U2634 (N_2634,N_1670,N_1319);
nor U2635 (N_2635,N_1637,N_1974);
and U2636 (N_2636,N_1641,N_1617);
nor U2637 (N_2637,N_1306,N_1655);
nor U2638 (N_2638,N_1223,N_1567);
nand U2639 (N_2639,N_1287,N_1392);
xor U2640 (N_2640,N_1167,N_1160);
nand U2641 (N_2641,N_1740,N_1127);
or U2642 (N_2642,N_1215,N_1902);
or U2643 (N_2643,N_1700,N_1088);
and U2644 (N_2644,N_1278,N_1764);
nor U2645 (N_2645,N_1625,N_1838);
or U2646 (N_2646,N_1749,N_1410);
nand U2647 (N_2647,N_1277,N_1556);
nor U2648 (N_2648,N_1242,N_1196);
or U2649 (N_2649,N_1941,N_1863);
nor U2650 (N_2650,N_1318,N_1533);
or U2651 (N_2651,N_1590,N_1884);
nand U2652 (N_2652,N_1039,N_1537);
nand U2653 (N_2653,N_1860,N_1283);
or U2654 (N_2654,N_1674,N_1325);
nand U2655 (N_2655,N_1931,N_1752);
or U2656 (N_2656,N_1969,N_1396);
and U2657 (N_2657,N_1221,N_1436);
xor U2658 (N_2658,N_1630,N_1465);
nor U2659 (N_2659,N_1359,N_1355);
and U2660 (N_2660,N_1949,N_1097);
nand U2661 (N_2661,N_1648,N_1381);
nand U2662 (N_2662,N_1150,N_1739);
nand U2663 (N_2663,N_1420,N_1515);
nand U2664 (N_2664,N_1273,N_1638);
nor U2665 (N_2665,N_1828,N_1451);
nand U2666 (N_2666,N_1634,N_1662);
and U2667 (N_2667,N_1642,N_1566);
nand U2668 (N_2668,N_1470,N_1955);
xnor U2669 (N_2669,N_1627,N_1497);
nand U2670 (N_2670,N_1615,N_1722);
xnor U2671 (N_2671,N_1002,N_1726);
or U2672 (N_2672,N_1685,N_1422);
nand U2673 (N_2673,N_1032,N_1842);
and U2674 (N_2674,N_1933,N_1850);
or U2675 (N_2675,N_1624,N_1681);
nor U2676 (N_2676,N_1699,N_1182);
and U2677 (N_2677,N_1188,N_1336);
or U2678 (N_2678,N_1236,N_1576);
nor U2679 (N_2679,N_1074,N_1188);
and U2680 (N_2680,N_1298,N_1708);
or U2681 (N_2681,N_1090,N_1554);
nand U2682 (N_2682,N_1709,N_1089);
and U2683 (N_2683,N_1545,N_1845);
xnor U2684 (N_2684,N_1853,N_1060);
nor U2685 (N_2685,N_1363,N_1421);
or U2686 (N_2686,N_1771,N_1913);
and U2687 (N_2687,N_1661,N_1305);
nor U2688 (N_2688,N_1819,N_1975);
and U2689 (N_2689,N_1336,N_1052);
nor U2690 (N_2690,N_1587,N_1252);
nand U2691 (N_2691,N_1447,N_1357);
or U2692 (N_2692,N_1347,N_1387);
nor U2693 (N_2693,N_1247,N_1148);
or U2694 (N_2694,N_1116,N_1979);
nand U2695 (N_2695,N_1952,N_1796);
or U2696 (N_2696,N_1107,N_1497);
nor U2697 (N_2697,N_1823,N_1779);
nand U2698 (N_2698,N_1605,N_1027);
or U2699 (N_2699,N_1834,N_1021);
nand U2700 (N_2700,N_1796,N_1543);
and U2701 (N_2701,N_1087,N_1468);
and U2702 (N_2702,N_1466,N_1402);
or U2703 (N_2703,N_1619,N_1008);
and U2704 (N_2704,N_1107,N_1529);
or U2705 (N_2705,N_1742,N_1200);
or U2706 (N_2706,N_1976,N_1460);
nor U2707 (N_2707,N_1477,N_1062);
and U2708 (N_2708,N_1387,N_1667);
and U2709 (N_2709,N_1950,N_1726);
nand U2710 (N_2710,N_1213,N_1638);
or U2711 (N_2711,N_1753,N_1342);
or U2712 (N_2712,N_1820,N_1769);
or U2713 (N_2713,N_1797,N_1864);
nand U2714 (N_2714,N_1003,N_1435);
xnor U2715 (N_2715,N_1245,N_1548);
nor U2716 (N_2716,N_1104,N_1118);
or U2717 (N_2717,N_1238,N_1312);
nand U2718 (N_2718,N_1194,N_1262);
or U2719 (N_2719,N_1069,N_1007);
or U2720 (N_2720,N_1849,N_1818);
nor U2721 (N_2721,N_1785,N_1086);
and U2722 (N_2722,N_1532,N_1132);
and U2723 (N_2723,N_1436,N_1263);
and U2724 (N_2724,N_1975,N_1360);
or U2725 (N_2725,N_1920,N_1892);
nand U2726 (N_2726,N_1671,N_1579);
nor U2727 (N_2727,N_1416,N_1807);
nand U2728 (N_2728,N_1766,N_1659);
nor U2729 (N_2729,N_1665,N_1664);
nor U2730 (N_2730,N_1509,N_1127);
nor U2731 (N_2731,N_1314,N_1245);
and U2732 (N_2732,N_1683,N_1789);
nor U2733 (N_2733,N_1062,N_1528);
or U2734 (N_2734,N_1422,N_1765);
nand U2735 (N_2735,N_1876,N_1018);
nor U2736 (N_2736,N_1400,N_1757);
nor U2737 (N_2737,N_1473,N_1895);
and U2738 (N_2738,N_1284,N_1639);
nand U2739 (N_2739,N_1187,N_1595);
nor U2740 (N_2740,N_1919,N_1935);
and U2741 (N_2741,N_1021,N_1606);
nor U2742 (N_2742,N_1588,N_1996);
nand U2743 (N_2743,N_1875,N_1142);
nand U2744 (N_2744,N_1676,N_1415);
and U2745 (N_2745,N_1662,N_1085);
and U2746 (N_2746,N_1988,N_1150);
nor U2747 (N_2747,N_1481,N_1435);
and U2748 (N_2748,N_1693,N_1807);
nor U2749 (N_2749,N_1497,N_1093);
and U2750 (N_2750,N_1818,N_1519);
and U2751 (N_2751,N_1060,N_1652);
nor U2752 (N_2752,N_1429,N_1117);
or U2753 (N_2753,N_1276,N_1900);
and U2754 (N_2754,N_1709,N_1044);
nor U2755 (N_2755,N_1637,N_1716);
or U2756 (N_2756,N_1099,N_1283);
nand U2757 (N_2757,N_1530,N_1688);
nor U2758 (N_2758,N_1246,N_1152);
xnor U2759 (N_2759,N_1883,N_1529);
nor U2760 (N_2760,N_1002,N_1649);
and U2761 (N_2761,N_1281,N_1091);
or U2762 (N_2762,N_1845,N_1771);
nor U2763 (N_2763,N_1413,N_1773);
nand U2764 (N_2764,N_1287,N_1446);
or U2765 (N_2765,N_1006,N_1339);
nand U2766 (N_2766,N_1028,N_1231);
nor U2767 (N_2767,N_1748,N_1892);
nor U2768 (N_2768,N_1604,N_1899);
nand U2769 (N_2769,N_1919,N_1188);
and U2770 (N_2770,N_1306,N_1376);
nor U2771 (N_2771,N_1723,N_1384);
or U2772 (N_2772,N_1033,N_1192);
xnor U2773 (N_2773,N_1051,N_1944);
nand U2774 (N_2774,N_1209,N_1808);
or U2775 (N_2775,N_1277,N_1671);
nand U2776 (N_2776,N_1376,N_1649);
nand U2777 (N_2777,N_1169,N_1739);
xnor U2778 (N_2778,N_1562,N_1710);
and U2779 (N_2779,N_1061,N_1512);
nor U2780 (N_2780,N_1641,N_1640);
nor U2781 (N_2781,N_1171,N_1577);
nand U2782 (N_2782,N_1787,N_1820);
nand U2783 (N_2783,N_1802,N_1630);
and U2784 (N_2784,N_1637,N_1583);
nand U2785 (N_2785,N_1884,N_1601);
nor U2786 (N_2786,N_1403,N_1195);
nor U2787 (N_2787,N_1361,N_1935);
nor U2788 (N_2788,N_1837,N_1047);
and U2789 (N_2789,N_1599,N_1053);
xor U2790 (N_2790,N_1053,N_1258);
nand U2791 (N_2791,N_1820,N_1784);
nor U2792 (N_2792,N_1778,N_1881);
and U2793 (N_2793,N_1356,N_1659);
nor U2794 (N_2794,N_1433,N_1078);
nand U2795 (N_2795,N_1520,N_1833);
and U2796 (N_2796,N_1130,N_1886);
nand U2797 (N_2797,N_1424,N_1074);
nand U2798 (N_2798,N_1315,N_1618);
xnor U2799 (N_2799,N_1757,N_1257);
or U2800 (N_2800,N_1791,N_1386);
and U2801 (N_2801,N_1027,N_1515);
nand U2802 (N_2802,N_1745,N_1257);
nor U2803 (N_2803,N_1756,N_1247);
nand U2804 (N_2804,N_1316,N_1607);
nand U2805 (N_2805,N_1392,N_1405);
nor U2806 (N_2806,N_1026,N_1544);
and U2807 (N_2807,N_1853,N_1113);
nor U2808 (N_2808,N_1586,N_1036);
nand U2809 (N_2809,N_1310,N_1187);
nand U2810 (N_2810,N_1501,N_1440);
and U2811 (N_2811,N_1157,N_1855);
nor U2812 (N_2812,N_1925,N_1618);
and U2813 (N_2813,N_1946,N_1060);
nor U2814 (N_2814,N_1577,N_1679);
or U2815 (N_2815,N_1177,N_1503);
nand U2816 (N_2816,N_1147,N_1457);
nor U2817 (N_2817,N_1353,N_1084);
or U2818 (N_2818,N_1628,N_1316);
or U2819 (N_2819,N_1308,N_1039);
and U2820 (N_2820,N_1610,N_1325);
xor U2821 (N_2821,N_1419,N_1604);
or U2822 (N_2822,N_1287,N_1355);
and U2823 (N_2823,N_1741,N_1234);
nand U2824 (N_2824,N_1971,N_1433);
nor U2825 (N_2825,N_1539,N_1052);
and U2826 (N_2826,N_1729,N_1211);
nand U2827 (N_2827,N_1006,N_1273);
and U2828 (N_2828,N_1211,N_1580);
and U2829 (N_2829,N_1465,N_1089);
or U2830 (N_2830,N_1482,N_1678);
and U2831 (N_2831,N_1784,N_1824);
or U2832 (N_2832,N_1869,N_1824);
and U2833 (N_2833,N_1799,N_1379);
and U2834 (N_2834,N_1048,N_1839);
and U2835 (N_2835,N_1609,N_1767);
nand U2836 (N_2836,N_1755,N_1068);
nand U2837 (N_2837,N_1669,N_1860);
nand U2838 (N_2838,N_1283,N_1345);
and U2839 (N_2839,N_1708,N_1485);
nand U2840 (N_2840,N_1650,N_1306);
and U2841 (N_2841,N_1401,N_1183);
nand U2842 (N_2842,N_1195,N_1612);
nor U2843 (N_2843,N_1946,N_1570);
nand U2844 (N_2844,N_1136,N_1019);
nor U2845 (N_2845,N_1533,N_1884);
nor U2846 (N_2846,N_1731,N_1993);
nor U2847 (N_2847,N_1233,N_1694);
or U2848 (N_2848,N_1301,N_1895);
nand U2849 (N_2849,N_1963,N_1642);
or U2850 (N_2850,N_1996,N_1404);
nor U2851 (N_2851,N_1522,N_1879);
nor U2852 (N_2852,N_1826,N_1347);
nand U2853 (N_2853,N_1070,N_1827);
nand U2854 (N_2854,N_1839,N_1405);
and U2855 (N_2855,N_1649,N_1996);
or U2856 (N_2856,N_1044,N_1690);
and U2857 (N_2857,N_1103,N_1132);
or U2858 (N_2858,N_1147,N_1195);
and U2859 (N_2859,N_1356,N_1982);
and U2860 (N_2860,N_1480,N_1055);
nand U2861 (N_2861,N_1376,N_1140);
or U2862 (N_2862,N_1983,N_1255);
nand U2863 (N_2863,N_1973,N_1260);
nor U2864 (N_2864,N_1970,N_1898);
and U2865 (N_2865,N_1166,N_1461);
and U2866 (N_2866,N_1194,N_1816);
or U2867 (N_2867,N_1678,N_1531);
nor U2868 (N_2868,N_1289,N_1393);
or U2869 (N_2869,N_1655,N_1417);
and U2870 (N_2870,N_1443,N_1365);
nand U2871 (N_2871,N_1083,N_1361);
xor U2872 (N_2872,N_1329,N_1211);
nand U2873 (N_2873,N_1558,N_1632);
and U2874 (N_2874,N_1821,N_1561);
or U2875 (N_2875,N_1012,N_1450);
or U2876 (N_2876,N_1912,N_1820);
or U2877 (N_2877,N_1956,N_1598);
nand U2878 (N_2878,N_1294,N_1483);
or U2879 (N_2879,N_1567,N_1913);
and U2880 (N_2880,N_1731,N_1991);
nor U2881 (N_2881,N_1836,N_1487);
or U2882 (N_2882,N_1908,N_1978);
or U2883 (N_2883,N_1883,N_1182);
and U2884 (N_2884,N_1656,N_1196);
nor U2885 (N_2885,N_1020,N_1247);
nand U2886 (N_2886,N_1766,N_1954);
nor U2887 (N_2887,N_1416,N_1003);
nand U2888 (N_2888,N_1353,N_1639);
nand U2889 (N_2889,N_1336,N_1701);
nand U2890 (N_2890,N_1907,N_1718);
and U2891 (N_2891,N_1253,N_1104);
nor U2892 (N_2892,N_1408,N_1584);
and U2893 (N_2893,N_1189,N_1125);
nor U2894 (N_2894,N_1103,N_1158);
and U2895 (N_2895,N_1525,N_1153);
or U2896 (N_2896,N_1317,N_1398);
or U2897 (N_2897,N_1646,N_1570);
nand U2898 (N_2898,N_1571,N_1722);
or U2899 (N_2899,N_1209,N_1940);
nor U2900 (N_2900,N_1806,N_1357);
nor U2901 (N_2901,N_1196,N_1395);
nor U2902 (N_2902,N_1109,N_1775);
nor U2903 (N_2903,N_1013,N_1402);
or U2904 (N_2904,N_1550,N_1635);
nor U2905 (N_2905,N_1403,N_1282);
or U2906 (N_2906,N_1827,N_1039);
nand U2907 (N_2907,N_1822,N_1111);
nand U2908 (N_2908,N_1094,N_1871);
and U2909 (N_2909,N_1066,N_1244);
or U2910 (N_2910,N_1392,N_1598);
and U2911 (N_2911,N_1203,N_1872);
nor U2912 (N_2912,N_1693,N_1066);
nand U2913 (N_2913,N_1911,N_1933);
xor U2914 (N_2914,N_1184,N_1076);
or U2915 (N_2915,N_1019,N_1068);
nor U2916 (N_2916,N_1063,N_1966);
or U2917 (N_2917,N_1311,N_1791);
nor U2918 (N_2918,N_1788,N_1746);
nand U2919 (N_2919,N_1596,N_1445);
and U2920 (N_2920,N_1069,N_1496);
or U2921 (N_2921,N_1350,N_1759);
nor U2922 (N_2922,N_1048,N_1364);
and U2923 (N_2923,N_1852,N_1141);
nand U2924 (N_2924,N_1174,N_1381);
or U2925 (N_2925,N_1535,N_1315);
nor U2926 (N_2926,N_1893,N_1501);
nor U2927 (N_2927,N_1860,N_1275);
and U2928 (N_2928,N_1148,N_1194);
or U2929 (N_2929,N_1119,N_1753);
xnor U2930 (N_2930,N_1665,N_1571);
and U2931 (N_2931,N_1868,N_1112);
nor U2932 (N_2932,N_1474,N_1795);
nand U2933 (N_2933,N_1199,N_1857);
nand U2934 (N_2934,N_1356,N_1588);
nand U2935 (N_2935,N_1466,N_1417);
nand U2936 (N_2936,N_1219,N_1306);
nor U2937 (N_2937,N_1779,N_1108);
and U2938 (N_2938,N_1231,N_1339);
and U2939 (N_2939,N_1062,N_1250);
and U2940 (N_2940,N_1087,N_1352);
nor U2941 (N_2941,N_1024,N_1124);
and U2942 (N_2942,N_1167,N_1212);
xor U2943 (N_2943,N_1550,N_1625);
nor U2944 (N_2944,N_1061,N_1342);
or U2945 (N_2945,N_1377,N_1554);
nand U2946 (N_2946,N_1184,N_1789);
nand U2947 (N_2947,N_1334,N_1527);
or U2948 (N_2948,N_1779,N_1094);
and U2949 (N_2949,N_1024,N_1603);
and U2950 (N_2950,N_1536,N_1468);
nand U2951 (N_2951,N_1981,N_1274);
or U2952 (N_2952,N_1535,N_1494);
nor U2953 (N_2953,N_1981,N_1478);
and U2954 (N_2954,N_1526,N_1415);
and U2955 (N_2955,N_1665,N_1342);
nand U2956 (N_2956,N_1971,N_1841);
nand U2957 (N_2957,N_1243,N_1074);
or U2958 (N_2958,N_1711,N_1503);
or U2959 (N_2959,N_1522,N_1837);
nand U2960 (N_2960,N_1442,N_1471);
nor U2961 (N_2961,N_1879,N_1493);
and U2962 (N_2962,N_1577,N_1712);
nand U2963 (N_2963,N_1507,N_1996);
nand U2964 (N_2964,N_1224,N_1585);
nand U2965 (N_2965,N_1020,N_1455);
nand U2966 (N_2966,N_1005,N_1836);
xnor U2967 (N_2967,N_1001,N_1760);
and U2968 (N_2968,N_1826,N_1317);
xor U2969 (N_2969,N_1384,N_1912);
and U2970 (N_2970,N_1408,N_1363);
nand U2971 (N_2971,N_1834,N_1980);
or U2972 (N_2972,N_1785,N_1788);
nand U2973 (N_2973,N_1664,N_1997);
and U2974 (N_2974,N_1891,N_1049);
or U2975 (N_2975,N_1721,N_1954);
nand U2976 (N_2976,N_1991,N_1550);
nor U2977 (N_2977,N_1989,N_1357);
nor U2978 (N_2978,N_1866,N_1640);
or U2979 (N_2979,N_1065,N_1921);
nor U2980 (N_2980,N_1384,N_1876);
and U2981 (N_2981,N_1767,N_1909);
and U2982 (N_2982,N_1691,N_1771);
nor U2983 (N_2983,N_1869,N_1283);
nor U2984 (N_2984,N_1801,N_1581);
nor U2985 (N_2985,N_1289,N_1921);
nor U2986 (N_2986,N_1108,N_1480);
and U2987 (N_2987,N_1491,N_1893);
and U2988 (N_2988,N_1187,N_1094);
or U2989 (N_2989,N_1617,N_1863);
and U2990 (N_2990,N_1260,N_1234);
or U2991 (N_2991,N_1861,N_1028);
and U2992 (N_2992,N_1312,N_1013);
or U2993 (N_2993,N_1358,N_1002);
nand U2994 (N_2994,N_1984,N_1352);
nand U2995 (N_2995,N_1740,N_1849);
and U2996 (N_2996,N_1496,N_1839);
nor U2997 (N_2997,N_1361,N_1579);
nor U2998 (N_2998,N_1085,N_1540);
or U2999 (N_2999,N_1623,N_1781);
nand UO_0 (O_0,N_2892,N_2286);
or UO_1 (O_1,N_2386,N_2314);
or UO_2 (O_2,N_2470,N_2742);
xor UO_3 (O_3,N_2917,N_2418);
nor UO_4 (O_4,N_2708,N_2489);
nand UO_5 (O_5,N_2010,N_2397);
nand UO_6 (O_6,N_2549,N_2529);
or UO_7 (O_7,N_2429,N_2838);
nand UO_8 (O_8,N_2372,N_2378);
or UO_9 (O_9,N_2180,N_2499);
and UO_10 (O_10,N_2756,N_2471);
nor UO_11 (O_11,N_2234,N_2951);
xnor UO_12 (O_12,N_2550,N_2704);
nor UO_13 (O_13,N_2814,N_2115);
nor UO_14 (O_14,N_2661,N_2349);
and UO_15 (O_15,N_2285,N_2227);
nor UO_16 (O_16,N_2518,N_2999);
and UO_17 (O_17,N_2943,N_2767);
or UO_18 (O_18,N_2051,N_2419);
nand UO_19 (O_19,N_2212,N_2982);
and UO_20 (O_20,N_2732,N_2241);
nand UO_21 (O_21,N_2639,N_2565);
nand UO_22 (O_22,N_2364,N_2843);
and UO_23 (O_23,N_2120,N_2213);
and UO_24 (O_24,N_2260,N_2291);
nand UO_25 (O_25,N_2510,N_2434);
and UO_26 (O_26,N_2146,N_2214);
nand UO_27 (O_27,N_2487,N_2857);
and UO_28 (O_28,N_2970,N_2840);
or UO_29 (O_29,N_2312,N_2348);
nand UO_30 (O_30,N_2083,N_2233);
or UO_31 (O_31,N_2566,N_2997);
and UO_32 (O_32,N_2346,N_2316);
nor UO_33 (O_33,N_2101,N_2779);
or UO_34 (O_34,N_2624,N_2579);
or UO_35 (O_35,N_2647,N_2939);
or UO_36 (O_36,N_2209,N_2502);
xnor UO_37 (O_37,N_2531,N_2297);
or UO_38 (O_38,N_2721,N_2652);
and UO_39 (O_39,N_2395,N_2517);
nor UO_40 (O_40,N_2469,N_2932);
or UO_41 (O_41,N_2221,N_2280);
and UO_42 (O_42,N_2793,N_2724);
and UO_43 (O_43,N_2203,N_2522);
or UO_44 (O_44,N_2025,N_2167);
nor UO_45 (O_45,N_2799,N_2050);
nand UO_46 (O_46,N_2005,N_2290);
nor UO_47 (O_47,N_2833,N_2466);
nand UO_48 (O_48,N_2757,N_2431);
nand UO_49 (O_49,N_2614,N_2974);
nand UO_50 (O_50,N_2995,N_2192);
and UO_51 (O_51,N_2141,N_2210);
xor UO_52 (O_52,N_2584,N_2946);
nor UO_53 (O_53,N_2926,N_2207);
and UO_54 (O_54,N_2353,N_2106);
and UO_55 (O_55,N_2244,N_2633);
and UO_56 (O_56,N_2889,N_2424);
or UO_57 (O_57,N_2636,N_2295);
and UO_58 (O_58,N_2491,N_2743);
or UO_59 (O_59,N_2069,N_2712);
and UO_60 (O_60,N_2407,N_2964);
nor UO_61 (O_61,N_2042,N_2271);
nor UO_62 (O_62,N_2139,N_2880);
or UO_63 (O_63,N_2899,N_2024);
or UO_64 (O_64,N_2329,N_2702);
nor UO_65 (O_65,N_2648,N_2119);
nand UO_66 (O_66,N_2805,N_2507);
and UO_67 (O_67,N_2334,N_2483);
or UO_68 (O_68,N_2947,N_2125);
nor UO_69 (O_69,N_2953,N_2354);
or UO_70 (O_70,N_2226,N_2055);
nor UO_71 (O_71,N_2933,N_2835);
nand UO_72 (O_72,N_2856,N_2384);
or UO_73 (O_73,N_2338,N_2012);
nor UO_74 (O_74,N_2655,N_2706);
nand UO_75 (O_75,N_2711,N_2422);
and UO_76 (O_76,N_2797,N_2401);
nor UO_77 (O_77,N_2519,N_2570);
xor UO_78 (O_78,N_2744,N_2156);
and UO_79 (O_79,N_2362,N_2243);
or UO_80 (O_80,N_2476,N_2077);
xor UO_81 (O_81,N_2006,N_2720);
nand UO_82 (O_82,N_2028,N_2102);
xor UO_83 (O_83,N_2788,N_2130);
xor UO_84 (O_84,N_2361,N_2199);
or UO_85 (O_85,N_2008,N_2668);
and UO_86 (O_86,N_2056,N_2701);
nand UO_87 (O_87,N_2147,N_2670);
nand UO_88 (O_88,N_2194,N_2099);
and UO_89 (O_89,N_2467,N_2906);
nor UO_90 (O_90,N_2071,N_2546);
nand UO_91 (O_91,N_2231,N_2446);
nor UO_92 (O_92,N_2820,N_2236);
nand UO_93 (O_93,N_2237,N_2317);
nand UO_94 (O_94,N_2060,N_2621);
xnor UO_95 (O_95,N_2311,N_2627);
or UO_96 (O_96,N_2664,N_2722);
or UO_97 (O_97,N_2760,N_2726);
or UO_98 (O_98,N_2681,N_2885);
nor UO_99 (O_99,N_2331,N_2924);
or UO_100 (O_100,N_2457,N_2490);
nor UO_101 (O_101,N_2861,N_2961);
and UO_102 (O_102,N_2406,N_2716);
nor UO_103 (O_103,N_2941,N_2078);
and UO_104 (O_104,N_2993,N_2642);
nor UO_105 (O_105,N_2343,N_2171);
nor UO_106 (O_106,N_2543,N_2504);
or UO_107 (O_107,N_2436,N_2088);
or UO_108 (O_108,N_2665,N_2275);
or UO_109 (O_109,N_2162,N_2200);
and UO_110 (O_110,N_2062,N_2766);
or UO_111 (O_111,N_2644,N_2693);
or UO_112 (O_112,N_2085,N_2765);
and UO_113 (O_113,N_2332,N_2414);
nand UO_114 (O_114,N_2195,N_2298);
xor UO_115 (O_115,N_2325,N_2018);
nor UO_116 (O_116,N_2268,N_2428);
xor UO_117 (O_117,N_2824,N_2834);
or UO_118 (O_118,N_2854,N_2986);
and UO_119 (O_119,N_2206,N_2293);
nor UO_120 (O_120,N_2448,N_2445);
and UO_121 (O_121,N_2780,N_2002);
nand UO_122 (O_122,N_2656,N_2092);
nor UO_123 (O_123,N_2294,N_2255);
nand UO_124 (O_124,N_2315,N_2505);
or UO_125 (O_125,N_2122,N_2322);
and UO_126 (O_126,N_2340,N_2968);
or UO_127 (O_127,N_2152,N_2117);
or UO_128 (O_128,N_2605,N_2021);
nand UO_129 (O_129,N_2931,N_2818);
nand UO_130 (O_130,N_2287,N_2450);
nor UO_131 (O_131,N_2278,N_2615);
nand UO_132 (O_132,N_2806,N_2279);
or UO_133 (O_133,N_2082,N_2155);
or UO_134 (O_134,N_2893,N_2442);
or UO_135 (O_135,N_2523,N_2262);
and UO_136 (O_136,N_2734,N_2815);
or UO_137 (O_137,N_2738,N_2411);
nor UO_138 (O_138,N_2859,N_2729);
or UO_139 (O_139,N_2913,N_2850);
or UO_140 (O_140,N_2011,N_2076);
or UO_141 (O_141,N_2950,N_2145);
nor UO_142 (O_142,N_2819,N_2219);
nand UO_143 (O_143,N_2020,N_2918);
and UO_144 (O_144,N_2687,N_2527);
and UO_145 (O_145,N_2230,N_2075);
nor UO_146 (O_146,N_2983,N_2925);
or UO_147 (O_147,N_2172,N_2555);
and UO_148 (O_148,N_2274,N_2870);
xor UO_149 (O_149,N_2852,N_2124);
and UO_150 (O_150,N_2173,N_2320);
and UO_151 (O_151,N_2336,N_2328);
nor UO_152 (O_152,N_2530,N_2136);
and UO_153 (O_153,N_2956,N_2126);
or UO_154 (O_154,N_2034,N_2848);
nor UO_155 (O_155,N_2508,N_2103);
or UO_156 (O_156,N_2225,N_2762);
xnor UO_157 (O_157,N_2758,N_2506);
or UO_158 (O_158,N_2169,N_2830);
or UO_159 (O_159,N_2067,N_2697);
nand UO_160 (O_160,N_2586,N_2773);
or UO_161 (O_161,N_2973,N_2065);
xnor UO_162 (O_162,N_2938,N_2360);
or UO_163 (O_163,N_2356,N_2532);
or UO_164 (O_164,N_2149,N_2984);
and UO_165 (O_165,N_2168,N_2193);
nand UO_166 (O_166,N_2501,N_2842);
nand UO_167 (O_167,N_2849,N_2321);
and UO_168 (O_168,N_2001,N_2402);
or UO_169 (O_169,N_2879,N_2868);
nand UO_170 (O_170,N_2571,N_2975);
and UO_171 (O_171,N_2560,N_2373);
nand UO_172 (O_172,N_2229,N_2417);
nand UO_173 (O_173,N_2447,N_2073);
and UO_174 (O_174,N_2715,N_2351);
nand UO_175 (O_175,N_2474,N_2405);
or UO_176 (O_176,N_2178,N_2239);
nor UO_177 (O_177,N_2710,N_2277);
and UO_178 (O_178,N_2463,N_2232);
and UO_179 (O_179,N_2427,N_2383);
or UO_180 (O_180,N_2461,N_2750);
nor UO_181 (O_181,N_2804,N_2246);
or UO_182 (O_182,N_2841,N_2914);
and UO_183 (O_183,N_2577,N_2632);
nand UO_184 (O_184,N_2503,N_2423);
nand UO_185 (O_185,N_2545,N_2536);
nor UO_186 (O_186,N_2540,N_2563);
and UO_187 (O_187,N_2904,N_2900);
or UO_188 (O_188,N_2719,N_2257);
nand UO_189 (O_189,N_2657,N_2377);
nor UO_190 (O_190,N_2735,N_2421);
and UO_191 (O_191,N_2304,N_2717);
or UO_192 (O_192,N_2683,N_2324);
and UO_193 (O_193,N_2572,N_2033);
or UO_194 (O_194,N_2537,N_2674);
or UO_195 (O_195,N_2971,N_2333);
nand UO_196 (O_196,N_2610,N_2086);
and UO_197 (O_197,N_2641,N_2435);
and UO_198 (O_198,N_2218,N_2177);
nor UO_199 (O_199,N_2408,N_2544);
or UO_200 (O_200,N_2190,N_2070);
nor UO_201 (O_201,N_2794,N_2616);
nor UO_202 (O_202,N_2630,N_2538);
and UO_203 (O_203,N_2238,N_2250);
and UO_204 (O_204,N_2955,N_2249);
nand UO_205 (O_205,N_2612,N_2969);
xor UO_206 (O_206,N_2705,N_2682);
and UO_207 (O_207,N_2035,N_2366);
and UO_208 (O_208,N_2525,N_2604);
or UO_209 (O_209,N_2201,N_2494);
or UO_210 (O_210,N_2910,N_2671);
or UO_211 (O_211,N_2748,N_2675);
and UO_212 (O_212,N_2980,N_2381);
nand UO_213 (O_213,N_2808,N_2666);
nor UO_214 (O_214,N_2266,N_2844);
nor UO_215 (O_215,N_2443,N_2022);
nor UO_216 (O_216,N_2363,N_2821);
nand UO_217 (O_217,N_2184,N_2942);
or UO_218 (O_218,N_2047,N_2521);
and UO_219 (O_219,N_2862,N_2472);
xnor UO_220 (O_220,N_2759,N_2622);
nand UO_221 (O_221,N_2134,N_2619);
nor UO_222 (O_222,N_2958,N_2617);
nand UO_223 (O_223,N_2396,N_2347);
or UO_224 (O_224,N_2387,N_2258);
nand UO_225 (O_225,N_2763,N_2030);
and UO_226 (O_226,N_2598,N_2599);
or UO_227 (O_227,N_2089,N_2380);
nor UO_228 (O_228,N_2137,N_2669);
or UO_229 (O_229,N_2928,N_2009);
nor UO_230 (O_230,N_2723,N_2822);
nor UO_231 (O_231,N_2595,N_2660);
nor UO_232 (O_232,N_2620,N_2151);
and UO_233 (O_233,N_2326,N_2772);
nor UO_234 (O_234,N_2945,N_2987);
nand UO_235 (O_235,N_2475,N_2394);
or UO_236 (O_236,N_2131,N_2851);
or UO_237 (O_237,N_2123,N_2662);
nor UO_238 (O_238,N_2198,N_2288);
nand UO_239 (O_239,N_2399,N_2063);
nand UO_240 (O_240,N_2509,N_2369);
nor UO_241 (O_241,N_2046,N_2118);
or UO_242 (O_242,N_2486,N_2409);
nor UO_243 (O_243,N_2651,N_2526);
nand UO_244 (O_244,N_2299,N_2189);
or UO_245 (O_245,N_2292,N_2004);
nand UO_246 (O_246,N_2860,N_2846);
nor UO_247 (O_247,N_2667,N_2553);
nand UO_248 (O_248,N_2342,N_2112);
nand UO_249 (O_249,N_2330,N_2144);
nor UO_250 (O_250,N_2684,N_2784);
nand UO_251 (O_251,N_2769,N_2157);
or UO_252 (O_252,N_2359,N_2204);
nor UO_253 (O_253,N_2916,N_2438);
nor UO_254 (O_254,N_2937,N_2400);
or UO_255 (O_255,N_2954,N_2680);
nand UO_256 (O_256,N_2658,N_2367);
nor UO_257 (O_257,N_2812,N_2220);
nand UO_258 (O_258,N_2875,N_2319);
or UO_259 (O_259,N_2026,N_2371);
or UO_260 (O_260,N_2912,N_2019);
and UO_261 (O_261,N_2302,N_2686);
or UO_262 (O_262,N_2464,N_2989);
or UO_263 (O_263,N_2003,N_2927);
or UO_264 (O_264,N_2618,N_2589);
nand UO_265 (O_265,N_2420,N_2044);
and UO_266 (O_266,N_2978,N_2810);
nor UO_267 (O_267,N_2813,N_2921);
nor UO_268 (O_268,N_2087,N_2495);
nor UO_269 (O_269,N_2606,N_2135);
and UO_270 (O_270,N_2388,N_2079);
and UO_271 (O_271,N_2375,N_2569);
nand UO_272 (O_272,N_2654,N_2393);
and UO_273 (O_273,N_2281,N_2211);
nand UO_274 (O_274,N_2497,N_2276);
or UO_275 (O_275,N_2175,N_2498);
and UO_276 (O_276,N_2263,N_2318);
nand UO_277 (O_277,N_2747,N_2777);
and UO_278 (O_278,N_2093,N_2480);
nor UO_279 (O_279,N_2223,N_2795);
and UO_280 (O_280,N_2803,N_2802);
or UO_281 (O_281,N_2901,N_2128);
and UO_282 (O_282,N_2873,N_2040);
and UO_283 (O_283,N_2897,N_2382);
or UO_284 (O_284,N_2404,N_2170);
nor UO_285 (O_285,N_2164,N_2344);
nor UO_286 (O_286,N_2864,N_2809);
and UO_287 (O_287,N_2037,N_2981);
nand UO_288 (O_288,N_2597,N_2609);
or UO_289 (O_289,N_2308,N_2301);
nor UO_290 (O_290,N_2825,N_2534);
and UO_291 (O_291,N_2695,N_2979);
or UO_292 (O_292,N_2269,N_2339);
nand UO_293 (O_293,N_2465,N_2049);
or UO_294 (O_294,N_2608,N_2098);
nor UO_295 (O_295,N_2064,N_2798);
xnor UO_296 (O_296,N_2165,N_2458);
and UO_297 (O_297,N_2478,N_2138);
or UO_298 (O_298,N_2965,N_2692);
and UO_299 (O_299,N_2068,N_2645);
and UO_300 (O_300,N_2273,N_2740);
and UO_301 (O_301,N_2129,N_2222);
nand UO_302 (O_302,N_2023,N_2245);
nand UO_303 (O_303,N_2548,N_2254);
nand UO_304 (O_304,N_2041,N_2628);
nor UO_305 (O_305,N_2453,N_2886);
or UO_306 (O_306,N_2554,N_2535);
nor UO_307 (O_307,N_2452,N_2057);
nor UO_308 (O_308,N_2588,N_2678);
or UO_309 (O_309,N_2385,N_2929);
xnor UO_310 (O_310,N_2725,N_2930);
nand UO_311 (O_311,N_2751,N_2307);
or UO_312 (O_312,N_2090,N_2878);
and UO_313 (O_313,N_2456,N_2186);
nor UO_314 (O_314,N_2728,N_2576);
and UO_315 (O_315,N_2966,N_2533);
nand UO_316 (O_316,N_2310,N_2948);
nor UO_317 (O_317,N_2876,N_2043);
nor UO_318 (O_318,N_2736,N_2185);
xnor UO_319 (O_319,N_2631,N_2365);
and UO_320 (O_320,N_2782,N_2659);
nand UO_321 (O_321,N_2855,N_2768);
nand UO_322 (O_322,N_2158,N_2058);
or UO_323 (O_323,N_2727,N_2413);
or UO_324 (O_324,N_2224,N_2066);
or UO_325 (O_325,N_2771,N_2593);
nand UO_326 (O_326,N_2646,N_2634);
and UO_327 (O_327,N_2160,N_2649);
nor UO_328 (O_328,N_2603,N_2585);
nor UO_329 (O_329,N_2996,N_2991);
or UO_330 (O_330,N_2872,N_2962);
nor UO_331 (O_331,N_2449,N_2564);
or UO_332 (O_332,N_2094,N_2764);
nand UO_333 (O_333,N_2568,N_2350);
and UO_334 (O_334,N_2080,N_2709);
and UO_335 (O_335,N_2036,N_2183);
and UO_336 (O_336,N_2866,N_2282);
nor UO_337 (O_337,N_2352,N_2836);
and UO_338 (O_338,N_2539,N_2888);
nand UO_339 (O_339,N_2561,N_2296);
and UO_340 (O_340,N_2988,N_2327);
and UO_341 (O_341,N_2944,N_2713);
xor UO_342 (O_342,N_2573,N_2635);
nand UO_343 (O_343,N_2679,N_2629);
nand UO_344 (O_344,N_2858,N_2473);
nor UO_345 (O_345,N_2052,N_2783);
nand UO_346 (O_346,N_2110,N_2454);
and UO_347 (O_347,N_2074,N_2267);
nand UO_348 (O_348,N_2638,N_2029);
nand UO_349 (O_349,N_2919,N_2908);
or UO_350 (O_350,N_2807,N_2903);
or UO_351 (O_351,N_2755,N_2992);
nand UO_352 (O_352,N_2007,N_2140);
xnor UO_353 (O_353,N_2559,N_2459);
nor UO_354 (O_354,N_2578,N_2240);
nand UO_355 (O_355,N_2541,N_2460);
nor UO_356 (O_356,N_2337,N_2789);
or UO_357 (O_357,N_2587,N_2884);
and UO_358 (O_358,N_2863,N_2081);
and UO_359 (O_359,N_2949,N_2444);
nand UO_360 (O_360,N_2557,N_2358);
and UO_361 (O_361,N_2785,N_2468);
nand UO_362 (O_362,N_2289,N_2994);
or UO_363 (O_363,N_2865,N_2514);
or UO_364 (O_364,N_2215,N_2831);
and UO_365 (O_365,N_2432,N_2677);
or UO_366 (O_366,N_2934,N_2196);
or UO_367 (O_367,N_2091,N_2694);
nor UO_368 (O_368,N_2500,N_2672);
nor UO_369 (O_369,N_2881,N_2492);
nor UO_370 (O_370,N_2776,N_2389);
or UO_371 (O_371,N_2580,N_2556);
or UO_372 (O_372,N_2095,N_2650);
and UO_373 (O_373,N_2967,N_2187);
and UO_374 (O_374,N_2781,N_2216);
nor UO_375 (O_375,N_2817,N_2714);
nor UO_376 (O_376,N_2261,N_2832);
nand UO_377 (O_377,N_2707,N_2515);
xor UO_378 (O_378,N_2013,N_2922);
or UO_379 (O_379,N_2513,N_2462);
or UO_380 (O_380,N_2935,N_2733);
and UO_381 (O_381,N_2217,N_2259);
or UO_382 (O_382,N_2582,N_2481);
nor UO_383 (O_383,N_2054,N_2496);
nand UO_384 (O_384,N_2703,N_2053);
nand UO_385 (O_385,N_2829,N_2017);
nor UO_386 (O_386,N_2826,N_2749);
xor UO_387 (O_387,N_2264,N_2567);
nor UO_388 (O_388,N_2084,N_2786);
or UO_389 (O_389,N_2096,N_2623);
nor UO_390 (O_390,N_2403,N_2109);
nor UO_391 (O_391,N_2309,N_2441);
nand UO_392 (O_392,N_2440,N_2611);
nor UO_393 (O_393,N_2528,N_2247);
nand UO_394 (O_394,N_2891,N_2883);
or UO_395 (O_395,N_2032,N_2031);
or UO_396 (O_396,N_2594,N_2552);
or UO_397 (O_397,N_2699,N_2796);
and UO_398 (O_398,N_2600,N_2113);
and UO_399 (O_399,N_2197,N_2700);
and UO_400 (O_400,N_2121,N_2920);
nand UO_401 (O_401,N_2575,N_2752);
nor UO_402 (O_402,N_2208,N_2256);
and UO_403 (O_403,N_2272,N_2248);
nand UO_404 (O_404,N_2691,N_2205);
and UO_405 (O_405,N_2590,N_2626);
nor UO_406 (O_406,N_2663,N_2283);
or UO_407 (O_407,N_2963,N_2038);
nor UO_408 (O_408,N_2990,N_2898);
nor UO_409 (O_409,N_2105,N_2801);
or UO_410 (O_410,N_2410,N_2602);
or UO_411 (O_411,N_2398,N_2368);
nor UO_412 (O_412,N_2390,N_2839);
xor UO_413 (O_413,N_2142,N_2300);
and UO_414 (O_414,N_2412,N_2048);
nand UO_415 (O_415,N_2355,N_2845);
nand UO_416 (O_416,N_2150,N_2972);
or UO_417 (O_417,N_2188,N_2376);
nor UO_418 (O_418,N_2143,N_2542);
and UO_419 (O_419,N_2437,N_2909);
nor UO_420 (O_420,N_2688,N_2323);
nor UO_421 (O_421,N_2161,N_2770);
nand UO_422 (O_422,N_2753,N_2015);
or UO_423 (O_423,N_2426,N_2640);
nand UO_424 (O_424,N_2718,N_2960);
nand UO_425 (O_425,N_2828,N_2191);
nor UO_426 (O_426,N_2811,N_2379);
or UO_427 (O_427,N_2847,N_2108);
nor UO_428 (O_428,N_2696,N_2775);
and UO_429 (O_429,N_2111,N_2558);
nand UO_430 (O_430,N_2653,N_2520);
xnor UO_431 (O_431,N_2698,N_2731);
xnor UO_432 (O_432,N_2416,N_2159);
or UO_433 (O_433,N_2730,N_2455);
nand UO_434 (O_434,N_2512,N_2202);
or UO_435 (O_435,N_2251,N_2132);
and UO_436 (O_436,N_2874,N_2341);
nor UO_437 (O_437,N_2867,N_2761);
or UO_438 (O_438,N_2270,N_2061);
or UO_439 (O_439,N_2228,N_2689);
nor UO_440 (O_440,N_2305,N_2415);
and UO_441 (O_441,N_2592,N_2039);
nand UO_442 (O_442,N_2345,N_2905);
or UO_443 (O_443,N_2792,N_2133);
or UO_444 (O_444,N_2059,N_2685);
nand UO_445 (O_445,N_2581,N_2127);
nor UO_446 (O_446,N_2911,N_2936);
nand UO_447 (O_447,N_2871,N_2511);
nor UO_448 (O_448,N_2000,N_2837);
nand UO_449 (O_449,N_2739,N_2016);
and UO_450 (O_450,N_2902,N_2998);
nor UO_451 (O_451,N_2100,N_2451);
and UO_452 (O_452,N_2303,N_2163);
nor UO_453 (O_453,N_2027,N_2745);
or UO_454 (O_454,N_2601,N_2923);
or UO_455 (O_455,N_2097,N_2551);
nor UO_456 (O_456,N_2976,N_2439);
and UO_457 (O_457,N_2562,N_2690);
or UO_458 (O_458,N_2607,N_2741);
or UO_459 (O_459,N_2433,N_2045);
nand UO_460 (O_460,N_2977,N_2253);
nor UO_461 (O_461,N_2370,N_2877);
and UO_462 (O_462,N_2425,N_2335);
nand UO_463 (O_463,N_2391,N_2153);
nor UO_464 (O_464,N_2235,N_2179);
and UO_465 (O_465,N_2181,N_2625);
nand UO_466 (O_466,N_2591,N_2583);
nor UO_467 (O_467,N_2896,N_2313);
nor UO_468 (O_468,N_2853,N_2104);
and UO_469 (O_469,N_2014,N_2107);
nand UO_470 (O_470,N_2643,N_2488);
nand UO_471 (O_471,N_2915,N_2306);
nand UO_472 (O_472,N_2737,N_2116);
nand UO_473 (O_473,N_2357,N_2252);
nand UO_474 (O_474,N_2072,N_2791);
nand UO_475 (O_475,N_2482,N_2754);
xnor UO_476 (O_476,N_2166,N_2676);
nor UO_477 (O_477,N_2148,N_2493);
nor UO_478 (O_478,N_2827,N_2882);
and UO_479 (O_479,N_2114,N_2673);
or UO_480 (O_480,N_2485,N_2374);
or UO_481 (O_481,N_2746,N_2869);
and UO_482 (O_482,N_2774,N_2637);
nor UO_483 (O_483,N_2154,N_2284);
nor UO_484 (O_484,N_2574,N_2894);
or UO_485 (O_485,N_2940,N_2800);
xor UO_486 (O_486,N_2816,N_2242);
and UO_487 (O_487,N_2547,N_2959);
and UO_488 (O_488,N_2524,N_2823);
nor UO_489 (O_489,N_2176,N_2778);
nor UO_490 (O_490,N_2890,N_2182);
or UO_491 (O_491,N_2596,N_2952);
or UO_492 (O_492,N_2479,N_2790);
nor UO_493 (O_493,N_2787,N_2484);
nor UO_494 (O_494,N_2265,N_2895);
and UO_495 (O_495,N_2392,N_2516);
nand UO_496 (O_496,N_2430,N_2613);
nand UO_497 (O_497,N_2887,N_2957);
nor UO_498 (O_498,N_2907,N_2174);
nor UO_499 (O_499,N_2985,N_2477);
endmodule