module basic_1500_15000_2000_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1419,In_773);
or U1 (N_1,In_691,In_317);
nand U2 (N_2,In_1014,In_868);
and U3 (N_3,In_390,In_174);
nor U4 (N_4,In_357,In_1411);
nand U5 (N_5,In_240,In_764);
nand U6 (N_6,In_507,In_61);
xor U7 (N_7,In_307,In_65);
nand U8 (N_8,In_314,In_1271);
nand U9 (N_9,In_690,In_1019);
or U10 (N_10,In_740,In_566);
nand U11 (N_11,In_342,In_1316);
xor U12 (N_12,In_45,In_1072);
or U13 (N_13,In_84,In_684);
nand U14 (N_14,In_47,In_1258);
xor U15 (N_15,In_523,In_771);
nor U16 (N_16,In_186,In_1191);
nand U17 (N_17,In_155,In_1209);
xor U18 (N_18,In_1284,In_1350);
nor U19 (N_19,In_1385,In_933);
nor U20 (N_20,In_264,In_511);
nand U21 (N_21,In_51,In_1043);
or U22 (N_22,In_774,In_1124);
nor U23 (N_23,In_949,In_1178);
and U24 (N_24,In_1206,In_1245);
or U25 (N_25,In_262,In_627);
nand U26 (N_26,In_896,In_945);
nand U27 (N_27,In_145,In_620);
and U28 (N_28,In_1467,In_369);
nor U29 (N_29,In_1370,In_501);
nor U30 (N_30,In_88,In_841);
or U31 (N_31,In_254,In_290);
and U32 (N_32,In_1255,In_237);
or U33 (N_33,In_1098,In_1495);
nor U34 (N_34,In_578,In_179);
or U35 (N_35,In_1488,In_15);
or U36 (N_36,In_1490,In_1464);
and U37 (N_37,In_499,In_1219);
nand U38 (N_38,In_1131,In_666);
and U39 (N_39,In_132,In_883);
xnor U40 (N_40,In_1094,In_696);
and U41 (N_41,In_834,In_862);
or U42 (N_42,In_393,In_635);
and U43 (N_43,In_99,In_746);
or U44 (N_44,In_1026,In_579);
nand U45 (N_45,In_376,In_1185);
or U46 (N_46,In_1189,In_526);
nand U47 (N_47,In_648,In_1149);
and U48 (N_48,In_1242,In_1067);
xnor U49 (N_49,In_1312,In_38);
nor U50 (N_50,In_1355,In_86);
nor U51 (N_51,In_412,In_1384);
or U52 (N_52,In_819,In_508);
nor U53 (N_53,In_983,In_1274);
and U54 (N_54,In_982,In_1166);
or U55 (N_55,In_599,In_1364);
nand U56 (N_56,In_612,In_426);
or U57 (N_57,In_812,In_46);
nand U58 (N_58,In_52,In_1346);
or U59 (N_59,In_717,In_815);
and U60 (N_60,In_611,In_1367);
nor U61 (N_61,In_276,In_960);
and U62 (N_62,In_1028,In_1273);
and U63 (N_63,In_795,In_1418);
or U64 (N_64,In_441,In_804);
nor U65 (N_65,In_452,In_233);
nand U66 (N_66,In_486,In_837);
nor U67 (N_67,In_1328,In_692);
or U68 (N_68,In_202,In_545);
nor U69 (N_69,In_655,In_1058);
nor U70 (N_70,In_1222,In_496);
or U71 (N_71,In_497,In_1243);
nand U72 (N_72,In_219,In_249);
or U73 (N_73,In_1008,In_225);
nand U74 (N_74,In_1290,In_1383);
nand U75 (N_75,In_586,In_934);
nand U76 (N_76,In_871,In_1204);
or U77 (N_77,In_251,In_451);
xnor U78 (N_78,In_208,In_852);
nor U79 (N_79,In_1237,In_1445);
and U80 (N_80,In_741,In_1382);
nor U81 (N_81,In_447,In_1038);
nand U82 (N_82,In_1494,In_1076);
or U83 (N_83,In_201,In_79);
nor U84 (N_84,In_543,In_114);
or U85 (N_85,In_955,In_1037);
nor U86 (N_86,In_198,In_231);
and U87 (N_87,In_1186,In_937);
or U88 (N_88,In_374,In_415);
nor U89 (N_89,In_260,In_600);
nor U90 (N_90,In_115,In_454);
nand U91 (N_91,In_414,In_375);
nor U92 (N_92,In_1205,In_1175);
nor U93 (N_93,In_978,In_320);
and U94 (N_94,In_1087,In_1184);
xnor U95 (N_95,In_844,In_652);
xor U96 (N_96,In_1121,In_793);
xnor U97 (N_97,In_248,In_222);
and U98 (N_98,In_1262,In_1250);
nand U99 (N_99,In_50,In_707);
and U100 (N_100,In_212,In_998);
nor U101 (N_101,In_918,In_1065);
and U102 (N_102,In_556,In_1128);
nor U103 (N_103,In_1403,In_1200);
nand U104 (N_104,In_1342,In_1196);
nor U105 (N_105,In_581,In_951);
or U106 (N_106,In_873,In_1224);
nand U107 (N_107,In_1289,In_3);
xnor U108 (N_108,In_784,In_345);
and U109 (N_109,In_801,In_528);
nand U110 (N_110,In_1305,In_197);
and U111 (N_111,In_990,In_1152);
or U112 (N_112,In_806,In_271);
nand U113 (N_113,In_498,In_1343);
or U114 (N_114,In_350,In_470);
nand U115 (N_115,In_823,In_568);
nand U116 (N_116,In_628,In_29);
nand U117 (N_117,In_794,In_619);
nor U118 (N_118,In_1122,In_298);
or U119 (N_119,In_365,In_129);
and U120 (N_120,In_433,In_985);
nand U121 (N_121,In_315,In_1260);
nand U122 (N_122,In_1077,In_825);
or U123 (N_123,In_1234,In_931);
nand U124 (N_124,In_884,In_1448);
or U125 (N_125,In_1107,In_716);
nand U126 (N_126,In_610,In_1127);
nand U127 (N_127,In_1155,In_58);
xor U128 (N_128,In_966,In_1414);
xor U129 (N_129,In_623,In_778);
nor U130 (N_130,In_100,In_495);
and U131 (N_131,In_370,In_1352);
or U132 (N_132,In_5,In_553);
nand U133 (N_133,In_941,In_89);
xor U134 (N_134,In_1060,In_954);
and U135 (N_135,In_1435,In_833);
xnor U136 (N_136,In_715,In_668);
or U137 (N_137,In_807,In_172);
and U138 (N_138,In_205,In_1432);
and U139 (N_139,In_190,In_1389);
and U140 (N_140,In_363,In_780);
and U141 (N_141,In_661,In_540);
or U142 (N_142,In_26,In_10);
xor U143 (N_143,In_324,In_762);
nand U144 (N_144,In_602,In_743);
and U145 (N_145,In_1375,In_232);
or U146 (N_146,In_269,In_171);
nand U147 (N_147,In_176,In_263);
and U148 (N_148,In_257,In_554);
nand U149 (N_149,In_798,In_953);
or U150 (N_150,In_1154,In_814);
or U151 (N_151,In_1463,In_512);
nand U152 (N_152,In_895,In_775);
or U153 (N_153,In_1397,In_1335);
xnor U154 (N_154,In_419,In_713);
xnor U155 (N_155,In_721,In_981);
and U156 (N_156,In_1169,In_1408);
or U157 (N_157,In_1079,In_428);
nor U158 (N_158,In_117,In_1442);
and U159 (N_159,In_1415,In_1459);
and U160 (N_160,In_407,In_702);
or U161 (N_161,In_988,In_548);
or U162 (N_162,In_195,In_322);
xor U163 (N_163,In_1150,In_538);
xnor U164 (N_164,In_241,In_1135);
nor U165 (N_165,In_289,In_1317);
xor U166 (N_166,In_1269,In_160);
nor U167 (N_167,In_1251,In_1130);
xnor U168 (N_168,In_353,In_323);
or U169 (N_169,In_855,In_976);
nand U170 (N_170,In_1226,In_653);
nor U171 (N_171,In_839,In_1091);
and U172 (N_172,In_1341,In_261);
xor U173 (N_173,In_1119,In_1147);
nand U174 (N_174,In_491,In_1171);
and U175 (N_175,In_539,In_166);
or U176 (N_176,In_911,In_239);
and U177 (N_177,In_1148,In_275);
xor U178 (N_178,In_564,In_20);
nand U179 (N_179,In_1410,In_1460);
and U180 (N_180,In_1322,In_1081);
nor U181 (N_181,In_96,In_877);
or U182 (N_182,In_1436,In_71);
nand U183 (N_183,In_126,In_1202);
or U184 (N_184,In_1301,In_316);
or U185 (N_185,In_971,In_584);
xnor U186 (N_186,In_141,In_673);
nand U187 (N_187,In_739,In_1314);
nand U188 (N_188,In_979,In_1489);
xor U189 (N_189,In_562,In_786);
xor U190 (N_190,In_722,In_1480);
nor U191 (N_191,In_676,In_1208);
xor U192 (N_192,In_223,In_1310);
and U193 (N_193,In_847,In_1444);
xnor U194 (N_194,In_207,In_9);
and U195 (N_195,In_1376,In_247);
or U196 (N_196,In_494,In_952);
nand U197 (N_197,In_1474,In_133);
nand U198 (N_198,In_519,In_296);
nor U199 (N_199,In_1032,In_1398);
nor U200 (N_200,In_1381,In_1159);
nor U201 (N_201,In_1438,In_1344);
or U202 (N_202,In_555,In_481);
or U203 (N_203,In_1306,In_885);
and U204 (N_204,In_905,In_607);
and U205 (N_205,In_1325,In_1421);
nand U206 (N_206,In_973,In_678);
or U207 (N_207,In_700,In_416);
xor U208 (N_208,In_351,In_476);
nand U209 (N_209,In_1017,In_1394);
xor U210 (N_210,In_980,In_752);
nor U211 (N_211,In_4,In_347);
nand U212 (N_212,In_387,In_464);
and U213 (N_213,In_1391,In_803);
xnor U214 (N_214,In_1327,In_425);
xnor U215 (N_215,In_518,In_14);
xnor U216 (N_216,In_1434,In_571);
xor U217 (N_217,In_704,In_790);
nor U218 (N_218,In_867,In_649);
nor U219 (N_219,In_992,In_457);
nand U220 (N_220,In_685,In_932);
nand U221 (N_221,In_354,In_760);
nand U222 (N_222,In_74,In_273);
xor U223 (N_223,In_295,In_1086);
nand U224 (N_224,In_448,In_1221);
xor U225 (N_225,In_392,In_1275);
nor U226 (N_226,In_708,In_339);
nor U227 (N_227,In_128,In_1496);
nor U228 (N_228,In_644,In_948);
or U229 (N_229,In_1347,In_1142);
nand U230 (N_230,In_604,In_1188);
nor U231 (N_231,In_1092,In_404);
nand U232 (N_232,In_1003,In_168);
or U233 (N_233,In_820,In_830);
xor U234 (N_234,In_621,In_977);
nand U235 (N_235,In_1264,In_206);
nor U236 (N_236,In_935,In_697);
and U237 (N_237,In_576,In_443);
or U238 (N_238,In_183,In_367);
xnor U239 (N_239,In_1299,In_791);
and U240 (N_240,In_626,In_410);
nor U241 (N_241,In_48,In_734);
or U242 (N_242,In_592,In_1272);
and U243 (N_243,In_349,In_1492);
nand U244 (N_244,In_974,In_736);
or U245 (N_245,In_32,In_882);
nand U246 (N_246,In_595,In_23);
nand U247 (N_247,In_1268,In_1084);
xor U248 (N_248,In_1104,In_1402);
nor U249 (N_249,In_1454,In_11);
and U250 (N_250,In_1493,In_665);
xnor U251 (N_251,In_1099,In_440);
and U252 (N_252,In_118,In_711);
xnor U253 (N_253,In_40,In_371);
nor U254 (N_254,In_881,In_487);
nand U255 (N_255,In_865,In_738);
nor U256 (N_256,In_259,In_570);
nand U257 (N_257,In_1074,In_783);
nor U258 (N_258,In_1416,In_929);
xor U259 (N_259,In_200,In_1198);
xor U260 (N_260,In_102,In_1471);
xnor U261 (N_261,In_1027,In_1180);
or U262 (N_262,In_104,In_1320);
xnor U263 (N_263,In_899,In_719);
xnor U264 (N_264,In_1238,In_897);
and U265 (N_265,In_593,In_334);
and U266 (N_266,In_28,In_1045);
or U267 (N_267,In_688,In_733);
nor U268 (N_268,In_1083,In_758);
or U269 (N_269,In_826,In_1283);
xnor U270 (N_270,In_56,In_116);
or U271 (N_271,In_327,In_16);
and U272 (N_272,In_1348,In_854);
or U273 (N_273,In_749,In_664);
xnor U274 (N_274,In_1151,In_348);
nor U275 (N_275,In_185,In_1024);
xnor U276 (N_276,In_1430,In_699);
nor U277 (N_277,In_891,In_710);
xor U278 (N_278,In_490,In_645);
and U279 (N_279,In_1117,In_1016);
xor U280 (N_280,In_226,In_557);
xnor U281 (N_281,In_777,In_583);
xor U282 (N_282,In_1143,In_1357);
nand U283 (N_283,In_1013,In_1109);
nand U284 (N_284,In_580,In_671);
xnor U285 (N_285,In_636,In_308);
and U286 (N_286,In_304,In_506);
xor U287 (N_287,In_106,In_912);
and U288 (N_288,In_377,In_1120);
nor U289 (N_289,In_1247,In_1168);
xor U290 (N_290,In_559,In_1007);
xor U291 (N_291,In_1363,In_164);
nand U292 (N_292,In_438,In_1177);
and U293 (N_293,In_196,In_389);
nor U294 (N_294,In_284,In_1176);
nor U295 (N_295,In_12,In_394);
nand U296 (N_296,In_516,In_714);
or U297 (N_297,In_277,In_41);
xor U298 (N_298,In_1270,In_679);
and U299 (N_299,In_1125,In_832);
nand U300 (N_300,N_292,N_80);
or U301 (N_301,N_91,N_84);
and U302 (N_302,In_787,In_1246);
or U303 (N_303,In_1484,N_182);
xnor U304 (N_304,In_329,N_221);
nor U305 (N_305,In_385,N_70);
or U306 (N_306,In_1052,In_890);
and U307 (N_307,In_1431,In_1387);
and U308 (N_308,N_126,In_422);
xor U309 (N_309,In_396,In_1374);
or U310 (N_310,In_169,In_913);
nand U311 (N_311,In_864,In_346);
or U312 (N_312,In_140,In_1473);
nor U313 (N_313,In_1164,In_95);
nor U314 (N_314,In_657,In_1211);
nor U315 (N_315,In_811,N_138);
xor U316 (N_316,N_115,In_565);
nor U317 (N_317,In_192,In_70);
nand U318 (N_318,In_544,N_67);
or U319 (N_319,N_106,In_417);
and U320 (N_320,In_55,N_108);
nand U321 (N_321,In_869,In_502);
xor U322 (N_322,N_242,In_1167);
nand U323 (N_323,In_472,N_142);
and U324 (N_324,In_962,In_1115);
xor U325 (N_325,In_361,N_119);
nand U326 (N_326,In_677,In_898);
nand U327 (N_327,In_1441,N_214);
nand U328 (N_328,In_154,In_845);
nor U329 (N_329,N_227,In_123);
or U330 (N_330,N_20,In_1009);
xnor U331 (N_331,In_378,In_789);
and U332 (N_332,In_744,In_359);
xor U333 (N_333,In_573,In_401);
xnor U334 (N_334,N_68,In_73);
nand U335 (N_335,In_191,In_936);
or U336 (N_336,In_991,In_1034);
xor U337 (N_337,In_770,In_513);
and U338 (N_338,In_1498,In_1059);
xor U339 (N_339,In_879,In_634);
and U340 (N_340,In_309,In_1371);
nand U341 (N_341,In_69,In_1068);
or U342 (N_342,N_52,In_87);
and U343 (N_343,In_996,In_282);
and U344 (N_344,In_799,In_1455);
nor U345 (N_345,In_330,N_192);
xnor U346 (N_346,In_310,In_875);
and U347 (N_347,N_45,In_624);
nor U348 (N_348,In_243,In_1422);
or U349 (N_349,In_1229,In_950);
nand U350 (N_350,N_161,In_221);
or U351 (N_351,In_209,N_27);
nor U352 (N_352,In_1427,In_689);
and U353 (N_353,In_31,In_432);
nor U354 (N_354,N_97,In_63);
xor U355 (N_355,In_1497,In_910);
or U356 (N_356,In_459,In_1302);
xor U357 (N_357,In_280,N_61);
or U358 (N_358,In_1349,N_36);
nor U359 (N_359,In_1286,N_87);
nand U360 (N_360,In_340,In_127);
nor U361 (N_361,In_13,N_240);
and U362 (N_362,In_1182,In_1042);
nor U363 (N_363,In_1281,In_999);
or U364 (N_364,In_737,N_195);
and U365 (N_365,In_8,N_265);
and U366 (N_366,In_542,In_928);
nand U367 (N_367,In_60,In_134);
and U368 (N_368,In_630,In_1409);
nor U369 (N_369,In_1136,In_1318);
xor U370 (N_370,In_917,N_260);
nor U371 (N_371,In_161,In_1429);
xor U372 (N_372,In_81,In_1323);
nor U373 (N_373,In_420,In_747);
or U374 (N_374,In_148,N_2);
or U375 (N_375,In_136,In_940);
or U376 (N_376,N_103,In_22);
and U377 (N_377,In_54,In_1071);
and U378 (N_378,In_816,N_187);
or U379 (N_379,In_616,In_1358);
nor U380 (N_380,In_19,In_1361);
nand U381 (N_381,N_213,In_1174);
or U382 (N_382,In_458,In_1156);
and U383 (N_383,In_442,In_1103);
and U384 (N_384,N_148,In_105);
nand U385 (N_385,In_533,In_838);
nor U386 (N_386,In_709,In_745);
and U387 (N_387,In_321,In_1025);
nand U388 (N_388,In_532,In_1362);
xor U389 (N_389,In_144,N_135);
nor U390 (N_390,In_1239,N_197);
and U391 (N_391,In_391,N_244);
and U392 (N_392,In_83,In_1187);
xor U393 (N_393,N_92,N_13);
and U394 (N_394,In_757,In_1468);
and U395 (N_395,In_124,In_587);
or U396 (N_396,N_122,N_226);
and U397 (N_397,N_280,N_165);
nand U398 (N_398,In_646,In_215);
or U399 (N_399,N_129,In_475);
nor U400 (N_400,In_510,In_1139);
nand U401 (N_401,N_58,N_145);
xnor U402 (N_402,In_255,N_180);
nor U403 (N_403,In_914,N_140);
nand U404 (N_404,In_920,In_731);
nor U405 (N_405,In_1388,N_35);
nor U406 (N_406,In_1378,N_210);
xnor U407 (N_407,In_843,In_776);
xor U408 (N_408,In_246,N_73);
or U409 (N_409,In_1292,In_480);
xor U410 (N_410,In_466,In_228);
and U411 (N_411,In_1450,In_1369);
nor U412 (N_412,In_229,N_201);
or U413 (N_413,N_264,In_1308);
and U414 (N_414,In_287,In_756);
xnor U415 (N_415,In_408,In_1257);
or U416 (N_416,In_449,In_68);
and U417 (N_417,N_37,In_1057);
or U418 (N_418,N_204,In_1088);
and U419 (N_419,In_887,In_1105);
or U420 (N_420,N_83,In_1424);
nor U421 (N_421,In_437,In_424);
nand U422 (N_422,In_159,In_1053);
nor U423 (N_423,N_215,In_325);
and U424 (N_424,In_362,N_263);
and U425 (N_425,In_633,In_529);
nor U426 (N_426,In_1102,In_641);
nor U427 (N_427,In_1232,In_266);
and U428 (N_428,In_1324,N_33);
and U429 (N_429,In_640,In_639);
or U430 (N_430,N_297,N_123);
nor U431 (N_431,N_271,In_109);
xnor U432 (N_432,In_384,N_205);
nor U433 (N_433,In_622,In_840);
and U434 (N_434,In_292,In_492);
or U435 (N_435,In_824,In_817);
nor U436 (N_436,N_216,In_1465);
xor U437 (N_437,In_101,In_1339);
nor U438 (N_438,In_268,In_1218);
xor U439 (N_439,In_629,N_171);
xnor U440 (N_440,In_66,In_561);
nor U441 (N_441,In_1303,In_1288);
and U442 (N_442,In_409,In_286);
xor U443 (N_443,In_1261,N_40);
xnor U444 (N_444,In_984,In_1080);
nor U445 (N_445,N_247,In_227);
nor U446 (N_446,In_379,In_683);
or U447 (N_447,In_503,N_34);
nor U448 (N_448,In_693,In_727);
or U449 (N_449,N_291,N_199);
nand U450 (N_450,In_444,N_189);
nor U451 (N_451,In_326,N_160);
nor U452 (N_452,In_318,N_232);
nor U453 (N_453,In_958,In_1108);
nand U454 (N_454,In_1210,In_1447);
and U455 (N_455,In_252,In_1356);
nor U456 (N_456,N_258,N_71);
and U457 (N_457,In_1417,In_366);
nor U458 (N_458,In_274,In_919);
nor U459 (N_459,N_253,In_767);
nor U460 (N_460,In_285,N_74);
xnor U461 (N_461,In_631,In_151);
xnor U462 (N_462,In_759,In_368);
nor U463 (N_463,In_1300,In_297);
and U464 (N_464,N_65,In_244);
xor U465 (N_465,N_136,In_1033);
or U466 (N_466,In_1138,In_849);
nand U467 (N_467,In_725,In_1097);
xnor U468 (N_468,In_6,In_1179);
and U469 (N_469,In_792,N_17);
or U470 (N_470,In_1070,In_1401);
or U471 (N_471,N_155,In_1157);
and U472 (N_472,In_352,In_1137);
and U473 (N_473,N_49,In_220);
and U474 (N_474,In_706,In_900);
or U475 (N_475,In_333,In_698);
or U476 (N_476,In_1276,In_1018);
xnor U477 (N_477,In_413,N_38);
or U478 (N_478,N_186,In_450);
xnor U479 (N_479,In_279,In_1100);
nand U480 (N_480,N_149,In_281);
xor U481 (N_481,N_235,N_29);
xor U482 (N_482,In_802,In_430);
xor U483 (N_483,In_1051,In_1332);
nand U484 (N_484,In_97,In_204);
xnor U485 (N_485,In_153,N_94);
or U486 (N_486,In_902,In_122);
nand U487 (N_487,In_1395,In_1153);
nand U488 (N_488,In_78,In_1015);
or U489 (N_489,N_162,N_273);
nand U490 (N_490,In_959,In_567);
nor U491 (N_491,In_563,In_146);
nor U492 (N_492,In_924,In_167);
nand U493 (N_493,In_1295,N_223);
xnor U494 (N_494,In_1047,In_360);
xor U495 (N_495,N_93,N_274);
and U496 (N_496,In_1129,N_241);
or U497 (N_497,In_575,In_720);
or U498 (N_498,N_151,In_1315);
xnor U499 (N_499,N_251,In_1066);
or U500 (N_500,In_1112,In_474);
or U501 (N_501,In_1197,In_1462);
nand U502 (N_502,In_1337,N_261);
nand U503 (N_503,N_64,N_218);
nor U504 (N_504,In_469,In_796);
nand U505 (N_505,In_779,In_866);
xor U506 (N_506,N_50,In_970);
and U507 (N_507,N_228,In_829);
xor U508 (N_508,N_219,In_788);
nand U509 (N_509,In_606,In_1050);
nor U510 (N_510,N_114,In_43);
nor U511 (N_511,In_894,In_637);
or U512 (N_512,In_1039,In_388);
nor U513 (N_513,In_1365,In_431);
and U514 (N_514,N_113,In_256);
nor U515 (N_515,In_312,In_654);
or U516 (N_516,In_1133,In_272);
or U517 (N_517,In_718,In_1475);
and U518 (N_518,In_111,In_730);
or U519 (N_519,In_582,In_601);
nor U520 (N_520,In_489,In_965);
xor U521 (N_521,In_1194,N_296);
and U522 (N_522,In_681,N_179);
nor U523 (N_523,In_288,In_1022);
and U524 (N_524,In_1160,In_597);
and U525 (N_525,N_238,In_44);
nand U526 (N_526,In_1297,In_467);
or U527 (N_527,In_957,N_30);
or U528 (N_528,In_380,In_76);
nand U529 (N_529,In_1114,In_33);
and U530 (N_530,In_372,In_300);
xor U531 (N_531,N_267,In_1440);
nand U532 (N_532,In_1291,In_230);
nor U533 (N_533,In_886,N_154);
and U534 (N_534,In_1172,In_520);
nand U535 (N_535,In_525,N_15);
or U536 (N_536,In_35,In_1005);
nor U537 (N_537,N_104,In_460);
nand U538 (N_538,In_1061,In_1330);
xnor U539 (N_539,In_1132,In_921);
or U540 (N_540,In_157,N_57);
nor U541 (N_541,In_1111,N_254);
nor U542 (N_542,In_1457,N_51);
nand U543 (N_543,In_850,In_1217);
nor U544 (N_544,In_1134,N_53);
nor U545 (N_545,In_113,In_427);
and U546 (N_546,In_180,In_1491);
and U547 (N_547,N_268,In_853);
nor U548 (N_548,In_1446,In_662);
or U549 (N_549,N_48,In_625);
nand U550 (N_550,In_1021,In_753);
or U551 (N_551,N_21,N_105);
nand U552 (N_552,In_613,In_1461);
or U553 (N_553,In_1011,In_1334);
nor U554 (N_554,In_37,In_436);
nand U555 (N_555,In_1235,In_483);
nand U556 (N_556,In_1449,In_930);
or U557 (N_557,In_986,In_963);
and U558 (N_558,In_828,In_1201);
xnor U559 (N_559,In_1340,In_1118);
and U560 (N_560,In_1307,In_1106);
nand U561 (N_561,N_159,In_1096);
nand U562 (N_562,N_281,N_252);
and U563 (N_563,In_1482,N_28);
and U564 (N_564,N_76,In_614);
xnor U565 (N_565,In_397,In_1478);
xnor U566 (N_566,N_42,In_336);
xnor U567 (N_567,In_944,In_1046);
nand U568 (N_568,In_165,In_1426);
nand U569 (N_569,N_172,N_157);
and U570 (N_570,N_224,In_993);
and U571 (N_571,In_1423,In_906);
nand U572 (N_572,In_1195,N_121);
or U573 (N_573,In_859,N_209);
nor U574 (N_574,In_210,In_943);
or U575 (N_575,In_1359,In_189);
nor U576 (N_576,In_909,In_478);
xor U577 (N_577,In_382,In_813);
nor U578 (N_578,In_1279,In_549);
nor U579 (N_579,In_735,N_112);
nand U580 (N_580,In_1095,N_208);
nand U581 (N_581,In_64,In_1486);
nor U582 (N_582,In_17,N_298);
nor U583 (N_583,N_118,N_134);
or U584 (N_584,In_632,In_1223);
and U585 (N_585,N_18,In_1101);
and U586 (N_586,In_400,N_8);
nand U587 (N_587,In_1123,In_972);
and U588 (N_588,In_669,In_1377);
and U589 (N_589,In_1,In_1145);
nor U590 (N_590,In_213,N_299);
xnor U591 (N_591,In_27,In_343);
nand U592 (N_592,In_1451,In_181);
nand U593 (N_593,In_62,N_288);
and U594 (N_594,In_7,In_103);
and U595 (N_595,In_822,In_585);
nor U596 (N_596,N_193,In_769);
xnor U597 (N_597,In_651,In_821);
or U598 (N_598,In_535,N_294);
and U599 (N_599,In_121,In_265);
or U600 (N_600,N_435,N_554);
nor U601 (N_601,In_728,N_438);
nand U602 (N_602,In_915,N_266);
nor U603 (N_603,In_732,N_545);
nand U604 (N_604,In_463,N_169);
and U605 (N_605,N_340,N_415);
xor U606 (N_606,N_414,In_650);
nor U607 (N_607,In_1386,In_541);
xor U608 (N_608,N_550,In_1207);
or U609 (N_609,N_31,N_315);
nor U610 (N_610,In_30,In_1085);
or U611 (N_611,N_525,N_400);
and U612 (N_612,N_124,In_618);
or U613 (N_613,In_617,In_199);
nand U614 (N_614,In_1165,In_435);
xor U615 (N_615,N_436,In_818);
and U616 (N_616,In_1041,In_997);
xnor U617 (N_617,In_1055,In_1393);
or U618 (N_618,In_291,In_551);
nand U619 (N_619,N_527,N_537);
xnor U620 (N_620,N_334,N_495);
xnor U621 (N_621,N_568,In_482);
xor U622 (N_622,In_218,N_546);
nor U623 (N_623,In_547,In_682);
or U624 (N_624,N_330,In_1230);
nor U625 (N_625,N_245,N_200);
nor U626 (N_626,In_406,N_146);
and U627 (N_627,In_1241,N_289);
or U628 (N_628,N_77,In_137);
xor U629 (N_629,N_499,N_358);
nand U630 (N_630,In_785,In_761);
or U631 (N_631,N_454,N_451);
or U632 (N_632,In_515,N_338);
and U633 (N_633,N_314,In_1090);
nand U634 (N_634,In_1485,N_99);
and U635 (N_635,In_615,In_294);
nand U636 (N_636,In_1333,In_1476);
or U637 (N_637,In_1063,In_1285);
xor U638 (N_638,In_465,N_5);
nor U639 (N_639,In_1287,In_34);
xnor U640 (N_640,In_1373,N_486);
and U641 (N_641,N_54,N_446);
xnor U642 (N_642,In_723,N_56);
nand U643 (N_643,N_236,N_379);
or U644 (N_644,In_1216,In_338);
xor U645 (N_645,In_80,In_1439);
nand U646 (N_646,In_1146,N_96);
xor U647 (N_647,N_455,N_86);
or U648 (N_648,In_946,N_353);
nor U649 (N_649,In_1470,N_403);
or U650 (N_650,In_1089,N_212);
or U651 (N_651,N_181,N_567);
nand U652 (N_652,N_89,In_1023);
nand U653 (N_653,N_540,In_302);
nand U654 (N_654,In_39,N_468);
xnor U655 (N_655,In_1437,N_283);
nor U656 (N_656,In_687,N_588);
xnor U657 (N_657,In_1256,In_1282);
nor U658 (N_658,N_392,N_395);
and U659 (N_659,In_552,In_178);
nor U660 (N_660,In_524,N_85);
or U661 (N_661,N_262,N_300);
and U662 (N_662,In_670,N_66);
nor U663 (N_663,In_589,In_994);
or U664 (N_664,N_375,N_331);
nor U665 (N_665,In_484,N_391);
nor U666 (N_666,N_350,N_198);
nor U667 (N_667,N_592,In_142);
or U668 (N_668,N_11,N_349);
or U669 (N_669,N_412,In_1183);
and U670 (N_670,N_307,N_0);
nor U671 (N_671,N_324,In_429);
and U672 (N_672,In_242,N_543);
or U673 (N_673,N_348,In_1040);
nor U674 (N_674,N_166,N_559);
nor U675 (N_675,In_125,In_119);
nor U676 (N_676,In_1469,In_139);
or U677 (N_677,N_257,N_459);
nand U678 (N_678,N_595,N_585);
and U679 (N_679,In_797,In_42);
or U680 (N_680,N_259,In_1002);
nand U681 (N_681,N_491,In_1294);
xor U682 (N_682,In_1048,N_481);
nor U683 (N_683,N_359,In_184);
nor U684 (N_684,N_557,N_335);
or U685 (N_685,N_81,N_323);
or U686 (N_686,N_466,N_98);
and U687 (N_687,In_311,In_305);
or U688 (N_688,In_927,In_726);
nor U689 (N_689,N_560,N_480);
nor U690 (N_690,In_577,In_110);
and U691 (N_691,In_1407,In_609);
nand U692 (N_692,N_143,N_561);
or U693 (N_693,N_482,In_782);
nor U694 (N_694,N_309,In_488);
nor U695 (N_695,N_7,N_164);
xor U696 (N_696,In_872,N_328);
nor U697 (N_697,N_347,In_203);
nand U698 (N_698,In_1392,In_1326);
nor U699 (N_699,N_490,In_1481);
nand U700 (N_700,N_133,In_1056);
xor U701 (N_701,N_426,In_1366);
nand U702 (N_702,N_329,In_901);
xnor U703 (N_703,N_575,N_471);
xor U704 (N_704,N_496,In_1190);
or U705 (N_705,In_835,In_860);
and U706 (N_706,In_194,In_1360);
xor U707 (N_707,In_893,N_423);
xor U708 (N_708,In_188,N_220);
or U709 (N_709,N_248,N_178);
or U710 (N_710,N_321,In_527);
and U711 (N_711,N_333,N_107);
or U712 (N_712,In_590,N_386);
and U713 (N_713,N_472,In_591);
or U714 (N_714,In_1400,N_470);
xnor U715 (N_715,N_336,N_373);
nor U716 (N_716,N_494,In_1263);
xor U717 (N_717,N_387,N_487);
and U718 (N_718,In_750,In_1173);
or U719 (N_719,N_111,In_926);
and U720 (N_720,N_581,N_357);
nand U721 (N_721,In_1331,In_162);
or U722 (N_722,N_552,N_507);
xnor U723 (N_723,N_249,In_303);
xor U724 (N_724,N_467,In_904);
nand U725 (N_725,In_358,N_553);
or U726 (N_726,In_674,N_492);
nor U727 (N_727,In_1472,N_312);
xor U728 (N_728,N_506,In_158);
nor U729 (N_729,N_246,In_91);
xnor U730 (N_730,N_463,N_429);
xnor U731 (N_731,In_1181,N_82);
xnor U732 (N_732,In_49,In_341);
nor U733 (N_733,N_449,In_1313);
nand U734 (N_734,N_305,N_32);
or U735 (N_735,N_503,In_594);
or U736 (N_736,N_41,In_82);
xnor U737 (N_737,N_302,In_331);
xor U738 (N_738,N_243,N_59);
or U739 (N_739,N_184,In_1144);
or U740 (N_740,N_410,N_176);
xnor U741 (N_741,N_341,In_439);
nand U742 (N_742,N_12,N_202);
nand U743 (N_743,In_143,In_1329);
xor U744 (N_744,In_182,N_275);
nor U745 (N_745,N_109,N_79);
nand U746 (N_746,N_548,N_422);
xor U747 (N_747,In_987,In_238);
and U748 (N_748,In_471,In_253);
or U749 (N_749,N_39,In_293);
or U750 (N_750,N_88,N_368);
or U751 (N_751,In_1227,In_92);
nor U752 (N_752,In_0,N_437);
or U753 (N_753,In_810,In_1477);
and U754 (N_754,In_1390,N_456);
nor U755 (N_755,In_656,N_117);
nor U756 (N_756,In_77,In_536);
xnor U757 (N_757,N_43,In_234);
or U758 (N_758,In_765,N_485);
nor U759 (N_759,In_135,N_318);
nor U760 (N_760,In_1254,In_1113);
or U761 (N_761,In_173,In_112);
or U762 (N_762,In_907,N_352);
or U763 (N_763,N_406,N_377);
nand U764 (N_764,N_389,N_397);
nor U765 (N_765,In_75,N_443);
nand U766 (N_766,N_19,In_1452);
xnor U767 (N_767,In_858,In_1345);
nand U768 (N_768,In_550,N_16);
or U769 (N_769,N_177,In_660);
nand U770 (N_770,N_308,N_398);
nor U771 (N_771,In_1428,N_120);
or U772 (N_772,N_256,In_72);
and U773 (N_773,In_537,N_519);
xnor U774 (N_774,N_295,In_445);
nor U775 (N_775,N_473,In_479);
or U776 (N_776,N_589,N_520);
nor U777 (N_777,In_964,In_574);
nand U778 (N_778,N_130,N_497);
nand U779 (N_779,N_69,N_380);
and U780 (N_780,In_1396,N_325);
nor U781 (N_781,In_505,In_1212);
xnor U782 (N_782,N_584,N_404);
nand U783 (N_783,N_322,N_234);
and U784 (N_784,In_751,N_441);
nand U785 (N_785,N_564,In_504);
nor U786 (N_786,In_1249,In_1420);
or U787 (N_787,N_206,N_277);
and U788 (N_788,In_1082,N_413);
nor U789 (N_789,N_222,In_1203);
nand U790 (N_790,In_968,N_382);
or U791 (N_791,N_425,N_371);
xor U792 (N_792,In_156,In_403);
or U793 (N_793,In_608,N_110);
xor U794 (N_794,N_346,In_521);
nand U795 (N_795,N_569,In_1244);
nand U796 (N_796,N_477,N_479);
and U797 (N_797,N_444,In_1433);
nor U798 (N_798,N_424,N_529);
nor U799 (N_799,In_364,N_378);
and U800 (N_800,N_583,In_1304);
or U801 (N_801,In_961,N_396);
and U802 (N_802,N_551,In_398);
nor U803 (N_803,N_326,N_526);
xnor U804 (N_804,N_282,N_229);
nor U805 (N_805,In_1252,In_851);
or U806 (N_806,In_938,N_465);
or U807 (N_807,In_546,N_417);
or U808 (N_808,In_1404,N_515);
nand U809 (N_809,In_1075,In_130);
and U810 (N_810,In_1029,In_663);
xnor U811 (N_811,In_373,N_116);
nand U812 (N_812,N_150,In_211);
nand U813 (N_813,In_1010,In_808);
nand U814 (N_814,In_1215,In_1240);
or U815 (N_815,In_1158,In_863);
nand U816 (N_816,In_381,N_539);
or U817 (N_817,In_236,N_90);
or U818 (N_818,In_455,N_365);
or U819 (N_819,In_1035,In_680);
xnor U820 (N_820,N_460,In_405);
and U821 (N_821,N_60,N_535);
nand U822 (N_822,In_170,N_174);
or U823 (N_823,N_284,N_279);
or U824 (N_824,In_1353,In_1162);
xnor U825 (N_825,In_337,In_908);
xnor U826 (N_826,N_319,N_469);
xor U827 (N_827,In_705,In_1253);
and U828 (N_828,N_390,N_144);
and U829 (N_829,In_861,In_24);
or U830 (N_830,In_831,In_1443);
or U831 (N_831,In_1110,In_878);
nand U832 (N_832,In_1266,In_313);
or U833 (N_833,In_108,N_303);
nor U834 (N_834,In_1012,N_316);
or U835 (N_835,In_344,In_500);
and U836 (N_836,N_139,N_44);
xor U837 (N_837,In_1406,In_596);
or U838 (N_838,In_1336,In_989);
and U839 (N_839,N_137,N_453);
or U840 (N_840,In_667,In_1458);
xnor U841 (N_841,N_131,N_225);
xor U842 (N_842,N_191,N_9);
nand U843 (N_843,In_947,In_1004);
and U844 (N_844,N_533,N_514);
nand U845 (N_845,In_755,In_995);
nand U846 (N_846,N_427,N_522);
xnor U847 (N_847,In_149,N_369);
nor U848 (N_848,In_395,N_163);
xnor U849 (N_849,N_489,N_419);
nor U850 (N_850,In_1380,In_922);
and U851 (N_851,In_1049,N_464);
xnor U852 (N_852,In_530,In_1487);
nor U853 (N_853,N_306,In_703);
xnor U854 (N_854,In_766,N_547);
or U855 (N_855,N_10,N_313);
nand U856 (N_856,In_418,N_597);
nor U857 (N_857,N_337,N_3);
nor U858 (N_858,N_332,N_428);
xnor U859 (N_859,N_183,In_772);
and U860 (N_860,In_1338,N_408);
nand U861 (N_861,N_293,In_1225);
or U862 (N_862,N_175,N_483);
or U863 (N_863,In_355,N_102);
nor U864 (N_864,N_518,In_572);
and U865 (N_865,N_141,N_211);
nand U866 (N_866,In_748,N_310);
or U867 (N_867,In_1031,In_848);
xnor U868 (N_868,N_230,N_433);
xnor U869 (N_869,N_528,In_107);
nand U870 (N_870,N_383,In_534);
xnor U871 (N_871,In_1479,In_421);
nand U872 (N_872,In_642,In_1228);
nor U873 (N_873,In_85,In_1265);
or U874 (N_874,In_175,N_6);
and U875 (N_875,N_538,In_306);
nand U876 (N_876,N_343,N_339);
nand U877 (N_877,In_456,N_311);
or U878 (N_878,N_278,N_147);
and U879 (N_879,In_163,In_57);
xor U880 (N_880,N_269,In_468);
nand U881 (N_881,In_216,In_874);
or U882 (N_882,N_563,In_270);
and U883 (N_883,In_187,N_362);
and U884 (N_884,In_659,N_62);
or U885 (N_885,In_1379,In_245);
nor U886 (N_886,In_332,In_423);
and U887 (N_887,N_100,N_598);
and U888 (N_888,N_364,N_388);
nand U889 (N_889,In_1483,N_448);
xnor U890 (N_890,N_301,N_558);
xor U891 (N_891,In_301,N_582);
nand U892 (N_892,In_846,In_1163);
or U893 (N_893,In_150,In_217);
nand U894 (N_894,N_153,N_447);
and U895 (N_895,N_95,In_724);
nand U896 (N_896,In_1368,In_1236);
and U897 (N_897,In_138,N_393);
and U898 (N_898,In_1233,N_272);
or U899 (N_899,N_591,In_712);
xor U900 (N_900,In_93,N_644);
or U901 (N_901,N_304,N_727);
nand U902 (N_902,N_648,In_319);
or U903 (N_903,N_721,N_669);
xor U904 (N_904,N_830,N_532);
xnor U905 (N_905,In_836,N_777);
nand U906 (N_906,In_1170,In_842);
xor U907 (N_907,N_634,N_445);
nor U908 (N_908,N_128,N_320);
or U909 (N_909,In_1116,N_844);
and U910 (N_910,N_651,N_723);
nand U911 (N_911,N_642,N_824);
and U912 (N_912,N_724,N_703);
xor U913 (N_913,N_190,N_342);
and U914 (N_914,N_718,N_394);
nand U915 (N_915,In_1073,N_851);
nor U916 (N_916,N_621,N_327);
nor U917 (N_917,N_806,N_861);
nand U918 (N_918,N_594,N_746);
or U919 (N_919,N_233,N_668);
and U920 (N_920,N_630,In_1412);
xnor U921 (N_921,N_510,In_514);
nand U922 (N_922,N_617,N_803);
nor U923 (N_923,N_679,In_1248);
and U924 (N_924,N_758,N_810);
xnor U925 (N_925,N_757,N_688);
xnor U926 (N_926,N_194,N_796);
nor U927 (N_927,In_558,In_21);
or U928 (N_928,In_658,N_749);
or U929 (N_929,In_916,N_608);
nor U930 (N_930,N_363,N_25);
and U931 (N_931,N_837,In_98);
xnor U932 (N_932,N_741,N_656);
nor U933 (N_933,N_873,N_654);
or U934 (N_934,N_680,In_299);
nor U935 (N_935,N_686,N_684);
xnor U936 (N_936,N_843,N_22);
nor U937 (N_937,In_94,N_512);
nor U938 (N_938,N_794,N_505);
and U939 (N_939,In_1259,N_576);
and U940 (N_940,N_681,N_484);
or U941 (N_941,N_541,In_975);
nor U942 (N_942,N_884,In_605);
nand U943 (N_943,N_168,In_531);
xor U944 (N_944,N_834,N_743);
nand U945 (N_945,N_287,N_734);
nor U946 (N_946,N_127,N_26);
or U947 (N_947,N_891,N_693);
nor U948 (N_948,In_1093,N_629);
nor U949 (N_949,N_841,N_747);
and U950 (N_950,N_638,N_689);
nor U951 (N_951,N_890,In_969);
nand U952 (N_952,N_894,N_670);
xnor U953 (N_953,In_1267,N_709);
nor U954 (N_954,N_763,N_361);
and U955 (N_955,N_461,In_53);
or U956 (N_956,N_536,N_697);
xor U957 (N_957,N_829,N_407);
nand U958 (N_958,N_699,N_674);
or U959 (N_959,N_24,In_335);
xnor U960 (N_960,N_63,N_577);
or U961 (N_961,N_587,N_524);
or U962 (N_962,In_701,N_893);
nor U963 (N_963,N_676,N_782);
nor U964 (N_964,N_671,In_1293);
xor U965 (N_965,N_868,N_354);
xnor U966 (N_966,N_628,In_1064);
or U967 (N_967,N_870,N_852);
and U968 (N_968,N_733,N_897);
xnor U969 (N_969,N_619,N_755);
xor U970 (N_970,In_1466,N_899);
xor U971 (N_971,N_623,N_786);
and U972 (N_972,N_875,In_889);
xor U973 (N_973,N_421,In_1413);
and U974 (N_974,N_647,N_729);
nand U975 (N_975,N_690,N_839);
xor U976 (N_976,In_967,N_372);
and U977 (N_977,In_522,In_1036);
xor U978 (N_978,N_799,N_695);
or U979 (N_979,In_193,N_687);
and U980 (N_980,In_1309,In_1277);
xor U981 (N_981,N_701,N_572);
or U982 (N_982,N_820,N_286);
nor U983 (N_983,N_815,N_55);
nand U984 (N_984,In_224,In_1278);
or U985 (N_985,N_579,N_748);
and U986 (N_986,N_847,N_788);
or U987 (N_987,N_611,N_883);
and U988 (N_988,N_791,N_498);
and U989 (N_989,N_661,In_1161);
or U990 (N_990,In_473,N_850);
nand U991 (N_991,N_766,N_886);
xor U992 (N_992,N_370,N_685);
xor U993 (N_993,N_573,N_203);
and U994 (N_994,N_887,N_874);
nor U995 (N_995,N_606,N_857);
nand U996 (N_996,N_667,N_167);
nand U997 (N_997,N_879,N_664);
and U998 (N_998,N_771,In_509);
nand U999 (N_999,In_1214,N_366);
and U1000 (N_1000,In_214,N_493);
and U1001 (N_1001,N_827,N_714);
nand U1002 (N_1002,N_826,In_386);
xor U1003 (N_1003,N_462,N_773);
nor U1004 (N_1004,N_722,N_880);
xnor U1005 (N_1005,N_620,N_663);
xnor U1006 (N_1006,N_823,N_633);
nand U1007 (N_1007,N_692,N_385);
nand U1008 (N_1008,N_675,N_170);
or U1009 (N_1009,N_374,N_317);
and U1010 (N_1010,N_158,N_645);
nor U1011 (N_1011,N_475,N_418);
or U1012 (N_1012,In_485,N_706);
xnor U1013 (N_1013,N_660,In_694);
nand U1014 (N_1014,N_420,In_1020);
or U1015 (N_1015,N_578,N_360);
and U1016 (N_1016,N_615,N_549);
nand U1017 (N_1017,In_925,In_1141);
and U1018 (N_1018,N_607,N_476);
or U1019 (N_1019,N_544,N_785);
xnor U1020 (N_1020,N_678,N_586);
and U1021 (N_1021,N_376,N_237);
xnor U1022 (N_1022,In_1354,N_736);
nand U1023 (N_1023,N_713,In_399);
or U1024 (N_1024,N_285,N_764);
xnor U1025 (N_1025,N_802,N_641);
or U1026 (N_1026,In_1078,N_556);
xor U1027 (N_1027,N_345,In_695);
nand U1028 (N_1028,In_809,N_627);
or U1029 (N_1029,N_892,N_715);
and U1030 (N_1030,N_752,N_566);
nand U1031 (N_1031,N_501,N_622);
or U1032 (N_1032,In_888,N_478);
nor U1033 (N_1033,In_461,In_383);
xnor U1034 (N_1034,N_858,In_939);
xnor U1035 (N_1035,N_542,N_737);
nor U1036 (N_1036,In_356,In_805);
nand U1037 (N_1037,N_778,N_800);
and U1038 (N_1038,N_770,In_36);
or U1039 (N_1039,N_655,N_132);
or U1040 (N_1040,In_729,N_725);
xnor U1041 (N_1041,N_818,N_571);
xnor U1042 (N_1042,N_761,N_658);
nor U1043 (N_1043,N_517,In_923);
xor U1044 (N_1044,N_650,N_759);
xor U1045 (N_1045,N_790,N_502);
nand U1046 (N_1046,N_603,N_784);
nor U1047 (N_1047,N_659,N_504);
or U1048 (N_1048,In_686,N_355);
xnor U1049 (N_1049,N_787,N_871);
xnor U1050 (N_1050,N_775,In_25);
nand U1051 (N_1051,N_700,N_819);
and U1052 (N_1052,In_742,In_90);
nand U1053 (N_1053,N_270,N_801);
and U1054 (N_1054,N_896,N_711);
nor U1055 (N_1055,In_517,N_665);
nand U1056 (N_1056,N_14,N_846);
and U1057 (N_1057,N_402,N_580);
or U1058 (N_1058,N_101,N_704);
or U1059 (N_1059,N_590,N_812);
nor U1060 (N_1060,N_239,N_173);
nor U1061 (N_1061,In_1405,N_367);
nand U1062 (N_1062,In_1044,In_1006);
or U1063 (N_1063,N_710,N_848);
xor U1064 (N_1064,N_838,N_523);
nand U1065 (N_1065,N_666,N_399);
nor U1066 (N_1066,In_1030,In_453);
or U1067 (N_1067,N_832,N_530);
nor U1068 (N_1068,N_637,N_513);
and U1069 (N_1069,N_509,In_942);
or U1070 (N_1070,In_675,N_866);
or U1071 (N_1071,In_638,In_131);
and U1072 (N_1072,N_632,N_636);
nor U1073 (N_1073,N_696,N_814);
nor U1074 (N_1074,N_762,N_565);
and U1075 (N_1075,N_756,N_876);
xor U1076 (N_1076,N_702,N_207);
nand U1077 (N_1077,N_842,N_653);
nand U1078 (N_1078,N_739,N_646);
nor U1079 (N_1079,In_603,N_624);
xor U1080 (N_1080,In_18,In_434);
and U1081 (N_1081,In_267,N_488);
or U1082 (N_1082,N_381,N_156);
and U1083 (N_1083,N_431,N_188);
xnor U1084 (N_1084,N_231,In_647);
nor U1085 (N_1085,N_185,In_1231);
nand U1086 (N_1086,In_477,In_892);
xor U1087 (N_1087,N_864,In_250);
nor U1088 (N_1088,In_1296,N_765);
xor U1089 (N_1089,In_1192,In_1351);
xnor U1090 (N_1090,In_152,N_411);
nand U1091 (N_1091,In_1372,N_780);
xnor U1092 (N_1092,N_776,N_450);
and U1093 (N_1093,In_1000,N_878);
xnor U1094 (N_1094,N_869,N_889);
nor U1095 (N_1095,N_439,N_673);
or U1096 (N_1096,N_849,N_250);
and U1097 (N_1097,N_442,N_885);
or U1098 (N_1098,In_956,N_640);
nand U1099 (N_1099,In_1062,N_831);
nor U1100 (N_1100,N_811,N_440);
nor U1101 (N_1101,In_278,In_763);
and U1102 (N_1102,In_1321,N_555);
nand U1103 (N_1103,In_1199,N_730);
nor U1104 (N_1104,In_1213,N_694);
nand U1105 (N_1105,In_283,N_859);
and U1106 (N_1106,In_411,N_570);
nor U1107 (N_1107,N_877,In_1298);
and U1108 (N_1108,N_768,N_860);
xor U1109 (N_1109,N_356,N_708);
xnor U1110 (N_1110,N_822,N_432);
and U1111 (N_1111,N_881,N_47);
nor U1112 (N_1112,N_772,In_1140);
and U1113 (N_1113,N_797,N_732);
nor U1114 (N_1114,N_738,N_344);
nand U1115 (N_1115,N_616,N_804);
and U1116 (N_1116,N_405,N_720);
or U1117 (N_1117,N_508,N_845);
or U1118 (N_1118,N_521,N_895);
xnor U1119 (N_1119,In_754,In_1499);
or U1120 (N_1120,In_857,N_652);
xnor U1121 (N_1121,N_840,N_601);
xnor U1122 (N_1122,N_789,N_662);
xor U1123 (N_1123,N_854,In_643);
nor U1124 (N_1124,N_716,N_78);
nor U1125 (N_1125,N_888,In_1220);
or U1126 (N_1126,N_740,In_903);
and U1127 (N_1127,N_351,In_1001);
or U1128 (N_1128,In_258,N_833);
xor U1129 (N_1129,N_516,N_872);
and U1130 (N_1130,N_774,N_683);
or U1131 (N_1131,N_75,N_255);
and U1132 (N_1132,N_434,N_474);
xnor U1133 (N_1133,N_807,N_817);
and U1134 (N_1134,N_793,In_1126);
or U1135 (N_1135,In_120,N_862);
nor U1136 (N_1136,N_836,N_853);
and U1137 (N_1137,N_534,N_682);
and U1138 (N_1138,N_698,N_596);
or U1139 (N_1139,N_657,N_500);
and U1140 (N_1140,In_1280,N_72);
nand U1141 (N_1141,N_795,N_783);
nor U1142 (N_1142,In_493,In_462);
xnor U1143 (N_1143,N_614,N_753);
nand U1144 (N_1144,N_856,N_562);
or U1145 (N_1145,N_691,N_769);
nand U1146 (N_1146,N_816,N_705);
nand U1147 (N_1147,N_767,N_643);
or U1148 (N_1148,N_760,N_409);
nand U1149 (N_1149,N_805,In_598);
nor U1150 (N_1150,N_609,N_23);
nor U1151 (N_1151,N_779,N_882);
nand U1152 (N_1152,N_457,In_1425);
nor U1153 (N_1153,N_726,N_639);
nor U1154 (N_1154,N_452,N_593);
or U1155 (N_1155,In_446,N_605);
and U1156 (N_1156,N_600,In_1399);
nor U1157 (N_1157,In_147,N_511);
nand U1158 (N_1158,In_1453,N_531);
xnor U1159 (N_1159,N_863,N_401);
nand U1160 (N_1160,N_618,N_798);
or U1161 (N_1161,N_745,N_649);
xor U1162 (N_1162,N_865,N_631);
nor U1163 (N_1163,N_46,N_430);
nand U1164 (N_1164,N_821,N_613);
nor U1165 (N_1165,In_1456,In_781);
xnor U1166 (N_1166,In_235,N_217);
nand U1167 (N_1167,N_867,N_625);
and U1168 (N_1168,N_751,N_809);
and U1169 (N_1169,N_731,In_1054);
and U1170 (N_1170,In_59,In_768);
or U1171 (N_1171,N_735,In_870);
or U1172 (N_1172,In_2,N_828);
xnor U1173 (N_1173,N_635,N_604);
nand U1174 (N_1174,N_813,N_792);
xor U1175 (N_1175,N_416,N_4);
or U1176 (N_1176,N_125,In_177);
or U1177 (N_1177,N_808,N_707);
nand U1178 (N_1178,N_855,N_825);
xnor U1179 (N_1179,In_588,N_712);
nor U1180 (N_1180,N_152,N_781);
nor U1181 (N_1181,N_742,In_1311);
nor U1182 (N_1182,In_67,N_574);
nand U1183 (N_1183,N_672,N_276);
nor U1184 (N_1184,N_835,N_196);
and U1185 (N_1185,In_800,N_458);
and U1186 (N_1186,N_898,N_610);
nor U1187 (N_1187,N_599,N_290);
nand U1188 (N_1188,In_1319,N_602);
or U1189 (N_1189,In_880,N_750);
nand U1190 (N_1190,In_1193,N_754);
or U1191 (N_1191,N_677,In_560);
or U1192 (N_1192,In_827,In_856);
nor U1193 (N_1193,N_1,N_384);
nor U1194 (N_1194,N_717,In_569);
or U1195 (N_1195,In_402,N_719);
or U1196 (N_1196,N_626,In_876);
and U1197 (N_1197,N_728,N_744);
nand U1198 (N_1198,N_612,In_328);
nand U1199 (N_1199,In_1069,In_672);
xor U1200 (N_1200,N_1070,N_1189);
nor U1201 (N_1201,N_1133,N_948);
nor U1202 (N_1202,N_917,N_1105);
nand U1203 (N_1203,N_924,N_1066);
nand U1204 (N_1204,N_1030,N_1161);
and U1205 (N_1205,N_929,N_921);
xnor U1206 (N_1206,N_1198,N_1121);
nor U1207 (N_1207,N_1104,N_1165);
nand U1208 (N_1208,N_930,N_1028);
and U1209 (N_1209,N_1085,N_1180);
nand U1210 (N_1210,N_1178,N_1118);
or U1211 (N_1211,N_1064,N_975);
nand U1212 (N_1212,N_1050,N_1142);
xor U1213 (N_1213,N_943,N_963);
and U1214 (N_1214,N_904,N_1128);
and U1215 (N_1215,N_1182,N_1194);
nor U1216 (N_1216,N_1075,N_1083);
nand U1217 (N_1217,N_1008,N_1037);
nor U1218 (N_1218,N_1143,N_1041);
or U1219 (N_1219,N_1038,N_964);
and U1220 (N_1220,N_906,N_1016);
xnor U1221 (N_1221,N_919,N_956);
or U1222 (N_1222,N_931,N_1036);
nand U1223 (N_1223,N_998,N_969);
or U1224 (N_1224,N_1102,N_997);
and U1225 (N_1225,N_979,N_984);
nor U1226 (N_1226,N_950,N_1170);
nor U1227 (N_1227,N_970,N_900);
nand U1228 (N_1228,N_1126,N_937);
xnor U1229 (N_1229,N_1112,N_1011);
or U1230 (N_1230,N_905,N_934);
nand U1231 (N_1231,N_974,N_1120);
or U1232 (N_1232,N_1012,N_1000);
or U1233 (N_1233,N_1057,N_1084);
nand U1234 (N_1234,N_1032,N_922);
nand U1235 (N_1235,N_1029,N_1122);
and U1236 (N_1236,N_911,N_1002);
and U1237 (N_1237,N_968,N_1107);
or U1238 (N_1238,N_1138,N_1145);
xor U1239 (N_1239,N_923,N_967);
xnor U1240 (N_1240,N_1049,N_939);
and U1241 (N_1241,N_992,N_962);
nand U1242 (N_1242,N_1046,N_1086);
nor U1243 (N_1243,N_1119,N_1051);
and U1244 (N_1244,N_910,N_1190);
or U1245 (N_1245,N_972,N_1171);
or U1246 (N_1246,N_1110,N_980);
nor U1247 (N_1247,N_996,N_1168);
xor U1248 (N_1248,N_936,N_1080);
or U1249 (N_1249,N_1092,N_1155);
nor U1250 (N_1250,N_1054,N_1106);
and U1251 (N_1251,N_1131,N_1117);
nand U1252 (N_1252,N_1088,N_1072);
nand U1253 (N_1253,N_1079,N_1132);
xnor U1254 (N_1254,N_1010,N_1044);
nor U1255 (N_1255,N_920,N_987);
xnor U1256 (N_1256,N_989,N_927);
nor U1257 (N_1257,N_1174,N_1159);
nand U1258 (N_1258,N_933,N_1141);
nor U1259 (N_1259,N_1087,N_1153);
nor U1260 (N_1260,N_1006,N_977);
xor U1261 (N_1261,N_990,N_1071);
nor U1262 (N_1262,N_1172,N_1196);
or U1263 (N_1263,N_1045,N_1160);
xnor U1264 (N_1264,N_1179,N_916);
nand U1265 (N_1265,N_1069,N_1094);
and U1266 (N_1266,N_909,N_1108);
nand U1267 (N_1267,N_1139,N_1033);
or U1268 (N_1268,N_951,N_1111);
nand U1269 (N_1269,N_1093,N_1146);
nor U1270 (N_1270,N_1137,N_935);
nand U1271 (N_1271,N_1048,N_952);
and U1272 (N_1272,N_957,N_1040);
nand U1273 (N_1273,N_1101,N_1115);
nand U1274 (N_1274,N_1167,N_1007);
or U1275 (N_1275,N_1024,N_1082);
and U1276 (N_1276,N_1148,N_1157);
nand U1277 (N_1277,N_949,N_994);
or U1278 (N_1278,N_1127,N_1125);
nor U1279 (N_1279,N_1150,N_1154);
nor U1280 (N_1280,N_1026,N_1097);
and U1281 (N_1281,N_1060,N_941);
nor U1282 (N_1282,N_901,N_1067);
nand U1283 (N_1283,N_1192,N_1034);
or U1284 (N_1284,N_1164,N_1039);
xnor U1285 (N_1285,N_1001,N_1042);
and U1286 (N_1286,N_961,N_1129);
nor U1287 (N_1287,N_946,N_1077);
nand U1288 (N_1288,N_926,N_958);
nor U1289 (N_1289,N_1052,N_1199);
or U1290 (N_1290,N_912,N_913);
nor U1291 (N_1291,N_1185,N_1173);
and U1292 (N_1292,N_1081,N_1158);
nor U1293 (N_1293,N_1156,N_1162);
nor U1294 (N_1294,N_985,N_940);
and U1295 (N_1295,N_1193,N_1035);
nand U1296 (N_1296,N_1056,N_944);
and U1297 (N_1297,N_1135,N_1022);
nand U1298 (N_1298,N_1191,N_971);
or U1299 (N_1299,N_1136,N_965);
xnor U1300 (N_1300,N_1096,N_1188);
nand U1301 (N_1301,N_902,N_955);
nand U1302 (N_1302,N_976,N_1103);
and U1303 (N_1303,N_1005,N_1065);
or U1304 (N_1304,N_1149,N_1187);
xnor U1305 (N_1305,N_959,N_1058);
xor U1306 (N_1306,N_938,N_982);
and U1307 (N_1307,N_1151,N_1099);
nor U1308 (N_1308,N_1144,N_918);
or U1309 (N_1309,N_1177,N_1014);
nand U1310 (N_1310,N_1089,N_908);
and U1311 (N_1311,N_1023,N_1100);
nand U1312 (N_1312,N_1095,N_1123);
nor U1313 (N_1313,N_1140,N_1166);
nor U1314 (N_1314,N_960,N_1090);
and U1315 (N_1315,N_999,N_1134);
xor U1316 (N_1316,N_1078,N_1109);
or U1317 (N_1317,N_914,N_988);
or U1318 (N_1318,N_991,N_1004);
nand U1319 (N_1319,N_1113,N_1147);
nor U1320 (N_1320,N_1184,N_953);
xnor U1321 (N_1321,N_986,N_1183);
nand U1322 (N_1322,N_1116,N_1098);
or U1323 (N_1323,N_1061,N_1009);
xor U1324 (N_1324,N_1031,N_1013);
nor U1325 (N_1325,N_915,N_1027);
nor U1326 (N_1326,N_966,N_1186);
nand U1327 (N_1327,N_1074,N_1176);
nor U1328 (N_1328,N_1130,N_1076);
nor U1329 (N_1329,N_1152,N_945);
nor U1330 (N_1330,N_1025,N_981);
nor U1331 (N_1331,N_1021,N_1169);
and U1332 (N_1332,N_1114,N_1197);
and U1333 (N_1333,N_1175,N_1091);
or U1334 (N_1334,N_925,N_1059);
and U1335 (N_1335,N_932,N_1068);
nor U1336 (N_1336,N_973,N_928);
nor U1337 (N_1337,N_978,N_1015);
or U1338 (N_1338,N_1003,N_1073);
or U1339 (N_1339,N_1063,N_993);
nand U1340 (N_1340,N_1055,N_1017);
or U1341 (N_1341,N_1047,N_1062);
xor U1342 (N_1342,N_903,N_1195);
xor U1343 (N_1343,N_1043,N_942);
and U1344 (N_1344,N_947,N_1163);
xnor U1345 (N_1345,N_1018,N_1019);
and U1346 (N_1346,N_954,N_1181);
and U1347 (N_1347,N_995,N_1053);
or U1348 (N_1348,N_983,N_1124);
nand U1349 (N_1349,N_907,N_1020);
or U1350 (N_1350,N_1103,N_1162);
nor U1351 (N_1351,N_1144,N_1142);
nor U1352 (N_1352,N_1004,N_1099);
and U1353 (N_1353,N_910,N_1119);
nor U1354 (N_1354,N_1156,N_1164);
nor U1355 (N_1355,N_1016,N_1199);
and U1356 (N_1356,N_972,N_1084);
or U1357 (N_1357,N_1157,N_974);
and U1358 (N_1358,N_1101,N_957);
nor U1359 (N_1359,N_1178,N_1010);
or U1360 (N_1360,N_1188,N_981);
xnor U1361 (N_1361,N_976,N_1052);
nand U1362 (N_1362,N_1171,N_928);
nand U1363 (N_1363,N_947,N_1079);
and U1364 (N_1364,N_946,N_934);
nand U1365 (N_1365,N_1160,N_1161);
xnor U1366 (N_1366,N_1087,N_1161);
nor U1367 (N_1367,N_1054,N_993);
nor U1368 (N_1368,N_954,N_1077);
nor U1369 (N_1369,N_1123,N_1134);
nand U1370 (N_1370,N_1028,N_980);
nor U1371 (N_1371,N_1188,N_1010);
xor U1372 (N_1372,N_993,N_1141);
nor U1373 (N_1373,N_947,N_1039);
nand U1374 (N_1374,N_1021,N_919);
or U1375 (N_1375,N_1101,N_1112);
and U1376 (N_1376,N_970,N_990);
xor U1377 (N_1377,N_999,N_1139);
nor U1378 (N_1378,N_920,N_1167);
nor U1379 (N_1379,N_1056,N_1106);
xor U1380 (N_1380,N_1154,N_981);
or U1381 (N_1381,N_1030,N_964);
or U1382 (N_1382,N_1123,N_945);
or U1383 (N_1383,N_1084,N_1030);
xnor U1384 (N_1384,N_1054,N_915);
or U1385 (N_1385,N_1197,N_1075);
nor U1386 (N_1386,N_957,N_1056);
and U1387 (N_1387,N_1012,N_1002);
nand U1388 (N_1388,N_1139,N_984);
nor U1389 (N_1389,N_1124,N_1166);
or U1390 (N_1390,N_954,N_968);
nand U1391 (N_1391,N_1022,N_1004);
xor U1392 (N_1392,N_1136,N_1197);
nor U1393 (N_1393,N_1137,N_1021);
or U1394 (N_1394,N_1010,N_1088);
xnor U1395 (N_1395,N_1036,N_999);
or U1396 (N_1396,N_1014,N_1099);
nor U1397 (N_1397,N_964,N_1056);
or U1398 (N_1398,N_1132,N_1047);
nor U1399 (N_1399,N_1190,N_1175);
nor U1400 (N_1400,N_1185,N_1068);
nor U1401 (N_1401,N_936,N_1010);
nand U1402 (N_1402,N_1168,N_1164);
nor U1403 (N_1403,N_1195,N_1138);
nand U1404 (N_1404,N_926,N_1156);
xnor U1405 (N_1405,N_902,N_971);
or U1406 (N_1406,N_1189,N_1006);
or U1407 (N_1407,N_941,N_1051);
xnor U1408 (N_1408,N_1119,N_1175);
xor U1409 (N_1409,N_1171,N_1094);
xor U1410 (N_1410,N_1056,N_916);
or U1411 (N_1411,N_984,N_972);
or U1412 (N_1412,N_935,N_1066);
xor U1413 (N_1413,N_1078,N_969);
xnor U1414 (N_1414,N_1068,N_1010);
and U1415 (N_1415,N_1018,N_975);
nor U1416 (N_1416,N_1087,N_1028);
nand U1417 (N_1417,N_1006,N_988);
and U1418 (N_1418,N_995,N_1132);
nand U1419 (N_1419,N_942,N_940);
xor U1420 (N_1420,N_904,N_1185);
nand U1421 (N_1421,N_988,N_1100);
or U1422 (N_1422,N_1040,N_1000);
or U1423 (N_1423,N_1170,N_1153);
nand U1424 (N_1424,N_1071,N_1087);
nand U1425 (N_1425,N_956,N_1046);
and U1426 (N_1426,N_1170,N_1159);
nor U1427 (N_1427,N_1088,N_1161);
xor U1428 (N_1428,N_1046,N_943);
nor U1429 (N_1429,N_1179,N_1108);
nand U1430 (N_1430,N_910,N_973);
nand U1431 (N_1431,N_946,N_1042);
and U1432 (N_1432,N_900,N_1048);
xnor U1433 (N_1433,N_910,N_1115);
or U1434 (N_1434,N_952,N_1101);
nor U1435 (N_1435,N_998,N_1047);
and U1436 (N_1436,N_980,N_998);
nand U1437 (N_1437,N_1127,N_1138);
xor U1438 (N_1438,N_967,N_1174);
and U1439 (N_1439,N_1181,N_1121);
or U1440 (N_1440,N_1099,N_924);
nor U1441 (N_1441,N_1147,N_1157);
nand U1442 (N_1442,N_1014,N_1180);
nor U1443 (N_1443,N_932,N_1015);
xor U1444 (N_1444,N_939,N_1028);
nand U1445 (N_1445,N_1007,N_1135);
or U1446 (N_1446,N_1149,N_1102);
nor U1447 (N_1447,N_967,N_1171);
xor U1448 (N_1448,N_934,N_970);
or U1449 (N_1449,N_998,N_1134);
nand U1450 (N_1450,N_971,N_962);
nand U1451 (N_1451,N_908,N_979);
or U1452 (N_1452,N_1193,N_1118);
and U1453 (N_1453,N_1132,N_1008);
nand U1454 (N_1454,N_1080,N_1082);
nand U1455 (N_1455,N_986,N_918);
nand U1456 (N_1456,N_903,N_1102);
nand U1457 (N_1457,N_1011,N_978);
nand U1458 (N_1458,N_934,N_1164);
or U1459 (N_1459,N_1061,N_1028);
or U1460 (N_1460,N_1168,N_1192);
or U1461 (N_1461,N_1173,N_1114);
or U1462 (N_1462,N_1190,N_973);
and U1463 (N_1463,N_1075,N_997);
and U1464 (N_1464,N_1091,N_1080);
xor U1465 (N_1465,N_1118,N_1130);
and U1466 (N_1466,N_1093,N_1046);
nor U1467 (N_1467,N_1021,N_1129);
nor U1468 (N_1468,N_1006,N_1140);
or U1469 (N_1469,N_979,N_974);
nand U1470 (N_1470,N_1056,N_900);
xnor U1471 (N_1471,N_1075,N_965);
and U1472 (N_1472,N_1082,N_1050);
nand U1473 (N_1473,N_1038,N_1069);
or U1474 (N_1474,N_979,N_960);
xnor U1475 (N_1475,N_1197,N_973);
nand U1476 (N_1476,N_1097,N_1130);
xnor U1477 (N_1477,N_1014,N_909);
or U1478 (N_1478,N_1048,N_1105);
nor U1479 (N_1479,N_958,N_1046);
xnor U1480 (N_1480,N_1125,N_1065);
nor U1481 (N_1481,N_1045,N_903);
xor U1482 (N_1482,N_1074,N_993);
nand U1483 (N_1483,N_1008,N_951);
or U1484 (N_1484,N_1091,N_1067);
nand U1485 (N_1485,N_1181,N_974);
and U1486 (N_1486,N_951,N_959);
xor U1487 (N_1487,N_1189,N_968);
nand U1488 (N_1488,N_1194,N_1012);
nor U1489 (N_1489,N_977,N_926);
and U1490 (N_1490,N_956,N_900);
nand U1491 (N_1491,N_1004,N_1090);
nand U1492 (N_1492,N_1026,N_1019);
nand U1493 (N_1493,N_1118,N_1006);
and U1494 (N_1494,N_978,N_967);
xor U1495 (N_1495,N_932,N_919);
xnor U1496 (N_1496,N_910,N_1173);
xor U1497 (N_1497,N_980,N_957);
and U1498 (N_1498,N_1075,N_1045);
nand U1499 (N_1499,N_963,N_1142);
and U1500 (N_1500,N_1216,N_1485);
nor U1501 (N_1501,N_1231,N_1475);
nand U1502 (N_1502,N_1337,N_1480);
xor U1503 (N_1503,N_1420,N_1398);
and U1504 (N_1504,N_1328,N_1213);
nor U1505 (N_1505,N_1302,N_1408);
and U1506 (N_1506,N_1498,N_1397);
nor U1507 (N_1507,N_1319,N_1441);
or U1508 (N_1508,N_1399,N_1376);
nand U1509 (N_1509,N_1276,N_1320);
xor U1510 (N_1510,N_1315,N_1332);
nand U1511 (N_1511,N_1338,N_1347);
and U1512 (N_1512,N_1422,N_1241);
or U1513 (N_1513,N_1250,N_1203);
nand U1514 (N_1514,N_1427,N_1488);
nor U1515 (N_1515,N_1421,N_1344);
nand U1516 (N_1516,N_1416,N_1371);
and U1517 (N_1517,N_1339,N_1379);
xor U1518 (N_1518,N_1278,N_1452);
nor U1519 (N_1519,N_1403,N_1303);
nand U1520 (N_1520,N_1340,N_1405);
xor U1521 (N_1521,N_1275,N_1486);
nand U1522 (N_1522,N_1410,N_1277);
or U1523 (N_1523,N_1419,N_1336);
nor U1524 (N_1524,N_1472,N_1459);
nor U1525 (N_1525,N_1362,N_1295);
xor U1526 (N_1526,N_1221,N_1451);
nand U1527 (N_1527,N_1254,N_1449);
nor U1528 (N_1528,N_1429,N_1274);
and U1529 (N_1529,N_1366,N_1359);
and U1530 (N_1530,N_1424,N_1490);
and U1531 (N_1531,N_1463,N_1365);
or U1532 (N_1532,N_1270,N_1477);
nor U1533 (N_1533,N_1330,N_1375);
nand U1534 (N_1534,N_1245,N_1364);
xnor U1535 (N_1535,N_1207,N_1282);
or U1536 (N_1536,N_1411,N_1391);
xnor U1537 (N_1537,N_1209,N_1307);
xnor U1538 (N_1538,N_1395,N_1466);
nand U1539 (N_1539,N_1292,N_1322);
and U1540 (N_1540,N_1235,N_1311);
or U1541 (N_1541,N_1210,N_1478);
nand U1542 (N_1542,N_1447,N_1226);
or U1543 (N_1543,N_1329,N_1325);
xor U1544 (N_1544,N_1438,N_1385);
xnor U1545 (N_1545,N_1426,N_1247);
xor U1546 (N_1546,N_1423,N_1285);
nand U1547 (N_1547,N_1239,N_1223);
or U1548 (N_1548,N_1234,N_1263);
or U1549 (N_1549,N_1308,N_1389);
nand U1550 (N_1550,N_1269,N_1467);
nand U1551 (N_1551,N_1412,N_1439);
xor U1552 (N_1552,N_1491,N_1446);
or U1553 (N_1553,N_1479,N_1266);
and U1554 (N_1554,N_1313,N_1256);
nand U1555 (N_1555,N_1394,N_1448);
xnor U1556 (N_1556,N_1415,N_1383);
nor U1557 (N_1557,N_1215,N_1255);
nor U1558 (N_1558,N_1346,N_1357);
and U1559 (N_1559,N_1233,N_1378);
nor U1560 (N_1560,N_1392,N_1253);
nor U1561 (N_1561,N_1211,N_1280);
nand U1562 (N_1562,N_1377,N_1374);
and U1563 (N_1563,N_1342,N_1281);
or U1564 (N_1564,N_1462,N_1200);
nand U1565 (N_1565,N_1458,N_1252);
nor U1566 (N_1566,N_1373,N_1316);
or U1567 (N_1567,N_1323,N_1413);
or U1568 (N_1568,N_1229,N_1492);
or U1569 (N_1569,N_1249,N_1232);
and U1570 (N_1570,N_1341,N_1361);
and U1571 (N_1571,N_1219,N_1387);
xor U1572 (N_1572,N_1318,N_1432);
or U1573 (N_1573,N_1294,N_1440);
or U1574 (N_1574,N_1264,N_1312);
xor U1575 (N_1575,N_1246,N_1431);
or U1576 (N_1576,N_1487,N_1224);
or U1577 (N_1577,N_1314,N_1272);
or U1578 (N_1578,N_1493,N_1434);
nor U1579 (N_1579,N_1442,N_1222);
or U1580 (N_1580,N_1414,N_1251);
nand U1581 (N_1581,N_1331,N_1217);
xnor U1582 (N_1582,N_1388,N_1236);
nor U1583 (N_1583,N_1297,N_1349);
nor U1584 (N_1584,N_1353,N_1237);
or U1585 (N_1585,N_1382,N_1481);
or U1586 (N_1586,N_1304,N_1474);
nor U1587 (N_1587,N_1284,N_1406);
nor U1588 (N_1588,N_1453,N_1370);
xor U1589 (N_1589,N_1321,N_1317);
nand U1590 (N_1590,N_1228,N_1372);
nand U1591 (N_1591,N_1286,N_1380);
nor U1592 (N_1592,N_1358,N_1214);
or U1593 (N_1593,N_1267,N_1227);
nand U1594 (N_1594,N_1218,N_1205);
xor U1595 (N_1595,N_1469,N_1268);
and U1596 (N_1596,N_1265,N_1326);
and U1597 (N_1597,N_1202,N_1327);
and U1598 (N_1598,N_1367,N_1273);
nor U1599 (N_1599,N_1455,N_1204);
nor U1600 (N_1600,N_1283,N_1417);
and U1601 (N_1601,N_1407,N_1243);
and U1602 (N_1602,N_1220,N_1296);
nor U1603 (N_1603,N_1454,N_1260);
nor U1604 (N_1604,N_1261,N_1354);
nor U1605 (N_1605,N_1460,N_1428);
nand U1606 (N_1606,N_1445,N_1206);
xor U1607 (N_1607,N_1298,N_1465);
nand U1608 (N_1608,N_1400,N_1360);
nor U1609 (N_1609,N_1238,N_1259);
and U1610 (N_1610,N_1457,N_1348);
nand U1611 (N_1611,N_1476,N_1293);
nand U1612 (N_1612,N_1262,N_1433);
nor U1613 (N_1613,N_1212,N_1456);
and U1614 (N_1614,N_1271,N_1495);
xor U1615 (N_1615,N_1242,N_1436);
or U1616 (N_1616,N_1381,N_1343);
xor U1617 (N_1617,N_1402,N_1418);
nand U1618 (N_1618,N_1345,N_1497);
or U1619 (N_1619,N_1287,N_1390);
and U1620 (N_1620,N_1494,N_1496);
and U1621 (N_1621,N_1450,N_1468);
or U1622 (N_1622,N_1333,N_1471);
or U1623 (N_1623,N_1310,N_1355);
and U1624 (N_1624,N_1386,N_1352);
or U1625 (N_1625,N_1305,N_1437);
xnor U1626 (N_1626,N_1461,N_1301);
nand U1627 (N_1627,N_1257,N_1289);
and U1628 (N_1628,N_1290,N_1473);
nand U1629 (N_1629,N_1484,N_1334);
and U1630 (N_1630,N_1368,N_1288);
nor U1631 (N_1631,N_1291,N_1409);
and U1632 (N_1632,N_1201,N_1444);
and U1633 (N_1633,N_1363,N_1324);
and U1634 (N_1634,N_1404,N_1299);
nand U1635 (N_1635,N_1384,N_1350);
nor U1636 (N_1636,N_1309,N_1393);
xnor U1637 (N_1637,N_1335,N_1401);
and U1638 (N_1638,N_1230,N_1435);
or U1639 (N_1639,N_1225,N_1489);
or U1640 (N_1640,N_1425,N_1240);
nand U1641 (N_1641,N_1356,N_1279);
nor U1642 (N_1642,N_1369,N_1464);
nor U1643 (N_1643,N_1248,N_1470);
or U1644 (N_1644,N_1244,N_1208);
or U1645 (N_1645,N_1300,N_1396);
nor U1646 (N_1646,N_1443,N_1258);
nand U1647 (N_1647,N_1306,N_1482);
xnor U1648 (N_1648,N_1430,N_1351);
nor U1649 (N_1649,N_1483,N_1499);
nor U1650 (N_1650,N_1414,N_1316);
nor U1651 (N_1651,N_1312,N_1338);
nand U1652 (N_1652,N_1487,N_1486);
xor U1653 (N_1653,N_1433,N_1314);
nor U1654 (N_1654,N_1358,N_1226);
or U1655 (N_1655,N_1489,N_1223);
nor U1656 (N_1656,N_1327,N_1278);
or U1657 (N_1657,N_1210,N_1334);
nor U1658 (N_1658,N_1320,N_1455);
xor U1659 (N_1659,N_1369,N_1411);
nand U1660 (N_1660,N_1359,N_1285);
nor U1661 (N_1661,N_1238,N_1353);
nor U1662 (N_1662,N_1241,N_1249);
or U1663 (N_1663,N_1489,N_1414);
xnor U1664 (N_1664,N_1225,N_1459);
nor U1665 (N_1665,N_1281,N_1456);
xor U1666 (N_1666,N_1458,N_1301);
or U1667 (N_1667,N_1383,N_1258);
nand U1668 (N_1668,N_1432,N_1481);
and U1669 (N_1669,N_1213,N_1301);
nand U1670 (N_1670,N_1324,N_1264);
xnor U1671 (N_1671,N_1397,N_1218);
nand U1672 (N_1672,N_1274,N_1238);
nor U1673 (N_1673,N_1481,N_1423);
or U1674 (N_1674,N_1481,N_1375);
xnor U1675 (N_1675,N_1273,N_1489);
xnor U1676 (N_1676,N_1296,N_1403);
or U1677 (N_1677,N_1231,N_1382);
xor U1678 (N_1678,N_1410,N_1218);
nor U1679 (N_1679,N_1255,N_1334);
and U1680 (N_1680,N_1436,N_1415);
xor U1681 (N_1681,N_1336,N_1306);
xor U1682 (N_1682,N_1447,N_1438);
nor U1683 (N_1683,N_1413,N_1328);
nand U1684 (N_1684,N_1212,N_1352);
and U1685 (N_1685,N_1229,N_1411);
and U1686 (N_1686,N_1459,N_1201);
xor U1687 (N_1687,N_1279,N_1236);
or U1688 (N_1688,N_1222,N_1258);
nor U1689 (N_1689,N_1320,N_1465);
or U1690 (N_1690,N_1359,N_1419);
nor U1691 (N_1691,N_1208,N_1200);
nor U1692 (N_1692,N_1333,N_1462);
nor U1693 (N_1693,N_1329,N_1399);
or U1694 (N_1694,N_1407,N_1406);
nor U1695 (N_1695,N_1256,N_1235);
nor U1696 (N_1696,N_1353,N_1386);
or U1697 (N_1697,N_1339,N_1220);
nand U1698 (N_1698,N_1467,N_1435);
xnor U1699 (N_1699,N_1427,N_1286);
and U1700 (N_1700,N_1282,N_1353);
nor U1701 (N_1701,N_1401,N_1362);
nand U1702 (N_1702,N_1373,N_1448);
and U1703 (N_1703,N_1333,N_1494);
and U1704 (N_1704,N_1457,N_1398);
and U1705 (N_1705,N_1418,N_1409);
xor U1706 (N_1706,N_1230,N_1432);
and U1707 (N_1707,N_1286,N_1313);
or U1708 (N_1708,N_1234,N_1498);
or U1709 (N_1709,N_1371,N_1477);
and U1710 (N_1710,N_1378,N_1200);
xnor U1711 (N_1711,N_1486,N_1220);
xnor U1712 (N_1712,N_1453,N_1316);
or U1713 (N_1713,N_1358,N_1494);
or U1714 (N_1714,N_1424,N_1406);
or U1715 (N_1715,N_1429,N_1307);
nand U1716 (N_1716,N_1474,N_1230);
xor U1717 (N_1717,N_1434,N_1421);
and U1718 (N_1718,N_1270,N_1273);
or U1719 (N_1719,N_1259,N_1336);
xnor U1720 (N_1720,N_1451,N_1431);
nand U1721 (N_1721,N_1448,N_1344);
and U1722 (N_1722,N_1373,N_1485);
nor U1723 (N_1723,N_1209,N_1475);
and U1724 (N_1724,N_1291,N_1292);
or U1725 (N_1725,N_1491,N_1256);
xor U1726 (N_1726,N_1406,N_1405);
nor U1727 (N_1727,N_1463,N_1383);
or U1728 (N_1728,N_1347,N_1346);
or U1729 (N_1729,N_1349,N_1435);
nor U1730 (N_1730,N_1384,N_1202);
or U1731 (N_1731,N_1281,N_1346);
nand U1732 (N_1732,N_1422,N_1311);
and U1733 (N_1733,N_1252,N_1302);
or U1734 (N_1734,N_1367,N_1420);
xor U1735 (N_1735,N_1372,N_1409);
or U1736 (N_1736,N_1255,N_1448);
nor U1737 (N_1737,N_1252,N_1208);
nor U1738 (N_1738,N_1315,N_1474);
nor U1739 (N_1739,N_1391,N_1453);
nor U1740 (N_1740,N_1226,N_1315);
xor U1741 (N_1741,N_1311,N_1202);
or U1742 (N_1742,N_1327,N_1456);
or U1743 (N_1743,N_1476,N_1208);
nor U1744 (N_1744,N_1380,N_1341);
or U1745 (N_1745,N_1362,N_1485);
or U1746 (N_1746,N_1207,N_1458);
and U1747 (N_1747,N_1362,N_1398);
and U1748 (N_1748,N_1219,N_1209);
nand U1749 (N_1749,N_1250,N_1285);
nand U1750 (N_1750,N_1388,N_1311);
xor U1751 (N_1751,N_1333,N_1441);
nor U1752 (N_1752,N_1498,N_1362);
and U1753 (N_1753,N_1344,N_1467);
and U1754 (N_1754,N_1366,N_1403);
and U1755 (N_1755,N_1271,N_1268);
and U1756 (N_1756,N_1249,N_1356);
nand U1757 (N_1757,N_1257,N_1261);
nand U1758 (N_1758,N_1405,N_1332);
and U1759 (N_1759,N_1290,N_1356);
or U1760 (N_1760,N_1244,N_1293);
and U1761 (N_1761,N_1365,N_1288);
and U1762 (N_1762,N_1466,N_1279);
or U1763 (N_1763,N_1411,N_1201);
and U1764 (N_1764,N_1395,N_1257);
xnor U1765 (N_1765,N_1473,N_1431);
nand U1766 (N_1766,N_1214,N_1263);
nand U1767 (N_1767,N_1227,N_1269);
and U1768 (N_1768,N_1380,N_1425);
and U1769 (N_1769,N_1484,N_1280);
xnor U1770 (N_1770,N_1206,N_1216);
nand U1771 (N_1771,N_1274,N_1356);
nor U1772 (N_1772,N_1458,N_1445);
or U1773 (N_1773,N_1461,N_1331);
or U1774 (N_1774,N_1441,N_1445);
and U1775 (N_1775,N_1312,N_1385);
and U1776 (N_1776,N_1341,N_1235);
nor U1777 (N_1777,N_1265,N_1363);
and U1778 (N_1778,N_1266,N_1243);
nor U1779 (N_1779,N_1299,N_1276);
nand U1780 (N_1780,N_1352,N_1417);
or U1781 (N_1781,N_1412,N_1287);
nor U1782 (N_1782,N_1212,N_1245);
nand U1783 (N_1783,N_1282,N_1212);
nor U1784 (N_1784,N_1463,N_1357);
or U1785 (N_1785,N_1256,N_1383);
or U1786 (N_1786,N_1320,N_1391);
and U1787 (N_1787,N_1213,N_1278);
xor U1788 (N_1788,N_1388,N_1467);
or U1789 (N_1789,N_1434,N_1309);
nor U1790 (N_1790,N_1219,N_1459);
and U1791 (N_1791,N_1430,N_1296);
xor U1792 (N_1792,N_1383,N_1350);
nand U1793 (N_1793,N_1473,N_1344);
nand U1794 (N_1794,N_1374,N_1286);
xor U1795 (N_1795,N_1205,N_1369);
xor U1796 (N_1796,N_1254,N_1393);
nand U1797 (N_1797,N_1305,N_1357);
nand U1798 (N_1798,N_1384,N_1459);
nand U1799 (N_1799,N_1419,N_1376);
and U1800 (N_1800,N_1634,N_1777);
nor U1801 (N_1801,N_1677,N_1590);
and U1802 (N_1802,N_1778,N_1592);
nor U1803 (N_1803,N_1760,N_1645);
or U1804 (N_1804,N_1669,N_1566);
xor U1805 (N_1805,N_1611,N_1723);
nand U1806 (N_1806,N_1773,N_1709);
xnor U1807 (N_1807,N_1516,N_1549);
or U1808 (N_1808,N_1730,N_1682);
or U1809 (N_1809,N_1787,N_1691);
or U1810 (N_1810,N_1714,N_1548);
or U1811 (N_1811,N_1716,N_1733);
xnor U1812 (N_1812,N_1593,N_1635);
nand U1813 (N_1813,N_1531,N_1776);
nor U1814 (N_1814,N_1704,N_1604);
xnor U1815 (N_1815,N_1613,N_1582);
or U1816 (N_1816,N_1581,N_1722);
nand U1817 (N_1817,N_1775,N_1553);
and U1818 (N_1818,N_1754,N_1732);
nor U1819 (N_1819,N_1622,N_1740);
xnor U1820 (N_1820,N_1711,N_1628);
xor U1821 (N_1821,N_1702,N_1794);
nor U1822 (N_1822,N_1657,N_1655);
or U1823 (N_1823,N_1623,N_1543);
nor U1824 (N_1824,N_1667,N_1699);
or U1825 (N_1825,N_1643,N_1560);
nand U1826 (N_1826,N_1675,N_1670);
nand U1827 (N_1827,N_1644,N_1523);
xnor U1828 (N_1828,N_1517,N_1743);
nand U1829 (N_1829,N_1719,N_1642);
xor U1830 (N_1830,N_1568,N_1756);
and U1831 (N_1831,N_1753,N_1551);
and U1832 (N_1832,N_1652,N_1511);
xor U1833 (N_1833,N_1701,N_1676);
and U1834 (N_1834,N_1533,N_1619);
nand U1835 (N_1835,N_1700,N_1735);
nor U1836 (N_1836,N_1665,N_1745);
and U1837 (N_1837,N_1569,N_1542);
or U1838 (N_1838,N_1561,N_1715);
xor U1839 (N_1839,N_1658,N_1651);
nand U1840 (N_1840,N_1736,N_1600);
nand U1841 (N_1841,N_1536,N_1605);
nor U1842 (N_1842,N_1638,N_1718);
xnor U1843 (N_1843,N_1510,N_1545);
or U1844 (N_1844,N_1640,N_1694);
xnor U1845 (N_1845,N_1692,N_1668);
nor U1846 (N_1846,N_1578,N_1693);
and U1847 (N_1847,N_1729,N_1526);
nor U1848 (N_1848,N_1564,N_1686);
nand U1849 (N_1849,N_1666,N_1507);
nor U1850 (N_1850,N_1724,N_1646);
or U1851 (N_1851,N_1552,N_1731);
nor U1852 (N_1852,N_1734,N_1575);
and U1853 (N_1853,N_1793,N_1664);
xnor U1854 (N_1854,N_1789,N_1779);
nor U1855 (N_1855,N_1620,N_1741);
xor U1856 (N_1856,N_1653,N_1795);
xor U1857 (N_1857,N_1601,N_1727);
nand U1858 (N_1858,N_1521,N_1504);
nor U1859 (N_1859,N_1746,N_1541);
nor U1860 (N_1860,N_1555,N_1608);
or U1861 (N_1861,N_1617,N_1757);
nand U1862 (N_1862,N_1728,N_1750);
or U1863 (N_1863,N_1609,N_1572);
nand U1864 (N_1864,N_1546,N_1559);
nand U1865 (N_1865,N_1500,N_1678);
or U1866 (N_1866,N_1720,N_1632);
nand U1867 (N_1867,N_1594,N_1796);
and U1868 (N_1868,N_1529,N_1766);
or U1869 (N_1869,N_1610,N_1544);
nand U1870 (N_1870,N_1607,N_1615);
nor U1871 (N_1871,N_1554,N_1573);
xor U1872 (N_1872,N_1621,N_1626);
nand U1873 (N_1873,N_1770,N_1528);
and U1874 (N_1874,N_1631,N_1637);
or U1875 (N_1875,N_1713,N_1788);
xor U1876 (N_1876,N_1574,N_1580);
nand U1877 (N_1877,N_1761,N_1616);
or U1878 (N_1878,N_1768,N_1749);
and U1879 (N_1879,N_1738,N_1527);
and U1880 (N_1880,N_1570,N_1707);
or U1881 (N_1881,N_1641,N_1703);
nand U1882 (N_1882,N_1647,N_1679);
xnor U1883 (N_1883,N_1625,N_1758);
and U1884 (N_1884,N_1649,N_1721);
nor U1885 (N_1885,N_1525,N_1774);
or U1886 (N_1886,N_1726,N_1747);
xnor U1887 (N_1887,N_1662,N_1509);
or U1888 (N_1888,N_1639,N_1712);
xor U1889 (N_1889,N_1587,N_1519);
xnor U1890 (N_1890,N_1614,N_1524);
nand U1891 (N_1891,N_1798,N_1556);
xor U1892 (N_1892,N_1764,N_1799);
nand U1893 (N_1893,N_1748,N_1576);
or U1894 (N_1894,N_1530,N_1739);
xnor U1895 (N_1895,N_1598,N_1690);
nand U1896 (N_1896,N_1629,N_1624);
or U1897 (N_1897,N_1599,N_1681);
and U1898 (N_1898,N_1636,N_1503);
and U1899 (N_1899,N_1661,N_1762);
or U1900 (N_1900,N_1537,N_1782);
nor U1901 (N_1901,N_1786,N_1680);
or U1902 (N_1902,N_1591,N_1520);
xor U1903 (N_1903,N_1742,N_1585);
nand U1904 (N_1904,N_1683,N_1538);
and U1905 (N_1905,N_1654,N_1535);
nor U1906 (N_1906,N_1577,N_1684);
and U1907 (N_1907,N_1596,N_1685);
and U1908 (N_1908,N_1648,N_1562);
nand U1909 (N_1909,N_1784,N_1797);
or U1910 (N_1910,N_1588,N_1563);
and U1911 (N_1911,N_1514,N_1558);
nor U1912 (N_1912,N_1759,N_1710);
xnor U1913 (N_1913,N_1790,N_1547);
or U1914 (N_1914,N_1671,N_1557);
and U1915 (N_1915,N_1717,N_1532);
and U1916 (N_1916,N_1705,N_1550);
nand U1917 (N_1917,N_1650,N_1744);
nor U1918 (N_1918,N_1505,N_1752);
nor U1919 (N_1919,N_1534,N_1763);
and U1920 (N_1920,N_1508,N_1755);
nor U1921 (N_1921,N_1674,N_1772);
and U1922 (N_1922,N_1771,N_1565);
or U1923 (N_1923,N_1571,N_1579);
xor U1924 (N_1924,N_1502,N_1780);
nand U1925 (N_1925,N_1540,N_1697);
or U1926 (N_1926,N_1751,N_1785);
nand U1927 (N_1927,N_1696,N_1501);
or U1928 (N_1928,N_1627,N_1737);
and U1929 (N_1929,N_1513,N_1688);
and U1930 (N_1930,N_1602,N_1708);
xor U1931 (N_1931,N_1695,N_1595);
and U1932 (N_1932,N_1583,N_1515);
nor U1933 (N_1933,N_1769,N_1586);
xor U1934 (N_1934,N_1512,N_1672);
nand U1935 (N_1935,N_1689,N_1603);
or U1936 (N_1936,N_1606,N_1589);
and U1937 (N_1937,N_1659,N_1618);
nand U1938 (N_1938,N_1660,N_1663);
xor U1939 (N_1939,N_1584,N_1522);
and U1940 (N_1940,N_1706,N_1792);
xnor U1941 (N_1941,N_1612,N_1698);
nor U1942 (N_1942,N_1725,N_1656);
and U1943 (N_1943,N_1506,N_1687);
or U1944 (N_1944,N_1767,N_1765);
and U1945 (N_1945,N_1633,N_1597);
nand U1946 (N_1946,N_1781,N_1783);
and U1947 (N_1947,N_1673,N_1630);
or U1948 (N_1948,N_1791,N_1518);
or U1949 (N_1949,N_1539,N_1567);
nand U1950 (N_1950,N_1594,N_1736);
and U1951 (N_1951,N_1724,N_1589);
and U1952 (N_1952,N_1548,N_1604);
nand U1953 (N_1953,N_1570,N_1526);
nand U1954 (N_1954,N_1737,N_1713);
and U1955 (N_1955,N_1521,N_1597);
nand U1956 (N_1956,N_1684,N_1548);
or U1957 (N_1957,N_1602,N_1765);
xor U1958 (N_1958,N_1592,N_1540);
xnor U1959 (N_1959,N_1610,N_1686);
and U1960 (N_1960,N_1669,N_1764);
xor U1961 (N_1961,N_1720,N_1537);
nand U1962 (N_1962,N_1544,N_1531);
or U1963 (N_1963,N_1770,N_1513);
xnor U1964 (N_1964,N_1650,N_1565);
nor U1965 (N_1965,N_1689,N_1794);
and U1966 (N_1966,N_1545,N_1658);
and U1967 (N_1967,N_1620,N_1645);
xor U1968 (N_1968,N_1598,N_1633);
and U1969 (N_1969,N_1601,N_1641);
and U1970 (N_1970,N_1707,N_1584);
nor U1971 (N_1971,N_1689,N_1686);
nor U1972 (N_1972,N_1782,N_1727);
and U1973 (N_1973,N_1771,N_1796);
nand U1974 (N_1974,N_1611,N_1516);
nand U1975 (N_1975,N_1727,N_1642);
nand U1976 (N_1976,N_1593,N_1547);
and U1977 (N_1977,N_1789,N_1559);
nor U1978 (N_1978,N_1752,N_1607);
xor U1979 (N_1979,N_1759,N_1521);
nor U1980 (N_1980,N_1555,N_1645);
nand U1981 (N_1981,N_1745,N_1541);
or U1982 (N_1982,N_1701,N_1720);
nor U1983 (N_1983,N_1725,N_1602);
xnor U1984 (N_1984,N_1594,N_1688);
or U1985 (N_1985,N_1668,N_1726);
nand U1986 (N_1986,N_1711,N_1569);
or U1987 (N_1987,N_1623,N_1673);
nand U1988 (N_1988,N_1770,N_1626);
nand U1989 (N_1989,N_1696,N_1702);
nor U1990 (N_1990,N_1799,N_1545);
and U1991 (N_1991,N_1674,N_1716);
and U1992 (N_1992,N_1598,N_1726);
nor U1993 (N_1993,N_1555,N_1743);
xnor U1994 (N_1994,N_1532,N_1618);
or U1995 (N_1995,N_1501,N_1554);
or U1996 (N_1996,N_1552,N_1637);
nor U1997 (N_1997,N_1794,N_1703);
or U1998 (N_1998,N_1739,N_1555);
nand U1999 (N_1999,N_1753,N_1653);
nor U2000 (N_2000,N_1571,N_1583);
xnor U2001 (N_2001,N_1687,N_1781);
xor U2002 (N_2002,N_1545,N_1704);
xnor U2003 (N_2003,N_1756,N_1785);
nand U2004 (N_2004,N_1633,N_1692);
or U2005 (N_2005,N_1610,N_1588);
xor U2006 (N_2006,N_1593,N_1648);
or U2007 (N_2007,N_1747,N_1571);
or U2008 (N_2008,N_1732,N_1781);
nand U2009 (N_2009,N_1733,N_1765);
and U2010 (N_2010,N_1728,N_1773);
and U2011 (N_2011,N_1681,N_1742);
and U2012 (N_2012,N_1549,N_1510);
or U2013 (N_2013,N_1699,N_1547);
xor U2014 (N_2014,N_1692,N_1591);
or U2015 (N_2015,N_1716,N_1671);
and U2016 (N_2016,N_1552,N_1794);
nand U2017 (N_2017,N_1719,N_1666);
and U2018 (N_2018,N_1714,N_1572);
or U2019 (N_2019,N_1691,N_1669);
nand U2020 (N_2020,N_1651,N_1557);
and U2021 (N_2021,N_1798,N_1769);
and U2022 (N_2022,N_1562,N_1554);
and U2023 (N_2023,N_1538,N_1690);
xor U2024 (N_2024,N_1718,N_1597);
or U2025 (N_2025,N_1560,N_1726);
nand U2026 (N_2026,N_1749,N_1726);
nand U2027 (N_2027,N_1665,N_1702);
nor U2028 (N_2028,N_1602,N_1606);
or U2029 (N_2029,N_1719,N_1531);
and U2030 (N_2030,N_1569,N_1683);
or U2031 (N_2031,N_1721,N_1578);
nand U2032 (N_2032,N_1786,N_1769);
and U2033 (N_2033,N_1504,N_1649);
nor U2034 (N_2034,N_1554,N_1520);
xor U2035 (N_2035,N_1760,N_1663);
xor U2036 (N_2036,N_1668,N_1708);
xnor U2037 (N_2037,N_1573,N_1567);
xor U2038 (N_2038,N_1653,N_1736);
nand U2039 (N_2039,N_1664,N_1545);
and U2040 (N_2040,N_1760,N_1761);
nand U2041 (N_2041,N_1574,N_1511);
and U2042 (N_2042,N_1673,N_1667);
nand U2043 (N_2043,N_1674,N_1775);
xnor U2044 (N_2044,N_1697,N_1745);
xnor U2045 (N_2045,N_1793,N_1583);
nand U2046 (N_2046,N_1689,N_1788);
or U2047 (N_2047,N_1734,N_1612);
or U2048 (N_2048,N_1686,N_1546);
or U2049 (N_2049,N_1721,N_1504);
or U2050 (N_2050,N_1548,N_1620);
and U2051 (N_2051,N_1769,N_1545);
xnor U2052 (N_2052,N_1518,N_1658);
nor U2053 (N_2053,N_1640,N_1606);
nor U2054 (N_2054,N_1742,N_1777);
and U2055 (N_2055,N_1757,N_1563);
or U2056 (N_2056,N_1766,N_1557);
and U2057 (N_2057,N_1577,N_1720);
or U2058 (N_2058,N_1505,N_1707);
or U2059 (N_2059,N_1761,N_1617);
nor U2060 (N_2060,N_1555,N_1554);
nand U2061 (N_2061,N_1616,N_1572);
nor U2062 (N_2062,N_1522,N_1625);
nand U2063 (N_2063,N_1641,N_1522);
xor U2064 (N_2064,N_1785,N_1589);
or U2065 (N_2065,N_1618,N_1670);
nor U2066 (N_2066,N_1539,N_1523);
xor U2067 (N_2067,N_1616,N_1629);
nor U2068 (N_2068,N_1637,N_1589);
nor U2069 (N_2069,N_1775,N_1602);
xnor U2070 (N_2070,N_1543,N_1569);
and U2071 (N_2071,N_1768,N_1598);
nor U2072 (N_2072,N_1573,N_1579);
nor U2073 (N_2073,N_1500,N_1756);
nand U2074 (N_2074,N_1691,N_1769);
or U2075 (N_2075,N_1561,N_1565);
nand U2076 (N_2076,N_1500,N_1653);
xor U2077 (N_2077,N_1541,N_1502);
nor U2078 (N_2078,N_1519,N_1764);
xnor U2079 (N_2079,N_1765,N_1530);
xnor U2080 (N_2080,N_1626,N_1731);
xnor U2081 (N_2081,N_1638,N_1774);
xnor U2082 (N_2082,N_1732,N_1524);
xor U2083 (N_2083,N_1705,N_1544);
xnor U2084 (N_2084,N_1747,N_1638);
nor U2085 (N_2085,N_1626,N_1559);
and U2086 (N_2086,N_1520,N_1692);
or U2087 (N_2087,N_1700,N_1572);
or U2088 (N_2088,N_1507,N_1770);
xnor U2089 (N_2089,N_1723,N_1674);
nor U2090 (N_2090,N_1537,N_1567);
nand U2091 (N_2091,N_1573,N_1756);
or U2092 (N_2092,N_1725,N_1731);
xnor U2093 (N_2093,N_1573,N_1590);
xor U2094 (N_2094,N_1501,N_1639);
nor U2095 (N_2095,N_1550,N_1684);
xor U2096 (N_2096,N_1754,N_1704);
or U2097 (N_2097,N_1576,N_1664);
xor U2098 (N_2098,N_1548,N_1744);
or U2099 (N_2099,N_1683,N_1691);
or U2100 (N_2100,N_2057,N_1904);
xor U2101 (N_2101,N_1810,N_1966);
xor U2102 (N_2102,N_2023,N_1940);
and U2103 (N_2103,N_2084,N_2063);
or U2104 (N_2104,N_1985,N_1854);
nor U2105 (N_2105,N_1884,N_1891);
nand U2106 (N_2106,N_1802,N_2049);
and U2107 (N_2107,N_1963,N_2008);
nand U2108 (N_2108,N_1961,N_1839);
and U2109 (N_2109,N_1995,N_2093);
or U2110 (N_2110,N_1820,N_1841);
nor U2111 (N_2111,N_2091,N_2012);
or U2112 (N_2112,N_1993,N_2036);
and U2113 (N_2113,N_1831,N_2058);
nand U2114 (N_2114,N_1875,N_1980);
nor U2115 (N_2115,N_1988,N_1885);
nand U2116 (N_2116,N_2086,N_1919);
nor U2117 (N_2117,N_1974,N_1941);
nand U2118 (N_2118,N_1912,N_1836);
and U2119 (N_2119,N_1860,N_1849);
or U2120 (N_2120,N_1967,N_2020);
or U2121 (N_2121,N_1817,N_2030);
or U2122 (N_2122,N_1943,N_1812);
nand U2123 (N_2123,N_2077,N_1942);
nor U2124 (N_2124,N_2015,N_1896);
nor U2125 (N_2125,N_1801,N_1981);
and U2126 (N_2126,N_1951,N_1892);
xor U2127 (N_2127,N_1999,N_1870);
nor U2128 (N_2128,N_2098,N_2089);
or U2129 (N_2129,N_2054,N_2074);
xnor U2130 (N_2130,N_1983,N_1960);
and U2131 (N_2131,N_1846,N_1856);
and U2132 (N_2132,N_1866,N_1970);
nand U2133 (N_2133,N_1857,N_2043);
xor U2134 (N_2134,N_1933,N_1872);
nand U2135 (N_2135,N_1911,N_1874);
nor U2136 (N_2136,N_2048,N_2018);
nand U2137 (N_2137,N_2067,N_2081);
xor U2138 (N_2138,N_2097,N_1957);
nor U2139 (N_2139,N_1805,N_1915);
nor U2140 (N_2140,N_2078,N_1806);
nand U2141 (N_2141,N_1989,N_1950);
and U2142 (N_2142,N_1962,N_1876);
xor U2143 (N_2143,N_2073,N_2062);
nand U2144 (N_2144,N_1869,N_2010);
xor U2145 (N_2145,N_1819,N_1845);
nand U2146 (N_2146,N_2050,N_1926);
or U2147 (N_2147,N_1882,N_1871);
or U2148 (N_2148,N_2006,N_2021);
xor U2149 (N_2149,N_2080,N_1852);
nor U2150 (N_2150,N_2072,N_2040);
and U2151 (N_2151,N_1978,N_1826);
or U2152 (N_2152,N_2019,N_2009);
or U2153 (N_2153,N_2029,N_1890);
xor U2154 (N_2154,N_2092,N_1979);
or U2155 (N_2155,N_1928,N_1982);
or U2156 (N_2156,N_1834,N_2033);
and U2157 (N_2157,N_1977,N_1828);
nor U2158 (N_2158,N_1865,N_2000);
xnor U2159 (N_2159,N_1991,N_2065);
xor U2160 (N_2160,N_2056,N_1868);
nand U2161 (N_2161,N_1804,N_1944);
or U2162 (N_2162,N_1996,N_2037);
nand U2163 (N_2163,N_1986,N_1863);
or U2164 (N_2164,N_1948,N_1922);
and U2165 (N_2165,N_1864,N_1968);
nor U2166 (N_2166,N_2053,N_2026);
xnor U2167 (N_2167,N_1908,N_2028);
and U2168 (N_2168,N_2014,N_1859);
nand U2169 (N_2169,N_2004,N_1842);
or U2170 (N_2170,N_2096,N_2007);
nand U2171 (N_2171,N_1910,N_1907);
and U2172 (N_2172,N_1814,N_2041);
and U2173 (N_2173,N_1965,N_2095);
nor U2174 (N_2174,N_2045,N_1822);
and U2175 (N_2175,N_1877,N_1920);
nor U2176 (N_2176,N_1843,N_2083);
nor U2177 (N_2177,N_2003,N_2085);
and U2178 (N_2178,N_2070,N_2090);
and U2179 (N_2179,N_1823,N_2076);
nor U2180 (N_2180,N_2046,N_1878);
or U2181 (N_2181,N_1830,N_2088);
and U2182 (N_2182,N_1815,N_1899);
and U2183 (N_2183,N_1809,N_1800);
or U2184 (N_2184,N_1909,N_2002);
xor U2185 (N_2185,N_1807,N_1946);
nand U2186 (N_2186,N_2059,N_2071);
and U2187 (N_2187,N_1903,N_1984);
nand U2188 (N_2188,N_1932,N_2017);
nor U2189 (N_2189,N_1927,N_1888);
and U2190 (N_2190,N_1976,N_1987);
xnor U2191 (N_2191,N_1808,N_1913);
xor U2192 (N_2192,N_1886,N_1959);
xnor U2193 (N_2193,N_2013,N_2005);
nor U2194 (N_2194,N_2027,N_1937);
xor U2195 (N_2195,N_1955,N_2034);
or U2196 (N_2196,N_2052,N_1825);
or U2197 (N_2197,N_1821,N_2016);
and U2198 (N_2198,N_1939,N_1952);
nand U2199 (N_2199,N_2038,N_1971);
nor U2200 (N_2200,N_1931,N_1853);
or U2201 (N_2201,N_1829,N_1850);
nor U2202 (N_2202,N_1835,N_1935);
or U2203 (N_2203,N_1900,N_1827);
nor U2204 (N_2204,N_1905,N_1969);
or U2205 (N_2205,N_1925,N_1918);
nand U2206 (N_2206,N_1883,N_1824);
and U2207 (N_2207,N_1880,N_1964);
xor U2208 (N_2208,N_1894,N_2022);
nand U2209 (N_2209,N_1945,N_1994);
or U2210 (N_2210,N_1897,N_2055);
nor U2211 (N_2211,N_1833,N_1923);
nor U2212 (N_2212,N_2066,N_1916);
xnor U2213 (N_2213,N_2060,N_1902);
nor U2214 (N_2214,N_1803,N_2082);
xor U2215 (N_2215,N_1848,N_1818);
nor U2216 (N_2216,N_1873,N_1816);
and U2217 (N_2217,N_2032,N_1956);
nand U2218 (N_2218,N_2087,N_1832);
nand U2219 (N_2219,N_2069,N_2064);
nand U2220 (N_2220,N_2035,N_2024);
nand U2221 (N_2221,N_1837,N_1917);
xnor U2222 (N_2222,N_2099,N_1858);
xnor U2223 (N_2223,N_1949,N_1975);
nand U2224 (N_2224,N_1893,N_1990);
xnor U2225 (N_2225,N_1898,N_2011);
xnor U2226 (N_2226,N_1914,N_2047);
nand U2227 (N_2227,N_1954,N_1838);
nor U2228 (N_2228,N_1879,N_1861);
nand U2229 (N_2229,N_1953,N_2079);
and U2230 (N_2230,N_1938,N_1881);
and U2231 (N_2231,N_2094,N_1887);
or U2232 (N_2232,N_2061,N_1847);
or U2233 (N_2233,N_1851,N_1992);
nand U2234 (N_2234,N_1972,N_1930);
nor U2235 (N_2235,N_1958,N_1867);
and U2236 (N_2236,N_1840,N_2051);
or U2237 (N_2237,N_2068,N_1947);
nand U2238 (N_2238,N_1889,N_2001);
xor U2239 (N_2239,N_1936,N_1973);
xor U2240 (N_2240,N_2025,N_1855);
nand U2241 (N_2241,N_2044,N_1906);
xnor U2242 (N_2242,N_2042,N_1901);
or U2243 (N_2243,N_1997,N_1924);
xor U2244 (N_2244,N_1844,N_1929);
xnor U2245 (N_2245,N_1813,N_1811);
nand U2246 (N_2246,N_1934,N_1921);
nor U2247 (N_2247,N_2039,N_1998);
nand U2248 (N_2248,N_2031,N_1895);
xor U2249 (N_2249,N_2075,N_1862);
nand U2250 (N_2250,N_1809,N_1801);
xor U2251 (N_2251,N_2093,N_2025);
and U2252 (N_2252,N_2065,N_2031);
or U2253 (N_2253,N_2026,N_1859);
or U2254 (N_2254,N_1891,N_1950);
nand U2255 (N_2255,N_1890,N_2040);
or U2256 (N_2256,N_1895,N_2065);
nor U2257 (N_2257,N_1824,N_1945);
nand U2258 (N_2258,N_2018,N_2036);
nand U2259 (N_2259,N_1938,N_2006);
nor U2260 (N_2260,N_2021,N_1834);
or U2261 (N_2261,N_1997,N_1953);
nand U2262 (N_2262,N_2061,N_1933);
nor U2263 (N_2263,N_1886,N_1905);
or U2264 (N_2264,N_1964,N_1864);
nand U2265 (N_2265,N_1818,N_1825);
nand U2266 (N_2266,N_2091,N_1978);
and U2267 (N_2267,N_1813,N_1957);
and U2268 (N_2268,N_2008,N_1957);
xnor U2269 (N_2269,N_1935,N_1846);
xnor U2270 (N_2270,N_1911,N_1906);
xor U2271 (N_2271,N_1916,N_1861);
nor U2272 (N_2272,N_1801,N_1910);
xnor U2273 (N_2273,N_1809,N_2066);
and U2274 (N_2274,N_1953,N_1947);
nand U2275 (N_2275,N_1948,N_2062);
and U2276 (N_2276,N_2035,N_2070);
nor U2277 (N_2277,N_1974,N_1922);
xor U2278 (N_2278,N_2034,N_1872);
nand U2279 (N_2279,N_1862,N_1890);
nand U2280 (N_2280,N_1841,N_1974);
xor U2281 (N_2281,N_1903,N_1915);
nand U2282 (N_2282,N_1994,N_2078);
and U2283 (N_2283,N_1895,N_1851);
nand U2284 (N_2284,N_2038,N_1827);
and U2285 (N_2285,N_1931,N_1998);
nand U2286 (N_2286,N_2049,N_2021);
nand U2287 (N_2287,N_1825,N_1815);
nand U2288 (N_2288,N_1960,N_1816);
or U2289 (N_2289,N_1996,N_1951);
nor U2290 (N_2290,N_2097,N_2066);
nand U2291 (N_2291,N_1998,N_1829);
nor U2292 (N_2292,N_1955,N_1996);
nand U2293 (N_2293,N_1803,N_1914);
nand U2294 (N_2294,N_2097,N_2036);
or U2295 (N_2295,N_1847,N_2063);
xnor U2296 (N_2296,N_1855,N_1891);
or U2297 (N_2297,N_1949,N_1895);
and U2298 (N_2298,N_1899,N_1803);
nand U2299 (N_2299,N_1972,N_2070);
and U2300 (N_2300,N_2068,N_1866);
or U2301 (N_2301,N_2036,N_1926);
and U2302 (N_2302,N_1822,N_1912);
or U2303 (N_2303,N_2004,N_1899);
nand U2304 (N_2304,N_1910,N_2076);
nand U2305 (N_2305,N_1918,N_2039);
xor U2306 (N_2306,N_1801,N_2093);
xor U2307 (N_2307,N_1818,N_1956);
and U2308 (N_2308,N_2082,N_1848);
xor U2309 (N_2309,N_1992,N_2014);
xor U2310 (N_2310,N_1923,N_1860);
xnor U2311 (N_2311,N_1937,N_1976);
nand U2312 (N_2312,N_2053,N_1885);
or U2313 (N_2313,N_1925,N_1840);
or U2314 (N_2314,N_2084,N_2078);
or U2315 (N_2315,N_1805,N_1824);
nor U2316 (N_2316,N_2065,N_2020);
nor U2317 (N_2317,N_2053,N_2056);
nor U2318 (N_2318,N_2066,N_2072);
nor U2319 (N_2319,N_1892,N_1933);
nor U2320 (N_2320,N_1902,N_1966);
nor U2321 (N_2321,N_1927,N_2096);
or U2322 (N_2322,N_1838,N_1826);
or U2323 (N_2323,N_1926,N_1871);
nand U2324 (N_2324,N_2074,N_1834);
nor U2325 (N_2325,N_2004,N_2066);
and U2326 (N_2326,N_2088,N_1897);
nor U2327 (N_2327,N_2023,N_1987);
nor U2328 (N_2328,N_1967,N_2040);
or U2329 (N_2329,N_2020,N_1912);
and U2330 (N_2330,N_1968,N_1954);
nor U2331 (N_2331,N_1983,N_1985);
or U2332 (N_2332,N_1982,N_1971);
nand U2333 (N_2333,N_1927,N_1904);
xor U2334 (N_2334,N_1807,N_1801);
xor U2335 (N_2335,N_2049,N_2069);
or U2336 (N_2336,N_1901,N_2011);
xnor U2337 (N_2337,N_1993,N_2004);
xor U2338 (N_2338,N_1969,N_1914);
nand U2339 (N_2339,N_2065,N_2063);
nor U2340 (N_2340,N_2095,N_1966);
or U2341 (N_2341,N_2044,N_1882);
nor U2342 (N_2342,N_1870,N_1952);
or U2343 (N_2343,N_1878,N_2004);
and U2344 (N_2344,N_1911,N_1892);
and U2345 (N_2345,N_1967,N_1860);
and U2346 (N_2346,N_2062,N_1922);
xnor U2347 (N_2347,N_1805,N_1899);
xor U2348 (N_2348,N_2041,N_1848);
xor U2349 (N_2349,N_2068,N_2053);
xnor U2350 (N_2350,N_1981,N_2098);
nor U2351 (N_2351,N_1947,N_1887);
nor U2352 (N_2352,N_2013,N_1936);
or U2353 (N_2353,N_2003,N_2058);
or U2354 (N_2354,N_1928,N_1960);
and U2355 (N_2355,N_2076,N_1853);
nand U2356 (N_2356,N_1809,N_1831);
and U2357 (N_2357,N_1955,N_1828);
and U2358 (N_2358,N_2014,N_2000);
xor U2359 (N_2359,N_1979,N_2062);
and U2360 (N_2360,N_2066,N_1956);
or U2361 (N_2361,N_1927,N_1953);
and U2362 (N_2362,N_1825,N_2028);
or U2363 (N_2363,N_1827,N_2071);
or U2364 (N_2364,N_1997,N_2042);
nor U2365 (N_2365,N_1812,N_1941);
xnor U2366 (N_2366,N_1936,N_1988);
or U2367 (N_2367,N_1826,N_2041);
xor U2368 (N_2368,N_2075,N_1922);
and U2369 (N_2369,N_1929,N_1966);
xor U2370 (N_2370,N_2005,N_1977);
nor U2371 (N_2371,N_1999,N_1920);
or U2372 (N_2372,N_2050,N_1955);
nor U2373 (N_2373,N_1914,N_2062);
and U2374 (N_2374,N_1977,N_1895);
nor U2375 (N_2375,N_1845,N_2087);
or U2376 (N_2376,N_1968,N_2007);
or U2377 (N_2377,N_2045,N_2030);
xnor U2378 (N_2378,N_2066,N_1901);
nand U2379 (N_2379,N_2047,N_2099);
or U2380 (N_2380,N_2003,N_1881);
and U2381 (N_2381,N_1977,N_2045);
and U2382 (N_2382,N_2081,N_2001);
or U2383 (N_2383,N_1874,N_2048);
or U2384 (N_2384,N_1982,N_1886);
nor U2385 (N_2385,N_2071,N_1888);
nand U2386 (N_2386,N_1944,N_1884);
xor U2387 (N_2387,N_2053,N_2015);
nor U2388 (N_2388,N_1902,N_2096);
or U2389 (N_2389,N_1997,N_2034);
or U2390 (N_2390,N_1967,N_2041);
or U2391 (N_2391,N_1912,N_1991);
nor U2392 (N_2392,N_1818,N_1943);
xnor U2393 (N_2393,N_1825,N_1951);
nand U2394 (N_2394,N_2027,N_1949);
nand U2395 (N_2395,N_1935,N_2026);
xnor U2396 (N_2396,N_1973,N_1922);
nand U2397 (N_2397,N_1885,N_1994);
xor U2398 (N_2398,N_2063,N_1985);
xor U2399 (N_2399,N_1937,N_1815);
xnor U2400 (N_2400,N_2259,N_2187);
and U2401 (N_2401,N_2194,N_2224);
nand U2402 (N_2402,N_2214,N_2385);
xor U2403 (N_2403,N_2206,N_2389);
nor U2404 (N_2404,N_2218,N_2268);
and U2405 (N_2405,N_2276,N_2273);
and U2406 (N_2406,N_2314,N_2195);
nand U2407 (N_2407,N_2118,N_2226);
nand U2408 (N_2408,N_2179,N_2184);
nor U2409 (N_2409,N_2333,N_2126);
nand U2410 (N_2410,N_2243,N_2166);
or U2411 (N_2411,N_2341,N_2233);
nand U2412 (N_2412,N_2147,N_2338);
nand U2413 (N_2413,N_2145,N_2327);
nor U2414 (N_2414,N_2294,N_2173);
or U2415 (N_2415,N_2161,N_2111);
and U2416 (N_2416,N_2134,N_2106);
nand U2417 (N_2417,N_2232,N_2177);
nand U2418 (N_2418,N_2277,N_2258);
xnor U2419 (N_2419,N_2307,N_2153);
nand U2420 (N_2420,N_2114,N_2352);
nor U2421 (N_2421,N_2304,N_2135);
nand U2422 (N_2422,N_2255,N_2183);
xnor U2423 (N_2423,N_2387,N_2140);
nand U2424 (N_2424,N_2119,N_2384);
nor U2425 (N_2425,N_2355,N_2128);
nand U2426 (N_2426,N_2246,N_2220);
or U2427 (N_2427,N_2347,N_2150);
nor U2428 (N_2428,N_2256,N_2160);
xor U2429 (N_2429,N_2320,N_2264);
xor U2430 (N_2430,N_2180,N_2104);
nand U2431 (N_2431,N_2289,N_2253);
nor U2432 (N_2432,N_2288,N_2275);
xnor U2433 (N_2433,N_2379,N_2337);
nand U2434 (N_2434,N_2348,N_2192);
and U2435 (N_2435,N_2241,N_2157);
and U2436 (N_2436,N_2269,N_2176);
nand U2437 (N_2437,N_2235,N_2170);
and U2438 (N_2438,N_2399,N_2281);
nand U2439 (N_2439,N_2371,N_2367);
xor U2440 (N_2440,N_2318,N_2132);
xnor U2441 (N_2441,N_2257,N_2356);
nand U2442 (N_2442,N_2182,N_2368);
xor U2443 (N_2443,N_2110,N_2383);
and U2444 (N_2444,N_2291,N_2357);
xor U2445 (N_2445,N_2321,N_2252);
nor U2446 (N_2446,N_2133,N_2155);
xnor U2447 (N_2447,N_2260,N_2373);
nor U2448 (N_2448,N_2390,N_2293);
nand U2449 (N_2449,N_2353,N_2196);
and U2450 (N_2450,N_2113,N_2237);
nand U2451 (N_2451,N_2365,N_2267);
xnor U2452 (N_2452,N_2181,N_2372);
nor U2453 (N_2453,N_2343,N_2370);
xor U2454 (N_2454,N_2167,N_2362);
or U2455 (N_2455,N_2162,N_2398);
nand U2456 (N_2456,N_2396,N_2199);
nor U2457 (N_2457,N_2397,N_2313);
nor U2458 (N_2458,N_2236,N_2139);
nand U2459 (N_2459,N_2100,N_2102);
or U2460 (N_2460,N_2244,N_2231);
or U2461 (N_2461,N_2363,N_2219);
nor U2462 (N_2462,N_2287,N_2301);
xor U2463 (N_2463,N_2223,N_2266);
or U2464 (N_2464,N_2250,N_2271);
or U2465 (N_2465,N_2221,N_2366);
xor U2466 (N_2466,N_2329,N_2361);
xnor U2467 (N_2467,N_2208,N_2358);
nand U2468 (N_2468,N_2107,N_2332);
nand U2469 (N_2469,N_2309,N_2229);
xnor U2470 (N_2470,N_2340,N_2350);
nor U2471 (N_2471,N_2178,N_2303);
or U2472 (N_2472,N_2212,N_2127);
and U2473 (N_2473,N_2283,N_2117);
nor U2474 (N_2474,N_2130,N_2225);
nand U2475 (N_2475,N_2322,N_2354);
xnor U2476 (N_2476,N_2315,N_2146);
and U2477 (N_2477,N_2164,N_2345);
and U2478 (N_2478,N_2349,N_2308);
and U2479 (N_2479,N_2175,N_2359);
or U2480 (N_2480,N_2109,N_2156);
nand U2481 (N_2481,N_2163,N_2121);
nor U2482 (N_2482,N_2284,N_2207);
xnor U2483 (N_2483,N_2278,N_2346);
or U2484 (N_2484,N_2108,N_2395);
and U2485 (N_2485,N_2136,N_2190);
nand U2486 (N_2486,N_2209,N_2274);
and U2487 (N_2487,N_2377,N_2115);
or U2488 (N_2488,N_2238,N_2201);
nand U2489 (N_2489,N_2272,N_2138);
and U2490 (N_2490,N_2120,N_2101);
or U2491 (N_2491,N_2171,N_2339);
xnor U2492 (N_2492,N_2137,N_2296);
and U2493 (N_2493,N_2311,N_2290);
nor U2494 (N_2494,N_2230,N_2213);
or U2495 (N_2495,N_2143,N_2248);
or U2496 (N_2496,N_2263,N_2205);
nand U2497 (N_2497,N_2103,N_2188);
nor U2498 (N_2498,N_2382,N_2215);
nand U2499 (N_2499,N_2391,N_2282);
nand U2500 (N_2500,N_2305,N_2328);
nor U2501 (N_2501,N_2154,N_2151);
and U2502 (N_2502,N_2388,N_2342);
or U2503 (N_2503,N_2351,N_2186);
or U2504 (N_2504,N_2394,N_2381);
nor U2505 (N_2505,N_2240,N_2189);
nand U2506 (N_2506,N_2112,N_2380);
or U2507 (N_2507,N_2203,N_2168);
nand U2508 (N_2508,N_2302,N_2317);
nand U2509 (N_2509,N_2142,N_2286);
nor U2510 (N_2510,N_2210,N_2265);
nand U2511 (N_2511,N_2280,N_2279);
nor U2512 (N_2512,N_2193,N_2295);
nor U2513 (N_2513,N_2191,N_2222);
and U2514 (N_2514,N_2234,N_2122);
and U2515 (N_2515,N_2262,N_2334);
and U2516 (N_2516,N_2105,N_2148);
and U2517 (N_2517,N_2299,N_2324);
nor U2518 (N_2518,N_2197,N_2141);
nand U2519 (N_2519,N_2227,N_2323);
and U2520 (N_2520,N_2306,N_2254);
nor U2521 (N_2521,N_2393,N_2217);
xor U2522 (N_2522,N_2242,N_2131);
and U2523 (N_2523,N_2316,N_2331);
nand U2524 (N_2524,N_2123,N_2336);
or U2525 (N_2525,N_2251,N_2369);
nor U2526 (N_2526,N_2386,N_2325);
nor U2527 (N_2527,N_2129,N_2198);
or U2528 (N_2528,N_2174,N_2310);
or U2529 (N_2529,N_2152,N_2261);
xor U2530 (N_2530,N_2312,N_2124);
xor U2531 (N_2531,N_2298,N_2185);
nor U2532 (N_2532,N_2330,N_2245);
xor U2533 (N_2533,N_2326,N_2247);
and U2534 (N_2534,N_2297,N_2158);
and U2535 (N_2535,N_2116,N_2335);
nor U2536 (N_2536,N_2364,N_2144);
xnor U2537 (N_2537,N_2204,N_2285);
nor U2538 (N_2538,N_2392,N_2374);
xnor U2539 (N_2539,N_2172,N_2211);
or U2540 (N_2540,N_2125,N_2200);
nand U2541 (N_2541,N_2344,N_2228);
and U2542 (N_2542,N_2249,N_2375);
nor U2543 (N_2543,N_2149,N_2360);
nand U2544 (N_2544,N_2202,N_2300);
nor U2545 (N_2545,N_2378,N_2376);
xnor U2546 (N_2546,N_2169,N_2292);
nand U2547 (N_2547,N_2239,N_2159);
or U2548 (N_2548,N_2216,N_2165);
xnor U2549 (N_2549,N_2270,N_2319);
and U2550 (N_2550,N_2365,N_2391);
nor U2551 (N_2551,N_2367,N_2246);
or U2552 (N_2552,N_2191,N_2131);
and U2553 (N_2553,N_2245,N_2335);
xnor U2554 (N_2554,N_2341,N_2163);
nor U2555 (N_2555,N_2161,N_2373);
nor U2556 (N_2556,N_2344,N_2332);
or U2557 (N_2557,N_2116,N_2174);
nand U2558 (N_2558,N_2213,N_2204);
and U2559 (N_2559,N_2364,N_2207);
and U2560 (N_2560,N_2358,N_2150);
and U2561 (N_2561,N_2233,N_2327);
nand U2562 (N_2562,N_2385,N_2245);
nor U2563 (N_2563,N_2183,N_2155);
and U2564 (N_2564,N_2100,N_2260);
nor U2565 (N_2565,N_2391,N_2256);
nor U2566 (N_2566,N_2204,N_2356);
nor U2567 (N_2567,N_2363,N_2126);
xor U2568 (N_2568,N_2392,N_2191);
nand U2569 (N_2569,N_2306,N_2382);
nor U2570 (N_2570,N_2240,N_2151);
and U2571 (N_2571,N_2129,N_2116);
nor U2572 (N_2572,N_2235,N_2137);
and U2573 (N_2573,N_2231,N_2336);
xnor U2574 (N_2574,N_2234,N_2110);
xor U2575 (N_2575,N_2251,N_2394);
xnor U2576 (N_2576,N_2169,N_2122);
and U2577 (N_2577,N_2328,N_2246);
xor U2578 (N_2578,N_2374,N_2355);
nand U2579 (N_2579,N_2161,N_2374);
nand U2580 (N_2580,N_2277,N_2236);
or U2581 (N_2581,N_2261,N_2385);
and U2582 (N_2582,N_2196,N_2179);
nand U2583 (N_2583,N_2354,N_2341);
and U2584 (N_2584,N_2314,N_2361);
nand U2585 (N_2585,N_2216,N_2241);
or U2586 (N_2586,N_2176,N_2222);
xnor U2587 (N_2587,N_2144,N_2220);
nand U2588 (N_2588,N_2192,N_2372);
and U2589 (N_2589,N_2274,N_2397);
nor U2590 (N_2590,N_2263,N_2192);
or U2591 (N_2591,N_2267,N_2117);
and U2592 (N_2592,N_2215,N_2321);
nand U2593 (N_2593,N_2123,N_2216);
and U2594 (N_2594,N_2371,N_2137);
or U2595 (N_2595,N_2194,N_2189);
nand U2596 (N_2596,N_2174,N_2300);
xor U2597 (N_2597,N_2381,N_2219);
and U2598 (N_2598,N_2253,N_2338);
nor U2599 (N_2599,N_2153,N_2395);
or U2600 (N_2600,N_2383,N_2334);
and U2601 (N_2601,N_2282,N_2383);
and U2602 (N_2602,N_2224,N_2172);
nand U2603 (N_2603,N_2327,N_2166);
nand U2604 (N_2604,N_2146,N_2245);
xor U2605 (N_2605,N_2380,N_2194);
or U2606 (N_2606,N_2333,N_2393);
xor U2607 (N_2607,N_2370,N_2306);
and U2608 (N_2608,N_2279,N_2383);
nor U2609 (N_2609,N_2325,N_2216);
or U2610 (N_2610,N_2181,N_2251);
and U2611 (N_2611,N_2164,N_2263);
nor U2612 (N_2612,N_2201,N_2100);
and U2613 (N_2613,N_2231,N_2377);
nand U2614 (N_2614,N_2343,N_2249);
and U2615 (N_2615,N_2246,N_2186);
nand U2616 (N_2616,N_2309,N_2316);
nand U2617 (N_2617,N_2374,N_2309);
nand U2618 (N_2618,N_2273,N_2157);
nor U2619 (N_2619,N_2389,N_2227);
nor U2620 (N_2620,N_2275,N_2151);
and U2621 (N_2621,N_2134,N_2369);
nand U2622 (N_2622,N_2310,N_2220);
xnor U2623 (N_2623,N_2132,N_2100);
and U2624 (N_2624,N_2226,N_2369);
or U2625 (N_2625,N_2235,N_2152);
nand U2626 (N_2626,N_2363,N_2200);
xnor U2627 (N_2627,N_2103,N_2180);
or U2628 (N_2628,N_2168,N_2243);
nor U2629 (N_2629,N_2221,N_2106);
and U2630 (N_2630,N_2220,N_2268);
nor U2631 (N_2631,N_2331,N_2356);
or U2632 (N_2632,N_2361,N_2163);
xnor U2633 (N_2633,N_2224,N_2335);
and U2634 (N_2634,N_2181,N_2339);
and U2635 (N_2635,N_2248,N_2187);
and U2636 (N_2636,N_2321,N_2281);
nor U2637 (N_2637,N_2253,N_2157);
xor U2638 (N_2638,N_2135,N_2204);
nor U2639 (N_2639,N_2258,N_2377);
or U2640 (N_2640,N_2110,N_2378);
nor U2641 (N_2641,N_2167,N_2230);
xor U2642 (N_2642,N_2231,N_2103);
or U2643 (N_2643,N_2129,N_2183);
xor U2644 (N_2644,N_2328,N_2184);
nand U2645 (N_2645,N_2311,N_2186);
xnor U2646 (N_2646,N_2283,N_2156);
xnor U2647 (N_2647,N_2325,N_2201);
xnor U2648 (N_2648,N_2180,N_2397);
nor U2649 (N_2649,N_2232,N_2122);
and U2650 (N_2650,N_2211,N_2393);
or U2651 (N_2651,N_2323,N_2129);
nand U2652 (N_2652,N_2352,N_2226);
nand U2653 (N_2653,N_2366,N_2111);
nor U2654 (N_2654,N_2386,N_2283);
or U2655 (N_2655,N_2294,N_2208);
nand U2656 (N_2656,N_2316,N_2202);
xnor U2657 (N_2657,N_2124,N_2148);
nor U2658 (N_2658,N_2234,N_2355);
nor U2659 (N_2659,N_2169,N_2393);
nor U2660 (N_2660,N_2178,N_2136);
xnor U2661 (N_2661,N_2253,N_2116);
and U2662 (N_2662,N_2114,N_2174);
and U2663 (N_2663,N_2358,N_2222);
xor U2664 (N_2664,N_2233,N_2268);
and U2665 (N_2665,N_2115,N_2154);
and U2666 (N_2666,N_2350,N_2267);
nand U2667 (N_2667,N_2159,N_2206);
and U2668 (N_2668,N_2142,N_2264);
nor U2669 (N_2669,N_2311,N_2195);
nor U2670 (N_2670,N_2300,N_2341);
or U2671 (N_2671,N_2350,N_2364);
nor U2672 (N_2672,N_2127,N_2114);
and U2673 (N_2673,N_2395,N_2258);
xnor U2674 (N_2674,N_2337,N_2388);
xor U2675 (N_2675,N_2287,N_2235);
and U2676 (N_2676,N_2231,N_2203);
or U2677 (N_2677,N_2175,N_2347);
nor U2678 (N_2678,N_2162,N_2111);
xnor U2679 (N_2679,N_2378,N_2228);
and U2680 (N_2680,N_2208,N_2276);
and U2681 (N_2681,N_2227,N_2156);
and U2682 (N_2682,N_2358,N_2399);
nor U2683 (N_2683,N_2223,N_2337);
nor U2684 (N_2684,N_2399,N_2297);
nand U2685 (N_2685,N_2315,N_2343);
and U2686 (N_2686,N_2301,N_2338);
nor U2687 (N_2687,N_2261,N_2344);
or U2688 (N_2688,N_2126,N_2165);
or U2689 (N_2689,N_2379,N_2110);
and U2690 (N_2690,N_2375,N_2188);
or U2691 (N_2691,N_2103,N_2145);
and U2692 (N_2692,N_2315,N_2194);
and U2693 (N_2693,N_2166,N_2278);
or U2694 (N_2694,N_2175,N_2376);
nor U2695 (N_2695,N_2164,N_2160);
xor U2696 (N_2696,N_2155,N_2127);
xor U2697 (N_2697,N_2112,N_2189);
nand U2698 (N_2698,N_2217,N_2272);
xnor U2699 (N_2699,N_2245,N_2233);
and U2700 (N_2700,N_2501,N_2448);
xor U2701 (N_2701,N_2576,N_2417);
xor U2702 (N_2702,N_2435,N_2480);
and U2703 (N_2703,N_2454,N_2525);
nor U2704 (N_2704,N_2656,N_2545);
or U2705 (N_2705,N_2442,N_2415);
or U2706 (N_2706,N_2542,N_2553);
or U2707 (N_2707,N_2532,N_2594);
nor U2708 (N_2708,N_2482,N_2648);
xnor U2709 (N_2709,N_2627,N_2565);
xnor U2710 (N_2710,N_2593,N_2643);
xnor U2711 (N_2711,N_2632,N_2492);
and U2712 (N_2712,N_2666,N_2430);
nor U2713 (N_2713,N_2628,N_2633);
nor U2714 (N_2714,N_2672,N_2581);
and U2715 (N_2715,N_2403,N_2412);
or U2716 (N_2716,N_2425,N_2572);
nor U2717 (N_2717,N_2625,N_2547);
and U2718 (N_2718,N_2683,N_2597);
nand U2719 (N_2719,N_2690,N_2543);
nor U2720 (N_2720,N_2538,N_2663);
nor U2721 (N_2721,N_2562,N_2526);
and U2722 (N_2722,N_2429,N_2408);
and U2723 (N_2723,N_2590,N_2401);
xnor U2724 (N_2724,N_2588,N_2601);
nor U2725 (N_2725,N_2517,N_2447);
nand U2726 (N_2726,N_2557,N_2661);
xor U2727 (N_2727,N_2537,N_2622);
nand U2728 (N_2728,N_2668,N_2694);
or U2729 (N_2729,N_2436,N_2522);
and U2730 (N_2730,N_2431,N_2418);
nand U2731 (N_2731,N_2437,N_2536);
xnor U2732 (N_2732,N_2696,N_2484);
or U2733 (N_2733,N_2680,N_2469);
nor U2734 (N_2734,N_2520,N_2498);
and U2735 (N_2735,N_2664,N_2607);
and U2736 (N_2736,N_2462,N_2585);
and U2737 (N_2737,N_2410,N_2560);
nand U2738 (N_2738,N_2596,N_2592);
and U2739 (N_2739,N_2695,N_2506);
nand U2740 (N_2740,N_2471,N_2580);
nor U2741 (N_2741,N_2478,N_2516);
nor U2742 (N_2742,N_2479,N_2551);
xnor U2743 (N_2743,N_2684,N_2402);
and U2744 (N_2744,N_2621,N_2600);
xor U2745 (N_2745,N_2400,N_2589);
nand U2746 (N_2746,N_2416,N_2515);
or U2747 (N_2747,N_2449,N_2455);
or U2748 (N_2748,N_2534,N_2645);
or U2749 (N_2749,N_2639,N_2495);
nand U2750 (N_2750,N_2634,N_2640);
nand U2751 (N_2751,N_2660,N_2673);
and U2752 (N_2752,N_2598,N_2667);
xor U2753 (N_2753,N_2421,N_2438);
nor U2754 (N_2754,N_2508,N_2411);
nor U2755 (N_2755,N_2599,N_2468);
xnor U2756 (N_2756,N_2630,N_2563);
nor U2757 (N_2757,N_2422,N_2567);
xnor U2758 (N_2758,N_2444,N_2615);
nor U2759 (N_2759,N_2552,N_2616);
xor U2760 (N_2760,N_2647,N_2513);
or U2761 (N_2761,N_2612,N_2671);
and U2762 (N_2762,N_2574,N_2496);
and U2763 (N_2763,N_2638,N_2414);
nand U2764 (N_2764,N_2531,N_2649);
and U2765 (N_2765,N_2461,N_2626);
or U2766 (N_2766,N_2558,N_2587);
xnor U2767 (N_2767,N_2657,N_2419);
nand U2768 (N_2768,N_2646,N_2573);
nor U2769 (N_2769,N_2655,N_2698);
xnor U2770 (N_2770,N_2529,N_2406);
or U2771 (N_2771,N_2618,N_2604);
nor U2772 (N_2772,N_2533,N_2477);
and U2773 (N_2773,N_2569,N_2682);
xnor U2774 (N_2774,N_2608,N_2650);
xnor U2775 (N_2775,N_2564,N_2504);
nor U2776 (N_2776,N_2609,N_2485);
or U2777 (N_2777,N_2464,N_2662);
nand U2778 (N_2778,N_2474,N_2404);
nor U2779 (N_2779,N_2554,N_2434);
or U2780 (N_2780,N_2490,N_2606);
and U2781 (N_2781,N_2584,N_2577);
or U2782 (N_2782,N_2610,N_2503);
xor U2783 (N_2783,N_2511,N_2505);
xnor U2784 (N_2784,N_2678,N_2441);
xor U2785 (N_2785,N_2652,N_2472);
and U2786 (N_2786,N_2654,N_2641);
or U2787 (N_2787,N_2463,N_2617);
and U2788 (N_2788,N_2460,N_2453);
xnor U2789 (N_2789,N_2540,N_2693);
nand U2790 (N_2790,N_2409,N_2475);
or U2791 (N_2791,N_2443,N_2575);
or U2792 (N_2792,N_2413,N_2681);
nor U2793 (N_2793,N_2691,N_2595);
nor U2794 (N_2794,N_2544,N_2549);
or U2795 (N_2795,N_2502,N_2424);
nor U2796 (N_2796,N_2602,N_2530);
nand U2797 (N_2797,N_2687,N_2620);
nand U2798 (N_2798,N_2689,N_2611);
nand U2799 (N_2799,N_2445,N_2458);
nor U2800 (N_2800,N_2582,N_2420);
and U2801 (N_2801,N_2405,N_2583);
xor U2802 (N_2802,N_2603,N_2619);
and U2803 (N_2803,N_2570,N_2555);
and U2804 (N_2804,N_2457,N_2676);
xor U2805 (N_2805,N_2499,N_2512);
nand U2806 (N_2806,N_2519,N_2561);
nor U2807 (N_2807,N_2423,N_2635);
nor U2808 (N_2808,N_2550,N_2473);
or U2809 (N_2809,N_2566,N_2653);
nor U2810 (N_2810,N_2446,N_2644);
nor U2811 (N_2811,N_2631,N_2579);
nor U2812 (N_2812,N_2636,N_2497);
nor U2813 (N_2813,N_2440,N_2528);
or U2814 (N_2814,N_2428,N_2613);
and U2815 (N_2815,N_2486,N_2679);
or U2816 (N_2816,N_2546,N_2688);
xor U2817 (N_2817,N_2491,N_2675);
xor U2818 (N_2818,N_2407,N_2439);
xnor U2819 (N_2819,N_2697,N_2623);
and U2820 (N_2820,N_2665,N_2489);
nand U2821 (N_2821,N_2692,N_2481);
xor U2822 (N_2822,N_2451,N_2433);
and U2823 (N_2823,N_2674,N_2614);
and U2824 (N_2824,N_2642,N_2629);
xor U2825 (N_2825,N_2432,N_2427);
and U2826 (N_2826,N_2677,N_2637);
nand U2827 (N_2827,N_2456,N_2670);
or U2828 (N_2828,N_2493,N_2658);
nand U2829 (N_2829,N_2571,N_2586);
xor U2830 (N_2830,N_2548,N_2527);
nand U2831 (N_2831,N_2459,N_2488);
nand U2832 (N_2832,N_2578,N_2500);
and U2833 (N_2833,N_2605,N_2466);
or U2834 (N_2834,N_2659,N_2494);
xor U2835 (N_2835,N_2426,N_2535);
and U2836 (N_2836,N_2452,N_2539);
and U2837 (N_2837,N_2559,N_2524);
or U2838 (N_2838,N_2624,N_2483);
nor U2839 (N_2839,N_2686,N_2465);
xnor U2840 (N_2840,N_2669,N_2470);
nand U2841 (N_2841,N_2514,N_2521);
and U2842 (N_2842,N_2541,N_2450);
nand U2843 (N_2843,N_2523,N_2699);
or U2844 (N_2844,N_2509,N_2476);
or U2845 (N_2845,N_2507,N_2510);
or U2846 (N_2846,N_2487,N_2467);
and U2847 (N_2847,N_2568,N_2685);
and U2848 (N_2848,N_2591,N_2518);
xor U2849 (N_2849,N_2556,N_2651);
and U2850 (N_2850,N_2415,N_2419);
or U2851 (N_2851,N_2499,N_2428);
nor U2852 (N_2852,N_2481,N_2614);
or U2853 (N_2853,N_2403,N_2535);
or U2854 (N_2854,N_2645,N_2634);
nand U2855 (N_2855,N_2563,N_2556);
xnor U2856 (N_2856,N_2420,N_2483);
nor U2857 (N_2857,N_2596,N_2405);
nor U2858 (N_2858,N_2507,N_2413);
and U2859 (N_2859,N_2426,N_2568);
and U2860 (N_2860,N_2629,N_2592);
nand U2861 (N_2861,N_2596,N_2504);
or U2862 (N_2862,N_2626,N_2684);
nor U2863 (N_2863,N_2591,N_2524);
or U2864 (N_2864,N_2593,N_2687);
xnor U2865 (N_2865,N_2657,N_2543);
or U2866 (N_2866,N_2674,N_2632);
xor U2867 (N_2867,N_2599,N_2655);
and U2868 (N_2868,N_2647,N_2671);
nor U2869 (N_2869,N_2408,N_2409);
nor U2870 (N_2870,N_2437,N_2697);
xnor U2871 (N_2871,N_2425,N_2506);
nor U2872 (N_2872,N_2668,N_2465);
nand U2873 (N_2873,N_2563,N_2548);
xnor U2874 (N_2874,N_2436,N_2496);
and U2875 (N_2875,N_2643,N_2424);
nor U2876 (N_2876,N_2591,N_2415);
xnor U2877 (N_2877,N_2417,N_2650);
and U2878 (N_2878,N_2430,N_2687);
xnor U2879 (N_2879,N_2609,N_2552);
xnor U2880 (N_2880,N_2579,N_2657);
xor U2881 (N_2881,N_2464,N_2577);
xnor U2882 (N_2882,N_2465,N_2400);
xor U2883 (N_2883,N_2442,N_2554);
or U2884 (N_2884,N_2440,N_2534);
nand U2885 (N_2885,N_2571,N_2467);
or U2886 (N_2886,N_2430,N_2599);
or U2887 (N_2887,N_2612,N_2606);
or U2888 (N_2888,N_2699,N_2589);
xor U2889 (N_2889,N_2458,N_2422);
or U2890 (N_2890,N_2502,N_2699);
xor U2891 (N_2891,N_2437,N_2554);
nor U2892 (N_2892,N_2606,N_2419);
or U2893 (N_2893,N_2531,N_2462);
or U2894 (N_2894,N_2688,N_2658);
nor U2895 (N_2895,N_2638,N_2627);
or U2896 (N_2896,N_2456,N_2667);
or U2897 (N_2897,N_2418,N_2593);
or U2898 (N_2898,N_2646,N_2603);
nor U2899 (N_2899,N_2536,N_2544);
nand U2900 (N_2900,N_2690,N_2481);
xnor U2901 (N_2901,N_2470,N_2479);
xnor U2902 (N_2902,N_2567,N_2511);
nand U2903 (N_2903,N_2512,N_2460);
or U2904 (N_2904,N_2622,N_2572);
nor U2905 (N_2905,N_2526,N_2502);
or U2906 (N_2906,N_2607,N_2636);
nand U2907 (N_2907,N_2429,N_2435);
xnor U2908 (N_2908,N_2410,N_2670);
xnor U2909 (N_2909,N_2431,N_2643);
xnor U2910 (N_2910,N_2546,N_2442);
nor U2911 (N_2911,N_2685,N_2417);
xnor U2912 (N_2912,N_2419,N_2570);
or U2913 (N_2913,N_2647,N_2576);
nor U2914 (N_2914,N_2676,N_2513);
nor U2915 (N_2915,N_2524,N_2644);
xnor U2916 (N_2916,N_2455,N_2624);
and U2917 (N_2917,N_2542,N_2516);
nor U2918 (N_2918,N_2675,N_2517);
xor U2919 (N_2919,N_2549,N_2680);
xnor U2920 (N_2920,N_2428,N_2543);
and U2921 (N_2921,N_2691,N_2511);
and U2922 (N_2922,N_2504,N_2478);
or U2923 (N_2923,N_2686,N_2485);
or U2924 (N_2924,N_2644,N_2637);
nand U2925 (N_2925,N_2520,N_2696);
xor U2926 (N_2926,N_2690,N_2408);
xor U2927 (N_2927,N_2438,N_2454);
xor U2928 (N_2928,N_2465,N_2682);
nand U2929 (N_2929,N_2674,N_2460);
or U2930 (N_2930,N_2439,N_2644);
or U2931 (N_2931,N_2680,N_2492);
xnor U2932 (N_2932,N_2413,N_2528);
or U2933 (N_2933,N_2488,N_2553);
and U2934 (N_2934,N_2484,N_2653);
or U2935 (N_2935,N_2624,N_2558);
nand U2936 (N_2936,N_2532,N_2577);
and U2937 (N_2937,N_2550,N_2600);
xor U2938 (N_2938,N_2408,N_2419);
xor U2939 (N_2939,N_2560,N_2654);
or U2940 (N_2940,N_2535,N_2618);
nor U2941 (N_2941,N_2607,N_2670);
nand U2942 (N_2942,N_2454,N_2582);
or U2943 (N_2943,N_2462,N_2667);
and U2944 (N_2944,N_2500,N_2660);
xnor U2945 (N_2945,N_2516,N_2628);
nor U2946 (N_2946,N_2440,N_2543);
nor U2947 (N_2947,N_2686,N_2682);
nand U2948 (N_2948,N_2533,N_2469);
and U2949 (N_2949,N_2668,N_2538);
nand U2950 (N_2950,N_2534,N_2544);
nand U2951 (N_2951,N_2472,N_2624);
and U2952 (N_2952,N_2496,N_2633);
nor U2953 (N_2953,N_2687,N_2629);
nor U2954 (N_2954,N_2605,N_2517);
and U2955 (N_2955,N_2640,N_2506);
and U2956 (N_2956,N_2634,N_2545);
or U2957 (N_2957,N_2431,N_2534);
xnor U2958 (N_2958,N_2410,N_2485);
xor U2959 (N_2959,N_2683,N_2437);
nor U2960 (N_2960,N_2416,N_2599);
or U2961 (N_2961,N_2528,N_2636);
nand U2962 (N_2962,N_2696,N_2599);
or U2963 (N_2963,N_2639,N_2689);
nor U2964 (N_2964,N_2518,N_2455);
nor U2965 (N_2965,N_2436,N_2490);
nand U2966 (N_2966,N_2525,N_2466);
nand U2967 (N_2967,N_2625,N_2541);
nor U2968 (N_2968,N_2653,N_2458);
nand U2969 (N_2969,N_2611,N_2501);
or U2970 (N_2970,N_2503,N_2689);
nor U2971 (N_2971,N_2685,N_2476);
nand U2972 (N_2972,N_2567,N_2435);
nand U2973 (N_2973,N_2405,N_2607);
nand U2974 (N_2974,N_2409,N_2484);
nand U2975 (N_2975,N_2577,N_2496);
nand U2976 (N_2976,N_2549,N_2577);
nor U2977 (N_2977,N_2598,N_2488);
or U2978 (N_2978,N_2625,N_2465);
nand U2979 (N_2979,N_2533,N_2646);
xor U2980 (N_2980,N_2545,N_2444);
nand U2981 (N_2981,N_2527,N_2659);
nor U2982 (N_2982,N_2500,N_2473);
or U2983 (N_2983,N_2687,N_2677);
xnor U2984 (N_2984,N_2689,N_2599);
nand U2985 (N_2985,N_2667,N_2480);
nand U2986 (N_2986,N_2490,N_2444);
xor U2987 (N_2987,N_2508,N_2419);
xor U2988 (N_2988,N_2697,N_2432);
and U2989 (N_2989,N_2621,N_2690);
nand U2990 (N_2990,N_2515,N_2495);
nor U2991 (N_2991,N_2549,N_2547);
and U2992 (N_2992,N_2477,N_2440);
nand U2993 (N_2993,N_2697,N_2501);
and U2994 (N_2994,N_2434,N_2542);
xor U2995 (N_2995,N_2502,N_2648);
and U2996 (N_2996,N_2656,N_2406);
xnor U2997 (N_2997,N_2679,N_2474);
or U2998 (N_2998,N_2618,N_2685);
or U2999 (N_2999,N_2410,N_2525);
and U3000 (N_3000,N_2973,N_2813);
or U3001 (N_3001,N_2822,N_2756);
nor U3002 (N_3002,N_2781,N_2774);
nor U3003 (N_3003,N_2759,N_2923);
or U3004 (N_3004,N_2811,N_2745);
xor U3005 (N_3005,N_2996,N_2993);
nor U3006 (N_3006,N_2875,N_2969);
and U3007 (N_3007,N_2730,N_2736);
and U3008 (N_3008,N_2825,N_2995);
xnor U3009 (N_3009,N_2773,N_2729);
or U3010 (N_3010,N_2937,N_2799);
xor U3011 (N_3011,N_2843,N_2830);
and U3012 (N_3012,N_2861,N_2944);
and U3013 (N_3013,N_2705,N_2960);
xor U3014 (N_3014,N_2867,N_2725);
xor U3015 (N_3015,N_2852,N_2785);
xnor U3016 (N_3016,N_2789,N_2855);
nor U3017 (N_3017,N_2800,N_2719);
nor U3018 (N_3018,N_2753,N_2744);
nand U3019 (N_3019,N_2915,N_2802);
xnor U3020 (N_3020,N_2888,N_2771);
nand U3021 (N_3021,N_2887,N_2720);
nand U3022 (N_3022,N_2893,N_2769);
xnor U3023 (N_3023,N_2770,N_2897);
xor U3024 (N_3024,N_2877,N_2924);
and U3025 (N_3025,N_2701,N_2979);
or U3026 (N_3026,N_2921,N_2732);
xor U3027 (N_3027,N_2863,N_2910);
or U3028 (N_3028,N_2872,N_2903);
nand U3029 (N_3029,N_2776,N_2715);
nor U3030 (N_3030,N_2871,N_2810);
xnor U3031 (N_3031,N_2900,N_2765);
nor U3032 (N_3032,N_2734,N_2768);
nand U3033 (N_3033,N_2832,N_2763);
and U3034 (N_3034,N_2869,N_2842);
and U3035 (N_3035,N_2901,N_2741);
and U3036 (N_3036,N_2928,N_2831);
xnor U3037 (N_3037,N_2777,N_2812);
and U3038 (N_3038,N_2828,N_2794);
or U3039 (N_3039,N_2807,N_2735);
and U3040 (N_3040,N_2837,N_2961);
xnor U3041 (N_3041,N_2747,N_2870);
nand U3042 (N_3042,N_2801,N_2762);
and U3043 (N_3043,N_2882,N_2788);
nand U3044 (N_3044,N_2964,N_2833);
and U3045 (N_3045,N_2819,N_2751);
or U3046 (N_3046,N_2755,N_2970);
nor U3047 (N_3047,N_2845,N_2879);
xor U3048 (N_3048,N_2880,N_2949);
nand U3049 (N_3049,N_2959,N_2980);
nor U3050 (N_3050,N_2815,N_2999);
and U3051 (N_3051,N_2823,N_2991);
xnor U3052 (N_3052,N_2841,N_2968);
or U3053 (N_3053,N_2906,N_2943);
nand U3054 (N_3054,N_2998,N_2975);
nor U3055 (N_3055,N_2983,N_2752);
and U3056 (N_3056,N_2866,N_2817);
and U3057 (N_3057,N_2723,N_2862);
nor U3058 (N_3058,N_2787,N_2898);
nor U3059 (N_3059,N_2894,N_2972);
nand U3060 (N_3060,N_2935,N_2782);
nor U3061 (N_3061,N_2865,N_2733);
nand U3062 (N_3062,N_2742,N_2764);
xor U3063 (N_3063,N_2724,N_2976);
xnor U3064 (N_3064,N_2748,N_2726);
and U3065 (N_3065,N_2707,N_2708);
and U3066 (N_3066,N_2848,N_2954);
xnor U3067 (N_3067,N_2876,N_2904);
or U3068 (N_3068,N_2712,N_2925);
and U3069 (N_3069,N_2760,N_2709);
xor U3070 (N_3070,N_2982,N_2739);
or U3071 (N_3071,N_2786,N_2849);
or U3072 (N_3072,N_2761,N_2783);
or U3073 (N_3073,N_2766,N_2891);
nand U3074 (N_3074,N_2728,N_2803);
and U3075 (N_3075,N_2918,N_2883);
nand U3076 (N_3076,N_2718,N_2860);
nand U3077 (N_3077,N_2881,N_2884);
nand U3078 (N_3078,N_2957,N_2919);
and U3079 (N_3079,N_2847,N_2962);
and U3080 (N_3080,N_2749,N_2941);
nor U3081 (N_3081,N_2814,N_2780);
nor U3082 (N_3082,N_2953,N_2933);
xnor U3083 (N_3083,N_2965,N_2738);
nor U3084 (N_3084,N_2985,N_2994);
xnor U3085 (N_3085,N_2727,N_2911);
nor U3086 (N_3086,N_2927,N_2790);
nor U3087 (N_3087,N_2938,N_2805);
nand U3088 (N_3088,N_2859,N_2950);
nor U3089 (N_3089,N_2806,N_2704);
xnor U3090 (N_3090,N_2834,N_2779);
and U3091 (N_3091,N_2988,N_2722);
nand U3092 (N_3092,N_2955,N_2710);
or U3093 (N_3093,N_2912,N_2854);
xor U3094 (N_3094,N_2716,N_2700);
xnor U3095 (N_3095,N_2936,N_2791);
nor U3096 (N_3096,N_2703,N_2914);
xor U3097 (N_3097,N_2731,N_2850);
xor U3098 (N_3098,N_2934,N_2892);
and U3099 (N_3099,N_2987,N_2907);
and U3100 (N_3100,N_2913,N_2793);
or U3101 (N_3101,N_2940,N_2835);
nor U3102 (N_3102,N_2885,N_2839);
or U3103 (N_3103,N_2902,N_2948);
nand U3104 (N_3104,N_2824,N_2856);
nand U3105 (N_3105,N_2990,N_2743);
or U3106 (N_3106,N_2796,N_2804);
nor U3107 (N_3107,N_2816,N_2952);
xor U3108 (N_3108,N_2963,N_2827);
nor U3109 (N_3109,N_2818,N_2890);
and U3110 (N_3110,N_2858,N_2997);
or U3111 (N_3111,N_2714,N_2853);
nor U3112 (N_3112,N_2951,N_2702);
or U3113 (N_3113,N_2945,N_2706);
and U3114 (N_3114,N_2851,N_2798);
nand U3115 (N_3115,N_2746,N_2864);
nand U3116 (N_3116,N_2721,N_2820);
nand U3117 (N_3117,N_2838,N_2922);
or U3118 (N_3118,N_2896,N_2947);
nand U3119 (N_3119,N_2920,N_2757);
nor U3120 (N_3120,N_2977,N_2930);
xor U3121 (N_3121,N_2737,N_2868);
and U3122 (N_3122,N_2795,N_2956);
and U3123 (N_3123,N_2784,N_2857);
xnor U3124 (N_3124,N_2966,N_2844);
nand U3125 (N_3125,N_2958,N_2984);
xor U3126 (N_3126,N_2758,N_2740);
nand U3127 (N_3127,N_2772,N_2836);
and U3128 (N_3128,N_2886,N_2778);
and U3129 (N_3129,N_2873,N_2971);
or U3130 (N_3130,N_2713,N_2917);
xnor U3131 (N_3131,N_2797,N_2899);
nand U3132 (N_3132,N_2978,N_2874);
xor U3133 (N_3133,N_2840,N_2767);
and U3134 (N_3134,N_2792,N_2750);
nand U3135 (N_3135,N_2826,N_2926);
or U3136 (N_3136,N_2754,N_2942);
xor U3137 (N_3137,N_2895,N_2808);
nor U3138 (N_3138,N_2929,N_2878);
and U3139 (N_3139,N_2889,N_2908);
and U3140 (N_3140,N_2916,N_2846);
nor U3141 (N_3141,N_2909,N_2939);
xnor U3142 (N_3142,N_2974,N_2717);
nand U3143 (N_3143,N_2775,N_2989);
xnor U3144 (N_3144,N_2905,N_2946);
and U3145 (N_3145,N_2711,N_2821);
and U3146 (N_3146,N_2967,N_2981);
and U3147 (N_3147,N_2992,N_2986);
nand U3148 (N_3148,N_2931,N_2809);
xor U3149 (N_3149,N_2932,N_2829);
and U3150 (N_3150,N_2933,N_2796);
and U3151 (N_3151,N_2913,N_2786);
nor U3152 (N_3152,N_2997,N_2716);
or U3153 (N_3153,N_2926,N_2931);
xor U3154 (N_3154,N_2702,N_2909);
nor U3155 (N_3155,N_2781,N_2832);
xor U3156 (N_3156,N_2825,N_2920);
or U3157 (N_3157,N_2773,N_2859);
nor U3158 (N_3158,N_2764,N_2767);
or U3159 (N_3159,N_2749,N_2996);
or U3160 (N_3160,N_2929,N_2770);
or U3161 (N_3161,N_2888,N_2901);
xor U3162 (N_3162,N_2861,N_2978);
xor U3163 (N_3163,N_2886,N_2782);
and U3164 (N_3164,N_2703,N_2829);
nor U3165 (N_3165,N_2735,N_2791);
nor U3166 (N_3166,N_2764,N_2711);
and U3167 (N_3167,N_2960,N_2797);
nor U3168 (N_3168,N_2821,N_2929);
xor U3169 (N_3169,N_2752,N_2828);
nand U3170 (N_3170,N_2767,N_2736);
xnor U3171 (N_3171,N_2934,N_2845);
xor U3172 (N_3172,N_2811,N_2714);
nor U3173 (N_3173,N_2956,N_2793);
nand U3174 (N_3174,N_2745,N_2765);
and U3175 (N_3175,N_2940,N_2937);
nor U3176 (N_3176,N_2926,N_2994);
nor U3177 (N_3177,N_2855,N_2861);
nand U3178 (N_3178,N_2995,N_2773);
nand U3179 (N_3179,N_2731,N_2751);
and U3180 (N_3180,N_2738,N_2821);
and U3181 (N_3181,N_2968,N_2732);
xnor U3182 (N_3182,N_2891,N_2937);
or U3183 (N_3183,N_2839,N_2752);
nand U3184 (N_3184,N_2838,N_2916);
xnor U3185 (N_3185,N_2900,N_2703);
xnor U3186 (N_3186,N_2978,N_2948);
nor U3187 (N_3187,N_2864,N_2825);
xnor U3188 (N_3188,N_2768,N_2793);
xor U3189 (N_3189,N_2899,N_2811);
and U3190 (N_3190,N_2938,N_2708);
or U3191 (N_3191,N_2867,N_2787);
nand U3192 (N_3192,N_2834,N_2839);
nand U3193 (N_3193,N_2852,N_2801);
or U3194 (N_3194,N_2837,N_2719);
and U3195 (N_3195,N_2881,N_2797);
nor U3196 (N_3196,N_2774,N_2868);
nor U3197 (N_3197,N_2742,N_2913);
xor U3198 (N_3198,N_2882,N_2971);
or U3199 (N_3199,N_2838,N_2800);
nand U3200 (N_3200,N_2705,N_2970);
or U3201 (N_3201,N_2945,N_2709);
nor U3202 (N_3202,N_2707,N_2889);
or U3203 (N_3203,N_2728,N_2859);
or U3204 (N_3204,N_2772,N_2829);
xor U3205 (N_3205,N_2734,N_2927);
nor U3206 (N_3206,N_2998,N_2932);
nand U3207 (N_3207,N_2720,N_2833);
xor U3208 (N_3208,N_2882,N_2835);
and U3209 (N_3209,N_2830,N_2917);
xor U3210 (N_3210,N_2743,N_2873);
xor U3211 (N_3211,N_2920,N_2775);
nand U3212 (N_3212,N_2861,N_2768);
xor U3213 (N_3213,N_2942,N_2915);
nand U3214 (N_3214,N_2925,N_2704);
nor U3215 (N_3215,N_2827,N_2975);
nand U3216 (N_3216,N_2995,N_2938);
or U3217 (N_3217,N_2715,N_2712);
or U3218 (N_3218,N_2750,N_2772);
xor U3219 (N_3219,N_2761,N_2885);
nor U3220 (N_3220,N_2833,N_2857);
and U3221 (N_3221,N_2808,N_2992);
xor U3222 (N_3222,N_2802,N_2726);
and U3223 (N_3223,N_2990,N_2808);
and U3224 (N_3224,N_2799,N_2981);
or U3225 (N_3225,N_2703,N_2873);
xor U3226 (N_3226,N_2771,N_2896);
and U3227 (N_3227,N_2836,N_2720);
nand U3228 (N_3228,N_2846,N_2877);
xnor U3229 (N_3229,N_2832,N_2944);
nor U3230 (N_3230,N_2825,N_2782);
nor U3231 (N_3231,N_2871,N_2791);
or U3232 (N_3232,N_2974,N_2889);
nand U3233 (N_3233,N_2763,N_2917);
xor U3234 (N_3234,N_2924,N_2825);
xor U3235 (N_3235,N_2746,N_2961);
and U3236 (N_3236,N_2756,N_2860);
nand U3237 (N_3237,N_2821,N_2842);
xnor U3238 (N_3238,N_2829,N_2940);
and U3239 (N_3239,N_2944,N_2702);
and U3240 (N_3240,N_2824,N_2836);
nor U3241 (N_3241,N_2874,N_2983);
nand U3242 (N_3242,N_2999,N_2708);
or U3243 (N_3243,N_2851,N_2864);
and U3244 (N_3244,N_2903,N_2883);
and U3245 (N_3245,N_2959,N_2978);
nand U3246 (N_3246,N_2930,N_2934);
and U3247 (N_3247,N_2915,N_2856);
and U3248 (N_3248,N_2985,N_2780);
or U3249 (N_3249,N_2968,N_2755);
nand U3250 (N_3250,N_2993,N_2856);
or U3251 (N_3251,N_2868,N_2842);
xor U3252 (N_3252,N_2953,N_2711);
and U3253 (N_3253,N_2842,N_2796);
nand U3254 (N_3254,N_2800,N_2730);
and U3255 (N_3255,N_2974,N_2978);
nor U3256 (N_3256,N_2824,N_2966);
nor U3257 (N_3257,N_2847,N_2997);
nand U3258 (N_3258,N_2770,N_2729);
nor U3259 (N_3259,N_2996,N_2800);
nand U3260 (N_3260,N_2891,N_2791);
nor U3261 (N_3261,N_2720,N_2991);
nand U3262 (N_3262,N_2904,N_2725);
or U3263 (N_3263,N_2765,N_2971);
or U3264 (N_3264,N_2832,N_2744);
and U3265 (N_3265,N_2872,N_2884);
or U3266 (N_3266,N_2712,N_2741);
xor U3267 (N_3267,N_2864,N_2734);
or U3268 (N_3268,N_2969,N_2714);
and U3269 (N_3269,N_2755,N_2706);
nand U3270 (N_3270,N_2770,N_2805);
nor U3271 (N_3271,N_2895,N_2897);
xor U3272 (N_3272,N_2898,N_2750);
nor U3273 (N_3273,N_2949,N_2787);
and U3274 (N_3274,N_2877,N_2765);
and U3275 (N_3275,N_2711,N_2979);
and U3276 (N_3276,N_2901,N_2936);
nand U3277 (N_3277,N_2891,N_2850);
nor U3278 (N_3278,N_2748,N_2936);
or U3279 (N_3279,N_2710,N_2816);
xor U3280 (N_3280,N_2781,N_2903);
xnor U3281 (N_3281,N_2756,N_2819);
nand U3282 (N_3282,N_2769,N_2899);
or U3283 (N_3283,N_2973,N_2933);
nand U3284 (N_3284,N_2968,N_2762);
nor U3285 (N_3285,N_2776,N_2890);
or U3286 (N_3286,N_2878,N_2911);
xnor U3287 (N_3287,N_2929,N_2948);
and U3288 (N_3288,N_2939,N_2788);
nand U3289 (N_3289,N_2849,N_2962);
xnor U3290 (N_3290,N_2801,N_2827);
and U3291 (N_3291,N_2751,N_2775);
nor U3292 (N_3292,N_2740,N_2725);
xor U3293 (N_3293,N_2857,N_2964);
nand U3294 (N_3294,N_2931,N_2824);
or U3295 (N_3295,N_2870,N_2787);
or U3296 (N_3296,N_2799,N_2994);
and U3297 (N_3297,N_2789,N_2818);
nor U3298 (N_3298,N_2842,N_2748);
nand U3299 (N_3299,N_2741,N_2976);
nand U3300 (N_3300,N_3123,N_3035);
nor U3301 (N_3301,N_3011,N_3218);
or U3302 (N_3302,N_3052,N_3226);
nor U3303 (N_3303,N_3041,N_3100);
nor U3304 (N_3304,N_3213,N_3276);
xor U3305 (N_3305,N_3282,N_3222);
nor U3306 (N_3306,N_3275,N_3018);
nand U3307 (N_3307,N_3074,N_3228);
nand U3308 (N_3308,N_3053,N_3201);
and U3309 (N_3309,N_3235,N_3159);
nor U3310 (N_3310,N_3081,N_3132);
or U3311 (N_3311,N_3192,N_3281);
or U3312 (N_3312,N_3188,N_3167);
nand U3313 (N_3313,N_3273,N_3238);
nand U3314 (N_3314,N_3070,N_3279);
nand U3315 (N_3315,N_3198,N_3102);
nand U3316 (N_3316,N_3203,N_3060);
and U3317 (N_3317,N_3250,N_3183);
or U3318 (N_3318,N_3189,N_3193);
nor U3319 (N_3319,N_3025,N_3175);
nor U3320 (N_3320,N_3297,N_3269);
or U3321 (N_3321,N_3169,N_3085);
xor U3322 (N_3322,N_3015,N_3013);
nand U3323 (N_3323,N_3099,N_3073);
xnor U3324 (N_3324,N_3002,N_3014);
nand U3325 (N_3325,N_3056,N_3178);
xor U3326 (N_3326,N_3215,N_3161);
or U3327 (N_3327,N_3146,N_3140);
or U3328 (N_3328,N_3150,N_3045);
and U3329 (N_3329,N_3229,N_3225);
or U3330 (N_3330,N_3144,N_3107);
xnor U3331 (N_3331,N_3176,N_3034);
xnor U3332 (N_3332,N_3026,N_3130);
and U3333 (N_3333,N_3143,N_3171);
and U3334 (N_3334,N_3135,N_3019);
nand U3335 (N_3335,N_3039,N_3072);
nand U3336 (N_3336,N_3098,N_3094);
or U3337 (N_3337,N_3048,N_3077);
nand U3338 (N_3338,N_3265,N_3010);
xnor U3339 (N_3339,N_3111,N_3196);
nand U3340 (N_3340,N_3017,N_3118);
and U3341 (N_3341,N_3214,N_3231);
or U3342 (N_3342,N_3202,N_3075);
xnor U3343 (N_3343,N_3270,N_3125);
and U3344 (N_3344,N_3272,N_3148);
xnor U3345 (N_3345,N_3028,N_3036);
and U3346 (N_3346,N_3126,N_3078);
nor U3347 (N_3347,N_3103,N_3106);
xnor U3348 (N_3348,N_3001,N_3037);
and U3349 (N_3349,N_3173,N_3128);
or U3350 (N_3350,N_3061,N_3115);
xor U3351 (N_3351,N_3021,N_3095);
nand U3352 (N_3352,N_3101,N_3223);
and U3353 (N_3353,N_3032,N_3168);
nand U3354 (N_3354,N_3137,N_3117);
nand U3355 (N_3355,N_3283,N_3163);
nand U3356 (N_3356,N_3058,N_3289);
and U3357 (N_3357,N_3108,N_3142);
nor U3358 (N_3358,N_3033,N_3112);
xor U3359 (N_3359,N_3155,N_3280);
xnor U3360 (N_3360,N_3113,N_3267);
or U3361 (N_3361,N_3199,N_3274);
and U3362 (N_3362,N_3005,N_3129);
xnor U3363 (N_3363,N_3063,N_3187);
nand U3364 (N_3364,N_3258,N_3029);
or U3365 (N_3365,N_3181,N_3047);
nor U3366 (N_3366,N_3295,N_3154);
or U3367 (N_3367,N_3030,N_3271);
or U3368 (N_3368,N_3162,N_3240);
nand U3369 (N_3369,N_3000,N_3241);
xor U3370 (N_3370,N_3285,N_3197);
nor U3371 (N_3371,N_3204,N_3200);
xor U3372 (N_3372,N_3180,N_3262);
and U3373 (N_3373,N_3170,N_3165);
nor U3374 (N_3374,N_3207,N_3206);
xor U3375 (N_3375,N_3082,N_3046);
xor U3376 (N_3376,N_3127,N_3020);
or U3377 (N_3377,N_3065,N_3191);
nor U3378 (N_3378,N_3293,N_3022);
and U3379 (N_3379,N_3217,N_3221);
nand U3380 (N_3380,N_3209,N_3208);
xor U3381 (N_3381,N_3261,N_3114);
xor U3382 (N_3382,N_3055,N_3008);
nor U3383 (N_3383,N_3012,N_3237);
nand U3384 (N_3384,N_3090,N_3219);
and U3385 (N_3385,N_3027,N_3230);
xnor U3386 (N_3386,N_3043,N_3184);
nor U3387 (N_3387,N_3212,N_3179);
xor U3388 (N_3388,N_3244,N_3044);
xor U3389 (N_3389,N_3151,N_3120);
and U3390 (N_3390,N_3245,N_3079);
and U3391 (N_3391,N_3249,N_3003);
and U3392 (N_3392,N_3185,N_3054);
and U3393 (N_3393,N_3186,N_3080);
nand U3394 (N_3394,N_3139,N_3284);
or U3395 (N_3395,N_3211,N_3253);
and U3396 (N_3396,N_3158,N_3177);
or U3397 (N_3397,N_3290,N_3243);
nor U3398 (N_3398,N_3156,N_3069);
or U3399 (N_3399,N_3134,N_3097);
xor U3400 (N_3400,N_3104,N_3174);
and U3401 (N_3401,N_3109,N_3057);
nor U3402 (N_3402,N_3210,N_3268);
or U3403 (N_3403,N_3145,N_3224);
nand U3404 (N_3404,N_3004,N_3236);
nand U3405 (N_3405,N_3216,N_3166);
nor U3406 (N_3406,N_3278,N_3255);
nor U3407 (N_3407,N_3149,N_3248);
xnor U3408 (N_3408,N_3089,N_3259);
nor U3409 (N_3409,N_3182,N_3092);
xor U3410 (N_3410,N_3131,N_3016);
nand U3411 (N_3411,N_3291,N_3007);
nand U3412 (N_3412,N_3059,N_3049);
nand U3413 (N_3413,N_3110,N_3287);
nor U3414 (N_3414,N_3286,N_3288);
nand U3415 (N_3415,N_3105,N_3122);
xnor U3416 (N_3416,N_3084,N_3299);
or U3417 (N_3417,N_3093,N_3292);
or U3418 (N_3418,N_3232,N_3009);
and U3419 (N_3419,N_3062,N_3083);
and U3420 (N_3420,N_3076,N_3233);
nor U3421 (N_3421,N_3042,N_3087);
nor U3422 (N_3422,N_3242,N_3068);
xnor U3423 (N_3423,N_3067,N_3160);
xor U3424 (N_3424,N_3066,N_3164);
xor U3425 (N_3425,N_3121,N_3194);
and U3426 (N_3426,N_3006,N_3172);
nor U3427 (N_3427,N_3116,N_3050);
or U3428 (N_3428,N_3257,N_3091);
xor U3429 (N_3429,N_3031,N_3071);
and U3430 (N_3430,N_3152,N_3040);
or U3431 (N_3431,N_3247,N_3086);
or U3432 (N_3432,N_3138,N_3119);
and U3433 (N_3433,N_3263,N_3064);
and U3434 (N_3434,N_3136,N_3256);
xor U3435 (N_3435,N_3147,N_3051);
nand U3436 (N_3436,N_3023,N_3195);
nand U3437 (N_3437,N_3266,N_3157);
or U3438 (N_3438,N_3190,N_3227);
nand U3439 (N_3439,N_3220,N_3133);
nor U3440 (N_3440,N_3277,N_3239);
nand U3441 (N_3441,N_3124,N_3153);
and U3442 (N_3442,N_3088,N_3296);
xor U3443 (N_3443,N_3205,N_3096);
or U3444 (N_3444,N_3254,N_3024);
nand U3445 (N_3445,N_3038,N_3260);
nand U3446 (N_3446,N_3234,N_3246);
and U3447 (N_3447,N_3252,N_3298);
or U3448 (N_3448,N_3294,N_3251);
and U3449 (N_3449,N_3264,N_3141);
and U3450 (N_3450,N_3232,N_3285);
nor U3451 (N_3451,N_3183,N_3247);
or U3452 (N_3452,N_3106,N_3114);
nand U3453 (N_3453,N_3175,N_3040);
or U3454 (N_3454,N_3137,N_3211);
xnor U3455 (N_3455,N_3050,N_3080);
or U3456 (N_3456,N_3076,N_3014);
nor U3457 (N_3457,N_3190,N_3252);
nand U3458 (N_3458,N_3264,N_3155);
and U3459 (N_3459,N_3037,N_3079);
or U3460 (N_3460,N_3214,N_3232);
xor U3461 (N_3461,N_3051,N_3101);
nor U3462 (N_3462,N_3254,N_3020);
nand U3463 (N_3463,N_3013,N_3160);
nor U3464 (N_3464,N_3291,N_3294);
xor U3465 (N_3465,N_3010,N_3038);
nand U3466 (N_3466,N_3196,N_3024);
or U3467 (N_3467,N_3193,N_3029);
nand U3468 (N_3468,N_3290,N_3168);
and U3469 (N_3469,N_3234,N_3013);
nand U3470 (N_3470,N_3043,N_3134);
nor U3471 (N_3471,N_3173,N_3197);
or U3472 (N_3472,N_3259,N_3071);
nand U3473 (N_3473,N_3169,N_3197);
nor U3474 (N_3474,N_3015,N_3007);
or U3475 (N_3475,N_3040,N_3145);
or U3476 (N_3476,N_3234,N_3029);
xor U3477 (N_3477,N_3145,N_3104);
nand U3478 (N_3478,N_3161,N_3206);
or U3479 (N_3479,N_3189,N_3174);
nand U3480 (N_3480,N_3052,N_3264);
and U3481 (N_3481,N_3119,N_3124);
and U3482 (N_3482,N_3086,N_3009);
xnor U3483 (N_3483,N_3078,N_3212);
nand U3484 (N_3484,N_3237,N_3202);
or U3485 (N_3485,N_3046,N_3074);
xnor U3486 (N_3486,N_3192,N_3268);
xor U3487 (N_3487,N_3069,N_3277);
nor U3488 (N_3488,N_3039,N_3265);
nand U3489 (N_3489,N_3068,N_3262);
nor U3490 (N_3490,N_3217,N_3252);
nor U3491 (N_3491,N_3034,N_3018);
nor U3492 (N_3492,N_3123,N_3239);
and U3493 (N_3493,N_3298,N_3133);
nand U3494 (N_3494,N_3144,N_3130);
nor U3495 (N_3495,N_3009,N_3079);
and U3496 (N_3496,N_3200,N_3084);
or U3497 (N_3497,N_3212,N_3081);
nor U3498 (N_3498,N_3174,N_3231);
nand U3499 (N_3499,N_3087,N_3145);
xor U3500 (N_3500,N_3055,N_3178);
nand U3501 (N_3501,N_3036,N_3152);
and U3502 (N_3502,N_3262,N_3061);
and U3503 (N_3503,N_3225,N_3011);
nor U3504 (N_3504,N_3164,N_3025);
nor U3505 (N_3505,N_3264,N_3089);
nor U3506 (N_3506,N_3223,N_3024);
nor U3507 (N_3507,N_3292,N_3057);
nor U3508 (N_3508,N_3065,N_3148);
nor U3509 (N_3509,N_3297,N_3169);
or U3510 (N_3510,N_3283,N_3061);
and U3511 (N_3511,N_3250,N_3039);
nand U3512 (N_3512,N_3073,N_3139);
nand U3513 (N_3513,N_3276,N_3240);
xnor U3514 (N_3514,N_3238,N_3116);
nand U3515 (N_3515,N_3208,N_3290);
or U3516 (N_3516,N_3139,N_3201);
xnor U3517 (N_3517,N_3081,N_3012);
xnor U3518 (N_3518,N_3259,N_3179);
nand U3519 (N_3519,N_3092,N_3293);
nor U3520 (N_3520,N_3008,N_3012);
xnor U3521 (N_3521,N_3077,N_3065);
nand U3522 (N_3522,N_3105,N_3085);
or U3523 (N_3523,N_3062,N_3187);
nor U3524 (N_3524,N_3227,N_3155);
or U3525 (N_3525,N_3016,N_3135);
xnor U3526 (N_3526,N_3165,N_3123);
nand U3527 (N_3527,N_3282,N_3100);
and U3528 (N_3528,N_3243,N_3021);
xnor U3529 (N_3529,N_3221,N_3077);
xnor U3530 (N_3530,N_3207,N_3272);
nor U3531 (N_3531,N_3185,N_3165);
or U3532 (N_3532,N_3078,N_3188);
nand U3533 (N_3533,N_3172,N_3117);
nand U3534 (N_3534,N_3012,N_3204);
and U3535 (N_3535,N_3273,N_3006);
and U3536 (N_3536,N_3212,N_3293);
nand U3537 (N_3537,N_3273,N_3181);
or U3538 (N_3538,N_3252,N_3254);
nand U3539 (N_3539,N_3058,N_3254);
nand U3540 (N_3540,N_3152,N_3212);
xor U3541 (N_3541,N_3252,N_3067);
and U3542 (N_3542,N_3029,N_3065);
and U3543 (N_3543,N_3134,N_3175);
and U3544 (N_3544,N_3019,N_3232);
or U3545 (N_3545,N_3030,N_3178);
or U3546 (N_3546,N_3149,N_3297);
nor U3547 (N_3547,N_3094,N_3072);
nor U3548 (N_3548,N_3056,N_3127);
nand U3549 (N_3549,N_3052,N_3199);
or U3550 (N_3550,N_3182,N_3181);
or U3551 (N_3551,N_3291,N_3048);
xnor U3552 (N_3552,N_3192,N_3060);
xor U3553 (N_3553,N_3178,N_3063);
nor U3554 (N_3554,N_3050,N_3261);
nor U3555 (N_3555,N_3259,N_3048);
xnor U3556 (N_3556,N_3049,N_3203);
nor U3557 (N_3557,N_3272,N_3146);
nor U3558 (N_3558,N_3069,N_3058);
nand U3559 (N_3559,N_3144,N_3146);
nor U3560 (N_3560,N_3275,N_3072);
and U3561 (N_3561,N_3240,N_3177);
or U3562 (N_3562,N_3189,N_3080);
xnor U3563 (N_3563,N_3291,N_3134);
nand U3564 (N_3564,N_3074,N_3140);
xnor U3565 (N_3565,N_3047,N_3194);
and U3566 (N_3566,N_3204,N_3130);
or U3567 (N_3567,N_3277,N_3273);
and U3568 (N_3568,N_3137,N_3125);
or U3569 (N_3569,N_3089,N_3296);
xnor U3570 (N_3570,N_3124,N_3000);
nand U3571 (N_3571,N_3213,N_3212);
nand U3572 (N_3572,N_3142,N_3094);
nand U3573 (N_3573,N_3097,N_3260);
and U3574 (N_3574,N_3185,N_3017);
nor U3575 (N_3575,N_3002,N_3249);
or U3576 (N_3576,N_3227,N_3173);
nand U3577 (N_3577,N_3115,N_3171);
xnor U3578 (N_3578,N_3225,N_3267);
nand U3579 (N_3579,N_3137,N_3140);
and U3580 (N_3580,N_3002,N_3288);
or U3581 (N_3581,N_3243,N_3183);
or U3582 (N_3582,N_3222,N_3120);
nand U3583 (N_3583,N_3089,N_3090);
nor U3584 (N_3584,N_3000,N_3079);
nand U3585 (N_3585,N_3198,N_3231);
xor U3586 (N_3586,N_3252,N_3172);
or U3587 (N_3587,N_3202,N_3116);
and U3588 (N_3588,N_3027,N_3035);
nand U3589 (N_3589,N_3111,N_3116);
and U3590 (N_3590,N_3164,N_3108);
and U3591 (N_3591,N_3043,N_3108);
and U3592 (N_3592,N_3206,N_3096);
and U3593 (N_3593,N_3110,N_3178);
and U3594 (N_3594,N_3223,N_3017);
xor U3595 (N_3595,N_3268,N_3113);
xor U3596 (N_3596,N_3101,N_3295);
xnor U3597 (N_3597,N_3153,N_3187);
xor U3598 (N_3598,N_3090,N_3007);
or U3599 (N_3599,N_3142,N_3060);
nor U3600 (N_3600,N_3309,N_3340);
nor U3601 (N_3601,N_3521,N_3398);
xor U3602 (N_3602,N_3424,N_3513);
xor U3603 (N_3603,N_3584,N_3300);
or U3604 (N_3604,N_3525,N_3515);
or U3605 (N_3605,N_3569,N_3532);
nor U3606 (N_3606,N_3465,N_3423);
nor U3607 (N_3607,N_3575,N_3481);
nand U3608 (N_3608,N_3301,N_3302);
nor U3609 (N_3609,N_3567,N_3374);
nand U3610 (N_3610,N_3583,N_3455);
nor U3611 (N_3611,N_3313,N_3528);
and U3612 (N_3612,N_3571,N_3323);
or U3613 (N_3613,N_3500,N_3328);
xor U3614 (N_3614,N_3557,N_3399);
and U3615 (N_3615,N_3482,N_3409);
or U3616 (N_3616,N_3509,N_3363);
or U3617 (N_3617,N_3450,N_3581);
nor U3618 (N_3618,N_3457,N_3582);
nand U3619 (N_3619,N_3344,N_3564);
nand U3620 (N_3620,N_3317,N_3568);
nand U3621 (N_3621,N_3308,N_3422);
xor U3622 (N_3622,N_3362,N_3458);
or U3623 (N_3623,N_3596,N_3572);
and U3624 (N_3624,N_3499,N_3342);
nand U3625 (N_3625,N_3442,N_3453);
or U3626 (N_3626,N_3512,N_3413);
xor U3627 (N_3627,N_3530,N_3590);
or U3628 (N_3628,N_3594,N_3314);
xor U3629 (N_3629,N_3303,N_3554);
and U3630 (N_3630,N_3373,N_3587);
or U3631 (N_3631,N_3452,N_3316);
and U3632 (N_3632,N_3484,N_3524);
nor U3633 (N_3633,N_3329,N_3561);
or U3634 (N_3634,N_3573,N_3527);
or U3635 (N_3635,N_3480,N_3425);
nor U3636 (N_3636,N_3326,N_3574);
xor U3637 (N_3637,N_3548,N_3531);
xor U3638 (N_3638,N_3400,N_3421);
or U3639 (N_3639,N_3580,N_3339);
and U3640 (N_3640,N_3321,N_3414);
or U3641 (N_3641,N_3334,N_3545);
and U3642 (N_3642,N_3537,N_3430);
nor U3643 (N_3643,N_3366,N_3438);
and U3644 (N_3644,N_3351,N_3419);
nor U3645 (N_3645,N_3553,N_3467);
and U3646 (N_3646,N_3379,N_3591);
and U3647 (N_3647,N_3497,N_3431);
nor U3648 (N_3648,N_3459,N_3377);
nand U3649 (N_3649,N_3353,N_3487);
or U3650 (N_3650,N_3320,N_3415);
nor U3651 (N_3651,N_3420,N_3395);
nor U3652 (N_3652,N_3350,N_3535);
and U3653 (N_3653,N_3307,N_3376);
xnor U3654 (N_3654,N_3389,N_3386);
xnor U3655 (N_3655,N_3519,N_3485);
nand U3656 (N_3656,N_3354,N_3390);
or U3657 (N_3657,N_3331,N_3370);
or U3658 (N_3658,N_3401,N_3526);
xor U3659 (N_3659,N_3489,N_3556);
or U3660 (N_3660,N_3396,N_3516);
or U3661 (N_3661,N_3387,N_3468);
xnor U3662 (N_3662,N_3598,N_3529);
and U3663 (N_3663,N_3547,N_3506);
nand U3664 (N_3664,N_3551,N_3483);
or U3665 (N_3665,N_3437,N_3358);
and U3666 (N_3666,N_3406,N_3416);
nand U3667 (N_3667,N_3562,N_3433);
or U3668 (N_3668,N_3470,N_3534);
nor U3669 (N_3669,N_3381,N_3552);
nand U3670 (N_3670,N_3349,N_3305);
xnor U3671 (N_3671,N_3510,N_3549);
or U3672 (N_3672,N_3394,N_3566);
and U3673 (N_3673,N_3368,N_3471);
and U3674 (N_3674,N_3410,N_3397);
nand U3675 (N_3675,N_3518,N_3476);
xor U3676 (N_3676,N_3443,N_3428);
nand U3677 (N_3677,N_3463,N_3536);
xnor U3678 (N_3678,N_3507,N_3599);
nor U3679 (N_3679,N_3523,N_3492);
nor U3680 (N_3680,N_3360,N_3446);
or U3681 (N_3681,N_3347,N_3348);
nand U3682 (N_3682,N_3336,N_3511);
and U3683 (N_3683,N_3462,N_3346);
or U3684 (N_3684,N_3322,N_3595);
xor U3685 (N_3685,N_3404,N_3495);
nand U3686 (N_3686,N_3585,N_3319);
nand U3687 (N_3687,N_3392,N_3417);
xor U3688 (N_3688,N_3345,N_3324);
nor U3689 (N_3689,N_3445,N_3456);
or U3690 (N_3690,N_3441,N_3361);
nand U3691 (N_3691,N_3550,N_3490);
nor U3692 (N_3692,N_3440,N_3447);
nor U3693 (N_3693,N_3586,N_3576);
and U3694 (N_3694,N_3543,N_3474);
and U3695 (N_3695,N_3477,N_3449);
nand U3696 (N_3696,N_3589,N_3408);
or U3697 (N_3697,N_3472,N_3411);
or U3698 (N_3698,N_3563,N_3382);
or U3699 (N_3699,N_3357,N_3356);
nand U3700 (N_3700,N_3502,N_3306);
nor U3701 (N_3701,N_3426,N_3337);
or U3702 (N_3702,N_3486,N_3435);
or U3703 (N_3703,N_3432,N_3375);
nand U3704 (N_3704,N_3384,N_3369);
nand U3705 (N_3705,N_3546,N_3315);
or U3706 (N_3706,N_3577,N_3365);
or U3707 (N_3707,N_3380,N_3407);
xnor U3708 (N_3708,N_3544,N_3517);
nand U3709 (N_3709,N_3318,N_3391);
nor U3710 (N_3710,N_3451,N_3520);
or U3711 (N_3711,N_3540,N_3388);
nor U3712 (N_3712,N_3460,N_3367);
or U3713 (N_3713,N_3372,N_3464);
nor U3714 (N_3714,N_3429,N_3555);
and U3715 (N_3715,N_3505,N_3558);
xor U3716 (N_3716,N_3393,N_3473);
nor U3717 (N_3717,N_3402,N_3559);
xor U3718 (N_3718,N_3496,N_3338);
nor U3719 (N_3719,N_3493,N_3427);
xnor U3720 (N_3720,N_3466,N_3341);
and U3721 (N_3721,N_3570,N_3578);
or U3722 (N_3722,N_3412,N_3359);
nor U3723 (N_3723,N_3352,N_3355);
or U3724 (N_3724,N_3593,N_3325);
nor U3725 (N_3725,N_3327,N_3504);
and U3726 (N_3726,N_3335,N_3597);
xor U3727 (N_3727,N_3461,N_3378);
nand U3728 (N_3728,N_3312,N_3383);
or U3729 (N_3729,N_3444,N_3439);
or U3730 (N_3730,N_3522,N_3514);
or U3731 (N_3731,N_3418,N_3371);
and U3732 (N_3732,N_3311,N_3330);
and U3733 (N_3733,N_3479,N_3454);
or U3734 (N_3734,N_3503,N_3436);
nor U3735 (N_3735,N_3592,N_3588);
nand U3736 (N_3736,N_3333,N_3488);
nor U3737 (N_3737,N_3434,N_3494);
nand U3738 (N_3738,N_3508,N_3560);
nor U3739 (N_3739,N_3541,N_3475);
xnor U3740 (N_3740,N_3533,N_3448);
and U3741 (N_3741,N_3469,N_3310);
and U3742 (N_3742,N_3403,N_3385);
nor U3743 (N_3743,N_3304,N_3364);
nand U3744 (N_3744,N_3478,N_3565);
xor U3745 (N_3745,N_3501,N_3579);
and U3746 (N_3746,N_3542,N_3539);
xor U3747 (N_3747,N_3498,N_3538);
xnor U3748 (N_3748,N_3343,N_3332);
or U3749 (N_3749,N_3405,N_3491);
or U3750 (N_3750,N_3479,N_3564);
nor U3751 (N_3751,N_3413,N_3496);
nand U3752 (N_3752,N_3574,N_3333);
nor U3753 (N_3753,N_3302,N_3324);
nor U3754 (N_3754,N_3367,N_3500);
nor U3755 (N_3755,N_3435,N_3492);
nand U3756 (N_3756,N_3345,N_3363);
xnor U3757 (N_3757,N_3417,N_3383);
or U3758 (N_3758,N_3311,N_3541);
nand U3759 (N_3759,N_3346,N_3417);
nand U3760 (N_3760,N_3443,N_3390);
and U3761 (N_3761,N_3568,N_3476);
nand U3762 (N_3762,N_3560,N_3488);
nand U3763 (N_3763,N_3408,N_3403);
xor U3764 (N_3764,N_3463,N_3548);
nor U3765 (N_3765,N_3446,N_3421);
nand U3766 (N_3766,N_3364,N_3392);
or U3767 (N_3767,N_3382,N_3408);
xor U3768 (N_3768,N_3510,N_3360);
nand U3769 (N_3769,N_3336,N_3345);
nor U3770 (N_3770,N_3330,N_3595);
nand U3771 (N_3771,N_3526,N_3354);
nor U3772 (N_3772,N_3535,N_3513);
xor U3773 (N_3773,N_3542,N_3448);
nor U3774 (N_3774,N_3580,N_3583);
xnor U3775 (N_3775,N_3551,N_3491);
xnor U3776 (N_3776,N_3490,N_3353);
xnor U3777 (N_3777,N_3561,N_3461);
nor U3778 (N_3778,N_3499,N_3366);
xnor U3779 (N_3779,N_3591,N_3380);
or U3780 (N_3780,N_3519,N_3340);
or U3781 (N_3781,N_3328,N_3538);
nor U3782 (N_3782,N_3561,N_3407);
nand U3783 (N_3783,N_3396,N_3538);
nor U3784 (N_3784,N_3348,N_3555);
xnor U3785 (N_3785,N_3306,N_3391);
xnor U3786 (N_3786,N_3460,N_3361);
and U3787 (N_3787,N_3570,N_3468);
and U3788 (N_3788,N_3484,N_3552);
nand U3789 (N_3789,N_3302,N_3344);
and U3790 (N_3790,N_3531,N_3570);
xnor U3791 (N_3791,N_3406,N_3320);
or U3792 (N_3792,N_3339,N_3454);
or U3793 (N_3793,N_3437,N_3518);
nor U3794 (N_3794,N_3335,N_3541);
nand U3795 (N_3795,N_3312,N_3497);
and U3796 (N_3796,N_3586,N_3354);
and U3797 (N_3797,N_3517,N_3467);
and U3798 (N_3798,N_3552,N_3465);
nand U3799 (N_3799,N_3581,N_3396);
or U3800 (N_3800,N_3310,N_3586);
nand U3801 (N_3801,N_3573,N_3425);
nor U3802 (N_3802,N_3486,N_3323);
nor U3803 (N_3803,N_3373,N_3480);
nand U3804 (N_3804,N_3496,N_3568);
nand U3805 (N_3805,N_3446,N_3430);
nor U3806 (N_3806,N_3367,N_3303);
or U3807 (N_3807,N_3384,N_3328);
xnor U3808 (N_3808,N_3510,N_3314);
nor U3809 (N_3809,N_3369,N_3399);
nor U3810 (N_3810,N_3554,N_3448);
nand U3811 (N_3811,N_3398,N_3350);
or U3812 (N_3812,N_3336,N_3488);
xor U3813 (N_3813,N_3318,N_3519);
and U3814 (N_3814,N_3390,N_3569);
nor U3815 (N_3815,N_3428,N_3344);
nand U3816 (N_3816,N_3505,N_3492);
or U3817 (N_3817,N_3581,N_3311);
and U3818 (N_3818,N_3515,N_3329);
xnor U3819 (N_3819,N_3307,N_3385);
and U3820 (N_3820,N_3569,N_3334);
and U3821 (N_3821,N_3341,N_3416);
nor U3822 (N_3822,N_3322,N_3580);
nand U3823 (N_3823,N_3539,N_3445);
nor U3824 (N_3824,N_3470,N_3400);
nand U3825 (N_3825,N_3476,N_3356);
xnor U3826 (N_3826,N_3514,N_3419);
or U3827 (N_3827,N_3384,N_3338);
xor U3828 (N_3828,N_3523,N_3395);
xor U3829 (N_3829,N_3567,N_3483);
nand U3830 (N_3830,N_3498,N_3518);
nor U3831 (N_3831,N_3455,N_3310);
nand U3832 (N_3832,N_3304,N_3346);
or U3833 (N_3833,N_3590,N_3314);
and U3834 (N_3834,N_3321,N_3404);
xnor U3835 (N_3835,N_3502,N_3497);
or U3836 (N_3836,N_3599,N_3388);
or U3837 (N_3837,N_3354,N_3463);
or U3838 (N_3838,N_3455,N_3356);
xor U3839 (N_3839,N_3397,N_3306);
nor U3840 (N_3840,N_3386,N_3350);
nand U3841 (N_3841,N_3450,N_3510);
or U3842 (N_3842,N_3553,N_3507);
nor U3843 (N_3843,N_3454,N_3315);
xor U3844 (N_3844,N_3553,N_3561);
xor U3845 (N_3845,N_3313,N_3571);
or U3846 (N_3846,N_3433,N_3371);
xor U3847 (N_3847,N_3538,N_3452);
or U3848 (N_3848,N_3393,N_3420);
and U3849 (N_3849,N_3376,N_3340);
and U3850 (N_3850,N_3385,N_3368);
xnor U3851 (N_3851,N_3451,N_3400);
nor U3852 (N_3852,N_3507,N_3406);
xnor U3853 (N_3853,N_3354,N_3583);
xnor U3854 (N_3854,N_3518,N_3352);
and U3855 (N_3855,N_3430,N_3473);
nand U3856 (N_3856,N_3473,N_3563);
and U3857 (N_3857,N_3388,N_3473);
xnor U3858 (N_3858,N_3457,N_3371);
xor U3859 (N_3859,N_3341,N_3582);
or U3860 (N_3860,N_3321,N_3322);
xor U3861 (N_3861,N_3588,N_3413);
xnor U3862 (N_3862,N_3509,N_3378);
and U3863 (N_3863,N_3406,N_3552);
or U3864 (N_3864,N_3586,N_3487);
or U3865 (N_3865,N_3402,N_3571);
or U3866 (N_3866,N_3307,N_3460);
xor U3867 (N_3867,N_3531,N_3449);
nand U3868 (N_3868,N_3513,N_3501);
xnor U3869 (N_3869,N_3407,N_3586);
and U3870 (N_3870,N_3516,N_3346);
or U3871 (N_3871,N_3392,N_3589);
nand U3872 (N_3872,N_3555,N_3527);
xnor U3873 (N_3873,N_3473,N_3456);
or U3874 (N_3874,N_3310,N_3494);
nand U3875 (N_3875,N_3555,N_3476);
xor U3876 (N_3876,N_3437,N_3504);
nand U3877 (N_3877,N_3443,N_3559);
or U3878 (N_3878,N_3429,N_3505);
xnor U3879 (N_3879,N_3379,N_3316);
and U3880 (N_3880,N_3577,N_3417);
nand U3881 (N_3881,N_3548,N_3428);
or U3882 (N_3882,N_3519,N_3320);
nand U3883 (N_3883,N_3410,N_3548);
xor U3884 (N_3884,N_3367,N_3451);
nand U3885 (N_3885,N_3395,N_3465);
and U3886 (N_3886,N_3555,N_3492);
nand U3887 (N_3887,N_3530,N_3319);
xor U3888 (N_3888,N_3443,N_3511);
xor U3889 (N_3889,N_3304,N_3560);
and U3890 (N_3890,N_3539,N_3444);
nand U3891 (N_3891,N_3564,N_3394);
nand U3892 (N_3892,N_3489,N_3563);
nand U3893 (N_3893,N_3461,N_3450);
and U3894 (N_3894,N_3404,N_3558);
or U3895 (N_3895,N_3593,N_3495);
nand U3896 (N_3896,N_3575,N_3379);
or U3897 (N_3897,N_3509,N_3332);
or U3898 (N_3898,N_3314,N_3433);
or U3899 (N_3899,N_3364,N_3445);
xnor U3900 (N_3900,N_3849,N_3884);
xor U3901 (N_3901,N_3638,N_3613);
or U3902 (N_3902,N_3674,N_3844);
nand U3903 (N_3903,N_3852,N_3856);
and U3904 (N_3904,N_3705,N_3714);
and U3905 (N_3905,N_3658,N_3748);
or U3906 (N_3906,N_3710,N_3707);
nand U3907 (N_3907,N_3729,N_3723);
nor U3908 (N_3908,N_3612,N_3814);
xnor U3909 (N_3909,N_3838,N_3894);
or U3910 (N_3910,N_3857,N_3810);
or U3911 (N_3911,N_3822,N_3864);
or U3912 (N_3912,N_3732,N_3731);
nor U3913 (N_3913,N_3833,N_3642);
nor U3914 (N_3914,N_3828,N_3618);
and U3915 (N_3915,N_3869,N_3881);
or U3916 (N_3916,N_3666,N_3791);
nand U3917 (N_3917,N_3850,N_3811);
or U3918 (N_3918,N_3626,N_3718);
or U3919 (N_3919,N_3848,N_3819);
or U3920 (N_3920,N_3720,N_3829);
and U3921 (N_3921,N_3773,N_3740);
or U3922 (N_3922,N_3756,N_3851);
nor U3923 (N_3923,N_3686,N_3641);
and U3924 (N_3924,N_3895,N_3725);
nand U3925 (N_3925,N_3661,N_3610);
and U3926 (N_3926,N_3633,N_3853);
or U3927 (N_3927,N_3687,N_3761);
or U3928 (N_3928,N_3805,N_3672);
xor U3929 (N_3929,N_3681,N_3632);
xnor U3930 (N_3930,N_3823,N_3649);
and U3931 (N_3931,N_3647,N_3860);
nor U3932 (N_3932,N_3751,N_3623);
nand U3933 (N_3933,N_3874,N_3676);
nand U3934 (N_3934,N_3817,N_3634);
and U3935 (N_3935,N_3889,N_3789);
nand U3936 (N_3936,N_3701,N_3772);
nand U3937 (N_3937,N_3809,N_3782);
or U3938 (N_3938,N_3709,N_3630);
or U3939 (N_3939,N_3893,N_3764);
xnor U3940 (N_3940,N_3797,N_3767);
nor U3941 (N_3941,N_3624,N_3898);
xor U3942 (N_3942,N_3667,N_3783);
xnor U3943 (N_3943,N_3818,N_3603);
nand U3944 (N_3944,N_3745,N_3801);
xor U3945 (N_3945,N_3719,N_3752);
or U3946 (N_3946,N_3741,N_3680);
xnor U3947 (N_3947,N_3816,N_3652);
xor U3948 (N_3948,N_3639,N_3836);
and U3949 (N_3949,N_3826,N_3615);
and U3950 (N_3950,N_3820,N_3616);
xnor U3951 (N_3951,N_3675,N_3700);
or U3952 (N_3952,N_3862,N_3795);
nand U3953 (N_3953,N_3769,N_3839);
nor U3954 (N_3954,N_3799,N_3770);
nand U3955 (N_3955,N_3722,N_3825);
nand U3956 (N_3956,N_3780,N_3713);
and U3957 (N_3957,N_3653,N_3673);
nor U3958 (N_3958,N_3854,N_3684);
xor U3959 (N_3959,N_3656,N_3785);
nor U3960 (N_3960,N_3754,N_3747);
xnor U3961 (N_3961,N_3694,N_3774);
nor U3962 (N_3962,N_3784,N_3662);
nand U3963 (N_3963,N_3885,N_3827);
or U3964 (N_3964,N_3891,N_3644);
xnor U3965 (N_3965,N_3878,N_3742);
or U3966 (N_3966,N_3629,N_3604);
nand U3967 (N_3967,N_3706,N_3762);
nand U3968 (N_3968,N_3688,N_3858);
and U3969 (N_3969,N_3602,N_3807);
nor U3970 (N_3970,N_3699,N_3728);
nand U3971 (N_3971,N_3883,N_3696);
nand U3972 (N_3972,N_3697,N_3779);
xor U3973 (N_3973,N_3620,N_3776);
and U3974 (N_3974,N_3685,N_3781);
or U3975 (N_3975,N_3708,N_3689);
nand U3976 (N_3976,N_3636,N_3736);
or U3977 (N_3977,N_3665,N_3771);
nand U3978 (N_3978,N_3601,N_3803);
and U3979 (N_3979,N_3733,N_3617);
nor U3980 (N_3980,N_3873,N_3608);
nand U3981 (N_3981,N_3765,N_3759);
nand U3982 (N_3982,N_3690,N_3808);
or U3983 (N_3983,N_3605,N_3875);
xor U3984 (N_3984,N_3715,N_3861);
nor U3985 (N_3985,N_3804,N_3755);
and U3986 (N_3986,N_3695,N_3835);
or U3987 (N_3987,N_3669,N_3812);
nor U3988 (N_3988,N_3778,N_3749);
nor U3989 (N_3989,N_3768,N_3668);
nor U3990 (N_3990,N_3683,N_3846);
nand U3991 (N_3991,N_3867,N_3787);
nand U3992 (N_3992,N_3793,N_3831);
xor U3993 (N_3993,N_3637,N_3794);
nand U3994 (N_3994,N_3703,N_3788);
xnor U3995 (N_3995,N_3888,N_3664);
nor U3996 (N_3996,N_3663,N_3786);
and U3997 (N_3997,N_3657,N_3744);
xor U3998 (N_3998,N_3607,N_3842);
nor U3999 (N_3999,N_3646,N_3868);
or U4000 (N_4000,N_3880,N_3611);
nor U4001 (N_4001,N_3671,N_3650);
and U4002 (N_4002,N_3739,N_3832);
or U4003 (N_4003,N_3872,N_3899);
and U4004 (N_4004,N_3830,N_3758);
nand U4005 (N_4005,N_3679,N_3753);
nor U4006 (N_4006,N_3843,N_3897);
xnor U4007 (N_4007,N_3628,N_3892);
xor U4008 (N_4008,N_3737,N_3704);
and U4009 (N_4009,N_3877,N_3845);
and U4010 (N_4010,N_3655,N_3651);
or U4011 (N_4011,N_3627,N_3760);
and U4012 (N_4012,N_3727,N_3757);
and U4013 (N_4013,N_3721,N_3859);
or U4014 (N_4014,N_3743,N_3600);
xnor U4015 (N_4015,N_3643,N_3802);
nor U4016 (N_4016,N_3625,N_3645);
and U4017 (N_4017,N_3640,N_3792);
nor U4018 (N_4018,N_3648,N_3717);
or U4019 (N_4019,N_3834,N_3670);
xnor U4020 (N_4020,N_3738,N_3896);
xnor U4021 (N_4021,N_3693,N_3824);
nor U4022 (N_4022,N_3614,N_3659);
and U4023 (N_4023,N_3886,N_3724);
and U4024 (N_4024,N_3735,N_3635);
and U4025 (N_4025,N_3682,N_3870);
and U4026 (N_4026,N_3815,N_3882);
or U4027 (N_4027,N_3866,N_3702);
or U4028 (N_4028,N_3766,N_3876);
nand U4029 (N_4029,N_3763,N_3606);
nand U4030 (N_4030,N_3726,N_3631);
nand U4031 (N_4031,N_3837,N_3678);
xor U4032 (N_4032,N_3887,N_3798);
nor U4033 (N_4033,N_3821,N_3865);
nor U4034 (N_4034,N_3660,N_3847);
or U4035 (N_4035,N_3855,N_3622);
or U4036 (N_4036,N_3698,N_3800);
nand U4037 (N_4037,N_3806,N_3841);
and U4038 (N_4038,N_3890,N_3871);
xor U4039 (N_4039,N_3730,N_3746);
nor U4040 (N_4040,N_3750,N_3692);
and U4041 (N_4041,N_3863,N_3716);
xnor U4042 (N_4042,N_3879,N_3621);
and U4043 (N_4043,N_3677,N_3796);
xnor U4044 (N_4044,N_3840,N_3609);
xor U4045 (N_4045,N_3691,N_3711);
nor U4046 (N_4046,N_3734,N_3790);
nor U4047 (N_4047,N_3775,N_3654);
nand U4048 (N_4048,N_3777,N_3712);
nor U4049 (N_4049,N_3619,N_3813);
nor U4050 (N_4050,N_3864,N_3818);
nor U4051 (N_4051,N_3699,N_3674);
nand U4052 (N_4052,N_3882,N_3648);
nor U4053 (N_4053,N_3791,N_3673);
or U4054 (N_4054,N_3755,N_3871);
nor U4055 (N_4055,N_3860,N_3866);
and U4056 (N_4056,N_3777,N_3605);
xnor U4057 (N_4057,N_3844,N_3615);
and U4058 (N_4058,N_3767,N_3851);
nor U4059 (N_4059,N_3607,N_3854);
nand U4060 (N_4060,N_3740,N_3769);
nor U4061 (N_4061,N_3723,N_3817);
and U4062 (N_4062,N_3712,N_3737);
or U4063 (N_4063,N_3747,N_3635);
and U4064 (N_4064,N_3846,N_3772);
xnor U4065 (N_4065,N_3705,N_3609);
nand U4066 (N_4066,N_3645,N_3715);
nand U4067 (N_4067,N_3677,N_3670);
nand U4068 (N_4068,N_3757,N_3697);
and U4069 (N_4069,N_3620,N_3629);
and U4070 (N_4070,N_3623,N_3733);
xnor U4071 (N_4071,N_3842,N_3852);
or U4072 (N_4072,N_3821,N_3778);
nand U4073 (N_4073,N_3889,N_3625);
nor U4074 (N_4074,N_3812,N_3845);
nor U4075 (N_4075,N_3898,N_3876);
nand U4076 (N_4076,N_3836,N_3633);
and U4077 (N_4077,N_3876,N_3869);
nand U4078 (N_4078,N_3850,N_3617);
nand U4079 (N_4079,N_3889,N_3704);
or U4080 (N_4080,N_3605,N_3723);
and U4081 (N_4081,N_3763,N_3838);
nor U4082 (N_4082,N_3821,N_3816);
or U4083 (N_4083,N_3887,N_3741);
nor U4084 (N_4084,N_3602,N_3682);
nor U4085 (N_4085,N_3850,N_3602);
nand U4086 (N_4086,N_3768,N_3613);
or U4087 (N_4087,N_3884,N_3626);
nor U4088 (N_4088,N_3617,N_3644);
and U4089 (N_4089,N_3682,N_3638);
xor U4090 (N_4090,N_3752,N_3758);
nor U4091 (N_4091,N_3821,N_3794);
nand U4092 (N_4092,N_3759,N_3675);
nand U4093 (N_4093,N_3789,N_3765);
or U4094 (N_4094,N_3668,N_3724);
or U4095 (N_4095,N_3849,N_3649);
xnor U4096 (N_4096,N_3681,N_3641);
and U4097 (N_4097,N_3874,N_3602);
nand U4098 (N_4098,N_3776,N_3653);
or U4099 (N_4099,N_3641,N_3818);
xor U4100 (N_4100,N_3654,N_3730);
nand U4101 (N_4101,N_3617,N_3763);
xor U4102 (N_4102,N_3680,N_3711);
or U4103 (N_4103,N_3888,N_3700);
xnor U4104 (N_4104,N_3837,N_3713);
and U4105 (N_4105,N_3675,N_3645);
xnor U4106 (N_4106,N_3626,N_3777);
nand U4107 (N_4107,N_3868,N_3670);
nor U4108 (N_4108,N_3633,N_3800);
and U4109 (N_4109,N_3691,N_3738);
nor U4110 (N_4110,N_3827,N_3814);
nand U4111 (N_4111,N_3699,N_3641);
or U4112 (N_4112,N_3737,N_3717);
and U4113 (N_4113,N_3651,N_3762);
xor U4114 (N_4114,N_3687,N_3829);
nand U4115 (N_4115,N_3707,N_3770);
nor U4116 (N_4116,N_3860,N_3832);
nand U4117 (N_4117,N_3873,N_3751);
or U4118 (N_4118,N_3636,N_3627);
xnor U4119 (N_4119,N_3883,N_3862);
xnor U4120 (N_4120,N_3863,N_3776);
or U4121 (N_4121,N_3827,N_3869);
or U4122 (N_4122,N_3853,N_3809);
or U4123 (N_4123,N_3862,N_3693);
and U4124 (N_4124,N_3823,N_3854);
nor U4125 (N_4125,N_3700,N_3813);
xnor U4126 (N_4126,N_3775,N_3781);
nand U4127 (N_4127,N_3645,N_3831);
nand U4128 (N_4128,N_3700,N_3734);
and U4129 (N_4129,N_3803,N_3666);
or U4130 (N_4130,N_3711,N_3794);
xnor U4131 (N_4131,N_3772,N_3776);
xnor U4132 (N_4132,N_3612,N_3655);
or U4133 (N_4133,N_3706,N_3686);
xnor U4134 (N_4134,N_3600,N_3736);
xnor U4135 (N_4135,N_3899,N_3889);
nor U4136 (N_4136,N_3614,N_3725);
and U4137 (N_4137,N_3718,N_3666);
nor U4138 (N_4138,N_3631,N_3750);
xor U4139 (N_4139,N_3884,N_3678);
nand U4140 (N_4140,N_3862,N_3736);
nand U4141 (N_4141,N_3790,N_3623);
or U4142 (N_4142,N_3702,N_3803);
or U4143 (N_4143,N_3833,N_3777);
xor U4144 (N_4144,N_3708,N_3897);
or U4145 (N_4145,N_3681,N_3614);
nand U4146 (N_4146,N_3761,N_3667);
nor U4147 (N_4147,N_3603,N_3606);
xnor U4148 (N_4148,N_3881,N_3655);
xnor U4149 (N_4149,N_3768,N_3601);
xor U4150 (N_4150,N_3690,N_3783);
xnor U4151 (N_4151,N_3813,N_3878);
xnor U4152 (N_4152,N_3703,N_3673);
or U4153 (N_4153,N_3607,N_3808);
nand U4154 (N_4154,N_3735,N_3746);
and U4155 (N_4155,N_3898,N_3604);
or U4156 (N_4156,N_3736,N_3830);
nor U4157 (N_4157,N_3618,N_3777);
nor U4158 (N_4158,N_3642,N_3837);
or U4159 (N_4159,N_3681,N_3638);
xnor U4160 (N_4160,N_3612,N_3626);
nand U4161 (N_4161,N_3612,N_3726);
xnor U4162 (N_4162,N_3825,N_3642);
or U4163 (N_4163,N_3894,N_3624);
and U4164 (N_4164,N_3701,N_3712);
or U4165 (N_4165,N_3647,N_3707);
or U4166 (N_4166,N_3824,N_3896);
xnor U4167 (N_4167,N_3772,N_3608);
nor U4168 (N_4168,N_3864,N_3891);
and U4169 (N_4169,N_3700,N_3860);
and U4170 (N_4170,N_3863,N_3809);
nor U4171 (N_4171,N_3865,N_3622);
nor U4172 (N_4172,N_3638,N_3898);
xor U4173 (N_4173,N_3792,N_3706);
and U4174 (N_4174,N_3738,N_3645);
xnor U4175 (N_4175,N_3728,N_3674);
nand U4176 (N_4176,N_3661,N_3640);
or U4177 (N_4177,N_3790,N_3660);
xor U4178 (N_4178,N_3808,N_3864);
or U4179 (N_4179,N_3714,N_3671);
xor U4180 (N_4180,N_3849,N_3624);
and U4181 (N_4181,N_3677,N_3690);
and U4182 (N_4182,N_3643,N_3744);
or U4183 (N_4183,N_3714,N_3674);
nand U4184 (N_4184,N_3737,N_3806);
or U4185 (N_4185,N_3800,N_3696);
nand U4186 (N_4186,N_3780,N_3826);
nand U4187 (N_4187,N_3652,N_3837);
nand U4188 (N_4188,N_3819,N_3801);
nor U4189 (N_4189,N_3725,N_3864);
or U4190 (N_4190,N_3629,N_3621);
xor U4191 (N_4191,N_3738,N_3723);
and U4192 (N_4192,N_3640,N_3872);
nand U4193 (N_4193,N_3778,N_3708);
nand U4194 (N_4194,N_3625,N_3607);
xor U4195 (N_4195,N_3883,N_3854);
and U4196 (N_4196,N_3753,N_3741);
nor U4197 (N_4197,N_3692,N_3746);
or U4198 (N_4198,N_3878,N_3699);
nand U4199 (N_4199,N_3761,N_3657);
or U4200 (N_4200,N_4164,N_4086);
and U4201 (N_4201,N_3988,N_4010);
or U4202 (N_4202,N_3985,N_4171);
nand U4203 (N_4203,N_4078,N_4153);
xor U4204 (N_4204,N_3986,N_4187);
xnor U4205 (N_4205,N_4012,N_3946);
nor U4206 (N_4206,N_4109,N_4160);
or U4207 (N_4207,N_4099,N_3936);
and U4208 (N_4208,N_3980,N_3914);
xor U4209 (N_4209,N_4147,N_3996);
nor U4210 (N_4210,N_3927,N_3991);
nand U4211 (N_4211,N_4047,N_4169);
nor U4212 (N_4212,N_3962,N_4141);
or U4213 (N_4213,N_3906,N_4123);
or U4214 (N_4214,N_4031,N_4124);
xor U4215 (N_4215,N_4129,N_4046);
or U4216 (N_4216,N_4176,N_4155);
nand U4217 (N_4217,N_3965,N_4112);
and U4218 (N_4218,N_4040,N_3930);
and U4219 (N_4219,N_4000,N_3922);
nor U4220 (N_4220,N_3970,N_4103);
xnor U4221 (N_4221,N_4068,N_3903);
xnor U4222 (N_4222,N_3960,N_4023);
xor U4223 (N_4223,N_3944,N_4036);
or U4224 (N_4224,N_4179,N_4093);
or U4225 (N_4225,N_4158,N_3997);
nand U4226 (N_4226,N_3901,N_4077);
nand U4227 (N_4227,N_4064,N_4161);
nand U4228 (N_4228,N_4101,N_3933);
xnor U4229 (N_4229,N_4095,N_3918);
nand U4230 (N_4230,N_3984,N_4066);
nand U4231 (N_4231,N_4128,N_4126);
and U4232 (N_4232,N_4042,N_4178);
nand U4233 (N_4233,N_4087,N_4165);
nand U4234 (N_4234,N_4132,N_3932);
or U4235 (N_4235,N_4037,N_4032);
xor U4236 (N_4236,N_4117,N_3940);
or U4237 (N_4237,N_4048,N_4102);
and U4238 (N_4238,N_4092,N_4177);
xnor U4239 (N_4239,N_4044,N_4130);
nand U4240 (N_4240,N_4106,N_3998);
or U4241 (N_4241,N_3993,N_4009);
xnor U4242 (N_4242,N_4030,N_3941);
and U4243 (N_4243,N_3956,N_3967);
or U4244 (N_4244,N_4175,N_3913);
nand U4245 (N_4245,N_4020,N_4073);
nor U4246 (N_4246,N_4198,N_4060);
xor U4247 (N_4247,N_3911,N_3923);
nand U4248 (N_4248,N_4172,N_4082);
nor U4249 (N_4249,N_4071,N_3950);
nand U4250 (N_4250,N_4026,N_4001);
nand U4251 (N_4251,N_3969,N_3915);
and U4252 (N_4252,N_3939,N_3953);
nor U4253 (N_4253,N_4015,N_3972);
or U4254 (N_4254,N_4003,N_4049);
or U4255 (N_4255,N_4067,N_4136);
or U4256 (N_4256,N_3977,N_4024);
or U4257 (N_4257,N_4045,N_4055);
nand U4258 (N_4258,N_3921,N_4006);
or U4259 (N_4259,N_3912,N_3916);
and U4260 (N_4260,N_3904,N_4193);
nand U4261 (N_4261,N_4190,N_3924);
nand U4262 (N_4262,N_4008,N_4167);
and U4263 (N_4263,N_3968,N_4180);
nand U4264 (N_4264,N_4070,N_3943);
xor U4265 (N_4265,N_4054,N_4021);
or U4266 (N_4266,N_3961,N_3958);
xor U4267 (N_4267,N_4138,N_4182);
or U4268 (N_4268,N_4196,N_4168);
nor U4269 (N_4269,N_3917,N_3975);
and U4270 (N_4270,N_4051,N_3909);
nor U4271 (N_4271,N_4111,N_4125);
or U4272 (N_4272,N_3987,N_4083);
xnor U4273 (N_4273,N_3992,N_4140);
and U4274 (N_4274,N_4120,N_3971);
nand U4275 (N_4275,N_3928,N_4018);
nand U4276 (N_4276,N_3905,N_4137);
nand U4277 (N_4277,N_3900,N_4025);
or U4278 (N_4278,N_3908,N_4076);
or U4279 (N_4279,N_4186,N_4056);
nand U4280 (N_4280,N_4152,N_3907);
nor U4281 (N_4281,N_4097,N_4151);
nor U4282 (N_4282,N_3954,N_4121);
nand U4283 (N_4283,N_4184,N_4118);
nor U4284 (N_4284,N_3937,N_4189);
nor U4285 (N_4285,N_3948,N_4199);
or U4286 (N_4286,N_3920,N_4033);
nor U4287 (N_4287,N_3979,N_4094);
or U4288 (N_4288,N_3910,N_3999);
and U4289 (N_4289,N_4191,N_3959);
or U4290 (N_4290,N_3976,N_4100);
xnor U4291 (N_4291,N_4091,N_3951);
and U4292 (N_4292,N_4113,N_4127);
and U4293 (N_4293,N_4072,N_4063);
or U4294 (N_4294,N_4053,N_4080);
nor U4295 (N_4295,N_4107,N_4144);
nor U4296 (N_4296,N_4079,N_3949);
nand U4297 (N_4297,N_4074,N_4005);
nand U4298 (N_4298,N_4004,N_4002);
nor U4299 (N_4299,N_3963,N_4038);
nand U4300 (N_4300,N_4089,N_4156);
or U4301 (N_4301,N_3919,N_4085);
xnor U4302 (N_4302,N_4007,N_4110);
nand U4303 (N_4303,N_4016,N_4133);
xor U4304 (N_4304,N_4043,N_3925);
xnor U4305 (N_4305,N_3982,N_3938);
nand U4306 (N_4306,N_4084,N_4057);
and U4307 (N_4307,N_3934,N_4163);
xor U4308 (N_4308,N_4058,N_4149);
xnor U4309 (N_4309,N_4088,N_3957);
or U4310 (N_4310,N_3981,N_4134);
nor U4311 (N_4311,N_4122,N_3989);
or U4312 (N_4312,N_4108,N_4148);
nor U4313 (N_4313,N_4105,N_4062);
nand U4314 (N_4314,N_3994,N_4022);
or U4315 (N_4315,N_4013,N_4135);
nor U4316 (N_4316,N_4145,N_3978);
xnor U4317 (N_4317,N_3929,N_4131);
xor U4318 (N_4318,N_4029,N_3974);
or U4319 (N_4319,N_3942,N_4146);
xor U4320 (N_4320,N_3966,N_4096);
nand U4321 (N_4321,N_4185,N_4011);
xnor U4322 (N_4322,N_4017,N_4162);
or U4323 (N_4323,N_4061,N_4019);
or U4324 (N_4324,N_4081,N_4142);
nor U4325 (N_4325,N_4041,N_4065);
and U4326 (N_4326,N_4192,N_4143);
and U4327 (N_4327,N_4195,N_4039);
or U4328 (N_4328,N_3931,N_3947);
nor U4329 (N_4329,N_4028,N_3964);
nand U4330 (N_4330,N_4059,N_4027);
xnor U4331 (N_4331,N_3935,N_3955);
or U4332 (N_4332,N_3995,N_4114);
nor U4333 (N_4333,N_4188,N_4154);
or U4334 (N_4334,N_4035,N_4075);
nor U4335 (N_4335,N_3983,N_3973);
xor U4336 (N_4336,N_4116,N_4173);
xor U4337 (N_4337,N_4157,N_4194);
nor U4338 (N_4338,N_4150,N_4159);
nand U4339 (N_4339,N_4183,N_4197);
nand U4340 (N_4340,N_3945,N_3926);
or U4341 (N_4341,N_4174,N_4166);
and U4342 (N_4342,N_4115,N_4069);
or U4343 (N_4343,N_3952,N_4104);
nand U4344 (N_4344,N_4052,N_4034);
xor U4345 (N_4345,N_3990,N_4170);
xnor U4346 (N_4346,N_4181,N_4050);
xnor U4347 (N_4347,N_3902,N_4090);
nand U4348 (N_4348,N_4098,N_4139);
xor U4349 (N_4349,N_4119,N_4014);
nor U4350 (N_4350,N_3995,N_3907);
nand U4351 (N_4351,N_4152,N_4145);
nor U4352 (N_4352,N_4102,N_4002);
xor U4353 (N_4353,N_3968,N_4066);
xnor U4354 (N_4354,N_4137,N_4087);
xnor U4355 (N_4355,N_3971,N_4199);
nand U4356 (N_4356,N_4088,N_3962);
or U4357 (N_4357,N_4028,N_3959);
nor U4358 (N_4358,N_4148,N_4194);
and U4359 (N_4359,N_4133,N_4005);
and U4360 (N_4360,N_3944,N_4111);
nor U4361 (N_4361,N_4059,N_4045);
and U4362 (N_4362,N_4180,N_4046);
xnor U4363 (N_4363,N_3953,N_4068);
and U4364 (N_4364,N_4138,N_4048);
xnor U4365 (N_4365,N_3902,N_4050);
or U4366 (N_4366,N_4130,N_4005);
or U4367 (N_4367,N_3975,N_3943);
or U4368 (N_4368,N_4171,N_4133);
nor U4369 (N_4369,N_4109,N_4136);
or U4370 (N_4370,N_3910,N_3982);
nand U4371 (N_4371,N_3928,N_4024);
and U4372 (N_4372,N_4057,N_4124);
nand U4373 (N_4373,N_3915,N_4177);
or U4374 (N_4374,N_4168,N_4102);
or U4375 (N_4375,N_4071,N_4063);
or U4376 (N_4376,N_3950,N_4183);
nor U4377 (N_4377,N_4147,N_4001);
and U4378 (N_4378,N_4173,N_4137);
and U4379 (N_4379,N_3957,N_4041);
and U4380 (N_4380,N_3907,N_4147);
nand U4381 (N_4381,N_3972,N_4085);
nor U4382 (N_4382,N_4198,N_4137);
or U4383 (N_4383,N_3936,N_3929);
nand U4384 (N_4384,N_4104,N_4138);
nor U4385 (N_4385,N_4178,N_4166);
and U4386 (N_4386,N_4145,N_4068);
nand U4387 (N_4387,N_4167,N_4198);
nor U4388 (N_4388,N_4054,N_4033);
or U4389 (N_4389,N_3941,N_3916);
nor U4390 (N_4390,N_3962,N_3919);
xor U4391 (N_4391,N_3928,N_4109);
and U4392 (N_4392,N_4049,N_3923);
nand U4393 (N_4393,N_4134,N_4068);
and U4394 (N_4394,N_4034,N_4162);
or U4395 (N_4395,N_3931,N_4169);
and U4396 (N_4396,N_3903,N_4093);
nand U4397 (N_4397,N_4142,N_3981);
and U4398 (N_4398,N_4010,N_4143);
xnor U4399 (N_4399,N_3984,N_4091);
or U4400 (N_4400,N_4180,N_4107);
xnor U4401 (N_4401,N_3952,N_4049);
xnor U4402 (N_4402,N_4082,N_4173);
and U4403 (N_4403,N_3912,N_4141);
nand U4404 (N_4404,N_3967,N_3927);
or U4405 (N_4405,N_4134,N_3988);
nor U4406 (N_4406,N_4034,N_4091);
and U4407 (N_4407,N_3912,N_3954);
nand U4408 (N_4408,N_4189,N_4032);
nand U4409 (N_4409,N_4190,N_4075);
nand U4410 (N_4410,N_3921,N_4171);
xor U4411 (N_4411,N_3970,N_4184);
and U4412 (N_4412,N_3900,N_4021);
or U4413 (N_4413,N_4109,N_4173);
or U4414 (N_4414,N_4056,N_3913);
and U4415 (N_4415,N_4038,N_4021);
nand U4416 (N_4416,N_4156,N_3935);
xnor U4417 (N_4417,N_4147,N_3978);
nand U4418 (N_4418,N_4001,N_4178);
xor U4419 (N_4419,N_4120,N_4191);
and U4420 (N_4420,N_4141,N_4055);
xor U4421 (N_4421,N_3978,N_4101);
nor U4422 (N_4422,N_4022,N_3964);
nand U4423 (N_4423,N_4044,N_3973);
nor U4424 (N_4424,N_4181,N_3954);
nand U4425 (N_4425,N_4048,N_3995);
and U4426 (N_4426,N_3979,N_4028);
nor U4427 (N_4427,N_4052,N_4128);
xnor U4428 (N_4428,N_4024,N_4004);
xnor U4429 (N_4429,N_4178,N_4112);
nand U4430 (N_4430,N_4047,N_4178);
nand U4431 (N_4431,N_3932,N_4104);
nor U4432 (N_4432,N_3927,N_4068);
nand U4433 (N_4433,N_4127,N_4188);
nand U4434 (N_4434,N_4027,N_3962);
xnor U4435 (N_4435,N_3907,N_4168);
nand U4436 (N_4436,N_4062,N_3983);
nand U4437 (N_4437,N_3964,N_4040);
and U4438 (N_4438,N_3928,N_4081);
nand U4439 (N_4439,N_4059,N_4023);
and U4440 (N_4440,N_3914,N_3995);
xor U4441 (N_4441,N_4182,N_3980);
xnor U4442 (N_4442,N_3923,N_3984);
nor U4443 (N_4443,N_4127,N_4117);
nor U4444 (N_4444,N_4181,N_3943);
nor U4445 (N_4445,N_4002,N_4036);
or U4446 (N_4446,N_4145,N_4101);
nand U4447 (N_4447,N_4145,N_4003);
xnor U4448 (N_4448,N_4158,N_4032);
or U4449 (N_4449,N_4140,N_4024);
xor U4450 (N_4450,N_4123,N_4086);
or U4451 (N_4451,N_4183,N_4032);
xor U4452 (N_4452,N_3912,N_3923);
and U4453 (N_4453,N_4162,N_3964);
nor U4454 (N_4454,N_4157,N_4197);
and U4455 (N_4455,N_4028,N_3906);
nand U4456 (N_4456,N_3950,N_3907);
nand U4457 (N_4457,N_4146,N_4154);
or U4458 (N_4458,N_4037,N_4061);
nand U4459 (N_4459,N_4110,N_3957);
and U4460 (N_4460,N_4096,N_3984);
nand U4461 (N_4461,N_4067,N_4034);
or U4462 (N_4462,N_4000,N_4008);
nand U4463 (N_4463,N_4181,N_4163);
nand U4464 (N_4464,N_3946,N_4151);
or U4465 (N_4465,N_4185,N_4159);
or U4466 (N_4466,N_3998,N_4001);
and U4467 (N_4467,N_4165,N_4118);
xnor U4468 (N_4468,N_4068,N_4090);
xor U4469 (N_4469,N_3977,N_3982);
nor U4470 (N_4470,N_4031,N_4151);
xor U4471 (N_4471,N_3959,N_3962);
nor U4472 (N_4472,N_3995,N_4152);
and U4473 (N_4473,N_3928,N_4038);
nor U4474 (N_4474,N_4153,N_3937);
nor U4475 (N_4475,N_4161,N_4012);
or U4476 (N_4476,N_3907,N_3954);
nor U4477 (N_4477,N_4084,N_3998);
or U4478 (N_4478,N_4110,N_3933);
xor U4479 (N_4479,N_3951,N_4094);
or U4480 (N_4480,N_3966,N_4195);
nand U4481 (N_4481,N_3979,N_4038);
nand U4482 (N_4482,N_4012,N_4077);
xor U4483 (N_4483,N_4161,N_4199);
or U4484 (N_4484,N_3943,N_3974);
xnor U4485 (N_4485,N_4124,N_4081);
or U4486 (N_4486,N_4146,N_4135);
nand U4487 (N_4487,N_4044,N_3919);
xor U4488 (N_4488,N_3918,N_3912);
nor U4489 (N_4489,N_4103,N_4015);
nand U4490 (N_4490,N_4096,N_4184);
nor U4491 (N_4491,N_4130,N_3986);
nand U4492 (N_4492,N_4092,N_3936);
nand U4493 (N_4493,N_3984,N_3913);
or U4494 (N_4494,N_4021,N_4188);
or U4495 (N_4495,N_4000,N_3911);
and U4496 (N_4496,N_4187,N_4170);
or U4497 (N_4497,N_3963,N_3949);
or U4498 (N_4498,N_4035,N_4146);
xnor U4499 (N_4499,N_3943,N_4083);
or U4500 (N_4500,N_4308,N_4491);
and U4501 (N_4501,N_4313,N_4224);
or U4502 (N_4502,N_4211,N_4366);
nand U4503 (N_4503,N_4424,N_4471);
nand U4504 (N_4504,N_4437,N_4425);
nor U4505 (N_4505,N_4311,N_4417);
and U4506 (N_4506,N_4497,N_4247);
or U4507 (N_4507,N_4264,N_4396);
nor U4508 (N_4508,N_4287,N_4331);
nor U4509 (N_4509,N_4475,N_4484);
or U4510 (N_4510,N_4350,N_4406);
nor U4511 (N_4511,N_4261,N_4352);
and U4512 (N_4512,N_4305,N_4387);
and U4513 (N_4513,N_4429,N_4320);
or U4514 (N_4514,N_4339,N_4218);
nor U4515 (N_4515,N_4451,N_4421);
and U4516 (N_4516,N_4299,N_4277);
xor U4517 (N_4517,N_4498,N_4363);
or U4518 (N_4518,N_4215,N_4259);
and U4519 (N_4519,N_4276,N_4252);
xor U4520 (N_4520,N_4342,N_4416);
nor U4521 (N_4521,N_4370,N_4435);
or U4522 (N_4522,N_4434,N_4426);
xor U4523 (N_4523,N_4258,N_4253);
or U4524 (N_4524,N_4405,N_4336);
or U4525 (N_4525,N_4290,N_4280);
xor U4526 (N_4526,N_4457,N_4244);
and U4527 (N_4527,N_4479,N_4268);
nor U4528 (N_4528,N_4213,N_4292);
nor U4529 (N_4529,N_4327,N_4481);
xor U4530 (N_4530,N_4375,N_4458);
and U4531 (N_4531,N_4409,N_4205);
or U4532 (N_4532,N_4315,N_4372);
or U4533 (N_4533,N_4303,N_4289);
xor U4534 (N_4534,N_4222,N_4419);
and U4535 (N_4535,N_4265,N_4376);
or U4536 (N_4536,N_4369,N_4354);
nand U4537 (N_4537,N_4243,N_4230);
nand U4538 (N_4538,N_4249,N_4492);
and U4539 (N_4539,N_4499,N_4441);
and U4540 (N_4540,N_4464,N_4490);
nor U4541 (N_4541,N_4494,N_4486);
or U4542 (N_4542,N_4422,N_4487);
nor U4543 (N_4543,N_4496,N_4242);
nor U4544 (N_4544,N_4225,N_4488);
or U4545 (N_4545,N_4465,N_4201);
nor U4546 (N_4546,N_4220,N_4232);
or U4547 (N_4547,N_4233,N_4389);
and U4548 (N_4548,N_4383,N_4365);
nand U4549 (N_4549,N_4391,N_4355);
or U4550 (N_4550,N_4361,N_4228);
xnor U4551 (N_4551,N_4283,N_4351);
xor U4552 (N_4552,N_4410,N_4467);
or U4553 (N_4553,N_4238,N_4343);
or U4554 (N_4554,N_4284,N_4325);
nor U4555 (N_4555,N_4371,N_4411);
nor U4556 (N_4556,N_4399,N_4209);
xor U4557 (N_4557,N_4239,N_4278);
or U4558 (N_4558,N_4346,N_4381);
xor U4559 (N_4559,N_4227,N_4468);
xor U4560 (N_4560,N_4357,N_4200);
xnor U4561 (N_4561,N_4374,N_4377);
nand U4562 (N_4562,N_4384,N_4348);
xor U4563 (N_4563,N_4314,N_4217);
nand U4564 (N_4564,N_4310,N_4340);
xor U4565 (N_4565,N_4447,N_4293);
xnor U4566 (N_4566,N_4203,N_4415);
or U4567 (N_4567,N_4295,N_4245);
and U4568 (N_4568,N_4248,N_4250);
and U4569 (N_4569,N_4380,N_4237);
nor U4570 (N_4570,N_4246,N_4298);
nor U4571 (N_4571,N_4466,N_4291);
xnor U4572 (N_4572,N_4463,N_4221);
nand U4573 (N_4573,N_4347,N_4312);
nor U4574 (N_4574,N_4286,N_4482);
nor U4575 (N_4575,N_4439,N_4260);
nand U4576 (N_4576,N_4328,N_4378);
xnor U4577 (N_4577,N_4418,N_4300);
or U4578 (N_4578,N_4321,N_4279);
xor U4579 (N_4579,N_4229,N_4404);
nand U4580 (N_4580,N_4386,N_4207);
nor U4581 (N_4581,N_4493,N_4401);
and U4582 (N_4582,N_4449,N_4373);
and U4583 (N_4583,N_4296,N_4433);
and U4584 (N_4584,N_4345,N_4359);
xor U4585 (N_4585,N_4453,N_4270);
and U4586 (N_4586,N_4263,N_4271);
or U4587 (N_4587,N_4362,N_4480);
nand U4588 (N_4588,N_4403,N_4326);
nor U4589 (N_4589,N_4323,N_4256);
or U4590 (N_4590,N_4335,N_4334);
or U4591 (N_4591,N_4316,N_4208);
nor U4592 (N_4592,N_4317,N_4304);
nand U4593 (N_4593,N_4294,N_4414);
or U4594 (N_4594,N_4428,N_4319);
and U4595 (N_4595,N_4269,N_4413);
nor U4596 (N_4596,N_4382,N_4454);
nand U4597 (N_4597,N_4450,N_4202);
nor U4598 (N_4598,N_4322,N_4367);
or U4599 (N_4599,N_4459,N_4306);
nand U4600 (N_4600,N_4204,N_4431);
xor U4601 (N_4601,N_4407,N_4379);
nand U4602 (N_4602,N_4338,N_4456);
and U4603 (N_4603,N_4356,N_4332);
nand U4604 (N_4604,N_4318,N_4273);
nor U4605 (N_4605,N_4251,N_4432);
or U4606 (N_4606,N_4223,N_4309);
nand U4607 (N_4607,N_4473,N_4255);
nor U4608 (N_4608,N_4333,N_4324);
or U4609 (N_4609,N_4329,N_4281);
or U4610 (N_4610,N_4274,N_4427);
nor U4611 (N_4611,N_4272,N_4443);
or U4612 (N_4612,N_4330,N_4349);
xnor U4613 (N_4613,N_4344,N_4301);
nand U4614 (N_4614,N_4282,N_4297);
nor U4615 (N_4615,N_4236,N_4240);
nand U4616 (N_4616,N_4397,N_4455);
nor U4617 (N_4617,N_4393,N_4469);
xor U4618 (N_4618,N_4388,N_4302);
nor U4619 (N_4619,N_4241,N_4485);
nor U4620 (N_4620,N_4438,N_4254);
xnor U4621 (N_4621,N_4219,N_4235);
xnor U4622 (N_4622,N_4275,N_4266);
and U4623 (N_4623,N_4390,N_4470);
xnor U4624 (N_4624,N_4412,N_4436);
nor U4625 (N_4625,N_4216,N_4420);
nand U4626 (N_4626,N_4400,N_4267);
xor U4627 (N_4627,N_4364,N_4226);
and U4628 (N_4628,N_4307,N_4408);
nor U4629 (N_4629,N_4210,N_4489);
nor U4630 (N_4630,N_4353,N_4442);
nand U4631 (N_4631,N_4460,N_4337);
nor U4632 (N_4632,N_4445,N_4392);
nor U4633 (N_4633,N_4368,N_4478);
nor U4634 (N_4634,N_4444,N_4212);
nor U4635 (N_4635,N_4395,N_4234);
and U4636 (N_4636,N_4360,N_4257);
nor U4637 (N_4637,N_4448,N_4452);
nor U4638 (N_4638,N_4495,N_4385);
nand U4639 (N_4639,N_4423,N_4440);
and U4640 (N_4640,N_4288,N_4214);
nand U4641 (N_4641,N_4430,N_4477);
nand U4642 (N_4642,N_4341,N_4358);
or U4643 (N_4643,N_4394,N_4461);
and U4644 (N_4644,N_4398,N_4206);
or U4645 (N_4645,N_4474,N_4231);
xnor U4646 (N_4646,N_4483,N_4462);
and U4647 (N_4647,N_4262,N_4476);
xor U4648 (N_4648,N_4285,N_4402);
and U4649 (N_4649,N_4446,N_4472);
nand U4650 (N_4650,N_4444,N_4221);
or U4651 (N_4651,N_4239,N_4487);
or U4652 (N_4652,N_4253,N_4415);
or U4653 (N_4653,N_4311,N_4332);
and U4654 (N_4654,N_4248,N_4312);
xnor U4655 (N_4655,N_4359,N_4351);
and U4656 (N_4656,N_4281,N_4258);
and U4657 (N_4657,N_4264,N_4303);
xor U4658 (N_4658,N_4335,N_4435);
nand U4659 (N_4659,N_4236,N_4388);
and U4660 (N_4660,N_4436,N_4434);
or U4661 (N_4661,N_4283,N_4336);
nand U4662 (N_4662,N_4354,N_4370);
xnor U4663 (N_4663,N_4261,N_4331);
nand U4664 (N_4664,N_4429,N_4316);
or U4665 (N_4665,N_4262,N_4371);
xnor U4666 (N_4666,N_4437,N_4404);
xnor U4667 (N_4667,N_4481,N_4208);
nand U4668 (N_4668,N_4355,N_4372);
nor U4669 (N_4669,N_4271,N_4369);
nor U4670 (N_4670,N_4267,N_4332);
nand U4671 (N_4671,N_4280,N_4420);
and U4672 (N_4672,N_4256,N_4245);
xor U4673 (N_4673,N_4268,N_4462);
xnor U4674 (N_4674,N_4329,N_4235);
nor U4675 (N_4675,N_4460,N_4260);
and U4676 (N_4676,N_4478,N_4480);
or U4677 (N_4677,N_4495,N_4451);
and U4678 (N_4678,N_4219,N_4327);
xnor U4679 (N_4679,N_4281,N_4225);
nor U4680 (N_4680,N_4468,N_4456);
and U4681 (N_4681,N_4352,N_4495);
nor U4682 (N_4682,N_4431,N_4472);
xor U4683 (N_4683,N_4243,N_4270);
nor U4684 (N_4684,N_4272,N_4473);
or U4685 (N_4685,N_4470,N_4226);
nor U4686 (N_4686,N_4379,N_4351);
and U4687 (N_4687,N_4370,N_4252);
or U4688 (N_4688,N_4405,N_4329);
or U4689 (N_4689,N_4432,N_4215);
and U4690 (N_4690,N_4335,N_4386);
and U4691 (N_4691,N_4408,N_4233);
nor U4692 (N_4692,N_4431,N_4325);
or U4693 (N_4693,N_4234,N_4411);
or U4694 (N_4694,N_4493,N_4216);
and U4695 (N_4695,N_4445,N_4326);
xor U4696 (N_4696,N_4412,N_4273);
and U4697 (N_4697,N_4312,N_4472);
and U4698 (N_4698,N_4387,N_4258);
nand U4699 (N_4699,N_4212,N_4441);
xnor U4700 (N_4700,N_4484,N_4433);
and U4701 (N_4701,N_4396,N_4209);
nor U4702 (N_4702,N_4268,N_4468);
nor U4703 (N_4703,N_4404,N_4334);
and U4704 (N_4704,N_4410,N_4251);
or U4705 (N_4705,N_4351,N_4428);
nor U4706 (N_4706,N_4203,N_4244);
nor U4707 (N_4707,N_4409,N_4343);
and U4708 (N_4708,N_4394,N_4294);
nor U4709 (N_4709,N_4480,N_4319);
or U4710 (N_4710,N_4369,N_4490);
xnor U4711 (N_4711,N_4411,N_4255);
and U4712 (N_4712,N_4304,N_4416);
xnor U4713 (N_4713,N_4287,N_4489);
nand U4714 (N_4714,N_4483,N_4437);
xnor U4715 (N_4715,N_4455,N_4200);
or U4716 (N_4716,N_4298,N_4371);
xor U4717 (N_4717,N_4243,N_4227);
nor U4718 (N_4718,N_4389,N_4265);
and U4719 (N_4719,N_4317,N_4286);
nor U4720 (N_4720,N_4497,N_4204);
xnor U4721 (N_4721,N_4450,N_4260);
nand U4722 (N_4722,N_4327,N_4357);
nor U4723 (N_4723,N_4405,N_4234);
nor U4724 (N_4724,N_4242,N_4378);
and U4725 (N_4725,N_4248,N_4388);
nor U4726 (N_4726,N_4326,N_4461);
and U4727 (N_4727,N_4499,N_4227);
or U4728 (N_4728,N_4299,N_4216);
or U4729 (N_4729,N_4204,N_4323);
nand U4730 (N_4730,N_4367,N_4223);
xnor U4731 (N_4731,N_4289,N_4207);
or U4732 (N_4732,N_4405,N_4413);
and U4733 (N_4733,N_4324,N_4417);
or U4734 (N_4734,N_4329,N_4280);
nor U4735 (N_4735,N_4434,N_4379);
nor U4736 (N_4736,N_4443,N_4417);
xor U4737 (N_4737,N_4347,N_4355);
xnor U4738 (N_4738,N_4461,N_4210);
nor U4739 (N_4739,N_4346,N_4430);
nand U4740 (N_4740,N_4254,N_4323);
xnor U4741 (N_4741,N_4321,N_4344);
and U4742 (N_4742,N_4287,N_4393);
or U4743 (N_4743,N_4394,N_4341);
xnor U4744 (N_4744,N_4456,N_4274);
nor U4745 (N_4745,N_4238,N_4383);
and U4746 (N_4746,N_4287,N_4365);
nor U4747 (N_4747,N_4208,N_4292);
or U4748 (N_4748,N_4304,N_4490);
nand U4749 (N_4749,N_4375,N_4235);
or U4750 (N_4750,N_4396,N_4308);
xor U4751 (N_4751,N_4360,N_4280);
and U4752 (N_4752,N_4469,N_4317);
nor U4753 (N_4753,N_4264,N_4440);
and U4754 (N_4754,N_4205,N_4449);
or U4755 (N_4755,N_4392,N_4438);
xnor U4756 (N_4756,N_4366,N_4434);
nand U4757 (N_4757,N_4231,N_4336);
xnor U4758 (N_4758,N_4388,N_4415);
nor U4759 (N_4759,N_4330,N_4246);
nor U4760 (N_4760,N_4273,N_4217);
nor U4761 (N_4761,N_4227,N_4457);
nand U4762 (N_4762,N_4262,N_4474);
or U4763 (N_4763,N_4325,N_4329);
nor U4764 (N_4764,N_4398,N_4458);
and U4765 (N_4765,N_4350,N_4480);
or U4766 (N_4766,N_4494,N_4475);
xor U4767 (N_4767,N_4401,N_4254);
or U4768 (N_4768,N_4304,N_4389);
or U4769 (N_4769,N_4418,N_4205);
nor U4770 (N_4770,N_4375,N_4204);
nor U4771 (N_4771,N_4325,N_4236);
and U4772 (N_4772,N_4291,N_4313);
or U4773 (N_4773,N_4286,N_4204);
nor U4774 (N_4774,N_4240,N_4216);
nor U4775 (N_4775,N_4313,N_4231);
and U4776 (N_4776,N_4259,N_4385);
or U4777 (N_4777,N_4381,N_4282);
and U4778 (N_4778,N_4399,N_4233);
or U4779 (N_4779,N_4462,N_4439);
nor U4780 (N_4780,N_4390,N_4409);
nand U4781 (N_4781,N_4237,N_4294);
or U4782 (N_4782,N_4337,N_4423);
or U4783 (N_4783,N_4494,N_4247);
xnor U4784 (N_4784,N_4295,N_4296);
nor U4785 (N_4785,N_4242,N_4418);
xnor U4786 (N_4786,N_4391,N_4419);
xnor U4787 (N_4787,N_4219,N_4378);
xor U4788 (N_4788,N_4380,N_4434);
nor U4789 (N_4789,N_4316,N_4278);
or U4790 (N_4790,N_4251,N_4319);
xor U4791 (N_4791,N_4449,N_4278);
nand U4792 (N_4792,N_4484,N_4201);
xnor U4793 (N_4793,N_4211,N_4233);
xor U4794 (N_4794,N_4377,N_4463);
or U4795 (N_4795,N_4219,N_4418);
or U4796 (N_4796,N_4405,N_4463);
or U4797 (N_4797,N_4432,N_4271);
or U4798 (N_4798,N_4211,N_4358);
xor U4799 (N_4799,N_4444,N_4490);
xnor U4800 (N_4800,N_4534,N_4685);
and U4801 (N_4801,N_4693,N_4708);
nand U4802 (N_4802,N_4625,N_4697);
nand U4803 (N_4803,N_4690,N_4672);
or U4804 (N_4804,N_4681,N_4595);
or U4805 (N_4805,N_4547,N_4719);
nand U4806 (N_4806,N_4639,N_4557);
nor U4807 (N_4807,N_4715,N_4751);
nor U4808 (N_4808,N_4793,N_4781);
nand U4809 (N_4809,N_4515,N_4579);
xnor U4810 (N_4810,N_4501,N_4775);
and U4811 (N_4811,N_4658,N_4559);
or U4812 (N_4812,N_4790,N_4524);
nor U4813 (N_4813,N_4759,N_4680);
nor U4814 (N_4814,N_4592,N_4564);
and U4815 (N_4815,N_4603,N_4568);
xor U4816 (N_4816,N_4587,N_4606);
xor U4817 (N_4817,N_4567,N_4782);
xor U4818 (N_4818,N_4588,N_4598);
nand U4819 (N_4819,N_4504,N_4623);
and U4820 (N_4820,N_4632,N_4613);
or U4821 (N_4821,N_4666,N_4754);
xor U4822 (N_4822,N_4514,N_4582);
nand U4823 (N_4823,N_4783,N_4718);
nor U4824 (N_4824,N_4798,N_4714);
and U4825 (N_4825,N_4585,N_4669);
nand U4826 (N_4826,N_4502,N_4566);
and U4827 (N_4827,N_4704,N_4655);
xnor U4828 (N_4828,N_4521,N_4739);
and U4829 (N_4829,N_4744,N_4784);
and U4830 (N_4830,N_4539,N_4788);
or U4831 (N_4831,N_4540,N_4601);
nor U4832 (N_4832,N_4770,N_4622);
xor U4833 (N_4833,N_4667,N_4607);
xnor U4834 (N_4834,N_4648,N_4611);
nand U4835 (N_4835,N_4549,N_4701);
or U4836 (N_4836,N_4779,N_4619);
and U4837 (N_4837,N_4679,N_4767);
nand U4838 (N_4838,N_4555,N_4508);
nor U4839 (N_4839,N_4721,N_4505);
nand U4840 (N_4840,N_4794,N_4664);
or U4841 (N_4841,N_4691,N_4635);
or U4842 (N_4842,N_4795,N_4758);
xor U4843 (N_4843,N_4671,N_4734);
nand U4844 (N_4844,N_4736,N_4705);
and U4845 (N_4845,N_4551,N_4706);
and U4846 (N_4846,N_4563,N_4668);
nand U4847 (N_4847,N_4799,N_4774);
xnor U4848 (N_4848,N_4560,N_4516);
or U4849 (N_4849,N_4576,N_4604);
xnor U4850 (N_4850,N_4762,N_4626);
nand U4851 (N_4851,N_4730,N_4650);
xor U4852 (N_4852,N_4766,N_4609);
nor U4853 (N_4853,N_4546,N_4586);
nor U4854 (N_4854,N_4593,N_4649);
and U4855 (N_4855,N_4670,N_4776);
or U4856 (N_4856,N_4537,N_4677);
and U4857 (N_4857,N_4688,N_4631);
nor U4858 (N_4858,N_4642,N_4500);
or U4859 (N_4859,N_4533,N_4692);
or U4860 (N_4860,N_4634,N_4678);
nor U4861 (N_4861,N_4663,N_4591);
or U4862 (N_4862,N_4780,N_4536);
nand U4863 (N_4863,N_4528,N_4532);
or U4864 (N_4864,N_4789,N_4610);
nand U4865 (N_4865,N_4746,N_4657);
and U4866 (N_4866,N_4561,N_4600);
nor U4867 (N_4867,N_4565,N_4506);
nand U4868 (N_4868,N_4574,N_4627);
and U4869 (N_4869,N_4553,N_4689);
or U4870 (N_4870,N_4787,N_4525);
xor U4871 (N_4871,N_4519,N_4575);
and U4872 (N_4872,N_4589,N_4755);
or U4873 (N_4873,N_4662,N_4527);
xor U4874 (N_4874,N_4554,N_4723);
nor U4875 (N_4875,N_4531,N_4530);
and U4876 (N_4876,N_4583,N_4637);
nand U4877 (N_4877,N_4526,N_4659);
or U4878 (N_4878,N_4643,N_4696);
or U4879 (N_4879,N_4699,N_4520);
nand U4880 (N_4880,N_4511,N_4542);
and U4881 (N_4881,N_4602,N_4641);
or U4882 (N_4882,N_4713,N_4552);
nor U4883 (N_4883,N_4518,N_4791);
xnor U4884 (N_4884,N_4503,N_4687);
and U4885 (N_4885,N_4571,N_4737);
xor U4886 (N_4886,N_4673,N_4596);
nor U4887 (N_4887,N_4717,N_4578);
and U4888 (N_4888,N_4683,N_4640);
nor U4889 (N_4889,N_4763,N_4522);
nor U4890 (N_4890,N_4628,N_4653);
nor U4891 (N_4891,N_4614,N_4761);
and U4892 (N_4892,N_4535,N_4581);
xnor U4893 (N_4893,N_4517,N_4562);
and U4894 (N_4894,N_4616,N_4633);
xnor U4895 (N_4895,N_4550,N_4740);
xor U4896 (N_4896,N_4510,N_4726);
nor U4897 (N_4897,N_4572,N_4538);
nor U4898 (N_4898,N_4590,N_4753);
or U4899 (N_4899,N_4764,N_4700);
xnor U4900 (N_4900,N_4765,N_4772);
nand U4901 (N_4901,N_4577,N_4725);
or U4902 (N_4902,N_4695,N_4676);
xor U4903 (N_4903,N_4612,N_4644);
or U4904 (N_4904,N_4729,N_4752);
nand U4905 (N_4905,N_4728,N_4580);
or U4906 (N_4906,N_4727,N_4749);
and U4907 (N_4907,N_4636,N_4665);
xnor U4908 (N_4908,N_4722,N_4512);
xor U4909 (N_4909,N_4797,N_4656);
or U4910 (N_4910,N_4682,N_4594);
xor U4911 (N_4911,N_4748,N_4735);
and U4912 (N_4912,N_4777,N_4621);
nand U4913 (N_4913,N_4674,N_4652);
and U4914 (N_4914,N_4698,N_4620);
and U4915 (N_4915,N_4720,N_4545);
xnor U4916 (N_4916,N_4638,N_4778);
or U4917 (N_4917,N_4733,N_4742);
or U4918 (N_4918,N_4709,N_4757);
nand U4919 (N_4919,N_4741,N_4745);
or U4920 (N_4920,N_4711,N_4684);
or U4921 (N_4921,N_4768,N_4675);
nand U4922 (N_4922,N_4660,N_4686);
and U4923 (N_4923,N_4509,N_4584);
xnor U4924 (N_4924,N_4750,N_4646);
xor U4925 (N_4925,N_4716,N_4796);
xnor U4926 (N_4926,N_4556,N_4732);
nand U4927 (N_4927,N_4570,N_4786);
or U4928 (N_4928,N_4513,N_4615);
or U4929 (N_4929,N_4785,N_4773);
and U4930 (N_4930,N_4617,N_4792);
and U4931 (N_4931,N_4712,N_4573);
nand U4932 (N_4932,N_4703,N_4654);
nand U4933 (N_4933,N_4548,N_4624);
and U4934 (N_4934,N_4618,N_4661);
nor U4935 (N_4935,N_4541,N_4645);
or U4936 (N_4936,N_4569,N_4747);
nor U4937 (N_4937,N_4756,N_4651);
nor U4938 (N_4938,N_4529,N_4605);
or U4939 (N_4939,N_4523,N_4544);
nand U4940 (N_4940,N_4738,N_4630);
nand U4941 (N_4941,N_4731,N_4507);
or U4942 (N_4942,N_4743,N_4702);
and U4943 (N_4943,N_4724,N_4710);
xnor U4944 (N_4944,N_4608,N_4694);
or U4945 (N_4945,N_4707,N_4597);
xor U4946 (N_4946,N_4647,N_4629);
xnor U4947 (N_4947,N_4558,N_4543);
xor U4948 (N_4948,N_4769,N_4771);
nand U4949 (N_4949,N_4599,N_4760);
nand U4950 (N_4950,N_4563,N_4535);
nand U4951 (N_4951,N_4538,N_4599);
xnor U4952 (N_4952,N_4717,N_4545);
nand U4953 (N_4953,N_4745,N_4622);
and U4954 (N_4954,N_4545,N_4634);
xor U4955 (N_4955,N_4659,N_4576);
nand U4956 (N_4956,N_4550,N_4584);
nor U4957 (N_4957,N_4763,N_4685);
xnor U4958 (N_4958,N_4741,N_4786);
nor U4959 (N_4959,N_4741,N_4756);
and U4960 (N_4960,N_4548,N_4788);
or U4961 (N_4961,N_4699,N_4527);
or U4962 (N_4962,N_4523,N_4603);
xnor U4963 (N_4963,N_4695,N_4503);
or U4964 (N_4964,N_4572,N_4757);
xor U4965 (N_4965,N_4575,N_4616);
nor U4966 (N_4966,N_4601,N_4697);
and U4967 (N_4967,N_4732,N_4516);
and U4968 (N_4968,N_4673,N_4692);
nand U4969 (N_4969,N_4595,N_4754);
xnor U4970 (N_4970,N_4558,N_4606);
and U4971 (N_4971,N_4796,N_4569);
xnor U4972 (N_4972,N_4784,N_4611);
or U4973 (N_4973,N_4532,N_4615);
and U4974 (N_4974,N_4547,N_4784);
and U4975 (N_4975,N_4706,N_4518);
nand U4976 (N_4976,N_4611,N_4736);
nand U4977 (N_4977,N_4693,N_4779);
nor U4978 (N_4978,N_4586,N_4587);
and U4979 (N_4979,N_4584,N_4537);
nand U4980 (N_4980,N_4772,N_4663);
nor U4981 (N_4981,N_4729,N_4653);
and U4982 (N_4982,N_4525,N_4782);
or U4983 (N_4983,N_4665,N_4536);
or U4984 (N_4984,N_4653,N_4630);
nor U4985 (N_4985,N_4731,N_4753);
and U4986 (N_4986,N_4500,N_4666);
and U4987 (N_4987,N_4505,N_4699);
xnor U4988 (N_4988,N_4556,N_4522);
nor U4989 (N_4989,N_4597,N_4789);
nor U4990 (N_4990,N_4730,N_4663);
xnor U4991 (N_4991,N_4690,N_4567);
xnor U4992 (N_4992,N_4565,N_4611);
xor U4993 (N_4993,N_4632,N_4593);
nor U4994 (N_4994,N_4605,N_4779);
and U4995 (N_4995,N_4680,N_4670);
or U4996 (N_4996,N_4673,N_4774);
and U4997 (N_4997,N_4729,N_4538);
nor U4998 (N_4998,N_4531,N_4653);
xnor U4999 (N_4999,N_4792,N_4612);
nand U5000 (N_5000,N_4633,N_4760);
xnor U5001 (N_5001,N_4527,N_4748);
xor U5002 (N_5002,N_4698,N_4581);
nand U5003 (N_5003,N_4773,N_4616);
nand U5004 (N_5004,N_4786,N_4618);
xor U5005 (N_5005,N_4682,N_4652);
and U5006 (N_5006,N_4777,N_4544);
or U5007 (N_5007,N_4570,N_4564);
xnor U5008 (N_5008,N_4796,N_4508);
nor U5009 (N_5009,N_4598,N_4574);
nor U5010 (N_5010,N_4796,N_4711);
and U5011 (N_5011,N_4717,N_4603);
or U5012 (N_5012,N_4591,N_4587);
nand U5013 (N_5013,N_4600,N_4735);
or U5014 (N_5014,N_4711,N_4642);
xnor U5015 (N_5015,N_4547,N_4539);
and U5016 (N_5016,N_4681,N_4653);
nand U5017 (N_5017,N_4537,N_4771);
and U5018 (N_5018,N_4542,N_4505);
nand U5019 (N_5019,N_4790,N_4794);
nand U5020 (N_5020,N_4526,N_4756);
and U5021 (N_5021,N_4673,N_4750);
and U5022 (N_5022,N_4609,N_4749);
xor U5023 (N_5023,N_4614,N_4763);
and U5024 (N_5024,N_4519,N_4724);
nand U5025 (N_5025,N_4775,N_4750);
or U5026 (N_5026,N_4511,N_4732);
or U5027 (N_5027,N_4658,N_4715);
or U5028 (N_5028,N_4504,N_4759);
nor U5029 (N_5029,N_4639,N_4785);
or U5030 (N_5030,N_4787,N_4709);
nor U5031 (N_5031,N_4661,N_4522);
or U5032 (N_5032,N_4619,N_4792);
or U5033 (N_5033,N_4604,N_4618);
xor U5034 (N_5034,N_4532,N_4502);
nand U5035 (N_5035,N_4611,N_4723);
and U5036 (N_5036,N_4735,N_4730);
xor U5037 (N_5037,N_4571,N_4578);
xnor U5038 (N_5038,N_4684,N_4691);
nand U5039 (N_5039,N_4568,N_4656);
xnor U5040 (N_5040,N_4623,N_4572);
and U5041 (N_5041,N_4686,N_4538);
xnor U5042 (N_5042,N_4649,N_4797);
or U5043 (N_5043,N_4659,N_4586);
nor U5044 (N_5044,N_4598,N_4656);
nor U5045 (N_5045,N_4653,N_4611);
and U5046 (N_5046,N_4714,N_4553);
and U5047 (N_5047,N_4703,N_4538);
nor U5048 (N_5048,N_4747,N_4527);
nor U5049 (N_5049,N_4508,N_4659);
and U5050 (N_5050,N_4509,N_4524);
nand U5051 (N_5051,N_4565,N_4696);
and U5052 (N_5052,N_4577,N_4735);
and U5053 (N_5053,N_4547,N_4581);
xor U5054 (N_5054,N_4670,N_4609);
xnor U5055 (N_5055,N_4679,N_4556);
and U5056 (N_5056,N_4526,N_4653);
nor U5057 (N_5057,N_4589,N_4731);
or U5058 (N_5058,N_4726,N_4540);
or U5059 (N_5059,N_4688,N_4604);
nor U5060 (N_5060,N_4696,N_4547);
nand U5061 (N_5061,N_4780,N_4529);
nor U5062 (N_5062,N_4630,N_4522);
and U5063 (N_5063,N_4504,N_4605);
nor U5064 (N_5064,N_4758,N_4541);
and U5065 (N_5065,N_4780,N_4648);
and U5066 (N_5066,N_4510,N_4605);
and U5067 (N_5067,N_4582,N_4699);
xor U5068 (N_5068,N_4550,N_4742);
and U5069 (N_5069,N_4792,N_4519);
xnor U5070 (N_5070,N_4689,N_4750);
nand U5071 (N_5071,N_4627,N_4789);
nand U5072 (N_5072,N_4536,N_4639);
nor U5073 (N_5073,N_4693,N_4619);
and U5074 (N_5074,N_4575,N_4522);
nor U5075 (N_5075,N_4503,N_4524);
or U5076 (N_5076,N_4661,N_4595);
xnor U5077 (N_5077,N_4576,N_4760);
xnor U5078 (N_5078,N_4741,N_4513);
and U5079 (N_5079,N_4708,N_4738);
nor U5080 (N_5080,N_4619,N_4719);
xor U5081 (N_5081,N_4646,N_4707);
nor U5082 (N_5082,N_4548,N_4743);
and U5083 (N_5083,N_4556,N_4697);
xnor U5084 (N_5084,N_4583,N_4594);
nor U5085 (N_5085,N_4509,N_4709);
xor U5086 (N_5086,N_4760,N_4657);
xor U5087 (N_5087,N_4666,N_4633);
nand U5088 (N_5088,N_4772,N_4617);
and U5089 (N_5089,N_4607,N_4697);
nand U5090 (N_5090,N_4562,N_4504);
or U5091 (N_5091,N_4663,N_4704);
nor U5092 (N_5092,N_4502,N_4742);
xnor U5093 (N_5093,N_4754,N_4665);
or U5094 (N_5094,N_4589,N_4762);
nor U5095 (N_5095,N_4694,N_4515);
or U5096 (N_5096,N_4592,N_4644);
and U5097 (N_5097,N_4594,N_4674);
nand U5098 (N_5098,N_4516,N_4542);
or U5099 (N_5099,N_4592,N_4547);
nor U5100 (N_5100,N_5074,N_5077);
nand U5101 (N_5101,N_5017,N_4846);
nand U5102 (N_5102,N_4918,N_5049);
nand U5103 (N_5103,N_4830,N_4962);
and U5104 (N_5104,N_4915,N_4957);
nor U5105 (N_5105,N_4824,N_4862);
nand U5106 (N_5106,N_4959,N_5079);
xnor U5107 (N_5107,N_4840,N_4903);
and U5108 (N_5108,N_5054,N_4917);
nor U5109 (N_5109,N_4999,N_4889);
xnor U5110 (N_5110,N_4910,N_4946);
xnor U5111 (N_5111,N_4905,N_4863);
nand U5112 (N_5112,N_4857,N_5024);
xor U5113 (N_5113,N_4956,N_5072);
and U5114 (N_5114,N_4966,N_5053);
nand U5115 (N_5115,N_5001,N_4943);
and U5116 (N_5116,N_4833,N_4850);
nand U5117 (N_5117,N_4994,N_5010);
or U5118 (N_5118,N_4931,N_4950);
or U5119 (N_5119,N_4981,N_4842);
nor U5120 (N_5120,N_4835,N_5011);
nor U5121 (N_5121,N_4933,N_4961);
nand U5122 (N_5122,N_4995,N_5009);
nor U5123 (N_5123,N_4935,N_4834);
nor U5124 (N_5124,N_4924,N_4828);
and U5125 (N_5125,N_4942,N_4890);
and U5126 (N_5126,N_5086,N_4986);
or U5127 (N_5127,N_4870,N_5038);
nand U5128 (N_5128,N_5035,N_5060);
or U5129 (N_5129,N_4976,N_4851);
nor U5130 (N_5130,N_4822,N_4978);
and U5131 (N_5131,N_4940,N_4939);
nand U5132 (N_5132,N_4934,N_4896);
nor U5133 (N_5133,N_4888,N_4816);
or U5134 (N_5134,N_5094,N_4987);
and U5135 (N_5135,N_5045,N_4998);
or U5136 (N_5136,N_5099,N_4843);
nor U5137 (N_5137,N_5052,N_4877);
nand U5138 (N_5138,N_5082,N_4813);
and U5139 (N_5139,N_5044,N_4875);
or U5140 (N_5140,N_4895,N_4974);
xor U5141 (N_5141,N_4911,N_5055);
nand U5142 (N_5142,N_5020,N_5036);
or U5143 (N_5143,N_4847,N_4901);
xnor U5144 (N_5144,N_5098,N_4839);
or U5145 (N_5145,N_5061,N_5025);
or U5146 (N_5146,N_5034,N_4804);
xor U5147 (N_5147,N_5084,N_4990);
xnor U5148 (N_5148,N_4849,N_5093);
nand U5149 (N_5149,N_4874,N_4945);
or U5150 (N_5150,N_4982,N_4873);
or U5151 (N_5151,N_5090,N_5087);
nor U5152 (N_5152,N_5068,N_5051);
nor U5153 (N_5153,N_5069,N_4807);
and U5154 (N_5154,N_4867,N_4872);
nand U5155 (N_5155,N_5027,N_5008);
or U5156 (N_5156,N_4810,N_4805);
xnor U5157 (N_5157,N_5089,N_4853);
xor U5158 (N_5158,N_4930,N_5016);
nor U5159 (N_5159,N_4878,N_5056);
xnor U5160 (N_5160,N_4909,N_4988);
nor U5161 (N_5161,N_4936,N_4977);
and U5162 (N_5162,N_4891,N_4993);
xnor U5163 (N_5163,N_4967,N_4984);
and U5164 (N_5164,N_5019,N_5071);
xor U5165 (N_5165,N_4838,N_5062);
nand U5166 (N_5166,N_4894,N_5033);
xnor U5167 (N_5167,N_4815,N_4949);
and U5168 (N_5168,N_5064,N_4825);
nand U5169 (N_5169,N_5075,N_5050);
and U5170 (N_5170,N_4958,N_5004);
nand U5171 (N_5171,N_4937,N_4919);
and U5172 (N_5172,N_4941,N_5031);
nand U5173 (N_5173,N_5003,N_5088);
xnor U5174 (N_5174,N_4876,N_4973);
xor U5175 (N_5175,N_4811,N_4912);
nor U5176 (N_5176,N_4823,N_4968);
nand U5177 (N_5177,N_4951,N_5058);
nand U5178 (N_5178,N_4898,N_4860);
or U5179 (N_5179,N_4921,N_4837);
nand U5180 (N_5180,N_4971,N_4882);
or U5181 (N_5181,N_4831,N_4892);
and U5182 (N_5182,N_5012,N_4887);
or U5183 (N_5183,N_5037,N_4920);
or U5184 (N_5184,N_4858,N_4880);
or U5185 (N_5185,N_5000,N_4812);
nor U5186 (N_5186,N_4868,N_5096);
xor U5187 (N_5187,N_5039,N_5046);
nor U5188 (N_5188,N_5065,N_5091);
nor U5189 (N_5189,N_4806,N_4879);
nand U5190 (N_5190,N_4922,N_4829);
nor U5191 (N_5191,N_4929,N_5022);
or U5192 (N_5192,N_5070,N_4881);
nor U5193 (N_5193,N_5047,N_5083);
and U5194 (N_5194,N_4820,N_4826);
nand U5195 (N_5195,N_4827,N_5063);
nor U5196 (N_5196,N_4944,N_4844);
or U5197 (N_5197,N_5026,N_5030);
nor U5198 (N_5198,N_4983,N_5057);
xnor U5199 (N_5199,N_4989,N_4855);
xor U5200 (N_5200,N_4818,N_5028);
or U5201 (N_5201,N_4904,N_5013);
and U5202 (N_5202,N_4883,N_4801);
nor U5203 (N_5203,N_4819,N_5085);
xor U5204 (N_5204,N_4885,N_4817);
xnor U5205 (N_5205,N_4985,N_5092);
and U5206 (N_5206,N_5002,N_5097);
xor U5207 (N_5207,N_4928,N_5018);
or U5208 (N_5208,N_4996,N_5043);
nand U5209 (N_5209,N_5014,N_5067);
and U5210 (N_5210,N_4832,N_4803);
xnor U5211 (N_5211,N_4980,N_4865);
and U5212 (N_5212,N_4869,N_4852);
or U5213 (N_5213,N_4884,N_4927);
nand U5214 (N_5214,N_4965,N_4897);
or U5215 (N_5215,N_4900,N_4841);
nand U5216 (N_5216,N_4854,N_4969);
nand U5217 (N_5217,N_5006,N_4926);
xor U5218 (N_5218,N_4992,N_4953);
xnor U5219 (N_5219,N_5005,N_4845);
and U5220 (N_5220,N_5048,N_5041);
nand U5221 (N_5221,N_4906,N_5076);
nor U5222 (N_5222,N_4960,N_4932);
and U5223 (N_5223,N_4925,N_5029);
and U5224 (N_5224,N_5078,N_4899);
and U5225 (N_5225,N_4800,N_4997);
or U5226 (N_5226,N_4836,N_4979);
and U5227 (N_5227,N_4916,N_4893);
xor U5228 (N_5228,N_5015,N_4871);
and U5229 (N_5229,N_5032,N_4975);
xnor U5230 (N_5230,N_4814,N_4972);
or U5231 (N_5231,N_5095,N_4908);
nand U5232 (N_5232,N_4808,N_4802);
xor U5233 (N_5233,N_4864,N_5081);
and U5234 (N_5234,N_4991,N_5042);
nand U5235 (N_5235,N_4914,N_4964);
xor U5236 (N_5236,N_4955,N_4947);
or U5237 (N_5237,N_5080,N_4886);
and U5238 (N_5238,N_5007,N_5023);
nor U5239 (N_5239,N_4821,N_4970);
nand U5240 (N_5240,N_5059,N_5021);
nand U5241 (N_5241,N_4948,N_4809);
or U5242 (N_5242,N_4848,N_4866);
or U5243 (N_5243,N_4902,N_4923);
xnor U5244 (N_5244,N_4954,N_4856);
xnor U5245 (N_5245,N_4861,N_4859);
nand U5246 (N_5246,N_5073,N_4952);
nor U5247 (N_5247,N_4963,N_5040);
or U5248 (N_5248,N_4913,N_4907);
nor U5249 (N_5249,N_5066,N_4938);
xor U5250 (N_5250,N_5050,N_4939);
nand U5251 (N_5251,N_4918,N_4899);
xor U5252 (N_5252,N_5060,N_4878);
or U5253 (N_5253,N_4811,N_4859);
and U5254 (N_5254,N_5040,N_4969);
nand U5255 (N_5255,N_4862,N_4962);
xnor U5256 (N_5256,N_5063,N_4831);
or U5257 (N_5257,N_4979,N_4868);
nand U5258 (N_5258,N_5012,N_4928);
or U5259 (N_5259,N_4802,N_4814);
xor U5260 (N_5260,N_5095,N_5081);
or U5261 (N_5261,N_5036,N_5082);
or U5262 (N_5262,N_4877,N_4890);
and U5263 (N_5263,N_4984,N_4801);
nor U5264 (N_5264,N_5026,N_4866);
and U5265 (N_5265,N_4992,N_4824);
nand U5266 (N_5266,N_5075,N_5055);
or U5267 (N_5267,N_4934,N_4976);
xnor U5268 (N_5268,N_5051,N_4963);
or U5269 (N_5269,N_4991,N_4900);
nor U5270 (N_5270,N_4934,N_4820);
xnor U5271 (N_5271,N_5040,N_5054);
xnor U5272 (N_5272,N_5035,N_5037);
and U5273 (N_5273,N_5041,N_5097);
and U5274 (N_5274,N_4915,N_4823);
nor U5275 (N_5275,N_5040,N_4906);
or U5276 (N_5276,N_5089,N_4866);
nor U5277 (N_5277,N_5032,N_4993);
xor U5278 (N_5278,N_5013,N_5018);
nand U5279 (N_5279,N_5040,N_4938);
nand U5280 (N_5280,N_4952,N_4931);
nand U5281 (N_5281,N_4929,N_5095);
xor U5282 (N_5282,N_5063,N_4900);
nand U5283 (N_5283,N_5045,N_4856);
or U5284 (N_5284,N_4907,N_4850);
xor U5285 (N_5285,N_5014,N_4835);
or U5286 (N_5286,N_4845,N_5083);
nand U5287 (N_5287,N_4987,N_4820);
nand U5288 (N_5288,N_4838,N_4947);
nor U5289 (N_5289,N_4841,N_4964);
nor U5290 (N_5290,N_5003,N_5031);
nor U5291 (N_5291,N_5081,N_4821);
and U5292 (N_5292,N_4998,N_4923);
nand U5293 (N_5293,N_4818,N_4826);
xor U5294 (N_5294,N_4916,N_4941);
and U5295 (N_5295,N_5024,N_5055);
or U5296 (N_5296,N_5064,N_5011);
nor U5297 (N_5297,N_4909,N_4992);
nand U5298 (N_5298,N_5040,N_4979);
and U5299 (N_5299,N_5004,N_5073);
nand U5300 (N_5300,N_4841,N_4965);
nor U5301 (N_5301,N_5005,N_4831);
nand U5302 (N_5302,N_4826,N_4863);
nand U5303 (N_5303,N_4978,N_5036);
nand U5304 (N_5304,N_4946,N_4872);
or U5305 (N_5305,N_4913,N_4813);
or U5306 (N_5306,N_4955,N_5002);
xnor U5307 (N_5307,N_4997,N_4850);
and U5308 (N_5308,N_4889,N_5036);
and U5309 (N_5309,N_5069,N_4955);
xnor U5310 (N_5310,N_4802,N_4860);
nand U5311 (N_5311,N_4922,N_4892);
or U5312 (N_5312,N_5053,N_4935);
or U5313 (N_5313,N_4922,N_4946);
and U5314 (N_5314,N_4973,N_4980);
nor U5315 (N_5315,N_4906,N_4959);
and U5316 (N_5316,N_5087,N_5076);
nor U5317 (N_5317,N_4828,N_5043);
nor U5318 (N_5318,N_4962,N_4999);
nand U5319 (N_5319,N_4968,N_5083);
nand U5320 (N_5320,N_4977,N_4914);
nor U5321 (N_5321,N_4820,N_4839);
nor U5322 (N_5322,N_5012,N_5089);
or U5323 (N_5323,N_4868,N_4827);
or U5324 (N_5324,N_4920,N_4975);
xnor U5325 (N_5325,N_4935,N_4841);
xor U5326 (N_5326,N_5028,N_5031);
nor U5327 (N_5327,N_4856,N_5069);
nand U5328 (N_5328,N_4910,N_4985);
xor U5329 (N_5329,N_4983,N_5056);
nand U5330 (N_5330,N_4805,N_5011);
and U5331 (N_5331,N_4895,N_4800);
and U5332 (N_5332,N_5002,N_5070);
nand U5333 (N_5333,N_4941,N_5043);
nor U5334 (N_5334,N_5018,N_4946);
nand U5335 (N_5335,N_5011,N_4886);
and U5336 (N_5336,N_4853,N_4991);
xor U5337 (N_5337,N_5021,N_5017);
or U5338 (N_5338,N_4891,N_5072);
and U5339 (N_5339,N_4905,N_5074);
and U5340 (N_5340,N_4898,N_5092);
nor U5341 (N_5341,N_5077,N_5052);
xor U5342 (N_5342,N_5099,N_4904);
xnor U5343 (N_5343,N_4969,N_4858);
or U5344 (N_5344,N_4964,N_5038);
or U5345 (N_5345,N_5027,N_4946);
or U5346 (N_5346,N_4920,N_4831);
nand U5347 (N_5347,N_5090,N_4910);
and U5348 (N_5348,N_5079,N_4929);
xnor U5349 (N_5349,N_4903,N_4805);
or U5350 (N_5350,N_4929,N_4881);
nand U5351 (N_5351,N_4897,N_5076);
or U5352 (N_5352,N_4998,N_4889);
or U5353 (N_5353,N_4900,N_4921);
nand U5354 (N_5354,N_5049,N_5013);
or U5355 (N_5355,N_5011,N_5022);
or U5356 (N_5356,N_5007,N_5001);
and U5357 (N_5357,N_5016,N_5026);
and U5358 (N_5358,N_5078,N_4820);
nor U5359 (N_5359,N_5055,N_4903);
xor U5360 (N_5360,N_5067,N_5044);
and U5361 (N_5361,N_4808,N_4905);
or U5362 (N_5362,N_4874,N_4904);
nor U5363 (N_5363,N_5008,N_5062);
xor U5364 (N_5364,N_4952,N_5087);
xnor U5365 (N_5365,N_5074,N_4968);
and U5366 (N_5366,N_4991,N_4856);
and U5367 (N_5367,N_4882,N_5074);
nand U5368 (N_5368,N_4945,N_4989);
or U5369 (N_5369,N_4846,N_4831);
nor U5370 (N_5370,N_5081,N_4988);
or U5371 (N_5371,N_5063,N_4998);
and U5372 (N_5372,N_5068,N_4879);
nor U5373 (N_5373,N_4968,N_4876);
or U5374 (N_5374,N_4886,N_4892);
nand U5375 (N_5375,N_4868,N_4991);
xor U5376 (N_5376,N_4839,N_4815);
or U5377 (N_5377,N_4927,N_4892);
xor U5378 (N_5378,N_5096,N_4819);
xor U5379 (N_5379,N_4838,N_4908);
or U5380 (N_5380,N_4902,N_4956);
nand U5381 (N_5381,N_4916,N_4947);
nand U5382 (N_5382,N_5051,N_4891);
nor U5383 (N_5383,N_5097,N_4974);
and U5384 (N_5384,N_4893,N_4814);
and U5385 (N_5385,N_4942,N_5025);
xnor U5386 (N_5386,N_4959,N_4912);
nand U5387 (N_5387,N_4923,N_5028);
nand U5388 (N_5388,N_4964,N_4935);
and U5389 (N_5389,N_5078,N_4944);
and U5390 (N_5390,N_4822,N_4882);
xor U5391 (N_5391,N_4821,N_4938);
nor U5392 (N_5392,N_4915,N_4849);
xnor U5393 (N_5393,N_4981,N_5038);
or U5394 (N_5394,N_5010,N_4989);
nor U5395 (N_5395,N_4940,N_4977);
and U5396 (N_5396,N_5096,N_4890);
nor U5397 (N_5397,N_4878,N_5021);
nand U5398 (N_5398,N_4985,N_5087);
xnor U5399 (N_5399,N_5097,N_4889);
xnor U5400 (N_5400,N_5168,N_5355);
nor U5401 (N_5401,N_5216,N_5154);
nor U5402 (N_5402,N_5156,N_5311);
nand U5403 (N_5403,N_5342,N_5368);
or U5404 (N_5404,N_5345,N_5150);
nand U5405 (N_5405,N_5143,N_5267);
xor U5406 (N_5406,N_5176,N_5278);
and U5407 (N_5407,N_5155,N_5292);
nand U5408 (N_5408,N_5268,N_5190);
xnor U5409 (N_5409,N_5281,N_5398);
xnor U5410 (N_5410,N_5274,N_5104);
xor U5411 (N_5411,N_5175,N_5298);
and U5412 (N_5412,N_5257,N_5297);
nand U5413 (N_5413,N_5126,N_5111);
nand U5414 (N_5414,N_5350,N_5386);
or U5415 (N_5415,N_5220,N_5204);
or U5416 (N_5416,N_5137,N_5361);
xor U5417 (N_5417,N_5210,N_5151);
and U5418 (N_5418,N_5337,N_5128);
xnor U5419 (N_5419,N_5189,N_5166);
or U5420 (N_5420,N_5142,N_5282);
xnor U5421 (N_5421,N_5197,N_5365);
or U5422 (N_5422,N_5188,N_5160);
nor U5423 (N_5423,N_5254,N_5370);
xor U5424 (N_5424,N_5113,N_5163);
nand U5425 (N_5425,N_5314,N_5325);
or U5426 (N_5426,N_5146,N_5393);
or U5427 (N_5427,N_5182,N_5385);
nor U5428 (N_5428,N_5346,N_5193);
xnor U5429 (N_5429,N_5273,N_5114);
or U5430 (N_5430,N_5392,N_5328);
nor U5431 (N_5431,N_5223,N_5148);
xor U5432 (N_5432,N_5103,N_5159);
or U5433 (N_5433,N_5318,N_5131);
nand U5434 (N_5434,N_5366,N_5394);
nor U5435 (N_5435,N_5222,N_5358);
and U5436 (N_5436,N_5390,N_5121);
xnor U5437 (N_5437,N_5240,N_5119);
or U5438 (N_5438,N_5315,N_5161);
and U5439 (N_5439,N_5213,N_5312);
nand U5440 (N_5440,N_5229,N_5141);
nand U5441 (N_5441,N_5139,N_5324);
and U5442 (N_5442,N_5209,N_5158);
nand U5443 (N_5443,N_5225,N_5250);
nand U5444 (N_5444,N_5291,N_5124);
nor U5445 (N_5445,N_5236,N_5301);
nand U5446 (N_5446,N_5299,N_5226);
nand U5447 (N_5447,N_5391,N_5251);
xnor U5448 (N_5448,N_5224,N_5264);
xnor U5449 (N_5449,N_5347,N_5302);
xor U5450 (N_5450,N_5169,N_5271);
nand U5451 (N_5451,N_5107,N_5349);
and U5452 (N_5452,N_5330,N_5186);
xnor U5453 (N_5453,N_5245,N_5164);
and U5454 (N_5454,N_5172,N_5375);
nor U5455 (N_5455,N_5363,N_5353);
nor U5456 (N_5456,N_5296,N_5332);
xor U5457 (N_5457,N_5183,N_5329);
and U5458 (N_5458,N_5322,N_5246);
or U5459 (N_5459,N_5259,N_5371);
xnor U5460 (N_5460,N_5389,N_5244);
nor U5461 (N_5461,N_5270,N_5201);
xnor U5462 (N_5462,N_5135,N_5351);
xnor U5463 (N_5463,N_5232,N_5374);
nand U5464 (N_5464,N_5369,N_5178);
xor U5465 (N_5465,N_5280,N_5293);
nor U5466 (N_5466,N_5202,N_5108);
nor U5467 (N_5467,N_5117,N_5106);
or U5468 (N_5468,N_5260,N_5290);
xor U5469 (N_5469,N_5344,N_5205);
xnor U5470 (N_5470,N_5272,N_5227);
or U5471 (N_5471,N_5147,N_5207);
nand U5472 (N_5472,N_5132,N_5321);
and U5473 (N_5473,N_5133,N_5287);
and U5474 (N_5474,N_5100,N_5253);
and U5475 (N_5475,N_5165,N_5115);
nor U5476 (N_5476,N_5170,N_5234);
and U5477 (N_5477,N_5383,N_5309);
xor U5478 (N_5478,N_5231,N_5249);
and U5479 (N_5479,N_5116,N_5294);
or U5480 (N_5480,N_5378,N_5360);
nand U5481 (N_5481,N_5179,N_5334);
xor U5482 (N_5482,N_5238,N_5211);
or U5483 (N_5483,N_5339,N_5110);
nand U5484 (N_5484,N_5194,N_5377);
and U5485 (N_5485,N_5379,N_5367);
and U5486 (N_5486,N_5313,N_5326);
nor U5487 (N_5487,N_5239,N_5228);
nor U5488 (N_5488,N_5295,N_5372);
and U5489 (N_5489,N_5208,N_5130);
and U5490 (N_5490,N_5275,N_5305);
and U5491 (N_5491,N_5215,N_5105);
and U5492 (N_5492,N_5219,N_5134);
or U5493 (N_5493,N_5196,N_5343);
xor U5494 (N_5494,N_5247,N_5102);
or U5495 (N_5495,N_5380,N_5283);
and U5496 (N_5496,N_5125,N_5187);
nor U5497 (N_5497,N_5206,N_5181);
nor U5498 (N_5498,N_5286,N_5340);
nand U5499 (N_5499,N_5396,N_5373);
or U5500 (N_5500,N_5306,N_5336);
xor U5501 (N_5501,N_5354,N_5387);
nor U5502 (N_5502,N_5303,N_5192);
and U5503 (N_5503,N_5256,N_5217);
and U5504 (N_5504,N_5269,N_5123);
nand U5505 (N_5505,N_5277,N_5284);
nor U5506 (N_5506,N_5191,N_5198);
and U5507 (N_5507,N_5352,N_5203);
xnor U5508 (N_5508,N_5320,N_5357);
nand U5509 (N_5509,N_5212,N_5288);
xnor U5510 (N_5510,N_5157,N_5289);
nor U5511 (N_5511,N_5112,N_5242);
nor U5512 (N_5512,N_5127,N_5258);
nand U5513 (N_5513,N_5397,N_5304);
and U5514 (N_5514,N_5279,N_5300);
nor U5515 (N_5515,N_5323,N_5265);
nor U5516 (N_5516,N_5307,N_5153);
or U5517 (N_5517,N_5162,N_5356);
nor U5518 (N_5518,N_5185,N_5152);
nand U5519 (N_5519,N_5180,N_5261);
or U5520 (N_5520,N_5214,N_5149);
nor U5521 (N_5521,N_5362,N_5248);
nand U5522 (N_5522,N_5140,N_5177);
nand U5523 (N_5523,N_5308,N_5262);
and U5524 (N_5524,N_5376,N_5171);
xor U5525 (N_5525,N_5120,N_5327);
xor U5526 (N_5526,N_5199,N_5381);
or U5527 (N_5527,N_5335,N_5319);
nand U5528 (N_5528,N_5136,N_5237);
xnor U5529 (N_5529,N_5266,N_5184);
or U5530 (N_5530,N_5109,N_5122);
and U5531 (N_5531,N_5399,N_5285);
or U5532 (N_5532,N_5241,N_5243);
and U5533 (N_5533,N_5359,N_5252);
and U5534 (N_5534,N_5101,N_5129);
nor U5535 (N_5535,N_5395,N_5333);
and U5536 (N_5536,N_5388,N_5331);
and U5537 (N_5537,N_5310,N_5276);
or U5538 (N_5538,N_5263,N_5145);
or U5539 (N_5539,N_5317,N_5221);
nand U5540 (N_5540,N_5167,N_5316);
or U5541 (N_5541,N_5173,N_5255);
nor U5542 (N_5542,N_5338,N_5138);
and U5543 (N_5543,N_5218,N_5174);
nand U5544 (N_5544,N_5348,N_5200);
nor U5545 (N_5545,N_5118,N_5233);
nor U5546 (N_5546,N_5144,N_5384);
and U5547 (N_5547,N_5382,N_5195);
or U5548 (N_5548,N_5230,N_5341);
and U5549 (N_5549,N_5364,N_5235);
xnor U5550 (N_5550,N_5157,N_5228);
xnor U5551 (N_5551,N_5365,N_5347);
or U5552 (N_5552,N_5126,N_5172);
or U5553 (N_5553,N_5223,N_5381);
xor U5554 (N_5554,N_5383,N_5124);
nand U5555 (N_5555,N_5237,N_5189);
xnor U5556 (N_5556,N_5188,N_5294);
xor U5557 (N_5557,N_5168,N_5357);
and U5558 (N_5558,N_5374,N_5306);
xnor U5559 (N_5559,N_5191,N_5363);
or U5560 (N_5560,N_5163,N_5245);
nor U5561 (N_5561,N_5365,N_5263);
nor U5562 (N_5562,N_5120,N_5316);
and U5563 (N_5563,N_5323,N_5331);
nand U5564 (N_5564,N_5397,N_5151);
nor U5565 (N_5565,N_5370,N_5192);
nor U5566 (N_5566,N_5287,N_5378);
and U5567 (N_5567,N_5158,N_5258);
xor U5568 (N_5568,N_5175,N_5317);
or U5569 (N_5569,N_5313,N_5142);
nor U5570 (N_5570,N_5327,N_5355);
or U5571 (N_5571,N_5116,N_5150);
or U5572 (N_5572,N_5138,N_5285);
nand U5573 (N_5573,N_5322,N_5297);
and U5574 (N_5574,N_5337,N_5361);
nor U5575 (N_5575,N_5247,N_5213);
nand U5576 (N_5576,N_5381,N_5191);
xor U5577 (N_5577,N_5160,N_5275);
and U5578 (N_5578,N_5170,N_5213);
or U5579 (N_5579,N_5369,N_5207);
nand U5580 (N_5580,N_5274,N_5180);
or U5581 (N_5581,N_5110,N_5293);
or U5582 (N_5582,N_5311,N_5302);
and U5583 (N_5583,N_5389,N_5259);
and U5584 (N_5584,N_5393,N_5269);
xnor U5585 (N_5585,N_5200,N_5367);
nand U5586 (N_5586,N_5380,N_5171);
nor U5587 (N_5587,N_5179,N_5109);
and U5588 (N_5588,N_5134,N_5175);
and U5589 (N_5589,N_5159,N_5168);
and U5590 (N_5590,N_5336,N_5240);
nor U5591 (N_5591,N_5199,N_5337);
nand U5592 (N_5592,N_5216,N_5329);
xor U5593 (N_5593,N_5377,N_5352);
nand U5594 (N_5594,N_5266,N_5173);
xor U5595 (N_5595,N_5388,N_5351);
nand U5596 (N_5596,N_5210,N_5261);
and U5597 (N_5597,N_5214,N_5324);
xor U5598 (N_5598,N_5268,N_5240);
or U5599 (N_5599,N_5188,N_5137);
nor U5600 (N_5600,N_5113,N_5307);
or U5601 (N_5601,N_5188,N_5375);
xnor U5602 (N_5602,N_5321,N_5229);
nor U5603 (N_5603,N_5329,N_5261);
nor U5604 (N_5604,N_5363,N_5344);
xnor U5605 (N_5605,N_5138,N_5383);
nand U5606 (N_5606,N_5147,N_5108);
nand U5607 (N_5607,N_5287,N_5302);
nand U5608 (N_5608,N_5134,N_5157);
or U5609 (N_5609,N_5113,N_5144);
nor U5610 (N_5610,N_5391,N_5109);
nand U5611 (N_5611,N_5385,N_5241);
xor U5612 (N_5612,N_5221,N_5358);
or U5613 (N_5613,N_5357,N_5176);
nand U5614 (N_5614,N_5353,N_5368);
nor U5615 (N_5615,N_5388,N_5116);
or U5616 (N_5616,N_5286,N_5250);
nor U5617 (N_5617,N_5341,N_5314);
nor U5618 (N_5618,N_5378,N_5256);
nor U5619 (N_5619,N_5295,N_5318);
and U5620 (N_5620,N_5239,N_5158);
nor U5621 (N_5621,N_5106,N_5257);
and U5622 (N_5622,N_5157,N_5105);
xnor U5623 (N_5623,N_5289,N_5334);
nor U5624 (N_5624,N_5273,N_5146);
nand U5625 (N_5625,N_5160,N_5334);
nand U5626 (N_5626,N_5194,N_5228);
or U5627 (N_5627,N_5168,N_5202);
nand U5628 (N_5628,N_5160,N_5330);
or U5629 (N_5629,N_5398,N_5246);
nor U5630 (N_5630,N_5278,N_5354);
xor U5631 (N_5631,N_5367,N_5347);
xor U5632 (N_5632,N_5104,N_5141);
xnor U5633 (N_5633,N_5166,N_5178);
xor U5634 (N_5634,N_5177,N_5307);
or U5635 (N_5635,N_5383,N_5371);
or U5636 (N_5636,N_5169,N_5177);
xor U5637 (N_5637,N_5197,N_5210);
nand U5638 (N_5638,N_5385,N_5230);
xor U5639 (N_5639,N_5189,N_5354);
nand U5640 (N_5640,N_5104,N_5225);
nor U5641 (N_5641,N_5233,N_5353);
or U5642 (N_5642,N_5291,N_5244);
and U5643 (N_5643,N_5109,N_5336);
xnor U5644 (N_5644,N_5133,N_5235);
nand U5645 (N_5645,N_5163,N_5179);
or U5646 (N_5646,N_5107,N_5194);
and U5647 (N_5647,N_5222,N_5283);
nor U5648 (N_5648,N_5321,N_5342);
nor U5649 (N_5649,N_5161,N_5115);
nor U5650 (N_5650,N_5309,N_5295);
and U5651 (N_5651,N_5199,N_5159);
nor U5652 (N_5652,N_5132,N_5319);
and U5653 (N_5653,N_5217,N_5331);
nor U5654 (N_5654,N_5125,N_5203);
and U5655 (N_5655,N_5184,N_5255);
or U5656 (N_5656,N_5259,N_5109);
and U5657 (N_5657,N_5259,N_5126);
or U5658 (N_5658,N_5375,N_5210);
nand U5659 (N_5659,N_5179,N_5237);
or U5660 (N_5660,N_5244,N_5153);
or U5661 (N_5661,N_5179,N_5155);
nand U5662 (N_5662,N_5129,N_5116);
or U5663 (N_5663,N_5360,N_5204);
nand U5664 (N_5664,N_5374,N_5299);
and U5665 (N_5665,N_5312,N_5393);
or U5666 (N_5666,N_5128,N_5260);
and U5667 (N_5667,N_5246,N_5116);
nor U5668 (N_5668,N_5355,N_5299);
nor U5669 (N_5669,N_5399,N_5140);
and U5670 (N_5670,N_5117,N_5394);
xnor U5671 (N_5671,N_5218,N_5123);
or U5672 (N_5672,N_5169,N_5355);
or U5673 (N_5673,N_5109,N_5173);
xnor U5674 (N_5674,N_5318,N_5188);
nor U5675 (N_5675,N_5266,N_5219);
or U5676 (N_5676,N_5148,N_5103);
and U5677 (N_5677,N_5222,N_5163);
nand U5678 (N_5678,N_5300,N_5241);
nor U5679 (N_5679,N_5110,N_5211);
or U5680 (N_5680,N_5169,N_5220);
and U5681 (N_5681,N_5108,N_5159);
xor U5682 (N_5682,N_5165,N_5325);
or U5683 (N_5683,N_5329,N_5375);
or U5684 (N_5684,N_5393,N_5246);
nor U5685 (N_5685,N_5120,N_5163);
or U5686 (N_5686,N_5149,N_5308);
nand U5687 (N_5687,N_5246,N_5138);
nor U5688 (N_5688,N_5153,N_5235);
and U5689 (N_5689,N_5394,N_5276);
nor U5690 (N_5690,N_5153,N_5320);
and U5691 (N_5691,N_5327,N_5148);
or U5692 (N_5692,N_5228,N_5395);
xnor U5693 (N_5693,N_5171,N_5101);
and U5694 (N_5694,N_5195,N_5123);
xnor U5695 (N_5695,N_5276,N_5337);
or U5696 (N_5696,N_5271,N_5301);
or U5697 (N_5697,N_5367,N_5305);
xor U5698 (N_5698,N_5113,N_5157);
xor U5699 (N_5699,N_5299,N_5315);
xor U5700 (N_5700,N_5440,N_5678);
and U5701 (N_5701,N_5614,N_5505);
xor U5702 (N_5702,N_5623,N_5500);
xnor U5703 (N_5703,N_5469,N_5599);
xnor U5704 (N_5704,N_5409,N_5687);
or U5705 (N_5705,N_5433,N_5400);
and U5706 (N_5706,N_5458,N_5693);
and U5707 (N_5707,N_5507,N_5629);
xor U5708 (N_5708,N_5624,N_5641);
nor U5709 (N_5709,N_5552,N_5424);
nand U5710 (N_5710,N_5631,N_5446);
xnor U5711 (N_5711,N_5537,N_5662);
and U5712 (N_5712,N_5546,N_5692);
and U5713 (N_5713,N_5575,N_5492);
nand U5714 (N_5714,N_5568,N_5444);
or U5715 (N_5715,N_5605,N_5561);
xnor U5716 (N_5716,N_5680,N_5612);
xnor U5717 (N_5717,N_5620,N_5659);
xnor U5718 (N_5718,N_5632,N_5633);
nor U5719 (N_5719,N_5661,N_5564);
xor U5720 (N_5720,N_5531,N_5472);
nor U5721 (N_5721,N_5423,N_5410);
and U5722 (N_5722,N_5617,N_5526);
nand U5723 (N_5723,N_5509,N_5562);
and U5724 (N_5724,N_5465,N_5411);
xor U5725 (N_5725,N_5412,N_5566);
nor U5726 (N_5726,N_5642,N_5443);
and U5727 (N_5727,N_5671,N_5518);
xnor U5728 (N_5728,N_5466,N_5688);
xnor U5729 (N_5729,N_5541,N_5570);
or U5730 (N_5730,N_5403,N_5674);
xnor U5731 (N_5731,N_5455,N_5666);
nand U5732 (N_5732,N_5499,N_5521);
or U5733 (N_5733,N_5598,N_5556);
and U5734 (N_5734,N_5407,N_5656);
and U5735 (N_5735,N_5585,N_5611);
xor U5736 (N_5736,N_5664,N_5698);
xnor U5737 (N_5737,N_5497,N_5544);
xnor U5738 (N_5738,N_5647,N_5595);
xnor U5739 (N_5739,N_5417,N_5580);
and U5740 (N_5740,N_5533,N_5447);
nor U5741 (N_5741,N_5451,N_5691);
xor U5742 (N_5742,N_5569,N_5559);
xor U5743 (N_5743,N_5622,N_5438);
nand U5744 (N_5744,N_5517,N_5578);
or U5745 (N_5745,N_5540,N_5405);
nor U5746 (N_5746,N_5439,N_5685);
nor U5747 (N_5747,N_5514,N_5450);
or U5748 (N_5748,N_5584,N_5426);
xor U5749 (N_5749,N_5606,N_5571);
nor U5750 (N_5750,N_5553,N_5592);
nand U5751 (N_5751,N_5463,N_5502);
and U5752 (N_5752,N_5532,N_5460);
or U5753 (N_5753,N_5689,N_5457);
or U5754 (N_5754,N_5496,N_5435);
nand U5755 (N_5755,N_5520,N_5652);
xor U5756 (N_5756,N_5513,N_5506);
and U5757 (N_5757,N_5486,N_5603);
and U5758 (N_5758,N_5525,N_5429);
nand U5759 (N_5759,N_5651,N_5485);
nand U5760 (N_5760,N_5468,N_5511);
or U5761 (N_5761,N_5697,N_5555);
xor U5762 (N_5762,N_5422,N_5655);
nand U5763 (N_5763,N_5473,N_5621);
or U5764 (N_5764,N_5418,N_5658);
nor U5765 (N_5765,N_5576,N_5660);
nor U5766 (N_5766,N_5483,N_5480);
xnor U5767 (N_5767,N_5510,N_5670);
and U5768 (N_5768,N_5588,N_5600);
nor U5769 (N_5769,N_5663,N_5625);
or U5770 (N_5770,N_5679,N_5668);
xnor U5771 (N_5771,N_5613,N_5653);
nand U5772 (N_5772,N_5536,N_5470);
nor U5773 (N_5773,N_5522,N_5610);
nand U5774 (N_5774,N_5650,N_5628);
or U5775 (N_5775,N_5638,N_5667);
and U5776 (N_5776,N_5547,N_5419);
nand U5777 (N_5777,N_5683,N_5452);
xor U5778 (N_5778,N_5459,N_5442);
nor U5779 (N_5779,N_5448,N_5487);
nor U5780 (N_5780,N_5649,N_5681);
and U5781 (N_5781,N_5574,N_5495);
nand U5782 (N_5782,N_5604,N_5626);
nor U5783 (N_5783,N_5437,N_5672);
or U5784 (N_5784,N_5609,N_5695);
or U5785 (N_5785,N_5669,N_5581);
and U5786 (N_5786,N_5528,N_5607);
nand U5787 (N_5787,N_5523,N_5636);
xor U5788 (N_5788,N_5456,N_5618);
nand U5789 (N_5789,N_5639,N_5476);
nor U5790 (N_5790,N_5503,N_5640);
or U5791 (N_5791,N_5535,N_5665);
nor U5792 (N_5792,N_5587,N_5579);
nand U5793 (N_5793,N_5589,N_5453);
nand U5794 (N_5794,N_5543,N_5551);
xor U5795 (N_5795,N_5696,N_5594);
and U5796 (N_5796,N_5413,N_5690);
nor U5797 (N_5797,N_5461,N_5432);
xor U5798 (N_5798,N_5637,N_5408);
or U5799 (N_5799,N_5644,N_5699);
nand U5800 (N_5800,N_5572,N_5482);
or U5801 (N_5801,N_5441,N_5449);
and U5802 (N_5802,N_5493,N_5591);
nand U5803 (N_5803,N_5530,N_5657);
nand U5804 (N_5804,N_5498,N_5554);
nor U5805 (N_5805,N_5560,N_5467);
nand U5806 (N_5806,N_5431,N_5445);
nor U5807 (N_5807,N_5421,N_5515);
and U5808 (N_5808,N_5434,N_5586);
or U5809 (N_5809,N_5645,N_5415);
or U5810 (N_5810,N_5558,N_5538);
or U5811 (N_5811,N_5406,N_5464);
and U5812 (N_5812,N_5542,N_5616);
and U5813 (N_5813,N_5627,N_5479);
nor U5814 (N_5814,N_5654,N_5501);
or U5815 (N_5815,N_5539,N_5549);
and U5816 (N_5816,N_5475,N_5488);
xnor U5817 (N_5817,N_5420,N_5694);
nor U5818 (N_5818,N_5436,N_5481);
nor U5819 (N_5819,N_5545,N_5430);
nor U5820 (N_5820,N_5677,N_5512);
nand U5821 (N_5821,N_5643,N_5471);
nand U5822 (N_5822,N_5489,N_5548);
or U5823 (N_5823,N_5401,N_5557);
nor U5824 (N_5824,N_5519,N_5648);
nor U5825 (N_5825,N_5478,N_5635);
nor U5826 (N_5826,N_5646,N_5524);
or U5827 (N_5827,N_5416,N_5615);
xor U5828 (N_5828,N_5504,N_5477);
or U5829 (N_5829,N_5563,N_5462);
or U5830 (N_5830,N_5404,N_5676);
nand U5831 (N_5831,N_5565,N_5474);
and U5832 (N_5832,N_5534,N_5428);
nand U5833 (N_5833,N_5583,N_5608);
nor U5834 (N_5834,N_5601,N_5550);
and U5835 (N_5835,N_5597,N_5516);
nor U5836 (N_5836,N_5527,N_5491);
xnor U5837 (N_5837,N_5454,N_5577);
nand U5838 (N_5838,N_5602,N_5682);
or U5839 (N_5839,N_5673,N_5686);
and U5840 (N_5840,N_5529,N_5427);
and U5841 (N_5841,N_5634,N_5402);
xnor U5842 (N_5842,N_5593,N_5573);
and U5843 (N_5843,N_5567,N_5590);
nand U5844 (N_5844,N_5596,N_5484);
nand U5845 (N_5845,N_5619,N_5494);
nor U5846 (N_5846,N_5414,N_5630);
nor U5847 (N_5847,N_5675,N_5508);
nand U5848 (N_5848,N_5684,N_5425);
xnor U5849 (N_5849,N_5490,N_5582);
nor U5850 (N_5850,N_5519,N_5679);
nand U5851 (N_5851,N_5685,N_5695);
xnor U5852 (N_5852,N_5652,N_5546);
or U5853 (N_5853,N_5669,N_5502);
nand U5854 (N_5854,N_5526,N_5508);
and U5855 (N_5855,N_5483,N_5532);
or U5856 (N_5856,N_5630,N_5509);
or U5857 (N_5857,N_5613,N_5572);
and U5858 (N_5858,N_5427,N_5425);
or U5859 (N_5859,N_5478,N_5440);
nand U5860 (N_5860,N_5617,N_5468);
nor U5861 (N_5861,N_5486,N_5500);
nor U5862 (N_5862,N_5477,N_5498);
and U5863 (N_5863,N_5423,N_5648);
nor U5864 (N_5864,N_5438,N_5557);
and U5865 (N_5865,N_5594,N_5412);
or U5866 (N_5866,N_5548,N_5430);
or U5867 (N_5867,N_5587,N_5601);
or U5868 (N_5868,N_5622,N_5620);
xor U5869 (N_5869,N_5617,N_5597);
xnor U5870 (N_5870,N_5523,N_5650);
xnor U5871 (N_5871,N_5436,N_5588);
nand U5872 (N_5872,N_5650,N_5577);
nor U5873 (N_5873,N_5696,N_5640);
nand U5874 (N_5874,N_5443,N_5404);
nand U5875 (N_5875,N_5627,N_5483);
xor U5876 (N_5876,N_5610,N_5645);
nor U5877 (N_5877,N_5449,N_5519);
nand U5878 (N_5878,N_5409,N_5533);
xor U5879 (N_5879,N_5676,N_5536);
xor U5880 (N_5880,N_5524,N_5448);
xor U5881 (N_5881,N_5506,N_5631);
and U5882 (N_5882,N_5462,N_5485);
nor U5883 (N_5883,N_5617,N_5670);
nand U5884 (N_5884,N_5684,N_5556);
xor U5885 (N_5885,N_5641,N_5433);
nand U5886 (N_5886,N_5566,N_5434);
or U5887 (N_5887,N_5537,N_5456);
nand U5888 (N_5888,N_5551,N_5550);
or U5889 (N_5889,N_5629,N_5662);
nand U5890 (N_5890,N_5427,N_5504);
xor U5891 (N_5891,N_5520,N_5432);
or U5892 (N_5892,N_5402,N_5596);
or U5893 (N_5893,N_5547,N_5433);
and U5894 (N_5894,N_5682,N_5657);
and U5895 (N_5895,N_5417,N_5693);
nand U5896 (N_5896,N_5689,N_5503);
nand U5897 (N_5897,N_5443,N_5520);
and U5898 (N_5898,N_5532,N_5494);
nand U5899 (N_5899,N_5572,N_5496);
nor U5900 (N_5900,N_5629,N_5436);
nor U5901 (N_5901,N_5495,N_5444);
or U5902 (N_5902,N_5691,N_5508);
or U5903 (N_5903,N_5693,N_5567);
xor U5904 (N_5904,N_5512,N_5470);
nor U5905 (N_5905,N_5473,N_5487);
nand U5906 (N_5906,N_5682,N_5473);
xnor U5907 (N_5907,N_5498,N_5518);
nand U5908 (N_5908,N_5416,N_5523);
nor U5909 (N_5909,N_5439,N_5646);
and U5910 (N_5910,N_5674,N_5428);
and U5911 (N_5911,N_5557,N_5608);
nand U5912 (N_5912,N_5643,N_5631);
nor U5913 (N_5913,N_5506,N_5487);
xor U5914 (N_5914,N_5692,N_5480);
nand U5915 (N_5915,N_5686,N_5594);
nor U5916 (N_5916,N_5546,N_5508);
nor U5917 (N_5917,N_5637,N_5641);
or U5918 (N_5918,N_5501,N_5577);
xnor U5919 (N_5919,N_5663,N_5570);
xor U5920 (N_5920,N_5477,N_5428);
nor U5921 (N_5921,N_5450,N_5684);
xnor U5922 (N_5922,N_5480,N_5468);
and U5923 (N_5923,N_5417,N_5466);
and U5924 (N_5924,N_5515,N_5542);
xor U5925 (N_5925,N_5651,N_5509);
nor U5926 (N_5926,N_5569,N_5581);
and U5927 (N_5927,N_5497,N_5523);
nor U5928 (N_5928,N_5465,N_5682);
xnor U5929 (N_5929,N_5559,N_5537);
xnor U5930 (N_5930,N_5526,N_5532);
xnor U5931 (N_5931,N_5515,N_5471);
nand U5932 (N_5932,N_5437,N_5421);
and U5933 (N_5933,N_5634,N_5428);
or U5934 (N_5934,N_5550,N_5489);
nor U5935 (N_5935,N_5518,N_5500);
and U5936 (N_5936,N_5432,N_5667);
nor U5937 (N_5937,N_5479,N_5527);
nand U5938 (N_5938,N_5592,N_5406);
nor U5939 (N_5939,N_5600,N_5638);
or U5940 (N_5940,N_5623,N_5481);
or U5941 (N_5941,N_5561,N_5579);
and U5942 (N_5942,N_5498,N_5450);
nand U5943 (N_5943,N_5592,N_5443);
xnor U5944 (N_5944,N_5437,N_5446);
xor U5945 (N_5945,N_5581,N_5610);
and U5946 (N_5946,N_5485,N_5471);
xnor U5947 (N_5947,N_5449,N_5489);
and U5948 (N_5948,N_5499,N_5667);
and U5949 (N_5949,N_5516,N_5654);
and U5950 (N_5950,N_5583,N_5603);
nor U5951 (N_5951,N_5659,N_5426);
nor U5952 (N_5952,N_5671,N_5500);
xnor U5953 (N_5953,N_5571,N_5553);
nor U5954 (N_5954,N_5694,N_5499);
nor U5955 (N_5955,N_5652,N_5502);
xor U5956 (N_5956,N_5666,N_5541);
xor U5957 (N_5957,N_5645,N_5684);
xnor U5958 (N_5958,N_5614,N_5543);
and U5959 (N_5959,N_5627,N_5695);
or U5960 (N_5960,N_5443,N_5503);
nand U5961 (N_5961,N_5620,N_5639);
xnor U5962 (N_5962,N_5480,N_5539);
nand U5963 (N_5963,N_5486,N_5546);
xnor U5964 (N_5964,N_5597,N_5539);
xor U5965 (N_5965,N_5402,N_5694);
or U5966 (N_5966,N_5464,N_5565);
and U5967 (N_5967,N_5605,N_5530);
xor U5968 (N_5968,N_5509,N_5517);
and U5969 (N_5969,N_5665,N_5667);
or U5970 (N_5970,N_5411,N_5446);
and U5971 (N_5971,N_5405,N_5605);
nand U5972 (N_5972,N_5432,N_5659);
and U5973 (N_5973,N_5577,N_5403);
nand U5974 (N_5974,N_5495,N_5481);
and U5975 (N_5975,N_5602,N_5600);
nor U5976 (N_5976,N_5687,N_5533);
or U5977 (N_5977,N_5636,N_5590);
nand U5978 (N_5978,N_5455,N_5545);
xor U5979 (N_5979,N_5449,N_5597);
nand U5980 (N_5980,N_5419,N_5628);
and U5981 (N_5981,N_5666,N_5424);
nand U5982 (N_5982,N_5482,N_5453);
or U5983 (N_5983,N_5688,N_5657);
or U5984 (N_5984,N_5405,N_5464);
xnor U5985 (N_5985,N_5695,N_5596);
nand U5986 (N_5986,N_5691,N_5649);
nand U5987 (N_5987,N_5686,N_5494);
or U5988 (N_5988,N_5559,N_5400);
nor U5989 (N_5989,N_5521,N_5409);
nand U5990 (N_5990,N_5630,N_5610);
nor U5991 (N_5991,N_5680,N_5403);
and U5992 (N_5992,N_5624,N_5668);
nor U5993 (N_5993,N_5495,N_5666);
xor U5994 (N_5994,N_5565,N_5553);
or U5995 (N_5995,N_5443,N_5569);
xor U5996 (N_5996,N_5679,N_5634);
nand U5997 (N_5997,N_5536,N_5527);
or U5998 (N_5998,N_5425,N_5431);
nor U5999 (N_5999,N_5548,N_5693);
nand U6000 (N_6000,N_5911,N_5772);
xor U6001 (N_6001,N_5724,N_5875);
nor U6002 (N_6002,N_5981,N_5942);
nor U6003 (N_6003,N_5700,N_5759);
or U6004 (N_6004,N_5872,N_5945);
nand U6005 (N_6005,N_5899,N_5971);
nand U6006 (N_6006,N_5932,N_5857);
nand U6007 (N_6007,N_5865,N_5780);
nor U6008 (N_6008,N_5866,N_5923);
nor U6009 (N_6009,N_5763,N_5821);
or U6010 (N_6010,N_5963,N_5917);
nand U6011 (N_6011,N_5705,N_5771);
xor U6012 (N_6012,N_5717,N_5831);
xor U6013 (N_6013,N_5855,N_5744);
nand U6014 (N_6014,N_5755,N_5944);
or U6015 (N_6015,N_5712,N_5834);
or U6016 (N_6016,N_5863,N_5869);
or U6017 (N_6017,N_5846,N_5853);
nor U6018 (N_6018,N_5843,N_5743);
nor U6019 (N_6019,N_5709,N_5829);
xor U6020 (N_6020,N_5747,N_5910);
or U6021 (N_6021,N_5902,N_5801);
nand U6022 (N_6022,N_5994,N_5882);
nand U6023 (N_6023,N_5803,N_5817);
nand U6024 (N_6024,N_5805,N_5970);
xor U6025 (N_6025,N_5977,N_5820);
or U6026 (N_6026,N_5986,N_5824);
xor U6027 (N_6027,N_5713,N_5833);
xnor U6028 (N_6028,N_5929,N_5782);
and U6029 (N_6029,N_5984,N_5720);
xor U6030 (N_6030,N_5761,N_5949);
and U6031 (N_6031,N_5969,N_5734);
or U6032 (N_6032,N_5785,N_5768);
nor U6033 (N_6033,N_5979,N_5876);
or U6034 (N_6034,N_5888,N_5922);
xnor U6035 (N_6035,N_5919,N_5773);
and U6036 (N_6036,N_5976,N_5731);
nor U6037 (N_6037,N_5806,N_5940);
and U6038 (N_6038,N_5725,N_5867);
or U6039 (N_6039,N_5729,N_5856);
xor U6040 (N_6040,N_5766,N_5930);
nor U6041 (N_6041,N_5873,N_5823);
or U6042 (N_6042,N_5726,N_5762);
or U6043 (N_6043,N_5914,N_5704);
and U6044 (N_6044,N_5958,N_5799);
xor U6045 (N_6045,N_5751,N_5972);
nand U6046 (N_6046,N_5752,N_5885);
xnor U6047 (N_6047,N_5775,N_5928);
nand U6048 (N_6048,N_5870,N_5999);
nand U6049 (N_6049,N_5800,N_5794);
nand U6050 (N_6050,N_5896,N_5826);
and U6051 (N_6051,N_5769,N_5907);
or U6052 (N_6052,N_5728,N_5813);
xnor U6053 (N_6053,N_5891,N_5965);
or U6054 (N_6054,N_5881,N_5842);
and U6055 (N_6055,N_5955,N_5931);
xnor U6056 (N_6056,N_5733,N_5739);
nand U6057 (N_6057,N_5741,N_5701);
and U6058 (N_6058,N_5992,N_5991);
nor U6059 (N_6059,N_5933,N_5921);
nand U6060 (N_6060,N_5850,N_5948);
xnor U6061 (N_6061,N_5974,N_5900);
or U6062 (N_6062,N_5721,N_5854);
nor U6063 (N_6063,N_5711,N_5987);
and U6064 (N_6064,N_5874,N_5934);
xnor U6065 (N_6065,N_5795,N_5749);
xnor U6066 (N_6066,N_5904,N_5997);
nand U6067 (N_6067,N_5860,N_5892);
nand U6068 (N_6068,N_5920,N_5748);
or U6069 (N_6069,N_5995,N_5774);
or U6070 (N_6070,N_5790,N_5953);
nor U6071 (N_6071,N_5753,N_5836);
nor U6072 (N_6072,N_5973,N_5784);
or U6073 (N_6073,N_5844,N_5758);
nor U6074 (N_6074,N_5760,N_5727);
and U6075 (N_6075,N_5830,N_5791);
nand U6076 (N_6076,N_5887,N_5990);
and U6077 (N_6077,N_5832,N_5783);
and U6078 (N_6078,N_5947,N_5980);
xnor U6079 (N_6079,N_5707,N_5737);
nand U6080 (N_6080,N_5941,N_5779);
nand U6081 (N_6081,N_5835,N_5819);
nor U6082 (N_6082,N_5989,N_5809);
nor U6083 (N_6083,N_5903,N_5786);
xnor U6084 (N_6084,N_5998,N_5877);
and U6085 (N_6085,N_5852,N_5909);
or U6086 (N_6086,N_5978,N_5880);
and U6087 (N_6087,N_5802,N_5943);
nor U6088 (N_6088,N_5871,N_5996);
and U6089 (N_6089,N_5982,N_5745);
xor U6090 (N_6090,N_5935,N_5730);
nand U6091 (N_6091,N_5905,N_5796);
nand U6092 (N_6092,N_5837,N_5862);
nor U6093 (N_6093,N_5898,N_5804);
or U6094 (N_6094,N_5719,N_5957);
nor U6095 (N_6095,N_5845,N_5723);
and U6096 (N_6096,N_5915,N_5946);
or U6097 (N_6097,N_5716,N_5841);
xor U6098 (N_6098,N_5849,N_5702);
or U6099 (N_6099,N_5735,N_5893);
or U6100 (N_6100,N_5889,N_5937);
and U6101 (N_6101,N_5967,N_5956);
nand U6102 (N_6102,N_5825,N_5722);
nand U6103 (N_6103,N_5788,N_5754);
nand U6104 (N_6104,N_5828,N_5859);
or U6105 (N_6105,N_5960,N_5706);
and U6106 (N_6106,N_5840,N_5818);
and U6107 (N_6107,N_5968,N_5810);
nor U6108 (N_6108,N_5797,N_5884);
nand U6109 (N_6109,N_5738,N_5811);
nand U6110 (N_6110,N_5848,N_5959);
nand U6111 (N_6111,N_5916,N_5770);
nand U6112 (N_6112,N_5985,N_5778);
xnor U6113 (N_6113,N_5886,N_5894);
nand U6114 (N_6114,N_5808,N_5792);
nor U6115 (N_6115,N_5757,N_5954);
nor U6116 (N_6116,N_5975,N_5764);
nor U6117 (N_6117,N_5993,N_5746);
xnor U6118 (N_6118,N_5951,N_5858);
nand U6119 (N_6119,N_5868,N_5847);
nand U6120 (N_6120,N_5777,N_5740);
and U6121 (N_6121,N_5913,N_5864);
xnor U6122 (N_6122,N_5906,N_5897);
or U6123 (N_6123,N_5708,N_5879);
or U6124 (N_6124,N_5750,N_5988);
xnor U6125 (N_6125,N_5961,N_5827);
or U6126 (N_6126,N_5952,N_5736);
nor U6127 (N_6127,N_5793,N_5962);
nand U6128 (N_6128,N_5816,N_5776);
nor U6129 (N_6129,N_5765,N_5927);
or U6130 (N_6130,N_5798,N_5966);
and U6131 (N_6131,N_5925,N_5807);
and U6132 (N_6132,N_5924,N_5822);
xnor U6133 (N_6133,N_5781,N_5964);
xnor U6134 (N_6134,N_5861,N_5878);
and U6135 (N_6135,N_5732,N_5912);
nor U6136 (N_6136,N_5787,N_5838);
nand U6137 (N_6137,N_5815,N_5883);
nor U6138 (N_6138,N_5718,N_5742);
xor U6139 (N_6139,N_5939,N_5715);
nand U6140 (N_6140,N_5895,N_5901);
nor U6141 (N_6141,N_5890,N_5936);
nand U6142 (N_6142,N_5926,N_5908);
nor U6143 (N_6143,N_5938,N_5789);
nor U6144 (N_6144,N_5756,N_5814);
and U6145 (N_6145,N_5767,N_5950);
or U6146 (N_6146,N_5983,N_5714);
and U6147 (N_6147,N_5812,N_5851);
nand U6148 (N_6148,N_5703,N_5918);
or U6149 (N_6149,N_5839,N_5710);
and U6150 (N_6150,N_5805,N_5896);
xor U6151 (N_6151,N_5879,N_5985);
nor U6152 (N_6152,N_5762,N_5970);
or U6153 (N_6153,N_5910,N_5843);
nor U6154 (N_6154,N_5837,N_5976);
and U6155 (N_6155,N_5995,N_5776);
nand U6156 (N_6156,N_5963,N_5928);
nor U6157 (N_6157,N_5716,N_5905);
or U6158 (N_6158,N_5802,N_5915);
nor U6159 (N_6159,N_5797,N_5984);
and U6160 (N_6160,N_5812,N_5849);
nor U6161 (N_6161,N_5820,N_5756);
xor U6162 (N_6162,N_5761,N_5860);
and U6163 (N_6163,N_5843,N_5800);
or U6164 (N_6164,N_5990,N_5828);
and U6165 (N_6165,N_5780,N_5986);
xor U6166 (N_6166,N_5801,N_5817);
and U6167 (N_6167,N_5770,N_5990);
xnor U6168 (N_6168,N_5746,N_5916);
and U6169 (N_6169,N_5947,N_5772);
xor U6170 (N_6170,N_5750,N_5798);
xnor U6171 (N_6171,N_5721,N_5919);
or U6172 (N_6172,N_5931,N_5728);
nor U6173 (N_6173,N_5962,N_5904);
or U6174 (N_6174,N_5831,N_5924);
nand U6175 (N_6175,N_5955,N_5913);
nor U6176 (N_6176,N_5870,N_5911);
nor U6177 (N_6177,N_5823,N_5933);
and U6178 (N_6178,N_5833,N_5901);
or U6179 (N_6179,N_5866,N_5751);
and U6180 (N_6180,N_5923,N_5712);
or U6181 (N_6181,N_5921,N_5761);
xnor U6182 (N_6182,N_5924,N_5800);
nand U6183 (N_6183,N_5747,N_5871);
and U6184 (N_6184,N_5928,N_5901);
and U6185 (N_6185,N_5974,N_5959);
nand U6186 (N_6186,N_5970,N_5946);
or U6187 (N_6187,N_5965,N_5751);
nand U6188 (N_6188,N_5737,N_5740);
nand U6189 (N_6189,N_5975,N_5854);
nor U6190 (N_6190,N_5710,N_5796);
nand U6191 (N_6191,N_5895,N_5811);
and U6192 (N_6192,N_5959,N_5866);
nand U6193 (N_6193,N_5807,N_5700);
nand U6194 (N_6194,N_5923,N_5931);
or U6195 (N_6195,N_5901,N_5732);
nand U6196 (N_6196,N_5835,N_5821);
and U6197 (N_6197,N_5746,N_5972);
or U6198 (N_6198,N_5972,N_5784);
and U6199 (N_6199,N_5974,N_5871);
nand U6200 (N_6200,N_5898,N_5796);
and U6201 (N_6201,N_5887,N_5733);
and U6202 (N_6202,N_5804,N_5800);
nand U6203 (N_6203,N_5738,N_5921);
or U6204 (N_6204,N_5833,N_5928);
nand U6205 (N_6205,N_5803,N_5830);
nand U6206 (N_6206,N_5827,N_5732);
xor U6207 (N_6207,N_5906,N_5996);
nor U6208 (N_6208,N_5799,N_5806);
or U6209 (N_6209,N_5758,N_5784);
nand U6210 (N_6210,N_5815,N_5801);
nand U6211 (N_6211,N_5834,N_5844);
nand U6212 (N_6212,N_5884,N_5879);
or U6213 (N_6213,N_5802,N_5838);
xnor U6214 (N_6214,N_5739,N_5977);
nand U6215 (N_6215,N_5935,N_5851);
or U6216 (N_6216,N_5948,N_5869);
xnor U6217 (N_6217,N_5733,N_5853);
nor U6218 (N_6218,N_5925,N_5950);
xor U6219 (N_6219,N_5841,N_5718);
nor U6220 (N_6220,N_5779,N_5969);
or U6221 (N_6221,N_5942,N_5833);
xnor U6222 (N_6222,N_5815,N_5982);
or U6223 (N_6223,N_5955,N_5989);
nor U6224 (N_6224,N_5792,N_5845);
nor U6225 (N_6225,N_5867,N_5830);
xor U6226 (N_6226,N_5866,N_5771);
nor U6227 (N_6227,N_5708,N_5976);
xor U6228 (N_6228,N_5706,N_5838);
or U6229 (N_6229,N_5709,N_5706);
nor U6230 (N_6230,N_5867,N_5834);
or U6231 (N_6231,N_5839,N_5910);
xor U6232 (N_6232,N_5739,N_5987);
and U6233 (N_6233,N_5870,N_5725);
nand U6234 (N_6234,N_5773,N_5779);
nor U6235 (N_6235,N_5710,N_5886);
and U6236 (N_6236,N_5772,N_5794);
nand U6237 (N_6237,N_5797,N_5702);
nor U6238 (N_6238,N_5805,N_5907);
and U6239 (N_6239,N_5838,N_5991);
nor U6240 (N_6240,N_5950,N_5722);
nor U6241 (N_6241,N_5811,N_5701);
xnor U6242 (N_6242,N_5943,N_5911);
and U6243 (N_6243,N_5914,N_5845);
nand U6244 (N_6244,N_5975,N_5870);
nand U6245 (N_6245,N_5853,N_5938);
or U6246 (N_6246,N_5959,N_5785);
nor U6247 (N_6247,N_5723,N_5737);
and U6248 (N_6248,N_5805,N_5842);
or U6249 (N_6249,N_5721,N_5740);
and U6250 (N_6250,N_5850,N_5814);
or U6251 (N_6251,N_5833,N_5745);
and U6252 (N_6252,N_5883,N_5726);
and U6253 (N_6253,N_5947,N_5862);
xnor U6254 (N_6254,N_5728,N_5804);
nand U6255 (N_6255,N_5942,N_5965);
or U6256 (N_6256,N_5737,N_5908);
or U6257 (N_6257,N_5892,N_5838);
nand U6258 (N_6258,N_5999,N_5963);
nand U6259 (N_6259,N_5957,N_5911);
nand U6260 (N_6260,N_5796,N_5797);
and U6261 (N_6261,N_5790,N_5947);
and U6262 (N_6262,N_5710,N_5783);
nor U6263 (N_6263,N_5905,N_5882);
or U6264 (N_6264,N_5794,N_5783);
nand U6265 (N_6265,N_5968,N_5786);
nand U6266 (N_6266,N_5780,N_5713);
nor U6267 (N_6267,N_5703,N_5769);
or U6268 (N_6268,N_5771,N_5752);
nand U6269 (N_6269,N_5975,N_5946);
xnor U6270 (N_6270,N_5757,N_5818);
nor U6271 (N_6271,N_5891,N_5849);
nand U6272 (N_6272,N_5871,N_5731);
nor U6273 (N_6273,N_5825,N_5729);
or U6274 (N_6274,N_5893,N_5754);
nor U6275 (N_6275,N_5973,N_5966);
and U6276 (N_6276,N_5814,N_5766);
xnor U6277 (N_6277,N_5956,N_5789);
nor U6278 (N_6278,N_5813,N_5833);
or U6279 (N_6279,N_5900,N_5842);
nand U6280 (N_6280,N_5833,N_5951);
and U6281 (N_6281,N_5723,N_5726);
or U6282 (N_6282,N_5939,N_5885);
xnor U6283 (N_6283,N_5972,N_5884);
and U6284 (N_6284,N_5930,N_5785);
nand U6285 (N_6285,N_5780,N_5752);
nand U6286 (N_6286,N_5818,N_5962);
or U6287 (N_6287,N_5762,N_5944);
nor U6288 (N_6288,N_5830,N_5868);
xnor U6289 (N_6289,N_5718,N_5821);
nand U6290 (N_6290,N_5778,N_5869);
xor U6291 (N_6291,N_5783,N_5891);
or U6292 (N_6292,N_5817,N_5846);
and U6293 (N_6293,N_5747,N_5810);
or U6294 (N_6294,N_5918,N_5818);
nor U6295 (N_6295,N_5903,N_5840);
and U6296 (N_6296,N_5988,N_5780);
nor U6297 (N_6297,N_5830,N_5940);
xnor U6298 (N_6298,N_5742,N_5797);
nor U6299 (N_6299,N_5899,N_5734);
nor U6300 (N_6300,N_6225,N_6222);
nor U6301 (N_6301,N_6193,N_6140);
or U6302 (N_6302,N_6262,N_6022);
nor U6303 (N_6303,N_6097,N_6171);
nor U6304 (N_6304,N_6054,N_6187);
nor U6305 (N_6305,N_6076,N_6045);
nand U6306 (N_6306,N_6294,N_6084);
nand U6307 (N_6307,N_6079,N_6100);
nor U6308 (N_6308,N_6166,N_6053);
or U6309 (N_6309,N_6024,N_6023);
xor U6310 (N_6310,N_6252,N_6108);
and U6311 (N_6311,N_6082,N_6243);
xor U6312 (N_6312,N_6133,N_6078);
or U6313 (N_6313,N_6035,N_6272);
or U6314 (N_6314,N_6107,N_6158);
and U6315 (N_6315,N_6293,N_6092);
xor U6316 (N_6316,N_6221,N_6261);
nor U6317 (N_6317,N_6014,N_6271);
nor U6318 (N_6318,N_6147,N_6275);
nand U6319 (N_6319,N_6167,N_6062);
nor U6320 (N_6320,N_6118,N_6051);
nand U6321 (N_6321,N_6138,N_6152);
nand U6322 (N_6322,N_6017,N_6223);
nand U6323 (N_6323,N_6257,N_6141);
xnor U6324 (N_6324,N_6292,N_6284);
and U6325 (N_6325,N_6037,N_6117);
and U6326 (N_6326,N_6049,N_6248);
xnor U6327 (N_6327,N_6273,N_6006);
nor U6328 (N_6328,N_6214,N_6011);
and U6329 (N_6329,N_6212,N_6266);
or U6330 (N_6330,N_6040,N_6186);
xor U6331 (N_6331,N_6299,N_6095);
or U6332 (N_6332,N_6025,N_6163);
xnor U6333 (N_6333,N_6020,N_6149);
or U6334 (N_6334,N_6148,N_6238);
xnor U6335 (N_6335,N_6285,N_6122);
and U6336 (N_6336,N_6150,N_6042);
xnor U6337 (N_6337,N_6044,N_6290);
nor U6338 (N_6338,N_6139,N_6204);
and U6339 (N_6339,N_6205,N_6200);
nand U6340 (N_6340,N_6111,N_6229);
and U6341 (N_6341,N_6227,N_6287);
nand U6342 (N_6342,N_6072,N_6192);
or U6343 (N_6343,N_6196,N_6159);
nor U6344 (N_6344,N_6016,N_6146);
and U6345 (N_6345,N_6086,N_6128);
nand U6346 (N_6346,N_6096,N_6197);
nor U6347 (N_6347,N_6098,N_6008);
xnor U6348 (N_6348,N_6109,N_6286);
xnor U6349 (N_6349,N_6208,N_6242);
and U6350 (N_6350,N_6274,N_6069);
nand U6351 (N_6351,N_6081,N_6104);
or U6352 (N_6352,N_6028,N_6291);
xor U6353 (N_6353,N_6009,N_6189);
nand U6354 (N_6354,N_6179,N_6094);
nor U6355 (N_6355,N_6241,N_6143);
and U6356 (N_6356,N_6256,N_6112);
nor U6357 (N_6357,N_6087,N_6001);
nor U6358 (N_6358,N_6090,N_6002);
or U6359 (N_6359,N_6185,N_6019);
or U6360 (N_6360,N_6151,N_6036);
and U6361 (N_6361,N_6047,N_6064);
or U6362 (N_6362,N_6032,N_6101);
xor U6363 (N_6363,N_6161,N_6178);
nand U6364 (N_6364,N_6153,N_6198);
and U6365 (N_6365,N_6177,N_6254);
or U6366 (N_6366,N_6067,N_6282);
and U6367 (N_6367,N_6074,N_6235);
and U6368 (N_6368,N_6211,N_6279);
and U6369 (N_6369,N_6247,N_6057);
or U6370 (N_6370,N_6270,N_6216);
nand U6371 (N_6371,N_6259,N_6199);
xor U6372 (N_6372,N_6168,N_6219);
nor U6373 (N_6373,N_6277,N_6137);
nand U6374 (N_6374,N_6236,N_6120);
nor U6375 (N_6375,N_6245,N_6134);
and U6376 (N_6376,N_6075,N_6065);
and U6377 (N_6377,N_6070,N_6220);
nor U6378 (N_6378,N_6055,N_6126);
nor U6379 (N_6379,N_6105,N_6142);
or U6380 (N_6380,N_6106,N_6056);
xnor U6381 (N_6381,N_6007,N_6066);
nor U6382 (N_6382,N_6155,N_6080);
and U6383 (N_6383,N_6224,N_6071);
xnor U6384 (N_6384,N_6253,N_6162);
and U6385 (N_6385,N_6131,N_6210);
and U6386 (N_6386,N_6052,N_6102);
nor U6387 (N_6387,N_6269,N_6046);
nand U6388 (N_6388,N_6154,N_6237);
and U6389 (N_6389,N_6175,N_6289);
nand U6390 (N_6390,N_6264,N_6113);
nand U6391 (N_6391,N_6012,N_6093);
nor U6392 (N_6392,N_6173,N_6207);
and U6393 (N_6393,N_6296,N_6181);
nor U6394 (N_6394,N_6201,N_6073);
xor U6395 (N_6395,N_6283,N_6295);
or U6396 (N_6396,N_6184,N_6050);
nor U6397 (N_6397,N_6145,N_6209);
or U6398 (N_6398,N_6156,N_6191);
nand U6399 (N_6399,N_6115,N_6135);
xor U6400 (N_6400,N_6132,N_6030);
or U6401 (N_6401,N_6061,N_6215);
xor U6402 (N_6402,N_6039,N_6041);
nand U6403 (N_6403,N_6232,N_6027);
and U6404 (N_6404,N_6015,N_6103);
and U6405 (N_6405,N_6240,N_6083);
xnor U6406 (N_6406,N_6249,N_6116);
or U6407 (N_6407,N_6060,N_6085);
xor U6408 (N_6408,N_6000,N_6182);
and U6409 (N_6409,N_6226,N_6206);
or U6410 (N_6410,N_6258,N_6038);
and U6411 (N_6411,N_6281,N_6130);
nor U6412 (N_6412,N_6034,N_6213);
xor U6413 (N_6413,N_6231,N_6121);
xor U6414 (N_6414,N_6031,N_6136);
or U6415 (N_6415,N_6088,N_6278);
or U6416 (N_6416,N_6129,N_6244);
nor U6417 (N_6417,N_6110,N_6033);
or U6418 (N_6418,N_6043,N_6260);
and U6419 (N_6419,N_6013,N_6063);
nor U6420 (N_6420,N_6288,N_6077);
nand U6421 (N_6421,N_6169,N_6125);
and U6422 (N_6422,N_6114,N_6202);
nand U6423 (N_6423,N_6228,N_6172);
nor U6424 (N_6424,N_6089,N_6251);
xnor U6425 (N_6425,N_6194,N_6003);
nand U6426 (N_6426,N_6010,N_6268);
or U6427 (N_6427,N_6180,N_6267);
and U6428 (N_6428,N_6176,N_6218);
and U6429 (N_6429,N_6119,N_6029);
or U6430 (N_6430,N_6018,N_6263);
or U6431 (N_6431,N_6127,N_6058);
or U6432 (N_6432,N_6048,N_6298);
or U6433 (N_6433,N_6276,N_6190);
or U6434 (N_6434,N_6174,N_6068);
or U6435 (N_6435,N_6230,N_6144);
and U6436 (N_6436,N_6157,N_6239);
nand U6437 (N_6437,N_6160,N_6026);
xnor U6438 (N_6438,N_6005,N_6170);
nor U6439 (N_6439,N_6195,N_6091);
nand U6440 (N_6440,N_6059,N_6297);
nand U6441 (N_6441,N_6099,N_6004);
or U6442 (N_6442,N_6164,N_6188);
or U6443 (N_6443,N_6124,N_6265);
or U6444 (N_6444,N_6203,N_6217);
nand U6445 (N_6445,N_6255,N_6021);
nor U6446 (N_6446,N_6246,N_6280);
and U6447 (N_6447,N_6183,N_6165);
nand U6448 (N_6448,N_6123,N_6233);
and U6449 (N_6449,N_6234,N_6250);
xor U6450 (N_6450,N_6235,N_6150);
xnor U6451 (N_6451,N_6184,N_6084);
nor U6452 (N_6452,N_6255,N_6068);
and U6453 (N_6453,N_6139,N_6266);
xnor U6454 (N_6454,N_6194,N_6128);
nor U6455 (N_6455,N_6197,N_6248);
xor U6456 (N_6456,N_6228,N_6251);
nor U6457 (N_6457,N_6008,N_6193);
nor U6458 (N_6458,N_6194,N_6094);
and U6459 (N_6459,N_6191,N_6102);
xor U6460 (N_6460,N_6190,N_6288);
nand U6461 (N_6461,N_6166,N_6226);
and U6462 (N_6462,N_6107,N_6245);
xnor U6463 (N_6463,N_6203,N_6033);
nor U6464 (N_6464,N_6270,N_6296);
or U6465 (N_6465,N_6299,N_6003);
nor U6466 (N_6466,N_6089,N_6086);
nand U6467 (N_6467,N_6235,N_6002);
or U6468 (N_6468,N_6034,N_6090);
nand U6469 (N_6469,N_6133,N_6229);
xor U6470 (N_6470,N_6006,N_6054);
or U6471 (N_6471,N_6209,N_6076);
or U6472 (N_6472,N_6101,N_6279);
nand U6473 (N_6473,N_6056,N_6123);
nand U6474 (N_6474,N_6018,N_6105);
or U6475 (N_6475,N_6186,N_6083);
xor U6476 (N_6476,N_6163,N_6097);
or U6477 (N_6477,N_6268,N_6124);
or U6478 (N_6478,N_6149,N_6015);
and U6479 (N_6479,N_6266,N_6206);
or U6480 (N_6480,N_6274,N_6143);
xor U6481 (N_6481,N_6167,N_6118);
nor U6482 (N_6482,N_6215,N_6175);
nor U6483 (N_6483,N_6060,N_6141);
and U6484 (N_6484,N_6264,N_6149);
and U6485 (N_6485,N_6071,N_6227);
xnor U6486 (N_6486,N_6119,N_6193);
nor U6487 (N_6487,N_6074,N_6169);
nand U6488 (N_6488,N_6021,N_6138);
nand U6489 (N_6489,N_6136,N_6173);
xnor U6490 (N_6490,N_6039,N_6273);
and U6491 (N_6491,N_6272,N_6242);
nand U6492 (N_6492,N_6213,N_6236);
xor U6493 (N_6493,N_6156,N_6256);
nand U6494 (N_6494,N_6274,N_6170);
and U6495 (N_6495,N_6049,N_6192);
and U6496 (N_6496,N_6249,N_6142);
and U6497 (N_6497,N_6154,N_6159);
or U6498 (N_6498,N_6042,N_6139);
xor U6499 (N_6499,N_6013,N_6236);
nand U6500 (N_6500,N_6106,N_6086);
nor U6501 (N_6501,N_6056,N_6177);
xor U6502 (N_6502,N_6151,N_6215);
xor U6503 (N_6503,N_6231,N_6286);
or U6504 (N_6504,N_6013,N_6196);
and U6505 (N_6505,N_6053,N_6297);
or U6506 (N_6506,N_6297,N_6185);
nand U6507 (N_6507,N_6180,N_6041);
xnor U6508 (N_6508,N_6226,N_6205);
nand U6509 (N_6509,N_6267,N_6140);
nand U6510 (N_6510,N_6288,N_6022);
or U6511 (N_6511,N_6116,N_6007);
and U6512 (N_6512,N_6079,N_6063);
or U6513 (N_6513,N_6169,N_6197);
nor U6514 (N_6514,N_6235,N_6112);
nand U6515 (N_6515,N_6159,N_6287);
or U6516 (N_6516,N_6036,N_6053);
and U6517 (N_6517,N_6165,N_6138);
or U6518 (N_6518,N_6240,N_6001);
xor U6519 (N_6519,N_6254,N_6007);
nor U6520 (N_6520,N_6120,N_6183);
nand U6521 (N_6521,N_6028,N_6007);
xor U6522 (N_6522,N_6113,N_6010);
xor U6523 (N_6523,N_6073,N_6243);
or U6524 (N_6524,N_6115,N_6164);
xnor U6525 (N_6525,N_6016,N_6057);
xnor U6526 (N_6526,N_6074,N_6119);
nand U6527 (N_6527,N_6202,N_6244);
or U6528 (N_6528,N_6129,N_6272);
nand U6529 (N_6529,N_6298,N_6173);
nand U6530 (N_6530,N_6041,N_6107);
nand U6531 (N_6531,N_6207,N_6042);
nor U6532 (N_6532,N_6107,N_6146);
xor U6533 (N_6533,N_6067,N_6154);
or U6534 (N_6534,N_6126,N_6118);
nor U6535 (N_6535,N_6257,N_6177);
and U6536 (N_6536,N_6188,N_6072);
nor U6537 (N_6537,N_6005,N_6299);
or U6538 (N_6538,N_6261,N_6128);
xnor U6539 (N_6539,N_6104,N_6218);
xnor U6540 (N_6540,N_6058,N_6014);
or U6541 (N_6541,N_6014,N_6250);
nor U6542 (N_6542,N_6095,N_6120);
nor U6543 (N_6543,N_6176,N_6026);
nand U6544 (N_6544,N_6240,N_6040);
or U6545 (N_6545,N_6163,N_6078);
and U6546 (N_6546,N_6031,N_6177);
or U6547 (N_6547,N_6011,N_6124);
nand U6548 (N_6548,N_6156,N_6081);
or U6549 (N_6549,N_6008,N_6096);
and U6550 (N_6550,N_6291,N_6161);
nand U6551 (N_6551,N_6299,N_6267);
or U6552 (N_6552,N_6041,N_6209);
or U6553 (N_6553,N_6059,N_6027);
nor U6554 (N_6554,N_6075,N_6228);
nor U6555 (N_6555,N_6270,N_6111);
and U6556 (N_6556,N_6108,N_6232);
or U6557 (N_6557,N_6132,N_6103);
xor U6558 (N_6558,N_6282,N_6245);
nand U6559 (N_6559,N_6265,N_6209);
or U6560 (N_6560,N_6177,N_6271);
and U6561 (N_6561,N_6263,N_6146);
and U6562 (N_6562,N_6262,N_6066);
and U6563 (N_6563,N_6037,N_6130);
or U6564 (N_6564,N_6196,N_6107);
or U6565 (N_6565,N_6242,N_6046);
or U6566 (N_6566,N_6255,N_6099);
nor U6567 (N_6567,N_6016,N_6291);
xor U6568 (N_6568,N_6097,N_6009);
or U6569 (N_6569,N_6205,N_6289);
or U6570 (N_6570,N_6084,N_6079);
nand U6571 (N_6571,N_6048,N_6172);
nor U6572 (N_6572,N_6079,N_6026);
xnor U6573 (N_6573,N_6192,N_6055);
or U6574 (N_6574,N_6209,N_6256);
or U6575 (N_6575,N_6032,N_6036);
or U6576 (N_6576,N_6013,N_6018);
and U6577 (N_6577,N_6134,N_6085);
nand U6578 (N_6578,N_6240,N_6093);
or U6579 (N_6579,N_6258,N_6168);
nand U6580 (N_6580,N_6286,N_6167);
nor U6581 (N_6581,N_6099,N_6224);
xor U6582 (N_6582,N_6247,N_6206);
nor U6583 (N_6583,N_6145,N_6052);
or U6584 (N_6584,N_6077,N_6210);
nor U6585 (N_6585,N_6167,N_6086);
nor U6586 (N_6586,N_6146,N_6203);
nor U6587 (N_6587,N_6039,N_6066);
or U6588 (N_6588,N_6105,N_6219);
xnor U6589 (N_6589,N_6161,N_6298);
nor U6590 (N_6590,N_6066,N_6241);
or U6591 (N_6591,N_6072,N_6229);
nor U6592 (N_6592,N_6299,N_6189);
or U6593 (N_6593,N_6253,N_6057);
or U6594 (N_6594,N_6154,N_6102);
or U6595 (N_6595,N_6102,N_6201);
xnor U6596 (N_6596,N_6121,N_6236);
or U6597 (N_6597,N_6232,N_6238);
or U6598 (N_6598,N_6163,N_6204);
and U6599 (N_6599,N_6044,N_6275);
xor U6600 (N_6600,N_6482,N_6580);
nand U6601 (N_6601,N_6418,N_6399);
nand U6602 (N_6602,N_6476,N_6367);
xnor U6603 (N_6603,N_6357,N_6471);
nand U6604 (N_6604,N_6431,N_6341);
nand U6605 (N_6605,N_6489,N_6304);
xor U6606 (N_6606,N_6344,N_6523);
and U6607 (N_6607,N_6402,N_6306);
nor U6608 (N_6608,N_6408,N_6562);
and U6609 (N_6609,N_6353,N_6345);
nand U6610 (N_6610,N_6438,N_6546);
nor U6611 (N_6611,N_6404,N_6444);
nor U6612 (N_6612,N_6316,N_6406);
and U6613 (N_6613,N_6330,N_6417);
or U6614 (N_6614,N_6588,N_6392);
nor U6615 (N_6615,N_6581,N_6387);
nand U6616 (N_6616,N_6323,N_6479);
nor U6617 (N_6617,N_6597,N_6544);
nor U6618 (N_6618,N_6383,N_6415);
and U6619 (N_6619,N_6394,N_6473);
xnor U6620 (N_6620,N_6366,N_6337);
or U6621 (N_6621,N_6401,N_6569);
nand U6622 (N_6622,N_6380,N_6339);
xor U6623 (N_6623,N_6371,N_6400);
or U6624 (N_6624,N_6559,N_6318);
or U6625 (N_6625,N_6589,N_6596);
xnor U6626 (N_6626,N_6551,N_6434);
or U6627 (N_6627,N_6556,N_6303);
xnor U6628 (N_6628,N_6501,N_6567);
or U6629 (N_6629,N_6511,N_6552);
or U6630 (N_6630,N_6319,N_6557);
nand U6631 (N_6631,N_6382,N_6469);
xor U6632 (N_6632,N_6419,N_6514);
xnor U6633 (N_6633,N_6350,N_6351);
nand U6634 (N_6634,N_6409,N_6592);
nand U6635 (N_6635,N_6381,N_6553);
or U6636 (N_6636,N_6472,N_6426);
nand U6637 (N_6637,N_6529,N_6453);
nor U6638 (N_6638,N_6590,N_6495);
nor U6639 (N_6639,N_6414,N_6445);
and U6640 (N_6640,N_6389,N_6550);
and U6641 (N_6641,N_6300,N_6522);
xor U6642 (N_6642,N_6458,N_6313);
xor U6643 (N_6643,N_6599,N_6346);
nor U6644 (N_6644,N_6416,N_6494);
xor U6645 (N_6645,N_6533,N_6595);
and U6646 (N_6646,N_6502,N_6428);
nor U6647 (N_6647,N_6365,N_6435);
and U6648 (N_6648,N_6439,N_6390);
xnor U6649 (N_6649,N_6375,N_6521);
nand U6650 (N_6650,N_6467,N_6311);
nor U6651 (N_6651,N_6541,N_6457);
nand U6652 (N_6652,N_6591,N_6448);
or U6653 (N_6653,N_6301,N_6310);
nor U6654 (N_6654,N_6496,N_6477);
nor U6655 (N_6655,N_6369,N_6446);
or U6656 (N_6656,N_6530,N_6432);
or U6657 (N_6657,N_6534,N_6585);
nand U6658 (N_6658,N_6430,N_6348);
or U6659 (N_6659,N_6542,N_6427);
xnor U6660 (N_6660,N_6520,N_6395);
nand U6661 (N_6661,N_6334,N_6566);
xnor U6662 (N_6662,N_6468,N_6425);
nor U6663 (N_6663,N_6437,N_6558);
or U6664 (N_6664,N_6504,N_6579);
and U6665 (N_6665,N_6487,N_6412);
xor U6666 (N_6666,N_6516,N_6362);
nor U6667 (N_6667,N_6583,N_6374);
xor U6668 (N_6668,N_6503,N_6547);
nor U6669 (N_6669,N_6574,N_6452);
and U6670 (N_6670,N_6584,N_6440);
nor U6671 (N_6671,N_6466,N_6568);
and U6672 (N_6672,N_6548,N_6407);
or U6673 (N_6673,N_6524,N_6535);
xnor U6674 (N_6674,N_6454,N_6309);
nor U6675 (N_6675,N_6498,N_6325);
xor U6676 (N_6676,N_6305,N_6436);
nor U6677 (N_6677,N_6460,N_6308);
and U6678 (N_6678,N_6450,N_6540);
and U6679 (N_6679,N_6526,N_6499);
nor U6680 (N_6680,N_6360,N_6485);
xnor U6681 (N_6681,N_6314,N_6361);
nand U6682 (N_6682,N_6384,N_6481);
nand U6683 (N_6683,N_6359,N_6328);
or U6684 (N_6684,N_6349,N_6320);
xor U6685 (N_6685,N_6488,N_6563);
nand U6686 (N_6686,N_6470,N_6449);
or U6687 (N_6687,N_6575,N_6528);
nor U6688 (N_6688,N_6391,N_6386);
nor U6689 (N_6689,N_6447,N_6411);
nor U6690 (N_6690,N_6517,N_6388);
nand U6691 (N_6691,N_6465,N_6587);
nor U6692 (N_6692,N_6582,N_6405);
nor U6693 (N_6693,N_6486,N_6474);
nor U6694 (N_6694,N_6463,N_6519);
xor U6695 (N_6695,N_6338,N_6385);
or U6696 (N_6696,N_6327,N_6397);
or U6697 (N_6697,N_6429,N_6598);
nor U6698 (N_6698,N_6594,N_6364);
and U6699 (N_6699,N_6370,N_6451);
xor U6700 (N_6700,N_6420,N_6377);
or U6701 (N_6701,N_6322,N_6537);
xnor U6702 (N_6702,N_6512,N_6342);
nand U6703 (N_6703,N_6549,N_6480);
or U6704 (N_6704,N_6363,N_6510);
nor U6705 (N_6705,N_6376,N_6393);
nor U6706 (N_6706,N_6356,N_6507);
xor U6707 (N_6707,N_6565,N_6459);
and U6708 (N_6708,N_6505,N_6332);
and U6709 (N_6709,N_6379,N_6561);
or U6710 (N_6710,N_6484,N_6492);
nor U6711 (N_6711,N_6413,N_6576);
or U6712 (N_6712,N_6573,N_6324);
xnor U6713 (N_6713,N_6586,N_6545);
nand U6714 (N_6714,N_6422,N_6478);
or U6715 (N_6715,N_6455,N_6536);
nor U6716 (N_6716,N_6321,N_6560);
nor U6717 (N_6717,N_6442,N_6372);
nand U6718 (N_6718,N_6424,N_6340);
or U6719 (N_6719,N_6302,N_6493);
and U6720 (N_6720,N_6532,N_6531);
nor U6721 (N_6721,N_6354,N_6497);
and U6722 (N_6722,N_6347,N_6315);
nor U6723 (N_6723,N_6491,N_6513);
nand U6724 (N_6724,N_6462,N_6464);
or U6725 (N_6725,N_6490,N_6396);
xor U6726 (N_6726,N_6355,N_6525);
or U6727 (N_6727,N_6403,N_6421);
nor U6728 (N_6728,N_6508,N_6433);
xnor U6729 (N_6729,N_6518,N_6515);
xnor U6730 (N_6730,N_6368,N_6506);
nor U6731 (N_6731,N_6326,N_6443);
xnor U6732 (N_6732,N_6441,N_6333);
nand U6733 (N_6733,N_6527,N_6538);
or U6734 (N_6734,N_6564,N_6329);
and U6735 (N_6735,N_6577,N_6410);
nand U6736 (N_6736,N_6500,N_6317);
nand U6737 (N_6737,N_6343,N_6312);
or U6738 (N_6738,N_6509,N_6593);
nand U6739 (N_6739,N_6539,N_6307);
and U6740 (N_6740,N_6398,N_6456);
nand U6741 (N_6741,N_6578,N_6461);
and U6742 (N_6742,N_6572,N_6570);
or U6743 (N_6743,N_6571,N_6475);
nand U6744 (N_6744,N_6378,N_6373);
xor U6745 (N_6745,N_6554,N_6331);
nor U6746 (N_6746,N_6352,N_6335);
nand U6747 (N_6747,N_6555,N_6543);
and U6748 (N_6748,N_6483,N_6423);
nor U6749 (N_6749,N_6336,N_6358);
nand U6750 (N_6750,N_6393,N_6371);
nand U6751 (N_6751,N_6372,N_6421);
xor U6752 (N_6752,N_6543,N_6551);
or U6753 (N_6753,N_6396,N_6403);
or U6754 (N_6754,N_6480,N_6522);
nor U6755 (N_6755,N_6337,N_6379);
xor U6756 (N_6756,N_6322,N_6433);
xor U6757 (N_6757,N_6391,N_6432);
and U6758 (N_6758,N_6338,N_6322);
xnor U6759 (N_6759,N_6372,N_6319);
xor U6760 (N_6760,N_6568,N_6583);
nor U6761 (N_6761,N_6525,N_6472);
xor U6762 (N_6762,N_6341,N_6522);
nor U6763 (N_6763,N_6449,N_6515);
or U6764 (N_6764,N_6359,N_6319);
nand U6765 (N_6765,N_6531,N_6506);
and U6766 (N_6766,N_6584,N_6375);
nor U6767 (N_6767,N_6406,N_6567);
and U6768 (N_6768,N_6567,N_6450);
nor U6769 (N_6769,N_6566,N_6556);
nand U6770 (N_6770,N_6521,N_6435);
nand U6771 (N_6771,N_6389,N_6521);
xor U6772 (N_6772,N_6506,N_6536);
and U6773 (N_6773,N_6377,N_6340);
nor U6774 (N_6774,N_6448,N_6507);
xnor U6775 (N_6775,N_6386,N_6318);
or U6776 (N_6776,N_6478,N_6449);
nand U6777 (N_6777,N_6555,N_6393);
or U6778 (N_6778,N_6462,N_6544);
xnor U6779 (N_6779,N_6508,N_6404);
or U6780 (N_6780,N_6347,N_6437);
or U6781 (N_6781,N_6582,N_6415);
nand U6782 (N_6782,N_6340,N_6427);
or U6783 (N_6783,N_6471,N_6374);
and U6784 (N_6784,N_6381,N_6597);
nand U6785 (N_6785,N_6597,N_6520);
or U6786 (N_6786,N_6544,N_6323);
nand U6787 (N_6787,N_6546,N_6591);
nand U6788 (N_6788,N_6536,N_6335);
or U6789 (N_6789,N_6461,N_6483);
or U6790 (N_6790,N_6598,N_6370);
xor U6791 (N_6791,N_6462,N_6586);
nor U6792 (N_6792,N_6345,N_6423);
nor U6793 (N_6793,N_6574,N_6591);
or U6794 (N_6794,N_6319,N_6428);
and U6795 (N_6795,N_6410,N_6366);
and U6796 (N_6796,N_6398,N_6365);
nand U6797 (N_6797,N_6340,N_6581);
nand U6798 (N_6798,N_6583,N_6419);
and U6799 (N_6799,N_6312,N_6495);
and U6800 (N_6800,N_6352,N_6497);
nor U6801 (N_6801,N_6305,N_6307);
and U6802 (N_6802,N_6564,N_6342);
xor U6803 (N_6803,N_6495,N_6586);
xnor U6804 (N_6804,N_6580,N_6571);
xor U6805 (N_6805,N_6310,N_6440);
xnor U6806 (N_6806,N_6341,N_6413);
nor U6807 (N_6807,N_6442,N_6571);
xnor U6808 (N_6808,N_6457,N_6563);
nor U6809 (N_6809,N_6435,N_6542);
and U6810 (N_6810,N_6531,N_6353);
and U6811 (N_6811,N_6522,N_6340);
nand U6812 (N_6812,N_6424,N_6393);
or U6813 (N_6813,N_6443,N_6521);
and U6814 (N_6814,N_6363,N_6390);
or U6815 (N_6815,N_6354,N_6460);
or U6816 (N_6816,N_6564,N_6344);
nand U6817 (N_6817,N_6330,N_6325);
and U6818 (N_6818,N_6585,N_6478);
nor U6819 (N_6819,N_6580,N_6325);
or U6820 (N_6820,N_6461,N_6449);
xor U6821 (N_6821,N_6348,N_6504);
nand U6822 (N_6822,N_6479,N_6393);
and U6823 (N_6823,N_6443,N_6579);
or U6824 (N_6824,N_6499,N_6407);
xor U6825 (N_6825,N_6595,N_6448);
or U6826 (N_6826,N_6473,N_6498);
nand U6827 (N_6827,N_6314,N_6436);
xor U6828 (N_6828,N_6413,N_6566);
and U6829 (N_6829,N_6530,N_6409);
nor U6830 (N_6830,N_6362,N_6468);
xor U6831 (N_6831,N_6333,N_6311);
and U6832 (N_6832,N_6345,N_6453);
and U6833 (N_6833,N_6526,N_6392);
or U6834 (N_6834,N_6456,N_6420);
nand U6835 (N_6835,N_6451,N_6506);
nor U6836 (N_6836,N_6365,N_6338);
or U6837 (N_6837,N_6306,N_6406);
nand U6838 (N_6838,N_6574,N_6568);
xnor U6839 (N_6839,N_6485,N_6308);
or U6840 (N_6840,N_6437,N_6404);
nand U6841 (N_6841,N_6533,N_6410);
and U6842 (N_6842,N_6372,N_6405);
and U6843 (N_6843,N_6349,N_6482);
or U6844 (N_6844,N_6340,N_6539);
and U6845 (N_6845,N_6485,N_6413);
and U6846 (N_6846,N_6425,N_6307);
nand U6847 (N_6847,N_6450,N_6430);
and U6848 (N_6848,N_6424,N_6331);
nor U6849 (N_6849,N_6572,N_6357);
xnor U6850 (N_6850,N_6446,N_6375);
nand U6851 (N_6851,N_6521,N_6466);
nand U6852 (N_6852,N_6335,N_6500);
xnor U6853 (N_6853,N_6422,N_6310);
nor U6854 (N_6854,N_6331,N_6448);
and U6855 (N_6855,N_6454,N_6541);
and U6856 (N_6856,N_6420,N_6464);
xor U6857 (N_6857,N_6506,N_6421);
and U6858 (N_6858,N_6306,N_6425);
xor U6859 (N_6859,N_6484,N_6488);
and U6860 (N_6860,N_6581,N_6300);
nor U6861 (N_6861,N_6419,N_6464);
nand U6862 (N_6862,N_6397,N_6484);
or U6863 (N_6863,N_6563,N_6423);
nor U6864 (N_6864,N_6445,N_6409);
and U6865 (N_6865,N_6401,N_6549);
nand U6866 (N_6866,N_6362,N_6543);
nand U6867 (N_6867,N_6383,N_6363);
xor U6868 (N_6868,N_6417,N_6465);
nor U6869 (N_6869,N_6544,N_6388);
nand U6870 (N_6870,N_6585,N_6535);
and U6871 (N_6871,N_6407,N_6446);
nor U6872 (N_6872,N_6365,N_6319);
xor U6873 (N_6873,N_6338,N_6508);
and U6874 (N_6874,N_6379,N_6319);
xor U6875 (N_6875,N_6388,N_6479);
nor U6876 (N_6876,N_6327,N_6407);
or U6877 (N_6877,N_6586,N_6555);
nor U6878 (N_6878,N_6512,N_6508);
nand U6879 (N_6879,N_6316,N_6566);
nor U6880 (N_6880,N_6504,N_6338);
xor U6881 (N_6881,N_6501,N_6517);
xnor U6882 (N_6882,N_6439,N_6578);
nand U6883 (N_6883,N_6378,N_6308);
nand U6884 (N_6884,N_6410,N_6575);
xnor U6885 (N_6885,N_6599,N_6497);
and U6886 (N_6886,N_6313,N_6598);
xor U6887 (N_6887,N_6350,N_6567);
xnor U6888 (N_6888,N_6545,N_6356);
and U6889 (N_6889,N_6321,N_6443);
nand U6890 (N_6890,N_6380,N_6449);
and U6891 (N_6891,N_6435,N_6544);
nand U6892 (N_6892,N_6549,N_6400);
nand U6893 (N_6893,N_6549,N_6478);
and U6894 (N_6894,N_6367,N_6508);
xnor U6895 (N_6895,N_6494,N_6485);
nor U6896 (N_6896,N_6566,N_6332);
nor U6897 (N_6897,N_6407,N_6305);
xor U6898 (N_6898,N_6460,N_6393);
nand U6899 (N_6899,N_6593,N_6458);
nand U6900 (N_6900,N_6669,N_6814);
and U6901 (N_6901,N_6619,N_6679);
nand U6902 (N_6902,N_6738,N_6848);
nand U6903 (N_6903,N_6745,N_6894);
and U6904 (N_6904,N_6634,N_6884);
and U6905 (N_6905,N_6655,N_6881);
xor U6906 (N_6906,N_6701,N_6761);
and U6907 (N_6907,N_6898,N_6660);
nand U6908 (N_6908,N_6739,N_6869);
nand U6909 (N_6909,N_6858,N_6711);
nor U6910 (N_6910,N_6702,N_6666);
nand U6911 (N_6911,N_6801,N_6715);
xnor U6912 (N_6912,N_6762,N_6888);
nand U6913 (N_6913,N_6747,N_6722);
nand U6914 (N_6914,N_6844,N_6657);
nand U6915 (N_6915,N_6718,N_6680);
or U6916 (N_6916,N_6854,N_6707);
nor U6917 (N_6917,N_6827,N_6890);
nor U6918 (N_6918,N_6710,N_6749);
nand U6919 (N_6919,N_6867,N_6704);
and U6920 (N_6920,N_6830,N_6819);
and U6921 (N_6921,N_6615,N_6777);
and U6922 (N_6922,N_6630,N_6729);
xnor U6923 (N_6923,N_6637,N_6682);
nand U6924 (N_6924,N_6863,N_6641);
nor U6925 (N_6925,N_6813,N_6826);
nor U6926 (N_6926,N_6638,N_6636);
xor U6927 (N_6927,N_6778,N_6652);
nand U6928 (N_6928,N_6610,N_6705);
xnor U6929 (N_6929,N_6767,N_6783);
nand U6930 (N_6930,N_6656,N_6732);
or U6931 (N_6931,N_6880,N_6727);
and U6932 (N_6932,N_6866,N_6623);
xor U6933 (N_6933,N_6845,N_6803);
xor U6934 (N_6934,N_6627,N_6720);
nor U6935 (N_6935,N_6784,N_6786);
nor U6936 (N_6936,N_6685,N_6790);
xnor U6937 (N_6937,N_6736,N_6769);
nor U6938 (N_6938,N_6811,N_6808);
or U6939 (N_6939,N_6741,N_6797);
nor U6940 (N_6940,N_6671,N_6649);
or U6941 (N_6941,N_6635,N_6675);
or U6942 (N_6942,N_6896,N_6795);
xnor U6943 (N_6943,N_6820,N_6658);
and U6944 (N_6944,N_6601,N_6686);
nor U6945 (N_6945,N_6735,N_6774);
nand U6946 (N_6946,N_6626,N_6792);
nor U6947 (N_6947,N_6763,N_6708);
and U6948 (N_6948,N_6677,N_6726);
nor U6949 (N_6949,N_6815,N_6743);
and U6950 (N_6950,N_6633,N_6640);
or U6951 (N_6951,N_6800,N_6841);
nor U6952 (N_6952,N_6843,N_6609);
or U6953 (N_6953,N_6746,N_6689);
nand U6954 (N_6954,N_6611,N_6837);
nor U6955 (N_6955,N_6628,N_6759);
xor U6956 (N_6956,N_6833,N_6676);
or U6957 (N_6957,N_6842,N_6629);
xor U6958 (N_6958,N_6737,N_6631);
nor U6959 (N_6959,N_6731,N_6799);
or U6960 (N_6960,N_6753,N_6852);
xor U6961 (N_6961,N_6603,N_6754);
nor U6962 (N_6962,N_6696,N_6807);
nand U6963 (N_6963,N_6796,N_6846);
or U6964 (N_6964,N_6706,N_6692);
or U6965 (N_6965,N_6836,N_6674);
nor U6966 (N_6966,N_6829,N_6771);
nand U6967 (N_6967,N_6804,N_6606);
and U6968 (N_6968,N_6703,N_6664);
or U6969 (N_6969,N_6895,N_6602);
or U6970 (N_6970,N_6768,N_6873);
nor U6971 (N_6971,N_6672,N_6639);
nor U6972 (N_6972,N_6622,N_6600);
or U6973 (N_6973,N_6748,N_6875);
and U6974 (N_6974,N_6782,N_6744);
or U6975 (N_6975,N_6750,N_6613);
and U6976 (N_6976,N_6770,N_6802);
nor U6977 (N_6977,N_6861,N_6607);
nor U6978 (N_6978,N_6690,N_6870);
xnor U6979 (N_6979,N_6766,N_6765);
nor U6980 (N_6980,N_6616,N_6724);
nor U6981 (N_6981,N_6709,N_6862);
xor U6982 (N_6982,N_6721,N_6728);
or U6983 (N_6983,N_6806,N_6693);
and U6984 (N_6984,N_6899,N_6828);
xor U6985 (N_6985,N_6825,N_6624);
and U6986 (N_6986,N_6835,N_6856);
and U6987 (N_6987,N_6699,N_6752);
nand U6988 (N_6988,N_6719,N_6642);
nand U6989 (N_6989,N_6772,N_6882);
nand U6990 (N_6990,N_6860,N_6687);
and U6991 (N_6991,N_6805,N_6662);
and U6992 (N_6992,N_6789,N_6618);
and U6993 (N_6993,N_6614,N_6876);
nand U6994 (N_6994,N_6822,N_6794);
and U6995 (N_6995,N_6716,N_6650);
or U6996 (N_6996,N_6647,N_6791);
nor U6997 (N_6997,N_6665,N_6612);
nor U6998 (N_6998,N_6868,N_6851);
nand U6999 (N_6999,N_6877,N_6648);
xor U7000 (N_7000,N_6700,N_6793);
nor U7001 (N_7001,N_6857,N_6779);
nand U7002 (N_7002,N_6646,N_6760);
nand U7003 (N_7003,N_6823,N_6834);
nand U7004 (N_7004,N_6764,N_6859);
nand U7005 (N_7005,N_6818,N_6824);
nand U7006 (N_7006,N_6809,N_6733);
nand U7007 (N_7007,N_6663,N_6751);
or U7008 (N_7008,N_6865,N_6812);
xor U7009 (N_7009,N_6864,N_6605);
nor U7010 (N_7010,N_6713,N_6872);
or U7011 (N_7011,N_6668,N_6821);
and U7012 (N_7012,N_6617,N_6853);
and U7013 (N_7013,N_6810,N_6740);
and U7014 (N_7014,N_6697,N_6885);
nand U7015 (N_7015,N_6698,N_6840);
or U7016 (N_7016,N_6776,N_6887);
and U7017 (N_7017,N_6678,N_6667);
nand U7018 (N_7018,N_6625,N_6742);
nand U7019 (N_7019,N_6781,N_6758);
nand U7020 (N_7020,N_6897,N_6798);
and U7021 (N_7021,N_6832,N_6608);
nand U7022 (N_7022,N_6757,N_6734);
and U7023 (N_7023,N_6816,N_6654);
or U7024 (N_7024,N_6714,N_6688);
xor U7025 (N_7025,N_6879,N_6847);
and U7026 (N_7026,N_6670,N_6785);
nor U7027 (N_7027,N_6695,N_6780);
nand U7028 (N_7028,N_6756,N_6883);
nor U7029 (N_7029,N_6838,N_6775);
nand U7030 (N_7030,N_6691,N_6694);
and U7031 (N_7031,N_6892,N_6681);
or U7032 (N_7032,N_6683,N_6730);
nand U7033 (N_7033,N_6817,N_6725);
xor U7034 (N_7034,N_6849,N_6893);
nand U7035 (N_7035,N_6788,N_6717);
or U7036 (N_7036,N_6604,N_6661);
nand U7037 (N_7037,N_6755,N_6653);
or U7038 (N_7038,N_6889,N_6850);
xor U7039 (N_7039,N_6644,N_6839);
nand U7040 (N_7040,N_6891,N_6643);
nand U7041 (N_7041,N_6773,N_6645);
nor U7042 (N_7042,N_6659,N_6723);
nand U7043 (N_7043,N_6673,N_6620);
nor U7044 (N_7044,N_6621,N_6874);
nor U7045 (N_7045,N_6684,N_6871);
nand U7046 (N_7046,N_6855,N_6878);
xnor U7047 (N_7047,N_6632,N_6831);
nor U7048 (N_7048,N_6712,N_6886);
nor U7049 (N_7049,N_6787,N_6651);
and U7050 (N_7050,N_6808,N_6635);
and U7051 (N_7051,N_6790,N_6888);
xor U7052 (N_7052,N_6681,N_6896);
nand U7053 (N_7053,N_6602,N_6859);
nand U7054 (N_7054,N_6773,N_6640);
nor U7055 (N_7055,N_6656,N_6810);
nor U7056 (N_7056,N_6885,N_6613);
nor U7057 (N_7057,N_6662,N_6762);
and U7058 (N_7058,N_6772,N_6667);
nand U7059 (N_7059,N_6841,N_6891);
nor U7060 (N_7060,N_6843,N_6803);
xnor U7061 (N_7061,N_6883,N_6781);
or U7062 (N_7062,N_6859,N_6653);
xor U7063 (N_7063,N_6638,N_6808);
or U7064 (N_7064,N_6656,N_6678);
nor U7065 (N_7065,N_6723,N_6764);
and U7066 (N_7066,N_6661,N_6718);
nor U7067 (N_7067,N_6877,N_6637);
and U7068 (N_7068,N_6849,N_6778);
xor U7069 (N_7069,N_6621,N_6701);
nor U7070 (N_7070,N_6603,N_6718);
and U7071 (N_7071,N_6845,N_6671);
or U7072 (N_7072,N_6645,N_6744);
or U7073 (N_7073,N_6699,N_6773);
nand U7074 (N_7074,N_6656,N_6637);
nand U7075 (N_7075,N_6816,N_6801);
nand U7076 (N_7076,N_6788,N_6619);
and U7077 (N_7077,N_6865,N_6837);
and U7078 (N_7078,N_6683,N_6668);
nand U7079 (N_7079,N_6795,N_6773);
xor U7080 (N_7080,N_6845,N_6713);
nand U7081 (N_7081,N_6867,N_6871);
xor U7082 (N_7082,N_6689,N_6606);
and U7083 (N_7083,N_6663,N_6661);
and U7084 (N_7084,N_6633,N_6787);
and U7085 (N_7085,N_6887,N_6663);
xnor U7086 (N_7086,N_6636,N_6623);
nand U7087 (N_7087,N_6826,N_6606);
xor U7088 (N_7088,N_6856,N_6740);
or U7089 (N_7089,N_6646,N_6703);
xnor U7090 (N_7090,N_6805,N_6775);
and U7091 (N_7091,N_6749,N_6688);
nand U7092 (N_7092,N_6631,N_6772);
and U7093 (N_7093,N_6791,N_6875);
or U7094 (N_7094,N_6799,N_6891);
or U7095 (N_7095,N_6896,N_6654);
or U7096 (N_7096,N_6854,N_6612);
and U7097 (N_7097,N_6818,N_6863);
and U7098 (N_7098,N_6712,N_6867);
xor U7099 (N_7099,N_6789,N_6823);
nand U7100 (N_7100,N_6743,N_6806);
nor U7101 (N_7101,N_6822,N_6709);
nand U7102 (N_7102,N_6790,N_6805);
and U7103 (N_7103,N_6788,N_6699);
xor U7104 (N_7104,N_6668,N_6763);
nor U7105 (N_7105,N_6880,N_6856);
xor U7106 (N_7106,N_6630,N_6879);
and U7107 (N_7107,N_6642,N_6704);
xor U7108 (N_7108,N_6641,N_6683);
nand U7109 (N_7109,N_6604,N_6727);
and U7110 (N_7110,N_6857,N_6626);
nand U7111 (N_7111,N_6749,N_6725);
nor U7112 (N_7112,N_6827,N_6882);
and U7113 (N_7113,N_6858,N_6645);
nand U7114 (N_7114,N_6828,N_6657);
nand U7115 (N_7115,N_6645,N_6822);
or U7116 (N_7116,N_6662,N_6658);
xor U7117 (N_7117,N_6739,N_6824);
xor U7118 (N_7118,N_6819,N_6766);
and U7119 (N_7119,N_6753,N_6880);
nand U7120 (N_7120,N_6756,N_6751);
or U7121 (N_7121,N_6886,N_6831);
xnor U7122 (N_7122,N_6716,N_6865);
or U7123 (N_7123,N_6857,N_6712);
xor U7124 (N_7124,N_6759,N_6719);
xnor U7125 (N_7125,N_6687,N_6652);
or U7126 (N_7126,N_6833,N_6858);
nor U7127 (N_7127,N_6841,N_6838);
or U7128 (N_7128,N_6847,N_6766);
and U7129 (N_7129,N_6715,N_6792);
or U7130 (N_7130,N_6711,N_6607);
nor U7131 (N_7131,N_6714,N_6897);
and U7132 (N_7132,N_6707,N_6804);
xnor U7133 (N_7133,N_6788,N_6848);
xor U7134 (N_7134,N_6883,N_6825);
xnor U7135 (N_7135,N_6664,N_6829);
xnor U7136 (N_7136,N_6600,N_6707);
and U7137 (N_7137,N_6735,N_6739);
xnor U7138 (N_7138,N_6874,N_6834);
or U7139 (N_7139,N_6693,N_6644);
xnor U7140 (N_7140,N_6707,N_6643);
and U7141 (N_7141,N_6752,N_6684);
nor U7142 (N_7142,N_6814,N_6655);
nand U7143 (N_7143,N_6821,N_6751);
xor U7144 (N_7144,N_6759,N_6732);
or U7145 (N_7145,N_6859,N_6844);
or U7146 (N_7146,N_6749,N_6839);
xor U7147 (N_7147,N_6852,N_6761);
nor U7148 (N_7148,N_6645,N_6621);
nand U7149 (N_7149,N_6801,N_6842);
or U7150 (N_7150,N_6768,N_6791);
or U7151 (N_7151,N_6607,N_6646);
and U7152 (N_7152,N_6829,N_6699);
nand U7153 (N_7153,N_6838,N_6766);
nand U7154 (N_7154,N_6762,N_6694);
nand U7155 (N_7155,N_6790,N_6625);
nor U7156 (N_7156,N_6892,N_6663);
and U7157 (N_7157,N_6779,N_6801);
nand U7158 (N_7158,N_6632,N_6660);
nor U7159 (N_7159,N_6695,N_6601);
nor U7160 (N_7160,N_6686,N_6767);
xnor U7161 (N_7161,N_6719,N_6819);
nand U7162 (N_7162,N_6650,N_6854);
or U7163 (N_7163,N_6715,N_6617);
nand U7164 (N_7164,N_6844,N_6639);
nor U7165 (N_7165,N_6690,N_6646);
xnor U7166 (N_7166,N_6659,N_6704);
or U7167 (N_7167,N_6613,N_6816);
or U7168 (N_7168,N_6862,N_6736);
and U7169 (N_7169,N_6716,N_6823);
xor U7170 (N_7170,N_6611,N_6734);
and U7171 (N_7171,N_6613,N_6655);
and U7172 (N_7172,N_6705,N_6688);
and U7173 (N_7173,N_6818,N_6719);
and U7174 (N_7174,N_6832,N_6750);
nand U7175 (N_7175,N_6850,N_6738);
xor U7176 (N_7176,N_6722,N_6605);
xnor U7177 (N_7177,N_6682,N_6734);
and U7178 (N_7178,N_6778,N_6879);
nand U7179 (N_7179,N_6898,N_6755);
or U7180 (N_7180,N_6666,N_6701);
xnor U7181 (N_7181,N_6638,N_6631);
nor U7182 (N_7182,N_6701,N_6655);
xor U7183 (N_7183,N_6825,N_6747);
or U7184 (N_7184,N_6757,N_6876);
or U7185 (N_7185,N_6864,N_6829);
and U7186 (N_7186,N_6824,N_6658);
nand U7187 (N_7187,N_6650,N_6798);
nand U7188 (N_7188,N_6779,N_6606);
xor U7189 (N_7189,N_6801,N_6866);
and U7190 (N_7190,N_6699,N_6842);
xnor U7191 (N_7191,N_6683,N_6799);
nand U7192 (N_7192,N_6765,N_6716);
or U7193 (N_7193,N_6769,N_6866);
nor U7194 (N_7194,N_6653,N_6713);
xnor U7195 (N_7195,N_6641,N_6820);
nor U7196 (N_7196,N_6803,N_6607);
or U7197 (N_7197,N_6703,N_6872);
or U7198 (N_7198,N_6658,N_6649);
nand U7199 (N_7199,N_6751,N_6879);
xnor U7200 (N_7200,N_7163,N_6934);
nor U7201 (N_7201,N_7170,N_6926);
nor U7202 (N_7202,N_6979,N_6918);
and U7203 (N_7203,N_6971,N_7083);
nor U7204 (N_7204,N_7092,N_7022);
xor U7205 (N_7205,N_7137,N_7065);
xor U7206 (N_7206,N_7082,N_7043);
or U7207 (N_7207,N_7101,N_6915);
nand U7208 (N_7208,N_6951,N_7139);
nor U7209 (N_7209,N_7070,N_7089);
nor U7210 (N_7210,N_7106,N_7013);
xnor U7211 (N_7211,N_7091,N_6916);
and U7212 (N_7212,N_7125,N_7141);
nand U7213 (N_7213,N_7186,N_6923);
nand U7214 (N_7214,N_7134,N_7105);
and U7215 (N_7215,N_7197,N_7059);
or U7216 (N_7216,N_7174,N_7066);
nor U7217 (N_7217,N_6922,N_7078);
or U7218 (N_7218,N_6983,N_6940);
nor U7219 (N_7219,N_7159,N_6938);
nor U7220 (N_7220,N_7138,N_6998);
nand U7221 (N_7221,N_6995,N_6921);
and U7222 (N_7222,N_7054,N_7171);
and U7223 (N_7223,N_7195,N_6949);
nor U7224 (N_7224,N_7148,N_7079);
or U7225 (N_7225,N_7098,N_7194);
nand U7226 (N_7226,N_6948,N_7072);
and U7227 (N_7227,N_6912,N_7073);
nor U7228 (N_7228,N_6978,N_6937);
or U7229 (N_7229,N_6989,N_7165);
and U7230 (N_7230,N_7085,N_7025);
and U7231 (N_7231,N_7129,N_6950);
or U7232 (N_7232,N_7113,N_7185);
or U7233 (N_7233,N_7011,N_7131);
xor U7234 (N_7234,N_7150,N_6906);
nand U7235 (N_7235,N_6924,N_7050);
nor U7236 (N_7236,N_7009,N_7180);
and U7237 (N_7237,N_6944,N_7031);
nor U7238 (N_7238,N_7177,N_7124);
xor U7239 (N_7239,N_7046,N_7107);
nand U7240 (N_7240,N_7119,N_7196);
and U7241 (N_7241,N_6980,N_7084);
xor U7242 (N_7242,N_7029,N_7051);
and U7243 (N_7243,N_7183,N_7127);
and U7244 (N_7244,N_6900,N_6975);
and U7245 (N_7245,N_6928,N_6930);
nand U7246 (N_7246,N_7087,N_7143);
nand U7247 (N_7247,N_7156,N_6917);
xnor U7248 (N_7248,N_6935,N_6919);
or U7249 (N_7249,N_6984,N_7169);
nor U7250 (N_7250,N_7023,N_6943);
nand U7251 (N_7251,N_7007,N_6972);
xor U7252 (N_7252,N_7077,N_7094);
nand U7253 (N_7253,N_6985,N_7162);
and U7254 (N_7254,N_6909,N_6960);
xor U7255 (N_7255,N_7118,N_7157);
nor U7256 (N_7256,N_7096,N_7088);
xor U7257 (N_7257,N_7151,N_6974);
and U7258 (N_7258,N_7116,N_7075);
xor U7259 (N_7259,N_7130,N_6902);
xor U7260 (N_7260,N_6920,N_6933);
or U7261 (N_7261,N_6999,N_7004);
and U7262 (N_7262,N_7112,N_7115);
or U7263 (N_7263,N_7018,N_6904);
nor U7264 (N_7264,N_6947,N_6908);
or U7265 (N_7265,N_7010,N_6970);
or U7266 (N_7266,N_7161,N_7049);
and U7267 (N_7267,N_7047,N_6955);
xor U7268 (N_7268,N_6941,N_7095);
xor U7269 (N_7269,N_7061,N_7190);
nor U7270 (N_7270,N_7037,N_7117);
or U7271 (N_7271,N_7027,N_7168);
nor U7272 (N_7272,N_7193,N_6976);
xor U7273 (N_7273,N_7048,N_6953);
xnor U7274 (N_7274,N_7060,N_7071);
nor U7275 (N_7275,N_7160,N_7142);
and U7276 (N_7276,N_6986,N_7104);
nor U7277 (N_7277,N_6961,N_7012);
nand U7278 (N_7278,N_7017,N_7015);
xor U7279 (N_7279,N_7145,N_7097);
or U7280 (N_7280,N_7053,N_7103);
nor U7281 (N_7281,N_7064,N_6992);
and U7282 (N_7282,N_7136,N_6965);
and U7283 (N_7283,N_7147,N_7020);
nand U7284 (N_7284,N_6942,N_7038);
or U7285 (N_7285,N_7099,N_7086);
or U7286 (N_7286,N_7149,N_7114);
and U7287 (N_7287,N_7080,N_6968);
nand U7288 (N_7288,N_7014,N_6996);
and U7289 (N_7289,N_7030,N_6959);
and U7290 (N_7290,N_7035,N_7006);
and U7291 (N_7291,N_7167,N_7155);
nand U7292 (N_7292,N_7135,N_6952);
and U7293 (N_7293,N_6997,N_7032);
nor U7294 (N_7294,N_7069,N_7172);
and U7295 (N_7295,N_7178,N_7121);
nand U7296 (N_7296,N_7001,N_7154);
or U7297 (N_7297,N_7021,N_6969);
or U7298 (N_7298,N_7179,N_7166);
nand U7299 (N_7299,N_7133,N_6977);
xor U7300 (N_7300,N_7000,N_6946);
and U7301 (N_7301,N_6962,N_7164);
xor U7302 (N_7302,N_6963,N_6987);
and U7303 (N_7303,N_6973,N_7074);
and U7304 (N_7304,N_6954,N_7120);
nand U7305 (N_7305,N_7040,N_6964);
and U7306 (N_7306,N_7144,N_7192);
nor U7307 (N_7307,N_7034,N_7184);
and U7308 (N_7308,N_7140,N_6931);
xor U7309 (N_7309,N_7005,N_6939);
nand U7310 (N_7310,N_7057,N_7076);
or U7311 (N_7311,N_7100,N_7056);
nand U7312 (N_7312,N_7052,N_7158);
nor U7313 (N_7313,N_7081,N_7126);
nand U7314 (N_7314,N_7041,N_7122);
or U7315 (N_7315,N_7039,N_6907);
nand U7316 (N_7316,N_6988,N_7090);
or U7317 (N_7317,N_7175,N_6967);
and U7318 (N_7318,N_7189,N_6910);
xnor U7319 (N_7319,N_7123,N_7068);
nor U7320 (N_7320,N_7062,N_7187);
nor U7321 (N_7321,N_7063,N_7199);
xnor U7322 (N_7322,N_7067,N_7191);
and U7323 (N_7323,N_7044,N_6903);
and U7324 (N_7324,N_7055,N_6993);
nand U7325 (N_7325,N_6945,N_7146);
nand U7326 (N_7326,N_7153,N_7033);
nand U7327 (N_7327,N_7111,N_6929);
or U7328 (N_7328,N_6925,N_6966);
or U7329 (N_7329,N_7024,N_7016);
nand U7330 (N_7330,N_6913,N_7019);
nand U7331 (N_7331,N_6911,N_6982);
or U7332 (N_7332,N_6994,N_6901);
or U7333 (N_7333,N_7093,N_7058);
xnor U7334 (N_7334,N_7182,N_7152);
nor U7335 (N_7335,N_7008,N_7042);
and U7336 (N_7336,N_7045,N_7109);
and U7337 (N_7337,N_7026,N_7173);
and U7338 (N_7338,N_7128,N_6905);
xor U7339 (N_7339,N_6932,N_6981);
nor U7340 (N_7340,N_7176,N_7132);
nor U7341 (N_7341,N_6927,N_7188);
xnor U7342 (N_7342,N_6914,N_7028);
or U7343 (N_7343,N_6991,N_6957);
nor U7344 (N_7344,N_6990,N_7198);
nand U7345 (N_7345,N_7108,N_7110);
and U7346 (N_7346,N_7002,N_6958);
and U7347 (N_7347,N_6956,N_7036);
nor U7348 (N_7348,N_7102,N_7003);
xnor U7349 (N_7349,N_6936,N_7181);
nor U7350 (N_7350,N_7154,N_6975);
and U7351 (N_7351,N_6989,N_6916);
xor U7352 (N_7352,N_7103,N_7164);
and U7353 (N_7353,N_7125,N_7171);
or U7354 (N_7354,N_7077,N_6946);
nor U7355 (N_7355,N_6934,N_6933);
nand U7356 (N_7356,N_6945,N_6994);
xnor U7357 (N_7357,N_6914,N_6985);
or U7358 (N_7358,N_6976,N_7070);
xor U7359 (N_7359,N_6912,N_7096);
xnor U7360 (N_7360,N_7104,N_7135);
xor U7361 (N_7361,N_7128,N_7181);
nand U7362 (N_7362,N_7068,N_7059);
nand U7363 (N_7363,N_7118,N_7145);
nor U7364 (N_7364,N_7151,N_7155);
nand U7365 (N_7365,N_7043,N_7171);
or U7366 (N_7366,N_6967,N_6983);
nor U7367 (N_7367,N_7092,N_6988);
or U7368 (N_7368,N_7189,N_7197);
and U7369 (N_7369,N_7120,N_6961);
or U7370 (N_7370,N_7090,N_7159);
nand U7371 (N_7371,N_6961,N_7014);
and U7372 (N_7372,N_7100,N_7084);
and U7373 (N_7373,N_7053,N_7086);
xnor U7374 (N_7374,N_7175,N_7144);
nand U7375 (N_7375,N_6973,N_7021);
nor U7376 (N_7376,N_7195,N_7041);
xnor U7377 (N_7377,N_6927,N_6962);
nand U7378 (N_7378,N_7049,N_7073);
nand U7379 (N_7379,N_6924,N_6967);
nor U7380 (N_7380,N_7039,N_6923);
and U7381 (N_7381,N_7042,N_7153);
nor U7382 (N_7382,N_6933,N_6984);
xor U7383 (N_7383,N_7007,N_7054);
xor U7384 (N_7384,N_7065,N_7026);
or U7385 (N_7385,N_7148,N_7063);
xor U7386 (N_7386,N_6909,N_7114);
nand U7387 (N_7387,N_7061,N_6906);
nand U7388 (N_7388,N_6919,N_7171);
nand U7389 (N_7389,N_7106,N_7119);
nor U7390 (N_7390,N_7097,N_6939);
nand U7391 (N_7391,N_7159,N_6902);
and U7392 (N_7392,N_7198,N_6954);
nor U7393 (N_7393,N_7187,N_7142);
and U7394 (N_7394,N_6969,N_7164);
and U7395 (N_7395,N_6926,N_7149);
and U7396 (N_7396,N_6900,N_7135);
xnor U7397 (N_7397,N_7030,N_7084);
xnor U7398 (N_7398,N_6913,N_7138);
nor U7399 (N_7399,N_7131,N_7165);
and U7400 (N_7400,N_7132,N_6947);
nand U7401 (N_7401,N_7142,N_7158);
nand U7402 (N_7402,N_7060,N_7150);
nor U7403 (N_7403,N_6919,N_7075);
nand U7404 (N_7404,N_7024,N_7051);
or U7405 (N_7405,N_6902,N_6968);
nand U7406 (N_7406,N_7194,N_7004);
and U7407 (N_7407,N_7036,N_7056);
and U7408 (N_7408,N_7106,N_7072);
nor U7409 (N_7409,N_6923,N_7104);
or U7410 (N_7410,N_7160,N_6992);
and U7411 (N_7411,N_6928,N_7067);
nand U7412 (N_7412,N_7046,N_7088);
nand U7413 (N_7413,N_6978,N_7140);
and U7414 (N_7414,N_7047,N_6903);
or U7415 (N_7415,N_6984,N_7187);
nand U7416 (N_7416,N_7045,N_6905);
xnor U7417 (N_7417,N_7150,N_7139);
nor U7418 (N_7418,N_7117,N_6908);
nand U7419 (N_7419,N_7186,N_7159);
and U7420 (N_7420,N_7071,N_7026);
and U7421 (N_7421,N_6912,N_6992);
nor U7422 (N_7422,N_7116,N_6972);
nor U7423 (N_7423,N_6932,N_7021);
nand U7424 (N_7424,N_7075,N_7155);
nor U7425 (N_7425,N_7007,N_6979);
nor U7426 (N_7426,N_7130,N_6903);
or U7427 (N_7427,N_7139,N_7028);
nand U7428 (N_7428,N_6930,N_6993);
or U7429 (N_7429,N_6973,N_6960);
nand U7430 (N_7430,N_7162,N_7197);
and U7431 (N_7431,N_6941,N_7171);
or U7432 (N_7432,N_7102,N_7013);
or U7433 (N_7433,N_6958,N_7082);
nand U7434 (N_7434,N_6981,N_6940);
nand U7435 (N_7435,N_6993,N_7059);
and U7436 (N_7436,N_7047,N_7033);
nand U7437 (N_7437,N_7051,N_7095);
xnor U7438 (N_7438,N_7102,N_7084);
xnor U7439 (N_7439,N_7128,N_6997);
xor U7440 (N_7440,N_7161,N_7045);
and U7441 (N_7441,N_6936,N_7048);
xor U7442 (N_7442,N_7022,N_7046);
or U7443 (N_7443,N_7070,N_7146);
xor U7444 (N_7444,N_7069,N_7132);
and U7445 (N_7445,N_7110,N_6914);
xor U7446 (N_7446,N_6932,N_7049);
nand U7447 (N_7447,N_7094,N_6960);
or U7448 (N_7448,N_7060,N_7033);
and U7449 (N_7449,N_7031,N_6987);
or U7450 (N_7450,N_7125,N_7074);
and U7451 (N_7451,N_7014,N_7193);
nand U7452 (N_7452,N_6941,N_7088);
xor U7453 (N_7453,N_7027,N_6950);
or U7454 (N_7454,N_6928,N_6963);
nand U7455 (N_7455,N_6987,N_6948);
xor U7456 (N_7456,N_6901,N_7145);
xor U7457 (N_7457,N_6983,N_7070);
xnor U7458 (N_7458,N_6951,N_7060);
and U7459 (N_7459,N_7114,N_7091);
and U7460 (N_7460,N_6971,N_7026);
nor U7461 (N_7461,N_7066,N_7172);
xor U7462 (N_7462,N_6974,N_7080);
xnor U7463 (N_7463,N_6921,N_7072);
nand U7464 (N_7464,N_7033,N_6919);
xor U7465 (N_7465,N_7106,N_7142);
or U7466 (N_7466,N_7011,N_6936);
nand U7467 (N_7467,N_6960,N_7113);
nor U7468 (N_7468,N_7041,N_7159);
xor U7469 (N_7469,N_7138,N_7043);
nor U7470 (N_7470,N_7114,N_6939);
nand U7471 (N_7471,N_7009,N_6966);
and U7472 (N_7472,N_7191,N_6953);
xor U7473 (N_7473,N_6923,N_7068);
or U7474 (N_7474,N_7075,N_6993);
nand U7475 (N_7475,N_7141,N_6934);
and U7476 (N_7476,N_7010,N_7090);
nor U7477 (N_7477,N_6930,N_7182);
or U7478 (N_7478,N_6981,N_6912);
xnor U7479 (N_7479,N_6938,N_7181);
nand U7480 (N_7480,N_6913,N_7157);
nand U7481 (N_7481,N_7188,N_6953);
nor U7482 (N_7482,N_7007,N_7089);
nor U7483 (N_7483,N_7026,N_7193);
nand U7484 (N_7484,N_7169,N_6996);
nand U7485 (N_7485,N_7106,N_7015);
and U7486 (N_7486,N_6990,N_6992);
nor U7487 (N_7487,N_7029,N_6907);
nand U7488 (N_7488,N_7143,N_6907);
or U7489 (N_7489,N_7109,N_7094);
and U7490 (N_7490,N_7155,N_7071);
nand U7491 (N_7491,N_7178,N_6987);
or U7492 (N_7492,N_7018,N_6965);
nand U7493 (N_7493,N_6999,N_7001);
nand U7494 (N_7494,N_7008,N_6964);
xor U7495 (N_7495,N_7051,N_6960);
nand U7496 (N_7496,N_7088,N_7140);
and U7497 (N_7497,N_6952,N_7165);
or U7498 (N_7498,N_7001,N_7070);
nand U7499 (N_7499,N_7158,N_6931);
xnor U7500 (N_7500,N_7287,N_7239);
xor U7501 (N_7501,N_7223,N_7251);
nor U7502 (N_7502,N_7237,N_7497);
and U7503 (N_7503,N_7387,N_7364);
nor U7504 (N_7504,N_7241,N_7461);
nor U7505 (N_7505,N_7398,N_7310);
nand U7506 (N_7506,N_7431,N_7325);
and U7507 (N_7507,N_7238,N_7205);
nor U7508 (N_7508,N_7372,N_7361);
nand U7509 (N_7509,N_7427,N_7301);
nor U7510 (N_7510,N_7424,N_7496);
nor U7511 (N_7511,N_7343,N_7475);
nand U7512 (N_7512,N_7440,N_7304);
nor U7513 (N_7513,N_7204,N_7377);
nor U7514 (N_7514,N_7299,N_7286);
or U7515 (N_7515,N_7344,N_7282);
xor U7516 (N_7516,N_7438,N_7315);
and U7517 (N_7517,N_7337,N_7406);
nor U7518 (N_7518,N_7484,N_7376);
nor U7519 (N_7519,N_7278,N_7249);
nor U7520 (N_7520,N_7303,N_7358);
xor U7521 (N_7521,N_7452,N_7355);
nand U7522 (N_7522,N_7467,N_7260);
xnor U7523 (N_7523,N_7378,N_7430);
xnor U7524 (N_7524,N_7384,N_7478);
nand U7525 (N_7525,N_7371,N_7367);
nor U7526 (N_7526,N_7397,N_7353);
or U7527 (N_7527,N_7492,N_7485);
nor U7528 (N_7528,N_7487,N_7422);
nor U7529 (N_7529,N_7225,N_7469);
and U7530 (N_7530,N_7476,N_7436);
and U7531 (N_7531,N_7334,N_7365);
or U7532 (N_7532,N_7449,N_7221);
nor U7533 (N_7533,N_7488,N_7292);
xnor U7534 (N_7534,N_7454,N_7414);
nor U7535 (N_7535,N_7354,N_7296);
and U7536 (N_7536,N_7336,N_7226);
nor U7537 (N_7537,N_7392,N_7255);
and U7538 (N_7538,N_7227,N_7470);
or U7539 (N_7539,N_7389,N_7335);
and U7540 (N_7540,N_7435,N_7493);
xnor U7541 (N_7541,N_7311,N_7274);
xnor U7542 (N_7542,N_7419,N_7222);
nand U7543 (N_7543,N_7284,N_7429);
or U7544 (N_7544,N_7434,N_7327);
or U7545 (N_7545,N_7349,N_7374);
and U7546 (N_7546,N_7236,N_7329);
xnor U7547 (N_7547,N_7481,N_7425);
nor U7548 (N_7548,N_7277,N_7402);
and U7549 (N_7549,N_7360,N_7230);
nor U7550 (N_7550,N_7348,N_7298);
and U7551 (N_7551,N_7441,N_7280);
and U7552 (N_7552,N_7499,N_7339);
nor U7553 (N_7553,N_7346,N_7331);
nor U7554 (N_7554,N_7391,N_7269);
xor U7555 (N_7555,N_7231,N_7285);
xor U7556 (N_7556,N_7258,N_7480);
or U7557 (N_7557,N_7482,N_7383);
or U7558 (N_7558,N_7347,N_7256);
nor U7559 (N_7559,N_7297,N_7432);
nor U7560 (N_7560,N_7279,N_7302);
nand U7561 (N_7561,N_7330,N_7243);
nor U7562 (N_7562,N_7382,N_7323);
xor U7563 (N_7563,N_7314,N_7240);
and U7564 (N_7564,N_7386,N_7345);
nand U7565 (N_7565,N_7291,N_7281);
or U7566 (N_7566,N_7445,N_7465);
xor U7567 (N_7567,N_7413,N_7201);
xor U7568 (N_7568,N_7443,N_7381);
or U7569 (N_7569,N_7477,N_7246);
xnor U7570 (N_7570,N_7217,N_7490);
or U7571 (N_7571,N_7351,N_7271);
nor U7572 (N_7572,N_7210,N_7459);
nand U7573 (N_7573,N_7234,N_7404);
xnor U7574 (N_7574,N_7312,N_7232);
xor U7575 (N_7575,N_7207,N_7228);
or U7576 (N_7576,N_7437,N_7316);
xor U7577 (N_7577,N_7396,N_7270);
nand U7578 (N_7578,N_7408,N_7261);
xnor U7579 (N_7579,N_7498,N_7420);
nand U7580 (N_7580,N_7211,N_7220);
xor U7581 (N_7581,N_7242,N_7446);
xor U7582 (N_7582,N_7410,N_7357);
and U7583 (N_7583,N_7495,N_7321);
nor U7584 (N_7584,N_7305,N_7244);
nor U7585 (N_7585,N_7341,N_7486);
xor U7586 (N_7586,N_7328,N_7268);
or U7587 (N_7587,N_7363,N_7411);
or U7588 (N_7588,N_7288,N_7473);
nand U7589 (N_7589,N_7373,N_7426);
xor U7590 (N_7590,N_7460,N_7313);
nor U7591 (N_7591,N_7380,N_7370);
and U7592 (N_7592,N_7368,N_7212);
nand U7593 (N_7593,N_7267,N_7324);
or U7594 (N_7594,N_7421,N_7252);
nor U7595 (N_7595,N_7474,N_7393);
nor U7596 (N_7596,N_7362,N_7448);
nor U7597 (N_7597,N_7338,N_7433);
nand U7598 (N_7598,N_7456,N_7253);
xnor U7599 (N_7599,N_7352,N_7293);
and U7600 (N_7600,N_7215,N_7333);
nor U7601 (N_7601,N_7219,N_7428);
nand U7602 (N_7602,N_7483,N_7289);
and U7603 (N_7603,N_7388,N_7214);
or U7604 (N_7604,N_7379,N_7229);
or U7605 (N_7605,N_7409,N_7203);
nand U7606 (N_7606,N_7359,N_7318);
and U7607 (N_7607,N_7218,N_7479);
or U7608 (N_7608,N_7290,N_7463);
and U7609 (N_7609,N_7444,N_7399);
and U7610 (N_7610,N_7472,N_7457);
nand U7611 (N_7611,N_7208,N_7202);
nor U7612 (N_7612,N_7262,N_7416);
or U7613 (N_7613,N_7447,N_7466);
nand U7614 (N_7614,N_7342,N_7322);
or U7615 (N_7615,N_7309,N_7412);
xnor U7616 (N_7616,N_7401,N_7400);
xnor U7617 (N_7617,N_7206,N_7350);
and U7618 (N_7618,N_7306,N_7453);
and U7619 (N_7619,N_7439,N_7209);
and U7620 (N_7620,N_7248,N_7369);
xnor U7621 (N_7621,N_7451,N_7471);
and U7622 (N_7622,N_7332,N_7455);
nand U7623 (N_7623,N_7403,N_7462);
xnor U7624 (N_7624,N_7375,N_7235);
and U7625 (N_7625,N_7407,N_7300);
nand U7626 (N_7626,N_7494,N_7319);
nor U7627 (N_7627,N_7307,N_7295);
and U7628 (N_7628,N_7458,N_7405);
and U7629 (N_7629,N_7265,N_7263);
or U7630 (N_7630,N_7200,N_7272);
or U7631 (N_7631,N_7264,N_7213);
nor U7632 (N_7632,N_7418,N_7394);
and U7633 (N_7633,N_7326,N_7395);
xor U7634 (N_7634,N_7250,N_7366);
or U7635 (N_7635,N_7356,N_7442);
and U7636 (N_7636,N_7468,N_7423);
or U7637 (N_7637,N_7275,N_7276);
or U7638 (N_7638,N_7308,N_7417);
xnor U7639 (N_7639,N_7233,N_7489);
nor U7640 (N_7640,N_7294,N_7266);
nand U7641 (N_7641,N_7340,N_7317);
or U7642 (N_7642,N_7390,N_7257);
and U7643 (N_7643,N_7216,N_7464);
xnor U7644 (N_7644,N_7491,N_7450);
nand U7645 (N_7645,N_7224,N_7385);
nor U7646 (N_7646,N_7247,N_7320);
nor U7647 (N_7647,N_7259,N_7415);
and U7648 (N_7648,N_7273,N_7245);
and U7649 (N_7649,N_7254,N_7283);
nor U7650 (N_7650,N_7429,N_7335);
nor U7651 (N_7651,N_7332,N_7493);
and U7652 (N_7652,N_7444,N_7348);
nor U7653 (N_7653,N_7207,N_7215);
or U7654 (N_7654,N_7401,N_7370);
or U7655 (N_7655,N_7347,N_7365);
or U7656 (N_7656,N_7435,N_7219);
or U7657 (N_7657,N_7359,N_7305);
nand U7658 (N_7658,N_7248,N_7271);
and U7659 (N_7659,N_7417,N_7467);
and U7660 (N_7660,N_7411,N_7282);
and U7661 (N_7661,N_7494,N_7233);
and U7662 (N_7662,N_7258,N_7309);
and U7663 (N_7663,N_7261,N_7257);
and U7664 (N_7664,N_7220,N_7372);
or U7665 (N_7665,N_7410,N_7293);
and U7666 (N_7666,N_7397,N_7234);
nand U7667 (N_7667,N_7457,N_7418);
xor U7668 (N_7668,N_7473,N_7309);
and U7669 (N_7669,N_7346,N_7257);
nand U7670 (N_7670,N_7367,N_7270);
and U7671 (N_7671,N_7392,N_7432);
nand U7672 (N_7672,N_7201,N_7282);
xnor U7673 (N_7673,N_7435,N_7394);
or U7674 (N_7674,N_7335,N_7266);
xnor U7675 (N_7675,N_7469,N_7291);
and U7676 (N_7676,N_7251,N_7326);
xnor U7677 (N_7677,N_7484,N_7377);
xnor U7678 (N_7678,N_7479,N_7387);
or U7679 (N_7679,N_7494,N_7343);
or U7680 (N_7680,N_7359,N_7447);
nor U7681 (N_7681,N_7254,N_7451);
nand U7682 (N_7682,N_7439,N_7425);
nor U7683 (N_7683,N_7249,N_7227);
xor U7684 (N_7684,N_7376,N_7458);
nand U7685 (N_7685,N_7276,N_7465);
nor U7686 (N_7686,N_7282,N_7309);
and U7687 (N_7687,N_7354,N_7387);
or U7688 (N_7688,N_7204,N_7357);
nand U7689 (N_7689,N_7447,N_7442);
nor U7690 (N_7690,N_7467,N_7294);
or U7691 (N_7691,N_7279,N_7213);
xor U7692 (N_7692,N_7412,N_7316);
and U7693 (N_7693,N_7374,N_7330);
and U7694 (N_7694,N_7432,N_7224);
xnor U7695 (N_7695,N_7415,N_7261);
or U7696 (N_7696,N_7460,N_7332);
and U7697 (N_7697,N_7296,N_7217);
nand U7698 (N_7698,N_7491,N_7455);
nor U7699 (N_7699,N_7306,N_7290);
xnor U7700 (N_7700,N_7371,N_7386);
or U7701 (N_7701,N_7484,N_7404);
nand U7702 (N_7702,N_7395,N_7324);
nor U7703 (N_7703,N_7389,N_7366);
and U7704 (N_7704,N_7412,N_7410);
or U7705 (N_7705,N_7264,N_7449);
xnor U7706 (N_7706,N_7415,N_7202);
xnor U7707 (N_7707,N_7375,N_7229);
xor U7708 (N_7708,N_7202,N_7372);
xor U7709 (N_7709,N_7296,N_7453);
or U7710 (N_7710,N_7453,N_7303);
nand U7711 (N_7711,N_7279,N_7338);
and U7712 (N_7712,N_7498,N_7390);
xnor U7713 (N_7713,N_7418,N_7212);
nand U7714 (N_7714,N_7295,N_7424);
nand U7715 (N_7715,N_7408,N_7476);
and U7716 (N_7716,N_7376,N_7469);
and U7717 (N_7717,N_7329,N_7408);
nor U7718 (N_7718,N_7498,N_7325);
nor U7719 (N_7719,N_7211,N_7292);
or U7720 (N_7720,N_7492,N_7495);
or U7721 (N_7721,N_7307,N_7242);
nor U7722 (N_7722,N_7408,N_7352);
or U7723 (N_7723,N_7291,N_7300);
xnor U7724 (N_7724,N_7448,N_7410);
xor U7725 (N_7725,N_7399,N_7443);
nor U7726 (N_7726,N_7205,N_7269);
and U7727 (N_7727,N_7429,N_7485);
and U7728 (N_7728,N_7429,N_7436);
and U7729 (N_7729,N_7474,N_7411);
nor U7730 (N_7730,N_7388,N_7385);
nand U7731 (N_7731,N_7301,N_7204);
xnor U7732 (N_7732,N_7267,N_7404);
or U7733 (N_7733,N_7208,N_7234);
nor U7734 (N_7734,N_7319,N_7417);
xnor U7735 (N_7735,N_7232,N_7292);
nand U7736 (N_7736,N_7471,N_7333);
nand U7737 (N_7737,N_7351,N_7439);
and U7738 (N_7738,N_7235,N_7465);
nand U7739 (N_7739,N_7312,N_7474);
and U7740 (N_7740,N_7370,N_7452);
nand U7741 (N_7741,N_7229,N_7228);
and U7742 (N_7742,N_7226,N_7398);
nor U7743 (N_7743,N_7484,N_7494);
nand U7744 (N_7744,N_7385,N_7240);
nor U7745 (N_7745,N_7471,N_7497);
or U7746 (N_7746,N_7397,N_7333);
and U7747 (N_7747,N_7221,N_7219);
xor U7748 (N_7748,N_7250,N_7494);
nor U7749 (N_7749,N_7429,N_7277);
or U7750 (N_7750,N_7403,N_7315);
xor U7751 (N_7751,N_7481,N_7491);
nor U7752 (N_7752,N_7461,N_7226);
and U7753 (N_7753,N_7397,N_7241);
nand U7754 (N_7754,N_7476,N_7421);
and U7755 (N_7755,N_7284,N_7214);
and U7756 (N_7756,N_7292,N_7214);
nor U7757 (N_7757,N_7305,N_7472);
or U7758 (N_7758,N_7402,N_7411);
nor U7759 (N_7759,N_7281,N_7257);
nor U7760 (N_7760,N_7252,N_7459);
or U7761 (N_7761,N_7251,N_7236);
xnor U7762 (N_7762,N_7261,N_7492);
xnor U7763 (N_7763,N_7437,N_7270);
nor U7764 (N_7764,N_7388,N_7290);
nor U7765 (N_7765,N_7364,N_7280);
or U7766 (N_7766,N_7433,N_7363);
nand U7767 (N_7767,N_7430,N_7343);
and U7768 (N_7768,N_7496,N_7450);
or U7769 (N_7769,N_7371,N_7296);
nand U7770 (N_7770,N_7372,N_7446);
nor U7771 (N_7771,N_7487,N_7377);
and U7772 (N_7772,N_7402,N_7226);
nand U7773 (N_7773,N_7379,N_7232);
xor U7774 (N_7774,N_7363,N_7356);
xnor U7775 (N_7775,N_7327,N_7250);
or U7776 (N_7776,N_7415,N_7235);
xnor U7777 (N_7777,N_7275,N_7412);
or U7778 (N_7778,N_7379,N_7411);
nand U7779 (N_7779,N_7402,N_7243);
xnor U7780 (N_7780,N_7272,N_7406);
or U7781 (N_7781,N_7201,N_7456);
and U7782 (N_7782,N_7334,N_7337);
nor U7783 (N_7783,N_7296,N_7437);
and U7784 (N_7784,N_7265,N_7436);
nand U7785 (N_7785,N_7372,N_7379);
nor U7786 (N_7786,N_7461,N_7454);
or U7787 (N_7787,N_7463,N_7300);
nor U7788 (N_7788,N_7441,N_7240);
nand U7789 (N_7789,N_7423,N_7243);
nand U7790 (N_7790,N_7440,N_7263);
or U7791 (N_7791,N_7341,N_7336);
nand U7792 (N_7792,N_7400,N_7357);
nor U7793 (N_7793,N_7340,N_7290);
and U7794 (N_7794,N_7216,N_7299);
and U7795 (N_7795,N_7313,N_7405);
xor U7796 (N_7796,N_7307,N_7429);
or U7797 (N_7797,N_7230,N_7459);
xnor U7798 (N_7798,N_7266,N_7395);
and U7799 (N_7799,N_7248,N_7445);
xnor U7800 (N_7800,N_7747,N_7696);
nand U7801 (N_7801,N_7719,N_7684);
or U7802 (N_7802,N_7725,N_7723);
nand U7803 (N_7803,N_7601,N_7667);
xor U7804 (N_7804,N_7654,N_7637);
and U7805 (N_7805,N_7670,N_7778);
nor U7806 (N_7806,N_7686,N_7539);
or U7807 (N_7807,N_7672,N_7739);
and U7808 (N_7808,N_7578,N_7768);
and U7809 (N_7809,N_7795,N_7634);
xnor U7810 (N_7810,N_7581,N_7512);
nor U7811 (N_7811,N_7614,N_7749);
and U7812 (N_7812,N_7732,N_7730);
xor U7813 (N_7813,N_7577,N_7527);
and U7814 (N_7814,N_7606,N_7751);
and U7815 (N_7815,N_7769,N_7733);
and U7816 (N_7816,N_7510,N_7628);
or U7817 (N_7817,N_7737,N_7515);
or U7818 (N_7818,N_7556,N_7573);
nand U7819 (N_7819,N_7558,N_7677);
and U7820 (N_7820,N_7596,N_7574);
nor U7821 (N_7821,N_7724,N_7655);
nor U7822 (N_7822,N_7509,N_7656);
nand U7823 (N_7823,N_7602,N_7584);
or U7824 (N_7824,N_7507,N_7593);
or U7825 (N_7825,N_7711,N_7542);
nor U7826 (N_7826,N_7715,N_7695);
nor U7827 (N_7827,N_7750,N_7781);
and U7828 (N_7828,N_7618,N_7799);
and U7829 (N_7829,N_7757,N_7566);
nand U7830 (N_7830,N_7666,N_7565);
and U7831 (N_7831,N_7718,N_7599);
nand U7832 (N_7832,N_7752,N_7632);
and U7833 (N_7833,N_7550,N_7740);
or U7834 (N_7834,N_7783,N_7549);
nand U7835 (N_7835,N_7505,N_7728);
nor U7836 (N_7836,N_7793,N_7640);
and U7837 (N_7837,N_7610,N_7533);
or U7838 (N_7838,N_7503,N_7589);
nor U7839 (N_7839,N_7635,N_7780);
nor U7840 (N_7840,N_7540,N_7513);
and U7841 (N_7841,N_7658,N_7561);
and U7842 (N_7842,N_7553,N_7664);
nand U7843 (N_7843,N_7645,N_7506);
nand U7844 (N_7844,N_7586,N_7536);
nand U7845 (N_7845,N_7772,N_7797);
nand U7846 (N_7846,N_7560,N_7544);
nand U7847 (N_7847,N_7671,N_7764);
nand U7848 (N_7848,N_7520,N_7519);
nand U7849 (N_7849,N_7551,N_7774);
xnor U7850 (N_7850,N_7771,N_7784);
or U7851 (N_7851,N_7570,N_7607);
nor U7852 (N_7852,N_7563,N_7644);
nor U7853 (N_7853,N_7526,N_7674);
nand U7854 (N_7854,N_7611,N_7625);
or U7855 (N_7855,N_7798,N_7703);
and U7856 (N_7856,N_7590,N_7704);
xor U7857 (N_7857,N_7609,N_7720);
nor U7858 (N_7858,N_7731,N_7525);
or U7859 (N_7859,N_7588,N_7500);
and U7860 (N_7860,N_7600,N_7736);
nor U7861 (N_7861,N_7652,N_7762);
and U7862 (N_7862,N_7766,N_7673);
or U7863 (N_7863,N_7663,N_7641);
nor U7864 (N_7864,N_7592,N_7518);
nand U7865 (N_7865,N_7594,N_7697);
or U7866 (N_7866,N_7782,N_7554);
xnor U7867 (N_7867,N_7534,N_7744);
xnor U7868 (N_7868,N_7562,N_7653);
xnor U7869 (N_7869,N_7692,N_7760);
and U7870 (N_7870,N_7546,N_7557);
xnor U7871 (N_7871,N_7531,N_7712);
nand U7872 (N_7872,N_7597,N_7657);
nand U7873 (N_7873,N_7761,N_7514);
and U7874 (N_7874,N_7676,N_7511);
xnor U7875 (N_7875,N_7791,N_7572);
nor U7876 (N_7876,N_7700,N_7575);
nor U7877 (N_7877,N_7693,N_7638);
or U7878 (N_7878,N_7608,N_7620);
nor U7879 (N_7879,N_7631,N_7660);
xor U7880 (N_7880,N_7708,N_7651);
or U7881 (N_7881,N_7538,N_7517);
nor U7882 (N_7882,N_7626,N_7685);
nand U7883 (N_7883,N_7547,N_7555);
nand U7884 (N_7884,N_7787,N_7636);
xor U7885 (N_7885,N_7659,N_7564);
nor U7886 (N_7886,N_7583,N_7706);
nand U7887 (N_7887,N_7707,N_7543);
nor U7888 (N_7888,N_7742,N_7694);
xor U7889 (N_7889,N_7776,N_7755);
nor U7890 (N_7890,N_7516,N_7710);
xnor U7891 (N_7891,N_7748,N_7587);
xor U7892 (N_7892,N_7786,N_7524);
nand U7893 (N_7893,N_7763,N_7770);
nand U7894 (N_7894,N_7759,N_7585);
nor U7895 (N_7895,N_7617,N_7691);
and U7896 (N_7896,N_7621,N_7698);
and U7897 (N_7897,N_7522,N_7643);
xor U7898 (N_7898,N_7649,N_7648);
nand U7899 (N_7899,N_7545,N_7675);
xnor U7900 (N_7900,N_7662,N_7745);
xor U7901 (N_7901,N_7502,N_7767);
xor U7902 (N_7902,N_7541,N_7647);
nor U7903 (N_7903,N_7702,N_7729);
xor U7904 (N_7904,N_7713,N_7559);
nand U7905 (N_7905,N_7548,N_7504);
xor U7906 (N_7906,N_7639,N_7688);
xnor U7907 (N_7907,N_7629,N_7624);
nand U7908 (N_7908,N_7630,N_7646);
xnor U7909 (N_7909,N_7753,N_7567);
and U7910 (N_7910,N_7619,N_7532);
nand U7911 (N_7911,N_7773,N_7616);
nand U7912 (N_7912,N_7790,N_7552);
or U7913 (N_7913,N_7537,N_7735);
nand U7914 (N_7914,N_7679,N_7678);
nor U7915 (N_7915,N_7754,N_7756);
nand U7916 (N_7916,N_7668,N_7582);
xnor U7917 (N_7917,N_7788,N_7579);
nor U7918 (N_7918,N_7612,N_7669);
nor U7919 (N_7919,N_7605,N_7705);
or U7920 (N_7920,N_7530,N_7613);
nor U7921 (N_7921,N_7521,N_7580);
nand U7922 (N_7922,N_7777,N_7535);
xnor U7923 (N_7923,N_7508,N_7683);
nand U7924 (N_7924,N_7689,N_7661);
xor U7925 (N_7925,N_7714,N_7741);
xor U7926 (N_7926,N_7765,N_7721);
and U7927 (N_7927,N_7789,N_7665);
nor U7928 (N_7928,N_7682,N_7785);
and U7929 (N_7929,N_7604,N_7738);
xnor U7930 (N_7930,N_7775,N_7690);
xor U7931 (N_7931,N_7623,N_7746);
xor U7932 (N_7932,N_7529,N_7687);
nor U7933 (N_7933,N_7627,N_7568);
or U7934 (N_7934,N_7650,N_7796);
nand U7935 (N_7935,N_7615,N_7569);
nand U7936 (N_7936,N_7726,N_7523);
nand U7937 (N_7937,N_7571,N_7633);
nand U7938 (N_7938,N_7699,N_7792);
nor U7939 (N_7939,N_7758,N_7681);
nor U7940 (N_7940,N_7794,N_7622);
xor U7941 (N_7941,N_7701,N_7576);
nand U7942 (N_7942,N_7743,N_7591);
or U7943 (N_7943,N_7734,N_7709);
nor U7944 (N_7944,N_7642,N_7501);
nor U7945 (N_7945,N_7595,N_7779);
xor U7946 (N_7946,N_7722,N_7598);
or U7947 (N_7947,N_7603,N_7680);
nor U7948 (N_7948,N_7716,N_7727);
and U7949 (N_7949,N_7717,N_7528);
xor U7950 (N_7950,N_7536,N_7565);
and U7951 (N_7951,N_7550,N_7743);
and U7952 (N_7952,N_7524,N_7676);
nand U7953 (N_7953,N_7682,N_7695);
or U7954 (N_7954,N_7779,N_7735);
nand U7955 (N_7955,N_7503,N_7643);
or U7956 (N_7956,N_7752,N_7700);
nor U7957 (N_7957,N_7795,N_7629);
and U7958 (N_7958,N_7719,N_7727);
xor U7959 (N_7959,N_7552,N_7558);
and U7960 (N_7960,N_7691,N_7793);
nor U7961 (N_7961,N_7561,N_7670);
and U7962 (N_7962,N_7633,N_7759);
xor U7963 (N_7963,N_7634,N_7547);
and U7964 (N_7964,N_7522,N_7591);
and U7965 (N_7965,N_7665,N_7746);
nor U7966 (N_7966,N_7526,N_7791);
and U7967 (N_7967,N_7699,N_7784);
or U7968 (N_7968,N_7693,N_7590);
nor U7969 (N_7969,N_7596,N_7657);
and U7970 (N_7970,N_7517,N_7646);
xor U7971 (N_7971,N_7733,N_7588);
or U7972 (N_7972,N_7536,N_7587);
and U7973 (N_7973,N_7610,N_7690);
xor U7974 (N_7974,N_7723,N_7797);
or U7975 (N_7975,N_7708,N_7777);
or U7976 (N_7976,N_7606,N_7720);
and U7977 (N_7977,N_7575,N_7669);
nor U7978 (N_7978,N_7526,N_7609);
nand U7979 (N_7979,N_7714,N_7636);
or U7980 (N_7980,N_7566,N_7752);
or U7981 (N_7981,N_7517,N_7583);
nand U7982 (N_7982,N_7694,N_7553);
and U7983 (N_7983,N_7750,N_7709);
nand U7984 (N_7984,N_7797,N_7546);
nand U7985 (N_7985,N_7559,N_7782);
nand U7986 (N_7986,N_7679,N_7719);
xor U7987 (N_7987,N_7795,N_7533);
or U7988 (N_7988,N_7646,N_7713);
or U7989 (N_7989,N_7760,N_7554);
and U7990 (N_7990,N_7636,N_7624);
or U7991 (N_7991,N_7777,N_7528);
nand U7992 (N_7992,N_7526,N_7523);
nand U7993 (N_7993,N_7666,N_7695);
and U7994 (N_7994,N_7517,N_7544);
and U7995 (N_7995,N_7766,N_7718);
xnor U7996 (N_7996,N_7569,N_7737);
and U7997 (N_7997,N_7519,N_7625);
xnor U7998 (N_7998,N_7647,N_7538);
or U7999 (N_7999,N_7502,N_7611);
or U8000 (N_8000,N_7551,N_7638);
nand U8001 (N_8001,N_7775,N_7599);
nand U8002 (N_8002,N_7765,N_7502);
or U8003 (N_8003,N_7526,N_7576);
or U8004 (N_8004,N_7618,N_7763);
or U8005 (N_8005,N_7531,N_7515);
and U8006 (N_8006,N_7742,N_7698);
or U8007 (N_8007,N_7621,N_7673);
nand U8008 (N_8008,N_7617,N_7544);
nand U8009 (N_8009,N_7731,N_7645);
nand U8010 (N_8010,N_7757,N_7736);
or U8011 (N_8011,N_7624,N_7674);
nor U8012 (N_8012,N_7652,N_7534);
or U8013 (N_8013,N_7603,N_7650);
nor U8014 (N_8014,N_7501,N_7781);
nand U8015 (N_8015,N_7639,N_7527);
xor U8016 (N_8016,N_7648,N_7724);
nor U8017 (N_8017,N_7528,N_7748);
nor U8018 (N_8018,N_7748,N_7699);
nor U8019 (N_8019,N_7584,N_7644);
or U8020 (N_8020,N_7699,N_7752);
or U8021 (N_8021,N_7771,N_7751);
nand U8022 (N_8022,N_7744,N_7777);
or U8023 (N_8023,N_7748,N_7736);
and U8024 (N_8024,N_7653,N_7599);
xnor U8025 (N_8025,N_7701,N_7654);
xnor U8026 (N_8026,N_7791,N_7646);
or U8027 (N_8027,N_7711,N_7610);
or U8028 (N_8028,N_7648,N_7646);
xnor U8029 (N_8029,N_7540,N_7676);
and U8030 (N_8030,N_7771,N_7787);
nor U8031 (N_8031,N_7731,N_7725);
or U8032 (N_8032,N_7519,N_7670);
nand U8033 (N_8033,N_7522,N_7564);
or U8034 (N_8034,N_7501,N_7606);
nand U8035 (N_8035,N_7734,N_7723);
xor U8036 (N_8036,N_7583,N_7607);
nor U8037 (N_8037,N_7523,N_7569);
nor U8038 (N_8038,N_7566,N_7715);
xor U8039 (N_8039,N_7501,N_7785);
nand U8040 (N_8040,N_7626,N_7742);
xor U8041 (N_8041,N_7566,N_7697);
nor U8042 (N_8042,N_7717,N_7650);
nor U8043 (N_8043,N_7737,N_7632);
xnor U8044 (N_8044,N_7641,N_7509);
nand U8045 (N_8045,N_7677,N_7512);
xnor U8046 (N_8046,N_7619,N_7520);
nand U8047 (N_8047,N_7694,N_7788);
nor U8048 (N_8048,N_7592,N_7677);
and U8049 (N_8049,N_7514,N_7791);
nor U8050 (N_8050,N_7678,N_7632);
nor U8051 (N_8051,N_7540,N_7670);
nor U8052 (N_8052,N_7777,N_7680);
nand U8053 (N_8053,N_7745,N_7695);
xnor U8054 (N_8054,N_7766,N_7753);
nand U8055 (N_8055,N_7525,N_7619);
xor U8056 (N_8056,N_7726,N_7709);
nand U8057 (N_8057,N_7687,N_7503);
nand U8058 (N_8058,N_7546,N_7653);
or U8059 (N_8059,N_7677,N_7598);
xnor U8060 (N_8060,N_7698,N_7514);
nor U8061 (N_8061,N_7504,N_7542);
or U8062 (N_8062,N_7764,N_7620);
nor U8063 (N_8063,N_7563,N_7704);
or U8064 (N_8064,N_7783,N_7714);
or U8065 (N_8065,N_7639,N_7570);
or U8066 (N_8066,N_7763,N_7594);
or U8067 (N_8067,N_7722,N_7736);
nor U8068 (N_8068,N_7737,N_7552);
nor U8069 (N_8069,N_7518,N_7724);
nand U8070 (N_8070,N_7543,N_7640);
or U8071 (N_8071,N_7794,N_7599);
xor U8072 (N_8072,N_7799,N_7690);
xor U8073 (N_8073,N_7638,N_7624);
or U8074 (N_8074,N_7709,N_7509);
or U8075 (N_8075,N_7556,N_7522);
or U8076 (N_8076,N_7696,N_7626);
xor U8077 (N_8077,N_7580,N_7555);
nor U8078 (N_8078,N_7780,N_7645);
nand U8079 (N_8079,N_7760,N_7574);
or U8080 (N_8080,N_7614,N_7704);
nor U8081 (N_8081,N_7507,N_7798);
nand U8082 (N_8082,N_7571,N_7735);
or U8083 (N_8083,N_7745,N_7565);
xor U8084 (N_8084,N_7685,N_7699);
and U8085 (N_8085,N_7722,N_7651);
nor U8086 (N_8086,N_7663,N_7527);
nor U8087 (N_8087,N_7602,N_7541);
xor U8088 (N_8088,N_7782,N_7726);
or U8089 (N_8089,N_7692,N_7504);
nand U8090 (N_8090,N_7507,N_7762);
xnor U8091 (N_8091,N_7686,N_7650);
xor U8092 (N_8092,N_7656,N_7780);
and U8093 (N_8093,N_7722,N_7765);
nand U8094 (N_8094,N_7628,N_7502);
and U8095 (N_8095,N_7505,N_7553);
and U8096 (N_8096,N_7634,N_7760);
xnor U8097 (N_8097,N_7658,N_7710);
xor U8098 (N_8098,N_7661,N_7585);
or U8099 (N_8099,N_7566,N_7713);
nor U8100 (N_8100,N_8098,N_8052);
or U8101 (N_8101,N_7802,N_8065);
nand U8102 (N_8102,N_7805,N_7957);
and U8103 (N_8103,N_8009,N_8030);
nor U8104 (N_8104,N_8056,N_8037);
xnor U8105 (N_8105,N_8034,N_8024);
and U8106 (N_8106,N_7974,N_7954);
nor U8107 (N_8107,N_8092,N_7949);
and U8108 (N_8108,N_8075,N_7851);
xnor U8109 (N_8109,N_7867,N_7860);
xnor U8110 (N_8110,N_7989,N_7864);
nand U8111 (N_8111,N_7882,N_7898);
nor U8112 (N_8112,N_8015,N_7857);
nand U8113 (N_8113,N_8051,N_7913);
nand U8114 (N_8114,N_8078,N_8069);
nand U8115 (N_8115,N_7810,N_8012);
nand U8116 (N_8116,N_8044,N_7958);
or U8117 (N_8117,N_7887,N_8083);
nor U8118 (N_8118,N_8026,N_8002);
and U8119 (N_8119,N_7827,N_7907);
or U8120 (N_8120,N_7987,N_8001);
nor U8121 (N_8121,N_7980,N_7978);
nand U8122 (N_8122,N_7896,N_8022);
nand U8123 (N_8123,N_7930,N_8021);
or U8124 (N_8124,N_7839,N_8080);
nor U8125 (N_8125,N_8074,N_7821);
or U8126 (N_8126,N_8084,N_7814);
or U8127 (N_8127,N_8059,N_7817);
nor U8128 (N_8128,N_8076,N_7942);
nand U8129 (N_8129,N_7933,N_7904);
nor U8130 (N_8130,N_8003,N_8082);
and U8131 (N_8131,N_8046,N_7916);
xnor U8132 (N_8132,N_7825,N_8063);
and U8133 (N_8133,N_7990,N_7973);
xor U8134 (N_8134,N_7955,N_7950);
or U8135 (N_8135,N_7931,N_7878);
xor U8136 (N_8136,N_8060,N_7861);
nand U8137 (N_8137,N_7844,N_7870);
nand U8138 (N_8138,N_7897,N_8087);
nor U8139 (N_8139,N_7981,N_7905);
nor U8140 (N_8140,N_7800,N_7853);
xnor U8141 (N_8141,N_7831,N_7856);
and U8142 (N_8142,N_8048,N_7935);
or U8143 (N_8143,N_7823,N_8004);
nand U8144 (N_8144,N_7952,N_7809);
nand U8145 (N_8145,N_7979,N_8047);
xor U8146 (N_8146,N_7837,N_7964);
xor U8147 (N_8147,N_7876,N_8073);
xor U8148 (N_8148,N_7858,N_7946);
and U8149 (N_8149,N_8099,N_8019);
xor U8150 (N_8150,N_7811,N_7885);
or U8151 (N_8151,N_8042,N_8011);
xor U8152 (N_8152,N_7908,N_7845);
nand U8153 (N_8153,N_7822,N_7919);
xnor U8154 (N_8154,N_8064,N_7863);
nor U8155 (N_8155,N_7871,N_8041);
or U8156 (N_8156,N_8007,N_7911);
nor U8157 (N_8157,N_7828,N_8097);
xnor U8158 (N_8158,N_7881,N_7884);
and U8159 (N_8159,N_7842,N_7994);
xor U8160 (N_8160,N_7912,N_7850);
nor U8161 (N_8161,N_8079,N_7862);
or U8162 (N_8162,N_7848,N_7932);
or U8163 (N_8163,N_7944,N_7874);
or U8164 (N_8164,N_7890,N_7961);
xor U8165 (N_8165,N_7895,N_8045);
or U8166 (N_8166,N_7824,N_7976);
nor U8167 (N_8167,N_7986,N_8013);
or U8168 (N_8168,N_7900,N_8008);
nor U8169 (N_8169,N_7807,N_7927);
xnor U8170 (N_8170,N_7923,N_7920);
nor U8171 (N_8171,N_7840,N_7801);
nor U8172 (N_8172,N_7906,N_7886);
xor U8173 (N_8173,N_7967,N_8043);
or U8174 (N_8174,N_8058,N_8033);
nor U8175 (N_8175,N_7838,N_7929);
or U8176 (N_8176,N_8014,N_8057);
and U8177 (N_8177,N_7934,N_7830);
or U8178 (N_8178,N_8072,N_7938);
nor U8179 (N_8179,N_8023,N_7962);
xor U8180 (N_8180,N_7915,N_7988);
nand U8181 (N_8181,N_7977,N_8054);
or U8182 (N_8182,N_8027,N_7922);
or U8183 (N_8183,N_8017,N_7866);
xor U8184 (N_8184,N_7993,N_7970);
and U8185 (N_8185,N_7879,N_7960);
nand U8186 (N_8186,N_7982,N_7940);
xor U8187 (N_8187,N_7836,N_7849);
nand U8188 (N_8188,N_8067,N_7996);
xor U8189 (N_8189,N_7984,N_7893);
xnor U8190 (N_8190,N_7924,N_8091);
and U8191 (N_8191,N_7926,N_7951);
nand U8192 (N_8192,N_7818,N_7936);
nand U8193 (N_8193,N_7855,N_7843);
or U8194 (N_8194,N_7941,N_7937);
and U8195 (N_8195,N_7903,N_7899);
xor U8196 (N_8196,N_7877,N_7852);
and U8197 (N_8197,N_8062,N_7925);
nor U8198 (N_8198,N_7854,N_7847);
nor U8199 (N_8199,N_7889,N_7815);
and U8200 (N_8200,N_8029,N_7972);
nand U8201 (N_8201,N_8032,N_8089);
and U8202 (N_8202,N_8010,N_7910);
and U8203 (N_8203,N_7969,N_8061);
nand U8204 (N_8204,N_7846,N_7868);
nor U8205 (N_8205,N_7869,N_8071);
or U8206 (N_8206,N_7959,N_7918);
nand U8207 (N_8207,N_8090,N_7914);
nand U8208 (N_8208,N_7921,N_7939);
or U8209 (N_8209,N_8000,N_8068);
nor U8210 (N_8210,N_8088,N_8086);
or U8211 (N_8211,N_7833,N_7894);
or U8212 (N_8212,N_8005,N_7991);
xor U8213 (N_8213,N_7813,N_7992);
nor U8214 (N_8214,N_7891,N_8035);
nor U8215 (N_8215,N_7812,N_8016);
or U8216 (N_8216,N_7947,N_7875);
or U8217 (N_8217,N_7971,N_7859);
nand U8218 (N_8218,N_8053,N_8006);
and U8219 (N_8219,N_7909,N_7928);
and U8220 (N_8220,N_8096,N_7995);
nand U8221 (N_8221,N_7945,N_7985);
xnor U8222 (N_8222,N_7804,N_8020);
and U8223 (N_8223,N_7826,N_8040);
nor U8224 (N_8224,N_8025,N_7819);
xor U8225 (N_8225,N_7808,N_7963);
nor U8226 (N_8226,N_8077,N_8028);
xor U8227 (N_8227,N_7948,N_8066);
or U8228 (N_8228,N_7873,N_7966);
or U8229 (N_8229,N_7999,N_7956);
and U8230 (N_8230,N_7841,N_8018);
nand U8231 (N_8231,N_8070,N_7902);
or U8232 (N_8232,N_7872,N_8093);
xnor U8233 (N_8233,N_7888,N_8039);
nor U8234 (N_8234,N_8050,N_7997);
nand U8235 (N_8235,N_7835,N_7829);
nand U8236 (N_8236,N_7816,N_7865);
and U8237 (N_8237,N_7943,N_8081);
nor U8238 (N_8238,N_7820,N_7953);
nand U8239 (N_8239,N_8036,N_8095);
nor U8240 (N_8240,N_8085,N_7968);
or U8241 (N_8241,N_8038,N_7901);
nand U8242 (N_8242,N_7832,N_7892);
and U8243 (N_8243,N_8055,N_8049);
xor U8244 (N_8244,N_8094,N_7803);
and U8245 (N_8245,N_7834,N_7965);
or U8246 (N_8246,N_7983,N_8031);
nand U8247 (N_8247,N_7998,N_7880);
nor U8248 (N_8248,N_7883,N_7917);
nor U8249 (N_8249,N_7806,N_7975);
and U8250 (N_8250,N_8020,N_7929);
nand U8251 (N_8251,N_7982,N_7823);
or U8252 (N_8252,N_7976,N_7942);
xnor U8253 (N_8253,N_7988,N_7820);
nand U8254 (N_8254,N_7810,N_8087);
and U8255 (N_8255,N_7932,N_8054);
or U8256 (N_8256,N_7803,N_8034);
nand U8257 (N_8257,N_7962,N_7979);
and U8258 (N_8258,N_8090,N_7915);
and U8259 (N_8259,N_7852,N_7907);
or U8260 (N_8260,N_8059,N_8076);
or U8261 (N_8261,N_8062,N_8008);
and U8262 (N_8262,N_7810,N_7853);
nand U8263 (N_8263,N_7838,N_7909);
and U8264 (N_8264,N_7812,N_7969);
or U8265 (N_8265,N_8046,N_8018);
or U8266 (N_8266,N_8028,N_7828);
xnor U8267 (N_8267,N_8048,N_8008);
and U8268 (N_8268,N_7806,N_7899);
or U8269 (N_8269,N_8086,N_7870);
nor U8270 (N_8270,N_7824,N_7914);
or U8271 (N_8271,N_7889,N_8007);
nor U8272 (N_8272,N_7810,N_8039);
xor U8273 (N_8273,N_7861,N_7857);
or U8274 (N_8274,N_7985,N_7977);
or U8275 (N_8275,N_8089,N_7980);
nand U8276 (N_8276,N_7840,N_7866);
or U8277 (N_8277,N_8003,N_7870);
xnor U8278 (N_8278,N_8067,N_8038);
or U8279 (N_8279,N_7800,N_7996);
and U8280 (N_8280,N_8037,N_7858);
and U8281 (N_8281,N_7886,N_7900);
xnor U8282 (N_8282,N_7890,N_8096);
nor U8283 (N_8283,N_7877,N_7867);
and U8284 (N_8284,N_8026,N_7967);
nand U8285 (N_8285,N_7898,N_7857);
nor U8286 (N_8286,N_7827,N_8091);
and U8287 (N_8287,N_7907,N_7916);
or U8288 (N_8288,N_7956,N_8069);
nor U8289 (N_8289,N_7818,N_7872);
nand U8290 (N_8290,N_7890,N_8031);
and U8291 (N_8291,N_7839,N_7832);
or U8292 (N_8292,N_7987,N_7964);
and U8293 (N_8293,N_7833,N_7928);
xnor U8294 (N_8294,N_7998,N_7861);
and U8295 (N_8295,N_8068,N_7875);
or U8296 (N_8296,N_8004,N_8023);
nor U8297 (N_8297,N_8060,N_7819);
nand U8298 (N_8298,N_7999,N_8079);
nand U8299 (N_8299,N_7956,N_7899);
nand U8300 (N_8300,N_7968,N_7925);
or U8301 (N_8301,N_8099,N_8031);
or U8302 (N_8302,N_8072,N_8023);
or U8303 (N_8303,N_8085,N_7922);
xor U8304 (N_8304,N_7870,N_7953);
or U8305 (N_8305,N_7985,N_8051);
nor U8306 (N_8306,N_8074,N_7909);
nor U8307 (N_8307,N_7921,N_7815);
xor U8308 (N_8308,N_7981,N_8024);
nor U8309 (N_8309,N_7826,N_8098);
nand U8310 (N_8310,N_7870,N_7912);
or U8311 (N_8311,N_8071,N_8034);
nand U8312 (N_8312,N_7827,N_7891);
xnor U8313 (N_8313,N_7925,N_7854);
and U8314 (N_8314,N_7949,N_7854);
nor U8315 (N_8315,N_7947,N_8028);
or U8316 (N_8316,N_8094,N_7863);
nor U8317 (N_8317,N_7832,N_8014);
xor U8318 (N_8318,N_7940,N_8028);
nand U8319 (N_8319,N_7981,N_8081);
and U8320 (N_8320,N_7893,N_8001);
and U8321 (N_8321,N_7847,N_7942);
and U8322 (N_8322,N_7801,N_7911);
or U8323 (N_8323,N_7892,N_7971);
nand U8324 (N_8324,N_7849,N_8077);
or U8325 (N_8325,N_7851,N_7874);
xnor U8326 (N_8326,N_7981,N_8017);
or U8327 (N_8327,N_7840,N_8044);
nand U8328 (N_8328,N_7988,N_7985);
nor U8329 (N_8329,N_7977,N_8065);
or U8330 (N_8330,N_7907,N_8073);
nor U8331 (N_8331,N_7962,N_8022);
nand U8332 (N_8332,N_7921,N_7996);
nand U8333 (N_8333,N_8017,N_7853);
nand U8334 (N_8334,N_7852,N_7867);
nor U8335 (N_8335,N_8045,N_7890);
and U8336 (N_8336,N_8004,N_7921);
nor U8337 (N_8337,N_8037,N_7930);
and U8338 (N_8338,N_8040,N_7850);
nand U8339 (N_8339,N_7948,N_8071);
nand U8340 (N_8340,N_7891,N_7841);
and U8341 (N_8341,N_7894,N_7958);
nand U8342 (N_8342,N_8081,N_7857);
xnor U8343 (N_8343,N_7916,N_8007);
or U8344 (N_8344,N_7994,N_8065);
nand U8345 (N_8345,N_8010,N_7959);
and U8346 (N_8346,N_7994,N_7908);
and U8347 (N_8347,N_7956,N_7803);
nand U8348 (N_8348,N_7803,N_7847);
or U8349 (N_8349,N_8091,N_7840);
or U8350 (N_8350,N_7807,N_8076);
xor U8351 (N_8351,N_7835,N_8069);
or U8352 (N_8352,N_7830,N_8040);
nand U8353 (N_8353,N_8096,N_7914);
or U8354 (N_8354,N_7957,N_8079);
nor U8355 (N_8355,N_8059,N_7927);
or U8356 (N_8356,N_8003,N_7940);
or U8357 (N_8357,N_8007,N_8072);
or U8358 (N_8358,N_7998,N_7941);
xor U8359 (N_8359,N_7993,N_8044);
and U8360 (N_8360,N_7852,N_7952);
nand U8361 (N_8361,N_7957,N_7858);
nand U8362 (N_8362,N_7989,N_7870);
xor U8363 (N_8363,N_7835,N_7818);
nor U8364 (N_8364,N_8085,N_8080);
nor U8365 (N_8365,N_7999,N_7811);
and U8366 (N_8366,N_8007,N_7885);
and U8367 (N_8367,N_8037,N_7801);
nor U8368 (N_8368,N_7986,N_7969);
nand U8369 (N_8369,N_8079,N_7970);
or U8370 (N_8370,N_7969,N_7989);
and U8371 (N_8371,N_8063,N_7994);
nand U8372 (N_8372,N_8074,N_8049);
and U8373 (N_8373,N_7842,N_8031);
or U8374 (N_8374,N_7970,N_7925);
xnor U8375 (N_8375,N_7842,N_8052);
nor U8376 (N_8376,N_7980,N_7839);
nand U8377 (N_8377,N_8061,N_8041);
and U8378 (N_8378,N_7833,N_8064);
nand U8379 (N_8379,N_8065,N_7913);
nand U8380 (N_8380,N_7875,N_8064);
or U8381 (N_8381,N_8048,N_7877);
and U8382 (N_8382,N_7848,N_7864);
and U8383 (N_8383,N_7891,N_7897);
or U8384 (N_8384,N_8079,N_7916);
xnor U8385 (N_8385,N_7817,N_8025);
or U8386 (N_8386,N_7867,N_8017);
and U8387 (N_8387,N_8055,N_8047);
nor U8388 (N_8388,N_7994,N_7800);
and U8389 (N_8389,N_7876,N_7920);
nand U8390 (N_8390,N_8094,N_7814);
nand U8391 (N_8391,N_7929,N_7950);
and U8392 (N_8392,N_7872,N_7906);
nand U8393 (N_8393,N_7965,N_7942);
xor U8394 (N_8394,N_7986,N_7946);
and U8395 (N_8395,N_7959,N_8008);
nor U8396 (N_8396,N_7956,N_8001);
or U8397 (N_8397,N_7880,N_7923);
nand U8398 (N_8398,N_8019,N_8053);
xor U8399 (N_8399,N_8046,N_7935);
xnor U8400 (N_8400,N_8397,N_8396);
nor U8401 (N_8401,N_8235,N_8221);
xnor U8402 (N_8402,N_8259,N_8108);
or U8403 (N_8403,N_8105,N_8191);
nor U8404 (N_8404,N_8146,N_8262);
xor U8405 (N_8405,N_8314,N_8303);
xor U8406 (N_8406,N_8237,N_8238);
and U8407 (N_8407,N_8112,N_8106);
nand U8408 (N_8408,N_8297,N_8305);
nand U8409 (N_8409,N_8242,N_8157);
or U8410 (N_8410,N_8289,N_8358);
nor U8411 (N_8411,N_8366,N_8180);
xnor U8412 (N_8412,N_8300,N_8275);
and U8413 (N_8413,N_8168,N_8308);
or U8414 (N_8414,N_8370,N_8362);
or U8415 (N_8415,N_8261,N_8376);
xnor U8416 (N_8416,N_8270,N_8188);
xnor U8417 (N_8417,N_8179,N_8109);
xor U8418 (N_8418,N_8239,N_8317);
xnor U8419 (N_8419,N_8390,N_8318);
xor U8420 (N_8420,N_8244,N_8380);
nor U8421 (N_8421,N_8125,N_8187);
nor U8422 (N_8422,N_8155,N_8296);
xor U8423 (N_8423,N_8383,N_8124);
xor U8424 (N_8424,N_8138,N_8233);
xor U8425 (N_8425,N_8208,N_8101);
or U8426 (N_8426,N_8194,N_8243);
nand U8427 (N_8427,N_8339,N_8373);
nor U8428 (N_8428,N_8241,N_8174);
xnor U8429 (N_8429,N_8272,N_8218);
nor U8430 (N_8430,N_8288,N_8126);
nand U8431 (N_8431,N_8120,N_8361);
and U8432 (N_8432,N_8398,N_8207);
nor U8433 (N_8433,N_8253,N_8193);
nand U8434 (N_8434,N_8331,N_8260);
or U8435 (N_8435,N_8395,N_8177);
or U8436 (N_8436,N_8224,N_8163);
or U8437 (N_8437,N_8330,N_8249);
nor U8438 (N_8438,N_8195,N_8309);
or U8439 (N_8439,N_8389,N_8319);
nor U8440 (N_8440,N_8315,N_8378);
xnor U8441 (N_8441,N_8332,N_8154);
or U8442 (N_8442,N_8178,N_8279);
and U8443 (N_8443,N_8290,N_8327);
or U8444 (N_8444,N_8387,N_8394);
and U8445 (N_8445,N_8113,N_8100);
nand U8446 (N_8446,N_8299,N_8333);
and U8447 (N_8447,N_8206,N_8159);
nor U8448 (N_8448,N_8137,N_8271);
nand U8449 (N_8449,N_8228,N_8165);
or U8450 (N_8450,N_8329,N_8252);
and U8451 (N_8451,N_8216,N_8255);
nand U8452 (N_8452,N_8250,N_8189);
xnor U8453 (N_8453,N_8246,N_8220);
nand U8454 (N_8454,N_8121,N_8236);
nand U8455 (N_8455,N_8198,N_8148);
or U8456 (N_8456,N_8222,N_8134);
nor U8457 (N_8457,N_8298,N_8136);
nor U8458 (N_8458,N_8215,N_8353);
xnor U8459 (N_8459,N_8133,N_8164);
or U8460 (N_8460,N_8377,N_8116);
or U8461 (N_8461,N_8213,N_8285);
nor U8462 (N_8462,N_8230,N_8254);
or U8463 (N_8463,N_8141,N_8161);
and U8464 (N_8464,N_8368,N_8247);
nor U8465 (N_8465,N_8104,N_8231);
nand U8466 (N_8466,N_8167,N_8278);
and U8467 (N_8467,N_8132,N_8349);
and U8468 (N_8468,N_8382,N_8140);
nor U8469 (N_8469,N_8123,N_8291);
or U8470 (N_8470,N_8355,N_8186);
nor U8471 (N_8471,N_8367,N_8313);
and U8472 (N_8472,N_8344,N_8284);
and U8473 (N_8473,N_8345,N_8268);
and U8474 (N_8474,N_8128,N_8149);
or U8475 (N_8475,N_8334,N_8201);
nand U8476 (N_8476,N_8365,N_8371);
xnor U8477 (N_8477,N_8185,N_8184);
xor U8478 (N_8478,N_8173,N_8384);
and U8479 (N_8479,N_8286,N_8274);
or U8480 (N_8480,N_8343,N_8266);
xnor U8481 (N_8481,N_8203,N_8114);
and U8482 (N_8482,N_8248,N_8356);
xnor U8483 (N_8483,N_8301,N_8338);
nor U8484 (N_8484,N_8111,N_8147);
and U8485 (N_8485,N_8166,N_8359);
nor U8486 (N_8486,N_8322,N_8229);
xnor U8487 (N_8487,N_8219,N_8304);
xor U8488 (N_8488,N_8281,N_8381);
and U8489 (N_8489,N_8341,N_8392);
nor U8490 (N_8490,N_8399,N_8360);
and U8491 (N_8491,N_8307,N_8131);
nand U8492 (N_8492,N_8379,N_8294);
or U8493 (N_8493,N_8139,N_8265);
nand U8494 (N_8494,N_8200,N_8282);
nand U8495 (N_8495,N_8202,N_8335);
and U8496 (N_8496,N_8267,N_8357);
or U8497 (N_8497,N_8227,N_8388);
xor U8498 (N_8498,N_8115,N_8119);
or U8499 (N_8499,N_8256,N_8199);
nand U8500 (N_8500,N_8372,N_8245);
and U8501 (N_8501,N_8293,N_8354);
or U8502 (N_8502,N_8336,N_8144);
xor U8503 (N_8503,N_8226,N_8302);
or U8504 (N_8504,N_8352,N_8183);
xnor U8505 (N_8505,N_8350,N_8171);
and U8506 (N_8506,N_8196,N_8156);
xnor U8507 (N_8507,N_8232,N_8192);
nand U8508 (N_8508,N_8351,N_8325);
and U8509 (N_8509,N_8385,N_8127);
nor U8510 (N_8510,N_8292,N_8150);
xnor U8511 (N_8511,N_8169,N_8240);
nand U8512 (N_8512,N_8295,N_8181);
or U8513 (N_8513,N_8182,N_8283);
or U8514 (N_8514,N_8211,N_8103);
xnor U8515 (N_8515,N_8264,N_8153);
nand U8516 (N_8516,N_8212,N_8209);
nand U8517 (N_8517,N_8323,N_8151);
and U8518 (N_8518,N_8160,N_8258);
nor U8519 (N_8519,N_8102,N_8287);
and U8520 (N_8520,N_8210,N_8328);
and U8521 (N_8521,N_8145,N_8234);
or U8522 (N_8522,N_8342,N_8277);
and U8523 (N_8523,N_8374,N_8152);
or U8524 (N_8524,N_8310,N_8269);
nor U8525 (N_8525,N_8273,N_8347);
nor U8526 (N_8526,N_8346,N_8257);
and U8527 (N_8527,N_8118,N_8312);
and U8528 (N_8528,N_8321,N_8337);
or U8529 (N_8529,N_8263,N_8214);
or U8530 (N_8530,N_8320,N_8251);
xnor U8531 (N_8531,N_8280,N_8158);
and U8532 (N_8532,N_8324,N_8340);
xnor U8533 (N_8533,N_8162,N_8117);
nor U8534 (N_8534,N_8375,N_8306);
and U8535 (N_8535,N_8223,N_8204);
and U8536 (N_8536,N_8393,N_8316);
nand U8537 (N_8537,N_8143,N_8107);
xnor U8538 (N_8538,N_8190,N_8176);
xnor U8539 (N_8539,N_8129,N_8130);
nand U8540 (N_8540,N_8326,N_8311);
or U8541 (N_8541,N_8170,N_8364);
or U8542 (N_8542,N_8217,N_8225);
or U8543 (N_8543,N_8197,N_8363);
xor U8544 (N_8544,N_8369,N_8386);
nand U8545 (N_8545,N_8142,N_8122);
nor U8546 (N_8546,N_8276,N_8205);
nand U8547 (N_8547,N_8110,N_8135);
nor U8548 (N_8548,N_8175,N_8172);
xnor U8549 (N_8549,N_8348,N_8391);
or U8550 (N_8550,N_8345,N_8167);
or U8551 (N_8551,N_8186,N_8246);
xnor U8552 (N_8552,N_8174,N_8395);
or U8553 (N_8553,N_8106,N_8385);
nand U8554 (N_8554,N_8181,N_8336);
nand U8555 (N_8555,N_8110,N_8333);
or U8556 (N_8556,N_8177,N_8363);
nor U8557 (N_8557,N_8328,N_8291);
and U8558 (N_8558,N_8259,N_8154);
or U8559 (N_8559,N_8160,N_8173);
and U8560 (N_8560,N_8386,N_8163);
and U8561 (N_8561,N_8107,N_8377);
or U8562 (N_8562,N_8397,N_8333);
and U8563 (N_8563,N_8212,N_8327);
nand U8564 (N_8564,N_8138,N_8142);
nand U8565 (N_8565,N_8151,N_8314);
and U8566 (N_8566,N_8346,N_8394);
or U8567 (N_8567,N_8349,N_8345);
and U8568 (N_8568,N_8283,N_8220);
and U8569 (N_8569,N_8213,N_8280);
nor U8570 (N_8570,N_8372,N_8286);
nor U8571 (N_8571,N_8228,N_8332);
or U8572 (N_8572,N_8341,N_8177);
xor U8573 (N_8573,N_8108,N_8121);
nor U8574 (N_8574,N_8342,N_8164);
xor U8575 (N_8575,N_8350,N_8347);
nand U8576 (N_8576,N_8266,N_8198);
xnor U8577 (N_8577,N_8325,N_8157);
or U8578 (N_8578,N_8197,N_8191);
and U8579 (N_8579,N_8132,N_8382);
nor U8580 (N_8580,N_8259,N_8256);
or U8581 (N_8581,N_8267,N_8332);
xnor U8582 (N_8582,N_8211,N_8244);
xnor U8583 (N_8583,N_8389,N_8265);
nor U8584 (N_8584,N_8248,N_8287);
nand U8585 (N_8585,N_8284,N_8195);
nand U8586 (N_8586,N_8152,N_8399);
and U8587 (N_8587,N_8191,N_8163);
xor U8588 (N_8588,N_8238,N_8166);
nand U8589 (N_8589,N_8213,N_8138);
and U8590 (N_8590,N_8395,N_8382);
and U8591 (N_8591,N_8124,N_8367);
and U8592 (N_8592,N_8164,N_8351);
nand U8593 (N_8593,N_8395,N_8217);
nand U8594 (N_8594,N_8130,N_8280);
nor U8595 (N_8595,N_8395,N_8242);
xor U8596 (N_8596,N_8349,N_8318);
nand U8597 (N_8597,N_8113,N_8383);
nor U8598 (N_8598,N_8292,N_8135);
and U8599 (N_8599,N_8133,N_8351);
or U8600 (N_8600,N_8290,N_8266);
or U8601 (N_8601,N_8225,N_8205);
xnor U8602 (N_8602,N_8132,N_8220);
and U8603 (N_8603,N_8292,N_8140);
nand U8604 (N_8604,N_8362,N_8372);
nand U8605 (N_8605,N_8112,N_8383);
or U8606 (N_8606,N_8189,N_8279);
or U8607 (N_8607,N_8392,N_8191);
nand U8608 (N_8608,N_8307,N_8249);
nand U8609 (N_8609,N_8259,N_8354);
nor U8610 (N_8610,N_8119,N_8349);
xor U8611 (N_8611,N_8330,N_8283);
or U8612 (N_8612,N_8297,N_8362);
or U8613 (N_8613,N_8196,N_8301);
and U8614 (N_8614,N_8295,N_8212);
xor U8615 (N_8615,N_8308,N_8103);
or U8616 (N_8616,N_8332,N_8340);
and U8617 (N_8617,N_8311,N_8203);
nor U8618 (N_8618,N_8191,N_8196);
and U8619 (N_8619,N_8266,N_8337);
nor U8620 (N_8620,N_8151,N_8327);
or U8621 (N_8621,N_8168,N_8224);
and U8622 (N_8622,N_8319,N_8263);
nor U8623 (N_8623,N_8251,N_8240);
xnor U8624 (N_8624,N_8221,N_8124);
or U8625 (N_8625,N_8116,N_8175);
nor U8626 (N_8626,N_8142,N_8379);
nor U8627 (N_8627,N_8108,N_8216);
or U8628 (N_8628,N_8369,N_8358);
and U8629 (N_8629,N_8376,N_8241);
nand U8630 (N_8630,N_8366,N_8136);
nand U8631 (N_8631,N_8302,N_8292);
and U8632 (N_8632,N_8276,N_8382);
nor U8633 (N_8633,N_8197,N_8129);
nand U8634 (N_8634,N_8281,N_8183);
nand U8635 (N_8635,N_8229,N_8325);
nor U8636 (N_8636,N_8332,N_8341);
nand U8637 (N_8637,N_8264,N_8287);
or U8638 (N_8638,N_8254,N_8323);
nand U8639 (N_8639,N_8169,N_8335);
or U8640 (N_8640,N_8289,N_8197);
xor U8641 (N_8641,N_8357,N_8378);
xor U8642 (N_8642,N_8128,N_8311);
or U8643 (N_8643,N_8282,N_8109);
xnor U8644 (N_8644,N_8341,N_8135);
nor U8645 (N_8645,N_8360,N_8219);
or U8646 (N_8646,N_8327,N_8147);
and U8647 (N_8647,N_8398,N_8342);
or U8648 (N_8648,N_8116,N_8188);
xnor U8649 (N_8649,N_8159,N_8251);
nor U8650 (N_8650,N_8334,N_8151);
nand U8651 (N_8651,N_8281,N_8332);
nand U8652 (N_8652,N_8262,N_8350);
xnor U8653 (N_8653,N_8158,N_8174);
and U8654 (N_8654,N_8193,N_8372);
xnor U8655 (N_8655,N_8397,N_8123);
and U8656 (N_8656,N_8242,N_8184);
and U8657 (N_8657,N_8189,N_8254);
nor U8658 (N_8658,N_8157,N_8318);
xnor U8659 (N_8659,N_8184,N_8172);
and U8660 (N_8660,N_8136,N_8285);
nand U8661 (N_8661,N_8230,N_8127);
or U8662 (N_8662,N_8133,N_8211);
nor U8663 (N_8663,N_8285,N_8359);
nor U8664 (N_8664,N_8380,N_8324);
xnor U8665 (N_8665,N_8264,N_8143);
nor U8666 (N_8666,N_8334,N_8222);
nand U8667 (N_8667,N_8255,N_8221);
nand U8668 (N_8668,N_8102,N_8198);
and U8669 (N_8669,N_8209,N_8251);
and U8670 (N_8670,N_8323,N_8338);
or U8671 (N_8671,N_8280,N_8121);
nor U8672 (N_8672,N_8175,N_8244);
xnor U8673 (N_8673,N_8175,N_8107);
nor U8674 (N_8674,N_8120,N_8186);
and U8675 (N_8675,N_8173,N_8130);
and U8676 (N_8676,N_8275,N_8377);
nand U8677 (N_8677,N_8212,N_8370);
nor U8678 (N_8678,N_8134,N_8105);
and U8679 (N_8679,N_8395,N_8106);
nor U8680 (N_8680,N_8280,N_8356);
nor U8681 (N_8681,N_8256,N_8147);
nand U8682 (N_8682,N_8312,N_8364);
and U8683 (N_8683,N_8245,N_8203);
nand U8684 (N_8684,N_8303,N_8368);
or U8685 (N_8685,N_8278,N_8179);
or U8686 (N_8686,N_8241,N_8121);
nor U8687 (N_8687,N_8169,N_8160);
xnor U8688 (N_8688,N_8145,N_8261);
xor U8689 (N_8689,N_8382,N_8203);
nor U8690 (N_8690,N_8160,N_8287);
nand U8691 (N_8691,N_8256,N_8146);
nand U8692 (N_8692,N_8139,N_8243);
and U8693 (N_8693,N_8162,N_8235);
or U8694 (N_8694,N_8386,N_8302);
or U8695 (N_8695,N_8207,N_8209);
and U8696 (N_8696,N_8102,N_8372);
nor U8697 (N_8697,N_8150,N_8141);
nor U8698 (N_8698,N_8137,N_8242);
xor U8699 (N_8699,N_8242,N_8213);
nor U8700 (N_8700,N_8636,N_8654);
or U8701 (N_8701,N_8504,N_8443);
xnor U8702 (N_8702,N_8439,N_8540);
xnor U8703 (N_8703,N_8586,N_8678);
xnor U8704 (N_8704,N_8520,N_8482);
nand U8705 (N_8705,N_8627,N_8566);
nor U8706 (N_8706,N_8557,N_8513);
and U8707 (N_8707,N_8537,N_8605);
xnor U8708 (N_8708,N_8653,N_8418);
or U8709 (N_8709,N_8624,N_8503);
or U8710 (N_8710,N_8663,N_8413);
or U8711 (N_8711,N_8519,N_8688);
and U8712 (N_8712,N_8623,N_8660);
or U8713 (N_8713,N_8526,N_8419);
nand U8714 (N_8714,N_8630,N_8544);
nand U8715 (N_8715,N_8489,N_8650);
nor U8716 (N_8716,N_8621,N_8631);
or U8717 (N_8717,N_8649,N_8569);
nor U8718 (N_8718,N_8615,N_8414);
nand U8719 (N_8719,N_8644,N_8656);
nor U8720 (N_8720,N_8416,N_8422);
nor U8721 (N_8721,N_8478,N_8558);
or U8722 (N_8722,N_8436,N_8610);
or U8723 (N_8723,N_8607,N_8588);
nor U8724 (N_8724,N_8480,N_8498);
nand U8725 (N_8725,N_8488,N_8635);
nand U8726 (N_8726,N_8677,N_8541);
or U8727 (N_8727,N_8449,N_8609);
xnor U8728 (N_8728,N_8451,N_8691);
and U8729 (N_8729,N_8538,N_8567);
nor U8730 (N_8730,N_8466,N_8611);
nand U8731 (N_8731,N_8666,N_8604);
xor U8732 (N_8732,N_8458,N_8594);
nand U8733 (N_8733,N_8589,N_8642);
or U8734 (N_8734,N_8561,N_8600);
xor U8735 (N_8735,N_8564,N_8477);
nor U8736 (N_8736,N_8501,N_8428);
xnor U8737 (N_8737,N_8463,N_8554);
nand U8738 (N_8738,N_8673,N_8618);
nand U8739 (N_8739,N_8536,N_8431);
xnor U8740 (N_8740,N_8555,N_8695);
nand U8741 (N_8741,N_8625,N_8619);
nand U8742 (N_8742,N_8486,N_8682);
nand U8743 (N_8743,N_8645,N_8499);
xnor U8744 (N_8744,N_8651,N_8505);
nor U8745 (N_8745,N_8612,N_8590);
and U8746 (N_8746,N_8493,N_8690);
nand U8747 (N_8747,N_8490,N_8514);
xor U8748 (N_8748,N_8510,N_8598);
xor U8749 (N_8749,N_8445,N_8405);
and U8750 (N_8750,N_8565,N_8652);
nand U8751 (N_8751,N_8582,N_8592);
or U8752 (N_8752,N_8496,N_8464);
or U8753 (N_8753,N_8447,N_8452);
nor U8754 (N_8754,N_8689,N_8597);
or U8755 (N_8755,N_8575,N_8495);
and U8756 (N_8756,N_8613,N_8670);
nand U8757 (N_8757,N_8577,N_8626);
xor U8758 (N_8758,N_8430,N_8429);
xor U8759 (N_8759,N_8664,N_8433);
nand U8760 (N_8760,N_8502,N_8442);
nand U8761 (N_8761,N_8438,N_8456);
nor U8762 (N_8762,N_8548,N_8553);
and U8763 (N_8763,N_8531,N_8539);
nand U8764 (N_8764,N_8601,N_8409);
xnor U8765 (N_8765,N_8484,N_8591);
and U8766 (N_8766,N_8687,N_8512);
and U8767 (N_8767,N_8667,N_8684);
or U8768 (N_8768,N_8455,N_8572);
xnor U8769 (N_8769,N_8596,N_8639);
and U8770 (N_8770,N_8622,N_8521);
xnor U8771 (N_8771,N_8475,N_8603);
nor U8772 (N_8772,N_8525,N_8560);
or U8773 (N_8773,N_8693,N_8699);
and U8774 (N_8774,N_8437,N_8574);
nor U8775 (N_8775,N_8628,N_8579);
xor U8776 (N_8776,N_8492,N_8400);
and U8777 (N_8777,N_8402,N_8543);
nand U8778 (N_8778,N_8435,N_8599);
and U8779 (N_8779,N_8646,N_8697);
nand U8780 (N_8780,N_8427,N_8406);
and U8781 (N_8781,N_8424,N_8508);
and U8782 (N_8782,N_8485,N_8529);
xor U8783 (N_8783,N_8655,N_8683);
nor U8784 (N_8784,N_8524,N_8608);
nor U8785 (N_8785,N_8542,N_8616);
and U8786 (N_8786,N_8685,N_8573);
or U8787 (N_8787,N_8665,N_8448);
nor U8788 (N_8788,N_8568,N_8509);
xnor U8789 (N_8789,N_8587,N_8412);
xor U8790 (N_8790,N_8675,N_8638);
nand U8791 (N_8791,N_8415,N_8551);
nand U8792 (N_8792,N_8491,N_8562);
or U8793 (N_8793,N_8634,N_8535);
or U8794 (N_8794,N_8473,N_8632);
nand U8795 (N_8795,N_8563,N_8545);
or U8796 (N_8796,N_8527,N_8669);
nor U8797 (N_8797,N_8500,N_8483);
nand U8798 (N_8798,N_8641,N_8547);
and U8799 (N_8799,N_8578,N_8640);
nor U8800 (N_8800,N_8668,N_8658);
and U8801 (N_8801,N_8516,N_8533);
nor U8802 (N_8802,N_8647,N_8518);
nor U8803 (N_8803,N_8401,N_8471);
nand U8804 (N_8804,N_8470,N_8417);
nand U8805 (N_8805,N_8585,N_8662);
and U8806 (N_8806,N_8549,N_8469);
nor U8807 (N_8807,N_8672,N_8459);
xnor U8808 (N_8808,N_8559,N_8583);
or U8809 (N_8809,N_8637,N_8465);
xnor U8810 (N_8810,N_8528,N_8648);
or U8811 (N_8811,N_8698,N_8457);
and U8812 (N_8812,N_8694,N_8481);
xor U8813 (N_8813,N_8494,N_8440);
or U8814 (N_8814,N_8606,N_8408);
or U8815 (N_8815,N_8454,N_8676);
and U8816 (N_8816,N_8659,N_8432);
xnor U8817 (N_8817,N_8423,N_8580);
and U8818 (N_8818,N_8534,N_8674);
xnor U8819 (N_8819,N_8444,N_8507);
and U8820 (N_8820,N_8461,N_8407);
and U8821 (N_8821,N_8515,N_8680);
or U8822 (N_8822,N_8671,N_8614);
or U8823 (N_8823,N_8556,N_8446);
xor U8824 (N_8824,N_8421,N_8629);
xor U8825 (N_8825,N_8462,N_8523);
nor U8826 (N_8826,N_8686,N_8532);
nor U8827 (N_8827,N_8570,N_8571);
nand U8828 (N_8828,N_8546,N_8595);
or U8829 (N_8829,N_8460,N_8434);
nand U8830 (N_8830,N_8552,N_8426);
xor U8831 (N_8831,N_8581,N_8602);
xnor U8832 (N_8832,N_8550,N_8522);
or U8833 (N_8833,N_8643,N_8633);
nor U8834 (N_8834,N_8661,N_8620);
nand U8835 (N_8835,N_8679,N_8474);
nand U8836 (N_8836,N_8453,N_8410);
xnor U8837 (N_8837,N_8506,N_8487);
nand U8838 (N_8838,N_8530,N_8441);
nor U8839 (N_8839,N_8692,N_8657);
xor U8840 (N_8840,N_8403,N_8467);
and U8841 (N_8841,N_8497,N_8593);
xor U8842 (N_8842,N_8411,N_8476);
and U8843 (N_8843,N_8450,N_8576);
nor U8844 (N_8844,N_8472,N_8517);
or U8845 (N_8845,N_8420,N_8617);
and U8846 (N_8846,N_8511,N_8681);
nor U8847 (N_8847,N_8404,N_8584);
xnor U8848 (N_8848,N_8468,N_8696);
nand U8849 (N_8849,N_8479,N_8425);
nand U8850 (N_8850,N_8626,N_8539);
nor U8851 (N_8851,N_8579,N_8650);
xor U8852 (N_8852,N_8625,N_8400);
nand U8853 (N_8853,N_8672,N_8435);
nand U8854 (N_8854,N_8467,N_8677);
or U8855 (N_8855,N_8549,N_8682);
nand U8856 (N_8856,N_8495,N_8596);
and U8857 (N_8857,N_8691,N_8480);
nor U8858 (N_8858,N_8576,N_8465);
nand U8859 (N_8859,N_8658,N_8609);
and U8860 (N_8860,N_8532,N_8643);
nor U8861 (N_8861,N_8501,N_8678);
nor U8862 (N_8862,N_8466,N_8640);
or U8863 (N_8863,N_8411,N_8554);
xor U8864 (N_8864,N_8423,N_8574);
or U8865 (N_8865,N_8550,N_8670);
nand U8866 (N_8866,N_8585,N_8493);
or U8867 (N_8867,N_8463,N_8409);
xor U8868 (N_8868,N_8555,N_8690);
xnor U8869 (N_8869,N_8511,N_8404);
xnor U8870 (N_8870,N_8527,N_8589);
and U8871 (N_8871,N_8560,N_8405);
and U8872 (N_8872,N_8453,N_8631);
and U8873 (N_8873,N_8614,N_8540);
or U8874 (N_8874,N_8582,N_8414);
nor U8875 (N_8875,N_8689,N_8611);
xor U8876 (N_8876,N_8503,N_8626);
xor U8877 (N_8877,N_8567,N_8666);
nor U8878 (N_8878,N_8615,N_8653);
nand U8879 (N_8879,N_8502,N_8529);
or U8880 (N_8880,N_8557,N_8502);
or U8881 (N_8881,N_8408,N_8599);
and U8882 (N_8882,N_8599,N_8644);
nor U8883 (N_8883,N_8491,N_8548);
xor U8884 (N_8884,N_8414,N_8446);
or U8885 (N_8885,N_8517,N_8551);
or U8886 (N_8886,N_8494,N_8677);
nand U8887 (N_8887,N_8531,N_8508);
nor U8888 (N_8888,N_8665,N_8643);
xor U8889 (N_8889,N_8444,N_8450);
nand U8890 (N_8890,N_8489,N_8557);
or U8891 (N_8891,N_8445,N_8621);
or U8892 (N_8892,N_8458,N_8509);
nand U8893 (N_8893,N_8477,N_8593);
nor U8894 (N_8894,N_8655,N_8501);
or U8895 (N_8895,N_8492,N_8557);
and U8896 (N_8896,N_8484,N_8698);
xor U8897 (N_8897,N_8547,N_8614);
and U8898 (N_8898,N_8443,N_8618);
nand U8899 (N_8899,N_8572,N_8515);
xnor U8900 (N_8900,N_8580,N_8565);
nor U8901 (N_8901,N_8644,N_8682);
nand U8902 (N_8902,N_8464,N_8435);
nor U8903 (N_8903,N_8665,N_8683);
xor U8904 (N_8904,N_8674,N_8487);
xnor U8905 (N_8905,N_8543,N_8420);
or U8906 (N_8906,N_8417,N_8670);
xor U8907 (N_8907,N_8588,N_8664);
and U8908 (N_8908,N_8511,N_8413);
nand U8909 (N_8909,N_8421,N_8664);
nor U8910 (N_8910,N_8650,N_8408);
xnor U8911 (N_8911,N_8581,N_8593);
or U8912 (N_8912,N_8504,N_8437);
and U8913 (N_8913,N_8658,N_8496);
nor U8914 (N_8914,N_8666,N_8435);
and U8915 (N_8915,N_8470,N_8557);
and U8916 (N_8916,N_8417,N_8599);
and U8917 (N_8917,N_8546,N_8697);
nor U8918 (N_8918,N_8586,N_8469);
xnor U8919 (N_8919,N_8521,N_8549);
nand U8920 (N_8920,N_8618,N_8495);
or U8921 (N_8921,N_8460,N_8518);
and U8922 (N_8922,N_8649,N_8514);
nand U8923 (N_8923,N_8593,N_8552);
nand U8924 (N_8924,N_8411,N_8569);
or U8925 (N_8925,N_8440,N_8508);
or U8926 (N_8926,N_8537,N_8557);
or U8927 (N_8927,N_8565,N_8698);
nand U8928 (N_8928,N_8489,N_8586);
and U8929 (N_8929,N_8582,N_8678);
or U8930 (N_8930,N_8470,N_8653);
xnor U8931 (N_8931,N_8577,N_8550);
nand U8932 (N_8932,N_8410,N_8534);
nor U8933 (N_8933,N_8527,N_8667);
xor U8934 (N_8934,N_8578,N_8401);
nor U8935 (N_8935,N_8451,N_8693);
xnor U8936 (N_8936,N_8668,N_8679);
or U8937 (N_8937,N_8588,N_8601);
or U8938 (N_8938,N_8481,N_8440);
or U8939 (N_8939,N_8470,N_8418);
xnor U8940 (N_8940,N_8537,N_8541);
nor U8941 (N_8941,N_8448,N_8625);
or U8942 (N_8942,N_8637,N_8459);
nand U8943 (N_8943,N_8621,N_8632);
and U8944 (N_8944,N_8615,N_8651);
and U8945 (N_8945,N_8466,N_8433);
or U8946 (N_8946,N_8632,N_8546);
or U8947 (N_8947,N_8578,N_8626);
xor U8948 (N_8948,N_8561,N_8500);
and U8949 (N_8949,N_8649,N_8455);
or U8950 (N_8950,N_8647,N_8625);
or U8951 (N_8951,N_8454,N_8586);
and U8952 (N_8952,N_8659,N_8481);
nor U8953 (N_8953,N_8435,N_8510);
nand U8954 (N_8954,N_8508,N_8429);
nand U8955 (N_8955,N_8564,N_8448);
nor U8956 (N_8956,N_8433,N_8425);
nand U8957 (N_8957,N_8693,N_8501);
nand U8958 (N_8958,N_8602,N_8639);
and U8959 (N_8959,N_8424,N_8687);
nand U8960 (N_8960,N_8553,N_8515);
xnor U8961 (N_8961,N_8601,N_8478);
and U8962 (N_8962,N_8570,N_8618);
and U8963 (N_8963,N_8432,N_8402);
or U8964 (N_8964,N_8537,N_8552);
nor U8965 (N_8965,N_8419,N_8563);
nand U8966 (N_8966,N_8526,N_8501);
nor U8967 (N_8967,N_8602,N_8409);
or U8968 (N_8968,N_8661,N_8642);
nor U8969 (N_8969,N_8466,N_8604);
and U8970 (N_8970,N_8595,N_8519);
and U8971 (N_8971,N_8543,N_8405);
and U8972 (N_8972,N_8501,N_8550);
nor U8973 (N_8973,N_8416,N_8603);
and U8974 (N_8974,N_8593,N_8536);
and U8975 (N_8975,N_8428,N_8639);
or U8976 (N_8976,N_8546,N_8492);
nor U8977 (N_8977,N_8409,N_8624);
nand U8978 (N_8978,N_8495,N_8582);
nor U8979 (N_8979,N_8662,N_8642);
and U8980 (N_8980,N_8561,N_8492);
nand U8981 (N_8981,N_8418,N_8671);
nand U8982 (N_8982,N_8479,N_8608);
or U8983 (N_8983,N_8412,N_8471);
and U8984 (N_8984,N_8566,N_8686);
nand U8985 (N_8985,N_8422,N_8536);
and U8986 (N_8986,N_8428,N_8523);
nor U8987 (N_8987,N_8589,N_8404);
nand U8988 (N_8988,N_8691,N_8533);
xnor U8989 (N_8989,N_8657,N_8581);
or U8990 (N_8990,N_8495,N_8511);
and U8991 (N_8991,N_8423,N_8506);
xnor U8992 (N_8992,N_8682,N_8480);
and U8993 (N_8993,N_8484,N_8466);
or U8994 (N_8994,N_8434,N_8588);
or U8995 (N_8995,N_8410,N_8666);
and U8996 (N_8996,N_8467,N_8692);
xnor U8997 (N_8997,N_8696,N_8612);
nand U8998 (N_8998,N_8544,N_8461);
nor U8999 (N_8999,N_8676,N_8677);
nand U9000 (N_9000,N_8866,N_8859);
nor U9001 (N_9001,N_8740,N_8850);
or U9002 (N_9002,N_8984,N_8817);
xnor U9003 (N_9003,N_8748,N_8733);
and U9004 (N_9004,N_8729,N_8713);
nand U9005 (N_9005,N_8821,N_8790);
nor U9006 (N_9006,N_8970,N_8929);
nand U9007 (N_9007,N_8775,N_8845);
xor U9008 (N_9008,N_8953,N_8760);
xnor U9009 (N_9009,N_8746,N_8924);
or U9010 (N_9010,N_8962,N_8876);
nand U9011 (N_9011,N_8855,N_8847);
and U9012 (N_9012,N_8762,N_8761);
and U9013 (N_9013,N_8884,N_8741);
or U9014 (N_9014,N_8702,N_8800);
or U9015 (N_9015,N_8710,N_8923);
nand U9016 (N_9016,N_8773,N_8808);
xor U9017 (N_9017,N_8933,N_8812);
and U9018 (N_9018,N_8901,N_8801);
nor U9019 (N_9019,N_8736,N_8872);
or U9020 (N_9020,N_8707,N_8827);
and U9021 (N_9021,N_8849,N_8758);
and U9022 (N_9022,N_8816,N_8788);
and U9023 (N_9023,N_8871,N_8907);
nor U9024 (N_9024,N_8873,N_8798);
nor U9025 (N_9025,N_8779,N_8753);
or U9026 (N_9026,N_8770,N_8759);
xnor U9027 (N_9027,N_8730,N_8720);
nor U9028 (N_9028,N_8774,N_8874);
nor U9029 (N_9029,N_8834,N_8910);
or U9030 (N_9030,N_8818,N_8882);
xor U9031 (N_9031,N_8795,N_8880);
nand U9032 (N_9032,N_8996,N_8757);
or U9033 (N_9033,N_8949,N_8714);
or U9034 (N_9034,N_8991,N_8727);
xor U9035 (N_9035,N_8947,N_8836);
or U9036 (N_9036,N_8703,N_8913);
or U9037 (N_9037,N_8792,N_8941);
and U9038 (N_9038,N_8771,N_8765);
xor U9039 (N_9039,N_8781,N_8886);
nor U9040 (N_9040,N_8930,N_8755);
xnor U9041 (N_9041,N_8980,N_8887);
nor U9042 (N_9042,N_8854,N_8749);
xnor U9043 (N_9043,N_8899,N_8701);
nand U9044 (N_9044,N_8853,N_8752);
nand U9045 (N_9045,N_8920,N_8868);
nor U9046 (N_9046,N_8903,N_8772);
xor U9047 (N_9047,N_8927,N_8754);
xnor U9048 (N_9048,N_8835,N_8785);
and U9049 (N_9049,N_8802,N_8909);
nor U9050 (N_9050,N_8906,N_8894);
and U9051 (N_9051,N_8726,N_8877);
nand U9052 (N_9052,N_8994,N_8968);
or U9053 (N_9053,N_8807,N_8964);
and U9054 (N_9054,N_8796,N_8756);
xnor U9055 (N_9055,N_8965,N_8922);
nor U9056 (N_9056,N_8857,N_8722);
and U9057 (N_9057,N_8958,N_8982);
and U9058 (N_9058,N_8926,N_8875);
and U9059 (N_9059,N_8879,N_8784);
or U9060 (N_9060,N_8969,N_8711);
nand U9061 (N_9061,N_8723,N_8916);
nor U9062 (N_9062,N_8799,N_8995);
nor U9063 (N_9063,N_8786,N_8981);
xor U9064 (N_9064,N_8938,N_8724);
nand U9065 (N_9065,N_8791,N_8700);
and U9066 (N_9066,N_8851,N_8731);
and U9067 (N_9067,N_8768,N_8867);
nor U9068 (N_9068,N_8750,N_8805);
and U9069 (N_9069,N_8833,N_8862);
nand U9070 (N_9070,N_8732,N_8946);
xnor U9071 (N_9071,N_8921,N_8815);
nor U9072 (N_9072,N_8937,N_8908);
xnor U9073 (N_9073,N_8863,N_8904);
nor U9074 (N_9074,N_8806,N_8888);
and U9075 (N_9075,N_8954,N_8897);
nor U9076 (N_9076,N_8979,N_8811);
nand U9077 (N_9077,N_8990,N_8870);
or U9078 (N_9078,N_8782,N_8989);
nor U9079 (N_9079,N_8764,N_8780);
xnor U9080 (N_9080,N_8900,N_8992);
or U9081 (N_9081,N_8842,N_8813);
or U9082 (N_9082,N_8824,N_8885);
nand U9083 (N_9083,N_8902,N_8721);
nand U9084 (N_9084,N_8844,N_8744);
and U9085 (N_9085,N_8819,N_8967);
xor U9086 (N_9086,N_8858,N_8919);
or U9087 (N_9087,N_8925,N_8794);
or U9088 (N_9088,N_8940,N_8956);
or U9089 (N_9089,N_8843,N_8715);
xnor U9090 (N_9090,N_8978,N_8963);
nor U9091 (N_9091,N_8735,N_8889);
nand U9092 (N_9092,N_8890,N_8892);
xnor U9093 (N_9093,N_8783,N_8972);
and U9094 (N_9094,N_8896,N_8828);
nor U9095 (N_9095,N_8942,N_8814);
nand U9096 (N_9096,N_8839,N_8777);
or U9097 (N_9097,N_8738,N_8955);
nor U9098 (N_9098,N_8999,N_8986);
or U9099 (N_9099,N_8905,N_8734);
xor U9100 (N_9100,N_8911,N_8831);
and U9101 (N_9101,N_8725,N_8705);
and U9102 (N_9102,N_8830,N_8763);
and U9103 (N_9103,N_8769,N_8932);
and U9104 (N_9104,N_8832,N_8966);
or U9105 (N_9105,N_8977,N_8829);
xor U9106 (N_9106,N_8718,N_8864);
nand U9107 (N_9107,N_8739,N_8914);
and U9108 (N_9108,N_8820,N_8883);
xnor U9109 (N_9109,N_8809,N_8993);
xor U9110 (N_9110,N_8934,N_8823);
xnor U9111 (N_9111,N_8975,N_8797);
and U9112 (N_9112,N_8944,N_8787);
nor U9113 (N_9113,N_8852,N_8895);
or U9114 (N_9114,N_8861,N_8767);
nand U9115 (N_9115,N_8959,N_8988);
and U9116 (N_9116,N_8743,N_8751);
or U9117 (N_9117,N_8745,N_8973);
or U9118 (N_9118,N_8793,N_8804);
nand U9119 (N_9119,N_8838,N_8974);
nand U9120 (N_9120,N_8840,N_8961);
nor U9121 (N_9121,N_8837,N_8825);
xnor U9122 (N_9122,N_8841,N_8860);
nor U9123 (N_9123,N_8960,N_8948);
xor U9124 (N_9124,N_8881,N_8865);
nand U9125 (N_9125,N_8951,N_8976);
xor U9126 (N_9126,N_8945,N_8848);
and U9127 (N_9127,N_8998,N_8737);
nand U9128 (N_9128,N_8822,N_8708);
nor U9129 (N_9129,N_8766,N_8931);
nand U9130 (N_9130,N_8846,N_8997);
or U9131 (N_9131,N_8912,N_8928);
nor U9132 (N_9132,N_8893,N_8987);
xor U9133 (N_9133,N_8898,N_8706);
nor U9134 (N_9134,N_8957,N_8728);
and U9135 (N_9135,N_8936,N_8935);
nand U9136 (N_9136,N_8789,N_8952);
xnor U9137 (N_9137,N_8826,N_8712);
xor U9138 (N_9138,N_8776,N_8803);
and U9139 (N_9139,N_8747,N_8742);
or U9140 (N_9140,N_8915,N_8971);
and U9141 (N_9141,N_8943,N_8950);
nand U9142 (N_9142,N_8891,N_8869);
and U9143 (N_9143,N_8810,N_8709);
or U9144 (N_9144,N_8878,N_8939);
xnor U9145 (N_9145,N_8985,N_8778);
or U9146 (N_9146,N_8918,N_8704);
xnor U9147 (N_9147,N_8856,N_8717);
xnor U9148 (N_9148,N_8917,N_8719);
or U9149 (N_9149,N_8716,N_8983);
and U9150 (N_9150,N_8829,N_8844);
nand U9151 (N_9151,N_8962,N_8735);
xnor U9152 (N_9152,N_8754,N_8922);
and U9153 (N_9153,N_8783,N_8744);
nand U9154 (N_9154,N_8884,N_8738);
nand U9155 (N_9155,N_8970,N_8721);
or U9156 (N_9156,N_8787,N_8871);
nand U9157 (N_9157,N_8875,N_8986);
nor U9158 (N_9158,N_8868,N_8805);
nor U9159 (N_9159,N_8800,N_8928);
nor U9160 (N_9160,N_8899,N_8836);
or U9161 (N_9161,N_8998,N_8889);
and U9162 (N_9162,N_8975,N_8833);
and U9163 (N_9163,N_8853,N_8885);
xor U9164 (N_9164,N_8987,N_8779);
nor U9165 (N_9165,N_8935,N_8791);
nor U9166 (N_9166,N_8900,N_8771);
and U9167 (N_9167,N_8902,N_8787);
and U9168 (N_9168,N_8908,N_8928);
xor U9169 (N_9169,N_8922,N_8931);
nand U9170 (N_9170,N_8964,N_8750);
or U9171 (N_9171,N_8931,N_8851);
nand U9172 (N_9172,N_8964,N_8836);
xnor U9173 (N_9173,N_8702,N_8908);
xnor U9174 (N_9174,N_8922,N_8912);
nand U9175 (N_9175,N_8960,N_8853);
or U9176 (N_9176,N_8729,N_8764);
xnor U9177 (N_9177,N_8874,N_8850);
and U9178 (N_9178,N_8816,N_8710);
or U9179 (N_9179,N_8819,N_8738);
and U9180 (N_9180,N_8738,N_8809);
xnor U9181 (N_9181,N_8926,N_8708);
nor U9182 (N_9182,N_8996,N_8744);
xor U9183 (N_9183,N_8909,N_8957);
or U9184 (N_9184,N_8797,N_8859);
xor U9185 (N_9185,N_8856,N_8862);
xor U9186 (N_9186,N_8972,N_8722);
or U9187 (N_9187,N_8737,N_8802);
xnor U9188 (N_9188,N_8952,N_8744);
xor U9189 (N_9189,N_8966,N_8987);
nand U9190 (N_9190,N_8776,N_8983);
xnor U9191 (N_9191,N_8883,N_8815);
or U9192 (N_9192,N_8922,N_8972);
nor U9193 (N_9193,N_8877,N_8786);
nor U9194 (N_9194,N_8986,N_8771);
nand U9195 (N_9195,N_8921,N_8821);
and U9196 (N_9196,N_8735,N_8829);
or U9197 (N_9197,N_8791,N_8895);
xnor U9198 (N_9198,N_8785,N_8715);
nand U9199 (N_9199,N_8892,N_8784);
and U9200 (N_9200,N_8866,N_8799);
or U9201 (N_9201,N_8970,N_8799);
or U9202 (N_9202,N_8776,N_8945);
nand U9203 (N_9203,N_8940,N_8820);
nand U9204 (N_9204,N_8942,N_8819);
nand U9205 (N_9205,N_8923,N_8967);
nand U9206 (N_9206,N_8918,N_8820);
or U9207 (N_9207,N_8814,N_8849);
or U9208 (N_9208,N_8771,N_8833);
or U9209 (N_9209,N_8773,N_8972);
nor U9210 (N_9210,N_8936,N_8991);
nand U9211 (N_9211,N_8721,N_8799);
xor U9212 (N_9212,N_8887,N_8877);
nand U9213 (N_9213,N_8710,N_8939);
or U9214 (N_9214,N_8940,N_8744);
nor U9215 (N_9215,N_8746,N_8984);
or U9216 (N_9216,N_8769,N_8974);
nor U9217 (N_9217,N_8932,N_8849);
or U9218 (N_9218,N_8765,N_8841);
xnor U9219 (N_9219,N_8962,N_8880);
or U9220 (N_9220,N_8724,N_8774);
and U9221 (N_9221,N_8836,N_8934);
xor U9222 (N_9222,N_8797,N_8983);
xor U9223 (N_9223,N_8972,N_8810);
nand U9224 (N_9224,N_8890,N_8862);
xnor U9225 (N_9225,N_8900,N_8918);
and U9226 (N_9226,N_8795,N_8711);
nand U9227 (N_9227,N_8859,N_8732);
nand U9228 (N_9228,N_8993,N_8734);
or U9229 (N_9229,N_8990,N_8874);
xnor U9230 (N_9230,N_8994,N_8835);
nand U9231 (N_9231,N_8750,N_8811);
nor U9232 (N_9232,N_8984,N_8794);
nor U9233 (N_9233,N_8981,N_8759);
nor U9234 (N_9234,N_8902,N_8725);
xor U9235 (N_9235,N_8958,N_8796);
and U9236 (N_9236,N_8738,N_8876);
nand U9237 (N_9237,N_8752,N_8892);
nor U9238 (N_9238,N_8964,N_8995);
xnor U9239 (N_9239,N_8749,N_8774);
or U9240 (N_9240,N_8743,N_8825);
or U9241 (N_9241,N_8942,N_8834);
and U9242 (N_9242,N_8957,N_8863);
nor U9243 (N_9243,N_8823,N_8767);
xnor U9244 (N_9244,N_8794,N_8766);
and U9245 (N_9245,N_8989,N_8927);
and U9246 (N_9246,N_8812,N_8833);
nor U9247 (N_9247,N_8869,N_8704);
or U9248 (N_9248,N_8902,N_8707);
nand U9249 (N_9249,N_8712,N_8900);
nand U9250 (N_9250,N_8735,N_8900);
and U9251 (N_9251,N_8704,N_8982);
nor U9252 (N_9252,N_8792,N_8868);
nor U9253 (N_9253,N_8793,N_8954);
xnor U9254 (N_9254,N_8907,N_8797);
nor U9255 (N_9255,N_8951,N_8776);
nor U9256 (N_9256,N_8811,N_8996);
nand U9257 (N_9257,N_8899,N_8869);
xnor U9258 (N_9258,N_8888,N_8847);
nand U9259 (N_9259,N_8822,N_8912);
or U9260 (N_9260,N_8991,N_8924);
nor U9261 (N_9261,N_8869,N_8731);
or U9262 (N_9262,N_8772,N_8704);
nand U9263 (N_9263,N_8785,N_8897);
nand U9264 (N_9264,N_8745,N_8887);
nand U9265 (N_9265,N_8970,N_8704);
and U9266 (N_9266,N_8761,N_8731);
and U9267 (N_9267,N_8713,N_8876);
nand U9268 (N_9268,N_8954,N_8935);
nand U9269 (N_9269,N_8958,N_8944);
and U9270 (N_9270,N_8885,N_8961);
nand U9271 (N_9271,N_8967,N_8766);
nor U9272 (N_9272,N_8853,N_8870);
or U9273 (N_9273,N_8948,N_8740);
xor U9274 (N_9274,N_8777,N_8701);
and U9275 (N_9275,N_8918,N_8734);
or U9276 (N_9276,N_8918,N_8851);
or U9277 (N_9277,N_8730,N_8774);
nand U9278 (N_9278,N_8798,N_8936);
nand U9279 (N_9279,N_8704,N_8908);
or U9280 (N_9280,N_8812,N_8886);
nor U9281 (N_9281,N_8744,N_8767);
and U9282 (N_9282,N_8921,N_8836);
nor U9283 (N_9283,N_8847,N_8933);
xnor U9284 (N_9284,N_8931,N_8910);
and U9285 (N_9285,N_8789,N_8723);
nand U9286 (N_9286,N_8804,N_8937);
or U9287 (N_9287,N_8899,N_8801);
xor U9288 (N_9288,N_8886,N_8844);
xnor U9289 (N_9289,N_8759,N_8848);
xor U9290 (N_9290,N_8779,N_8790);
or U9291 (N_9291,N_8802,N_8947);
and U9292 (N_9292,N_8862,N_8726);
and U9293 (N_9293,N_8950,N_8995);
xor U9294 (N_9294,N_8733,N_8864);
xnor U9295 (N_9295,N_8785,N_8779);
and U9296 (N_9296,N_8734,N_8833);
nor U9297 (N_9297,N_8845,N_8808);
and U9298 (N_9298,N_8930,N_8921);
and U9299 (N_9299,N_8795,N_8709);
xnor U9300 (N_9300,N_9076,N_9090);
xnor U9301 (N_9301,N_9271,N_9080);
nor U9302 (N_9302,N_9246,N_9206);
xor U9303 (N_9303,N_9019,N_9263);
or U9304 (N_9304,N_9038,N_9216);
nor U9305 (N_9305,N_9033,N_9297);
xnor U9306 (N_9306,N_9266,N_9186);
nand U9307 (N_9307,N_9183,N_9131);
nor U9308 (N_9308,N_9064,N_9047);
nor U9309 (N_9309,N_9114,N_9022);
nor U9310 (N_9310,N_9168,N_9095);
or U9311 (N_9311,N_9214,N_9036);
xnor U9312 (N_9312,N_9145,N_9283);
or U9313 (N_9313,N_9065,N_9136);
nor U9314 (N_9314,N_9202,N_9282);
and U9315 (N_9315,N_9225,N_9166);
and U9316 (N_9316,N_9151,N_9245);
nand U9317 (N_9317,N_9226,N_9133);
and U9318 (N_9318,N_9107,N_9143);
nor U9319 (N_9319,N_9296,N_9024);
xor U9320 (N_9320,N_9199,N_9190);
xor U9321 (N_9321,N_9126,N_9005);
xnor U9322 (N_9322,N_9039,N_9244);
xnor U9323 (N_9323,N_9258,N_9276);
nor U9324 (N_9324,N_9123,N_9121);
nand U9325 (N_9325,N_9285,N_9068);
xor U9326 (N_9326,N_9072,N_9223);
or U9327 (N_9327,N_9178,N_9132);
nor U9328 (N_9328,N_9012,N_9164);
or U9329 (N_9329,N_9015,N_9293);
xor U9330 (N_9330,N_9008,N_9248);
or U9331 (N_9331,N_9141,N_9144);
nor U9332 (N_9332,N_9174,N_9254);
nor U9333 (N_9333,N_9086,N_9111);
xnor U9334 (N_9334,N_9270,N_9099);
nand U9335 (N_9335,N_9284,N_9208);
or U9336 (N_9336,N_9235,N_9070);
xnor U9337 (N_9337,N_9085,N_9273);
nand U9338 (N_9338,N_9063,N_9057);
xnor U9339 (N_9339,N_9045,N_9134);
or U9340 (N_9340,N_9120,N_9105);
or U9341 (N_9341,N_9148,N_9251);
and U9342 (N_9342,N_9295,N_9272);
and U9343 (N_9343,N_9067,N_9156);
nor U9344 (N_9344,N_9212,N_9058);
nor U9345 (N_9345,N_9221,N_9103);
or U9346 (N_9346,N_9259,N_9192);
nand U9347 (N_9347,N_9138,N_9147);
nor U9348 (N_9348,N_9053,N_9242);
and U9349 (N_9349,N_9205,N_9098);
and U9350 (N_9350,N_9219,N_9267);
nor U9351 (N_9351,N_9004,N_9243);
or U9352 (N_9352,N_9218,N_9016);
nand U9353 (N_9353,N_9287,N_9171);
nor U9354 (N_9354,N_9001,N_9298);
nand U9355 (N_9355,N_9239,N_9207);
nor U9356 (N_9356,N_9288,N_9021);
or U9357 (N_9357,N_9203,N_9083);
nand U9358 (N_9358,N_9055,N_9198);
or U9359 (N_9359,N_9250,N_9152);
and U9360 (N_9360,N_9130,N_9092);
xor U9361 (N_9361,N_9277,N_9252);
and U9362 (N_9362,N_9172,N_9112);
or U9363 (N_9363,N_9094,N_9142);
xor U9364 (N_9364,N_9281,N_9291);
or U9365 (N_9365,N_9265,N_9052);
nand U9366 (N_9366,N_9180,N_9169);
and U9367 (N_9367,N_9191,N_9135);
nand U9368 (N_9368,N_9255,N_9077);
and U9369 (N_9369,N_9071,N_9153);
or U9370 (N_9370,N_9179,N_9013);
and U9371 (N_9371,N_9034,N_9173);
or U9372 (N_9372,N_9032,N_9200);
xor U9373 (N_9373,N_9149,N_9014);
nand U9374 (N_9374,N_9238,N_9280);
and U9375 (N_9375,N_9049,N_9119);
and U9376 (N_9376,N_9247,N_9158);
and U9377 (N_9377,N_9232,N_9162);
and U9378 (N_9378,N_9035,N_9117);
and U9379 (N_9379,N_9177,N_9181);
nand U9380 (N_9380,N_9044,N_9011);
or U9381 (N_9381,N_9220,N_9194);
or U9382 (N_9382,N_9066,N_9006);
or U9383 (N_9383,N_9050,N_9222);
or U9384 (N_9384,N_9185,N_9118);
and U9385 (N_9385,N_9201,N_9278);
xnor U9386 (N_9386,N_9028,N_9184);
xnor U9387 (N_9387,N_9088,N_9160);
and U9388 (N_9388,N_9017,N_9213);
nand U9389 (N_9389,N_9182,N_9228);
xor U9390 (N_9390,N_9079,N_9127);
xnor U9391 (N_9391,N_9087,N_9110);
nor U9392 (N_9392,N_9292,N_9150);
nor U9393 (N_9393,N_9018,N_9204);
or U9394 (N_9394,N_9093,N_9078);
nand U9395 (N_9395,N_9230,N_9262);
or U9396 (N_9396,N_9188,N_9109);
xnor U9397 (N_9397,N_9101,N_9268);
or U9398 (N_9398,N_9189,N_9187);
xor U9399 (N_9399,N_9113,N_9040);
xnor U9400 (N_9400,N_9031,N_9196);
or U9401 (N_9401,N_9037,N_9211);
nand U9402 (N_9402,N_9003,N_9096);
nor U9403 (N_9403,N_9157,N_9124);
or U9404 (N_9404,N_9020,N_9089);
nor U9405 (N_9405,N_9240,N_9106);
nand U9406 (N_9406,N_9261,N_9163);
xnor U9407 (N_9407,N_9227,N_9299);
xnor U9408 (N_9408,N_9084,N_9069);
and U9409 (N_9409,N_9061,N_9217);
or U9410 (N_9410,N_9074,N_9215);
or U9411 (N_9411,N_9231,N_9116);
or U9412 (N_9412,N_9275,N_9073);
nor U9413 (N_9413,N_9193,N_9097);
xor U9414 (N_9414,N_9002,N_9146);
or U9415 (N_9415,N_9026,N_9048);
and U9416 (N_9416,N_9170,N_9023);
and U9417 (N_9417,N_9054,N_9104);
xor U9418 (N_9418,N_9286,N_9294);
or U9419 (N_9419,N_9102,N_9122);
nor U9420 (N_9420,N_9241,N_9269);
or U9421 (N_9421,N_9140,N_9257);
nand U9422 (N_9422,N_9009,N_9091);
or U9423 (N_9423,N_9056,N_9210);
nand U9424 (N_9424,N_9042,N_9165);
nor U9425 (N_9425,N_9197,N_9253);
xnor U9426 (N_9426,N_9115,N_9233);
or U9427 (N_9427,N_9025,N_9161);
and U9428 (N_9428,N_9081,N_9125);
xor U9429 (N_9429,N_9229,N_9029);
or U9430 (N_9430,N_9137,N_9129);
xnor U9431 (N_9431,N_9224,N_9100);
nand U9432 (N_9432,N_9051,N_9256);
or U9433 (N_9433,N_9060,N_9236);
and U9434 (N_9434,N_9128,N_9139);
xor U9435 (N_9435,N_9159,N_9167);
or U9436 (N_9436,N_9249,N_9154);
and U9437 (N_9437,N_9176,N_9279);
xor U9438 (N_9438,N_9062,N_9209);
nand U9439 (N_9439,N_9264,N_9289);
or U9440 (N_9440,N_9290,N_9108);
or U9441 (N_9441,N_9234,N_9059);
nor U9442 (N_9442,N_9274,N_9010);
or U9443 (N_9443,N_9041,N_9260);
nand U9444 (N_9444,N_9195,N_9155);
or U9445 (N_9445,N_9046,N_9030);
and U9446 (N_9446,N_9043,N_9000);
nor U9447 (N_9447,N_9082,N_9027);
or U9448 (N_9448,N_9075,N_9175);
xnor U9449 (N_9449,N_9237,N_9007);
xor U9450 (N_9450,N_9069,N_9269);
nand U9451 (N_9451,N_9255,N_9182);
nor U9452 (N_9452,N_9078,N_9121);
xor U9453 (N_9453,N_9012,N_9131);
xor U9454 (N_9454,N_9203,N_9037);
nor U9455 (N_9455,N_9242,N_9009);
xnor U9456 (N_9456,N_9194,N_9236);
nor U9457 (N_9457,N_9225,N_9170);
xor U9458 (N_9458,N_9244,N_9066);
nor U9459 (N_9459,N_9268,N_9207);
nand U9460 (N_9460,N_9082,N_9111);
and U9461 (N_9461,N_9194,N_9055);
nor U9462 (N_9462,N_9070,N_9206);
xor U9463 (N_9463,N_9163,N_9081);
nor U9464 (N_9464,N_9222,N_9209);
nand U9465 (N_9465,N_9200,N_9093);
nand U9466 (N_9466,N_9155,N_9234);
nand U9467 (N_9467,N_9078,N_9034);
nand U9468 (N_9468,N_9206,N_9047);
nor U9469 (N_9469,N_9285,N_9132);
or U9470 (N_9470,N_9030,N_9119);
xnor U9471 (N_9471,N_9178,N_9054);
and U9472 (N_9472,N_9197,N_9213);
or U9473 (N_9473,N_9246,N_9213);
or U9474 (N_9474,N_9160,N_9236);
and U9475 (N_9475,N_9179,N_9014);
and U9476 (N_9476,N_9006,N_9027);
xnor U9477 (N_9477,N_9200,N_9262);
nand U9478 (N_9478,N_9149,N_9208);
nor U9479 (N_9479,N_9263,N_9169);
nor U9480 (N_9480,N_9044,N_9132);
nand U9481 (N_9481,N_9290,N_9063);
xnor U9482 (N_9482,N_9002,N_9014);
or U9483 (N_9483,N_9213,N_9097);
or U9484 (N_9484,N_9270,N_9155);
and U9485 (N_9485,N_9195,N_9128);
xor U9486 (N_9486,N_9072,N_9130);
nand U9487 (N_9487,N_9099,N_9017);
and U9488 (N_9488,N_9198,N_9234);
nor U9489 (N_9489,N_9174,N_9000);
nor U9490 (N_9490,N_9149,N_9250);
nand U9491 (N_9491,N_9074,N_9055);
nand U9492 (N_9492,N_9151,N_9109);
nand U9493 (N_9493,N_9174,N_9290);
nor U9494 (N_9494,N_9253,N_9121);
nand U9495 (N_9495,N_9011,N_9050);
xnor U9496 (N_9496,N_9260,N_9142);
nand U9497 (N_9497,N_9053,N_9237);
xor U9498 (N_9498,N_9236,N_9013);
nor U9499 (N_9499,N_9209,N_9032);
or U9500 (N_9500,N_9168,N_9159);
nand U9501 (N_9501,N_9277,N_9201);
nand U9502 (N_9502,N_9174,N_9054);
and U9503 (N_9503,N_9016,N_9101);
nor U9504 (N_9504,N_9176,N_9087);
nor U9505 (N_9505,N_9012,N_9066);
nor U9506 (N_9506,N_9131,N_9197);
xnor U9507 (N_9507,N_9007,N_9299);
nor U9508 (N_9508,N_9238,N_9203);
and U9509 (N_9509,N_9157,N_9126);
nand U9510 (N_9510,N_9021,N_9136);
or U9511 (N_9511,N_9129,N_9191);
nand U9512 (N_9512,N_9210,N_9032);
and U9513 (N_9513,N_9091,N_9253);
xnor U9514 (N_9514,N_9131,N_9243);
nor U9515 (N_9515,N_9203,N_9021);
nand U9516 (N_9516,N_9156,N_9120);
nor U9517 (N_9517,N_9004,N_9089);
and U9518 (N_9518,N_9185,N_9233);
nand U9519 (N_9519,N_9208,N_9141);
nor U9520 (N_9520,N_9096,N_9066);
xor U9521 (N_9521,N_9265,N_9298);
and U9522 (N_9522,N_9089,N_9159);
nand U9523 (N_9523,N_9285,N_9120);
xor U9524 (N_9524,N_9259,N_9297);
nand U9525 (N_9525,N_9210,N_9214);
and U9526 (N_9526,N_9238,N_9049);
nand U9527 (N_9527,N_9211,N_9223);
or U9528 (N_9528,N_9176,N_9139);
and U9529 (N_9529,N_9210,N_9159);
xnor U9530 (N_9530,N_9095,N_9167);
nand U9531 (N_9531,N_9117,N_9262);
nand U9532 (N_9532,N_9228,N_9177);
nand U9533 (N_9533,N_9214,N_9240);
and U9534 (N_9534,N_9046,N_9020);
xnor U9535 (N_9535,N_9072,N_9294);
and U9536 (N_9536,N_9167,N_9089);
nand U9537 (N_9537,N_9091,N_9163);
and U9538 (N_9538,N_9089,N_9258);
nand U9539 (N_9539,N_9181,N_9288);
xnor U9540 (N_9540,N_9015,N_9134);
xor U9541 (N_9541,N_9157,N_9174);
and U9542 (N_9542,N_9082,N_9135);
or U9543 (N_9543,N_9249,N_9299);
or U9544 (N_9544,N_9042,N_9265);
xor U9545 (N_9545,N_9232,N_9229);
xor U9546 (N_9546,N_9103,N_9117);
nand U9547 (N_9547,N_9131,N_9255);
or U9548 (N_9548,N_9266,N_9171);
or U9549 (N_9549,N_9210,N_9080);
or U9550 (N_9550,N_9213,N_9107);
or U9551 (N_9551,N_9004,N_9286);
nor U9552 (N_9552,N_9096,N_9158);
and U9553 (N_9553,N_9122,N_9236);
nand U9554 (N_9554,N_9056,N_9003);
xnor U9555 (N_9555,N_9004,N_9100);
and U9556 (N_9556,N_9197,N_9034);
nand U9557 (N_9557,N_9091,N_9155);
nand U9558 (N_9558,N_9219,N_9164);
xor U9559 (N_9559,N_9287,N_9258);
nand U9560 (N_9560,N_9142,N_9084);
or U9561 (N_9561,N_9015,N_9022);
or U9562 (N_9562,N_9199,N_9043);
and U9563 (N_9563,N_9219,N_9258);
nor U9564 (N_9564,N_9005,N_9233);
nand U9565 (N_9565,N_9263,N_9218);
xnor U9566 (N_9566,N_9226,N_9270);
xor U9567 (N_9567,N_9288,N_9262);
nor U9568 (N_9568,N_9278,N_9142);
nor U9569 (N_9569,N_9098,N_9155);
and U9570 (N_9570,N_9128,N_9118);
nand U9571 (N_9571,N_9211,N_9298);
nand U9572 (N_9572,N_9254,N_9165);
or U9573 (N_9573,N_9007,N_9056);
and U9574 (N_9574,N_9048,N_9146);
or U9575 (N_9575,N_9018,N_9065);
and U9576 (N_9576,N_9109,N_9217);
and U9577 (N_9577,N_9120,N_9264);
xnor U9578 (N_9578,N_9078,N_9271);
xor U9579 (N_9579,N_9042,N_9253);
and U9580 (N_9580,N_9005,N_9031);
or U9581 (N_9581,N_9045,N_9279);
or U9582 (N_9582,N_9081,N_9227);
xor U9583 (N_9583,N_9161,N_9230);
and U9584 (N_9584,N_9103,N_9020);
and U9585 (N_9585,N_9071,N_9050);
xor U9586 (N_9586,N_9102,N_9118);
nor U9587 (N_9587,N_9236,N_9225);
and U9588 (N_9588,N_9151,N_9285);
or U9589 (N_9589,N_9170,N_9296);
nand U9590 (N_9590,N_9034,N_9144);
nor U9591 (N_9591,N_9228,N_9003);
or U9592 (N_9592,N_9140,N_9234);
nor U9593 (N_9593,N_9142,N_9284);
nor U9594 (N_9594,N_9277,N_9288);
nand U9595 (N_9595,N_9147,N_9188);
nor U9596 (N_9596,N_9096,N_9036);
and U9597 (N_9597,N_9015,N_9282);
nor U9598 (N_9598,N_9240,N_9096);
or U9599 (N_9599,N_9282,N_9018);
and U9600 (N_9600,N_9315,N_9415);
nand U9601 (N_9601,N_9596,N_9494);
nand U9602 (N_9602,N_9312,N_9443);
or U9603 (N_9603,N_9322,N_9481);
nor U9604 (N_9604,N_9462,N_9525);
nand U9605 (N_9605,N_9377,N_9498);
or U9606 (N_9606,N_9533,N_9516);
nand U9607 (N_9607,N_9334,N_9382);
and U9608 (N_9608,N_9590,N_9486);
nor U9609 (N_9609,N_9302,N_9563);
and U9610 (N_9610,N_9501,N_9305);
or U9611 (N_9611,N_9544,N_9562);
nand U9612 (N_9612,N_9364,N_9500);
nor U9613 (N_9613,N_9450,N_9509);
nand U9614 (N_9614,N_9300,N_9582);
xor U9615 (N_9615,N_9507,N_9348);
or U9616 (N_9616,N_9577,N_9327);
nor U9617 (N_9617,N_9513,N_9461);
and U9618 (N_9618,N_9362,N_9324);
nor U9619 (N_9619,N_9502,N_9354);
nand U9620 (N_9620,N_9424,N_9534);
or U9621 (N_9621,N_9381,N_9579);
nor U9622 (N_9622,N_9587,N_9369);
nor U9623 (N_9623,N_9361,N_9368);
nand U9624 (N_9624,N_9447,N_9379);
and U9625 (N_9625,N_9313,N_9426);
xnor U9626 (N_9626,N_9521,N_9431);
nor U9627 (N_9627,N_9331,N_9458);
nor U9628 (N_9628,N_9383,N_9565);
nor U9629 (N_9629,N_9482,N_9335);
and U9630 (N_9630,N_9531,N_9572);
nand U9631 (N_9631,N_9540,N_9551);
nand U9632 (N_9632,N_9319,N_9597);
and U9633 (N_9633,N_9445,N_9575);
nor U9634 (N_9634,N_9375,N_9398);
or U9635 (N_9635,N_9317,N_9396);
and U9636 (N_9636,N_9373,N_9439);
nor U9637 (N_9637,N_9469,N_9366);
and U9638 (N_9638,N_9592,N_9511);
nor U9639 (N_9639,N_9350,N_9400);
xor U9640 (N_9640,N_9359,N_9473);
xor U9641 (N_9641,N_9491,N_9515);
nand U9642 (N_9642,N_9490,N_9423);
and U9643 (N_9643,N_9337,N_9588);
xor U9644 (N_9644,N_9306,N_9474);
or U9645 (N_9645,N_9430,N_9332);
nand U9646 (N_9646,N_9310,N_9455);
nor U9647 (N_9647,N_9344,N_9391);
xnor U9648 (N_9648,N_9476,N_9320);
or U9649 (N_9649,N_9360,N_9550);
and U9650 (N_9650,N_9546,N_9330);
nand U9651 (N_9651,N_9496,N_9438);
or U9652 (N_9652,N_9387,N_9418);
nor U9653 (N_9653,N_9542,N_9479);
nor U9654 (N_9654,N_9311,N_9304);
nor U9655 (N_9655,N_9417,N_9483);
nor U9656 (N_9656,N_9598,N_9411);
nor U9657 (N_9657,N_9386,N_9409);
and U9658 (N_9658,N_9547,N_9471);
and U9659 (N_9659,N_9558,N_9584);
nand U9660 (N_9660,N_9341,N_9301);
xnor U9661 (N_9661,N_9349,N_9539);
xnor U9662 (N_9662,N_9543,N_9535);
nor U9663 (N_9663,N_9399,N_9347);
xnor U9664 (N_9664,N_9492,N_9388);
xnor U9665 (N_9665,N_9466,N_9329);
nand U9666 (N_9666,N_9545,N_9568);
nand U9667 (N_9667,N_9581,N_9394);
nand U9668 (N_9668,N_9326,N_9460);
or U9669 (N_9669,N_9356,N_9395);
and U9670 (N_9670,N_9448,N_9374);
nand U9671 (N_9671,N_9453,N_9371);
nand U9672 (N_9672,N_9380,N_9524);
nor U9673 (N_9673,N_9338,N_9555);
and U9674 (N_9674,N_9484,N_9464);
nor U9675 (N_9675,N_9428,N_9487);
nand U9676 (N_9676,N_9336,N_9595);
or U9677 (N_9677,N_9510,N_9569);
and U9678 (N_9678,N_9328,N_9357);
nand U9679 (N_9679,N_9452,N_9316);
xor U9680 (N_9680,N_9591,N_9561);
or U9681 (N_9681,N_9427,N_9342);
or U9682 (N_9682,N_9407,N_9333);
xnor U9683 (N_9683,N_9594,N_9467);
or U9684 (N_9684,N_9422,N_9508);
and U9685 (N_9685,N_9526,N_9583);
xnor U9686 (N_9686,N_9472,N_9536);
xnor U9687 (N_9687,N_9429,N_9389);
nand U9688 (N_9688,N_9570,N_9308);
nand U9689 (N_9689,N_9571,N_9519);
or U9690 (N_9690,N_9573,N_9435);
and U9691 (N_9691,N_9325,N_9378);
xor U9692 (N_9692,N_9437,N_9530);
and U9693 (N_9693,N_9318,N_9390);
and U9694 (N_9694,N_9321,N_9365);
xnor U9695 (N_9695,N_9580,N_9444);
xor U9696 (N_9696,N_9440,N_9537);
nand U9697 (N_9697,N_9557,N_9477);
nor U9698 (N_9698,N_9419,N_9420);
or U9699 (N_9699,N_9401,N_9576);
nor U9700 (N_9700,N_9470,N_9499);
and U9701 (N_9701,N_9505,N_9522);
nor U9702 (N_9702,N_9367,N_9493);
and U9703 (N_9703,N_9463,N_9412);
xnor U9704 (N_9704,N_9434,N_9475);
and U9705 (N_9705,N_9370,N_9345);
xor U9706 (N_9706,N_9405,N_9538);
nor U9707 (N_9707,N_9497,N_9456);
and U9708 (N_9708,N_9413,N_9457);
xor U9709 (N_9709,N_9503,N_9517);
or U9710 (N_9710,N_9441,N_9552);
nor U9711 (N_9711,N_9459,N_9512);
or U9712 (N_9712,N_9346,N_9425);
nor U9713 (N_9713,N_9504,N_9564);
xor U9714 (N_9714,N_9560,N_9323);
nor U9715 (N_9715,N_9410,N_9353);
xnor U9716 (N_9716,N_9397,N_9589);
nor U9717 (N_9717,N_9449,N_9485);
xnor U9718 (N_9718,N_9527,N_9586);
and U9719 (N_9719,N_9355,N_9559);
nand U9720 (N_9720,N_9529,N_9518);
nor U9721 (N_9721,N_9393,N_9436);
xor U9722 (N_9722,N_9451,N_9303);
or U9723 (N_9723,N_9548,N_9480);
nor U9724 (N_9724,N_9468,N_9385);
or U9725 (N_9725,N_9340,N_9556);
xnor U9726 (N_9726,N_9433,N_9372);
or U9727 (N_9727,N_9314,N_9351);
xor U9728 (N_9728,N_9578,N_9309);
nor U9729 (N_9729,N_9532,N_9421);
nor U9730 (N_9730,N_9488,N_9478);
or U9731 (N_9731,N_9432,N_9414);
nand U9732 (N_9732,N_9454,N_9567);
and U9733 (N_9733,N_9402,N_9358);
and U9734 (N_9734,N_9352,N_9593);
xor U9735 (N_9735,N_9343,N_9528);
nor U9736 (N_9736,N_9446,N_9553);
nor U9737 (N_9737,N_9339,N_9566);
nand U9738 (N_9738,N_9599,N_9523);
or U9739 (N_9739,N_9384,N_9406);
or U9740 (N_9740,N_9514,N_9408);
xor U9741 (N_9741,N_9392,N_9541);
and U9742 (N_9742,N_9416,N_9495);
xnor U9743 (N_9743,N_9442,N_9489);
nand U9744 (N_9744,N_9307,N_9554);
xnor U9745 (N_9745,N_9465,N_9403);
nor U9746 (N_9746,N_9376,N_9549);
and U9747 (N_9747,N_9506,N_9404);
nand U9748 (N_9748,N_9363,N_9585);
xor U9749 (N_9749,N_9520,N_9574);
nor U9750 (N_9750,N_9566,N_9553);
and U9751 (N_9751,N_9598,N_9584);
and U9752 (N_9752,N_9541,N_9461);
nor U9753 (N_9753,N_9496,N_9482);
nor U9754 (N_9754,N_9515,N_9554);
and U9755 (N_9755,N_9400,N_9470);
nand U9756 (N_9756,N_9300,N_9586);
and U9757 (N_9757,N_9484,N_9352);
nor U9758 (N_9758,N_9578,N_9446);
xnor U9759 (N_9759,N_9428,N_9458);
xnor U9760 (N_9760,N_9525,N_9592);
or U9761 (N_9761,N_9446,N_9561);
nor U9762 (N_9762,N_9392,N_9367);
or U9763 (N_9763,N_9522,N_9500);
nand U9764 (N_9764,N_9313,N_9321);
xor U9765 (N_9765,N_9517,N_9518);
nand U9766 (N_9766,N_9459,N_9391);
nor U9767 (N_9767,N_9508,N_9580);
and U9768 (N_9768,N_9372,N_9546);
nand U9769 (N_9769,N_9540,N_9438);
and U9770 (N_9770,N_9547,N_9399);
and U9771 (N_9771,N_9450,N_9371);
nor U9772 (N_9772,N_9537,N_9523);
xnor U9773 (N_9773,N_9401,N_9446);
nand U9774 (N_9774,N_9551,N_9536);
and U9775 (N_9775,N_9313,N_9315);
nor U9776 (N_9776,N_9311,N_9307);
nand U9777 (N_9777,N_9467,N_9373);
nor U9778 (N_9778,N_9407,N_9330);
nor U9779 (N_9779,N_9522,N_9536);
nor U9780 (N_9780,N_9539,N_9465);
or U9781 (N_9781,N_9340,N_9424);
xor U9782 (N_9782,N_9392,N_9559);
xor U9783 (N_9783,N_9377,N_9525);
nand U9784 (N_9784,N_9541,N_9489);
and U9785 (N_9785,N_9327,N_9595);
nand U9786 (N_9786,N_9579,N_9491);
nand U9787 (N_9787,N_9400,N_9436);
or U9788 (N_9788,N_9334,N_9392);
nor U9789 (N_9789,N_9571,N_9359);
or U9790 (N_9790,N_9581,N_9481);
nand U9791 (N_9791,N_9375,N_9505);
nand U9792 (N_9792,N_9491,N_9496);
nor U9793 (N_9793,N_9587,N_9368);
nor U9794 (N_9794,N_9471,N_9513);
or U9795 (N_9795,N_9586,N_9457);
nor U9796 (N_9796,N_9370,N_9473);
xnor U9797 (N_9797,N_9522,N_9581);
or U9798 (N_9798,N_9464,N_9350);
nand U9799 (N_9799,N_9579,N_9509);
nor U9800 (N_9800,N_9502,N_9359);
or U9801 (N_9801,N_9586,N_9578);
or U9802 (N_9802,N_9435,N_9587);
or U9803 (N_9803,N_9488,N_9441);
xnor U9804 (N_9804,N_9574,N_9360);
and U9805 (N_9805,N_9551,N_9480);
xnor U9806 (N_9806,N_9557,N_9540);
or U9807 (N_9807,N_9504,N_9374);
nand U9808 (N_9808,N_9410,N_9309);
xnor U9809 (N_9809,N_9526,N_9358);
nor U9810 (N_9810,N_9345,N_9343);
xnor U9811 (N_9811,N_9357,N_9517);
nor U9812 (N_9812,N_9322,N_9438);
and U9813 (N_9813,N_9557,N_9508);
and U9814 (N_9814,N_9598,N_9586);
nand U9815 (N_9815,N_9475,N_9461);
and U9816 (N_9816,N_9596,N_9526);
or U9817 (N_9817,N_9455,N_9542);
and U9818 (N_9818,N_9537,N_9594);
nor U9819 (N_9819,N_9427,N_9316);
nor U9820 (N_9820,N_9596,N_9313);
and U9821 (N_9821,N_9312,N_9301);
xnor U9822 (N_9822,N_9302,N_9475);
nand U9823 (N_9823,N_9301,N_9447);
and U9824 (N_9824,N_9461,N_9445);
or U9825 (N_9825,N_9570,N_9524);
or U9826 (N_9826,N_9499,N_9401);
nand U9827 (N_9827,N_9386,N_9505);
and U9828 (N_9828,N_9460,N_9389);
or U9829 (N_9829,N_9305,N_9360);
xor U9830 (N_9830,N_9309,N_9434);
nor U9831 (N_9831,N_9503,N_9423);
or U9832 (N_9832,N_9370,N_9413);
nand U9833 (N_9833,N_9343,N_9347);
xnor U9834 (N_9834,N_9434,N_9343);
xnor U9835 (N_9835,N_9412,N_9537);
or U9836 (N_9836,N_9568,N_9325);
nor U9837 (N_9837,N_9493,N_9520);
xnor U9838 (N_9838,N_9570,N_9462);
xor U9839 (N_9839,N_9563,N_9536);
xor U9840 (N_9840,N_9545,N_9302);
or U9841 (N_9841,N_9364,N_9566);
or U9842 (N_9842,N_9485,N_9461);
nand U9843 (N_9843,N_9357,N_9547);
nor U9844 (N_9844,N_9403,N_9424);
xnor U9845 (N_9845,N_9348,N_9552);
xnor U9846 (N_9846,N_9323,N_9570);
xor U9847 (N_9847,N_9342,N_9309);
or U9848 (N_9848,N_9399,N_9374);
or U9849 (N_9849,N_9534,N_9435);
xor U9850 (N_9850,N_9347,N_9408);
or U9851 (N_9851,N_9585,N_9406);
nor U9852 (N_9852,N_9586,N_9310);
nor U9853 (N_9853,N_9567,N_9301);
xnor U9854 (N_9854,N_9559,N_9374);
and U9855 (N_9855,N_9379,N_9446);
nor U9856 (N_9856,N_9380,N_9410);
and U9857 (N_9857,N_9481,N_9358);
and U9858 (N_9858,N_9472,N_9411);
or U9859 (N_9859,N_9306,N_9578);
xor U9860 (N_9860,N_9443,N_9558);
and U9861 (N_9861,N_9512,N_9596);
nand U9862 (N_9862,N_9531,N_9566);
nand U9863 (N_9863,N_9306,N_9364);
xnor U9864 (N_9864,N_9453,N_9531);
nor U9865 (N_9865,N_9351,N_9491);
xor U9866 (N_9866,N_9301,N_9339);
or U9867 (N_9867,N_9307,N_9495);
xnor U9868 (N_9868,N_9340,N_9360);
nor U9869 (N_9869,N_9482,N_9411);
and U9870 (N_9870,N_9304,N_9570);
or U9871 (N_9871,N_9562,N_9590);
nor U9872 (N_9872,N_9357,N_9596);
or U9873 (N_9873,N_9467,N_9318);
xor U9874 (N_9874,N_9327,N_9593);
xnor U9875 (N_9875,N_9465,N_9560);
or U9876 (N_9876,N_9302,N_9595);
or U9877 (N_9877,N_9310,N_9428);
nand U9878 (N_9878,N_9535,N_9372);
and U9879 (N_9879,N_9418,N_9542);
xor U9880 (N_9880,N_9320,N_9385);
or U9881 (N_9881,N_9461,N_9586);
nand U9882 (N_9882,N_9455,N_9304);
or U9883 (N_9883,N_9591,N_9487);
or U9884 (N_9884,N_9335,N_9507);
or U9885 (N_9885,N_9511,N_9339);
and U9886 (N_9886,N_9371,N_9341);
nand U9887 (N_9887,N_9342,N_9381);
nand U9888 (N_9888,N_9589,N_9492);
and U9889 (N_9889,N_9497,N_9562);
nor U9890 (N_9890,N_9328,N_9594);
xor U9891 (N_9891,N_9301,N_9527);
nand U9892 (N_9892,N_9468,N_9549);
nand U9893 (N_9893,N_9518,N_9411);
and U9894 (N_9894,N_9424,N_9407);
or U9895 (N_9895,N_9355,N_9475);
and U9896 (N_9896,N_9388,N_9518);
and U9897 (N_9897,N_9331,N_9443);
xor U9898 (N_9898,N_9400,N_9388);
xor U9899 (N_9899,N_9549,N_9479);
nor U9900 (N_9900,N_9897,N_9616);
nor U9901 (N_9901,N_9723,N_9657);
nand U9902 (N_9902,N_9762,N_9670);
nand U9903 (N_9903,N_9649,N_9824);
nand U9904 (N_9904,N_9655,N_9642);
and U9905 (N_9905,N_9730,N_9620);
nor U9906 (N_9906,N_9878,N_9740);
nor U9907 (N_9907,N_9608,N_9892);
xor U9908 (N_9908,N_9708,N_9875);
and U9909 (N_9909,N_9802,N_9782);
nor U9910 (N_9910,N_9725,N_9832);
and U9911 (N_9911,N_9738,N_9793);
nor U9912 (N_9912,N_9803,N_9746);
xor U9913 (N_9913,N_9715,N_9799);
nor U9914 (N_9914,N_9704,N_9894);
nand U9915 (N_9915,N_9646,N_9609);
and U9916 (N_9916,N_9860,N_9805);
or U9917 (N_9917,N_9717,N_9747);
or U9918 (N_9918,N_9656,N_9870);
xor U9919 (N_9919,N_9874,N_9871);
xor U9920 (N_9920,N_9741,N_9882);
nand U9921 (N_9921,N_9696,N_9710);
or U9922 (N_9922,N_9822,N_9893);
nand U9923 (N_9923,N_9677,N_9776);
or U9924 (N_9924,N_9714,N_9823);
nor U9925 (N_9925,N_9669,N_9791);
and U9926 (N_9926,N_9817,N_9826);
and U9927 (N_9927,N_9754,N_9764);
nor U9928 (N_9928,N_9778,N_9682);
nand U9929 (N_9929,N_9859,N_9739);
nor U9930 (N_9930,N_9631,N_9683);
nor U9931 (N_9931,N_9829,N_9775);
and U9932 (N_9932,N_9648,N_9612);
nor U9933 (N_9933,N_9600,N_9872);
xor U9934 (N_9934,N_9877,N_9783);
or U9935 (N_9935,N_9659,N_9852);
nor U9936 (N_9936,N_9667,N_9702);
nand U9937 (N_9937,N_9816,N_9638);
and U9938 (N_9938,N_9845,N_9731);
and U9939 (N_9939,N_9868,N_9804);
xor U9940 (N_9940,N_9774,N_9844);
nand U9941 (N_9941,N_9622,N_9691);
nor U9942 (N_9942,N_9849,N_9742);
and U9943 (N_9943,N_9671,N_9626);
nand U9944 (N_9944,N_9830,N_9607);
or U9945 (N_9945,N_9606,N_9707);
xnor U9946 (N_9946,N_9837,N_9718);
xnor U9947 (N_9947,N_9701,N_9692);
nand U9948 (N_9948,N_9848,N_9767);
or U9949 (N_9949,N_9815,N_9729);
nand U9950 (N_9950,N_9673,N_9780);
nor U9951 (N_9951,N_9760,N_9650);
and U9952 (N_9952,N_9653,N_9895);
nand U9953 (N_9953,N_9689,N_9769);
and U9954 (N_9954,N_9668,N_9621);
nor U9955 (N_9955,N_9821,N_9732);
nand U9956 (N_9956,N_9758,N_9632);
xor U9957 (N_9957,N_9834,N_9685);
and U9958 (N_9958,N_9716,N_9801);
nor U9959 (N_9959,N_9755,N_9627);
and U9960 (N_9960,N_9726,N_9831);
nor U9961 (N_9961,N_9679,N_9789);
xor U9962 (N_9962,N_9863,N_9734);
or U9963 (N_9963,N_9750,N_9820);
and U9964 (N_9964,N_9751,N_9886);
and U9965 (N_9965,N_9641,N_9773);
xor U9966 (N_9966,N_9623,N_9722);
nor U9967 (N_9967,N_9749,N_9856);
nand U9968 (N_9968,N_9675,N_9680);
or U9969 (N_9969,N_9752,N_9633);
and U9970 (N_9970,N_9810,N_9819);
nand U9971 (N_9971,N_9880,N_9744);
xnor U9972 (N_9972,N_9853,N_9728);
or U9973 (N_9973,N_9664,N_9737);
nor U9974 (N_9974,N_9887,N_9881);
xor U9975 (N_9975,N_9889,N_9629);
nand U9976 (N_9976,N_9634,N_9818);
and U9977 (N_9977,N_9809,N_9651);
xor U9978 (N_9978,N_9625,N_9888);
nand U9979 (N_9979,N_9645,N_9765);
or U9980 (N_9980,N_9806,N_9637);
nor U9981 (N_9981,N_9613,N_9727);
and U9982 (N_9982,N_9733,N_9647);
xnor U9983 (N_9983,N_9869,N_9743);
nand U9984 (N_9984,N_9772,N_9858);
xor U9985 (N_9985,N_9720,N_9786);
or U9986 (N_9986,N_9601,N_9896);
nor U9987 (N_9987,N_9687,N_9891);
and U9988 (N_9988,N_9839,N_9784);
xnor U9989 (N_9989,N_9697,N_9867);
xor U9990 (N_9990,N_9624,N_9757);
nor U9991 (N_9991,N_9652,N_9756);
xnor U9992 (N_9992,N_9753,N_9628);
nand U9993 (N_9993,N_9899,N_9636);
or U9994 (N_9994,N_9662,N_9605);
and U9995 (N_9995,N_9879,N_9611);
nor U9996 (N_9996,N_9795,N_9861);
nor U9997 (N_9997,N_9811,N_9604);
or U9998 (N_9998,N_9862,N_9854);
xnor U9999 (N_9999,N_9630,N_9766);
and U10000 (N_10000,N_9865,N_9615);
and U10001 (N_10001,N_9681,N_9676);
and U10002 (N_10002,N_9761,N_9694);
nand U10003 (N_10003,N_9736,N_9855);
and U10004 (N_10004,N_9705,N_9794);
and U10005 (N_10005,N_9808,N_9768);
and U10006 (N_10006,N_9639,N_9851);
or U10007 (N_10007,N_9898,N_9644);
nor U10008 (N_10008,N_9843,N_9807);
nor U10009 (N_10009,N_9686,N_9602);
or U10010 (N_10010,N_9812,N_9721);
xnor U10011 (N_10011,N_9827,N_9790);
xnor U10012 (N_10012,N_9666,N_9660);
or U10013 (N_10013,N_9864,N_9785);
nor U10014 (N_10014,N_9603,N_9693);
and U10015 (N_10015,N_9800,N_9690);
nand U10016 (N_10016,N_9838,N_9763);
xor U10017 (N_10017,N_9828,N_9711);
nor U10018 (N_10018,N_9796,N_9719);
xnor U10019 (N_10019,N_9709,N_9777);
and U10020 (N_10020,N_9890,N_9713);
or U10021 (N_10021,N_9857,N_9835);
nor U10022 (N_10022,N_9813,N_9640);
nor U10023 (N_10023,N_9695,N_9661);
nand U10024 (N_10024,N_9643,N_9814);
nand U10025 (N_10025,N_9745,N_9678);
or U10026 (N_10026,N_9665,N_9842);
or U10027 (N_10027,N_9850,N_9654);
or U10028 (N_10028,N_9840,N_9699);
xnor U10029 (N_10029,N_9825,N_9779);
nand U10030 (N_10030,N_9866,N_9846);
and U10031 (N_10031,N_9674,N_9833);
or U10032 (N_10032,N_9712,N_9748);
xor U10033 (N_10033,N_9797,N_9884);
or U10034 (N_10034,N_9698,N_9617);
xor U10035 (N_10035,N_9610,N_9614);
nor U10036 (N_10036,N_9873,N_9841);
or U10037 (N_10037,N_9788,N_9883);
nand U10038 (N_10038,N_9619,N_9663);
nor U10039 (N_10039,N_9771,N_9658);
nor U10040 (N_10040,N_9770,N_9706);
and U10041 (N_10041,N_9876,N_9703);
and U10042 (N_10042,N_9618,N_9700);
or U10043 (N_10043,N_9635,N_9684);
xnor U10044 (N_10044,N_9836,N_9885);
xnor U10045 (N_10045,N_9792,N_9787);
or U10046 (N_10046,N_9798,N_9735);
nor U10047 (N_10047,N_9847,N_9781);
nor U10048 (N_10048,N_9688,N_9672);
and U10049 (N_10049,N_9724,N_9759);
nor U10050 (N_10050,N_9785,N_9631);
and U10051 (N_10051,N_9764,N_9610);
xor U10052 (N_10052,N_9729,N_9601);
xnor U10053 (N_10053,N_9851,N_9838);
nand U10054 (N_10054,N_9664,N_9640);
xnor U10055 (N_10055,N_9680,N_9737);
xnor U10056 (N_10056,N_9778,N_9641);
or U10057 (N_10057,N_9670,N_9614);
or U10058 (N_10058,N_9874,N_9889);
xnor U10059 (N_10059,N_9881,N_9886);
nand U10060 (N_10060,N_9609,N_9767);
xnor U10061 (N_10061,N_9784,N_9744);
and U10062 (N_10062,N_9826,N_9840);
nand U10063 (N_10063,N_9654,N_9771);
nor U10064 (N_10064,N_9861,N_9804);
nand U10065 (N_10065,N_9761,N_9745);
or U10066 (N_10066,N_9762,N_9649);
nand U10067 (N_10067,N_9765,N_9846);
nor U10068 (N_10068,N_9872,N_9827);
nand U10069 (N_10069,N_9785,N_9786);
nor U10070 (N_10070,N_9749,N_9725);
nor U10071 (N_10071,N_9600,N_9747);
nand U10072 (N_10072,N_9734,N_9670);
and U10073 (N_10073,N_9612,N_9640);
nor U10074 (N_10074,N_9813,N_9658);
nor U10075 (N_10075,N_9755,N_9678);
xnor U10076 (N_10076,N_9674,N_9849);
xor U10077 (N_10077,N_9788,N_9846);
nor U10078 (N_10078,N_9621,N_9788);
xor U10079 (N_10079,N_9638,N_9683);
and U10080 (N_10080,N_9729,N_9684);
nor U10081 (N_10081,N_9723,N_9785);
xnor U10082 (N_10082,N_9650,N_9888);
nand U10083 (N_10083,N_9809,N_9743);
or U10084 (N_10084,N_9874,N_9793);
nand U10085 (N_10085,N_9727,N_9638);
or U10086 (N_10086,N_9665,N_9687);
or U10087 (N_10087,N_9787,N_9837);
and U10088 (N_10088,N_9727,N_9797);
or U10089 (N_10089,N_9809,N_9765);
and U10090 (N_10090,N_9606,N_9677);
or U10091 (N_10091,N_9688,N_9731);
nand U10092 (N_10092,N_9693,N_9654);
and U10093 (N_10093,N_9884,N_9619);
xor U10094 (N_10094,N_9740,N_9682);
and U10095 (N_10095,N_9853,N_9897);
or U10096 (N_10096,N_9748,N_9607);
nand U10097 (N_10097,N_9704,N_9688);
or U10098 (N_10098,N_9889,N_9668);
and U10099 (N_10099,N_9796,N_9824);
nand U10100 (N_10100,N_9861,N_9712);
nand U10101 (N_10101,N_9669,N_9624);
xnor U10102 (N_10102,N_9768,N_9846);
xor U10103 (N_10103,N_9703,N_9648);
and U10104 (N_10104,N_9679,N_9607);
xnor U10105 (N_10105,N_9740,N_9749);
and U10106 (N_10106,N_9668,N_9809);
or U10107 (N_10107,N_9824,N_9668);
nand U10108 (N_10108,N_9750,N_9800);
nand U10109 (N_10109,N_9624,N_9738);
or U10110 (N_10110,N_9664,N_9711);
and U10111 (N_10111,N_9664,N_9771);
nand U10112 (N_10112,N_9620,N_9643);
or U10113 (N_10113,N_9753,N_9745);
and U10114 (N_10114,N_9861,N_9680);
and U10115 (N_10115,N_9680,N_9706);
nand U10116 (N_10116,N_9769,N_9720);
nand U10117 (N_10117,N_9867,N_9727);
or U10118 (N_10118,N_9678,N_9672);
nor U10119 (N_10119,N_9849,N_9817);
nor U10120 (N_10120,N_9737,N_9812);
or U10121 (N_10121,N_9822,N_9666);
nor U10122 (N_10122,N_9788,N_9881);
nor U10123 (N_10123,N_9684,N_9791);
and U10124 (N_10124,N_9699,N_9655);
nor U10125 (N_10125,N_9687,N_9624);
or U10126 (N_10126,N_9633,N_9634);
nor U10127 (N_10127,N_9612,N_9647);
nor U10128 (N_10128,N_9737,N_9631);
nand U10129 (N_10129,N_9650,N_9660);
nor U10130 (N_10130,N_9893,N_9695);
or U10131 (N_10131,N_9698,N_9896);
or U10132 (N_10132,N_9742,N_9832);
xor U10133 (N_10133,N_9766,N_9723);
xor U10134 (N_10134,N_9616,N_9822);
or U10135 (N_10135,N_9784,N_9687);
xnor U10136 (N_10136,N_9606,N_9660);
and U10137 (N_10137,N_9694,N_9671);
nand U10138 (N_10138,N_9619,N_9609);
and U10139 (N_10139,N_9750,N_9653);
nor U10140 (N_10140,N_9846,N_9878);
or U10141 (N_10141,N_9648,N_9705);
and U10142 (N_10142,N_9613,N_9851);
nand U10143 (N_10143,N_9764,N_9642);
nand U10144 (N_10144,N_9786,N_9709);
xnor U10145 (N_10145,N_9850,N_9885);
or U10146 (N_10146,N_9670,N_9629);
nor U10147 (N_10147,N_9721,N_9685);
nand U10148 (N_10148,N_9782,N_9813);
nand U10149 (N_10149,N_9612,N_9683);
or U10150 (N_10150,N_9740,N_9713);
or U10151 (N_10151,N_9660,N_9878);
nand U10152 (N_10152,N_9605,N_9637);
nor U10153 (N_10153,N_9604,N_9744);
or U10154 (N_10154,N_9767,N_9676);
nand U10155 (N_10155,N_9736,N_9614);
and U10156 (N_10156,N_9733,N_9793);
nand U10157 (N_10157,N_9721,N_9835);
nand U10158 (N_10158,N_9697,N_9692);
nor U10159 (N_10159,N_9793,N_9806);
or U10160 (N_10160,N_9825,N_9882);
and U10161 (N_10161,N_9879,N_9659);
or U10162 (N_10162,N_9675,N_9718);
or U10163 (N_10163,N_9767,N_9872);
or U10164 (N_10164,N_9785,N_9642);
or U10165 (N_10165,N_9807,N_9842);
and U10166 (N_10166,N_9785,N_9695);
xnor U10167 (N_10167,N_9685,N_9840);
or U10168 (N_10168,N_9885,N_9837);
xnor U10169 (N_10169,N_9612,N_9808);
nor U10170 (N_10170,N_9801,N_9765);
and U10171 (N_10171,N_9818,N_9860);
nor U10172 (N_10172,N_9687,N_9820);
nand U10173 (N_10173,N_9846,N_9725);
and U10174 (N_10174,N_9870,N_9890);
nor U10175 (N_10175,N_9875,N_9827);
xor U10176 (N_10176,N_9758,N_9847);
nand U10177 (N_10177,N_9813,N_9719);
xor U10178 (N_10178,N_9866,N_9701);
or U10179 (N_10179,N_9653,N_9600);
or U10180 (N_10180,N_9697,N_9853);
or U10181 (N_10181,N_9668,N_9848);
or U10182 (N_10182,N_9768,N_9831);
xor U10183 (N_10183,N_9838,N_9667);
or U10184 (N_10184,N_9726,N_9692);
nor U10185 (N_10185,N_9797,N_9753);
xnor U10186 (N_10186,N_9671,N_9736);
or U10187 (N_10187,N_9807,N_9850);
nor U10188 (N_10188,N_9738,N_9652);
and U10189 (N_10189,N_9884,N_9682);
or U10190 (N_10190,N_9695,N_9762);
and U10191 (N_10191,N_9884,N_9621);
and U10192 (N_10192,N_9784,N_9747);
and U10193 (N_10193,N_9799,N_9639);
nor U10194 (N_10194,N_9628,N_9897);
xor U10195 (N_10195,N_9792,N_9817);
nor U10196 (N_10196,N_9613,N_9703);
nor U10197 (N_10197,N_9635,N_9899);
or U10198 (N_10198,N_9834,N_9634);
nand U10199 (N_10199,N_9725,N_9624);
xor U10200 (N_10200,N_10109,N_9940);
and U10201 (N_10201,N_10060,N_9966);
or U10202 (N_10202,N_10020,N_9965);
nand U10203 (N_10203,N_10038,N_10129);
nor U10204 (N_10204,N_10193,N_10098);
nand U10205 (N_10205,N_10077,N_9971);
nor U10206 (N_10206,N_10127,N_10057);
xor U10207 (N_10207,N_10171,N_9923);
or U10208 (N_10208,N_10143,N_10004);
xor U10209 (N_10209,N_10067,N_9949);
or U10210 (N_10210,N_9911,N_10173);
nor U10211 (N_10211,N_9972,N_9989);
nand U10212 (N_10212,N_10022,N_9948);
or U10213 (N_10213,N_10012,N_10006);
and U10214 (N_10214,N_9995,N_10072);
nand U10215 (N_10215,N_10187,N_9950);
or U10216 (N_10216,N_10030,N_10066);
nor U10217 (N_10217,N_10011,N_10157);
xnor U10218 (N_10218,N_10176,N_10005);
nor U10219 (N_10219,N_10100,N_9922);
nand U10220 (N_10220,N_9918,N_9928);
or U10221 (N_10221,N_10055,N_10002);
or U10222 (N_10222,N_9954,N_10069);
nor U10223 (N_10223,N_9976,N_9946);
or U10224 (N_10224,N_10045,N_10120);
and U10225 (N_10225,N_10059,N_10039);
nand U10226 (N_10226,N_10191,N_10138);
nor U10227 (N_10227,N_10140,N_9904);
nor U10228 (N_10228,N_10037,N_10051);
nor U10229 (N_10229,N_9991,N_10056);
nand U10230 (N_10230,N_9981,N_9975);
and U10231 (N_10231,N_10093,N_10048);
nand U10232 (N_10232,N_10184,N_10085);
nor U10233 (N_10233,N_9934,N_10159);
or U10234 (N_10234,N_10008,N_10145);
nor U10235 (N_10235,N_10024,N_9993);
nand U10236 (N_10236,N_10076,N_9912);
and U10237 (N_10237,N_10174,N_9900);
nand U10238 (N_10238,N_9947,N_9969);
nand U10239 (N_10239,N_9935,N_10155);
nor U10240 (N_10240,N_10121,N_10168);
nor U10241 (N_10241,N_9951,N_10035);
nand U10242 (N_10242,N_10156,N_10130);
nor U10243 (N_10243,N_9945,N_10108);
and U10244 (N_10244,N_9978,N_9970);
xor U10245 (N_10245,N_9973,N_9987);
nor U10246 (N_10246,N_9983,N_10190);
or U10247 (N_10247,N_10040,N_10009);
or U10248 (N_10248,N_10046,N_10199);
xnor U10249 (N_10249,N_9903,N_10000);
and U10250 (N_10250,N_9936,N_9913);
and U10251 (N_10251,N_10158,N_10122);
and U10252 (N_10252,N_10189,N_10131);
or U10253 (N_10253,N_10153,N_10135);
nand U10254 (N_10254,N_9957,N_10170);
or U10255 (N_10255,N_10142,N_10188);
and U10256 (N_10256,N_10194,N_9941);
xor U10257 (N_10257,N_10021,N_10034);
nand U10258 (N_10258,N_10062,N_10179);
and U10259 (N_10259,N_10061,N_10063);
xor U10260 (N_10260,N_10036,N_10095);
or U10261 (N_10261,N_9917,N_10103);
or U10262 (N_10262,N_10115,N_9927);
nor U10263 (N_10263,N_10125,N_10075);
and U10264 (N_10264,N_10086,N_9906);
and U10265 (N_10265,N_10087,N_10016);
and U10266 (N_10266,N_10041,N_9932);
nor U10267 (N_10267,N_10118,N_9980);
nand U10268 (N_10268,N_10096,N_10148);
and U10269 (N_10269,N_10003,N_9990);
nand U10270 (N_10270,N_10042,N_10132);
nand U10271 (N_10271,N_9999,N_9974);
nand U10272 (N_10272,N_9907,N_9943);
nor U10273 (N_10273,N_10113,N_10097);
and U10274 (N_10274,N_10044,N_9988);
nand U10275 (N_10275,N_10149,N_10074);
or U10276 (N_10276,N_10106,N_10169);
xnor U10277 (N_10277,N_10198,N_10026);
and U10278 (N_10278,N_10081,N_9920);
nor U10279 (N_10279,N_9901,N_9924);
nor U10280 (N_10280,N_9929,N_10114);
or U10281 (N_10281,N_9908,N_10028);
or U10282 (N_10282,N_10141,N_10017);
nor U10283 (N_10283,N_10082,N_10025);
or U10284 (N_10284,N_10110,N_10018);
nand U10285 (N_10285,N_10101,N_10134);
nor U10286 (N_10286,N_9956,N_10105);
and U10287 (N_10287,N_10137,N_10154);
or U10288 (N_10288,N_10123,N_10071);
nand U10289 (N_10289,N_9919,N_10073);
nor U10290 (N_10290,N_10172,N_9905);
nand U10291 (N_10291,N_10197,N_10107);
xnor U10292 (N_10292,N_9942,N_10104);
nor U10293 (N_10293,N_10052,N_9992);
xnor U10294 (N_10294,N_9984,N_9964);
or U10295 (N_10295,N_10080,N_10050);
or U10296 (N_10296,N_9921,N_10124);
or U10297 (N_10297,N_10180,N_10068);
xor U10298 (N_10298,N_10058,N_9925);
or U10299 (N_10299,N_10083,N_10007);
nor U10300 (N_10300,N_10013,N_10043);
nor U10301 (N_10301,N_9982,N_10182);
xnor U10302 (N_10302,N_10031,N_10139);
nor U10303 (N_10303,N_10112,N_10160);
and U10304 (N_10304,N_10054,N_10094);
nor U10305 (N_10305,N_9955,N_9931);
nand U10306 (N_10306,N_9997,N_9977);
nand U10307 (N_10307,N_10053,N_10163);
xnor U10308 (N_10308,N_9959,N_10049);
nand U10309 (N_10309,N_10078,N_9960);
nand U10310 (N_10310,N_10161,N_10047);
nand U10311 (N_10311,N_9968,N_10102);
and U10312 (N_10312,N_9914,N_10165);
xnor U10313 (N_10313,N_10032,N_10164);
nor U10314 (N_10314,N_10175,N_10178);
xnor U10315 (N_10315,N_10177,N_9996);
xnor U10316 (N_10316,N_10001,N_10167);
nor U10317 (N_10317,N_10019,N_9985);
and U10318 (N_10318,N_10091,N_10183);
nand U10319 (N_10319,N_10027,N_10150);
and U10320 (N_10320,N_9962,N_9986);
or U10321 (N_10321,N_10133,N_9926);
xnor U10322 (N_10322,N_10084,N_10152);
nor U10323 (N_10323,N_9910,N_10128);
xnor U10324 (N_10324,N_10151,N_10014);
and U10325 (N_10325,N_9958,N_10092);
xor U10326 (N_10326,N_10136,N_9916);
or U10327 (N_10327,N_9967,N_10015);
xnor U10328 (N_10328,N_9933,N_9952);
nand U10329 (N_10329,N_10166,N_10010);
nor U10330 (N_10330,N_10146,N_10079);
and U10331 (N_10331,N_10196,N_9909);
xor U10332 (N_10332,N_9939,N_10029);
xnor U10333 (N_10333,N_10192,N_10090);
or U10334 (N_10334,N_9938,N_10070);
or U10335 (N_10335,N_10144,N_9994);
xor U10336 (N_10336,N_10147,N_10064);
and U10337 (N_10337,N_9953,N_10065);
xnor U10338 (N_10338,N_9930,N_10111);
and U10339 (N_10339,N_10119,N_10186);
nand U10340 (N_10340,N_9915,N_10088);
or U10341 (N_10341,N_10023,N_10126);
nor U10342 (N_10342,N_9998,N_10089);
xor U10343 (N_10343,N_9961,N_10099);
and U10344 (N_10344,N_10117,N_10185);
and U10345 (N_10345,N_10116,N_9937);
and U10346 (N_10346,N_9979,N_10181);
and U10347 (N_10347,N_10033,N_9944);
or U10348 (N_10348,N_9902,N_10162);
nor U10349 (N_10349,N_10195,N_9963);
nand U10350 (N_10350,N_9957,N_10163);
nor U10351 (N_10351,N_10158,N_9968);
nor U10352 (N_10352,N_10167,N_10143);
or U10353 (N_10353,N_10032,N_9978);
nand U10354 (N_10354,N_10091,N_9937);
nand U10355 (N_10355,N_10114,N_10084);
or U10356 (N_10356,N_10013,N_10042);
xor U10357 (N_10357,N_10017,N_9900);
or U10358 (N_10358,N_10048,N_9923);
or U10359 (N_10359,N_9948,N_10088);
nand U10360 (N_10360,N_10102,N_9917);
xor U10361 (N_10361,N_9990,N_9944);
or U10362 (N_10362,N_10053,N_10044);
nor U10363 (N_10363,N_9991,N_10118);
xor U10364 (N_10364,N_10199,N_10107);
and U10365 (N_10365,N_9939,N_10175);
or U10366 (N_10366,N_9929,N_10067);
nor U10367 (N_10367,N_9986,N_10052);
or U10368 (N_10368,N_9924,N_10114);
nand U10369 (N_10369,N_10006,N_9909);
or U10370 (N_10370,N_10100,N_10042);
nor U10371 (N_10371,N_10194,N_10042);
nand U10372 (N_10372,N_10074,N_10055);
nand U10373 (N_10373,N_9950,N_9953);
and U10374 (N_10374,N_10152,N_9991);
or U10375 (N_10375,N_10079,N_9931);
nand U10376 (N_10376,N_10157,N_10068);
xor U10377 (N_10377,N_9954,N_9913);
xor U10378 (N_10378,N_10010,N_10093);
nor U10379 (N_10379,N_10012,N_10185);
xnor U10380 (N_10380,N_9997,N_9900);
or U10381 (N_10381,N_9934,N_10001);
xor U10382 (N_10382,N_10055,N_9997);
nand U10383 (N_10383,N_10010,N_10059);
and U10384 (N_10384,N_9924,N_10165);
nand U10385 (N_10385,N_10144,N_9934);
xnor U10386 (N_10386,N_10173,N_10165);
nand U10387 (N_10387,N_9969,N_10043);
or U10388 (N_10388,N_10030,N_10180);
nor U10389 (N_10389,N_10123,N_10119);
nand U10390 (N_10390,N_9958,N_9962);
xor U10391 (N_10391,N_10083,N_10039);
xnor U10392 (N_10392,N_9947,N_10152);
nand U10393 (N_10393,N_10021,N_10074);
and U10394 (N_10394,N_9962,N_9981);
nor U10395 (N_10395,N_9930,N_9901);
nand U10396 (N_10396,N_10016,N_10176);
nand U10397 (N_10397,N_10059,N_10168);
nor U10398 (N_10398,N_10173,N_10090);
nand U10399 (N_10399,N_10173,N_9958);
nand U10400 (N_10400,N_10071,N_10128);
nor U10401 (N_10401,N_10192,N_9989);
nand U10402 (N_10402,N_10112,N_9926);
nand U10403 (N_10403,N_9901,N_10102);
nand U10404 (N_10404,N_10185,N_10162);
or U10405 (N_10405,N_9959,N_10058);
or U10406 (N_10406,N_9995,N_10165);
xor U10407 (N_10407,N_9978,N_10116);
nor U10408 (N_10408,N_10161,N_10077);
nand U10409 (N_10409,N_10095,N_10035);
nor U10410 (N_10410,N_9974,N_10049);
xnor U10411 (N_10411,N_9928,N_9947);
and U10412 (N_10412,N_10002,N_9902);
and U10413 (N_10413,N_10193,N_10031);
and U10414 (N_10414,N_9994,N_10023);
xnor U10415 (N_10415,N_10041,N_10029);
xor U10416 (N_10416,N_9971,N_10181);
or U10417 (N_10417,N_10184,N_9966);
and U10418 (N_10418,N_9920,N_10164);
and U10419 (N_10419,N_10145,N_10104);
and U10420 (N_10420,N_10139,N_9972);
or U10421 (N_10421,N_10168,N_10071);
nor U10422 (N_10422,N_9933,N_9983);
nor U10423 (N_10423,N_9978,N_10093);
and U10424 (N_10424,N_10193,N_10053);
and U10425 (N_10425,N_10176,N_10127);
nor U10426 (N_10426,N_10079,N_9960);
or U10427 (N_10427,N_10043,N_9919);
and U10428 (N_10428,N_10115,N_10026);
nand U10429 (N_10429,N_10146,N_10093);
or U10430 (N_10430,N_10077,N_9956);
or U10431 (N_10431,N_9906,N_10129);
or U10432 (N_10432,N_10100,N_9915);
nand U10433 (N_10433,N_10136,N_9930);
or U10434 (N_10434,N_9934,N_9951);
and U10435 (N_10435,N_10010,N_9997);
or U10436 (N_10436,N_10159,N_10118);
or U10437 (N_10437,N_10002,N_9978);
or U10438 (N_10438,N_10144,N_9979);
or U10439 (N_10439,N_10107,N_10039);
or U10440 (N_10440,N_10147,N_9928);
and U10441 (N_10441,N_9976,N_10076);
nand U10442 (N_10442,N_10131,N_10057);
or U10443 (N_10443,N_10164,N_10051);
and U10444 (N_10444,N_9986,N_9912);
nand U10445 (N_10445,N_10067,N_10082);
and U10446 (N_10446,N_10143,N_10180);
or U10447 (N_10447,N_9901,N_9908);
xor U10448 (N_10448,N_10155,N_10115);
or U10449 (N_10449,N_9966,N_10056);
nor U10450 (N_10450,N_10018,N_9997);
nand U10451 (N_10451,N_10069,N_10071);
nor U10452 (N_10452,N_9984,N_10052);
or U10453 (N_10453,N_9957,N_10041);
or U10454 (N_10454,N_10130,N_9935);
nand U10455 (N_10455,N_10075,N_9912);
nand U10456 (N_10456,N_10002,N_9984);
and U10457 (N_10457,N_9912,N_10159);
nand U10458 (N_10458,N_10182,N_10179);
xnor U10459 (N_10459,N_9903,N_10156);
xor U10460 (N_10460,N_10047,N_10173);
nand U10461 (N_10461,N_9990,N_10110);
nor U10462 (N_10462,N_9963,N_10183);
nor U10463 (N_10463,N_10179,N_10082);
xnor U10464 (N_10464,N_10175,N_9965);
and U10465 (N_10465,N_10046,N_9966);
nand U10466 (N_10466,N_10056,N_10046);
or U10467 (N_10467,N_10018,N_10126);
nor U10468 (N_10468,N_10104,N_10099);
nand U10469 (N_10469,N_10002,N_9986);
or U10470 (N_10470,N_10179,N_10148);
or U10471 (N_10471,N_10016,N_9956);
nor U10472 (N_10472,N_9931,N_9926);
and U10473 (N_10473,N_9936,N_10043);
xnor U10474 (N_10474,N_10190,N_9906);
and U10475 (N_10475,N_9938,N_10156);
xnor U10476 (N_10476,N_9940,N_10078);
and U10477 (N_10477,N_9901,N_10105);
xor U10478 (N_10478,N_10123,N_10177);
nor U10479 (N_10479,N_10192,N_10046);
and U10480 (N_10480,N_9943,N_10147);
xnor U10481 (N_10481,N_10139,N_9951);
nand U10482 (N_10482,N_10172,N_9971);
nand U10483 (N_10483,N_9981,N_9996);
and U10484 (N_10484,N_10054,N_10152);
and U10485 (N_10485,N_10004,N_9967);
nand U10486 (N_10486,N_9980,N_9913);
xor U10487 (N_10487,N_10101,N_10168);
or U10488 (N_10488,N_10194,N_10025);
xor U10489 (N_10489,N_10077,N_10012);
or U10490 (N_10490,N_10032,N_10105);
nand U10491 (N_10491,N_10175,N_10027);
and U10492 (N_10492,N_10025,N_9930);
nor U10493 (N_10493,N_9909,N_10088);
nand U10494 (N_10494,N_10103,N_10063);
nor U10495 (N_10495,N_10052,N_9991);
nor U10496 (N_10496,N_9930,N_10163);
xor U10497 (N_10497,N_9964,N_9900);
xnor U10498 (N_10498,N_10114,N_9977);
or U10499 (N_10499,N_10013,N_10064);
xnor U10500 (N_10500,N_10238,N_10374);
or U10501 (N_10501,N_10499,N_10360);
or U10502 (N_10502,N_10477,N_10312);
or U10503 (N_10503,N_10316,N_10419);
or U10504 (N_10504,N_10211,N_10420);
nor U10505 (N_10505,N_10288,N_10320);
nor U10506 (N_10506,N_10247,N_10232);
and U10507 (N_10507,N_10381,N_10457);
nor U10508 (N_10508,N_10239,N_10336);
nor U10509 (N_10509,N_10251,N_10344);
xnor U10510 (N_10510,N_10350,N_10340);
xor U10511 (N_10511,N_10482,N_10405);
and U10512 (N_10512,N_10400,N_10302);
nor U10513 (N_10513,N_10416,N_10326);
xor U10514 (N_10514,N_10235,N_10276);
and U10515 (N_10515,N_10286,N_10334);
xor U10516 (N_10516,N_10339,N_10496);
xnor U10517 (N_10517,N_10364,N_10266);
or U10518 (N_10518,N_10230,N_10231);
nand U10519 (N_10519,N_10281,N_10367);
xnor U10520 (N_10520,N_10476,N_10462);
nand U10521 (N_10521,N_10327,N_10332);
xnor U10522 (N_10522,N_10423,N_10269);
and U10523 (N_10523,N_10427,N_10282);
and U10524 (N_10524,N_10328,N_10324);
nand U10525 (N_10525,N_10395,N_10446);
nor U10526 (N_10526,N_10305,N_10439);
xor U10527 (N_10527,N_10268,N_10382);
xor U10528 (N_10528,N_10293,N_10438);
or U10529 (N_10529,N_10223,N_10410);
and U10530 (N_10530,N_10489,N_10347);
or U10531 (N_10531,N_10474,N_10204);
xor U10532 (N_10532,N_10297,N_10253);
or U10533 (N_10533,N_10484,N_10299);
nor U10534 (N_10534,N_10463,N_10319);
or U10535 (N_10535,N_10404,N_10338);
nor U10536 (N_10536,N_10263,N_10387);
xnor U10537 (N_10537,N_10373,N_10418);
nand U10538 (N_10538,N_10412,N_10244);
nand U10539 (N_10539,N_10274,N_10415);
and U10540 (N_10540,N_10435,N_10362);
and U10541 (N_10541,N_10468,N_10424);
or U10542 (N_10542,N_10478,N_10240);
xor U10543 (N_10543,N_10358,N_10466);
nor U10544 (N_10544,N_10426,N_10366);
xor U10545 (N_10545,N_10242,N_10330);
nor U10546 (N_10546,N_10498,N_10413);
nand U10547 (N_10547,N_10308,N_10451);
nand U10548 (N_10548,N_10385,N_10214);
nor U10549 (N_10549,N_10252,N_10406);
or U10550 (N_10550,N_10434,N_10351);
or U10551 (N_10551,N_10490,N_10272);
nor U10552 (N_10552,N_10264,N_10453);
nor U10553 (N_10553,N_10398,N_10261);
nand U10554 (N_10554,N_10256,N_10488);
or U10555 (N_10555,N_10225,N_10245);
and U10556 (N_10556,N_10445,N_10201);
and U10557 (N_10557,N_10295,N_10206);
nor U10558 (N_10558,N_10375,N_10459);
or U10559 (N_10559,N_10409,N_10356);
nor U10560 (N_10560,N_10296,N_10370);
xnor U10561 (N_10561,N_10255,N_10321);
and U10562 (N_10562,N_10310,N_10289);
nand U10563 (N_10563,N_10383,N_10421);
and U10564 (N_10564,N_10294,N_10487);
nor U10565 (N_10565,N_10265,N_10202);
and U10566 (N_10566,N_10307,N_10250);
xnor U10567 (N_10567,N_10229,N_10280);
and U10568 (N_10568,N_10443,N_10391);
nand U10569 (N_10569,N_10470,N_10254);
or U10570 (N_10570,N_10411,N_10436);
nand U10571 (N_10571,N_10393,N_10472);
nor U10572 (N_10572,N_10348,N_10432);
nor U10573 (N_10573,N_10376,N_10311);
or U10574 (N_10574,N_10292,N_10323);
nand U10575 (N_10575,N_10301,N_10368);
nand U10576 (N_10576,N_10273,N_10441);
nor U10577 (N_10577,N_10258,N_10361);
nand U10578 (N_10578,N_10303,N_10341);
xor U10579 (N_10579,N_10497,N_10236);
and U10580 (N_10580,N_10473,N_10493);
and U10581 (N_10581,N_10318,N_10315);
and U10582 (N_10582,N_10218,N_10259);
nor U10583 (N_10583,N_10335,N_10458);
and U10584 (N_10584,N_10414,N_10207);
nand U10585 (N_10585,N_10352,N_10283);
nand U10586 (N_10586,N_10212,N_10392);
or U10587 (N_10587,N_10452,N_10461);
nand U10588 (N_10588,N_10379,N_10467);
or U10589 (N_10589,N_10278,N_10216);
nand U10590 (N_10590,N_10249,N_10275);
nor U10591 (N_10591,N_10354,N_10353);
or U10592 (N_10592,N_10454,N_10215);
nand U10593 (N_10593,N_10329,N_10433);
or U10594 (N_10594,N_10456,N_10304);
nor U10595 (N_10595,N_10349,N_10396);
nor U10596 (N_10596,N_10343,N_10217);
nand U10597 (N_10597,N_10380,N_10408);
and U10598 (N_10598,N_10460,N_10495);
and U10599 (N_10599,N_10437,N_10429);
xnor U10600 (N_10600,N_10222,N_10425);
or U10601 (N_10601,N_10449,N_10442);
or U10602 (N_10602,N_10345,N_10399);
and U10603 (N_10603,N_10270,N_10260);
nand U10604 (N_10604,N_10221,N_10233);
nor U10605 (N_10605,N_10300,N_10226);
nand U10606 (N_10606,N_10492,N_10219);
or U10607 (N_10607,N_10479,N_10203);
nor U10608 (N_10608,N_10234,N_10298);
nor U10609 (N_10609,N_10390,N_10448);
xnor U10610 (N_10610,N_10333,N_10237);
nand U10611 (N_10611,N_10363,N_10402);
or U10612 (N_10612,N_10365,N_10209);
and U10613 (N_10613,N_10309,N_10314);
xnor U10614 (N_10614,N_10450,N_10371);
nor U10615 (N_10615,N_10359,N_10322);
nand U10616 (N_10616,N_10485,N_10243);
nand U10617 (N_10617,N_10213,N_10291);
or U10618 (N_10618,N_10306,N_10417);
or U10619 (N_10619,N_10471,N_10494);
and U10620 (N_10620,N_10208,N_10369);
nand U10621 (N_10621,N_10200,N_10357);
nand U10622 (N_10622,N_10285,N_10355);
nand U10623 (N_10623,N_10224,N_10469);
nand U10624 (N_10624,N_10388,N_10257);
xor U10625 (N_10625,N_10475,N_10455);
and U10626 (N_10626,N_10389,N_10220);
xor U10627 (N_10627,N_10271,N_10447);
and U10628 (N_10628,N_10210,N_10480);
nor U10629 (N_10629,N_10284,N_10325);
and U10630 (N_10630,N_10262,N_10267);
nand U10631 (N_10631,N_10384,N_10279);
and U10632 (N_10632,N_10313,N_10486);
or U10633 (N_10633,N_10403,N_10422);
nor U10634 (N_10634,N_10464,N_10378);
nand U10635 (N_10635,N_10491,N_10337);
nor U10636 (N_10636,N_10372,N_10428);
or U10637 (N_10637,N_10444,N_10481);
nand U10638 (N_10638,N_10431,N_10290);
nor U10639 (N_10639,N_10248,N_10407);
and U10640 (N_10640,N_10205,N_10287);
and U10641 (N_10641,N_10430,N_10397);
or U10642 (N_10642,N_10277,N_10317);
nor U10643 (N_10643,N_10394,N_10401);
and U10644 (N_10644,N_10377,N_10440);
or U10645 (N_10645,N_10246,N_10331);
or U10646 (N_10646,N_10465,N_10228);
and U10647 (N_10647,N_10346,N_10342);
nand U10648 (N_10648,N_10386,N_10483);
or U10649 (N_10649,N_10227,N_10241);
or U10650 (N_10650,N_10206,N_10416);
xor U10651 (N_10651,N_10472,N_10490);
nand U10652 (N_10652,N_10458,N_10348);
and U10653 (N_10653,N_10465,N_10455);
nand U10654 (N_10654,N_10461,N_10350);
nor U10655 (N_10655,N_10220,N_10471);
and U10656 (N_10656,N_10363,N_10420);
or U10657 (N_10657,N_10439,N_10302);
and U10658 (N_10658,N_10427,N_10220);
xor U10659 (N_10659,N_10496,N_10377);
xor U10660 (N_10660,N_10309,N_10282);
and U10661 (N_10661,N_10381,N_10209);
nand U10662 (N_10662,N_10233,N_10223);
or U10663 (N_10663,N_10321,N_10203);
nand U10664 (N_10664,N_10291,N_10330);
nor U10665 (N_10665,N_10221,N_10491);
xor U10666 (N_10666,N_10480,N_10290);
and U10667 (N_10667,N_10293,N_10365);
nand U10668 (N_10668,N_10385,N_10470);
nand U10669 (N_10669,N_10446,N_10347);
nor U10670 (N_10670,N_10245,N_10356);
nand U10671 (N_10671,N_10375,N_10330);
nand U10672 (N_10672,N_10304,N_10290);
or U10673 (N_10673,N_10472,N_10338);
nand U10674 (N_10674,N_10491,N_10378);
nand U10675 (N_10675,N_10440,N_10347);
nand U10676 (N_10676,N_10468,N_10361);
nor U10677 (N_10677,N_10498,N_10379);
or U10678 (N_10678,N_10328,N_10435);
nand U10679 (N_10679,N_10360,N_10327);
nor U10680 (N_10680,N_10309,N_10463);
nor U10681 (N_10681,N_10216,N_10326);
nand U10682 (N_10682,N_10248,N_10356);
nand U10683 (N_10683,N_10487,N_10389);
and U10684 (N_10684,N_10239,N_10497);
xor U10685 (N_10685,N_10475,N_10391);
nor U10686 (N_10686,N_10463,N_10248);
nor U10687 (N_10687,N_10411,N_10443);
or U10688 (N_10688,N_10495,N_10298);
xor U10689 (N_10689,N_10376,N_10398);
or U10690 (N_10690,N_10422,N_10454);
and U10691 (N_10691,N_10261,N_10246);
nor U10692 (N_10692,N_10253,N_10290);
or U10693 (N_10693,N_10315,N_10249);
nand U10694 (N_10694,N_10201,N_10312);
nor U10695 (N_10695,N_10354,N_10473);
xor U10696 (N_10696,N_10476,N_10437);
xnor U10697 (N_10697,N_10430,N_10485);
xnor U10698 (N_10698,N_10335,N_10492);
xor U10699 (N_10699,N_10403,N_10262);
or U10700 (N_10700,N_10202,N_10207);
nand U10701 (N_10701,N_10275,N_10262);
and U10702 (N_10702,N_10371,N_10282);
xor U10703 (N_10703,N_10451,N_10379);
nor U10704 (N_10704,N_10468,N_10340);
and U10705 (N_10705,N_10244,N_10239);
and U10706 (N_10706,N_10217,N_10335);
xnor U10707 (N_10707,N_10468,N_10242);
xor U10708 (N_10708,N_10372,N_10285);
or U10709 (N_10709,N_10345,N_10475);
xnor U10710 (N_10710,N_10299,N_10218);
nor U10711 (N_10711,N_10314,N_10444);
or U10712 (N_10712,N_10243,N_10313);
and U10713 (N_10713,N_10253,N_10220);
or U10714 (N_10714,N_10483,N_10412);
nand U10715 (N_10715,N_10460,N_10434);
nand U10716 (N_10716,N_10302,N_10419);
and U10717 (N_10717,N_10394,N_10456);
nor U10718 (N_10718,N_10371,N_10243);
nor U10719 (N_10719,N_10377,N_10439);
xor U10720 (N_10720,N_10417,N_10241);
nand U10721 (N_10721,N_10256,N_10330);
nor U10722 (N_10722,N_10267,N_10280);
or U10723 (N_10723,N_10209,N_10256);
nor U10724 (N_10724,N_10485,N_10264);
nand U10725 (N_10725,N_10387,N_10462);
nand U10726 (N_10726,N_10361,N_10423);
or U10727 (N_10727,N_10376,N_10342);
nand U10728 (N_10728,N_10326,N_10274);
nor U10729 (N_10729,N_10404,N_10314);
and U10730 (N_10730,N_10369,N_10243);
nor U10731 (N_10731,N_10379,N_10424);
nand U10732 (N_10732,N_10254,N_10458);
and U10733 (N_10733,N_10487,N_10440);
and U10734 (N_10734,N_10354,N_10294);
nor U10735 (N_10735,N_10324,N_10388);
nor U10736 (N_10736,N_10310,N_10319);
xor U10737 (N_10737,N_10201,N_10326);
nand U10738 (N_10738,N_10256,N_10451);
or U10739 (N_10739,N_10219,N_10216);
and U10740 (N_10740,N_10276,N_10425);
nor U10741 (N_10741,N_10363,N_10322);
and U10742 (N_10742,N_10496,N_10220);
nor U10743 (N_10743,N_10326,N_10419);
nor U10744 (N_10744,N_10303,N_10309);
xnor U10745 (N_10745,N_10288,N_10417);
nand U10746 (N_10746,N_10274,N_10418);
nor U10747 (N_10747,N_10306,N_10412);
or U10748 (N_10748,N_10460,N_10262);
nor U10749 (N_10749,N_10203,N_10410);
and U10750 (N_10750,N_10333,N_10480);
nand U10751 (N_10751,N_10339,N_10334);
xor U10752 (N_10752,N_10331,N_10452);
xor U10753 (N_10753,N_10453,N_10281);
nor U10754 (N_10754,N_10335,N_10433);
or U10755 (N_10755,N_10477,N_10311);
nand U10756 (N_10756,N_10418,N_10309);
nor U10757 (N_10757,N_10292,N_10253);
xnor U10758 (N_10758,N_10298,N_10271);
or U10759 (N_10759,N_10300,N_10295);
xor U10760 (N_10760,N_10221,N_10227);
nor U10761 (N_10761,N_10359,N_10354);
or U10762 (N_10762,N_10397,N_10499);
nand U10763 (N_10763,N_10452,N_10426);
xor U10764 (N_10764,N_10279,N_10401);
nor U10765 (N_10765,N_10389,N_10413);
and U10766 (N_10766,N_10236,N_10446);
or U10767 (N_10767,N_10462,N_10389);
nand U10768 (N_10768,N_10388,N_10372);
and U10769 (N_10769,N_10394,N_10300);
and U10770 (N_10770,N_10211,N_10353);
xor U10771 (N_10771,N_10444,N_10320);
xnor U10772 (N_10772,N_10353,N_10242);
and U10773 (N_10773,N_10200,N_10283);
nand U10774 (N_10774,N_10311,N_10439);
nor U10775 (N_10775,N_10409,N_10327);
nor U10776 (N_10776,N_10347,N_10245);
or U10777 (N_10777,N_10283,N_10343);
and U10778 (N_10778,N_10297,N_10301);
and U10779 (N_10779,N_10227,N_10312);
xor U10780 (N_10780,N_10236,N_10476);
xnor U10781 (N_10781,N_10261,N_10339);
nand U10782 (N_10782,N_10486,N_10260);
nand U10783 (N_10783,N_10312,N_10275);
nor U10784 (N_10784,N_10241,N_10254);
nor U10785 (N_10785,N_10420,N_10494);
or U10786 (N_10786,N_10290,N_10364);
nand U10787 (N_10787,N_10387,N_10358);
xor U10788 (N_10788,N_10263,N_10312);
and U10789 (N_10789,N_10496,N_10211);
nor U10790 (N_10790,N_10478,N_10329);
xnor U10791 (N_10791,N_10349,N_10449);
and U10792 (N_10792,N_10306,N_10456);
and U10793 (N_10793,N_10295,N_10455);
nand U10794 (N_10794,N_10482,N_10428);
xnor U10795 (N_10795,N_10373,N_10348);
nor U10796 (N_10796,N_10332,N_10454);
nand U10797 (N_10797,N_10447,N_10421);
and U10798 (N_10798,N_10265,N_10282);
nor U10799 (N_10799,N_10318,N_10420);
nor U10800 (N_10800,N_10556,N_10788);
xor U10801 (N_10801,N_10750,N_10647);
xnor U10802 (N_10802,N_10623,N_10607);
or U10803 (N_10803,N_10586,N_10536);
nand U10804 (N_10804,N_10729,N_10567);
xor U10805 (N_10805,N_10662,N_10694);
or U10806 (N_10806,N_10686,N_10568);
xnor U10807 (N_10807,N_10786,N_10504);
nor U10808 (N_10808,N_10538,N_10722);
nor U10809 (N_10809,N_10582,N_10798);
nand U10810 (N_10810,N_10508,N_10572);
nand U10811 (N_10811,N_10604,N_10770);
and U10812 (N_10812,N_10502,N_10551);
or U10813 (N_10813,N_10636,N_10558);
xnor U10814 (N_10814,N_10571,N_10783);
nor U10815 (N_10815,N_10544,N_10775);
nand U10816 (N_10816,N_10642,N_10796);
nand U10817 (N_10817,N_10673,N_10619);
xor U10818 (N_10818,N_10717,N_10580);
and U10819 (N_10819,N_10660,N_10697);
nor U10820 (N_10820,N_10659,N_10521);
and U10821 (N_10821,N_10579,N_10577);
and U10822 (N_10822,N_10707,N_10670);
or U10823 (N_10823,N_10738,N_10599);
or U10824 (N_10824,N_10581,N_10736);
xnor U10825 (N_10825,N_10528,N_10732);
xnor U10826 (N_10826,N_10737,N_10693);
xor U10827 (N_10827,N_10573,N_10741);
nand U10828 (N_10828,N_10688,N_10759);
nor U10829 (N_10829,N_10704,N_10757);
or U10830 (N_10830,N_10630,N_10758);
and U10831 (N_10831,N_10540,N_10709);
xor U10832 (N_10832,N_10598,N_10681);
nand U10833 (N_10833,N_10641,N_10531);
nand U10834 (N_10834,N_10525,N_10595);
xor U10835 (N_10835,N_10596,N_10637);
xor U10836 (N_10836,N_10516,N_10601);
nor U10837 (N_10837,N_10629,N_10679);
and U10838 (N_10838,N_10734,N_10554);
or U10839 (N_10839,N_10773,N_10767);
xnor U10840 (N_10840,N_10651,N_10576);
nor U10841 (N_10841,N_10588,N_10663);
and U10842 (N_10842,N_10726,N_10523);
xnor U10843 (N_10843,N_10534,N_10746);
and U10844 (N_10844,N_10511,N_10677);
xor U10845 (N_10845,N_10570,N_10515);
xor U10846 (N_10846,N_10763,N_10638);
and U10847 (N_10847,N_10622,N_10626);
or U10848 (N_10848,N_10761,N_10618);
xor U10849 (N_10849,N_10644,N_10505);
and U10850 (N_10850,N_10631,N_10735);
or U10851 (N_10851,N_10676,N_10678);
xnor U10852 (N_10852,N_10780,N_10587);
and U10853 (N_10853,N_10716,N_10503);
nor U10854 (N_10854,N_10683,N_10699);
or U10855 (N_10855,N_10777,N_10654);
and U10856 (N_10856,N_10698,N_10616);
nor U10857 (N_10857,N_10721,N_10774);
and U10858 (N_10858,N_10633,N_10723);
and U10859 (N_10859,N_10743,N_10564);
nor U10860 (N_10860,N_10539,N_10550);
nand U10861 (N_10861,N_10532,N_10522);
nor U10862 (N_10862,N_10615,N_10546);
nand U10863 (N_10863,N_10712,N_10575);
nor U10864 (N_10864,N_10684,N_10744);
xnor U10865 (N_10865,N_10537,N_10795);
xor U10866 (N_10866,N_10594,N_10668);
or U10867 (N_10867,N_10574,N_10666);
nand U10868 (N_10868,N_10714,N_10760);
and U10869 (N_10869,N_10793,N_10789);
or U10870 (N_10870,N_10650,N_10643);
or U10871 (N_10871,N_10628,N_10782);
and U10872 (N_10872,N_10614,N_10555);
nor U10873 (N_10873,N_10702,N_10509);
or U10874 (N_10874,N_10545,N_10589);
xnor U10875 (N_10875,N_10590,N_10778);
nor U10876 (N_10876,N_10785,N_10613);
or U10877 (N_10877,N_10790,N_10687);
xnor U10878 (N_10878,N_10609,N_10605);
nand U10879 (N_10879,N_10752,N_10675);
nand U10880 (N_10880,N_10606,N_10724);
nor U10881 (N_10881,N_10611,N_10500);
nand U10882 (N_10882,N_10725,N_10624);
and U10883 (N_10883,N_10768,N_10745);
and U10884 (N_10884,N_10612,N_10602);
nand U10885 (N_10885,N_10731,N_10603);
and U10886 (N_10886,N_10563,N_10680);
nor U10887 (N_10887,N_10787,N_10655);
or U10888 (N_10888,N_10740,N_10640);
and U10889 (N_10889,N_10639,N_10527);
nand U10890 (N_10890,N_10583,N_10771);
or U10891 (N_10891,N_10627,N_10764);
nor U10892 (N_10892,N_10560,N_10569);
xor U10893 (N_10893,N_10674,N_10762);
or U10894 (N_10894,N_10781,N_10549);
xor U10895 (N_10895,N_10542,N_10658);
nor U10896 (N_10896,N_10715,N_10747);
xnor U10897 (N_10897,N_10518,N_10719);
xnor U10898 (N_10898,N_10703,N_10530);
nand U10899 (N_10899,N_10772,N_10608);
or U10900 (N_10900,N_10705,N_10794);
and U10901 (N_10901,N_10566,N_10672);
nand U10902 (N_10902,N_10685,N_10548);
or U10903 (N_10903,N_10652,N_10617);
nand U10904 (N_10904,N_10656,N_10784);
nor U10905 (N_10905,N_10755,N_10720);
and U10906 (N_10906,N_10562,N_10748);
or U10907 (N_10907,N_10506,N_10671);
or U10908 (N_10908,N_10541,N_10751);
xor U10909 (N_10909,N_10730,N_10621);
or U10910 (N_10910,N_10776,N_10620);
or U10911 (N_10911,N_10520,N_10792);
nand U10912 (N_10912,N_10552,N_10754);
xnor U10913 (N_10913,N_10559,N_10529);
nor U10914 (N_10914,N_10635,N_10718);
or U10915 (N_10915,N_10739,N_10634);
and U10916 (N_10916,N_10661,N_10756);
or U10917 (N_10917,N_10691,N_10713);
nor U10918 (N_10918,N_10701,N_10667);
or U10919 (N_10919,N_10728,N_10799);
nor U10920 (N_10920,N_10791,N_10543);
nor U10921 (N_10921,N_10696,N_10547);
or U10922 (N_10922,N_10669,N_10501);
xor U10923 (N_10923,N_10665,N_10524);
and U10924 (N_10924,N_10653,N_10690);
xnor U10925 (N_10925,N_10610,N_10689);
or U10926 (N_10926,N_10657,N_10711);
nor U10927 (N_10927,N_10710,N_10706);
nor U10928 (N_10928,N_10592,N_10645);
or U10929 (N_10929,N_10514,N_10700);
xnor U10930 (N_10930,N_10535,N_10733);
nand U10931 (N_10931,N_10585,N_10593);
or U10932 (N_10932,N_10765,N_10779);
nor U10933 (N_10933,N_10507,N_10510);
and U10934 (N_10934,N_10766,N_10578);
or U10935 (N_10935,N_10649,N_10513);
or U10936 (N_10936,N_10512,N_10648);
and U10937 (N_10937,N_10533,N_10664);
or U10938 (N_10938,N_10519,N_10591);
or U10939 (N_10939,N_10753,N_10749);
nand U10940 (N_10940,N_10632,N_10557);
nor U10941 (N_10941,N_10708,N_10597);
nand U10942 (N_10942,N_10565,N_10646);
or U10943 (N_10943,N_10682,N_10553);
xnor U10944 (N_10944,N_10692,N_10797);
xnor U10945 (N_10945,N_10742,N_10769);
xnor U10946 (N_10946,N_10526,N_10561);
xnor U10947 (N_10947,N_10625,N_10584);
xnor U10948 (N_10948,N_10600,N_10695);
nand U10949 (N_10949,N_10727,N_10517);
xor U10950 (N_10950,N_10707,N_10563);
and U10951 (N_10951,N_10577,N_10626);
and U10952 (N_10952,N_10701,N_10775);
or U10953 (N_10953,N_10691,N_10770);
xnor U10954 (N_10954,N_10564,N_10535);
nor U10955 (N_10955,N_10732,N_10634);
nand U10956 (N_10956,N_10628,N_10658);
xnor U10957 (N_10957,N_10554,N_10605);
or U10958 (N_10958,N_10756,N_10542);
nor U10959 (N_10959,N_10659,N_10751);
or U10960 (N_10960,N_10669,N_10549);
xor U10961 (N_10961,N_10524,N_10712);
nand U10962 (N_10962,N_10724,N_10795);
xnor U10963 (N_10963,N_10613,N_10547);
xnor U10964 (N_10964,N_10556,N_10781);
and U10965 (N_10965,N_10545,N_10574);
xor U10966 (N_10966,N_10552,N_10734);
xnor U10967 (N_10967,N_10639,N_10776);
and U10968 (N_10968,N_10600,N_10636);
and U10969 (N_10969,N_10588,N_10619);
nand U10970 (N_10970,N_10556,N_10606);
and U10971 (N_10971,N_10679,N_10524);
and U10972 (N_10972,N_10543,N_10507);
or U10973 (N_10973,N_10563,N_10571);
and U10974 (N_10974,N_10779,N_10715);
or U10975 (N_10975,N_10533,N_10684);
and U10976 (N_10976,N_10621,N_10508);
nor U10977 (N_10977,N_10767,N_10592);
xor U10978 (N_10978,N_10610,N_10636);
nand U10979 (N_10979,N_10570,N_10651);
xnor U10980 (N_10980,N_10675,N_10725);
or U10981 (N_10981,N_10721,N_10647);
and U10982 (N_10982,N_10572,N_10663);
and U10983 (N_10983,N_10685,N_10649);
xnor U10984 (N_10984,N_10739,N_10599);
nand U10985 (N_10985,N_10682,N_10660);
and U10986 (N_10986,N_10759,N_10599);
or U10987 (N_10987,N_10782,N_10702);
or U10988 (N_10988,N_10725,N_10620);
xnor U10989 (N_10989,N_10711,N_10715);
and U10990 (N_10990,N_10649,N_10556);
nand U10991 (N_10991,N_10568,N_10598);
nor U10992 (N_10992,N_10743,N_10515);
nor U10993 (N_10993,N_10690,N_10717);
xor U10994 (N_10994,N_10798,N_10794);
nor U10995 (N_10995,N_10778,N_10561);
xor U10996 (N_10996,N_10770,N_10602);
and U10997 (N_10997,N_10660,N_10586);
xnor U10998 (N_10998,N_10635,N_10557);
nand U10999 (N_10999,N_10517,N_10586);
or U11000 (N_11000,N_10646,N_10762);
nand U11001 (N_11001,N_10701,N_10628);
xor U11002 (N_11002,N_10773,N_10618);
and U11003 (N_11003,N_10688,N_10704);
nor U11004 (N_11004,N_10566,N_10633);
and U11005 (N_11005,N_10620,N_10727);
or U11006 (N_11006,N_10647,N_10691);
nor U11007 (N_11007,N_10612,N_10653);
nor U11008 (N_11008,N_10737,N_10625);
or U11009 (N_11009,N_10688,N_10577);
or U11010 (N_11010,N_10631,N_10763);
nand U11011 (N_11011,N_10683,N_10788);
nand U11012 (N_11012,N_10694,N_10575);
nor U11013 (N_11013,N_10530,N_10745);
xnor U11014 (N_11014,N_10774,N_10602);
nor U11015 (N_11015,N_10536,N_10781);
nand U11016 (N_11016,N_10584,N_10602);
xor U11017 (N_11017,N_10792,N_10659);
nand U11018 (N_11018,N_10545,N_10667);
nor U11019 (N_11019,N_10633,N_10782);
nand U11020 (N_11020,N_10752,N_10652);
or U11021 (N_11021,N_10550,N_10503);
xor U11022 (N_11022,N_10681,N_10626);
or U11023 (N_11023,N_10702,N_10718);
or U11024 (N_11024,N_10771,N_10642);
and U11025 (N_11025,N_10712,N_10702);
nand U11026 (N_11026,N_10524,N_10505);
nor U11027 (N_11027,N_10586,N_10630);
and U11028 (N_11028,N_10554,N_10666);
or U11029 (N_11029,N_10692,N_10562);
xnor U11030 (N_11030,N_10684,N_10615);
nor U11031 (N_11031,N_10545,N_10793);
or U11032 (N_11032,N_10668,N_10615);
nand U11033 (N_11033,N_10738,N_10680);
xnor U11034 (N_11034,N_10506,N_10551);
xnor U11035 (N_11035,N_10745,N_10700);
nand U11036 (N_11036,N_10549,N_10566);
and U11037 (N_11037,N_10758,N_10705);
or U11038 (N_11038,N_10514,N_10783);
nand U11039 (N_11039,N_10544,N_10647);
xnor U11040 (N_11040,N_10524,N_10652);
nor U11041 (N_11041,N_10789,N_10638);
xnor U11042 (N_11042,N_10648,N_10745);
nor U11043 (N_11043,N_10751,N_10543);
and U11044 (N_11044,N_10514,N_10695);
and U11045 (N_11045,N_10662,N_10583);
xor U11046 (N_11046,N_10789,N_10773);
and U11047 (N_11047,N_10556,N_10671);
nand U11048 (N_11048,N_10686,N_10734);
nand U11049 (N_11049,N_10702,N_10720);
xnor U11050 (N_11050,N_10505,N_10685);
xnor U11051 (N_11051,N_10660,N_10514);
xnor U11052 (N_11052,N_10701,N_10643);
nor U11053 (N_11053,N_10606,N_10630);
xor U11054 (N_11054,N_10744,N_10667);
and U11055 (N_11055,N_10742,N_10534);
or U11056 (N_11056,N_10614,N_10706);
or U11057 (N_11057,N_10586,N_10777);
nor U11058 (N_11058,N_10759,N_10566);
and U11059 (N_11059,N_10702,N_10599);
and U11060 (N_11060,N_10778,N_10710);
xnor U11061 (N_11061,N_10719,N_10534);
nand U11062 (N_11062,N_10698,N_10641);
and U11063 (N_11063,N_10787,N_10686);
xnor U11064 (N_11064,N_10553,N_10556);
nand U11065 (N_11065,N_10551,N_10752);
or U11066 (N_11066,N_10676,N_10505);
or U11067 (N_11067,N_10719,N_10627);
or U11068 (N_11068,N_10672,N_10796);
xnor U11069 (N_11069,N_10580,N_10576);
nor U11070 (N_11070,N_10741,N_10755);
xnor U11071 (N_11071,N_10720,N_10561);
xor U11072 (N_11072,N_10747,N_10501);
xnor U11073 (N_11073,N_10695,N_10616);
and U11074 (N_11074,N_10618,N_10540);
nor U11075 (N_11075,N_10608,N_10545);
and U11076 (N_11076,N_10551,N_10679);
or U11077 (N_11077,N_10735,N_10737);
or U11078 (N_11078,N_10580,N_10536);
nand U11079 (N_11079,N_10533,N_10741);
and U11080 (N_11080,N_10620,N_10634);
or U11081 (N_11081,N_10627,N_10621);
and U11082 (N_11082,N_10716,N_10544);
xnor U11083 (N_11083,N_10519,N_10529);
or U11084 (N_11084,N_10791,N_10622);
nor U11085 (N_11085,N_10528,N_10598);
or U11086 (N_11086,N_10735,N_10721);
nor U11087 (N_11087,N_10580,N_10544);
nor U11088 (N_11088,N_10747,N_10527);
nor U11089 (N_11089,N_10579,N_10643);
nand U11090 (N_11090,N_10768,N_10700);
xnor U11091 (N_11091,N_10571,N_10508);
nand U11092 (N_11092,N_10697,N_10549);
nand U11093 (N_11093,N_10533,N_10579);
or U11094 (N_11094,N_10711,N_10654);
nor U11095 (N_11095,N_10779,N_10520);
and U11096 (N_11096,N_10528,N_10620);
xnor U11097 (N_11097,N_10664,N_10572);
nand U11098 (N_11098,N_10622,N_10588);
xnor U11099 (N_11099,N_10562,N_10694);
xnor U11100 (N_11100,N_10829,N_11062);
nand U11101 (N_11101,N_10999,N_11091);
xnor U11102 (N_11102,N_10863,N_11044);
or U11103 (N_11103,N_10869,N_11040);
nor U11104 (N_11104,N_10926,N_10940);
and U11105 (N_11105,N_10824,N_11002);
nor U11106 (N_11106,N_10996,N_10850);
nor U11107 (N_11107,N_10929,N_10836);
nand U11108 (N_11108,N_10963,N_11011);
and U11109 (N_11109,N_10826,N_10902);
and U11110 (N_11110,N_10942,N_10965);
nor U11111 (N_11111,N_10854,N_11050);
xnor U11112 (N_11112,N_10953,N_11046);
nor U11113 (N_11113,N_10847,N_10807);
or U11114 (N_11114,N_10907,N_10886);
nand U11115 (N_11115,N_10858,N_10835);
or U11116 (N_11116,N_10985,N_11007);
or U11117 (N_11117,N_10892,N_11003);
xnor U11118 (N_11118,N_11070,N_11090);
and U11119 (N_11119,N_10859,N_10843);
nor U11120 (N_11120,N_10832,N_10805);
nand U11121 (N_11121,N_11028,N_10846);
xor U11122 (N_11122,N_10868,N_10816);
nor U11123 (N_11123,N_10825,N_10918);
xnor U11124 (N_11124,N_11025,N_11030);
xor U11125 (N_11125,N_11076,N_10899);
or U11126 (N_11126,N_10975,N_10870);
nand U11127 (N_11127,N_10877,N_10928);
nand U11128 (N_11128,N_11072,N_10946);
or U11129 (N_11129,N_11022,N_10900);
nor U11130 (N_11130,N_10806,N_10849);
and U11131 (N_11131,N_11010,N_10984);
nand U11132 (N_11132,N_11019,N_11052);
or U11133 (N_11133,N_11066,N_10920);
nand U11134 (N_11134,N_10915,N_11001);
and U11135 (N_11135,N_10973,N_10980);
or U11136 (N_11136,N_10954,N_11012);
and U11137 (N_11137,N_10943,N_10864);
or U11138 (N_11138,N_10947,N_11094);
or U11139 (N_11139,N_10887,N_10823);
or U11140 (N_11140,N_10983,N_11021);
and U11141 (N_11141,N_11027,N_10866);
or U11142 (N_11142,N_10960,N_10917);
and U11143 (N_11143,N_10951,N_11031);
nor U11144 (N_11144,N_11055,N_11064);
or U11145 (N_11145,N_10974,N_10851);
nor U11146 (N_11146,N_10803,N_10867);
xor U11147 (N_11147,N_11075,N_11005);
and U11148 (N_11148,N_10986,N_10989);
nor U11149 (N_11149,N_10971,N_10898);
nor U11150 (N_11150,N_11054,N_11000);
xnor U11151 (N_11151,N_10922,N_11089);
xor U11152 (N_11152,N_10968,N_11071);
nand U11153 (N_11153,N_11018,N_10873);
nand U11154 (N_11154,N_10855,N_10978);
nor U11155 (N_11155,N_11082,N_10879);
nand U11156 (N_11156,N_10895,N_10821);
nor U11157 (N_11157,N_10876,N_11015);
nor U11158 (N_11158,N_10959,N_10808);
xor U11159 (N_11159,N_11096,N_10995);
nand U11160 (N_11160,N_11098,N_10813);
nand U11161 (N_11161,N_10802,N_10828);
xor U11162 (N_11162,N_11006,N_11093);
xnor U11163 (N_11163,N_10822,N_10804);
nand U11164 (N_11164,N_10830,N_10931);
or U11165 (N_11165,N_10890,N_10800);
nand U11166 (N_11166,N_11061,N_10982);
nor U11167 (N_11167,N_10815,N_10927);
nor U11168 (N_11168,N_10941,N_10871);
nor U11169 (N_11169,N_10919,N_10993);
and U11170 (N_11170,N_10812,N_11074);
xnor U11171 (N_11171,N_10834,N_11014);
and U11172 (N_11172,N_10932,N_11058);
nand U11173 (N_11173,N_10938,N_11016);
or U11174 (N_11174,N_11023,N_11037);
and U11175 (N_11175,N_10820,N_10958);
nand U11176 (N_11176,N_11029,N_11097);
or U11177 (N_11177,N_11095,N_10930);
nor U11178 (N_11178,N_10911,N_10889);
nand U11179 (N_11179,N_11048,N_11083);
xnor U11180 (N_11180,N_10934,N_10981);
xor U11181 (N_11181,N_11073,N_10909);
and U11182 (N_11182,N_10977,N_10833);
xnor U11183 (N_11183,N_11063,N_11041);
nand U11184 (N_11184,N_10979,N_10914);
nand U11185 (N_11185,N_10924,N_11068);
and U11186 (N_11186,N_11065,N_10969);
or U11187 (N_11187,N_10861,N_11035);
or U11188 (N_11188,N_10970,N_10976);
nand U11189 (N_11189,N_10881,N_10857);
and U11190 (N_11190,N_10801,N_10841);
nor U11191 (N_11191,N_10860,N_11008);
nand U11192 (N_11192,N_10883,N_10901);
nor U11193 (N_11193,N_10818,N_11056);
and U11194 (N_11194,N_11045,N_10945);
nor U11195 (N_11195,N_10937,N_11034);
nand U11196 (N_11196,N_10988,N_11099);
xor U11197 (N_11197,N_10809,N_11077);
nor U11198 (N_11198,N_10852,N_10967);
and U11199 (N_11199,N_10888,N_10956);
nand U11200 (N_11200,N_11042,N_10961);
nor U11201 (N_11201,N_10831,N_10839);
and U11202 (N_11202,N_11043,N_10936);
xnor U11203 (N_11203,N_10935,N_10882);
nor U11204 (N_11204,N_10811,N_10904);
xor U11205 (N_11205,N_11078,N_10933);
and U11206 (N_11206,N_10819,N_10842);
nand U11207 (N_11207,N_10905,N_11024);
and U11208 (N_11208,N_10908,N_10952);
nor U11209 (N_11209,N_11081,N_11051);
nand U11210 (N_11210,N_10878,N_11033);
nor U11211 (N_11211,N_10817,N_11038);
xor U11212 (N_11212,N_10923,N_11088);
xor U11213 (N_11213,N_10991,N_10994);
nor U11214 (N_11214,N_11026,N_10948);
nor U11215 (N_11215,N_11013,N_11036);
or U11216 (N_11216,N_10827,N_10955);
and U11217 (N_11217,N_10875,N_10957);
or U11218 (N_11218,N_10972,N_10862);
or U11219 (N_11219,N_10998,N_11087);
or U11220 (N_11220,N_10939,N_11020);
nor U11221 (N_11221,N_11009,N_10853);
nor U11222 (N_11222,N_11069,N_10894);
and U11223 (N_11223,N_11047,N_10814);
and U11224 (N_11224,N_10949,N_10872);
nand U11225 (N_11225,N_10912,N_10885);
nand U11226 (N_11226,N_10838,N_10840);
nand U11227 (N_11227,N_11084,N_11080);
xor U11228 (N_11228,N_11085,N_10845);
nand U11229 (N_11229,N_10990,N_10896);
or U11230 (N_11230,N_10966,N_10964);
and U11231 (N_11231,N_10884,N_10880);
and U11232 (N_11232,N_11086,N_11059);
nor U11233 (N_11233,N_10903,N_10865);
and U11234 (N_11234,N_10944,N_11049);
nor U11235 (N_11235,N_10910,N_10987);
nor U11236 (N_11236,N_10913,N_10856);
nand U11237 (N_11237,N_11053,N_10810);
or U11238 (N_11238,N_11004,N_10837);
or U11239 (N_11239,N_11067,N_10874);
and U11240 (N_11240,N_11032,N_10897);
xor U11241 (N_11241,N_10962,N_10916);
or U11242 (N_11242,N_10950,N_10925);
nor U11243 (N_11243,N_10997,N_11092);
nand U11244 (N_11244,N_10921,N_11039);
nor U11245 (N_11245,N_10893,N_10992);
nor U11246 (N_11246,N_10891,N_10844);
xnor U11247 (N_11247,N_11017,N_10906);
or U11248 (N_11248,N_11060,N_11079);
xnor U11249 (N_11249,N_10848,N_11057);
nand U11250 (N_11250,N_10866,N_10971);
and U11251 (N_11251,N_11003,N_11067);
xor U11252 (N_11252,N_11053,N_10913);
or U11253 (N_11253,N_11067,N_10802);
nand U11254 (N_11254,N_10904,N_10885);
nor U11255 (N_11255,N_11081,N_10893);
and U11256 (N_11256,N_10926,N_10959);
and U11257 (N_11257,N_10929,N_11065);
and U11258 (N_11258,N_10918,N_10960);
nor U11259 (N_11259,N_10821,N_11053);
nand U11260 (N_11260,N_10909,N_11003);
and U11261 (N_11261,N_10979,N_11072);
or U11262 (N_11262,N_11068,N_11020);
xor U11263 (N_11263,N_11075,N_10830);
nand U11264 (N_11264,N_10922,N_10982);
xor U11265 (N_11265,N_11046,N_10948);
or U11266 (N_11266,N_10976,N_11078);
and U11267 (N_11267,N_11052,N_11095);
and U11268 (N_11268,N_10890,N_10906);
xnor U11269 (N_11269,N_10972,N_10886);
xnor U11270 (N_11270,N_10980,N_10992);
xor U11271 (N_11271,N_10910,N_10902);
nor U11272 (N_11272,N_10910,N_11073);
xor U11273 (N_11273,N_11014,N_10868);
nor U11274 (N_11274,N_11052,N_10973);
or U11275 (N_11275,N_10895,N_10917);
or U11276 (N_11276,N_10811,N_11050);
xor U11277 (N_11277,N_11098,N_10914);
nand U11278 (N_11278,N_11059,N_10884);
nand U11279 (N_11279,N_10889,N_10996);
or U11280 (N_11280,N_10841,N_10851);
or U11281 (N_11281,N_10942,N_10828);
or U11282 (N_11282,N_11073,N_10816);
xor U11283 (N_11283,N_11057,N_10899);
nand U11284 (N_11284,N_10933,N_11081);
and U11285 (N_11285,N_11047,N_11084);
xnor U11286 (N_11286,N_10960,N_11099);
nand U11287 (N_11287,N_10997,N_11064);
or U11288 (N_11288,N_10860,N_11052);
xor U11289 (N_11289,N_10835,N_10965);
and U11290 (N_11290,N_11068,N_11039);
and U11291 (N_11291,N_10964,N_10988);
xor U11292 (N_11292,N_11027,N_11033);
nor U11293 (N_11293,N_11053,N_10811);
nor U11294 (N_11294,N_11046,N_11037);
nand U11295 (N_11295,N_11069,N_10931);
or U11296 (N_11296,N_10877,N_10843);
nor U11297 (N_11297,N_11095,N_10883);
xor U11298 (N_11298,N_11029,N_11038);
nor U11299 (N_11299,N_11068,N_10808);
xor U11300 (N_11300,N_10952,N_10847);
nor U11301 (N_11301,N_10809,N_10985);
or U11302 (N_11302,N_10975,N_11054);
or U11303 (N_11303,N_11065,N_10917);
nor U11304 (N_11304,N_10888,N_10931);
or U11305 (N_11305,N_11047,N_10987);
or U11306 (N_11306,N_10966,N_11070);
nand U11307 (N_11307,N_11061,N_10981);
nand U11308 (N_11308,N_11064,N_11017);
or U11309 (N_11309,N_11089,N_10856);
and U11310 (N_11310,N_10881,N_10870);
nand U11311 (N_11311,N_11029,N_11065);
xor U11312 (N_11312,N_11072,N_11058);
or U11313 (N_11313,N_10866,N_10856);
nand U11314 (N_11314,N_10917,N_11010);
nor U11315 (N_11315,N_10972,N_11063);
nor U11316 (N_11316,N_10919,N_10882);
xnor U11317 (N_11317,N_10973,N_11042);
or U11318 (N_11318,N_10912,N_11049);
and U11319 (N_11319,N_10954,N_11055);
and U11320 (N_11320,N_10834,N_10822);
nor U11321 (N_11321,N_10975,N_10807);
and U11322 (N_11322,N_11096,N_11092);
nand U11323 (N_11323,N_11015,N_11087);
xnor U11324 (N_11324,N_10913,N_10861);
nor U11325 (N_11325,N_10915,N_10812);
and U11326 (N_11326,N_10905,N_10881);
nand U11327 (N_11327,N_11091,N_10895);
or U11328 (N_11328,N_10893,N_10957);
xnor U11329 (N_11329,N_10869,N_11033);
xor U11330 (N_11330,N_10852,N_10814);
and U11331 (N_11331,N_10972,N_10866);
xor U11332 (N_11332,N_10932,N_11060);
nand U11333 (N_11333,N_10863,N_10878);
xnor U11334 (N_11334,N_10812,N_11019);
and U11335 (N_11335,N_10851,N_11089);
xnor U11336 (N_11336,N_10906,N_10824);
nor U11337 (N_11337,N_11042,N_10937);
xnor U11338 (N_11338,N_11051,N_10825);
xnor U11339 (N_11339,N_10839,N_10893);
nor U11340 (N_11340,N_10855,N_10859);
and U11341 (N_11341,N_10952,N_10949);
and U11342 (N_11342,N_11031,N_10924);
nand U11343 (N_11343,N_11016,N_10944);
xor U11344 (N_11344,N_11040,N_11066);
and U11345 (N_11345,N_10967,N_10956);
or U11346 (N_11346,N_11072,N_10862);
xor U11347 (N_11347,N_10869,N_10990);
nor U11348 (N_11348,N_11022,N_10899);
or U11349 (N_11349,N_10834,N_10803);
or U11350 (N_11350,N_10804,N_10895);
or U11351 (N_11351,N_10815,N_11017);
nor U11352 (N_11352,N_10858,N_10982);
and U11353 (N_11353,N_11046,N_11052);
or U11354 (N_11354,N_10908,N_10902);
and U11355 (N_11355,N_11044,N_11082);
and U11356 (N_11356,N_10902,N_10974);
nand U11357 (N_11357,N_11097,N_11096);
or U11358 (N_11358,N_10844,N_10893);
and U11359 (N_11359,N_11017,N_10924);
xnor U11360 (N_11360,N_10946,N_10819);
nor U11361 (N_11361,N_11090,N_10994);
nand U11362 (N_11362,N_10801,N_11014);
nor U11363 (N_11363,N_10916,N_10986);
nand U11364 (N_11364,N_10947,N_10996);
nand U11365 (N_11365,N_10899,N_10864);
nand U11366 (N_11366,N_11099,N_10807);
xnor U11367 (N_11367,N_10889,N_11072);
or U11368 (N_11368,N_10966,N_10908);
or U11369 (N_11369,N_10818,N_11005);
or U11370 (N_11370,N_10868,N_10843);
nor U11371 (N_11371,N_11039,N_11051);
xor U11372 (N_11372,N_10971,N_10810);
and U11373 (N_11373,N_11096,N_10905);
xnor U11374 (N_11374,N_11024,N_10820);
nand U11375 (N_11375,N_11019,N_10816);
nor U11376 (N_11376,N_10863,N_10908);
xnor U11377 (N_11377,N_10878,N_10859);
nor U11378 (N_11378,N_11033,N_10877);
and U11379 (N_11379,N_10900,N_10982);
or U11380 (N_11380,N_10864,N_11074);
xnor U11381 (N_11381,N_10962,N_11070);
and U11382 (N_11382,N_10814,N_10842);
and U11383 (N_11383,N_11019,N_10840);
xnor U11384 (N_11384,N_10810,N_10825);
xor U11385 (N_11385,N_10900,N_10907);
or U11386 (N_11386,N_11038,N_10851);
nand U11387 (N_11387,N_11046,N_11065);
or U11388 (N_11388,N_10877,N_10958);
nand U11389 (N_11389,N_10831,N_10969);
or U11390 (N_11390,N_10990,N_11096);
and U11391 (N_11391,N_11059,N_11072);
nand U11392 (N_11392,N_11006,N_11087);
and U11393 (N_11393,N_10803,N_10980);
xnor U11394 (N_11394,N_10953,N_10869);
nor U11395 (N_11395,N_10865,N_10814);
nand U11396 (N_11396,N_10843,N_10810);
nor U11397 (N_11397,N_11071,N_10809);
or U11398 (N_11398,N_10982,N_11015);
or U11399 (N_11399,N_11036,N_10993);
or U11400 (N_11400,N_11181,N_11254);
or U11401 (N_11401,N_11284,N_11331);
nand U11402 (N_11402,N_11103,N_11380);
and U11403 (N_11403,N_11269,N_11348);
nand U11404 (N_11404,N_11264,N_11302);
and U11405 (N_11405,N_11190,N_11147);
or U11406 (N_11406,N_11305,N_11385);
xor U11407 (N_11407,N_11361,N_11393);
nor U11408 (N_11408,N_11364,N_11358);
nand U11409 (N_11409,N_11367,N_11298);
or U11410 (N_11410,N_11225,N_11363);
nor U11411 (N_11411,N_11198,N_11274);
nand U11412 (N_11412,N_11160,N_11194);
or U11413 (N_11413,N_11262,N_11118);
nand U11414 (N_11414,N_11365,N_11180);
and U11415 (N_11415,N_11143,N_11173);
nor U11416 (N_11416,N_11316,N_11148);
xor U11417 (N_11417,N_11165,N_11244);
nand U11418 (N_11418,N_11170,N_11294);
nand U11419 (N_11419,N_11359,N_11101);
nand U11420 (N_11420,N_11155,N_11395);
and U11421 (N_11421,N_11205,N_11119);
nand U11422 (N_11422,N_11326,N_11357);
xor U11423 (N_11423,N_11156,N_11166);
xor U11424 (N_11424,N_11212,N_11164);
nand U11425 (N_11425,N_11292,N_11152);
xor U11426 (N_11426,N_11209,N_11340);
or U11427 (N_11427,N_11157,N_11182);
or U11428 (N_11428,N_11246,N_11161);
and U11429 (N_11429,N_11261,N_11347);
or U11430 (N_11430,N_11153,N_11311);
and U11431 (N_11431,N_11231,N_11237);
nand U11432 (N_11432,N_11317,N_11123);
or U11433 (N_11433,N_11250,N_11360);
or U11434 (N_11434,N_11336,N_11247);
nand U11435 (N_11435,N_11169,N_11323);
nand U11436 (N_11436,N_11189,N_11200);
or U11437 (N_11437,N_11276,N_11120);
nand U11438 (N_11438,N_11343,N_11327);
nor U11439 (N_11439,N_11381,N_11228);
nand U11440 (N_11440,N_11187,N_11387);
nand U11441 (N_11441,N_11211,N_11345);
nand U11442 (N_11442,N_11279,N_11272);
nand U11443 (N_11443,N_11275,N_11158);
or U11444 (N_11444,N_11337,N_11307);
or U11445 (N_11445,N_11122,N_11174);
and U11446 (N_11446,N_11328,N_11146);
and U11447 (N_11447,N_11203,N_11338);
or U11448 (N_11448,N_11290,N_11249);
or U11449 (N_11449,N_11133,N_11273);
or U11450 (N_11450,N_11396,N_11135);
or U11451 (N_11451,N_11177,N_11121);
or U11452 (N_11452,N_11176,N_11139);
and U11453 (N_11453,N_11394,N_11219);
or U11454 (N_11454,N_11356,N_11382);
nand U11455 (N_11455,N_11224,N_11255);
nand U11456 (N_11456,N_11227,N_11350);
and U11457 (N_11457,N_11389,N_11130);
nand U11458 (N_11458,N_11131,N_11397);
nand U11459 (N_11459,N_11142,N_11287);
or U11460 (N_11460,N_11339,N_11222);
or U11461 (N_11461,N_11217,N_11175);
nand U11462 (N_11462,N_11334,N_11283);
nand U11463 (N_11463,N_11301,N_11253);
xor U11464 (N_11464,N_11304,N_11383);
nor U11465 (N_11465,N_11377,N_11293);
nor U11466 (N_11466,N_11235,N_11313);
nor U11467 (N_11467,N_11234,N_11391);
nor U11468 (N_11468,N_11163,N_11136);
nor U11469 (N_11469,N_11168,N_11116);
or U11470 (N_11470,N_11353,N_11315);
or U11471 (N_11471,N_11221,N_11126);
or U11472 (N_11472,N_11109,N_11243);
xor U11473 (N_11473,N_11240,N_11236);
nor U11474 (N_11474,N_11127,N_11266);
xnor U11475 (N_11475,N_11330,N_11325);
nand U11476 (N_11476,N_11199,N_11207);
or U11477 (N_11477,N_11281,N_11320);
xor U11478 (N_11478,N_11151,N_11218);
or U11479 (N_11479,N_11329,N_11140);
or U11480 (N_11480,N_11312,N_11179);
nand U11481 (N_11481,N_11132,N_11223);
or U11482 (N_11482,N_11362,N_11251);
or U11483 (N_11483,N_11270,N_11300);
or U11484 (N_11484,N_11289,N_11260);
xor U11485 (N_11485,N_11178,N_11378);
or U11486 (N_11486,N_11241,N_11271);
nand U11487 (N_11487,N_11355,N_11319);
and U11488 (N_11488,N_11303,N_11159);
nand U11489 (N_11489,N_11308,N_11333);
xnor U11490 (N_11490,N_11242,N_11332);
xnor U11491 (N_11491,N_11280,N_11117);
and U11492 (N_11492,N_11299,N_11215);
or U11493 (N_11493,N_11149,N_11196);
nor U11494 (N_11494,N_11105,N_11229);
nand U11495 (N_11495,N_11233,N_11314);
or U11496 (N_11496,N_11351,N_11171);
nor U11497 (N_11497,N_11318,N_11386);
nor U11498 (N_11498,N_11115,N_11112);
xor U11499 (N_11499,N_11296,N_11193);
or U11500 (N_11500,N_11108,N_11384);
nor U11501 (N_11501,N_11344,N_11100);
and U11502 (N_11502,N_11369,N_11232);
nand U11503 (N_11503,N_11341,N_11259);
and U11504 (N_11504,N_11214,N_11192);
nor U11505 (N_11505,N_11376,N_11278);
nand U11506 (N_11506,N_11322,N_11398);
or U11507 (N_11507,N_11371,N_11107);
and U11508 (N_11508,N_11388,N_11286);
and U11509 (N_11509,N_11210,N_11113);
xnor U11510 (N_11510,N_11238,N_11288);
and U11511 (N_11511,N_11372,N_11102);
and U11512 (N_11512,N_11216,N_11268);
or U11513 (N_11513,N_11134,N_11206);
xnor U11514 (N_11514,N_11342,N_11125);
nand U11515 (N_11515,N_11208,N_11129);
xor U11516 (N_11516,N_11368,N_11267);
nand U11517 (N_11517,N_11263,N_11110);
nand U11518 (N_11518,N_11295,N_11201);
xor U11519 (N_11519,N_11309,N_11213);
nand U11520 (N_11520,N_11186,N_11252);
xor U11521 (N_11521,N_11310,N_11366);
nand U11522 (N_11522,N_11204,N_11144);
nor U11523 (N_11523,N_11154,N_11258);
or U11524 (N_11524,N_11124,N_11202);
xnor U11525 (N_11525,N_11162,N_11306);
or U11526 (N_11526,N_11245,N_11197);
or U11527 (N_11527,N_11230,N_11373);
and U11528 (N_11528,N_11277,N_11141);
xnor U11529 (N_11529,N_11150,N_11335);
nand U11530 (N_11530,N_11137,N_11167);
and U11531 (N_11531,N_11172,N_11248);
and U11532 (N_11532,N_11185,N_11379);
nand U11533 (N_11533,N_11282,N_11354);
nand U11534 (N_11534,N_11375,N_11352);
nand U11535 (N_11535,N_11184,N_11257);
nand U11536 (N_11536,N_11239,N_11138);
or U11537 (N_11537,N_11111,N_11128);
or U11538 (N_11538,N_11346,N_11285);
or U11539 (N_11539,N_11374,N_11256);
nand U11540 (N_11540,N_11265,N_11220);
or U11541 (N_11541,N_11349,N_11226);
or U11542 (N_11542,N_11392,N_11104);
nand U11543 (N_11543,N_11321,N_11114);
nand U11544 (N_11544,N_11106,N_11183);
nand U11545 (N_11545,N_11145,N_11291);
xor U11546 (N_11546,N_11191,N_11188);
nor U11547 (N_11547,N_11370,N_11399);
nor U11548 (N_11548,N_11324,N_11195);
and U11549 (N_11549,N_11297,N_11390);
xnor U11550 (N_11550,N_11315,N_11381);
nor U11551 (N_11551,N_11397,N_11313);
nand U11552 (N_11552,N_11279,N_11343);
nand U11553 (N_11553,N_11212,N_11261);
and U11554 (N_11554,N_11241,N_11276);
xor U11555 (N_11555,N_11349,N_11257);
xor U11556 (N_11556,N_11195,N_11197);
nor U11557 (N_11557,N_11287,N_11378);
and U11558 (N_11558,N_11329,N_11143);
xnor U11559 (N_11559,N_11216,N_11293);
xnor U11560 (N_11560,N_11128,N_11305);
nor U11561 (N_11561,N_11321,N_11278);
or U11562 (N_11562,N_11102,N_11232);
or U11563 (N_11563,N_11398,N_11314);
or U11564 (N_11564,N_11263,N_11160);
xor U11565 (N_11565,N_11167,N_11103);
nand U11566 (N_11566,N_11105,N_11367);
nand U11567 (N_11567,N_11379,N_11368);
nand U11568 (N_11568,N_11394,N_11170);
and U11569 (N_11569,N_11173,N_11207);
nand U11570 (N_11570,N_11209,N_11213);
nand U11571 (N_11571,N_11174,N_11279);
nand U11572 (N_11572,N_11111,N_11372);
and U11573 (N_11573,N_11286,N_11265);
nand U11574 (N_11574,N_11174,N_11119);
nand U11575 (N_11575,N_11292,N_11185);
or U11576 (N_11576,N_11245,N_11153);
or U11577 (N_11577,N_11334,N_11254);
nor U11578 (N_11578,N_11161,N_11111);
nand U11579 (N_11579,N_11231,N_11132);
and U11580 (N_11580,N_11281,N_11392);
xnor U11581 (N_11581,N_11397,N_11321);
nor U11582 (N_11582,N_11310,N_11176);
and U11583 (N_11583,N_11136,N_11241);
nor U11584 (N_11584,N_11302,N_11191);
or U11585 (N_11585,N_11220,N_11322);
nor U11586 (N_11586,N_11341,N_11311);
nor U11587 (N_11587,N_11314,N_11369);
xor U11588 (N_11588,N_11152,N_11377);
nand U11589 (N_11589,N_11133,N_11398);
nand U11590 (N_11590,N_11102,N_11389);
or U11591 (N_11591,N_11194,N_11126);
or U11592 (N_11592,N_11142,N_11240);
xnor U11593 (N_11593,N_11221,N_11361);
and U11594 (N_11594,N_11137,N_11135);
or U11595 (N_11595,N_11216,N_11353);
and U11596 (N_11596,N_11164,N_11286);
xor U11597 (N_11597,N_11342,N_11379);
xnor U11598 (N_11598,N_11263,N_11120);
nor U11599 (N_11599,N_11229,N_11387);
and U11600 (N_11600,N_11333,N_11226);
and U11601 (N_11601,N_11327,N_11108);
xnor U11602 (N_11602,N_11146,N_11200);
and U11603 (N_11603,N_11284,N_11371);
or U11604 (N_11604,N_11278,N_11398);
nor U11605 (N_11605,N_11298,N_11126);
or U11606 (N_11606,N_11242,N_11202);
nand U11607 (N_11607,N_11358,N_11241);
nor U11608 (N_11608,N_11264,N_11155);
nor U11609 (N_11609,N_11100,N_11335);
nor U11610 (N_11610,N_11319,N_11340);
nor U11611 (N_11611,N_11256,N_11120);
or U11612 (N_11612,N_11156,N_11130);
and U11613 (N_11613,N_11227,N_11165);
nor U11614 (N_11614,N_11203,N_11316);
nor U11615 (N_11615,N_11398,N_11137);
nor U11616 (N_11616,N_11351,N_11374);
xor U11617 (N_11617,N_11370,N_11174);
xor U11618 (N_11618,N_11193,N_11163);
or U11619 (N_11619,N_11285,N_11148);
xnor U11620 (N_11620,N_11311,N_11353);
xor U11621 (N_11621,N_11162,N_11123);
nor U11622 (N_11622,N_11315,N_11195);
xor U11623 (N_11623,N_11268,N_11122);
nor U11624 (N_11624,N_11100,N_11325);
nor U11625 (N_11625,N_11285,N_11121);
nand U11626 (N_11626,N_11216,N_11388);
or U11627 (N_11627,N_11249,N_11157);
nand U11628 (N_11628,N_11208,N_11309);
or U11629 (N_11629,N_11269,N_11329);
and U11630 (N_11630,N_11184,N_11120);
nand U11631 (N_11631,N_11393,N_11323);
or U11632 (N_11632,N_11302,N_11119);
nor U11633 (N_11633,N_11398,N_11223);
or U11634 (N_11634,N_11102,N_11134);
nor U11635 (N_11635,N_11121,N_11357);
nor U11636 (N_11636,N_11306,N_11300);
xnor U11637 (N_11637,N_11204,N_11223);
or U11638 (N_11638,N_11129,N_11373);
xor U11639 (N_11639,N_11138,N_11135);
or U11640 (N_11640,N_11359,N_11172);
nand U11641 (N_11641,N_11195,N_11261);
or U11642 (N_11642,N_11267,N_11392);
and U11643 (N_11643,N_11108,N_11132);
and U11644 (N_11644,N_11381,N_11395);
nand U11645 (N_11645,N_11225,N_11227);
or U11646 (N_11646,N_11392,N_11166);
nor U11647 (N_11647,N_11224,N_11143);
and U11648 (N_11648,N_11187,N_11112);
xor U11649 (N_11649,N_11289,N_11110);
and U11650 (N_11650,N_11185,N_11107);
or U11651 (N_11651,N_11189,N_11299);
and U11652 (N_11652,N_11209,N_11304);
xor U11653 (N_11653,N_11281,N_11131);
nand U11654 (N_11654,N_11171,N_11214);
xnor U11655 (N_11655,N_11106,N_11240);
or U11656 (N_11656,N_11221,N_11343);
nor U11657 (N_11657,N_11131,N_11199);
xor U11658 (N_11658,N_11124,N_11187);
nor U11659 (N_11659,N_11275,N_11246);
xnor U11660 (N_11660,N_11341,N_11115);
nand U11661 (N_11661,N_11235,N_11270);
and U11662 (N_11662,N_11139,N_11350);
nor U11663 (N_11663,N_11295,N_11103);
and U11664 (N_11664,N_11181,N_11207);
xor U11665 (N_11665,N_11333,N_11276);
and U11666 (N_11666,N_11382,N_11359);
or U11667 (N_11667,N_11137,N_11305);
and U11668 (N_11668,N_11100,N_11179);
nand U11669 (N_11669,N_11273,N_11318);
or U11670 (N_11670,N_11375,N_11317);
nor U11671 (N_11671,N_11305,N_11302);
nand U11672 (N_11672,N_11121,N_11201);
and U11673 (N_11673,N_11391,N_11319);
and U11674 (N_11674,N_11181,N_11107);
and U11675 (N_11675,N_11388,N_11256);
nor U11676 (N_11676,N_11330,N_11163);
nor U11677 (N_11677,N_11267,N_11396);
and U11678 (N_11678,N_11215,N_11194);
xor U11679 (N_11679,N_11252,N_11368);
nand U11680 (N_11680,N_11123,N_11236);
and U11681 (N_11681,N_11252,N_11331);
or U11682 (N_11682,N_11210,N_11341);
or U11683 (N_11683,N_11292,N_11124);
and U11684 (N_11684,N_11265,N_11103);
xor U11685 (N_11685,N_11242,N_11178);
or U11686 (N_11686,N_11213,N_11297);
nand U11687 (N_11687,N_11191,N_11248);
nor U11688 (N_11688,N_11217,N_11138);
xor U11689 (N_11689,N_11308,N_11290);
nor U11690 (N_11690,N_11264,N_11112);
or U11691 (N_11691,N_11154,N_11246);
xnor U11692 (N_11692,N_11182,N_11385);
nand U11693 (N_11693,N_11263,N_11187);
xor U11694 (N_11694,N_11162,N_11141);
nor U11695 (N_11695,N_11136,N_11230);
or U11696 (N_11696,N_11366,N_11275);
and U11697 (N_11697,N_11116,N_11281);
nand U11698 (N_11698,N_11333,N_11374);
and U11699 (N_11699,N_11116,N_11127);
or U11700 (N_11700,N_11649,N_11410);
xor U11701 (N_11701,N_11476,N_11551);
nand U11702 (N_11702,N_11627,N_11662);
nor U11703 (N_11703,N_11565,N_11496);
or U11704 (N_11704,N_11464,N_11610);
xor U11705 (N_11705,N_11698,N_11626);
and U11706 (N_11706,N_11575,N_11600);
nand U11707 (N_11707,N_11606,N_11446);
and U11708 (N_11708,N_11584,N_11502);
nand U11709 (N_11709,N_11460,N_11424);
xor U11710 (N_11710,N_11517,N_11532);
and U11711 (N_11711,N_11695,N_11455);
xnor U11712 (N_11712,N_11435,N_11580);
or U11713 (N_11713,N_11548,N_11540);
nor U11714 (N_11714,N_11433,N_11545);
and U11715 (N_11715,N_11522,N_11482);
nand U11716 (N_11716,N_11594,N_11526);
nand U11717 (N_11717,N_11509,N_11590);
and U11718 (N_11718,N_11596,N_11592);
and U11719 (N_11719,N_11426,N_11541);
and U11720 (N_11720,N_11549,N_11625);
and U11721 (N_11721,N_11642,N_11572);
or U11722 (N_11722,N_11680,N_11574);
or U11723 (N_11723,N_11688,N_11648);
nor U11724 (N_11724,N_11653,N_11402);
or U11725 (N_11725,N_11501,N_11519);
xor U11726 (N_11726,N_11576,N_11515);
xor U11727 (N_11727,N_11593,N_11524);
and U11728 (N_11728,N_11619,N_11673);
nor U11729 (N_11729,N_11414,N_11440);
nor U11730 (N_11730,N_11454,N_11546);
xor U11731 (N_11731,N_11559,N_11678);
nand U11732 (N_11732,N_11542,N_11666);
and U11733 (N_11733,N_11483,N_11437);
nand U11734 (N_11734,N_11462,N_11489);
nor U11735 (N_11735,N_11422,N_11612);
nand U11736 (N_11736,N_11658,N_11506);
and U11737 (N_11737,N_11553,N_11432);
nor U11738 (N_11738,N_11628,N_11487);
or U11739 (N_11739,N_11550,N_11652);
and U11740 (N_11740,N_11504,N_11685);
and U11741 (N_11741,N_11693,N_11493);
and U11742 (N_11742,N_11495,N_11692);
or U11743 (N_11743,N_11635,N_11566);
xor U11744 (N_11744,N_11654,N_11557);
and U11745 (N_11745,N_11441,N_11534);
nand U11746 (N_11746,N_11556,N_11547);
or U11747 (N_11747,N_11475,N_11529);
nor U11748 (N_11748,N_11633,N_11412);
nand U11749 (N_11749,N_11536,N_11639);
nand U11750 (N_11750,N_11578,N_11492);
or U11751 (N_11751,N_11671,N_11516);
and U11752 (N_11752,N_11521,N_11663);
nand U11753 (N_11753,N_11563,N_11603);
or U11754 (N_11754,N_11461,N_11668);
nand U11755 (N_11755,N_11687,N_11651);
and U11756 (N_11756,N_11456,N_11561);
nor U11757 (N_11757,N_11413,N_11511);
or U11758 (N_11758,N_11525,N_11416);
xnor U11759 (N_11759,N_11684,N_11469);
nor U11760 (N_11760,N_11676,N_11555);
xnor U11761 (N_11761,N_11677,N_11638);
and U11762 (N_11762,N_11417,N_11468);
nand U11763 (N_11763,N_11568,N_11405);
or U11764 (N_11764,N_11699,N_11491);
xnor U11765 (N_11765,N_11477,N_11444);
nand U11766 (N_11766,N_11484,N_11623);
xor U11767 (N_11767,N_11505,N_11466);
xor U11768 (N_11768,N_11602,N_11494);
xor U11769 (N_11769,N_11558,N_11616);
nor U11770 (N_11770,N_11421,N_11431);
or U11771 (N_11771,N_11429,N_11400);
and U11772 (N_11772,N_11457,N_11404);
or U11773 (N_11773,N_11473,N_11514);
xor U11774 (N_11774,N_11503,N_11497);
nor U11775 (N_11775,N_11443,N_11630);
nor U11776 (N_11776,N_11442,N_11609);
and U11777 (N_11777,N_11579,N_11523);
xor U11778 (N_11778,N_11571,N_11694);
or U11779 (N_11779,N_11560,N_11598);
xor U11780 (N_11780,N_11588,N_11595);
nor U11781 (N_11781,N_11528,N_11543);
and U11782 (N_11782,N_11647,N_11659);
or U11783 (N_11783,N_11617,N_11644);
nor U11784 (N_11784,N_11428,N_11645);
nand U11785 (N_11785,N_11488,N_11690);
nand U11786 (N_11786,N_11531,N_11445);
nand U11787 (N_11787,N_11537,N_11618);
xnor U11788 (N_11788,N_11527,N_11641);
or U11789 (N_11789,N_11518,N_11408);
xnor U11790 (N_11790,N_11530,N_11407);
or U11791 (N_11791,N_11544,N_11490);
nand U11792 (N_11792,N_11567,N_11679);
xnor U11793 (N_11793,N_11539,N_11611);
and U11794 (N_11794,N_11669,N_11452);
or U11795 (N_11795,N_11599,N_11697);
xnor U11796 (N_11796,N_11683,N_11447);
xnor U11797 (N_11797,N_11661,N_11589);
and U11798 (N_11798,N_11664,N_11569);
nor U11799 (N_11799,N_11479,N_11419);
or U11800 (N_11800,N_11450,N_11478);
or U11801 (N_11801,N_11583,N_11637);
xor U11802 (N_11802,N_11481,N_11562);
xor U11803 (N_11803,N_11581,N_11434);
nor U11804 (N_11804,N_11657,N_11554);
or U11805 (N_11805,N_11453,N_11471);
nand U11806 (N_11806,N_11689,N_11449);
and U11807 (N_11807,N_11535,N_11467);
xnor U11808 (N_11808,N_11585,N_11538);
or U11809 (N_11809,N_11552,N_11420);
xnor U11810 (N_11810,N_11520,N_11409);
nor U11811 (N_11811,N_11427,N_11607);
nand U11812 (N_11812,N_11670,N_11513);
or U11813 (N_11813,N_11650,N_11401);
and U11814 (N_11814,N_11624,N_11458);
and U11815 (N_11815,N_11672,N_11508);
xnor U11816 (N_11816,N_11629,N_11499);
and U11817 (N_11817,N_11570,N_11622);
or U11818 (N_11818,N_11634,N_11640);
nand U11819 (N_11819,N_11691,N_11436);
xor U11820 (N_11820,N_11591,N_11667);
nand U11821 (N_11821,N_11696,N_11486);
and U11822 (N_11822,N_11614,N_11465);
or U11823 (N_11823,N_11485,N_11665);
or U11824 (N_11824,N_11620,N_11500);
nor U11825 (N_11825,N_11587,N_11615);
xnor U11826 (N_11826,N_11582,N_11681);
nand U11827 (N_11827,N_11448,N_11474);
xor U11828 (N_11828,N_11564,N_11430);
and U11829 (N_11829,N_11415,N_11577);
nand U11830 (N_11830,N_11423,N_11643);
xnor U11831 (N_11831,N_11403,N_11686);
or U11832 (N_11832,N_11613,N_11605);
and U11833 (N_11833,N_11510,N_11507);
or U11834 (N_11834,N_11636,N_11411);
nand U11835 (N_11835,N_11472,N_11512);
or U11836 (N_11836,N_11646,N_11675);
xor U11837 (N_11837,N_11655,N_11439);
nor U11838 (N_11838,N_11597,N_11660);
xnor U11839 (N_11839,N_11470,N_11674);
xor U11840 (N_11840,N_11656,N_11604);
and U11841 (N_11841,N_11533,N_11632);
nand U11842 (N_11842,N_11438,N_11418);
xnor U11843 (N_11843,N_11480,N_11406);
xnor U11844 (N_11844,N_11682,N_11425);
nand U11845 (N_11845,N_11601,N_11498);
or U11846 (N_11846,N_11608,N_11586);
and U11847 (N_11847,N_11463,N_11459);
xnor U11848 (N_11848,N_11631,N_11573);
nor U11849 (N_11849,N_11621,N_11451);
nor U11850 (N_11850,N_11410,N_11697);
and U11851 (N_11851,N_11664,N_11570);
xor U11852 (N_11852,N_11422,N_11443);
and U11853 (N_11853,N_11671,N_11672);
or U11854 (N_11854,N_11578,N_11630);
xnor U11855 (N_11855,N_11542,N_11482);
and U11856 (N_11856,N_11655,N_11446);
or U11857 (N_11857,N_11419,N_11565);
xor U11858 (N_11858,N_11426,N_11638);
xnor U11859 (N_11859,N_11514,N_11557);
nor U11860 (N_11860,N_11597,N_11530);
and U11861 (N_11861,N_11461,N_11655);
and U11862 (N_11862,N_11401,N_11413);
xor U11863 (N_11863,N_11617,N_11666);
or U11864 (N_11864,N_11472,N_11639);
nor U11865 (N_11865,N_11655,N_11478);
nand U11866 (N_11866,N_11494,N_11620);
or U11867 (N_11867,N_11617,N_11475);
nor U11868 (N_11868,N_11487,N_11663);
xor U11869 (N_11869,N_11630,N_11626);
and U11870 (N_11870,N_11613,N_11565);
xor U11871 (N_11871,N_11467,N_11409);
nand U11872 (N_11872,N_11676,N_11451);
or U11873 (N_11873,N_11641,N_11473);
and U11874 (N_11874,N_11490,N_11475);
nand U11875 (N_11875,N_11602,N_11627);
nor U11876 (N_11876,N_11642,N_11684);
and U11877 (N_11877,N_11577,N_11684);
or U11878 (N_11878,N_11634,N_11642);
xnor U11879 (N_11879,N_11691,N_11683);
or U11880 (N_11880,N_11501,N_11619);
nand U11881 (N_11881,N_11535,N_11572);
or U11882 (N_11882,N_11461,N_11455);
or U11883 (N_11883,N_11595,N_11458);
and U11884 (N_11884,N_11661,N_11448);
nor U11885 (N_11885,N_11414,N_11415);
or U11886 (N_11886,N_11658,N_11405);
nor U11887 (N_11887,N_11545,N_11640);
nor U11888 (N_11888,N_11535,N_11411);
nand U11889 (N_11889,N_11442,N_11563);
xnor U11890 (N_11890,N_11606,N_11417);
nand U11891 (N_11891,N_11666,N_11425);
nand U11892 (N_11892,N_11481,N_11565);
xnor U11893 (N_11893,N_11561,N_11683);
nor U11894 (N_11894,N_11656,N_11568);
and U11895 (N_11895,N_11619,N_11657);
nand U11896 (N_11896,N_11415,N_11402);
and U11897 (N_11897,N_11586,N_11632);
or U11898 (N_11898,N_11643,N_11420);
nor U11899 (N_11899,N_11406,N_11632);
xnor U11900 (N_11900,N_11629,N_11642);
xnor U11901 (N_11901,N_11523,N_11455);
or U11902 (N_11902,N_11600,N_11405);
nand U11903 (N_11903,N_11504,N_11589);
nor U11904 (N_11904,N_11431,N_11658);
and U11905 (N_11905,N_11545,N_11611);
nor U11906 (N_11906,N_11433,N_11684);
and U11907 (N_11907,N_11430,N_11460);
nor U11908 (N_11908,N_11691,N_11686);
and U11909 (N_11909,N_11462,N_11400);
nor U11910 (N_11910,N_11472,N_11407);
or U11911 (N_11911,N_11662,N_11606);
and U11912 (N_11912,N_11613,N_11558);
and U11913 (N_11913,N_11619,N_11429);
nor U11914 (N_11914,N_11424,N_11570);
nand U11915 (N_11915,N_11470,N_11512);
nand U11916 (N_11916,N_11577,N_11576);
xnor U11917 (N_11917,N_11583,N_11534);
nand U11918 (N_11918,N_11623,N_11403);
nand U11919 (N_11919,N_11575,N_11524);
or U11920 (N_11920,N_11539,N_11661);
or U11921 (N_11921,N_11690,N_11689);
or U11922 (N_11922,N_11498,N_11629);
xnor U11923 (N_11923,N_11568,N_11544);
nand U11924 (N_11924,N_11561,N_11443);
and U11925 (N_11925,N_11667,N_11534);
or U11926 (N_11926,N_11629,N_11666);
or U11927 (N_11927,N_11563,N_11525);
and U11928 (N_11928,N_11613,N_11651);
xor U11929 (N_11929,N_11575,N_11680);
and U11930 (N_11930,N_11400,N_11503);
or U11931 (N_11931,N_11656,N_11419);
nand U11932 (N_11932,N_11607,N_11518);
nand U11933 (N_11933,N_11465,N_11632);
nand U11934 (N_11934,N_11495,N_11506);
or U11935 (N_11935,N_11617,N_11581);
nand U11936 (N_11936,N_11651,N_11565);
nand U11937 (N_11937,N_11670,N_11688);
or U11938 (N_11938,N_11602,N_11514);
and U11939 (N_11939,N_11582,N_11673);
xnor U11940 (N_11940,N_11479,N_11640);
nand U11941 (N_11941,N_11538,N_11572);
nand U11942 (N_11942,N_11491,N_11473);
nand U11943 (N_11943,N_11653,N_11411);
and U11944 (N_11944,N_11473,N_11442);
and U11945 (N_11945,N_11481,N_11424);
xnor U11946 (N_11946,N_11589,N_11580);
nand U11947 (N_11947,N_11628,N_11445);
or U11948 (N_11948,N_11560,N_11406);
nand U11949 (N_11949,N_11448,N_11410);
nor U11950 (N_11950,N_11632,N_11463);
nor U11951 (N_11951,N_11417,N_11477);
and U11952 (N_11952,N_11632,N_11426);
nor U11953 (N_11953,N_11619,N_11559);
nor U11954 (N_11954,N_11424,N_11446);
xnor U11955 (N_11955,N_11516,N_11692);
or U11956 (N_11956,N_11441,N_11506);
nand U11957 (N_11957,N_11643,N_11609);
nor U11958 (N_11958,N_11527,N_11617);
or U11959 (N_11959,N_11490,N_11585);
xnor U11960 (N_11960,N_11675,N_11491);
xnor U11961 (N_11961,N_11510,N_11435);
xnor U11962 (N_11962,N_11494,N_11509);
or U11963 (N_11963,N_11478,N_11555);
and U11964 (N_11964,N_11574,N_11674);
nand U11965 (N_11965,N_11640,N_11476);
and U11966 (N_11966,N_11483,N_11467);
and U11967 (N_11967,N_11410,N_11654);
nor U11968 (N_11968,N_11468,N_11529);
nand U11969 (N_11969,N_11452,N_11661);
xor U11970 (N_11970,N_11680,N_11469);
xnor U11971 (N_11971,N_11662,N_11695);
nand U11972 (N_11972,N_11554,N_11475);
and U11973 (N_11973,N_11429,N_11531);
nand U11974 (N_11974,N_11565,N_11633);
xnor U11975 (N_11975,N_11417,N_11506);
and U11976 (N_11976,N_11479,N_11630);
nand U11977 (N_11977,N_11448,N_11458);
xnor U11978 (N_11978,N_11496,N_11624);
nor U11979 (N_11979,N_11607,N_11484);
and U11980 (N_11980,N_11485,N_11427);
and U11981 (N_11981,N_11476,N_11622);
or U11982 (N_11982,N_11586,N_11571);
or U11983 (N_11983,N_11654,N_11605);
or U11984 (N_11984,N_11663,N_11488);
nor U11985 (N_11985,N_11663,N_11584);
nand U11986 (N_11986,N_11693,N_11622);
nand U11987 (N_11987,N_11628,N_11651);
xnor U11988 (N_11988,N_11585,N_11646);
nand U11989 (N_11989,N_11487,N_11668);
or U11990 (N_11990,N_11691,N_11560);
or U11991 (N_11991,N_11411,N_11663);
xnor U11992 (N_11992,N_11421,N_11434);
or U11993 (N_11993,N_11516,N_11666);
or U11994 (N_11994,N_11495,N_11436);
xnor U11995 (N_11995,N_11534,N_11483);
and U11996 (N_11996,N_11470,N_11453);
nor U11997 (N_11997,N_11580,N_11475);
and U11998 (N_11998,N_11610,N_11410);
nand U11999 (N_11999,N_11514,N_11580);
nand U12000 (N_12000,N_11919,N_11880);
and U12001 (N_12001,N_11837,N_11759);
or U12002 (N_12002,N_11765,N_11995);
and U12003 (N_12003,N_11928,N_11804);
nor U12004 (N_12004,N_11879,N_11877);
nand U12005 (N_12005,N_11772,N_11985);
xnor U12006 (N_12006,N_11706,N_11718);
and U12007 (N_12007,N_11813,N_11744);
or U12008 (N_12008,N_11730,N_11974);
nor U12009 (N_12009,N_11956,N_11717);
nor U12010 (N_12010,N_11723,N_11904);
nand U12011 (N_12011,N_11854,N_11705);
xnor U12012 (N_12012,N_11917,N_11777);
nor U12013 (N_12013,N_11859,N_11841);
nor U12014 (N_12014,N_11756,N_11794);
nand U12015 (N_12015,N_11967,N_11834);
and U12016 (N_12016,N_11884,N_11999);
nor U12017 (N_12017,N_11910,N_11832);
nand U12018 (N_12018,N_11865,N_11779);
xnor U12019 (N_12019,N_11932,N_11811);
and U12020 (N_12020,N_11856,N_11761);
nand U12021 (N_12021,N_11711,N_11736);
nor U12022 (N_12022,N_11805,N_11776);
nand U12023 (N_12023,N_11826,N_11943);
and U12024 (N_12024,N_11984,N_11975);
nand U12025 (N_12025,N_11857,N_11762);
or U12026 (N_12026,N_11976,N_11861);
and U12027 (N_12027,N_11712,N_11864);
and U12028 (N_12028,N_11977,N_11838);
xnor U12029 (N_12029,N_11815,N_11728);
and U12030 (N_12030,N_11710,N_11828);
nor U12031 (N_12031,N_11923,N_11930);
xnor U12032 (N_12032,N_11862,N_11790);
nor U12033 (N_12033,N_11979,N_11781);
and U12034 (N_12034,N_11746,N_11969);
nor U12035 (N_12035,N_11822,N_11853);
xnor U12036 (N_12036,N_11780,N_11793);
or U12037 (N_12037,N_11770,N_11849);
xnor U12038 (N_12038,N_11745,N_11949);
xnor U12039 (N_12039,N_11876,N_11993);
nand U12040 (N_12040,N_11972,N_11818);
nor U12041 (N_12041,N_11725,N_11959);
nand U12042 (N_12042,N_11885,N_11992);
nor U12043 (N_12043,N_11960,N_11792);
and U12044 (N_12044,N_11986,N_11817);
nand U12045 (N_12045,N_11931,N_11807);
xor U12046 (N_12046,N_11878,N_11937);
and U12047 (N_12047,N_11737,N_11897);
xnor U12048 (N_12048,N_11748,N_11795);
and U12049 (N_12049,N_11741,N_11947);
xnor U12050 (N_12050,N_11842,N_11808);
nor U12051 (N_12051,N_11866,N_11901);
and U12052 (N_12052,N_11767,N_11982);
nor U12053 (N_12053,N_11915,N_11708);
and U12054 (N_12054,N_11913,N_11830);
xnor U12055 (N_12055,N_11774,N_11890);
nand U12056 (N_12056,N_11755,N_11800);
nor U12057 (N_12057,N_11952,N_11852);
xor U12058 (N_12058,N_11988,N_11844);
nand U12059 (N_12059,N_11860,N_11953);
nand U12060 (N_12060,N_11806,N_11843);
xor U12061 (N_12061,N_11700,N_11934);
nor U12062 (N_12062,N_11751,N_11942);
nand U12063 (N_12063,N_11820,N_11922);
nand U12064 (N_12064,N_11905,N_11875);
nand U12065 (N_12065,N_11733,N_11791);
or U12066 (N_12066,N_11933,N_11892);
and U12067 (N_12067,N_11929,N_11749);
nand U12068 (N_12068,N_11920,N_11720);
nor U12069 (N_12069,N_11824,N_11734);
xor U12070 (N_12070,N_11991,N_11978);
nor U12071 (N_12071,N_11889,N_11845);
and U12072 (N_12072,N_11764,N_11958);
nor U12073 (N_12073,N_11742,N_11768);
nand U12074 (N_12074,N_11703,N_11850);
xnor U12075 (N_12075,N_11848,N_11716);
and U12076 (N_12076,N_11753,N_11927);
nand U12077 (N_12077,N_11970,N_11973);
and U12078 (N_12078,N_11938,N_11945);
xor U12079 (N_12079,N_11738,N_11722);
nor U12080 (N_12080,N_11964,N_11758);
nand U12081 (N_12081,N_11729,N_11771);
nor U12082 (N_12082,N_11788,N_11916);
and U12083 (N_12083,N_11951,N_11874);
or U12084 (N_12084,N_11810,N_11921);
nand U12085 (N_12085,N_11996,N_11990);
or U12086 (N_12086,N_11721,N_11833);
nand U12087 (N_12087,N_11763,N_11957);
nor U12088 (N_12088,N_11769,N_11819);
and U12089 (N_12089,N_11909,N_11714);
nor U12090 (N_12090,N_11831,N_11903);
nand U12091 (N_12091,N_11871,N_11707);
xnor U12092 (N_12092,N_11882,N_11899);
and U12093 (N_12093,N_11719,N_11987);
or U12094 (N_12094,N_11896,N_11887);
and U12095 (N_12095,N_11925,N_11908);
xnor U12096 (N_12096,N_11918,N_11911);
and U12097 (N_12097,N_11963,N_11981);
nor U12098 (N_12098,N_11912,N_11868);
nand U12099 (N_12099,N_11731,N_11935);
and U12100 (N_12100,N_11840,N_11778);
nor U12101 (N_12101,N_11702,N_11948);
xor U12102 (N_12102,N_11914,N_11962);
and U12103 (N_12103,N_11786,N_11907);
nor U12104 (N_12104,N_11869,N_11883);
or U12105 (N_12105,N_11829,N_11825);
and U12106 (N_12106,N_11735,N_11814);
and U12107 (N_12107,N_11867,N_11750);
or U12108 (N_12108,N_11863,N_11966);
nor U12109 (N_12109,N_11802,N_11936);
nor U12110 (N_12110,N_11946,N_11858);
nor U12111 (N_12111,N_11747,N_11739);
or U12112 (N_12112,N_11809,N_11855);
nand U12113 (N_12113,N_11839,N_11950);
nor U12114 (N_12114,N_11752,N_11941);
nand U12115 (N_12115,N_11939,N_11796);
xor U12116 (N_12116,N_11881,N_11872);
or U12117 (N_12117,N_11989,N_11726);
nand U12118 (N_12118,N_11955,N_11965);
xnor U12119 (N_12119,N_11799,N_11783);
xnor U12120 (N_12120,N_11900,N_11998);
nor U12121 (N_12121,N_11732,N_11954);
or U12122 (N_12122,N_11798,N_11983);
xnor U12123 (N_12123,N_11847,N_11787);
nand U12124 (N_12124,N_11902,N_11926);
or U12125 (N_12125,N_11961,N_11797);
or U12126 (N_12126,N_11968,N_11784);
nor U12127 (N_12127,N_11835,N_11766);
xnor U12128 (N_12128,N_11827,N_11715);
and U12129 (N_12129,N_11823,N_11944);
nor U12130 (N_12130,N_11836,N_11870);
xor U12131 (N_12131,N_11851,N_11727);
and U12132 (N_12132,N_11886,N_11775);
nor U12133 (N_12133,N_11701,N_11980);
and U12134 (N_12134,N_11906,N_11894);
and U12135 (N_12135,N_11789,N_11704);
xor U12136 (N_12136,N_11740,N_11803);
xor U12137 (N_12137,N_11801,N_11782);
or U12138 (N_12138,N_11757,N_11713);
and U12139 (N_12139,N_11760,N_11893);
nor U12140 (N_12140,N_11895,N_11997);
and U12141 (N_12141,N_11971,N_11891);
or U12142 (N_12142,N_11773,N_11821);
or U12143 (N_12143,N_11846,N_11816);
nand U12144 (N_12144,N_11724,N_11709);
nor U12145 (N_12145,N_11940,N_11785);
and U12146 (N_12146,N_11888,N_11743);
and U12147 (N_12147,N_11754,N_11898);
and U12148 (N_12148,N_11873,N_11924);
and U12149 (N_12149,N_11812,N_11994);
nor U12150 (N_12150,N_11713,N_11933);
xnor U12151 (N_12151,N_11757,N_11813);
or U12152 (N_12152,N_11887,N_11889);
or U12153 (N_12153,N_11965,N_11741);
xnor U12154 (N_12154,N_11760,N_11955);
nand U12155 (N_12155,N_11755,N_11745);
nand U12156 (N_12156,N_11952,N_11979);
and U12157 (N_12157,N_11747,N_11807);
nand U12158 (N_12158,N_11909,N_11757);
xnor U12159 (N_12159,N_11830,N_11739);
or U12160 (N_12160,N_11719,N_11958);
nor U12161 (N_12161,N_11712,N_11756);
or U12162 (N_12162,N_11742,N_11931);
or U12163 (N_12163,N_11904,N_11796);
nor U12164 (N_12164,N_11773,N_11952);
xor U12165 (N_12165,N_11874,N_11742);
nor U12166 (N_12166,N_11909,N_11974);
or U12167 (N_12167,N_11879,N_11733);
nand U12168 (N_12168,N_11966,N_11780);
nand U12169 (N_12169,N_11811,N_11930);
or U12170 (N_12170,N_11747,N_11722);
or U12171 (N_12171,N_11733,N_11704);
or U12172 (N_12172,N_11958,N_11979);
and U12173 (N_12173,N_11813,N_11947);
nand U12174 (N_12174,N_11921,N_11755);
nor U12175 (N_12175,N_11793,N_11770);
and U12176 (N_12176,N_11710,N_11939);
xnor U12177 (N_12177,N_11914,N_11846);
and U12178 (N_12178,N_11846,N_11856);
or U12179 (N_12179,N_11939,N_11944);
xnor U12180 (N_12180,N_11924,N_11998);
nand U12181 (N_12181,N_11835,N_11978);
nand U12182 (N_12182,N_11899,N_11812);
nand U12183 (N_12183,N_11810,N_11911);
nor U12184 (N_12184,N_11804,N_11955);
nand U12185 (N_12185,N_11807,N_11866);
nand U12186 (N_12186,N_11920,N_11933);
or U12187 (N_12187,N_11846,N_11872);
and U12188 (N_12188,N_11863,N_11890);
nor U12189 (N_12189,N_11889,N_11950);
or U12190 (N_12190,N_11809,N_11959);
nand U12191 (N_12191,N_11775,N_11885);
nor U12192 (N_12192,N_11971,N_11785);
xor U12193 (N_12193,N_11943,N_11991);
nand U12194 (N_12194,N_11814,N_11959);
or U12195 (N_12195,N_11737,N_11703);
and U12196 (N_12196,N_11815,N_11790);
xnor U12197 (N_12197,N_11781,N_11763);
nand U12198 (N_12198,N_11707,N_11824);
xnor U12199 (N_12199,N_11794,N_11739);
or U12200 (N_12200,N_11807,N_11839);
nand U12201 (N_12201,N_11737,N_11781);
and U12202 (N_12202,N_11703,N_11989);
or U12203 (N_12203,N_11957,N_11943);
nor U12204 (N_12204,N_11969,N_11894);
xnor U12205 (N_12205,N_11800,N_11714);
nand U12206 (N_12206,N_11896,N_11814);
or U12207 (N_12207,N_11994,N_11852);
or U12208 (N_12208,N_11806,N_11756);
nand U12209 (N_12209,N_11809,N_11997);
nor U12210 (N_12210,N_11825,N_11888);
nor U12211 (N_12211,N_11729,N_11966);
and U12212 (N_12212,N_11839,N_11796);
or U12213 (N_12213,N_11862,N_11766);
nor U12214 (N_12214,N_11934,N_11844);
xnor U12215 (N_12215,N_11782,N_11838);
or U12216 (N_12216,N_11960,N_11703);
and U12217 (N_12217,N_11982,N_11934);
and U12218 (N_12218,N_11735,N_11897);
or U12219 (N_12219,N_11757,N_11868);
xor U12220 (N_12220,N_11904,N_11852);
nor U12221 (N_12221,N_11916,N_11747);
nand U12222 (N_12222,N_11882,N_11773);
xnor U12223 (N_12223,N_11900,N_11972);
xor U12224 (N_12224,N_11804,N_11789);
nor U12225 (N_12225,N_11769,N_11864);
or U12226 (N_12226,N_11941,N_11732);
and U12227 (N_12227,N_11798,N_11741);
nand U12228 (N_12228,N_11718,N_11897);
nand U12229 (N_12229,N_11804,N_11959);
and U12230 (N_12230,N_11937,N_11897);
and U12231 (N_12231,N_11824,N_11916);
xor U12232 (N_12232,N_11777,N_11852);
xnor U12233 (N_12233,N_11894,N_11874);
or U12234 (N_12234,N_11789,N_11963);
or U12235 (N_12235,N_11874,N_11924);
nand U12236 (N_12236,N_11749,N_11719);
nand U12237 (N_12237,N_11936,N_11754);
nor U12238 (N_12238,N_11875,N_11959);
xor U12239 (N_12239,N_11847,N_11854);
and U12240 (N_12240,N_11705,N_11832);
or U12241 (N_12241,N_11759,N_11980);
nor U12242 (N_12242,N_11813,N_11789);
and U12243 (N_12243,N_11719,N_11838);
nor U12244 (N_12244,N_11744,N_11812);
nor U12245 (N_12245,N_11897,N_11732);
nor U12246 (N_12246,N_11913,N_11719);
nor U12247 (N_12247,N_11701,N_11870);
and U12248 (N_12248,N_11701,N_11936);
nor U12249 (N_12249,N_11750,N_11809);
nor U12250 (N_12250,N_11701,N_11741);
nand U12251 (N_12251,N_11903,N_11962);
or U12252 (N_12252,N_11811,N_11915);
nand U12253 (N_12253,N_11905,N_11839);
nor U12254 (N_12254,N_11831,N_11897);
nand U12255 (N_12255,N_11858,N_11708);
or U12256 (N_12256,N_11820,N_11790);
or U12257 (N_12257,N_11821,N_11917);
nand U12258 (N_12258,N_11960,N_11818);
and U12259 (N_12259,N_11914,N_11986);
and U12260 (N_12260,N_11706,N_11997);
and U12261 (N_12261,N_11750,N_11978);
or U12262 (N_12262,N_11810,N_11718);
or U12263 (N_12263,N_11959,N_11891);
xnor U12264 (N_12264,N_11776,N_11730);
nand U12265 (N_12265,N_11998,N_11768);
nor U12266 (N_12266,N_11866,N_11984);
and U12267 (N_12267,N_11847,N_11969);
and U12268 (N_12268,N_11809,N_11905);
nand U12269 (N_12269,N_11853,N_11733);
nor U12270 (N_12270,N_11736,N_11728);
and U12271 (N_12271,N_11829,N_11821);
nor U12272 (N_12272,N_11846,N_11912);
nand U12273 (N_12273,N_11938,N_11887);
nor U12274 (N_12274,N_11820,N_11856);
or U12275 (N_12275,N_11749,N_11827);
nor U12276 (N_12276,N_11770,N_11763);
nand U12277 (N_12277,N_11963,N_11912);
nand U12278 (N_12278,N_11970,N_11935);
or U12279 (N_12279,N_11868,N_11973);
nor U12280 (N_12280,N_11711,N_11932);
and U12281 (N_12281,N_11861,N_11719);
nor U12282 (N_12282,N_11810,N_11855);
or U12283 (N_12283,N_11800,N_11826);
and U12284 (N_12284,N_11824,N_11944);
and U12285 (N_12285,N_11981,N_11955);
nor U12286 (N_12286,N_11860,N_11956);
and U12287 (N_12287,N_11900,N_11802);
nand U12288 (N_12288,N_11756,N_11852);
nand U12289 (N_12289,N_11977,N_11832);
nand U12290 (N_12290,N_11768,N_11849);
xnor U12291 (N_12291,N_11982,N_11793);
nand U12292 (N_12292,N_11922,N_11723);
nand U12293 (N_12293,N_11771,N_11857);
nor U12294 (N_12294,N_11838,N_11956);
nor U12295 (N_12295,N_11929,N_11882);
or U12296 (N_12296,N_11735,N_11969);
xnor U12297 (N_12297,N_11729,N_11727);
and U12298 (N_12298,N_11795,N_11765);
nand U12299 (N_12299,N_11801,N_11832);
or U12300 (N_12300,N_12234,N_12052);
and U12301 (N_12301,N_12231,N_12202);
nand U12302 (N_12302,N_12181,N_12046);
nor U12303 (N_12303,N_12049,N_12008);
nand U12304 (N_12304,N_12289,N_12056);
xor U12305 (N_12305,N_12042,N_12237);
nor U12306 (N_12306,N_12146,N_12028);
nor U12307 (N_12307,N_12216,N_12058);
nor U12308 (N_12308,N_12043,N_12064);
xor U12309 (N_12309,N_12271,N_12149);
or U12310 (N_12310,N_12014,N_12243);
xor U12311 (N_12311,N_12118,N_12245);
nor U12312 (N_12312,N_12195,N_12132);
xnor U12313 (N_12313,N_12179,N_12018);
xor U12314 (N_12314,N_12083,N_12148);
nand U12315 (N_12315,N_12189,N_12062);
or U12316 (N_12316,N_12205,N_12248);
and U12317 (N_12317,N_12044,N_12225);
and U12318 (N_12318,N_12136,N_12096);
xnor U12319 (N_12319,N_12178,N_12298);
nand U12320 (N_12320,N_12113,N_12278);
and U12321 (N_12321,N_12280,N_12218);
nand U12322 (N_12322,N_12254,N_12251);
and U12323 (N_12323,N_12232,N_12286);
or U12324 (N_12324,N_12077,N_12228);
and U12325 (N_12325,N_12107,N_12025);
xor U12326 (N_12326,N_12168,N_12033);
nor U12327 (N_12327,N_12227,N_12082);
xnor U12328 (N_12328,N_12264,N_12050);
xnor U12329 (N_12329,N_12021,N_12063);
nand U12330 (N_12330,N_12172,N_12000);
nor U12331 (N_12331,N_12193,N_12102);
or U12332 (N_12332,N_12069,N_12079);
or U12333 (N_12333,N_12258,N_12210);
xor U12334 (N_12334,N_12233,N_12104);
and U12335 (N_12335,N_12284,N_12186);
and U12336 (N_12336,N_12017,N_12203);
and U12337 (N_12337,N_12217,N_12045);
nand U12338 (N_12338,N_12222,N_12260);
nand U12339 (N_12339,N_12273,N_12122);
nor U12340 (N_12340,N_12097,N_12282);
and U12341 (N_12341,N_12038,N_12211);
nand U12342 (N_12342,N_12139,N_12229);
and U12343 (N_12343,N_12117,N_12263);
or U12344 (N_12344,N_12199,N_12295);
and U12345 (N_12345,N_12085,N_12027);
or U12346 (N_12346,N_12037,N_12007);
xnor U12347 (N_12347,N_12110,N_12130);
nor U12348 (N_12348,N_12268,N_12125);
and U12349 (N_12349,N_12170,N_12187);
nor U12350 (N_12350,N_12004,N_12214);
nor U12351 (N_12351,N_12005,N_12240);
nor U12352 (N_12352,N_12200,N_12274);
nor U12353 (N_12353,N_12212,N_12283);
nor U12354 (N_12354,N_12088,N_12140);
and U12355 (N_12355,N_12030,N_12105);
xor U12356 (N_12356,N_12055,N_12003);
nor U12357 (N_12357,N_12215,N_12023);
nor U12358 (N_12358,N_12279,N_12171);
and U12359 (N_12359,N_12092,N_12255);
nor U12360 (N_12360,N_12256,N_12031);
and U12361 (N_12361,N_12126,N_12197);
nand U12362 (N_12362,N_12169,N_12120);
or U12363 (N_12363,N_12142,N_12154);
xnor U12364 (N_12364,N_12138,N_12124);
and U12365 (N_12365,N_12164,N_12059);
or U12366 (N_12366,N_12161,N_12272);
nand U12367 (N_12367,N_12269,N_12065);
nand U12368 (N_12368,N_12297,N_12158);
nand U12369 (N_12369,N_12127,N_12134);
nand U12370 (N_12370,N_12155,N_12277);
and U12371 (N_12371,N_12247,N_12198);
nand U12372 (N_12372,N_12119,N_12048);
nand U12373 (N_12373,N_12188,N_12201);
nor U12374 (N_12374,N_12246,N_12292);
nand U12375 (N_12375,N_12133,N_12241);
nand U12376 (N_12376,N_12177,N_12001);
nor U12377 (N_12377,N_12180,N_12144);
and U12378 (N_12378,N_12294,N_12054);
nand U12379 (N_12379,N_12147,N_12039);
or U12380 (N_12380,N_12173,N_12115);
or U12381 (N_12381,N_12236,N_12242);
or U12382 (N_12382,N_12190,N_12160);
and U12383 (N_12383,N_12207,N_12143);
xor U12384 (N_12384,N_12182,N_12265);
and U12385 (N_12385,N_12275,N_12116);
xor U12386 (N_12386,N_12047,N_12219);
xor U12387 (N_12387,N_12296,N_12267);
xor U12388 (N_12388,N_12076,N_12192);
or U12389 (N_12389,N_12183,N_12270);
nor U12390 (N_12390,N_12066,N_12253);
nor U12391 (N_12391,N_12016,N_12184);
nand U12392 (N_12392,N_12262,N_12153);
xnor U12393 (N_12393,N_12165,N_12167);
and U12394 (N_12394,N_12250,N_12226);
xor U12395 (N_12395,N_12121,N_12108);
xnor U12396 (N_12396,N_12206,N_12159);
xor U12397 (N_12397,N_12093,N_12141);
or U12398 (N_12398,N_12091,N_12029);
xnor U12399 (N_12399,N_12224,N_12162);
xor U12400 (N_12400,N_12145,N_12061);
xnor U12401 (N_12401,N_12087,N_12259);
and U12402 (N_12402,N_12002,N_12261);
xnor U12403 (N_12403,N_12191,N_12128);
or U12404 (N_12404,N_12239,N_12244);
xor U12405 (N_12405,N_12230,N_12078);
nor U12406 (N_12406,N_12137,N_12213);
nand U12407 (N_12407,N_12081,N_12106);
nor U12408 (N_12408,N_12026,N_12011);
and U12409 (N_12409,N_12114,N_12015);
or U12410 (N_12410,N_12094,N_12035);
nor U12411 (N_12411,N_12073,N_12086);
nand U12412 (N_12412,N_12013,N_12156);
or U12413 (N_12413,N_12006,N_12157);
nor U12414 (N_12414,N_12075,N_12131);
or U12415 (N_12415,N_12223,N_12204);
xor U12416 (N_12416,N_12287,N_12101);
xor U12417 (N_12417,N_12070,N_12009);
or U12418 (N_12418,N_12238,N_12024);
nand U12419 (N_12419,N_12266,N_12185);
and U12420 (N_12420,N_12068,N_12020);
xor U12421 (N_12421,N_12196,N_12285);
nor U12422 (N_12422,N_12293,N_12067);
and U12423 (N_12423,N_12041,N_12053);
nand U12424 (N_12424,N_12209,N_12249);
nand U12425 (N_12425,N_12099,N_12123);
nor U12426 (N_12426,N_12135,N_12150);
or U12427 (N_12427,N_12022,N_12257);
nor U12428 (N_12428,N_12290,N_12276);
nand U12429 (N_12429,N_12084,N_12089);
or U12430 (N_12430,N_12072,N_12152);
and U12431 (N_12431,N_12220,N_12111);
and U12432 (N_12432,N_12112,N_12299);
nor U12433 (N_12433,N_12032,N_12151);
xor U12434 (N_12434,N_12090,N_12100);
nand U12435 (N_12435,N_12010,N_12175);
or U12436 (N_12436,N_12034,N_12166);
nand U12437 (N_12437,N_12163,N_12051);
nor U12438 (N_12438,N_12036,N_12176);
or U12439 (N_12439,N_12098,N_12019);
nor U12440 (N_12440,N_12040,N_12074);
nand U12441 (N_12441,N_12103,N_12281);
nand U12442 (N_12442,N_12129,N_12012);
nand U12443 (N_12443,N_12194,N_12288);
nor U12444 (N_12444,N_12252,N_12095);
nor U12445 (N_12445,N_12071,N_12080);
nor U12446 (N_12446,N_12221,N_12057);
xnor U12447 (N_12447,N_12291,N_12235);
nor U12448 (N_12448,N_12060,N_12208);
nand U12449 (N_12449,N_12174,N_12109);
nor U12450 (N_12450,N_12023,N_12136);
and U12451 (N_12451,N_12287,N_12031);
xnor U12452 (N_12452,N_12165,N_12123);
and U12453 (N_12453,N_12231,N_12270);
and U12454 (N_12454,N_12012,N_12143);
nand U12455 (N_12455,N_12282,N_12187);
and U12456 (N_12456,N_12059,N_12100);
and U12457 (N_12457,N_12183,N_12268);
xnor U12458 (N_12458,N_12160,N_12221);
and U12459 (N_12459,N_12258,N_12097);
and U12460 (N_12460,N_12127,N_12012);
nor U12461 (N_12461,N_12030,N_12236);
nand U12462 (N_12462,N_12128,N_12101);
nand U12463 (N_12463,N_12220,N_12078);
and U12464 (N_12464,N_12175,N_12178);
or U12465 (N_12465,N_12165,N_12094);
and U12466 (N_12466,N_12128,N_12248);
nand U12467 (N_12467,N_12249,N_12288);
xor U12468 (N_12468,N_12187,N_12154);
or U12469 (N_12469,N_12080,N_12134);
nand U12470 (N_12470,N_12162,N_12133);
and U12471 (N_12471,N_12053,N_12048);
xnor U12472 (N_12472,N_12224,N_12074);
and U12473 (N_12473,N_12272,N_12108);
nor U12474 (N_12474,N_12163,N_12244);
or U12475 (N_12475,N_12158,N_12124);
or U12476 (N_12476,N_12183,N_12195);
nor U12477 (N_12477,N_12097,N_12250);
nand U12478 (N_12478,N_12240,N_12231);
nand U12479 (N_12479,N_12026,N_12237);
nand U12480 (N_12480,N_12136,N_12197);
nor U12481 (N_12481,N_12106,N_12090);
nand U12482 (N_12482,N_12083,N_12177);
and U12483 (N_12483,N_12086,N_12192);
and U12484 (N_12484,N_12142,N_12019);
or U12485 (N_12485,N_12075,N_12168);
nor U12486 (N_12486,N_12285,N_12157);
xor U12487 (N_12487,N_12190,N_12256);
xnor U12488 (N_12488,N_12235,N_12116);
nor U12489 (N_12489,N_12200,N_12248);
and U12490 (N_12490,N_12223,N_12093);
xor U12491 (N_12491,N_12183,N_12225);
xnor U12492 (N_12492,N_12274,N_12089);
and U12493 (N_12493,N_12216,N_12160);
nor U12494 (N_12494,N_12030,N_12009);
nor U12495 (N_12495,N_12188,N_12145);
or U12496 (N_12496,N_12247,N_12053);
xor U12497 (N_12497,N_12049,N_12155);
or U12498 (N_12498,N_12105,N_12061);
or U12499 (N_12499,N_12214,N_12273);
and U12500 (N_12500,N_12044,N_12210);
and U12501 (N_12501,N_12194,N_12068);
and U12502 (N_12502,N_12015,N_12156);
nor U12503 (N_12503,N_12013,N_12059);
and U12504 (N_12504,N_12249,N_12167);
xnor U12505 (N_12505,N_12008,N_12070);
nor U12506 (N_12506,N_12091,N_12125);
xor U12507 (N_12507,N_12249,N_12143);
nand U12508 (N_12508,N_12080,N_12246);
nand U12509 (N_12509,N_12020,N_12058);
and U12510 (N_12510,N_12121,N_12050);
and U12511 (N_12511,N_12298,N_12156);
nor U12512 (N_12512,N_12198,N_12013);
and U12513 (N_12513,N_12060,N_12137);
nand U12514 (N_12514,N_12060,N_12168);
or U12515 (N_12515,N_12255,N_12190);
or U12516 (N_12516,N_12035,N_12202);
and U12517 (N_12517,N_12032,N_12178);
xor U12518 (N_12518,N_12063,N_12136);
and U12519 (N_12519,N_12247,N_12021);
xnor U12520 (N_12520,N_12134,N_12280);
nor U12521 (N_12521,N_12015,N_12049);
or U12522 (N_12522,N_12233,N_12062);
and U12523 (N_12523,N_12085,N_12060);
nand U12524 (N_12524,N_12128,N_12271);
or U12525 (N_12525,N_12283,N_12037);
and U12526 (N_12526,N_12295,N_12027);
or U12527 (N_12527,N_12144,N_12127);
xnor U12528 (N_12528,N_12013,N_12240);
nand U12529 (N_12529,N_12133,N_12148);
nor U12530 (N_12530,N_12113,N_12040);
xor U12531 (N_12531,N_12186,N_12020);
or U12532 (N_12532,N_12196,N_12291);
nand U12533 (N_12533,N_12148,N_12151);
and U12534 (N_12534,N_12144,N_12182);
xor U12535 (N_12535,N_12165,N_12121);
nor U12536 (N_12536,N_12105,N_12204);
or U12537 (N_12537,N_12188,N_12224);
nand U12538 (N_12538,N_12260,N_12239);
or U12539 (N_12539,N_12015,N_12280);
or U12540 (N_12540,N_12188,N_12118);
or U12541 (N_12541,N_12292,N_12128);
or U12542 (N_12542,N_12163,N_12024);
nand U12543 (N_12543,N_12097,N_12144);
or U12544 (N_12544,N_12181,N_12136);
xor U12545 (N_12545,N_12210,N_12092);
and U12546 (N_12546,N_12240,N_12174);
nor U12547 (N_12547,N_12048,N_12245);
and U12548 (N_12548,N_12033,N_12137);
and U12549 (N_12549,N_12044,N_12118);
nor U12550 (N_12550,N_12007,N_12000);
nor U12551 (N_12551,N_12265,N_12066);
or U12552 (N_12552,N_12299,N_12108);
xnor U12553 (N_12553,N_12278,N_12029);
nand U12554 (N_12554,N_12236,N_12162);
xnor U12555 (N_12555,N_12268,N_12264);
nor U12556 (N_12556,N_12089,N_12078);
xor U12557 (N_12557,N_12207,N_12139);
nor U12558 (N_12558,N_12253,N_12281);
xnor U12559 (N_12559,N_12009,N_12131);
and U12560 (N_12560,N_12241,N_12212);
xnor U12561 (N_12561,N_12144,N_12244);
xor U12562 (N_12562,N_12201,N_12232);
nor U12563 (N_12563,N_12153,N_12217);
or U12564 (N_12564,N_12216,N_12182);
xor U12565 (N_12565,N_12141,N_12249);
nor U12566 (N_12566,N_12084,N_12256);
nand U12567 (N_12567,N_12064,N_12117);
nor U12568 (N_12568,N_12294,N_12043);
or U12569 (N_12569,N_12059,N_12193);
or U12570 (N_12570,N_12045,N_12120);
nand U12571 (N_12571,N_12131,N_12063);
and U12572 (N_12572,N_12282,N_12159);
xor U12573 (N_12573,N_12149,N_12003);
and U12574 (N_12574,N_12203,N_12117);
nor U12575 (N_12575,N_12236,N_12120);
nor U12576 (N_12576,N_12004,N_12162);
nand U12577 (N_12577,N_12065,N_12081);
xor U12578 (N_12578,N_12065,N_12151);
nand U12579 (N_12579,N_12015,N_12239);
xor U12580 (N_12580,N_12150,N_12244);
nand U12581 (N_12581,N_12211,N_12195);
or U12582 (N_12582,N_12233,N_12084);
nor U12583 (N_12583,N_12207,N_12195);
nand U12584 (N_12584,N_12080,N_12233);
nor U12585 (N_12585,N_12044,N_12234);
nand U12586 (N_12586,N_12263,N_12013);
or U12587 (N_12587,N_12220,N_12170);
or U12588 (N_12588,N_12197,N_12159);
xor U12589 (N_12589,N_12248,N_12122);
nand U12590 (N_12590,N_12105,N_12125);
xor U12591 (N_12591,N_12161,N_12232);
or U12592 (N_12592,N_12295,N_12162);
nand U12593 (N_12593,N_12234,N_12152);
xnor U12594 (N_12594,N_12099,N_12130);
and U12595 (N_12595,N_12005,N_12147);
and U12596 (N_12596,N_12243,N_12227);
and U12597 (N_12597,N_12244,N_12157);
xor U12598 (N_12598,N_12252,N_12215);
nor U12599 (N_12599,N_12195,N_12256);
xor U12600 (N_12600,N_12321,N_12481);
nand U12601 (N_12601,N_12379,N_12490);
nand U12602 (N_12602,N_12366,N_12476);
and U12603 (N_12603,N_12505,N_12463);
and U12604 (N_12604,N_12347,N_12363);
and U12605 (N_12605,N_12351,N_12587);
and U12606 (N_12606,N_12525,N_12445);
xnor U12607 (N_12607,N_12548,N_12342);
nand U12608 (N_12608,N_12338,N_12494);
nand U12609 (N_12609,N_12408,N_12407);
and U12610 (N_12610,N_12499,N_12323);
nand U12611 (N_12611,N_12496,N_12550);
xnor U12612 (N_12612,N_12521,N_12566);
xnor U12613 (N_12613,N_12329,N_12564);
and U12614 (N_12614,N_12325,N_12447);
nor U12615 (N_12615,N_12393,N_12568);
or U12616 (N_12616,N_12519,N_12560);
or U12617 (N_12617,N_12511,N_12343);
or U12618 (N_12618,N_12431,N_12387);
nor U12619 (N_12619,N_12561,N_12554);
nor U12620 (N_12620,N_12535,N_12444);
nand U12621 (N_12621,N_12355,N_12576);
xor U12622 (N_12622,N_12312,N_12544);
nand U12623 (N_12623,N_12435,N_12324);
nand U12624 (N_12624,N_12388,N_12482);
or U12625 (N_12625,N_12436,N_12516);
xor U12626 (N_12626,N_12417,N_12359);
and U12627 (N_12627,N_12501,N_12491);
nor U12628 (N_12628,N_12339,N_12441);
and U12629 (N_12629,N_12307,N_12365);
xor U12630 (N_12630,N_12429,N_12372);
or U12631 (N_12631,N_12493,N_12327);
and U12632 (N_12632,N_12396,N_12461);
xor U12633 (N_12633,N_12403,N_12598);
or U12634 (N_12634,N_12410,N_12562);
and U12635 (N_12635,N_12506,N_12328);
or U12636 (N_12636,N_12440,N_12402);
and U12637 (N_12637,N_12424,N_12585);
nand U12638 (N_12638,N_12427,N_12563);
nand U12639 (N_12639,N_12474,N_12534);
xor U12640 (N_12640,N_12477,N_12446);
or U12641 (N_12641,N_12483,N_12421);
or U12642 (N_12642,N_12306,N_12539);
nand U12643 (N_12643,N_12443,N_12460);
nand U12644 (N_12644,N_12442,N_12599);
and U12645 (N_12645,N_12449,N_12570);
nand U12646 (N_12646,N_12466,N_12318);
xor U12647 (N_12647,N_12378,N_12553);
nand U12648 (N_12648,N_12345,N_12597);
nor U12649 (N_12649,N_12594,N_12334);
or U12650 (N_12650,N_12352,N_12502);
nand U12651 (N_12651,N_12484,N_12551);
nand U12652 (N_12652,N_12565,N_12391);
nand U12653 (N_12653,N_12361,N_12405);
or U12654 (N_12654,N_12572,N_12357);
and U12655 (N_12655,N_12448,N_12302);
xor U12656 (N_12656,N_12386,N_12376);
xnor U12657 (N_12657,N_12344,N_12577);
or U12658 (N_12658,N_12320,N_12542);
or U12659 (N_12659,N_12520,N_12541);
xor U12660 (N_12660,N_12303,N_12454);
and U12661 (N_12661,N_12335,N_12308);
or U12662 (N_12662,N_12371,N_12510);
nand U12663 (N_12663,N_12438,N_12336);
nand U12664 (N_12664,N_12399,N_12558);
xnor U12665 (N_12665,N_12559,N_12332);
nor U12666 (N_12666,N_12341,N_12508);
nand U12667 (N_12667,N_12432,N_12479);
and U12668 (N_12668,N_12513,N_12579);
or U12669 (N_12669,N_12540,N_12588);
xor U12670 (N_12670,N_12547,N_12418);
xnor U12671 (N_12671,N_12348,N_12375);
xnor U12672 (N_12672,N_12313,N_12364);
or U12673 (N_12673,N_12582,N_12314);
xor U12674 (N_12674,N_12575,N_12409);
nand U12675 (N_12675,N_12422,N_12404);
and U12676 (N_12676,N_12526,N_12395);
or U12677 (N_12677,N_12475,N_12381);
nand U12678 (N_12678,N_12549,N_12392);
nor U12679 (N_12679,N_12349,N_12412);
xnor U12680 (N_12680,N_12353,N_12414);
nand U12681 (N_12681,N_12420,N_12380);
and U12682 (N_12682,N_12552,N_12319);
nand U12683 (N_12683,N_12531,N_12437);
xnor U12684 (N_12684,N_12425,N_12589);
xor U12685 (N_12685,N_12331,N_12413);
xor U12686 (N_12686,N_12428,N_12337);
or U12687 (N_12687,N_12310,N_12368);
nand U12688 (N_12688,N_12301,N_12583);
or U12689 (N_12689,N_12528,N_12369);
nor U12690 (N_12690,N_12543,N_12584);
xnor U12691 (N_12691,N_12362,N_12382);
xor U12692 (N_12692,N_12469,N_12517);
or U12693 (N_12693,N_12459,N_12488);
nor U12694 (N_12694,N_12545,N_12567);
nor U12695 (N_12695,N_12497,N_12573);
xor U12696 (N_12696,N_12370,N_12512);
and U12697 (N_12697,N_12557,N_12423);
and U12698 (N_12698,N_12500,N_12596);
xnor U12699 (N_12699,N_12415,N_12555);
or U12700 (N_12700,N_12453,N_12530);
nor U12701 (N_12701,N_12305,N_12406);
or U12702 (N_12702,N_12581,N_12580);
nor U12703 (N_12703,N_12346,N_12401);
or U12704 (N_12704,N_12471,N_12489);
xnor U12705 (N_12705,N_12592,N_12467);
xnor U12706 (N_12706,N_12456,N_12509);
and U12707 (N_12707,N_12383,N_12518);
or U12708 (N_12708,N_12486,N_12394);
or U12709 (N_12709,N_12590,N_12574);
nand U12710 (N_12710,N_12457,N_12333);
nor U12711 (N_12711,N_12411,N_12350);
nor U12712 (N_12712,N_12398,N_12400);
nand U12713 (N_12713,N_12356,N_12311);
nor U12714 (N_12714,N_12485,N_12522);
or U12715 (N_12715,N_12586,N_12593);
nand U12716 (N_12716,N_12495,N_12529);
nor U12717 (N_12717,N_12373,N_12472);
and U12718 (N_12718,N_12492,N_12309);
xor U12719 (N_12719,N_12468,N_12300);
or U12720 (N_12720,N_12464,N_12462);
or U12721 (N_12721,N_12470,N_12384);
xnor U12722 (N_12722,N_12434,N_12533);
nand U12723 (N_12723,N_12397,N_12451);
nand U12724 (N_12724,N_12374,N_12536);
nand U12725 (N_12725,N_12316,N_12367);
or U12726 (N_12726,N_12419,N_12538);
xor U12727 (N_12727,N_12487,N_12317);
or U12728 (N_12728,N_12439,N_12455);
xor U12729 (N_12729,N_12473,N_12571);
xnor U12730 (N_12730,N_12304,N_12452);
nand U12731 (N_12731,N_12527,N_12578);
nand U12732 (N_12732,N_12450,N_12426);
xor U12733 (N_12733,N_12515,N_12480);
or U12734 (N_12734,N_12478,N_12377);
xor U12735 (N_12735,N_12358,N_12322);
nor U12736 (N_12736,N_12430,N_12532);
xnor U12737 (N_12737,N_12514,N_12556);
nand U12738 (N_12738,N_12433,N_12595);
nor U12739 (N_12739,N_12546,N_12340);
and U12740 (N_12740,N_12591,N_12416);
and U12741 (N_12741,N_12507,N_12504);
or U12742 (N_12742,N_12498,N_12385);
nand U12743 (N_12743,N_12390,N_12330);
or U12744 (N_12744,N_12523,N_12354);
nand U12745 (N_12745,N_12360,N_12458);
nor U12746 (N_12746,N_12389,N_12524);
xor U12747 (N_12747,N_12569,N_12315);
xnor U12748 (N_12748,N_12503,N_12326);
xor U12749 (N_12749,N_12537,N_12465);
or U12750 (N_12750,N_12425,N_12324);
nor U12751 (N_12751,N_12487,N_12464);
nor U12752 (N_12752,N_12482,N_12427);
xor U12753 (N_12753,N_12335,N_12527);
and U12754 (N_12754,N_12583,N_12427);
or U12755 (N_12755,N_12347,N_12460);
nor U12756 (N_12756,N_12453,N_12589);
nor U12757 (N_12757,N_12477,N_12471);
or U12758 (N_12758,N_12517,N_12432);
nor U12759 (N_12759,N_12501,N_12379);
nand U12760 (N_12760,N_12342,N_12359);
or U12761 (N_12761,N_12387,N_12426);
and U12762 (N_12762,N_12551,N_12457);
nor U12763 (N_12763,N_12522,N_12330);
or U12764 (N_12764,N_12452,N_12432);
and U12765 (N_12765,N_12460,N_12358);
and U12766 (N_12766,N_12401,N_12386);
nand U12767 (N_12767,N_12392,N_12525);
xor U12768 (N_12768,N_12335,N_12586);
nand U12769 (N_12769,N_12556,N_12500);
nand U12770 (N_12770,N_12490,N_12423);
xor U12771 (N_12771,N_12444,N_12303);
and U12772 (N_12772,N_12398,N_12482);
and U12773 (N_12773,N_12333,N_12409);
and U12774 (N_12774,N_12484,N_12335);
nor U12775 (N_12775,N_12378,N_12574);
xor U12776 (N_12776,N_12451,N_12541);
nor U12777 (N_12777,N_12361,N_12334);
and U12778 (N_12778,N_12308,N_12499);
and U12779 (N_12779,N_12507,N_12343);
nor U12780 (N_12780,N_12434,N_12323);
nand U12781 (N_12781,N_12513,N_12463);
and U12782 (N_12782,N_12404,N_12556);
or U12783 (N_12783,N_12437,N_12597);
or U12784 (N_12784,N_12477,N_12430);
xnor U12785 (N_12785,N_12373,N_12505);
nor U12786 (N_12786,N_12393,N_12523);
or U12787 (N_12787,N_12321,N_12398);
nor U12788 (N_12788,N_12378,N_12479);
and U12789 (N_12789,N_12346,N_12533);
xnor U12790 (N_12790,N_12392,N_12436);
nor U12791 (N_12791,N_12342,N_12331);
nand U12792 (N_12792,N_12427,N_12348);
nand U12793 (N_12793,N_12337,N_12520);
xor U12794 (N_12794,N_12467,N_12532);
and U12795 (N_12795,N_12345,N_12340);
nand U12796 (N_12796,N_12409,N_12368);
nand U12797 (N_12797,N_12543,N_12368);
and U12798 (N_12798,N_12338,N_12570);
nor U12799 (N_12799,N_12331,N_12457);
and U12800 (N_12800,N_12371,N_12542);
and U12801 (N_12801,N_12587,N_12480);
or U12802 (N_12802,N_12450,N_12447);
nand U12803 (N_12803,N_12321,N_12571);
xnor U12804 (N_12804,N_12464,N_12575);
xor U12805 (N_12805,N_12316,N_12382);
nand U12806 (N_12806,N_12332,N_12539);
and U12807 (N_12807,N_12470,N_12369);
and U12808 (N_12808,N_12367,N_12402);
and U12809 (N_12809,N_12491,N_12322);
nand U12810 (N_12810,N_12531,N_12358);
xnor U12811 (N_12811,N_12400,N_12537);
and U12812 (N_12812,N_12478,N_12447);
or U12813 (N_12813,N_12378,N_12504);
nor U12814 (N_12814,N_12358,N_12503);
xnor U12815 (N_12815,N_12502,N_12464);
xnor U12816 (N_12816,N_12315,N_12333);
nand U12817 (N_12817,N_12470,N_12393);
or U12818 (N_12818,N_12526,N_12371);
nor U12819 (N_12819,N_12493,N_12594);
nand U12820 (N_12820,N_12584,N_12578);
nand U12821 (N_12821,N_12462,N_12380);
or U12822 (N_12822,N_12393,N_12576);
and U12823 (N_12823,N_12429,N_12421);
nand U12824 (N_12824,N_12330,N_12447);
nand U12825 (N_12825,N_12518,N_12362);
nor U12826 (N_12826,N_12566,N_12540);
xnor U12827 (N_12827,N_12400,N_12567);
nor U12828 (N_12828,N_12587,N_12414);
nand U12829 (N_12829,N_12356,N_12532);
nand U12830 (N_12830,N_12585,N_12448);
nand U12831 (N_12831,N_12368,N_12430);
xor U12832 (N_12832,N_12479,N_12514);
xnor U12833 (N_12833,N_12564,N_12331);
nor U12834 (N_12834,N_12341,N_12407);
nor U12835 (N_12835,N_12413,N_12591);
nor U12836 (N_12836,N_12396,N_12367);
xor U12837 (N_12837,N_12338,N_12372);
nand U12838 (N_12838,N_12357,N_12348);
nor U12839 (N_12839,N_12433,N_12392);
and U12840 (N_12840,N_12505,N_12454);
nor U12841 (N_12841,N_12376,N_12404);
and U12842 (N_12842,N_12559,N_12386);
nor U12843 (N_12843,N_12436,N_12384);
nand U12844 (N_12844,N_12513,N_12385);
xnor U12845 (N_12845,N_12303,N_12568);
and U12846 (N_12846,N_12531,N_12466);
xor U12847 (N_12847,N_12454,N_12506);
nand U12848 (N_12848,N_12436,N_12354);
nor U12849 (N_12849,N_12318,N_12306);
nor U12850 (N_12850,N_12563,N_12417);
nor U12851 (N_12851,N_12359,N_12419);
xor U12852 (N_12852,N_12474,N_12513);
xor U12853 (N_12853,N_12361,N_12459);
xor U12854 (N_12854,N_12452,N_12333);
or U12855 (N_12855,N_12415,N_12512);
nor U12856 (N_12856,N_12428,N_12598);
xor U12857 (N_12857,N_12422,N_12504);
nand U12858 (N_12858,N_12560,N_12599);
nor U12859 (N_12859,N_12505,N_12432);
nand U12860 (N_12860,N_12402,N_12472);
nand U12861 (N_12861,N_12525,N_12407);
xor U12862 (N_12862,N_12519,N_12370);
nor U12863 (N_12863,N_12500,N_12480);
nor U12864 (N_12864,N_12555,N_12351);
nor U12865 (N_12865,N_12493,N_12380);
and U12866 (N_12866,N_12558,N_12383);
nand U12867 (N_12867,N_12575,N_12544);
or U12868 (N_12868,N_12333,N_12306);
xor U12869 (N_12869,N_12402,N_12493);
and U12870 (N_12870,N_12341,N_12406);
or U12871 (N_12871,N_12509,N_12392);
nand U12872 (N_12872,N_12311,N_12541);
nor U12873 (N_12873,N_12356,N_12592);
and U12874 (N_12874,N_12371,N_12469);
and U12875 (N_12875,N_12417,N_12578);
or U12876 (N_12876,N_12427,N_12526);
xor U12877 (N_12877,N_12547,N_12303);
nand U12878 (N_12878,N_12395,N_12328);
nand U12879 (N_12879,N_12408,N_12360);
xor U12880 (N_12880,N_12539,N_12372);
nand U12881 (N_12881,N_12587,N_12599);
nor U12882 (N_12882,N_12597,N_12402);
or U12883 (N_12883,N_12534,N_12539);
nor U12884 (N_12884,N_12456,N_12332);
nand U12885 (N_12885,N_12416,N_12565);
nor U12886 (N_12886,N_12375,N_12467);
or U12887 (N_12887,N_12371,N_12406);
or U12888 (N_12888,N_12311,N_12464);
nand U12889 (N_12889,N_12574,N_12327);
nand U12890 (N_12890,N_12317,N_12370);
and U12891 (N_12891,N_12401,N_12530);
nand U12892 (N_12892,N_12377,N_12474);
nand U12893 (N_12893,N_12491,N_12399);
nand U12894 (N_12894,N_12515,N_12390);
xor U12895 (N_12895,N_12468,N_12464);
or U12896 (N_12896,N_12313,N_12311);
nand U12897 (N_12897,N_12417,N_12499);
nand U12898 (N_12898,N_12518,N_12331);
nand U12899 (N_12899,N_12574,N_12330);
nor U12900 (N_12900,N_12770,N_12887);
nor U12901 (N_12901,N_12752,N_12796);
and U12902 (N_12902,N_12619,N_12762);
or U12903 (N_12903,N_12607,N_12795);
nand U12904 (N_12904,N_12755,N_12773);
xnor U12905 (N_12905,N_12705,N_12726);
and U12906 (N_12906,N_12818,N_12868);
nor U12907 (N_12907,N_12636,N_12841);
nand U12908 (N_12908,N_12661,N_12806);
nor U12909 (N_12909,N_12675,N_12882);
or U12910 (N_12910,N_12878,N_12898);
nand U12911 (N_12911,N_12814,N_12648);
or U12912 (N_12912,N_12679,N_12828);
or U12913 (N_12913,N_12876,N_12712);
or U12914 (N_12914,N_12644,N_12824);
or U12915 (N_12915,N_12608,N_12685);
and U12916 (N_12916,N_12823,N_12757);
nand U12917 (N_12917,N_12670,N_12656);
or U12918 (N_12918,N_12885,N_12689);
xor U12919 (N_12919,N_12849,N_12838);
nor U12920 (N_12920,N_12682,N_12810);
nand U12921 (N_12921,N_12746,N_12719);
xnor U12922 (N_12922,N_12664,N_12684);
or U12923 (N_12923,N_12758,N_12729);
nor U12924 (N_12924,N_12804,N_12601);
and U12925 (N_12925,N_12869,N_12693);
and U12926 (N_12926,N_12843,N_12788);
xor U12927 (N_12927,N_12884,N_12723);
and U12928 (N_12928,N_12650,N_12744);
nand U12929 (N_12929,N_12750,N_12791);
xnor U12930 (N_12930,N_12753,N_12618);
nand U12931 (N_12931,N_12674,N_12658);
xor U12932 (N_12932,N_12751,N_12771);
xnor U12933 (N_12933,N_12604,N_12812);
nor U12934 (N_12934,N_12735,N_12805);
xnor U12935 (N_12935,N_12766,N_12802);
and U12936 (N_12936,N_12842,N_12688);
nand U12937 (N_12937,N_12799,N_12890);
and U12938 (N_12938,N_12700,N_12754);
and U12939 (N_12939,N_12867,N_12653);
nand U12940 (N_12940,N_12871,N_12769);
or U12941 (N_12941,N_12739,N_12774);
or U12942 (N_12942,N_12632,N_12895);
and U12943 (N_12943,N_12809,N_12780);
xor U12944 (N_12944,N_12612,N_12819);
and U12945 (N_12945,N_12800,N_12870);
or U12946 (N_12946,N_12775,N_12781);
nand U12947 (N_12947,N_12764,N_12654);
nand U12948 (N_12948,N_12856,N_12732);
xnor U12949 (N_12949,N_12865,N_12695);
and U12950 (N_12950,N_12629,N_12665);
and U12951 (N_12951,N_12738,N_12696);
nand U12952 (N_12952,N_12850,N_12760);
xnor U12953 (N_12953,N_12657,N_12829);
xor U12954 (N_12954,N_12763,N_12733);
nand U12955 (N_12955,N_12896,N_12745);
xnor U12956 (N_12956,N_12721,N_12645);
and U12957 (N_12957,N_12702,N_12718);
nor U12958 (N_12958,N_12892,N_12639);
and U12959 (N_12959,N_12697,N_12894);
nor U12960 (N_12960,N_12724,N_12741);
nand U12961 (N_12961,N_12672,N_12704);
or U12962 (N_12962,N_12787,N_12826);
and U12963 (N_12963,N_12680,N_12606);
and U12964 (N_12964,N_12866,N_12716);
nand U12965 (N_12965,N_12853,N_12840);
or U12966 (N_12966,N_12649,N_12813);
and U12967 (N_12967,N_12715,N_12625);
or U12968 (N_12968,N_12683,N_12839);
and U12969 (N_12969,N_12893,N_12634);
nand U12970 (N_12970,N_12877,N_12628);
and U12971 (N_12971,N_12662,N_12659);
nor U12972 (N_12972,N_12633,N_12666);
and U12973 (N_12973,N_12671,N_12709);
and U12974 (N_12974,N_12873,N_12891);
or U12975 (N_12975,N_12631,N_12861);
and U12976 (N_12976,N_12779,N_12616);
nor U12977 (N_12977,N_12827,N_12785);
and U12978 (N_12978,N_12831,N_12707);
nand U12979 (N_12979,N_12797,N_12711);
xnor U12980 (N_12980,N_12730,N_12848);
nand U12981 (N_12981,N_12815,N_12889);
or U12982 (N_12982,N_12832,N_12691);
nor U12983 (N_12983,N_12742,N_12676);
nand U12984 (N_12984,N_12782,N_12825);
nor U12985 (N_12985,N_12647,N_12860);
and U12986 (N_12986,N_12611,N_12602);
nor U12987 (N_12987,N_12765,N_12710);
and U12988 (N_12988,N_12678,N_12655);
nand U12989 (N_12989,N_12880,N_12743);
and U12990 (N_12990,N_12673,N_12652);
nand U12991 (N_12991,N_12600,N_12845);
nor U12992 (N_12992,N_12722,N_12899);
xnor U12993 (N_12993,N_12792,N_12635);
nor U12994 (N_12994,N_12663,N_12759);
or U12995 (N_12995,N_12640,N_12690);
nand U12996 (N_12996,N_12784,N_12835);
nand U12997 (N_12997,N_12768,N_12807);
and U12998 (N_12998,N_12669,N_12725);
nand U12999 (N_12999,N_12816,N_12811);
and U13000 (N_13000,N_12677,N_12660);
xor U13001 (N_13001,N_12615,N_12778);
or U13002 (N_13002,N_12864,N_12605);
or U13003 (N_13003,N_12803,N_12681);
nand U13004 (N_13004,N_12874,N_12687);
nand U13005 (N_13005,N_12881,N_12855);
nor U13006 (N_13006,N_12621,N_12630);
nor U13007 (N_13007,N_12830,N_12613);
xor U13008 (N_13008,N_12699,N_12767);
nor U13009 (N_13009,N_12668,N_12610);
xnor U13010 (N_13010,N_12609,N_12728);
or U13011 (N_13011,N_12620,N_12638);
and U13012 (N_13012,N_12777,N_12617);
xnor U13013 (N_13013,N_12761,N_12720);
and U13014 (N_13014,N_12651,N_12789);
xnor U13015 (N_13015,N_12667,N_12614);
and U13016 (N_13016,N_12886,N_12794);
xor U13017 (N_13017,N_12749,N_12772);
or U13018 (N_13018,N_12747,N_12851);
nand U13019 (N_13019,N_12736,N_12686);
nand U13020 (N_13020,N_12833,N_12740);
nand U13021 (N_13021,N_12737,N_12820);
nor U13022 (N_13022,N_12646,N_12879);
nand U13023 (N_13023,N_12862,N_12626);
and U13024 (N_13024,N_12852,N_12847);
and U13025 (N_13025,N_12821,N_12748);
and U13026 (N_13026,N_12854,N_12883);
and U13027 (N_13027,N_12808,N_12857);
nand U13028 (N_13028,N_12844,N_12703);
xnor U13029 (N_13029,N_12713,N_12706);
or U13030 (N_13030,N_12623,N_12786);
or U13031 (N_13031,N_12714,N_12834);
nand U13032 (N_13032,N_12817,N_12642);
or U13033 (N_13033,N_12837,N_12888);
or U13034 (N_13034,N_12783,N_12822);
xnor U13035 (N_13035,N_12624,N_12727);
nand U13036 (N_13036,N_12643,N_12798);
and U13037 (N_13037,N_12603,N_12734);
nand U13038 (N_13038,N_12872,N_12793);
xnor U13039 (N_13039,N_12846,N_12641);
or U13040 (N_13040,N_12897,N_12717);
nor U13041 (N_13041,N_12858,N_12875);
and U13042 (N_13042,N_12698,N_12731);
and U13043 (N_13043,N_12622,N_12637);
nand U13044 (N_13044,N_12708,N_12756);
nor U13045 (N_13045,N_12627,N_12694);
nor U13046 (N_13046,N_12863,N_12859);
and U13047 (N_13047,N_12801,N_12836);
nor U13048 (N_13048,N_12701,N_12790);
and U13049 (N_13049,N_12692,N_12776);
xnor U13050 (N_13050,N_12787,N_12896);
nand U13051 (N_13051,N_12737,N_12824);
or U13052 (N_13052,N_12864,N_12636);
and U13053 (N_13053,N_12756,N_12813);
nand U13054 (N_13054,N_12725,N_12768);
nand U13055 (N_13055,N_12868,N_12643);
xnor U13056 (N_13056,N_12621,N_12710);
or U13057 (N_13057,N_12673,N_12882);
or U13058 (N_13058,N_12662,N_12832);
and U13059 (N_13059,N_12765,N_12726);
or U13060 (N_13060,N_12601,N_12666);
or U13061 (N_13061,N_12616,N_12770);
xnor U13062 (N_13062,N_12782,N_12731);
or U13063 (N_13063,N_12615,N_12678);
and U13064 (N_13064,N_12809,N_12737);
nor U13065 (N_13065,N_12719,N_12676);
nor U13066 (N_13066,N_12807,N_12779);
and U13067 (N_13067,N_12611,N_12846);
and U13068 (N_13068,N_12854,N_12657);
or U13069 (N_13069,N_12872,N_12707);
nor U13070 (N_13070,N_12714,N_12823);
or U13071 (N_13071,N_12872,N_12692);
nand U13072 (N_13072,N_12849,N_12804);
nand U13073 (N_13073,N_12685,N_12640);
or U13074 (N_13074,N_12800,N_12832);
nand U13075 (N_13075,N_12718,N_12712);
nand U13076 (N_13076,N_12746,N_12607);
and U13077 (N_13077,N_12618,N_12896);
xor U13078 (N_13078,N_12616,N_12867);
xnor U13079 (N_13079,N_12662,N_12788);
nand U13080 (N_13080,N_12764,N_12628);
xor U13081 (N_13081,N_12781,N_12696);
or U13082 (N_13082,N_12898,N_12707);
xnor U13083 (N_13083,N_12761,N_12829);
and U13084 (N_13084,N_12807,N_12811);
xnor U13085 (N_13085,N_12653,N_12715);
or U13086 (N_13086,N_12696,N_12739);
nor U13087 (N_13087,N_12638,N_12774);
xnor U13088 (N_13088,N_12705,N_12885);
and U13089 (N_13089,N_12883,N_12715);
xnor U13090 (N_13090,N_12779,N_12731);
and U13091 (N_13091,N_12655,N_12828);
xnor U13092 (N_13092,N_12807,N_12788);
nand U13093 (N_13093,N_12780,N_12833);
nor U13094 (N_13094,N_12789,N_12876);
xor U13095 (N_13095,N_12727,N_12781);
and U13096 (N_13096,N_12725,N_12637);
nor U13097 (N_13097,N_12766,N_12869);
xnor U13098 (N_13098,N_12603,N_12844);
and U13099 (N_13099,N_12637,N_12712);
xor U13100 (N_13100,N_12722,N_12647);
xor U13101 (N_13101,N_12725,N_12742);
xor U13102 (N_13102,N_12808,N_12660);
nor U13103 (N_13103,N_12671,N_12744);
nand U13104 (N_13104,N_12672,N_12614);
nand U13105 (N_13105,N_12840,N_12835);
and U13106 (N_13106,N_12743,N_12633);
nor U13107 (N_13107,N_12707,N_12722);
xor U13108 (N_13108,N_12815,N_12887);
or U13109 (N_13109,N_12729,N_12886);
nand U13110 (N_13110,N_12800,N_12621);
or U13111 (N_13111,N_12802,N_12630);
nor U13112 (N_13112,N_12742,N_12855);
nor U13113 (N_13113,N_12679,N_12687);
or U13114 (N_13114,N_12848,N_12753);
or U13115 (N_13115,N_12602,N_12603);
nor U13116 (N_13116,N_12770,N_12620);
or U13117 (N_13117,N_12851,N_12679);
nor U13118 (N_13118,N_12714,N_12829);
or U13119 (N_13119,N_12734,N_12728);
nand U13120 (N_13120,N_12678,N_12872);
and U13121 (N_13121,N_12779,N_12667);
nor U13122 (N_13122,N_12865,N_12748);
or U13123 (N_13123,N_12679,N_12886);
or U13124 (N_13124,N_12832,N_12636);
and U13125 (N_13125,N_12654,N_12892);
or U13126 (N_13126,N_12871,N_12712);
nand U13127 (N_13127,N_12839,N_12613);
xnor U13128 (N_13128,N_12752,N_12823);
nor U13129 (N_13129,N_12610,N_12626);
xor U13130 (N_13130,N_12838,N_12696);
and U13131 (N_13131,N_12731,N_12711);
or U13132 (N_13132,N_12743,N_12832);
xnor U13133 (N_13133,N_12821,N_12740);
nand U13134 (N_13134,N_12844,N_12853);
nor U13135 (N_13135,N_12897,N_12755);
or U13136 (N_13136,N_12600,N_12616);
nand U13137 (N_13137,N_12634,N_12616);
or U13138 (N_13138,N_12843,N_12889);
nor U13139 (N_13139,N_12778,N_12672);
nand U13140 (N_13140,N_12794,N_12755);
or U13141 (N_13141,N_12845,N_12834);
or U13142 (N_13142,N_12672,N_12737);
and U13143 (N_13143,N_12823,N_12600);
xor U13144 (N_13144,N_12636,N_12701);
nor U13145 (N_13145,N_12813,N_12747);
and U13146 (N_13146,N_12859,N_12646);
or U13147 (N_13147,N_12748,N_12832);
nor U13148 (N_13148,N_12698,N_12789);
and U13149 (N_13149,N_12882,N_12801);
nand U13150 (N_13150,N_12756,N_12705);
nor U13151 (N_13151,N_12895,N_12733);
nor U13152 (N_13152,N_12719,N_12639);
or U13153 (N_13153,N_12869,N_12728);
or U13154 (N_13154,N_12740,N_12700);
xnor U13155 (N_13155,N_12690,N_12777);
and U13156 (N_13156,N_12735,N_12642);
and U13157 (N_13157,N_12712,N_12794);
nand U13158 (N_13158,N_12841,N_12721);
xnor U13159 (N_13159,N_12858,N_12743);
or U13160 (N_13160,N_12620,N_12703);
nand U13161 (N_13161,N_12635,N_12888);
xor U13162 (N_13162,N_12803,N_12880);
or U13163 (N_13163,N_12639,N_12854);
nand U13164 (N_13164,N_12693,N_12626);
or U13165 (N_13165,N_12690,N_12785);
nand U13166 (N_13166,N_12662,N_12704);
nor U13167 (N_13167,N_12639,N_12805);
and U13168 (N_13168,N_12871,N_12625);
nand U13169 (N_13169,N_12838,N_12841);
or U13170 (N_13170,N_12736,N_12669);
nor U13171 (N_13171,N_12703,N_12624);
nor U13172 (N_13172,N_12834,N_12610);
xor U13173 (N_13173,N_12605,N_12841);
and U13174 (N_13174,N_12604,N_12870);
and U13175 (N_13175,N_12886,N_12691);
xor U13176 (N_13176,N_12611,N_12783);
and U13177 (N_13177,N_12732,N_12705);
nand U13178 (N_13178,N_12646,N_12873);
or U13179 (N_13179,N_12823,N_12825);
or U13180 (N_13180,N_12852,N_12830);
and U13181 (N_13181,N_12771,N_12767);
or U13182 (N_13182,N_12738,N_12602);
and U13183 (N_13183,N_12676,N_12770);
xnor U13184 (N_13184,N_12823,N_12607);
and U13185 (N_13185,N_12655,N_12681);
nand U13186 (N_13186,N_12670,N_12794);
nor U13187 (N_13187,N_12780,N_12633);
xor U13188 (N_13188,N_12720,N_12786);
nor U13189 (N_13189,N_12803,N_12873);
nor U13190 (N_13190,N_12675,N_12826);
xor U13191 (N_13191,N_12640,N_12670);
nand U13192 (N_13192,N_12840,N_12818);
xnor U13193 (N_13193,N_12648,N_12766);
nand U13194 (N_13194,N_12787,N_12858);
nand U13195 (N_13195,N_12860,N_12697);
nand U13196 (N_13196,N_12702,N_12843);
nor U13197 (N_13197,N_12615,N_12899);
nor U13198 (N_13198,N_12711,N_12709);
xor U13199 (N_13199,N_12899,N_12842);
or U13200 (N_13200,N_13139,N_13175);
xnor U13201 (N_13201,N_12960,N_13089);
nand U13202 (N_13202,N_13077,N_12996);
or U13203 (N_13203,N_13073,N_13143);
or U13204 (N_13204,N_13045,N_13162);
or U13205 (N_13205,N_12910,N_13066);
nand U13206 (N_13206,N_12972,N_13093);
or U13207 (N_13207,N_13053,N_13178);
or U13208 (N_13208,N_13019,N_13122);
nor U13209 (N_13209,N_13003,N_13188);
nand U13210 (N_13210,N_13186,N_13080);
xnor U13211 (N_13211,N_12952,N_13129);
nand U13212 (N_13212,N_12942,N_13123);
xor U13213 (N_13213,N_13159,N_12905);
and U13214 (N_13214,N_12947,N_13191);
nand U13215 (N_13215,N_12975,N_13114);
nor U13216 (N_13216,N_13033,N_13108);
or U13217 (N_13217,N_13124,N_13150);
and U13218 (N_13218,N_13136,N_13034);
nand U13219 (N_13219,N_13095,N_13144);
nand U13220 (N_13220,N_13088,N_12948);
nand U13221 (N_13221,N_13086,N_12982);
and U13222 (N_13222,N_13098,N_12980);
xnor U13223 (N_13223,N_12904,N_13107);
nor U13224 (N_13224,N_12930,N_13177);
or U13225 (N_13225,N_13041,N_13063);
and U13226 (N_13226,N_12915,N_13010);
and U13227 (N_13227,N_13052,N_13085);
or U13228 (N_13228,N_13040,N_12959);
nand U13229 (N_13229,N_13047,N_13110);
nand U13230 (N_13230,N_13198,N_13035);
xor U13231 (N_13231,N_13069,N_12953);
nand U13232 (N_13232,N_13032,N_12964);
xnor U13233 (N_13233,N_13071,N_12977);
and U13234 (N_13234,N_12974,N_12936);
nor U13235 (N_13235,N_13149,N_13082);
xor U13236 (N_13236,N_12920,N_13091);
nand U13237 (N_13237,N_12968,N_13015);
and U13238 (N_13238,N_12950,N_12916);
nand U13239 (N_13239,N_13100,N_13044);
and U13240 (N_13240,N_13163,N_12967);
or U13241 (N_13241,N_13170,N_13043);
and U13242 (N_13242,N_13151,N_12945);
or U13243 (N_13243,N_13038,N_13103);
or U13244 (N_13244,N_13167,N_13017);
nor U13245 (N_13245,N_13018,N_13160);
nor U13246 (N_13246,N_12971,N_13014);
nand U13247 (N_13247,N_13116,N_12956);
and U13248 (N_13248,N_13172,N_13070);
nand U13249 (N_13249,N_13078,N_12925);
nand U13250 (N_13250,N_12913,N_13193);
xnor U13251 (N_13251,N_12909,N_12966);
or U13252 (N_13252,N_13007,N_13011);
and U13253 (N_13253,N_13026,N_13120);
nor U13254 (N_13254,N_13106,N_12938);
nand U13255 (N_13255,N_12903,N_13101);
nor U13256 (N_13256,N_12932,N_12976);
nand U13257 (N_13257,N_12935,N_13165);
nand U13258 (N_13258,N_12984,N_13059);
nand U13259 (N_13259,N_12970,N_13031);
nand U13260 (N_13260,N_13128,N_13174);
nand U13261 (N_13261,N_13176,N_12918);
nand U13262 (N_13262,N_12919,N_13183);
or U13263 (N_13263,N_13060,N_12988);
nor U13264 (N_13264,N_13061,N_12902);
or U13265 (N_13265,N_13154,N_12986);
or U13266 (N_13266,N_13083,N_13084);
or U13267 (N_13267,N_13147,N_12954);
and U13268 (N_13268,N_12963,N_13072);
nor U13269 (N_13269,N_12969,N_13016);
or U13270 (N_13270,N_13008,N_13117);
nor U13271 (N_13271,N_13037,N_13006);
or U13272 (N_13272,N_13009,N_13002);
nor U13273 (N_13273,N_12989,N_13197);
xnor U13274 (N_13274,N_13046,N_12939);
nor U13275 (N_13275,N_12979,N_13153);
and U13276 (N_13276,N_13079,N_12957);
nor U13277 (N_13277,N_12985,N_13161);
xor U13278 (N_13278,N_13028,N_13109);
or U13279 (N_13279,N_12900,N_13022);
or U13280 (N_13280,N_13187,N_12994);
xnor U13281 (N_13281,N_13104,N_13118);
nand U13282 (N_13282,N_12907,N_13181);
nand U13283 (N_13283,N_13048,N_13168);
nand U13284 (N_13284,N_13051,N_12981);
nand U13285 (N_13285,N_12962,N_13194);
xnor U13286 (N_13286,N_12992,N_13189);
or U13287 (N_13287,N_12928,N_13020);
xor U13288 (N_13288,N_12973,N_13097);
and U13289 (N_13289,N_12990,N_13087);
xor U13290 (N_13290,N_13199,N_13021);
and U13291 (N_13291,N_12991,N_13173);
or U13292 (N_13292,N_12965,N_12934);
nor U13293 (N_13293,N_13125,N_13001);
xor U13294 (N_13294,N_12951,N_13130);
xnor U13295 (N_13295,N_12901,N_13075);
nor U13296 (N_13296,N_13024,N_13164);
and U13297 (N_13297,N_13025,N_13190);
nand U13298 (N_13298,N_13005,N_12944);
or U13299 (N_13299,N_13099,N_13064);
xnor U13300 (N_13300,N_12923,N_13179);
nor U13301 (N_13301,N_13180,N_13081);
nand U13302 (N_13302,N_13145,N_12912);
or U13303 (N_13303,N_12987,N_12908);
nand U13304 (N_13304,N_13134,N_12941);
nand U13305 (N_13305,N_12998,N_12937);
nand U13306 (N_13306,N_13036,N_12921);
nor U13307 (N_13307,N_13094,N_13113);
or U13308 (N_13308,N_13142,N_13039);
or U13309 (N_13309,N_12927,N_13049);
and U13310 (N_13310,N_13127,N_13105);
nand U13311 (N_13311,N_13133,N_13192);
xnor U13312 (N_13312,N_13030,N_13119);
xnor U13313 (N_13313,N_12993,N_13121);
nor U13314 (N_13314,N_13090,N_13102);
nand U13315 (N_13315,N_12958,N_13027);
and U13316 (N_13316,N_12924,N_13138);
or U13317 (N_13317,N_13195,N_13042);
or U13318 (N_13318,N_13065,N_13004);
xor U13319 (N_13319,N_12999,N_13132);
xor U13320 (N_13320,N_13112,N_13000);
or U13321 (N_13321,N_13171,N_12949);
nor U13322 (N_13322,N_13169,N_13050);
or U13323 (N_13323,N_13141,N_13062);
nand U13324 (N_13324,N_13068,N_12955);
nor U13325 (N_13325,N_13166,N_13184);
and U13326 (N_13326,N_13013,N_12943);
xor U13327 (N_13327,N_13137,N_12911);
xor U13328 (N_13328,N_13135,N_13157);
or U13329 (N_13329,N_13058,N_13182);
or U13330 (N_13330,N_12940,N_13152);
nand U13331 (N_13331,N_13111,N_13156);
nor U13332 (N_13332,N_12929,N_13131);
and U13333 (N_13333,N_12933,N_13140);
and U13334 (N_13334,N_12931,N_13055);
or U13335 (N_13335,N_13092,N_12983);
nor U13336 (N_13336,N_13185,N_12906);
and U13337 (N_13337,N_13023,N_13056);
or U13338 (N_13338,N_12946,N_12922);
and U13339 (N_13339,N_12914,N_12995);
and U13340 (N_13340,N_13096,N_13146);
xor U13341 (N_13341,N_13126,N_13115);
nor U13342 (N_13342,N_12961,N_12926);
nand U13343 (N_13343,N_13158,N_13057);
or U13344 (N_13344,N_13054,N_13148);
nor U13345 (N_13345,N_13012,N_13196);
xnor U13346 (N_13346,N_12997,N_13074);
nor U13347 (N_13347,N_12978,N_13067);
xnor U13348 (N_13348,N_13029,N_13076);
or U13349 (N_13349,N_12917,N_13155);
nand U13350 (N_13350,N_13160,N_13177);
nand U13351 (N_13351,N_13118,N_13029);
or U13352 (N_13352,N_13167,N_13101);
nor U13353 (N_13353,N_13054,N_13144);
or U13354 (N_13354,N_12920,N_12977);
and U13355 (N_13355,N_13182,N_12951);
xnor U13356 (N_13356,N_13198,N_13078);
or U13357 (N_13357,N_13037,N_12915);
or U13358 (N_13358,N_12980,N_12903);
xor U13359 (N_13359,N_12937,N_13163);
nor U13360 (N_13360,N_13074,N_12959);
nor U13361 (N_13361,N_13153,N_12915);
xnor U13362 (N_13362,N_12933,N_13086);
xor U13363 (N_13363,N_12980,N_13151);
xnor U13364 (N_13364,N_13121,N_13102);
or U13365 (N_13365,N_13174,N_13015);
xnor U13366 (N_13366,N_12917,N_13137);
nand U13367 (N_13367,N_13038,N_13175);
or U13368 (N_13368,N_13058,N_13030);
xnor U13369 (N_13369,N_12942,N_13165);
xnor U13370 (N_13370,N_13163,N_13034);
nor U13371 (N_13371,N_13129,N_12993);
xnor U13372 (N_13372,N_12910,N_13153);
and U13373 (N_13373,N_12999,N_12921);
xor U13374 (N_13374,N_13152,N_13113);
xor U13375 (N_13375,N_13059,N_13196);
and U13376 (N_13376,N_13108,N_12966);
xnor U13377 (N_13377,N_12922,N_13157);
xor U13378 (N_13378,N_13001,N_12912);
and U13379 (N_13379,N_13027,N_12993);
and U13380 (N_13380,N_13163,N_13138);
nor U13381 (N_13381,N_13162,N_13153);
or U13382 (N_13382,N_12943,N_13128);
or U13383 (N_13383,N_13010,N_13132);
nor U13384 (N_13384,N_13165,N_13196);
nor U13385 (N_13385,N_13079,N_13180);
xor U13386 (N_13386,N_13186,N_12994);
nor U13387 (N_13387,N_13141,N_13182);
xnor U13388 (N_13388,N_13178,N_13192);
nand U13389 (N_13389,N_13087,N_12903);
xor U13390 (N_13390,N_12908,N_13097);
xor U13391 (N_13391,N_12906,N_13143);
xor U13392 (N_13392,N_13136,N_13019);
or U13393 (N_13393,N_12962,N_13008);
or U13394 (N_13394,N_13180,N_13023);
nand U13395 (N_13395,N_13112,N_13073);
nor U13396 (N_13396,N_13150,N_12922);
and U13397 (N_13397,N_13026,N_13138);
or U13398 (N_13398,N_13170,N_12904);
xor U13399 (N_13399,N_12900,N_13080);
or U13400 (N_13400,N_12971,N_13155);
nor U13401 (N_13401,N_13119,N_13186);
nand U13402 (N_13402,N_12970,N_13055);
nand U13403 (N_13403,N_12957,N_13170);
xor U13404 (N_13404,N_12927,N_12907);
or U13405 (N_13405,N_12915,N_13072);
nor U13406 (N_13406,N_13168,N_13133);
xor U13407 (N_13407,N_13002,N_13010);
xor U13408 (N_13408,N_13068,N_13019);
xnor U13409 (N_13409,N_12947,N_13186);
xor U13410 (N_13410,N_13050,N_12987);
or U13411 (N_13411,N_12971,N_13044);
nand U13412 (N_13412,N_13072,N_13025);
or U13413 (N_13413,N_13151,N_13055);
nor U13414 (N_13414,N_12918,N_13049);
nand U13415 (N_13415,N_13122,N_13075);
or U13416 (N_13416,N_13187,N_13011);
and U13417 (N_13417,N_12974,N_13170);
or U13418 (N_13418,N_12940,N_12933);
xnor U13419 (N_13419,N_13137,N_13107);
nor U13420 (N_13420,N_12940,N_13035);
and U13421 (N_13421,N_13031,N_13139);
nand U13422 (N_13422,N_13001,N_13014);
or U13423 (N_13423,N_12964,N_13005);
nor U13424 (N_13424,N_13066,N_13186);
nor U13425 (N_13425,N_12908,N_13129);
or U13426 (N_13426,N_13075,N_13165);
nor U13427 (N_13427,N_13037,N_13137);
nand U13428 (N_13428,N_13035,N_13086);
and U13429 (N_13429,N_12921,N_12956);
and U13430 (N_13430,N_13149,N_13044);
nand U13431 (N_13431,N_13096,N_13071);
xnor U13432 (N_13432,N_13035,N_13038);
or U13433 (N_13433,N_13149,N_13143);
nand U13434 (N_13434,N_13105,N_13112);
or U13435 (N_13435,N_13171,N_12928);
xor U13436 (N_13436,N_13187,N_13094);
nand U13437 (N_13437,N_12969,N_12966);
nand U13438 (N_13438,N_13041,N_13108);
and U13439 (N_13439,N_13026,N_12959);
nand U13440 (N_13440,N_13192,N_12907);
nand U13441 (N_13441,N_12916,N_13004);
and U13442 (N_13442,N_13155,N_12953);
nor U13443 (N_13443,N_13142,N_12918);
nand U13444 (N_13444,N_13157,N_13144);
nor U13445 (N_13445,N_13044,N_12965);
and U13446 (N_13446,N_13038,N_13158);
or U13447 (N_13447,N_13028,N_13006);
or U13448 (N_13448,N_13019,N_13171);
and U13449 (N_13449,N_13023,N_13087);
xor U13450 (N_13450,N_13075,N_13104);
and U13451 (N_13451,N_12954,N_13198);
and U13452 (N_13452,N_13067,N_13084);
and U13453 (N_13453,N_13019,N_13067);
or U13454 (N_13454,N_12962,N_12943);
nand U13455 (N_13455,N_12922,N_13067);
nand U13456 (N_13456,N_13130,N_12969);
nor U13457 (N_13457,N_13016,N_12934);
xor U13458 (N_13458,N_13019,N_13094);
and U13459 (N_13459,N_12943,N_13100);
nor U13460 (N_13460,N_13051,N_13025);
nand U13461 (N_13461,N_13093,N_13080);
nand U13462 (N_13462,N_13147,N_13105);
or U13463 (N_13463,N_12967,N_12917);
nor U13464 (N_13464,N_13189,N_12945);
and U13465 (N_13465,N_12965,N_12981);
nor U13466 (N_13466,N_13195,N_13041);
nor U13467 (N_13467,N_12940,N_13077);
xor U13468 (N_13468,N_13126,N_13154);
or U13469 (N_13469,N_13140,N_13138);
xnor U13470 (N_13470,N_13105,N_12903);
nor U13471 (N_13471,N_13083,N_13061);
and U13472 (N_13472,N_13100,N_13071);
nor U13473 (N_13473,N_12943,N_13012);
nor U13474 (N_13474,N_13108,N_12997);
xor U13475 (N_13475,N_13032,N_13151);
nand U13476 (N_13476,N_12929,N_13105);
nor U13477 (N_13477,N_13085,N_13076);
xnor U13478 (N_13478,N_13061,N_13088);
and U13479 (N_13479,N_12988,N_13167);
nor U13480 (N_13480,N_13087,N_12922);
nor U13481 (N_13481,N_13093,N_13109);
xnor U13482 (N_13482,N_13039,N_13133);
and U13483 (N_13483,N_12998,N_13052);
nand U13484 (N_13484,N_13010,N_13058);
and U13485 (N_13485,N_13122,N_13149);
xor U13486 (N_13486,N_13121,N_13113);
and U13487 (N_13487,N_13086,N_13148);
and U13488 (N_13488,N_12928,N_13009);
or U13489 (N_13489,N_13016,N_13053);
nor U13490 (N_13490,N_13032,N_13170);
nor U13491 (N_13491,N_13032,N_12968);
xor U13492 (N_13492,N_12949,N_13134);
nor U13493 (N_13493,N_13089,N_13162);
and U13494 (N_13494,N_13093,N_13132);
or U13495 (N_13495,N_13150,N_12962);
and U13496 (N_13496,N_12993,N_12962);
and U13497 (N_13497,N_12959,N_12952);
nand U13498 (N_13498,N_13010,N_13099);
and U13499 (N_13499,N_13184,N_13047);
nor U13500 (N_13500,N_13433,N_13251);
and U13501 (N_13501,N_13217,N_13229);
nor U13502 (N_13502,N_13237,N_13289);
xor U13503 (N_13503,N_13452,N_13282);
xor U13504 (N_13504,N_13419,N_13395);
xor U13505 (N_13505,N_13252,N_13448);
or U13506 (N_13506,N_13353,N_13284);
nand U13507 (N_13507,N_13455,N_13478);
nor U13508 (N_13508,N_13427,N_13440);
nor U13509 (N_13509,N_13241,N_13230);
nor U13510 (N_13510,N_13285,N_13415);
and U13511 (N_13511,N_13441,N_13363);
and U13512 (N_13512,N_13403,N_13453);
and U13513 (N_13513,N_13393,N_13439);
and U13514 (N_13514,N_13208,N_13288);
xor U13515 (N_13515,N_13343,N_13316);
nor U13516 (N_13516,N_13220,N_13374);
xnor U13517 (N_13517,N_13221,N_13405);
nand U13518 (N_13518,N_13400,N_13386);
nor U13519 (N_13519,N_13227,N_13224);
or U13520 (N_13520,N_13368,N_13218);
xnor U13521 (N_13521,N_13246,N_13488);
nor U13522 (N_13522,N_13387,N_13454);
xnor U13523 (N_13523,N_13333,N_13490);
and U13524 (N_13524,N_13260,N_13381);
or U13525 (N_13525,N_13446,N_13347);
nor U13526 (N_13526,N_13301,N_13264);
nor U13527 (N_13527,N_13366,N_13384);
nand U13528 (N_13528,N_13329,N_13385);
and U13529 (N_13529,N_13402,N_13444);
nand U13530 (N_13530,N_13468,N_13323);
and U13531 (N_13531,N_13438,N_13349);
and U13532 (N_13532,N_13355,N_13397);
nand U13533 (N_13533,N_13437,N_13473);
and U13534 (N_13534,N_13216,N_13272);
nand U13535 (N_13535,N_13350,N_13319);
or U13536 (N_13536,N_13352,N_13201);
nor U13537 (N_13537,N_13461,N_13431);
and U13538 (N_13538,N_13327,N_13214);
or U13539 (N_13539,N_13481,N_13424);
and U13540 (N_13540,N_13408,N_13429);
nand U13541 (N_13541,N_13476,N_13362);
and U13542 (N_13542,N_13256,N_13339);
nor U13543 (N_13543,N_13497,N_13228);
xnor U13544 (N_13544,N_13257,N_13213);
or U13545 (N_13545,N_13279,N_13344);
or U13546 (N_13546,N_13268,N_13411);
nor U13547 (N_13547,N_13425,N_13430);
nor U13548 (N_13548,N_13434,N_13462);
xor U13549 (N_13549,N_13239,N_13467);
xor U13550 (N_13550,N_13428,N_13372);
nor U13551 (N_13551,N_13296,N_13360);
and U13552 (N_13552,N_13249,N_13305);
nand U13553 (N_13553,N_13435,N_13370);
nor U13554 (N_13554,N_13234,N_13298);
xnor U13555 (N_13555,N_13326,N_13270);
nor U13556 (N_13556,N_13422,N_13259);
xor U13557 (N_13557,N_13447,N_13375);
nand U13558 (N_13558,N_13223,N_13315);
xnor U13559 (N_13559,N_13331,N_13283);
xnor U13560 (N_13560,N_13255,N_13358);
nand U13561 (N_13561,N_13314,N_13348);
nor U13562 (N_13562,N_13373,N_13474);
and U13563 (N_13563,N_13342,N_13483);
nor U13564 (N_13564,N_13292,N_13410);
xnor U13565 (N_13565,N_13276,N_13231);
nand U13566 (N_13566,N_13357,N_13294);
and U13567 (N_13567,N_13426,N_13317);
nor U13568 (N_13568,N_13311,N_13328);
nor U13569 (N_13569,N_13356,N_13369);
or U13570 (N_13570,N_13258,N_13281);
nor U13571 (N_13571,N_13240,N_13253);
nand U13572 (N_13572,N_13287,N_13421);
or U13573 (N_13573,N_13377,N_13280);
nand U13574 (N_13574,N_13489,N_13345);
nand U13575 (N_13575,N_13307,N_13392);
nand U13576 (N_13576,N_13320,N_13406);
or U13577 (N_13577,N_13409,N_13267);
xnor U13578 (N_13578,N_13436,N_13340);
or U13579 (N_13579,N_13383,N_13236);
nand U13580 (N_13580,N_13376,N_13203);
nor U13581 (N_13581,N_13457,N_13226);
nand U13582 (N_13582,N_13346,N_13404);
xnor U13583 (N_13583,N_13337,N_13202);
and U13584 (N_13584,N_13493,N_13472);
nand U13585 (N_13585,N_13388,N_13456);
or U13586 (N_13586,N_13396,N_13313);
xor U13587 (N_13587,N_13361,N_13238);
or U13588 (N_13588,N_13443,N_13266);
xnor U13589 (N_13589,N_13277,N_13309);
nor U13590 (N_13590,N_13495,N_13354);
nor U13591 (N_13591,N_13359,N_13460);
nand U13592 (N_13592,N_13336,N_13451);
or U13593 (N_13593,N_13449,N_13338);
nor U13594 (N_13594,N_13243,N_13498);
and U13595 (N_13595,N_13310,N_13232);
nor U13596 (N_13596,N_13209,N_13269);
xor U13597 (N_13597,N_13245,N_13261);
nand U13598 (N_13598,N_13250,N_13263);
xor U13599 (N_13599,N_13205,N_13445);
and U13600 (N_13600,N_13412,N_13390);
nor U13601 (N_13601,N_13297,N_13432);
or U13602 (N_13602,N_13487,N_13278);
nand U13603 (N_13603,N_13416,N_13471);
nor U13604 (N_13604,N_13394,N_13306);
xnor U13605 (N_13605,N_13254,N_13389);
or U13606 (N_13606,N_13332,N_13450);
nand U13607 (N_13607,N_13420,N_13334);
nand U13608 (N_13608,N_13210,N_13371);
nor U13609 (N_13609,N_13423,N_13321);
and U13610 (N_13610,N_13484,N_13364);
xor U13611 (N_13611,N_13262,N_13274);
or U13612 (N_13612,N_13244,N_13464);
nor U13613 (N_13613,N_13211,N_13200);
xor U13614 (N_13614,N_13458,N_13401);
or U13615 (N_13615,N_13318,N_13414);
or U13616 (N_13616,N_13469,N_13391);
nand U13617 (N_13617,N_13293,N_13325);
nor U13618 (N_13618,N_13486,N_13499);
nand U13619 (N_13619,N_13465,N_13302);
and U13620 (N_13620,N_13398,N_13482);
xnor U13621 (N_13621,N_13379,N_13378);
xor U13622 (N_13622,N_13304,N_13242);
nor U13623 (N_13623,N_13413,N_13291);
nor U13624 (N_13624,N_13207,N_13273);
xnor U13625 (N_13625,N_13418,N_13248);
or U13626 (N_13626,N_13295,N_13417);
or U13627 (N_13627,N_13475,N_13222);
and U13628 (N_13628,N_13204,N_13496);
xnor U13629 (N_13629,N_13470,N_13480);
xor U13630 (N_13630,N_13365,N_13367);
nor U13631 (N_13631,N_13247,N_13271);
and U13632 (N_13632,N_13312,N_13300);
nor U13633 (N_13633,N_13494,N_13290);
xor U13634 (N_13634,N_13219,N_13233);
nor U13635 (N_13635,N_13206,N_13407);
nand U13636 (N_13636,N_13299,N_13442);
nand U13637 (N_13637,N_13212,N_13265);
or U13638 (N_13638,N_13330,N_13235);
nor U13639 (N_13639,N_13479,N_13322);
nand U13640 (N_13640,N_13225,N_13382);
nand U13641 (N_13641,N_13351,N_13485);
nor U13642 (N_13642,N_13275,N_13459);
or U13643 (N_13643,N_13463,N_13303);
xor U13644 (N_13644,N_13466,N_13215);
xnor U13645 (N_13645,N_13324,N_13399);
nor U13646 (N_13646,N_13477,N_13286);
nand U13647 (N_13647,N_13335,N_13308);
and U13648 (N_13648,N_13492,N_13491);
or U13649 (N_13649,N_13380,N_13341);
or U13650 (N_13650,N_13445,N_13256);
and U13651 (N_13651,N_13450,N_13294);
or U13652 (N_13652,N_13231,N_13245);
or U13653 (N_13653,N_13367,N_13385);
nor U13654 (N_13654,N_13335,N_13203);
and U13655 (N_13655,N_13336,N_13246);
or U13656 (N_13656,N_13306,N_13364);
nand U13657 (N_13657,N_13368,N_13369);
nor U13658 (N_13658,N_13360,N_13227);
or U13659 (N_13659,N_13458,N_13461);
nand U13660 (N_13660,N_13333,N_13252);
and U13661 (N_13661,N_13346,N_13348);
and U13662 (N_13662,N_13369,N_13440);
xnor U13663 (N_13663,N_13320,N_13330);
or U13664 (N_13664,N_13302,N_13392);
nor U13665 (N_13665,N_13344,N_13259);
nand U13666 (N_13666,N_13356,N_13399);
nor U13667 (N_13667,N_13414,N_13496);
and U13668 (N_13668,N_13453,N_13294);
and U13669 (N_13669,N_13295,N_13443);
or U13670 (N_13670,N_13462,N_13222);
xnor U13671 (N_13671,N_13445,N_13251);
or U13672 (N_13672,N_13227,N_13408);
and U13673 (N_13673,N_13464,N_13343);
xor U13674 (N_13674,N_13220,N_13392);
xnor U13675 (N_13675,N_13291,N_13379);
nor U13676 (N_13676,N_13362,N_13360);
xnor U13677 (N_13677,N_13461,N_13220);
nor U13678 (N_13678,N_13282,N_13398);
and U13679 (N_13679,N_13461,N_13415);
xor U13680 (N_13680,N_13481,N_13378);
xnor U13681 (N_13681,N_13286,N_13288);
nor U13682 (N_13682,N_13303,N_13367);
xor U13683 (N_13683,N_13347,N_13391);
nand U13684 (N_13684,N_13351,N_13234);
nand U13685 (N_13685,N_13450,N_13321);
xor U13686 (N_13686,N_13370,N_13265);
nand U13687 (N_13687,N_13447,N_13398);
xor U13688 (N_13688,N_13237,N_13291);
nand U13689 (N_13689,N_13315,N_13376);
or U13690 (N_13690,N_13274,N_13254);
xnor U13691 (N_13691,N_13246,N_13282);
nand U13692 (N_13692,N_13330,N_13331);
nor U13693 (N_13693,N_13458,N_13241);
nand U13694 (N_13694,N_13477,N_13335);
xnor U13695 (N_13695,N_13302,N_13263);
and U13696 (N_13696,N_13226,N_13253);
and U13697 (N_13697,N_13203,N_13314);
or U13698 (N_13698,N_13479,N_13358);
xnor U13699 (N_13699,N_13226,N_13378);
and U13700 (N_13700,N_13238,N_13208);
and U13701 (N_13701,N_13483,N_13311);
nand U13702 (N_13702,N_13484,N_13467);
or U13703 (N_13703,N_13222,N_13482);
or U13704 (N_13704,N_13414,N_13380);
or U13705 (N_13705,N_13366,N_13287);
or U13706 (N_13706,N_13357,N_13378);
and U13707 (N_13707,N_13365,N_13283);
or U13708 (N_13708,N_13269,N_13276);
nor U13709 (N_13709,N_13354,N_13365);
nor U13710 (N_13710,N_13483,N_13295);
or U13711 (N_13711,N_13380,N_13303);
xnor U13712 (N_13712,N_13456,N_13417);
nor U13713 (N_13713,N_13245,N_13454);
and U13714 (N_13714,N_13411,N_13473);
nand U13715 (N_13715,N_13336,N_13218);
nor U13716 (N_13716,N_13216,N_13442);
nand U13717 (N_13717,N_13216,N_13206);
and U13718 (N_13718,N_13435,N_13366);
xor U13719 (N_13719,N_13316,N_13390);
xnor U13720 (N_13720,N_13206,N_13385);
and U13721 (N_13721,N_13471,N_13336);
and U13722 (N_13722,N_13497,N_13287);
xor U13723 (N_13723,N_13364,N_13203);
nand U13724 (N_13724,N_13386,N_13357);
and U13725 (N_13725,N_13474,N_13457);
and U13726 (N_13726,N_13215,N_13451);
nor U13727 (N_13727,N_13408,N_13289);
nand U13728 (N_13728,N_13292,N_13337);
xnor U13729 (N_13729,N_13431,N_13498);
xnor U13730 (N_13730,N_13405,N_13437);
and U13731 (N_13731,N_13295,N_13310);
xor U13732 (N_13732,N_13304,N_13236);
nand U13733 (N_13733,N_13231,N_13371);
xor U13734 (N_13734,N_13350,N_13486);
xor U13735 (N_13735,N_13477,N_13345);
nor U13736 (N_13736,N_13427,N_13422);
xnor U13737 (N_13737,N_13335,N_13242);
nor U13738 (N_13738,N_13362,N_13214);
nor U13739 (N_13739,N_13452,N_13460);
nand U13740 (N_13740,N_13265,N_13394);
or U13741 (N_13741,N_13281,N_13369);
or U13742 (N_13742,N_13248,N_13465);
nor U13743 (N_13743,N_13271,N_13489);
or U13744 (N_13744,N_13378,N_13325);
nand U13745 (N_13745,N_13482,N_13445);
or U13746 (N_13746,N_13337,N_13396);
or U13747 (N_13747,N_13217,N_13447);
nor U13748 (N_13748,N_13312,N_13455);
nand U13749 (N_13749,N_13473,N_13399);
xor U13750 (N_13750,N_13359,N_13286);
or U13751 (N_13751,N_13372,N_13426);
or U13752 (N_13752,N_13460,N_13313);
nand U13753 (N_13753,N_13467,N_13325);
xnor U13754 (N_13754,N_13420,N_13321);
or U13755 (N_13755,N_13362,N_13220);
nor U13756 (N_13756,N_13394,N_13379);
or U13757 (N_13757,N_13209,N_13361);
and U13758 (N_13758,N_13375,N_13476);
xnor U13759 (N_13759,N_13293,N_13462);
nor U13760 (N_13760,N_13272,N_13277);
and U13761 (N_13761,N_13220,N_13279);
xor U13762 (N_13762,N_13470,N_13476);
and U13763 (N_13763,N_13298,N_13395);
xnor U13764 (N_13764,N_13205,N_13375);
xor U13765 (N_13765,N_13259,N_13489);
or U13766 (N_13766,N_13348,N_13326);
xnor U13767 (N_13767,N_13377,N_13283);
nand U13768 (N_13768,N_13368,N_13276);
or U13769 (N_13769,N_13249,N_13420);
or U13770 (N_13770,N_13483,N_13482);
and U13771 (N_13771,N_13476,N_13361);
and U13772 (N_13772,N_13263,N_13211);
nor U13773 (N_13773,N_13409,N_13315);
nor U13774 (N_13774,N_13460,N_13289);
nor U13775 (N_13775,N_13251,N_13417);
and U13776 (N_13776,N_13450,N_13446);
nor U13777 (N_13777,N_13455,N_13217);
nand U13778 (N_13778,N_13374,N_13229);
nand U13779 (N_13779,N_13416,N_13460);
nand U13780 (N_13780,N_13272,N_13256);
nor U13781 (N_13781,N_13417,N_13233);
nand U13782 (N_13782,N_13322,N_13472);
xnor U13783 (N_13783,N_13478,N_13246);
or U13784 (N_13784,N_13272,N_13339);
xnor U13785 (N_13785,N_13259,N_13310);
or U13786 (N_13786,N_13439,N_13310);
and U13787 (N_13787,N_13274,N_13475);
nand U13788 (N_13788,N_13256,N_13474);
nand U13789 (N_13789,N_13273,N_13230);
nand U13790 (N_13790,N_13220,N_13248);
xor U13791 (N_13791,N_13244,N_13340);
and U13792 (N_13792,N_13413,N_13384);
nor U13793 (N_13793,N_13335,N_13433);
or U13794 (N_13794,N_13212,N_13448);
xnor U13795 (N_13795,N_13423,N_13382);
or U13796 (N_13796,N_13222,N_13266);
xor U13797 (N_13797,N_13452,N_13272);
nor U13798 (N_13798,N_13330,N_13305);
or U13799 (N_13799,N_13367,N_13432);
and U13800 (N_13800,N_13632,N_13536);
and U13801 (N_13801,N_13791,N_13630);
or U13802 (N_13802,N_13571,N_13564);
and U13803 (N_13803,N_13595,N_13750);
and U13804 (N_13804,N_13514,N_13534);
nand U13805 (N_13805,N_13749,N_13792);
nand U13806 (N_13806,N_13707,N_13610);
nand U13807 (N_13807,N_13565,N_13548);
and U13808 (N_13808,N_13515,N_13686);
nor U13809 (N_13809,N_13611,N_13679);
nand U13810 (N_13810,N_13789,N_13698);
or U13811 (N_13811,N_13763,N_13641);
and U13812 (N_13812,N_13502,N_13725);
nand U13813 (N_13813,N_13708,N_13702);
xnor U13814 (N_13814,N_13547,N_13695);
nand U13815 (N_13815,N_13524,N_13798);
and U13816 (N_13816,N_13648,N_13793);
or U13817 (N_13817,N_13776,N_13522);
xor U13818 (N_13818,N_13628,N_13652);
nand U13819 (N_13819,N_13600,N_13533);
and U13820 (N_13820,N_13623,N_13584);
nor U13821 (N_13821,N_13604,N_13631);
and U13822 (N_13822,N_13764,N_13538);
nand U13823 (N_13823,N_13657,N_13511);
and U13824 (N_13824,N_13768,N_13517);
xor U13825 (N_13825,N_13519,N_13532);
nand U13826 (N_13826,N_13753,N_13799);
or U13827 (N_13827,N_13527,N_13762);
xor U13828 (N_13828,N_13561,N_13599);
nor U13829 (N_13829,N_13715,N_13575);
xor U13830 (N_13830,N_13562,N_13615);
or U13831 (N_13831,N_13658,N_13556);
nor U13832 (N_13832,N_13795,N_13516);
nand U13833 (N_13833,N_13784,N_13693);
nor U13834 (N_13834,N_13523,N_13714);
nor U13835 (N_13835,N_13582,N_13663);
or U13836 (N_13836,N_13744,N_13752);
or U13837 (N_13837,N_13757,N_13782);
xor U13838 (N_13838,N_13691,N_13659);
and U13839 (N_13839,N_13700,N_13509);
xnor U13840 (N_13840,N_13772,N_13669);
or U13841 (N_13841,N_13609,N_13594);
nand U13842 (N_13842,N_13797,N_13726);
nor U13843 (N_13843,N_13688,N_13718);
or U13844 (N_13844,N_13638,N_13597);
nand U13845 (N_13845,N_13767,N_13655);
nor U13846 (N_13846,N_13553,N_13760);
nand U13847 (N_13847,N_13775,N_13704);
nor U13848 (N_13848,N_13587,N_13660);
or U13849 (N_13849,N_13520,N_13625);
xor U13850 (N_13850,N_13647,N_13559);
or U13851 (N_13851,N_13709,N_13684);
nand U13852 (N_13852,N_13670,N_13745);
and U13853 (N_13853,N_13640,N_13566);
xor U13854 (N_13854,N_13737,N_13633);
and U13855 (N_13855,N_13539,N_13614);
and U13856 (N_13856,N_13560,N_13552);
nand U13857 (N_13857,N_13689,N_13579);
nand U13858 (N_13858,N_13606,N_13755);
and U13859 (N_13859,N_13507,N_13501);
or U13860 (N_13860,N_13568,N_13712);
and U13861 (N_13861,N_13710,N_13613);
and U13862 (N_13862,N_13537,N_13549);
nor U13863 (N_13863,N_13642,N_13619);
and U13864 (N_13864,N_13616,N_13621);
xnor U13865 (N_13865,N_13783,N_13681);
or U13866 (N_13866,N_13588,N_13618);
or U13867 (N_13867,N_13790,N_13774);
and U13868 (N_13868,N_13738,N_13719);
and U13869 (N_13869,N_13518,N_13504);
and U13870 (N_13870,N_13662,N_13721);
xnor U13871 (N_13871,N_13627,N_13531);
nor U13872 (N_13872,N_13730,N_13529);
nand U13873 (N_13873,N_13735,N_13664);
nand U13874 (N_13874,N_13622,N_13781);
nor U13875 (N_13875,N_13653,N_13722);
nand U13876 (N_13876,N_13505,N_13770);
and U13877 (N_13877,N_13736,N_13761);
nor U13878 (N_13878,N_13580,N_13654);
nor U13879 (N_13879,N_13794,N_13683);
xnor U13880 (N_13880,N_13777,N_13785);
nand U13881 (N_13881,N_13671,N_13593);
xnor U13882 (N_13882,N_13626,N_13605);
nor U13883 (N_13883,N_13699,N_13687);
nand U13884 (N_13884,N_13541,N_13742);
xnor U13885 (N_13885,N_13766,N_13503);
or U13886 (N_13886,N_13703,N_13754);
xnor U13887 (N_13887,N_13581,N_13577);
xnor U13888 (N_13888,N_13666,N_13747);
or U13889 (N_13889,N_13578,N_13673);
xnor U13890 (N_13890,N_13512,N_13500);
xnor U13891 (N_13891,N_13508,N_13685);
nand U13892 (N_13892,N_13780,N_13690);
xor U13893 (N_13893,N_13675,N_13574);
nand U13894 (N_13894,N_13651,N_13591);
and U13895 (N_13895,N_13724,N_13543);
nand U13896 (N_13896,N_13717,N_13680);
or U13897 (N_13897,N_13713,N_13786);
nand U13898 (N_13898,N_13546,N_13701);
or U13899 (N_13899,N_13706,N_13540);
and U13900 (N_13900,N_13567,N_13590);
nand U13901 (N_13901,N_13734,N_13759);
xor U13902 (N_13902,N_13697,N_13740);
nand U13903 (N_13903,N_13592,N_13733);
xnor U13904 (N_13904,N_13555,N_13525);
or U13905 (N_13905,N_13643,N_13674);
or U13906 (N_13906,N_13506,N_13676);
and U13907 (N_13907,N_13602,N_13526);
nor U13908 (N_13908,N_13535,N_13758);
or U13909 (N_13909,N_13765,N_13743);
or U13910 (N_13910,N_13668,N_13645);
and U13911 (N_13911,N_13544,N_13650);
and U13912 (N_13912,N_13723,N_13705);
xnor U13913 (N_13913,N_13771,N_13569);
or U13914 (N_13914,N_13731,N_13573);
nor U13915 (N_13915,N_13557,N_13661);
xnor U13916 (N_13916,N_13624,N_13696);
nand U13917 (N_13917,N_13530,N_13551);
and U13918 (N_13918,N_13741,N_13639);
nand U13919 (N_13919,N_13598,N_13550);
nand U13920 (N_13920,N_13629,N_13711);
or U13921 (N_13921,N_13672,N_13644);
nor U13922 (N_13922,N_13788,N_13589);
nand U13923 (N_13923,N_13558,N_13528);
xnor U13924 (N_13924,N_13656,N_13545);
xor U13925 (N_13925,N_13583,N_13513);
nor U13926 (N_13926,N_13635,N_13727);
and U13927 (N_13927,N_13751,N_13612);
or U13928 (N_13928,N_13510,N_13596);
xor U13929 (N_13929,N_13720,N_13521);
or U13930 (N_13930,N_13694,N_13787);
or U13931 (N_13931,N_13634,N_13617);
nor U13932 (N_13932,N_13620,N_13769);
and U13933 (N_13933,N_13779,N_13746);
and U13934 (N_13934,N_13716,N_13756);
and U13935 (N_13935,N_13554,N_13677);
or U13936 (N_13936,N_13692,N_13570);
nor U13937 (N_13937,N_13586,N_13748);
nand U13938 (N_13938,N_13778,N_13576);
xor U13939 (N_13939,N_13607,N_13603);
or U13940 (N_13940,N_13682,N_13665);
nand U13941 (N_13941,N_13796,N_13773);
nand U13942 (N_13942,N_13563,N_13739);
or U13943 (N_13943,N_13601,N_13729);
and U13944 (N_13944,N_13637,N_13646);
nor U13945 (N_13945,N_13542,N_13678);
nand U13946 (N_13946,N_13572,N_13585);
nand U13947 (N_13947,N_13636,N_13649);
or U13948 (N_13948,N_13608,N_13732);
and U13949 (N_13949,N_13667,N_13728);
or U13950 (N_13950,N_13686,N_13749);
nor U13951 (N_13951,N_13789,N_13787);
nand U13952 (N_13952,N_13623,N_13743);
nand U13953 (N_13953,N_13697,N_13774);
and U13954 (N_13954,N_13699,N_13778);
nor U13955 (N_13955,N_13694,N_13723);
and U13956 (N_13956,N_13729,N_13574);
xnor U13957 (N_13957,N_13794,N_13582);
xnor U13958 (N_13958,N_13671,N_13796);
and U13959 (N_13959,N_13514,N_13703);
and U13960 (N_13960,N_13766,N_13616);
and U13961 (N_13961,N_13667,N_13716);
nand U13962 (N_13962,N_13564,N_13789);
nor U13963 (N_13963,N_13746,N_13773);
and U13964 (N_13964,N_13569,N_13719);
and U13965 (N_13965,N_13607,N_13578);
nor U13966 (N_13966,N_13682,N_13625);
xor U13967 (N_13967,N_13755,N_13620);
nor U13968 (N_13968,N_13645,N_13793);
nand U13969 (N_13969,N_13771,N_13581);
and U13970 (N_13970,N_13661,N_13511);
nand U13971 (N_13971,N_13640,N_13586);
xnor U13972 (N_13972,N_13543,N_13740);
nor U13973 (N_13973,N_13745,N_13581);
nand U13974 (N_13974,N_13581,N_13736);
nor U13975 (N_13975,N_13642,N_13550);
or U13976 (N_13976,N_13652,N_13527);
nor U13977 (N_13977,N_13756,N_13701);
xor U13978 (N_13978,N_13506,N_13602);
and U13979 (N_13979,N_13774,N_13701);
or U13980 (N_13980,N_13746,N_13612);
and U13981 (N_13981,N_13758,N_13730);
nand U13982 (N_13982,N_13613,N_13602);
nand U13983 (N_13983,N_13500,N_13577);
xnor U13984 (N_13984,N_13741,N_13623);
nor U13985 (N_13985,N_13536,N_13652);
and U13986 (N_13986,N_13789,N_13794);
xor U13987 (N_13987,N_13538,N_13748);
nand U13988 (N_13988,N_13537,N_13513);
nand U13989 (N_13989,N_13557,N_13692);
nand U13990 (N_13990,N_13691,N_13675);
xnor U13991 (N_13991,N_13711,N_13578);
xnor U13992 (N_13992,N_13554,N_13585);
and U13993 (N_13993,N_13589,N_13611);
and U13994 (N_13994,N_13609,N_13755);
and U13995 (N_13995,N_13555,N_13594);
and U13996 (N_13996,N_13790,N_13586);
xnor U13997 (N_13997,N_13779,N_13651);
nand U13998 (N_13998,N_13610,N_13736);
xor U13999 (N_13999,N_13757,N_13559);
and U14000 (N_14000,N_13560,N_13640);
xnor U14001 (N_14001,N_13619,N_13656);
nor U14002 (N_14002,N_13698,N_13758);
and U14003 (N_14003,N_13697,N_13769);
and U14004 (N_14004,N_13639,N_13507);
or U14005 (N_14005,N_13539,N_13623);
nand U14006 (N_14006,N_13696,N_13600);
nor U14007 (N_14007,N_13710,N_13760);
xnor U14008 (N_14008,N_13657,N_13697);
nor U14009 (N_14009,N_13505,N_13797);
and U14010 (N_14010,N_13607,N_13712);
nand U14011 (N_14011,N_13639,N_13637);
or U14012 (N_14012,N_13571,N_13570);
xor U14013 (N_14013,N_13576,N_13796);
nand U14014 (N_14014,N_13564,N_13787);
or U14015 (N_14015,N_13697,N_13636);
or U14016 (N_14016,N_13701,N_13758);
and U14017 (N_14017,N_13588,N_13548);
nor U14018 (N_14018,N_13797,N_13547);
nand U14019 (N_14019,N_13651,N_13698);
and U14020 (N_14020,N_13670,N_13618);
xnor U14021 (N_14021,N_13779,N_13689);
or U14022 (N_14022,N_13664,N_13744);
nor U14023 (N_14023,N_13651,N_13668);
or U14024 (N_14024,N_13570,N_13730);
or U14025 (N_14025,N_13707,N_13787);
nor U14026 (N_14026,N_13677,N_13507);
or U14027 (N_14027,N_13532,N_13686);
nor U14028 (N_14028,N_13533,N_13556);
nand U14029 (N_14029,N_13719,N_13595);
nor U14030 (N_14030,N_13609,N_13507);
or U14031 (N_14031,N_13788,N_13773);
nand U14032 (N_14032,N_13715,N_13776);
nand U14033 (N_14033,N_13502,N_13595);
xor U14034 (N_14034,N_13632,N_13578);
nand U14035 (N_14035,N_13736,N_13534);
or U14036 (N_14036,N_13525,N_13650);
nand U14037 (N_14037,N_13515,N_13597);
and U14038 (N_14038,N_13596,N_13625);
xor U14039 (N_14039,N_13631,N_13743);
nor U14040 (N_14040,N_13533,N_13595);
or U14041 (N_14041,N_13670,N_13699);
nand U14042 (N_14042,N_13510,N_13672);
xnor U14043 (N_14043,N_13588,N_13676);
and U14044 (N_14044,N_13651,N_13773);
and U14045 (N_14045,N_13758,N_13774);
or U14046 (N_14046,N_13597,N_13518);
or U14047 (N_14047,N_13633,N_13700);
nor U14048 (N_14048,N_13622,N_13783);
or U14049 (N_14049,N_13586,N_13783);
and U14050 (N_14050,N_13656,N_13677);
xor U14051 (N_14051,N_13772,N_13537);
nor U14052 (N_14052,N_13681,N_13612);
or U14053 (N_14053,N_13793,N_13625);
and U14054 (N_14054,N_13607,N_13669);
xor U14055 (N_14055,N_13739,N_13567);
or U14056 (N_14056,N_13505,N_13748);
or U14057 (N_14057,N_13731,N_13635);
or U14058 (N_14058,N_13623,N_13552);
or U14059 (N_14059,N_13779,N_13668);
or U14060 (N_14060,N_13739,N_13609);
and U14061 (N_14061,N_13789,N_13776);
nor U14062 (N_14062,N_13703,N_13522);
and U14063 (N_14063,N_13599,N_13506);
nor U14064 (N_14064,N_13728,N_13683);
or U14065 (N_14065,N_13795,N_13645);
nand U14066 (N_14066,N_13606,N_13745);
or U14067 (N_14067,N_13509,N_13726);
and U14068 (N_14068,N_13632,N_13537);
nand U14069 (N_14069,N_13678,N_13739);
or U14070 (N_14070,N_13543,N_13609);
nand U14071 (N_14071,N_13679,N_13757);
nand U14072 (N_14072,N_13553,N_13500);
or U14073 (N_14073,N_13783,N_13671);
xnor U14074 (N_14074,N_13668,N_13725);
nand U14075 (N_14075,N_13776,N_13704);
nand U14076 (N_14076,N_13578,N_13692);
xnor U14077 (N_14077,N_13569,N_13640);
xnor U14078 (N_14078,N_13759,N_13669);
and U14079 (N_14079,N_13657,N_13644);
nand U14080 (N_14080,N_13578,N_13570);
and U14081 (N_14081,N_13647,N_13737);
or U14082 (N_14082,N_13730,N_13560);
and U14083 (N_14083,N_13621,N_13679);
nor U14084 (N_14084,N_13710,N_13606);
or U14085 (N_14085,N_13634,N_13512);
and U14086 (N_14086,N_13564,N_13716);
nor U14087 (N_14087,N_13620,N_13500);
nand U14088 (N_14088,N_13723,N_13649);
xnor U14089 (N_14089,N_13575,N_13675);
xor U14090 (N_14090,N_13517,N_13641);
nand U14091 (N_14091,N_13605,N_13736);
or U14092 (N_14092,N_13543,N_13523);
and U14093 (N_14093,N_13618,N_13666);
xnor U14094 (N_14094,N_13556,N_13599);
or U14095 (N_14095,N_13668,N_13763);
or U14096 (N_14096,N_13703,N_13797);
nand U14097 (N_14097,N_13725,N_13742);
xor U14098 (N_14098,N_13756,N_13691);
nand U14099 (N_14099,N_13763,N_13727);
or U14100 (N_14100,N_13998,N_14058);
and U14101 (N_14101,N_14034,N_13896);
and U14102 (N_14102,N_14078,N_13868);
xnor U14103 (N_14103,N_13826,N_14094);
or U14104 (N_14104,N_13899,N_14037);
nand U14105 (N_14105,N_13855,N_13966);
or U14106 (N_14106,N_13957,N_14067);
nor U14107 (N_14107,N_14048,N_13928);
xnor U14108 (N_14108,N_13932,N_13838);
and U14109 (N_14109,N_13940,N_14080);
nand U14110 (N_14110,N_14065,N_13997);
and U14111 (N_14111,N_13829,N_13802);
nand U14112 (N_14112,N_13999,N_14056);
or U14113 (N_14113,N_14028,N_14092);
and U14114 (N_14114,N_14042,N_13807);
and U14115 (N_14115,N_14044,N_14026);
nor U14116 (N_14116,N_13922,N_14091);
nand U14117 (N_14117,N_13936,N_13901);
xnor U14118 (N_14118,N_13929,N_13842);
nand U14119 (N_14119,N_14079,N_14033);
nor U14120 (N_14120,N_13965,N_13923);
and U14121 (N_14121,N_14064,N_13810);
and U14122 (N_14122,N_14084,N_13971);
xnor U14123 (N_14123,N_13918,N_14027);
nand U14124 (N_14124,N_13809,N_13836);
nand U14125 (N_14125,N_13849,N_13992);
nor U14126 (N_14126,N_13964,N_13900);
nand U14127 (N_14127,N_14063,N_13801);
nand U14128 (N_14128,N_14030,N_13821);
xor U14129 (N_14129,N_13831,N_14035);
xor U14130 (N_14130,N_13840,N_13917);
xor U14131 (N_14131,N_14017,N_13871);
xnor U14132 (N_14132,N_14050,N_14022);
xor U14133 (N_14133,N_13939,N_13911);
nor U14134 (N_14134,N_13956,N_13869);
nand U14135 (N_14135,N_13914,N_13908);
nor U14136 (N_14136,N_14066,N_14016);
nand U14137 (N_14137,N_13866,N_13882);
nor U14138 (N_14138,N_13806,N_13909);
xnor U14139 (N_14139,N_13843,N_13990);
nor U14140 (N_14140,N_13867,N_14020);
nor U14141 (N_14141,N_13820,N_13972);
or U14142 (N_14142,N_14073,N_13979);
and U14143 (N_14143,N_13920,N_13891);
nand U14144 (N_14144,N_13904,N_14013);
and U14145 (N_14145,N_13950,N_14051);
nand U14146 (N_14146,N_13839,N_13879);
xor U14147 (N_14147,N_13814,N_13994);
or U14148 (N_14148,N_14006,N_14015);
xor U14149 (N_14149,N_14099,N_14062);
nand U14150 (N_14150,N_13969,N_14086);
nand U14151 (N_14151,N_13827,N_13945);
or U14152 (N_14152,N_13958,N_13895);
nor U14153 (N_14153,N_13986,N_13984);
and U14154 (N_14154,N_13991,N_14089);
nand U14155 (N_14155,N_13851,N_13805);
or U14156 (N_14156,N_13877,N_13937);
and U14157 (N_14157,N_13906,N_13872);
and U14158 (N_14158,N_13980,N_13876);
nor U14159 (N_14159,N_14003,N_13886);
nor U14160 (N_14160,N_13856,N_13907);
nand U14161 (N_14161,N_14008,N_13847);
nand U14162 (N_14162,N_13925,N_14085);
xnor U14163 (N_14163,N_13853,N_13949);
xor U14164 (N_14164,N_14096,N_13861);
xor U14165 (N_14165,N_14031,N_13863);
xnor U14166 (N_14166,N_14018,N_13926);
and U14167 (N_14167,N_13915,N_13808);
nand U14168 (N_14168,N_14081,N_14002);
and U14169 (N_14169,N_14069,N_13995);
and U14170 (N_14170,N_13976,N_13977);
or U14171 (N_14171,N_13996,N_13848);
nor U14172 (N_14172,N_14093,N_13864);
and U14173 (N_14173,N_14040,N_14074);
or U14174 (N_14174,N_13817,N_13973);
nand U14175 (N_14175,N_14047,N_14041);
nand U14176 (N_14176,N_13874,N_14024);
xor U14177 (N_14177,N_13852,N_13883);
nand U14178 (N_14178,N_13885,N_14057);
and U14179 (N_14179,N_13968,N_14010);
nor U14180 (N_14180,N_13858,N_14049);
and U14181 (N_14181,N_13884,N_13850);
nand U14182 (N_14182,N_14097,N_13963);
or U14183 (N_14183,N_14083,N_13913);
nand U14184 (N_14184,N_13889,N_13832);
nand U14185 (N_14185,N_13897,N_14001);
nor U14186 (N_14186,N_13961,N_14023);
and U14187 (N_14187,N_13955,N_14004);
or U14188 (N_14188,N_13875,N_13919);
or U14189 (N_14189,N_14068,N_13934);
nor U14190 (N_14190,N_14087,N_13844);
and U14191 (N_14191,N_14070,N_13902);
nand U14192 (N_14192,N_13892,N_13974);
or U14193 (N_14193,N_13824,N_13878);
xor U14194 (N_14194,N_14007,N_13951);
nand U14195 (N_14195,N_13845,N_13981);
nor U14196 (N_14196,N_13888,N_13912);
or U14197 (N_14197,N_13816,N_13818);
nand U14198 (N_14198,N_13825,N_13947);
or U14199 (N_14199,N_14019,N_13959);
nand U14200 (N_14200,N_13975,N_13946);
or U14201 (N_14201,N_13983,N_14025);
nand U14202 (N_14202,N_13828,N_13989);
or U14203 (N_14203,N_13930,N_13887);
nand U14204 (N_14204,N_13948,N_14055);
nand U14205 (N_14205,N_13938,N_13860);
nor U14206 (N_14206,N_13835,N_13812);
and U14207 (N_14207,N_13944,N_13987);
or U14208 (N_14208,N_14098,N_14052);
or U14209 (N_14209,N_13837,N_14000);
nand U14210 (N_14210,N_14009,N_13881);
nand U14211 (N_14211,N_14012,N_14077);
xor U14212 (N_14212,N_14095,N_13880);
or U14213 (N_14213,N_13953,N_14021);
or U14214 (N_14214,N_13873,N_13931);
or U14215 (N_14215,N_13985,N_13903);
xnor U14216 (N_14216,N_14029,N_14082);
and U14217 (N_14217,N_13833,N_13846);
or U14218 (N_14218,N_13962,N_13830);
or U14219 (N_14219,N_13890,N_13927);
or U14220 (N_14220,N_13822,N_14038);
nor U14221 (N_14221,N_13854,N_13910);
or U14222 (N_14222,N_13815,N_13811);
nand U14223 (N_14223,N_13935,N_14090);
nand U14224 (N_14224,N_13803,N_14043);
xor U14225 (N_14225,N_13819,N_13941);
xnor U14226 (N_14226,N_13933,N_14060);
nor U14227 (N_14227,N_14045,N_14014);
and U14228 (N_14228,N_14072,N_13859);
and U14229 (N_14229,N_14088,N_13894);
or U14230 (N_14230,N_13982,N_13841);
xor U14231 (N_14231,N_13988,N_13857);
nand U14232 (N_14232,N_13967,N_13800);
and U14233 (N_14233,N_13865,N_13954);
nand U14234 (N_14234,N_13960,N_13916);
xor U14235 (N_14235,N_13898,N_14011);
xor U14236 (N_14236,N_13862,N_13834);
xnor U14237 (N_14237,N_13978,N_13823);
xnor U14238 (N_14238,N_14071,N_13993);
nor U14239 (N_14239,N_13804,N_13924);
nor U14240 (N_14240,N_13893,N_14061);
nor U14241 (N_14241,N_13942,N_14053);
nor U14242 (N_14242,N_13943,N_13952);
xor U14243 (N_14243,N_14076,N_14036);
nor U14244 (N_14244,N_14005,N_13970);
nand U14245 (N_14245,N_14075,N_13921);
or U14246 (N_14246,N_13813,N_13905);
nand U14247 (N_14247,N_14054,N_14059);
nand U14248 (N_14248,N_14046,N_14032);
xor U14249 (N_14249,N_13870,N_14039);
or U14250 (N_14250,N_13943,N_13904);
nand U14251 (N_14251,N_13831,N_13965);
and U14252 (N_14252,N_13834,N_13892);
nor U14253 (N_14253,N_14050,N_13984);
nor U14254 (N_14254,N_13967,N_13958);
xor U14255 (N_14255,N_13900,N_14081);
nand U14256 (N_14256,N_13889,N_13860);
xor U14257 (N_14257,N_13944,N_13985);
nand U14258 (N_14258,N_13813,N_14012);
and U14259 (N_14259,N_13937,N_13846);
xor U14260 (N_14260,N_13999,N_13964);
or U14261 (N_14261,N_13803,N_14032);
or U14262 (N_14262,N_14084,N_13892);
nand U14263 (N_14263,N_13839,N_13908);
nand U14264 (N_14264,N_13816,N_13882);
nor U14265 (N_14265,N_13974,N_14086);
nand U14266 (N_14266,N_13844,N_13886);
or U14267 (N_14267,N_13990,N_13909);
or U14268 (N_14268,N_13974,N_14040);
and U14269 (N_14269,N_13847,N_13818);
nor U14270 (N_14270,N_13904,N_14027);
nor U14271 (N_14271,N_13875,N_13944);
or U14272 (N_14272,N_13882,N_13822);
or U14273 (N_14273,N_13909,N_14024);
nor U14274 (N_14274,N_13819,N_14012);
and U14275 (N_14275,N_14092,N_13881);
nor U14276 (N_14276,N_13939,N_13833);
xnor U14277 (N_14277,N_13861,N_13821);
xnor U14278 (N_14278,N_13959,N_13943);
nand U14279 (N_14279,N_14043,N_13889);
and U14280 (N_14280,N_13815,N_13985);
nand U14281 (N_14281,N_13995,N_13857);
xnor U14282 (N_14282,N_14034,N_14025);
and U14283 (N_14283,N_14016,N_13903);
nor U14284 (N_14284,N_13935,N_14075);
nor U14285 (N_14285,N_14005,N_13954);
or U14286 (N_14286,N_13926,N_13871);
nand U14287 (N_14287,N_13822,N_14024);
nor U14288 (N_14288,N_13995,N_14008);
nor U14289 (N_14289,N_13985,N_13892);
nand U14290 (N_14290,N_13958,N_13925);
nand U14291 (N_14291,N_14086,N_13815);
or U14292 (N_14292,N_13825,N_14042);
xnor U14293 (N_14293,N_13920,N_14048);
or U14294 (N_14294,N_13869,N_14031);
nand U14295 (N_14295,N_13800,N_13966);
xor U14296 (N_14296,N_13880,N_14093);
nor U14297 (N_14297,N_13889,N_14082);
nand U14298 (N_14298,N_13841,N_14081);
nor U14299 (N_14299,N_13957,N_13819);
nor U14300 (N_14300,N_13843,N_13955);
or U14301 (N_14301,N_13960,N_13838);
and U14302 (N_14302,N_13856,N_14086);
or U14303 (N_14303,N_14056,N_14008);
nand U14304 (N_14304,N_13920,N_14083);
and U14305 (N_14305,N_13830,N_13831);
nor U14306 (N_14306,N_13877,N_13802);
and U14307 (N_14307,N_13993,N_13972);
xor U14308 (N_14308,N_13899,N_13967);
nor U14309 (N_14309,N_13825,N_13840);
and U14310 (N_14310,N_13871,N_13902);
or U14311 (N_14311,N_13887,N_13873);
and U14312 (N_14312,N_13856,N_13924);
and U14313 (N_14313,N_14021,N_13987);
or U14314 (N_14314,N_13981,N_13918);
nand U14315 (N_14315,N_13881,N_14013);
nand U14316 (N_14316,N_13940,N_13849);
xnor U14317 (N_14317,N_13883,N_13931);
nor U14318 (N_14318,N_13842,N_13970);
nor U14319 (N_14319,N_13870,N_13946);
xnor U14320 (N_14320,N_13945,N_14040);
or U14321 (N_14321,N_13826,N_14077);
and U14322 (N_14322,N_13929,N_13936);
xnor U14323 (N_14323,N_13924,N_13890);
nand U14324 (N_14324,N_13943,N_13933);
nand U14325 (N_14325,N_14016,N_13832);
and U14326 (N_14326,N_14037,N_13846);
and U14327 (N_14327,N_13832,N_13834);
xor U14328 (N_14328,N_13895,N_14005);
nand U14329 (N_14329,N_14038,N_13927);
xor U14330 (N_14330,N_13867,N_14016);
nor U14331 (N_14331,N_13828,N_13844);
nand U14332 (N_14332,N_13993,N_13872);
nand U14333 (N_14333,N_13843,N_13879);
xnor U14334 (N_14334,N_13978,N_14052);
nand U14335 (N_14335,N_14055,N_13985);
or U14336 (N_14336,N_14037,N_13971);
or U14337 (N_14337,N_14024,N_13966);
or U14338 (N_14338,N_13957,N_13847);
or U14339 (N_14339,N_14045,N_13964);
nand U14340 (N_14340,N_13836,N_13969);
xor U14341 (N_14341,N_14033,N_13901);
nor U14342 (N_14342,N_13909,N_14082);
xor U14343 (N_14343,N_14047,N_14003);
and U14344 (N_14344,N_13980,N_13862);
or U14345 (N_14345,N_13806,N_13991);
nand U14346 (N_14346,N_14079,N_13987);
xor U14347 (N_14347,N_14094,N_13843);
and U14348 (N_14348,N_13970,N_14015);
or U14349 (N_14349,N_13873,N_13962);
or U14350 (N_14350,N_13892,N_13940);
and U14351 (N_14351,N_13873,N_13899);
nand U14352 (N_14352,N_14042,N_13969);
nand U14353 (N_14353,N_13879,N_13940);
or U14354 (N_14354,N_14098,N_13950);
nand U14355 (N_14355,N_14009,N_13871);
xor U14356 (N_14356,N_13926,N_13911);
or U14357 (N_14357,N_13838,N_13840);
nor U14358 (N_14358,N_13854,N_13919);
or U14359 (N_14359,N_13869,N_13950);
and U14360 (N_14360,N_13928,N_14077);
and U14361 (N_14361,N_14082,N_14022);
nand U14362 (N_14362,N_13919,N_13820);
or U14363 (N_14363,N_13812,N_13816);
or U14364 (N_14364,N_13820,N_13977);
xor U14365 (N_14365,N_13896,N_13933);
xor U14366 (N_14366,N_14074,N_13854);
or U14367 (N_14367,N_13966,N_13880);
or U14368 (N_14368,N_13813,N_13961);
nand U14369 (N_14369,N_13838,N_13820);
xor U14370 (N_14370,N_13833,N_13845);
xnor U14371 (N_14371,N_13850,N_13995);
and U14372 (N_14372,N_13992,N_13855);
nand U14373 (N_14373,N_14052,N_13882);
nor U14374 (N_14374,N_14071,N_13928);
or U14375 (N_14375,N_13948,N_13942);
xnor U14376 (N_14376,N_14037,N_13860);
nand U14377 (N_14377,N_14007,N_14066);
and U14378 (N_14378,N_13858,N_13966);
and U14379 (N_14379,N_13965,N_13985);
or U14380 (N_14380,N_14043,N_14059);
nand U14381 (N_14381,N_13829,N_13997);
or U14382 (N_14382,N_13988,N_13822);
xor U14383 (N_14383,N_13975,N_13813);
or U14384 (N_14384,N_13884,N_13959);
xnor U14385 (N_14385,N_14096,N_13815);
xnor U14386 (N_14386,N_14080,N_13858);
nand U14387 (N_14387,N_13823,N_13809);
or U14388 (N_14388,N_13961,N_14061);
nand U14389 (N_14389,N_13867,N_14036);
nand U14390 (N_14390,N_13827,N_13934);
and U14391 (N_14391,N_14015,N_13865);
nor U14392 (N_14392,N_14082,N_13991);
xnor U14393 (N_14393,N_14078,N_13839);
nand U14394 (N_14394,N_14002,N_14006);
and U14395 (N_14395,N_13856,N_13817);
nand U14396 (N_14396,N_13934,N_14061);
and U14397 (N_14397,N_13863,N_14083);
xor U14398 (N_14398,N_14064,N_13833);
nor U14399 (N_14399,N_13882,N_14084);
xnor U14400 (N_14400,N_14156,N_14366);
xor U14401 (N_14401,N_14354,N_14157);
nor U14402 (N_14402,N_14172,N_14103);
nand U14403 (N_14403,N_14260,N_14137);
nor U14404 (N_14404,N_14146,N_14292);
and U14405 (N_14405,N_14198,N_14286);
nor U14406 (N_14406,N_14100,N_14193);
xnor U14407 (N_14407,N_14110,N_14296);
or U14408 (N_14408,N_14135,N_14192);
or U14409 (N_14409,N_14186,N_14324);
xor U14410 (N_14410,N_14267,N_14302);
nor U14411 (N_14411,N_14344,N_14180);
xor U14412 (N_14412,N_14177,N_14219);
and U14413 (N_14413,N_14250,N_14353);
or U14414 (N_14414,N_14212,N_14343);
nand U14415 (N_14415,N_14358,N_14339);
nor U14416 (N_14416,N_14317,N_14216);
nor U14417 (N_14417,N_14380,N_14308);
nor U14418 (N_14418,N_14179,N_14159);
and U14419 (N_14419,N_14351,N_14230);
nand U14420 (N_14420,N_14112,N_14222);
and U14421 (N_14421,N_14106,N_14122);
nand U14422 (N_14422,N_14356,N_14300);
nand U14423 (N_14423,N_14322,N_14334);
nor U14424 (N_14424,N_14151,N_14191);
and U14425 (N_14425,N_14117,N_14301);
or U14426 (N_14426,N_14252,N_14272);
or U14427 (N_14427,N_14237,N_14357);
xnor U14428 (N_14428,N_14297,N_14349);
and U14429 (N_14429,N_14384,N_14347);
and U14430 (N_14430,N_14206,N_14285);
and U14431 (N_14431,N_14398,N_14383);
xor U14432 (N_14432,N_14160,N_14319);
xor U14433 (N_14433,N_14367,N_14214);
xnor U14434 (N_14434,N_14305,N_14276);
nor U14435 (N_14435,N_14239,N_14107);
or U14436 (N_14436,N_14229,N_14119);
nand U14437 (N_14437,N_14217,N_14307);
nand U14438 (N_14438,N_14251,N_14105);
and U14439 (N_14439,N_14310,N_14150);
nand U14440 (N_14440,N_14277,N_14389);
xnor U14441 (N_14441,N_14234,N_14364);
and U14442 (N_14442,N_14218,N_14371);
nor U14443 (N_14443,N_14397,N_14162);
nand U14444 (N_14444,N_14329,N_14320);
nand U14445 (N_14445,N_14393,N_14265);
or U14446 (N_14446,N_14153,N_14326);
xnor U14447 (N_14447,N_14164,N_14295);
and U14448 (N_14448,N_14205,N_14166);
xnor U14449 (N_14449,N_14221,N_14182);
nor U14450 (N_14450,N_14394,N_14256);
nand U14451 (N_14451,N_14130,N_14184);
and U14452 (N_14452,N_14174,N_14284);
nor U14453 (N_14453,N_14176,N_14139);
and U14454 (N_14454,N_14323,N_14138);
or U14455 (N_14455,N_14315,N_14396);
nor U14456 (N_14456,N_14104,N_14243);
xnor U14457 (N_14457,N_14126,N_14152);
or U14458 (N_14458,N_14111,N_14370);
and U14459 (N_14459,N_14224,N_14211);
xor U14460 (N_14460,N_14312,N_14361);
or U14461 (N_14461,N_14337,N_14376);
xor U14462 (N_14462,N_14365,N_14269);
and U14463 (N_14463,N_14227,N_14259);
nand U14464 (N_14464,N_14142,N_14262);
xor U14465 (N_14465,N_14318,N_14147);
nand U14466 (N_14466,N_14289,N_14283);
nor U14467 (N_14467,N_14330,N_14125);
or U14468 (N_14468,N_14258,N_14145);
and U14469 (N_14469,N_14309,N_14209);
or U14470 (N_14470,N_14321,N_14197);
and U14471 (N_14471,N_14187,N_14331);
xor U14472 (N_14472,N_14228,N_14399);
xnor U14473 (N_14473,N_14195,N_14378);
nand U14474 (N_14474,N_14253,N_14175);
nand U14475 (N_14475,N_14379,N_14372);
nor U14476 (N_14476,N_14332,N_14141);
and U14477 (N_14477,N_14304,N_14368);
or U14478 (N_14478,N_14140,N_14223);
or U14479 (N_14479,N_14385,N_14255);
or U14480 (N_14480,N_14220,N_14345);
xnor U14481 (N_14481,N_14133,N_14363);
nor U14482 (N_14482,N_14204,N_14185);
and U14483 (N_14483,N_14178,N_14254);
nand U14484 (N_14484,N_14116,N_14173);
nand U14485 (N_14485,N_14248,N_14278);
and U14486 (N_14486,N_14266,N_14226);
and U14487 (N_14487,N_14240,N_14327);
or U14488 (N_14488,N_14294,N_14114);
xnor U14489 (N_14489,N_14281,N_14246);
xnor U14490 (N_14490,N_14121,N_14355);
nand U14491 (N_14491,N_14293,N_14338);
or U14492 (N_14492,N_14275,N_14168);
and U14493 (N_14493,N_14188,N_14148);
nor U14494 (N_14494,N_14328,N_14313);
xor U14495 (N_14495,N_14316,N_14369);
or U14496 (N_14496,N_14291,N_14333);
or U14497 (N_14497,N_14348,N_14299);
xnor U14498 (N_14498,N_14123,N_14392);
or U14499 (N_14499,N_14245,N_14249);
or U14500 (N_14500,N_14235,N_14196);
and U14501 (N_14501,N_14274,N_14388);
and U14502 (N_14502,N_14203,N_14233);
nand U14503 (N_14503,N_14264,N_14390);
and U14504 (N_14504,N_14163,N_14181);
nand U14505 (N_14505,N_14215,N_14335);
and U14506 (N_14506,N_14108,N_14341);
nand U14507 (N_14507,N_14238,N_14134);
nor U14508 (N_14508,N_14136,N_14287);
and U14509 (N_14509,N_14336,N_14381);
xor U14510 (N_14510,N_14382,N_14373);
xor U14511 (N_14511,N_14201,N_14167);
nand U14512 (N_14512,N_14387,N_14242);
nand U14513 (N_14513,N_14377,N_14340);
nor U14514 (N_14514,N_14247,N_14360);
nor U14515 (N_14515,N_14257,N_14231);
or U14516 (N_14516,N_14132,N_14325);
nor U14517 (N_14517,N_14158,N_14165);
nand U14518 (N_14518,N_14261,N_14194);
nand U14519 (N_14519,N_14189,N_14359);
nor U14520 (N_14520,N_14352,N_14118);
nor U14521 (N_14521,N_14200,N_14115);
or U14522 (N_14522,N_14346,N_14244);
and U14523 (N_14523,N_14311,N_14109);
or U14524 (N_14524,N_14171,N_14155);
nor U14525 (N_14525,N_14232,N_14350);
or U14526 (N_14526,N_14131,N_14386);
nand U14527 (N_14527,N_14213,N_14273);
nor U14528 (N_14528,N_14236,N_14270);
nor U14529 (N_14529,N_14170,N_14263);
xnor U14530 (N_14530,N_14101,N_14144);
nand U14531 (N_14531,N_14303,N_14342);
or U14532 (N_14532,N_14225,N_14102);
xor U14533 (N_14533,N_14143,N_14290);
or U14534 (N_14534,N_14161,N_14314);
or U14535 (N_14535,N_14395,N_14183);
nor U14536 (N_14536,N_14120,N_14374);
nor U14537 (N_14537,N_14154,N_14288);
and U14538 (N_14538,N_14210,N_14241);
nor U14539 (N_14539,N_14124,N_14375);
nand U14540 (N_14540,N_14190,N_14282);
or U14541 (N_14541,N_14149,N_14129);
nand U14542 (N_14542,N_14362,N_14268);
and U14543 (N_14543,N_14208,N_14202);
and U14544 (N_14544,N_14271,N_14298);
or U14545 (N_14545,N_14169,N_14128);
nand U14546 (N_14546,N_14279,N_14280);
nand U14547 (N_14547,N_14306,N_14207);
or U14548 (N_14548,N_14199,N_14113);
nor U14549 (N_14549,N_14127,N_14391);
xnor U14550 (N_14550,N_14209,N_14389);
nor U14551 (N_14551,N_14316,N_14382);
or U14552 (N_14552,N_14327,N_14123);
nor U14553 (N_14553,N_14288,N_14389);
xnor U14554 (N_14554,N_14340,N_14252);
nand U14555 (N_14555,N_14226,N_14282);
nor U14556 (N_14556,N_14231,N_14166);
nand U14557 (N_14557,N_14286,N_14258);
nor U14558 (N_14558,N_14187,N_14267);
nor U14559 (N_14559,N_14163,N_14178);
nor U14560 (N_14560,N_14329,N_14367);
nor U14561 (N_14561,N_14116,N_14168);
or U14562 (N_14562,N_14351,N_14343);
or U14563 (N_14563,N_14334,N_14141);
nand U14564 (N_14564,N_14147,N_14365);
xor U14565 (N_14565,N_14343,N_14120);
or U14566 (N_14566,N_14351,N_14332);
xnor U14567 (N_14567,N_14182,N_14370);
nor U14568 (N_14568,N_14118,N_14136);
or U14569 (N_14569,N_14331,N_14372);
nand U14570 (N_14570,N_14341,N_14154);
nand U14571 (N_14571,N_14326,N_14285);
and U14572 (N_14572,N_14395,N_14158);
xnor U14573 (N_14573,N_14225,N_14203);
nand U14574 (N_14574,N_14161,N_14276);
nor U14575 (N_14575,N_14186,N_14252);
xor U14576 (N_14576,N_14383,N_14219);
xnor U14577 (N_14577,N_14109,N_14172);
xnor U14578 (N_14578,N_14144,N_14124);
xor U14579 (N_14579,N_14232,N_14137);
or U14580 (N_14580,N_14207,N_14394);
and U14581 (N_14581,N_14386,N_14390);
and U14582 (N_14582,N_14285,N_14338);
and U14583 (N_14583,N_14357,N_14210);
nand U14584 (N_14584,N_14258,N_14278);
and U14585 (N_14585,N_14246,N_14111);
nand U14586 (N_14586,N_14138,N_14300);
and U14587 (N_14587,N_14100,N_14366);
or U14588 (N_14588,N_14304,N_14151);
nor U14589 (N_14589,N_14145,N_14142);
or U14590 (N_14590,N_14392,N_14108);
and U14591 (N_14591,N_14345,N_14392);
or U14592 (N_14592,N_14172,N_14233);
and U14593 (N_14593,N_14353,N_14334);
or U14594 (N_14594,N_14194,N_14227);
xor U14595 (N_14595,N_14302,N_14329);
nor U14596 (N_14596,N_14162,N_14307);
and U14597 (N_14597,N_14150,N_14261);
or U14598 (N_14598,N_14225,N_14262);
nand U14599 (N_14599,N_14321,N_14161);
nand U14600 (N_14600,N_14152,N_14384);
xor U14601 (N_14601,N_14306,N_14398);
nor U14602 (N_14602,N_14148,N_14144);
xor U14603 (N_14603,N_14172,N_14346);
nor U14604 (N_14604,N_14100,N_14290);
xor U14605 (N_14605,N_14262,N_14299);
nand U14606 (N_14606,N_14143,N_14370);
xnor U14607 (N_14607,N_14170,N_14249);
xor U14608 (N_14608,N_14356,N_14117);
xor U14609 (N_14609,N_14331,N_14170);
and U14610 (N_14610,N_14273,N_14336);
xor U14611 (N_14611,N_14284,N_14118);
nor U14612 (N_14612,N_14336,N_14356);
and U14613 (N_14613,N_14173,N_14374);
xnor U14614 (N_14614,N_14100,N_14163);
and U14615 (N_14615,N_14154,N_14389);
or U14616 (N_14616,N_14242,N_14137);
nand U14617 (N_14617,N_14297,N_14129);
xnor U14618 (N_14618,N_14264,N_14298);
and U14619 (N_14619,N_14177,N_14336);
or U14620 (N_14620,N_14169,N_14373);
nor U14621 (N_14621,N_14278,N_14360);
and U14622 (N_14622,N_14150,N_14133);
or U14623 (N_14623,N_14203,N_14372);
nor U14624 (N_14624,N_14329,N_14395);
nor U14625 (N_14625,N_14245,N_14190);
nor U14626 (N_14626,N_14307,N_14296);
xor U14627 (N_14627,N_14392,N_14105);
nand U14628 (N_14628,N_14148,N_14334);
and U14629 (N_14629,N_14116,N_14224);
xor U14630 (N_14630,N_14348,N_14300);
nor U14631 (N_14631,N_14144,N_14216);
nor U14632 (N_14632,N_14248,N_14194);
xor U14633 (N_14633,N_14362,N_14390);
nor U14634 (N_14634,N_14367,N_14264);
nor U14635 (N_14635,N_14389,N_14246);
or U14636 (N_14636,N_14128,N_14240);
and U14637 (N_14637,N_14217,N_14291);
nand U14638 (N_14638,N_14334,N_14314);
nor U14639 (N_14639,N_14216,N_14292);
nor U14640 (N_14640,N_14391,N_14343);
and U14641 (N_14641,N_14246,N_14211);
xnor U14642 (N_14642,N_14273,N_14225);
and U14643 (N_14643,N_14151,N_14196);
and U14644 (N_14644,N_14208,N_14368);
xnor U14645 (N_14645,N_14150,N_14202);
nand U14646 (N_14646,N_14335,N_14116);
xnor U14647 (N_14647,N_14200,N_14218);
xnor U14648 (N_14648,N_14104,N_14257);
and U14649 (N_14649,N_14347,N_14363);
or U14650 (N_14650,N_14104,N_14265);
xnor U14651 (N_14651,N_14274,N_14225);
nand U14652 (N_14652,N_14148,N_14332);
nor U14653 (N_14653,N_14128,N_14353);
and U14654 (N_14654,N_14354,N_14190);
or U14655 (N_14655,N_14197,N_14107);
and U14656 (N_14656,N_14130,N_14245);
and U14657 (N_14657,N_14208,N_14266);
xor U14658 (N_14658,N_14163,N_14116);
nor U14659 (N_14659,N_14232,N_14191);
nor U14660 (N_14660,N_14204,N_14297);
xnor U14661 (N_14661,N_14334,N_14236);
xnor U14662 (N_14662,N_14342,N_14328);
nor U14663 (N_14663,N_14305,N_14242);
and U14664 (N_14664,N_14277,N_14354);
and U14665 (N_14665,N_14204,N_14352);
or U14666 (N_14666,N_14339,N_14379);
nor U14667 (N_14667,N_14268,N_14110);
xor U14668 (N_14668,N_14371,N_14360);
nor U14669 (N_14669,N_14289,N_14294);
nand U14670 (N_14670,N_14290,N_14397);
or U14671 (N_14671,N_14368,N_14371);
or U14672 (N_14672,N_14258,N_14180);
nand U14673 (N_14673,N_14303,N_14240);
and U14674 (N_14674,N_14243,N_14324);
or U14675 (N_14675,N_14294,N_14164);
and U14676 (N_14676,N_14364,N_14173);
nor U14677 (N_14677,N_14145,N_14390);
nand U14678 (N_14678,N_14292,N_14352);
and U14679 (N_14679,N_14128,N_14382);
xnor U14680 (N_14680,N_14363,N_14250);
xnor U14681 (N_14681,N_14361,N_14174);
nor U14682 (N_14682,N_14149,N_14154);
nor U14683 (N_14683,N_14185,N_14102);
and U14684 (N_14684,N_14302,N_14299);
xor U14685 (N_14685,N_14349,N_14397);
xnor U14686 (N_14686,N_14242,N_14254);
or U14687 (N_14687,N_14123,N_14112);
or U14688 (N_14688,N_14192,N_14113);
or U14689 (N_14689,N_14292,N_14328);
and U14690 (N_14690,N_14271,N_14283);
or U14691 (N_14691,N_14313,N_14185);
and U14692 (N_14692,N_14184,N_14158);
and U14693 (N_14693,N_14309,N_14128);
and U14694 (N_14694,N_14325,N_14347);
nor U14695 (N_14695,N_14390,N_14246);
nor U14696 (N_14696,N_14112,N_14106);
xor U14697 (N_14697,N_14312,N_14376);
nor U14698 (N_14698,N_14383,N_14164);
and U14699 (N_14699,N_14266,N_14142);
nor U14700 (N_14700,N_14694,N_14546);
xnor U14701 (N_14701,N_14418,N_14548);
or U14702 (N_14702,N_14522,N_14699);
nand U14703 (N_14703,N_14494,N_14611);
nand U14704 (N_14704,N_14527,N_14486);
nand U14705 (N_14705,N_14503,N_14679);
nand U14706 (N_14706,N_14666,N_14554);
nand U14707 (N_14707,N_14448,N_14691);
xnor U14708 (N_14708,N_14533,N_14595);
nand U14709 (N_14709,N_14464,N_14453);
or U14710 (N_14710,N_14617,N_14447);
and U14711 (N_14711,N_14521,N_14463);
xnor U14712 (N_14712,N_14585,N_14683);
xnor U14713 (N_14713,N_14504,N_14639);
nor U14714 (N_14714,N_14460,N_14698);
xor U14715 (N_14715,N_14506,N_14583);
xor U14716 (N_14716,N_14584,N_14695);
xor U14717 (N_14717,N_14515,N_14541);
xor U14718 (N_14718,N_14559,N_14627);
and U14719 (N_14719,N_14400,N_14629);
or U14720 (N_14720,N_14470,N_14525);
nor U14721 (N_14721,N_14567,N_14661);
or U14722 (N_14722,N_14674,N_14543);
and U14723 (N_14723,N_14653,N_14651);
nand U14724 (N_14724,N_14454,N_14602);
and U14725 (N_14725,N_14539,N_14505);
nand U14726 (N_14726,N_14552,N_14440);
xor U14727 (N_14727,N_14413,N_14477);
nor U14728 (N_14728,N_14474,N_14437);
nand U14729 (N_14729,N_14623,N_14451);
xor U14730 (N_14730,N_14622,N_14626);
and U14731 (N_14731,N_14564,N_14618);
or U14732 (N_14732,N_14631,N_14646);
xnor U14733 (N_14733,N_14576,N_14652);
nand U14734 (N_14734,N_14480,N_14513);
or U14735 (N_14735,N_14406,N_14607);
xor U14736 (N_14736,N_14417,N_14571);
and U14737 (N_14737,N_14514,N_14680);
or U14738 (N_14738,N_14500,N_14671);
nand U14739 (N_14739,N_14545,N_14439);
and U14740 (N_14740,N_14508,N_14697);
or U14741 (N_14741,N_14484,N_14569);
and U14742 (N_14742,N_14491,N_14628);
or U14743 (N_14743,N_14673,N_14647);
or U14744 (N_14744,N_14690,N_14497);
nand U14745 (N_14745,N_14598,N_14613);
nand U14746 (N_14746,N_14632,N_14426);
nand U14747 (N_14747,N_14416,N_14452);
or U14748 (N_14748,N_14685,N_14605);
nor U14749 (N_14749,N_14578,N_14668);
nand U14750 (N_14750,N_14434,N_14662);
nand U14751 (N_14751,N_14549,N_14458);
and U14752 (N_14752,N_14510,N_14550);
and U14753 (N_14753,N_14524,N_14502);
nand U14754 (N_14754,N_14526,N_14431);
nor U14755 (N_14755,N_14473,N_14635);
nand U14756 (N_14756,N_14696,N_14446);
or U14757 (N_14757,N_14637,N_14441);
and U14758 (N_14758,N_14620,N_14411);
nor U14759 (N_14759,N_14650,N_14475);
nor U14760 (N_14760,N_14443,N_14608);
nand U14761 (N_14761,N_14401,N_14414);
nand U14762 (N_14762,N_14444,N_14609);
xnor U14763 (N_14763,N_14459,N_14672);
xor U14764 (N_14764,N_14472,N_14469);
and U14765 (N_14765,N_14681,N_14512);
or U14766 (N_14766,N_14498,N_14540);
or U14767 (N_14767,N_14537,N_14555);
or U14768 (N_14768,N_14432,N_14493);
and U14769 (N_14769,N_14574,N_14421);
and U14770 (N_14770,N_14573,N_14656);
and U14771 (N_14771,N_14495,N_14408);
xnor U14772 (N_14772,N_14660,N_14572);
xor U14773 (N_14773,N_14509,N_14588);
xor U14774 (N_14774,N_14517,N_14667);
nor U14775 (N_14775,N_14520,N_14478);
xor U14776 (N_14776,N_14592,N_14670);
or U14777 (N_14777,N_14511,N_14496);
xnor U14778 (N_14778,N_14676,N_14445);
xnor U14779 (N_14779,N_14530,N_14677);
nand U14780 (N_14780,N_14684,N_14556);
xor U14781 (N_14781,N_14604,N_14642);
xnor U14782 (N_14782,N_14558,N_14489);
xnor U14783 (N_14783,N_14471,N_14579);
nor U14784 (N_14784,N_14577,N_14658);
nor U14785 (N_14785,N_14675,N_14553);
nor U14786 (N_14786,N_14640,N_14600);
nand U14787 (N_14787,N_14430,N_14507);
and U14788 (N_14788,N_14435,N_14534);
and U14789 (N_14789,N_14612,N_14427);
xnor U14790 (N_14790,N_14479,N_14420);
and U14791 (N_14791,N_14570,N_14467);
and U14792 (N_14792,N_14449,N_14424);
xnor U14793 (N_14793,N_14654,N_14466);
nand U14794 (N_14794,N_14663,N_14633);
nand U14795 (N_14795,N_14423,N_14538);
xor U14796 (N_14796,N_14518,N_14442);
nor U14797 (N_14797,N_14648,N_14422);
nand U14798 (N_14798,N_14415,N_14412);
nor U14799 (N_14799,N_14580,N_14641);
xor U14800 (N_14800,N_14481,N_14565);
nand U14801 (N_14801,N_14560,N_14687);
or U14802 (N_14802,N_14490,N_14410);
xor U14803 (N_14803,N_14659,N_14455);
or U14804 (N_14804,N_14566,N_14457);
nor U14805 (N_14805,N_14610,N_14599);
and U14806 (N_14806,N_14615,N_14616);
xor U14807 (N_14807,N_14499,N_14601);
or U14808 (N_14808,N_14428,N_14596);
nor U14809 (N_14809,N_14485,N_14465);
xor U14810 (N_14810,N_14531,N_14606);
or U14811 (N_14811,N_14582,N_14450);
and U14812 (N_14812,N_14678,N_14634);
and U14813 (N_14813,N_14587,N_14483);
nor U14814 (N_14814,N_14551,N_14523);
nand U14815 (N_14815,N_14542,N_14468);
and U14816 (N_14816,N_14568,N_14563);
nand U14817 (N_14817,N_14621,N_14575);
xnor U14818 (N_14818,N_14689,N_14532);
nor U14819 (N_14819,N_14589,N_14535);
nor U14820 (N_14820,N_14669,N_14603);
nor U14821 (N_14821,N_14619,N_14625);
xnor U14822 (N_14822,N_14429,N_14544);
or U14823 (N_14823,N_14593,N_14425);
xor U14824 (N_14824,N_14557,N_14492);
or U14825 (N_14825,N_14686,N_14462);
nand U14826 (N_14826,N_14402,N_14649);
xnor U14827 (N_14827,N_14403,N_14409);
and U14828 (N_14828,N_14419,N_14519);
nor U14829 (N_14829,N_14405,N_14488);
or U14830 (N_14830,N_14664,N_14645);
or U14831 (N_14831,N_14436,N_14682);
and U14832 (N_14832,N_14590,N_14614);
or U14833 (N_14833,N_14597,N_14438);
nand U14834 (N_14834,N_14636,N_14561);
nand U14835 (N_14835,N_14528,N_14536);
nor U14836 (N_14836,N_14501,N_14476);
nand U14837 (N_14837,N_14586,N_14624);
xnor U14838 (N_14838,N_14692,N_14487);
nand U14839 (N_14839,N_14594,N_14638);
xnor U14840 (N_14840,N_14482,N_14562);
nor U14841 (N_14841,N_14581,N_14657);
nand U14842 (N_14842,N_14404,N_14461);
nand U14843 (N_14843,N_14529,N_14433);
or U14844 (N_14844,N_14644,N_14643);
or U14845 (N_14845,N_14655,N_14693);
xnor U14846 (N_14846,N_14547,N_14665);
nand U14847 (N_14847,N_14407,N_14630);
or U14848 (N_14848,N_14516,N_14688);
nor U14849 (N_14849,N_14591,N_14456);
and U14850 (N_14850,N_14670,N_14533);
or U14851 (N_14851,N_14552,N_14623);
nand U14852 (N_14852,N_14669,N_14502);
nor U14853 (N_14853,N_14613,N_14661);
xor U14854 (N_14854,N_14515,N_14626);
nand U14855 (N_14855,N_14653,N_14507);
or U14856 (N_14856,N_14654,N_14600);
or U14857 (N_14857,N_14495,N_14687);
nor U14858 (N_14858,N_14544,N_14534);
or U14859 (N_14859,N_14656,N_14465);
or U14860 (N_14860,N_14497,N_14475);
nor U14861 (N_14861,N_14651,N_14692);
nor U14862 (N_14862,N_14663,N_14463);
nand U14863 (N_14863,N_14506,N_14551);
nand U14864 (N_14864,N_14478,N_14492);
nor U14865 (N_14865,N_14429,N_14445);
and U14866 (N_14866,N_14555,N_14461);
xnor U14867 (N_14867,N_14566,N_14448);
nand U14868 (N_14868,N_14683,N_14508);
or U14869 (N_14869,N_14693,N_14522);
or U14870 (N_14870,N_14576,N_14653);
and U14871 (N_14871,N_14564,N_14451);
or U14872 (N_14872,N_14638,N_14531);
or U14873 (N_14873,N_14418,N_14620);
and U14874 (N_14874,N_14601,N_14424);
nor U14875 (N_14875,N_14532,N_14435);
xnor U14876 (N_14876,N_14599,N_14675);
xor U14877 (N_14877,N_14593,N_14589);
and U14878 (N_14878,N_14667,N_14498);
nand U14879 (N_14879,N_14468,N_14474);
xor U14880 (N_14880,N_14429,N_14452);
nor U14881 (N_14881,N_14589,N_14406);
nand U14882 (N_14882,N_14650,N_14551);
nor U14883 (N_14883,N_14429,N_14562);
xnor U14884 (N_14884,N_14408,N_14516);
and U14885 (N_14885,N_14649,N_14445);
xor U14886 (N_14886,N_14421,N_14418);
and U14887 (N_14887,N_14536,N_14515);
xnor U14888 (N_14888,N_14411,N_14466);
or U14889 (N_14889,N_14674,N_14589);
nor U14890 (N_14890,N_14536,N_14538);
nand U14891 (N_14891,N_14498,N_14693);
xor U14892 (N_14892,N_14581,N_14449);
or U14893 (N_14893,N_14667,N_14478);
or U14894 (N_14894,N_14521,N_14542);
xnor U14895 (N_14895,N_14418,N_14450);
xnor U14896 (N_14896,N_14451,N_14604);
nor U14897 (N_14897,N_14650,N_14519);
nor U14898 (N_14898,N_14686,N_14605);
nand U14899 (N_14899,N_14431,N_14474);
or U14900 (N_14900,N_14460,N_14687);
and U14901 (N_14901,N_14568,N_14586);
nor U14902 (N_14902,N_14625,N_14517);
nand U14903 (N_14903,N_14495,N_14420);
or U14904 (N_14904,N_14409,N_14625);
or U14905 (N_14905,N_14699,N_14524);
and U14906 (N_14906,N_14490,N_14647);
nand U14907 (N_14907,N_14630,N_14670);
or U14908 (N_14908,N_14539,N_14503);
and U14909 (N_14909,N_14419,N_14586);
and U14910 (N_14910,N_14622,N_14636);
or U14911 (N_14911,N_14647,N_14502);
and U14912 (N_14912,N_14404,N_14437);
xnor U14913 (N_14913,N_14517,N_14525);
and U14914 (N_14914,N_14494,N_14419);
or U14915 (N_14915,N_14521,N_14686);
or U14916 (N_14916,N_14428,N_14423);
or U14917 (N_14917,N_14668,N_14583);
or U14918 (N_14918,N_14665,N_14632);
xnor U14919 (N_14919,N_14560,N_14553);
or U14920 (N_14920,N_14456,N_14410);
and U14921 (N_14921,N_14420,N_14667);
and U14922 (N_14922,N_14410,N_14557);
and U14923 (N_14923,N_14640,N_14606);
nor U14924 (N_14924,N_14434,N_14613);
nand U14925 (N_14925,N_14525,N_14581);
xor U14926 (N_14926,N_14444,N_14554);
or U14927 (N_14927,N_14484,N_14513);
or U14928 (N_14928,N_14523,N_14647);
nor U14929 (N_14929,N_14535,N_14484);
nor U14930 (N_14930,N_14576,N_14414);
nand U14931 (N_14931,N_14664,N_14445);
and U14932 (N_14932,N_14554,N_14612);
nor U14933 (N_14933,N_14429,N_14468);
nand U14934 (N_14934,N_14496,N_14596);
nor U14935 (N_14935,N_14431,N_14422);
nor U14936 (N_14936,N_14441,N_14448);
nor U14937 (N_14937,N_14509,N_14506);
or U14938 (N_14938,N_14425,N_14651);
nand U14939 (N_14939,N_14422,N_14642);
xnor U14940 (N_14940,N_14557,N_14678);
and U14941 (N_14941,N_14582,N_14548);
and U14942 (N_14942,N_14427,N_14483);
and U14943 (N_14943,N_14658,N_14481);
or U14944 (N_14944,N_14515,N_14519);
nor U14945 (N_14945,N_14683,N_14686);
nand U14946 (N_14946,N_14554,N_14517);
xnor U14947 (N_14947,N_14676,N_14485);
or U14948 (N_14948,N_14497,N_14406);
xnor U14949 (N_14949,N_14671,N_14415);
nor U14950 (N_14950,N_14522,N_14564);
nor U14951 (N_14951,N_14547,N_14416);
or U14952 (N_14952,N_14612,N_14401);
and U14953 (N_14953,N_14563,N_14616);
xnor U14954 (N_14954,N_14585,N_14475);
and U14955 (N_14955,N_14695,N_14653);
nand U14956 (N_14956,N_14491,N_14677);
or U14957 (N_14957,N_14576,N_14674);
nand U14958 (N_14958,N_14537,N_14638);
nand U14959 (N_14959,N_14509,N_14564);
nand U14960 (N_14960,N_14454,N_14651);
nor U14961 (N_14961,N_14652,N_14518);
and U14962 (N_14962,N_14462,N_14593);
xor U14963 (N_14963,N_14428,N_14481);
or U14964 (N_14964,N_14546,N_14663);
xnor U14965 (N_14965,N_14659,N_14686);
or U14966 (N_14966,N_14636,N_14431);
xnor U14967 (N_14967,N_14565,N_14468);
nand U14968 (N_14968,N_14501,N_14624);
and U14969 (N_14969,N_14629,N_14489);
and U14970 (N_14970,N_14483,N_14656);
or U14971 (N_14971,N_14587,N_14639);
or U14972 (N_14972,N_14631,N_14570);
xor U14973 (N_14973,N_14568,N_14679);
nand U14974 (N_14974,N_14617,N_14581);
or U14975 (N_14975,N_14564,N_14446);
and U14976 (N_14976,N_14578,N_14409);
nor U14977 (N_14977,N_14622,N_14421);
and U14978 (N_14978,N_14424,N_14470);
nor U14979 (N_14979,N_14525,N_14439);
nand U14980 (N_14980,N_14478,N_14505);
nand U14981 (N_14981,N_14477,N_14534);
or U14982 (N_14982,N_14433,N_14688);
or U14983 (N_14983,N_14628,N_14567);
nand U14984 (N_14984,N_14513,N_14591);
xnor U14985 (N_14985,N_14539,N_14692);
or U14986 (N_14986,N_14617,N_14562);
and U14987 (N_14987,N_14521,N_14637);
nor U14988 (N_14988,N_14598,N_14545);
and U14989 (N_14989,N_14524,N_14694);
or U14990 (N_14990,N_14405,N_14433);
nor U14991 (N_14991,N_14592,N_14561);
or U14992 (N_14992,N_14679,N_14612);
nor U14993 (N_14993,N_14682,N_14480);
nand U14994 (N_14994,N_14540,N_14678);
or U14995 (N_14995,N_14589,N_14644);
nand U14996 (N_14996,N_14468,N_14415);
and U14997 (N_14997,N_14438,N_14531);
and U14998 (N_14998,N_14461,N_14559);
nor U14999 (N_14999,N_14403,N_14430);
xnor UO_0 (O_0,N_14790,N_14779);
nand UO_1 (O_1,N_14929,N_14870);
xnor UO_2 (O_2,N_14946,N_14859);
nand UO_3 (O_3,N_14727,N_14723);
and UO_4 (O_4,N_14710,N_14954);
nor UO_5 (O_5,N_14732,N_14967);
nor UO_6 (O_6,N_14939,N_14905);
or UO_7 (O_7,N_14825,N_14973);
nor UO_8 (O_8,N_14902,N_14777);
or UO_9 (O_9,N_14826,N_14885);
and UO_10 (O_10,N_14718,N_14700);
and UO_11 (O_11,N_14972,N_14838);
and UO_12 (O_12,N_14763,N_14752);
or UO_13 (O_13,N_14913,N_14909);
xnor UO_14 (O_14,N_14915,N_14994);
xnor UO_15 (O_15,N_14864,N_14962);
nand UO_16 (O_16,N_14977,N_14767);
nand UO_17 (O_17,N_14774,N_14823);
nor UO_18 (O_18,N_14854,N_14809);
nand UO_19 (O_19,N_14999,N_14773);
nor UO_20 (O_20,N_14730,N_14742);
nor UO_21 (O_21,N_14755,N_14768);
and UO_22 (O_22,N_14862,N_14898);
xnor UO_23 (O_23,N_14795,N_14948);
nor UO_24 (O_24,N_14841,N_14829);
nor UO_25 (O_25,N_14981,N_14754);
and UO_26 (O_26,N_14974,N_14934);
nand UO_27 (O_27,N_14997,N_14705);
nor UO_28 (O_28,N_14951,N_14960);
xnor UO_29 (O_29,N_14928,N_14814);
or UO_30 (O_30,N_14897,N_14964);
xnor UO_31 (O_31,N_14881,N_14764);
xnor UO_32 (O_32,N_14808,N_14707);
and UO_33 (O_33,N_14780,N_14861);
nor UO_34 (O_34,N_14832,N_14759);
or UO_35 (O_35,N_14706,N_14728);
nor UO_36 (O_36,N_14761,N_14886);
xnor UO_37 (O_37,N_14863,N_14801);
nand UO_38 (O_38,N_14800,N_14865);
xor UO_39 (O_39,N_14950,N_14855);
and UO_40 (O_40,N_14922,N_14804);
xnor UO_41 (O_41,N_14711,N_14729);
or UO_42 (O_42,N_14911,N_14715);
and UO_43 (O_43,N_14836,N_14858);
nand UO_44 (O_44,N_14724,N_14961);
xor UO_45 (O_45,N_14982,N_14888);
or UO_46 (O_46,N_14867,N_14975);
xnor UO_47 (O_47,N_14907,N_14787);
nand UO_48 (O_48,N_14916,N_14757);
xor UO_49 (O_49,N_14810,N_14903);
nor UO_50 (O_50,N_14957,N_14949);
nand UO_51 (O_51,N_14766,N_14938);
and UO_52 (O_52,N_14741,N_14802);
and UO_53 (O_53,N_14708,N_14990);
xor UO_54 (O_54,N_14896,N_14714);
and UO_55 (O_55,N_14822,N_14959);
or UO_56 (O_56,N_14993,N_14871);
or UO_57 (O_57,N_14873,N_14709);
nor UO_58 (O_58,N_14983,N_14857);
xnor UO_59 (O_59,N_14797,N_14877);
or UO_60 (O_60,N_14771,N_14904);
or UO_61 (O_61,N_14856,N_14748);
nor UO_62 (O_62,N_14936,N_14914);
or UO_63 (O_63,N_14917,N_14756);
nor UO_64 (O_64,N_14806,N_14875);
xor UO_65 (O_65,N_14783,N_14988);
nor UO_66 (O_66,N_14813,N_14719);
and UO_67 (O_67,N_14745,N_14762);
nor UO_68 (O_68,N_14733,N_14812);
or UO_69 (O_69,N_14924,N_14831);
xnor UO_70 (O_70,N_14844,N_14799);
nor UO_71 (O_71,N_14758,N_14874);
nand UO_72 (O_72,N_14891,N_14811);
nor UO_73 (O_73,N_14720,N_14930);
xor UO_74 (O_74,N_14899,N_14895);
and UO_75 (O_75,N_14869,N_14991);
or UO_76 (O_76,N_14940,N_14726);
nand UO_77 (O_77,N_14995,N_14717);
or UO_78 (O_78,N_14703,N_14821);
nor UO_79 (O_79,N_14918,N_14986);
and UO_80 (O_80,N_14743,N_14842);
xnor UO_81 (O_81,N_14912,N_14893);
nand UO_82 (O_82,N_14878,N_14947);
or UO_83 (O_83,N_14906,N_14834);
nand UO_84 (O_84,N_14933,N_14776);
and UO_85 (O_85,N_14944,N_14956);
and UO_86 (O_86,N_14910,N_14945);
xor UO_87 (O_87,N_14963,N_14998);
xnor UO_88 (O_88,N_14852,N_14704);
xnor UO_89 (O_89,N_14846,N_14890);
and UO_90 (O_90,N_14937,N_14819);
xnor UO_91 (O_91,N_14853,N_14935);
or UO_92 (O_92,N_14817,N_14750);
or UO_93 (O_93,N_14850,N_14920);
or UO_94 (O_94,N_14722,N_14820);
nand UO_95 (O_95,N_14765,N_14747);
xnor UO_96 (O_96,N_14781,N_14984);
nor UO_97 (O_97,N_14953,N_14835);
nand UO_98 (O_98,N_14721,N_14833);
nor UO_99 (O_99,N_14716,N_14943);
or UO_100 (O_100,N_14996,N_14816);
and UO_101 (O_101,N_14824,N_14968);
or UO_102 (O_102,N_14840,N_14866);
xnor UO_103 (O_103,N_14803,N_14879);
nand UO_104 (O_104,N_14839,N_14713);
nand UO_105 (O_105,N_14848,N_14805);
xor UO_106 (O_106,N_14894,N_14712);
nand UO_107 (O_107,N_14828,N_14769);
nand UO_108 (O_108,N_14753,N_14989);
and UO_109 (O_109,N_14785,N_14979);
or UO_110 (O_110,N_14900,N_14772);
xnor UO_111 (O_111,N_14749,N_14784);
nor UO_112 (O_112,N_14740,N_14731);
nor UO_113 (O_113,N_14985,N_14952);
nor UO_114 (O_114,N_14901,N_14793);
nand UO_115 (O_115,N_14889,N_14860);
nor UO_116 (O_116,N_14782,N_14966);
or UO_117 (O_117,N_14970,N_14789);
and UO_118 (O_118,N_14987,N_14791);
and UO_119 (O_119,N_14892,N_14872);
and UO_120 (O_120,N_14701,N_14926);
xor UO_121 (O_121,N_14737,N_14775);
xor UO_122 (O_122,N_14830,N_14925);
or UO_123 (O_123,N_14955,N_14978);
or UO_124 (O_124,N_14980,N_14736);
nor UO_125 (O_125,N_14843,N_14798);
nor UO_126 (O_126,N_14786,N_14851);
xor UO_127 (O_127,N_14932,N_14976);
and UO_128 (O_128,N_14969,N_14746);
nand UO_129 (O_129,N_14965,N_14734);
and UO_130 (O_130,N_14796,N_14908);
nor UO_131 (O_131,N_14792,N_14958);
nor UO_132 (O_132,N_14992,N_14849);
nor UO_133 (O_133,N_14837,N_14738);
or UO_134 (O_134,N_14794,N_14845);
or UO_135 (O_135,N_14876,N_14818);
nand UO_136 (O_136,N_14847,N_14883);
nand UO_137 (O_137,N_14887,N_14942);
and UO_138 (O_138,N_14702,N_14921);
or UO_139 (O_139,N_14868,N_14807);
xnor UO_140 (O_140,N_14770,N_14751);
or UO_141 (O_141,N_14919,N_14827);
xnor UO_142 (O_142,N_14735,N_14744);
and UO_143 (O_143,N_14725,N_14760);
and UO_144 (O_144,N_14778,N_14815);
and UO_145 (O_145,N_14931,N_14882);
or UO_146 (O_146,N_14971,N_14884);
nor UO_147 (O_147,N_14927,N_14739);
and UO_148 (O_148,N_14880,N_14923);
xnor UO_149 (O_149,N_14941,N_14788);
or UO_150 (O_150,N_14763,N_14931);
nand UO_151 (O_151,N_14708,N_14911);
and UO_152 (O_152,N_14935,N_14873);
nand UO_153 (O_153,N_14757,N_14885);
and UO_154 (O_154,N_14820,N_14700);
or UO_155 (O_155,N_14964,N_14827);
xnor UO_156 (O_156,N_14830,N_14952);
and UO_157 (O_157,N_14718,N_14770);
or UO_158 (O_158,N_14900,N_14748);
xnor UO_159 (O_159,N_14985,N_14754);
nand UO_160 (O_160,N_14966,N_14896);
and UO_161 (O_161,N_14787,N_14768);
xor UO_162 (O_162,N_14715,N_14840);
or UO_163 (O_163,N_14918,N_14980);
nor UO_164 (O_164,N_14936,N_14821);
nand UO_165 (O_165,N_14947,N_14891);
xor UO_166 (O_166,N_14743,N_14937);
nor UO_167 (O_167,N_14895,N_14835);
and UO_168 (O_168,N_14929,N_14889);
and UO_169 (O_169,N_14792,N_14732);
nor UO_170 (O_170,N_14910,N_14751);
and UO_171 (O_171,N_14876,N_14728);
xor UO_172 (O_172,N_14874,N_14888);
xnor UO_173 (O_173,N_14774,N_14891);
and UO_174 (O_174,N_14911,N_14724);
and UO_175 (O_175,N_14848,N_14958);
nor UO_176 (O_176,N_14935,N_14951);
nor UO_177 (O_177,N_14775,N_14909);
xnor UO_178 (O_178,N_14917,N_14846);
xnor UO_179 (O_179,N_14979,N_14717);
and UO_180 (O_180,N_14870,N_14864);
xor UO_181 (O_181,N_14875,N_14928);
nor UO_182 (O_182,N_14717,N_14895);
nand UO_183 (O_183,N_14763,N_14994);
or UO_184 (O_184,N_14770,N_14987);
nand UO_185 (O_185,N_14802,N_14966);
or UO_186 (O_186,N_14709,N_14788);
nor UO_187 (O_187,N_14972,N_14821);
nor UO_188 (O_188,N_14971,N_14860);
xnor UO_189 (O_189,N_14804,N_14783);
and UO_190 (O_190,N_14830,N_14953);
or UO_191 (O_191,N_14957,N_14869);
and UO_192 (O_192,N_14918,N_14788);
and UO_193 (O_193,N_14943,N_14845);
xnor UO_194 (O_194,N_14773,N_14893);
nand UO_195 (O_195,N_14940,N_14886);
and UO_196 (O_196,N_14832,N_14984);
or UO_197 (O_197,N_14722,N_14952);
xnor UO_198 (O_198,N_14885,N_14930);
xor UO_199 (O_199,N_14796,N_14911);
or UO_200 (O_200,N_14727,N_14981);
xnor UO_201 (O_201,N_14741,N_14922);
and UO_202 (O_202,N_14882,N_14974);
or UO_203 (O_203,N_14949,N_14879);
or UO_204 (O_204,N_14736,N_14838);
or UO_205 (O_205,N_14746,N_14976);
and UO_206 (O_206,N_14836,N_14776);
or UO_207 (O_207,N_14835,N_14725);
nor UO_208 (O_208,N_14730,N_14822);
nand UO_209 (O_209,N_14774,N_14840);
xor UO_210 (O_210,N_14912,N_14907);
or UO_211 (O_211,N_14884,N_14734);
and UO_212 (O_212,N_14897,N_14715);
and UO_213 (O_213,N_14865,N_14956);
nand UO_214 (O_214,N_14962,N_14876);
and UO_215 (O_215,N_14809,N_14931);
and UO_216 (O_216,N_14956,N_14704);
and UO_217 (O_217,N_14775,N_14821);
or UO_218 (O_218,N_14964,N_14993);
xnor UO_219 (O_219,N_14848,N_14788);
and UO_220 (O_220,N_14847,N_14951);
nor UO_221 (O_221,N_14825,N_14864);
nor UO_222 (O_222,N_14864,N_14952);
xnor UO_223 (O_223,N_14812,N_14983);
nand UO_224 (O_224,N_14923,N_14872);
nor UO_225 (O_225,N_14948,N_14782);
or UO_226 (O_226,N_14861,N_14762);
nor UO_227 (O_227,N_14873,N_14754);
nor UO_228 (O_228,N_14717,N_14936);
and UO_229 (O_229,N_14723,N_14825);
nand UO_230 (O_230,N_14761,N_14912);
xnor UO_231 (O_231,N_14888,N_14901);
nand UO_232 (O_232,N_14976,N_14856);
xor UO_233 (O_233,N_14903,N_14785);
nand UO_234 (O_234,N_14868,N_14878);
nand UO_235 (O_235,N_14836,N_14909);
xor UO_236 (O_236,N_14852,N_14749);
nor UO_237 (O_237,N_14841,N_14983);
nand UO_238 (O_238,N_14705,N_14983);
and UO_239 (O_239,N_14875,N_14776);
or UO_240 (O_240,N_14988,N_14835);
and UO_241 (O_241,N_14847,N_14773);
nor UO_242 (O_242,N_14814,N_14822);
nor UO_243 (O_243,N_14890,N_14960);
or UO_244 (O_244,N_14973,N_14950);
xor UO_245 (O_245,N_14756,N_14707);
xnor UO_246 (O_246,N_14815,N_14728);
or UO_247 (O_247,N_14896,N_14942);
nor UO_248 (O_248,N_14843,N_14945);
xor UO_249 (O_249,N_14900,N_14747);
and UO_250 (O_250,N_14744,N_14962);
xor UO_251 (O_251,N_14761,N_14720);
nor UO_252 (O_252,N_14947,N_14791);
nor UO_253 (O_253,N_14954,N_14793);
xor UO_254 (O_254,N_14967,N_14971);
xnor UO_255 (O_255,N_14882,N_14958);
and UO_256 (O_256,N_14949,N_14814);
nand UO_257 (O_257,N_14983,N_14984);
or UO_258 (O_258,N_14828,N_14919);
and UO_259 (O_259,N_14908,N_14963);
xnor UO_260 (O_260,N_14821,N_14878);
and UO_261 (O_261,N_14897,N_14928);
xor UO_262 (O_262,N_14950,N_14930);
and UO_263 (O_263,N_14834,N_14826);
and UO_264 (O_264,N_14971,N_14886);
and UO_265 (O_265,N_14771,N_14700);
and UO_266 (O_266,N_14861,N_14998);
xor UO_267 (O_267,N_14866,N_14797);
xnor UO_268 (O_268,N_14855,N_14889);
nand UO_269 (O_269,N_14700,N_14967);
nand UO_270 (O_270,N_14941,N_14759);
nand UO_271 (O_271,N_14936,N_14902);
nor UO_272 (O_272,N_14705,N_14954);
or UO_273 (O_273,N_14933,N_14826);
nand UO_274 (O_274,N_14892,N_14842);
nand UO_275 (O_275,N_14768,N_14858);
xnor UO_276 (O_276,N_14761,N_14777);
nor UO_277 (O_277,N_14896,N_14981);
nand UO_278 (O_278,N_14795,N_14860);
xnor UO_279 (O_279,N_14830,N_14995);
or UO_280 (O_280,N_14895,N_14707);
nor UO_281 (O_281,N_14896,N_14843);
nor UO_282 (O_282,N_14716,N_14724);
nor UO_283 (O_283,N_14964,N_14782);
or UO_284 (O_284,N_14700,N_14742);
xor UO_285 (O_285,N_14788,N_14865);
nor UO_286 (O_286,N_14980,N_14896);
or UO_287 (O_287,N_14927,N_14827);
nor UO_288 (O_288,N_14890,N_14790);
nor UO_289 (O_289,N_14981,N_14831);
and UO_290 (O_290,N_14935,N_14784);
nor UO_291 (O_291,N_14993,N_14973);
nand UO_292 (O_292,N_14936,N_14755);
nor UO_293 (O_293,N_14780,N_14954);
and UO_294 (O_294,N_14758,N_14916);
nand UO_295 (O_295,N_14925,N_14964);
or UO_296 (O_296,N_14821,N_14977);
or UO_297 (O_297,N_14821,N_14843);
and UO_298 (O_298,N_14731,N_14801);
nand UO_299 (O_299,N_14990,N_14834);
xor UO_300 (O_300,N_14908,N_14825);
nor UO_301 (O_301,N_14961,N_14777);
and UO_302 (O_302,N_14719,N_14887);
or UO_303 (O_303,N_14879,N_14750);
nand UO_304 (O_304,N_14756,N_14866);
nand UO_305 (O_305,N_14997,N_14981);
nand UO_306 (O_306,N_14917,N_14778);
nor UO_307 (O_307,N_14701,N_14801);
nand UO_308 (O_308,N_14962,N_14701);
nand UO_309 (O_309,N_14702,N_14721);
or UO_310 (O_310,N_14975,N_14778);
and UO_311 (O_311,N_14812,N_14737);
xnor UO_312 (O_312,N_14755,N_14700);
and UO_313 (O_313,N_14832,N_14953);
or UO_314 (O_314,N_14915,N_14763);
nor UO_315 (O_315,N_14826,N_14845);
nand UO_316 (O_316,N_14703,N_14838);
xor UO_317 (O_317,N_14715,N_14776);
xnor UO_318 (O_318,N_14989,N_14959);
nand UO_319 (O_319,N_14911,N_14773);
nand UO_320 (O_320,N_14819,N_14702);
or UO_321 (O_321,N_14964,N_14842);
and UO_322 (O_322,N_14781,N_14714);
xor UO_323 (O_323,N_14714,N_14996);
nor UO_324 (O_324,N_14844,N_14918);
nor UO_325 (O_325,N_14849,N_14889);
and UO_326 (O_326,N_14988,N_14785);
or UO_327 (O_327,N_14700,N_14808);
xor UO_328 (O_328,N_14735,N_14994);
and UO_329 (O_329,N_14899,N_14857);
or UO_330 (O_330,N_14755,N_14719);
xnor UO_331 (O_331,N_14727,N_14778);
or UO_332 (O_332,N_14750,N_14793);
or UO_333 (O_333,N_14789,N_14810);
or UO_334 (O_334,N_14933,N_14986);
nand UO_335 (O_335,N_14711,N_14702);
xnor UO_336 (O_336,N_14943,N_14731);
xor UO_337 (O_337,N_14704,N_14780);
xnor UO_338 (O_338,N_14705,N_14821);
nor UO_339 (O_339,N_14884,N_14759);
xnor UO_340 (O_340,N_14739,N_14817);
or UO_341 (O_341,N_14782,N_14992);
and UO_342 (O_342,N_14991,N_14787);
nor UO_343 (O_343,N_14956,N_14757);
nand UO_344 (O_344,N_14923,N_14778);
xnor UO_345 (O_345,N_14955,N_14808);
xor UO_346 (O_346,N_14970,N_14703);
nor UO_347 (O_347,N_14859,N_14970);
xnor UO_348 (O_348,N_14848,N_14965);
nor UO_349 (O_349,N_14884,N_14924);
nand UO_350 (O_350,N_14910,N_14813);
nand UO_351 (O_351,N_14722,N_14898);
xnor UO_352 (O_352,N_14850,N_14745);
nor UO_353 (O_353,N_14930,N_14957);
nor UO_354 (O_354,N_14831,N_14833);
xnor UO_355 (O_355,N_14788,N_14955);
nand UO_356 (O_356,N_14966,N_14926);
nor UO_357 (O_357,N_14882,N_14985);
nor UO_358 (O_358,N_14877,N_14856);
and UO_359 (O_359,N_14705,N_14892);
nand UO_360 (O_360,N_14861,N_14718);
and UO_361 (O_361,N_14987,N_14813);
nor UO_362 (O_362,N_14988,N_14805);
and UO_363 (O_363,N_14725,N_14832);
and UO_364 (O_364,N_14962,N_14982);
nand UO_365 (O_365,N_14921,N_14780);
nand UO_366 (O_366,N_14837,N_14925);
or UO_367 (O_367,N_14799,N_14825);
nand UO_368 (O_368,N_14769,N_14992);
nand UO_369 (O_369,N_14917,N_14795);
or UO_370 (O_370,N_14708,N_14927);
xor UO_371 (O_371,N_14910,N_14860);
and UO_372 (O_372,N_14832,N_14751);
xnor UO_373 (O_373,N_14908,N_14992);
nor UO_374 (O_374,N_14959,N_14919);
nand UO_375 (O_375,N_14894,N_14969);
nor UO_376 (O_376,N_14996,N_14961);
nand UO_377 (O_377,N_14901,N_14715);
xnor UO_378 (O_378,N_14888,N_14961);
and UO_379 (O_379,N_14900,N_14752);
xor UO_380 (O_380,N_14834,N_14714);
or UO_381 (O_381,N_14886,N_14873);
xor UO_382 (O_382,N_14743,N_14725);
and UO_383 (O_383,N_14728,N_14913);
nor UO_384 (O_384,N_14949,N_14735);
nor UO_385 (O_385,N_14934,N_14700);
and UO_386 (O_386,N_14759,N_14835);
and UO_387 (O_387,N_14829,N_14849);
xnor UO_388 (O_388,N_14838,N_14868);
nor UO_389 (O_389,N_14856,N_14907);
and UO_390 (O_390,N_14812,N_14745);
xnor UO_391 (O_391,N_14800,N_14867);
xor UO_392 (O_392,N_14758,N_14786);
and UO_393 (O_393,N_14941,N_14981);
and UO_394 (O_394,N_14855,N_14777);
nand UO_395 (O_395,N_14774,N_14719);
and UO_396 (O_396,N_14901,N_14777);
nand UO_397 (O_397,N_14867,N_14892);
and UO_398 (O_398,N_14826,N_14897);
xor UO_399 (O_399,N_14970,N_14940);
and UO_400 (O_400,N_14872,N_14851);
nor UO_401 (O_401,N_14750,N_14902);
or UO_402 (O_402,N_14994,N_14732);
nor UO_403 (O_403,N_14760,N_14998);
nor UO_404 (O_404,N_14757,N_14987);
nor UO_405 (O_405,N_14894,N_14796);
or UO_406 (O_406,N_14960,N_14962);
xnor UO_407 (O_407,N_14864,N_14905);
nand UO_408 (O_408,N_14858,N_14876);
nand UO_409 (O_409,N_14886,N_14956);
or UO_410 (O_410,N_14746,N_14701);
and UO_411 (O_411,N_14965,N_14808);
and UO_412 (O_412,N_14914,N_14736);
and UO_413 (O_413,N_14730,N_14832);
or UO_414 (O_414,N_14897,N_14831);
nor UO_415 (O_415,N_14945,N_14774);
nor UO_416 (O_416,N_14933,N_14701);
nand UO_417 (O_417,N_14955,N_14975);
nor UO_418 (O_418,N_14750,N_14727);
nand UO_419 (O_419,N_14780,N_14952);
and UO_420 (O_420,N_14836,N_14961);
nand UO_421 (O_421,N_14979,N_14756);
nand UO_422 (O_422,N_14973,N_14775);
and UO_423 (O_423,N_14829,N_14755);
xor UO_424 (O_424,N_14954,N_14911);
nand UO_425 (O_425,N_14907,N_14987);
nand UO_426 (O_426,N_14773,N_14876);
nor UO_427 (O_427,N_14973,N_14936);
nand UO_428 (O_428,N_14909,N_14925);
and UO_429 (O_429,N_14757,N_14745);
xor UO_430 (O_430,N_14931,N_14912);
nand UO_431 (O_431,N_14941,N_14921);
and UO_432 (O_432,N_14855,N_14839);
xnor UO_433 (O_433,N_14824,N_14725);
nor UO_434 (O_434,N_14744,N_14831);
nor UO_435 (O_435,N_14982,N_14759);
and UO_436 (O_436,N_14821,N_14875);
or UO_437 (O_437,N_14819,N_14869);
or UO_438 (O_438,N_14899,N_14737);
nand UO_439 (O_439,N_14706,N_14990);
and UO_440 (O_440,N_14794,N_14829);
and UO_441 (O_441,N_14877,N_14746);
or UO_442 (O_442,N_14869,N_14863);
or UO_443 (O_443,N_14830,N_14824);
or UO_444 (O_444,N_14874,N_14839);
or UO_445 (O_445,N_14923,N_14903);
and UO_446 (O_446,N_14736,N_14889);
nor UO_447 (O_447,N_14981,N_14915);
xor UO_448 (O_448,N_14994,N_14805);
nor UO_449 (O_449,N_14883,N_14845);
and UO_450 (O_450,N_14720,N_14881);
nor UO_451 (O_451,N_14757,N_14710);
xnor UO_452 (O_452,N_14949,N_14795);
or UO_453 (O_453,N_14746,N_14801);
nand UO_454 (O_454,N_14806,N_14810);
or UO_455 (O_455,N_14784,N_14787);
and UO_456 (O_456,N_14726,N_14973);
nor UO_457 (O_457,N_14958,N_14954);
nand UO_458 (O_458,N_14919,N_14703);
and UO_459 (O_459,N_14898,N_14979);
nor UO_460 (O_460,N_14862,N_14780);
nor UO_461 (O_461,N_14775,N_14947);
nor UO_462 (O_462,N_14985,N_14797);
xnor UO_463 (O_463,N_14844,N_14744);
xor UO_464 (O_464,N_14723,N_14949);
nor UO_465 (O_465,N_14969,N_14895);
xor UO_466 (O_466,N_14715,N_14727);
nor UO_467 (O_467,N_14947,N_14865);
or UO_468 (O_468,N_14801,N_14725);
nand UO_469 (O_469,N_14876,N_14826);
nor UO_470 (O_470,N_14975,N_14719);
nand UO_471 (O_471,N_14778,N_14999);
nor UO_472 (O_472,N_14980,N_14838);
or UO_473 (O_473,N_14707,N_14768);
or UO_474 (O_474,N_14808,N_14999);
xnor UO_475 (O_475,N_14959,N_14862);
nand UO_476 (O_476,N_14908,N_14971);
or UO_477 (O_477,N_14798,N_14719);
nand UO_478 (O_478,N_14736,N_14709);
nor UO_479 (O_479,N_14704,N_14725);
and UO_480 (O_480,N_14821,N_14757);
and UO_481 (O_481,N_14775,N_14774);
nand UO_482 (O_482,N_14928,N_14822);
or UO_483 (O_483,N_14843,N_14909);
xnor UO_484 (O_484,N_14754,N_14751);
or UO_485 (O_485,N_14887,N_14999);
nand UO_486 (O_486,N_14887,N_14701);
or UO_487 (O_487,N_14820,N_14866);
and UO_488 (O_488,N_14955,N_14921);
and UO_489 (O_489,N_14836,N_14886);
and UO_490 (O_490,N_14887,N_14789);
or UO_491 (O_491,N_14802,N_14830);
nor UO_492 (O_492,N_14788,N_14964);
xor UO_493 (O_493,N_14782,N_14773);
nand UO_494 (O_494,N_14981,N_14776);
or UO_495 (O_495,N_14759,N_14747);
nor UO_496 (O_496,N_14708,N_14945);
xnor UO_497 (O_497,N_14772,N_14736);
nand UO_498 (O_498,N_14860,N_14993);
xor UO_499 (O_499,N_14973,N_14758);
or UO_500 (O_500,N_14985,N_14892);
and UO_501 (O_501,N_14869,N_14968);
nand UO_502 (O_502,N_14758,N_14974);
xnor UO_503 (O_503,N_14823,N_14931);
or UO_504 (O_504,N_14726,N_14976);
xor UO_505 (O_505,N_14830,N_14823);
nor UO_506 (O_506,N_14771,N_14848);
nand UO_507 (O_507,N_14917,N_14872);
nor UO_508 (O_508,N_14974,N_14768);
nor UO_509 (O_509,N_14857,N_14754);
nand UO_510 (O_510,N_14909,N_14963);
xor UO_511 (O_511,N_14741,N_14983);
nor UO_512 (O_512,N_14724,N_14887);
or UO_513 (O_513,N_14750,N_14895);
nor UO_514 (O_514,N_14944,N_14703);
and UO_515 (O_515,N_14781,N_14893);
xnor UO_516 (O_516,N_14982,N_14923);
and UO_517 (O_517,N_14830,N_14731);
nand UO_518 (O_518,N_14778,N_14837);
nor UO_519 (O_519,N_14926,N_14778);
nand UO_520 (O_520,N_14733,N_14983);
nand UO_521 (O_521,N_14753,N_14841);
or UO_522 (O_522,N_14883,N_14800);
nor UO_523 (O_523,N_14921,N_14881);
xor UO_524 (O_524,N_14785,N_14802);
nor UO_525 (O_525,N_14762,N_14778);
nor UO_526 (O_526,N_14968,N_14961);
or UO_527 (O_527,N_14751,N_14983);
xor UO_528 (O_528,N_14972,N_14728);
nor UO_529 (O_529,N_14937,N_14863);
nor UO_530 (O_530,N_14831,N_14753);
nand UO_531 (O_531,N_14880,N_14911);
nand UO_532 (O_532,N_14743,N_14932);
or UO_533 (O_533,N_14915,N_14943);
or UO_534 (O_534,N_14851,N_14815);
nor UO_535 (O_535,N_14824,N_14878);
and UO_536 (O_536,N_14914,N_14897);
and UO_537 (O_537,N_14803,N_14865);
xor UO_538 (O_538,N_14937,N_14988);
nor UO_539 (O_539,N_14894,N_14739);
xnor UO_540 (O_540,N_14930,N_14804);
or UO_541 (O_541,N_14995,N_14706);
and UO_542 (O_542,N_14960,N_14947);
or UO_543 (O_543,N_14776,N_14869);
or UO_544 (O_544,N_14824,N_14937);
or UO_545 (O_545,N_14965,N_14833);
xor UO_546 (O_546,N_14833,N_14853);
or UO_547 (O_547,N_14875,N_14925);
nor UO_548 (O_548,N_14885,N_14855);
and UO_549 (O_549,N_14810,N_14770);
or UO_550 (O_550,N_14885,N_14839);
and UO_551 (O_551,N_14787,N_14945);
nor UO_552 (O_552,N_14800,N_14757);
or UO_553 (O_553,N_14906,N_14920);
xnor UO_554 (O_554,N_14772,N_14799);
and UO_555 (O_555,N_14995,N_14880);
nor UO_556 (O_556,N_14937,N_14729);
nand UO_557 (O_557,N_14879,N_14761);
and UO_558 (O_558,N_14861,N_14818);
or UO_559 (O_559,N_14972,N_14703);
nand UO_560 (O_560,N_14969,N_14815);
xnor UO_561 (O_561,N_14853,N_14871);
or UO_562 (O_562,N_14893,N_14825);
nand UO_563 (O_563,N_14936,N_14907);
xnor UO_564 (O_564,N_14861,N_14830);
and UO_565 (O_565,N_14968,N_14802);
or UO_566 (O_566,N_14842,N_14969);
nand UO_567 (O_567,N_14849,N_14938);
xnor UO_568 (O_568,N_14923,N_14893);
xnor UO_569 (O_569,N_14946,N_14901);
or UO_570 (O_570,N_14900,N_14885);
nor UO_571 (O_571,N_14853,N_14794);
xnor UO_572 (O_572,N_14926,N_14956);
nor UO_573 (O_573,N_14729,N_14751);
nor UO_574 (O_574,N_14948,N_14881);
xnor UO_575 (O_575,N_14797,N_14720);
or UO_576 (O_576,N_14788,N_14902);
nand UO_577 (O_577,N_14797,N_14913);
nand UO_578 (O_578,N_14790,N_14787);
or UO_579 (O_579,N_14874,N_14814);
nor UO_580 (O_580,N_14705,N_14995);
or UO_581 (O_581,N_14953,N_14759);
xor UO_582 (O_582,N_14919,N_14776);
xnor UO_583 (O_583,N_14934,N_14939);
nor UO_584 (O_584,N_14763,N_14950);
and UO_585 (O_585,N_14815,N_14722);
xnor UO_586 (O_586,N_14839,N_14947);
and UO_587 (O_587,N_14819,N_14709);
and UO_588 (O_588,N_14806,N_14998);
and UO_589 (O_589,N_14734,N_14805);
or UO_590 (O_590,N_14775,N_14817);
nor UO_591 (O_591,N_14859,N_14984);
or UO_592 (O_592,N_14713,N_14770);
nor UO_593 (O_593,N_14956,N_14842);
nor UO_594 (O_594,N_14801,N_14855);
nand UO_595 (O_595,N_14710,N_14713);
or UO_596 (O_596,N_14862,N_14982);
or UO_597 (O_597,N_14749,N_14949);
and UO_598 (O_598,N_14820,N_14875);
and UO_599 (O_599,N_14785,N_14823);
and UO_600 (O_600,N_14931,N_14841);
nand UO_601 (O_601,N_14993,N_14992);
xor UO_602 (O_602,N_14804,N_14752);
and UO_603 (O_603,N_14997,N_14859);
nor UO_604 (O_604,N_14923,N_14760);
or UO_605 (O_605,N_14937,N_14944);
nand UO_606 (O_606,N_14825,N_14986);
and UO_607 (O_607,N_14856,N_14851);
and UO_608 (O_608,N_14767,N_14737);
or UO_609 (O_609,N_14817,N_14937);
nor UO_610 (O_610,N_14831,N_14759);
nor UO_611 (O_611,N_14947,N_14824);
nand UO_612 (O_612,N_14727,N_14959);
or UO_613 (O_613,N_14846,N_14791);
nand UO_614 (O_614,N_14805,N_14725);
nand UO_615 (O_615,N_14890,N_14899);
and UO_616 (O_616,N_14999,N_14986);
xor UO_617 (O_617,N_14995,N_14869);
nand UO_618 (O_618,N_14764,N_14811);
nor UO_619 (O_619,N_14764,N_14860);
nand UO_620 (O_620,N_14912,N_14808);
or UO_621 (O_621,N_14708,N_14857);
and UO_622 (O_622,N_14702,N_14844);
and UO_623 (O_623,N_14832,N_14910);
and UO_624 (O_624,N_14707,N_14776);
or UO_625 (O_625,N_14861,N_14739);
nand UO_626 (O_626,N_14884,N_14732);
xnor UO_627 (O_627,N_14727,N_14900);
and UO_628 (O_628,N_14841,N_14849);
xor UO_629 (O_629,N_14868,N_14893);
nand UO_630 (O_630,N_14879,N_14956);
xor UO_631 (O_631,N_14849,N_14798);
nand UO_632 (O_632,N_14744,N_14993);
nor UO_633 (O_633,N_14874,N_14923);
and UO_634 (O_634,N_14718,N_14865);
xor UO_635 (O_635,N_14770,N_14771);
or UO_636 (O_636,N_14923,N_14921);
or UO_637 (O_637,N_14983,N_14814);
or UO_638 (O_638,N_14905,N_14904);
xnor UO_639 (O_639,N_14847,N_14764);
or UO_640 (O_640,N_14995,N_14862);
and UO_641 (O_641,N_14891,N_14710);
xor UO_642 (O_642,N_14887,N_14807);
nor UO_643 (O_643,N_14826,N_14881);
xor UO_644 (O_644,N_14890,N_14968);
and UO_645 (O_645,N_14915,N_14920);
or UO_646 (O_646,N_14965,N_14781);
xnor UO_647 (O_647,N_14722,N_14865);
xnor UO_648 (O_648,N_14722,N_14910);
nand UO_649 (O_649,N_14791,N_14882);
or UO_650 (O_650,N_14721,N_14729);
nor UO_651 (O_651,N_14700,N_14781);
xor UO_652 (O_652,N_14759,N_14958);
nand UO_653 (O_653,N_14741,N_14723);
or UO_654 (O_654,N_14950,N_14924);
and UO_655 (O_655,N_14919,N_14864);
nor UO_656 (O_656,N_14724,N_14806);
nor UO_657 (O_657,N_14947,N_14782);
or UO_658 (O_658,N_14990,N_14865);
xnor UO_659 (O_659,N_14993,N_14745);
nor UO_660 (O_660,N_14762,N_14878);
nor UO_661 (O_661,N_14840,N_14754);
and UO_662 (O_662,N_14929,N_14762);
nor UO_663 (O_663,N_14878,N_14944);
nand UO_664 (O_664,N_14729,N_14926);
nand UO_665 (O_665,N_14990,N_14928);
nor UO_666 (O_666,N_14712,N_14724);
nor UO_667 (O_667,N_14718,N_14725);
and UO_668 (O_668,N_14836,N_14854);
and UO_669 (O_669,N_14954,N_14717);
or UO_670 (O_670,N_14808,N_14759);
nor UO_671 (O_671,N_14850,N_14826);
nand UO_672 (O_672,N_14768,N_14747);
nand UO_673 (O_673,N_14844,N_14709);
or UO_674 (O_674,N_14877,N_14816);
xnor UO_675 (O_675,N_14893,N_14753);
nor UO_676 (O_676,N_14952,N_14837);
or UO_677 (O_677,N_14835,N_14855);
nand UO_678 (O_678,N_14781,N_14935);
nor UO_679 (O_679,N_14850,N_14945);
and UO_680 (O_680,N_14870,N_14916);
or UO_681 (O_681,N_14896,N_14726);
nor UO_682 (O_682,N_14794,N_14935);
nor UO_683 (O_683,N_14727,N_14728);
xor UO_684 (O_684,N_14983,N_14771);
nand UO_685 (O_685,N_14809,N_14733);
nor UO_686 (O_686,N_14711,N_14842);
nor UO_687 (O_687,N_14990,N_14750);
nand UO_688 (O_688,N_14901,N_14862);
xnor UO_689 (O_689,N_14907,N_14798);
xor UO_690 (O_690,N_14865,N_14721);
xor UO_691 (O_691,N_14765,N_14729);
xnor UO_692 (O_692,N_14993,N_14869);
nand UO_693 (O_693,N_14748,N_14778);
and UO_694 (O_694,N_14797,N_14719);
or UO_695 (O_695,N_14997,N_14830);
or UO_696 (O_696,N_14965,N_14716);
or UO_697 (O_697,N_14912,N_14975);
nor UO_698 (O_698,N_14851,N_14738);
nand UO_699 (O_699,N_14977,N_14743);
nand UO_700 (O_700,N_14903,N_14761);
nor UO_701 (O_701,N_14941,N_14911);
nor UO_702 (O_702,N_14849,N_14900);
xor UO_703 (O_703,N_14832,N_14937);
and UO_704 (O_704,N_14808,N_14799);
or UO_705 (O_705,N_14707,N_14736);
xor UO_706 (O_706,N_14952,N_14703);
xnor UO_707 (O_707,N_14904,N_14854);
nor UO_708 (O_708,N_14929,N_14868);
nand UO_709 (O_709,N_14835,N_14958);
or UO_710 (O_710,N_14990,N_14896);
xor UO_711 (O_711,N_14873,N_14766);
nor UO_712 (O_712,N_14744,N_14752);
and UO_713 (O_713,N_14976,N_14804);
or UO_714 (O_714,N_14865,N_14972);
nand UO_715 (O_715,N_14959,N_14907);
xor UO_716 (O_716,N_14909,N_14917);
nor UO_717 (O_717,N_14891,N_14979);
nand UO_718 (O_718,N_14929,N_14773);
or UO_719 (O_719,N_14919,N_14820);
or UO_720 (O_720,N_14842,N_14907);
nor UO_721 (O_721,N_14832,N_14911);
and UO_722 (O_722,N_14799,N_14967);
and UO_723 (O_723,N_14880,N_14820);
nor UO_724 (O_724,N_14978,N_14876);
nand UO_725 (O_725,N_14896,N_14935);
and UO_726 (O_726,N_14761,N_14955);
nand UO_727 (O_727,N_14718,N_14788);
nor UO_728 (O_728,N_14849,N_14974);
nor UO_729 (O_729,N_14742,N_14835);
and UO_730 (O_730,N_14754,N_14735);
nor UO_731 (O_731,N_14991,N_14830);
xnor UO_732 (O_732,N_14995,N_14823);
or UO_733 (O_733,N_14846,N_14886);
or UO_734 (O_734,N_14860,N_14768);
nand UO_735 (O_735,N_14942,N_14945);
nor UO_736 (O_736,N_14795,N_14957);
and UO_737 (O_737,N_14935,N_14868);
xnor UO_738 (O_738,N_14824,N_14862);
or UO_739 (O_739,N_14855,N_14989);
or UO_740 (O_740,N_14960,N_14903);
or UO_741 (O_741,N_14912,N_14956);
and UO_742 (O_742,N_14786,N_14749);
or UO_743 (O_743,N_14925,N_14760);
nand UO_744 (O_744,N_14743,N_14957);
nand UO_745 (O_745,N_14944,N_14748);
nor UO_746 (O_746,N_14909,N_14914);
nand UO_747 (O_747,N_14812,N_14836);
nor UO_748 (O_748,N_14989,N_14934);
and UO_749 (O_749,N_14751,N_14711);
or UO_750 (O_750,N_14714,N_14757);
nor UO_751 (O_751,N_14821,N_14748);
nor UO_752 (O_752,N_14856,N_14755);
or UO_753 (O_753,N_14700,N_14734);
or UO_754 (O_754,N_14754,N_14894);
and UO_755 (O_755,N_14885,N_14978);
nand UO_756 (O_756,N_14845,N_14966);
and UO_757 (O_757,N_14861,N_14722);
nor UO_758 (O_758,N_14833,N_14947);
and UO_759 (O_759,N_14710,N_14726);
nor UO_760 (O_760,N_14919,N_14793);
and UO_761 (O_761,N_14850,N_14701);
and UO_762 (O_762,N_14790,N_14851);
nor UO_763 (O_763,N_14963,N_14906);
nand UO_764 (O_764,N_14980,N_14938);
nor UO_765 (O_765,N_14773,N_14836);
and UO_766 (O_766,N_14733,N_14797);
nand UO_767 (O_767,N_14960,N_14764);
and UO_768 (O_768,N_14899,N_14738);
xor UO_769 (O_769,N_14899,N_14741);
nand UO_770 (O_770,N_14743,N_14701);
nand UO_771 (O_771,N_14762,N_14828);
or UO_772 (O_772,N_14968,N_14709);
nand UO_773 (O_773,N_14889,N_14735);
xor UO_774 (O_774,N_14934,N_14709);
and UO_775 (O_775,N_14874,N_14945);
nor UO_776 (O_776,N_14778,N_14700);
nor UO_777 (O_777,N_14735,N_14797);
xnor UO_778 (O_778,N_14733,N_14978);
xor UO_779 (O_779,N_14910,N_14715);
nor UO_780 (O_780,N_14821,N_14869);
and UO_781 (O_781,N_14867,N_14886);
nor UO_782 (O_782,N_14763,N_14940);
or UO_783 (O_783,N_14924,N_14939);
nand UO_784 (O_784,N_14821,N_14947);
nand UO_785 (O_785,N_14871,N_14840);
nand UO_786 (O_786,N_14717,N_14767);
nand UO_787 (O_787,N_14948,N_14898);
nand UO_788 (O_788,N_14722,N_14805);
nor UO_789 (O_789,N_14734,N_14825);
nor UO_790 (O_790,N_14862,N_14867);
nand UO_791 (O_791,N_14853,N_14957);
or UO_792 (O_792,N_14842,N_14808);
nor UO_793 (O_793,N_14860,N_14893);
xor UO_794 (O_794,N_14716,N_14915);
and UO_795 (O_795,N_14959,N_14723);
xor UO_796 (O_796,N_14836,N_14726);
or UO_797 (O_797,N_14730,N_14954);
or UO_798 (O_798,N_14722,N_14866);
xor UO_799 (O_799,N_14760,N_14917);
xnor UO_800 (O_800,N_14950,N_14905);
nand UO_801 (O_801,N_14719,N_14806);
xor UO_802 (O_802,N_14912,N_14768);
xor UO_803 (O_803,N_14943,N_14937);
or UO_804 (O_804,N_14807,N_14700);
nor UO_805 (O_805,N_14778,N_14868);
nor UO_806 (O_806,N_14790,N_14863);
or UO_807 (O_807,N_14838,N_14852);
xnor UO_808 (O_808,N_14720,N_14728);
xor UO_809 (O_809,N_14963,N_14802);
or UO_810 (O_810,N_14968,N_14863);
nor UO_811 (O_811,N_14925,N_14746);
and UO_812 (O_812,N_14922,N_14866);
nor UO_813 (O_813,N_14714,N_14823);
nand UO_814 (O_814,N_14911,N_14978);
and UO_815 (O_815,N_14888,N_14995);
nor UO_816 (O_816,N_14947,N_14743);
xnor UO_817 (O_817,N_14840,N_14848);
or UO_818 (O_818,N_14901,N_14863);
and UO_819 (O_819,N_14711,N_14866);
nor UO_820 (O_820,N_14946,N_14734);
xor UO_821 (O_821,N_14986,N_14755);
nand UO_822 (O_822,N_14951,N_14944);
xor UO_823 (O_823,N_14821,N_14717);
nor UO_824 (O_824,N_14848,N_14948);
nand UO_825 (O_825,N_14964,N_14838);
nand UO_826 (O_826,N_14986,N_14882);
nor UO_827 (O_827,N_14978,N_14743);
xnor UO_828 (O_828,N_14845,N_14850);
nor UO_829 (O_829,N_14733,N_14905);
xnor UO_830 (O_830,N_14938,N_14898);
nor UO_831 (O_831,N_14921,N_14997);
and UO_832 (O_832,N_14845,N_14861);
nand UO_833 (O_833,N_14802,N_14767);
or UO_834 (O_834,N_14817,N_14875);
nor UO_835 (O_835,N_14852,N_14842);
nor UO_836 (O_836,N_14859,N_14906);
nand UO_837 (O_837,N_14808,N_14911);
or UO_838 (O_838,N_14739,N_14837);
and UO_839 (O_839,N_14884,N_14861);
nand UO_840 (O_840,N_14928,N_14761);
xor UO_841 (O_841,N_14856,N_14770);
or UO_842 (O_842,N_14933,N_14831);
xor UO_843 (O_843,N_14717,N_14806);
nand UO_844 (O_844,N_14875,N_14968);
nor UO_845 (O_845,N_14968,N_14907);
or UO_846 (O_846,N_14866,N_14990);
nand UO_847 (O_847,N_14746,N_14807);
and UO_848 (O_848,N_14708,N_14811);
nor UO_849 (O_849,N_14808,N_14794);
nor UO_850 (O_850,N_14828,N_14795);
nand UO_851 (O_851,N_14886,N_14779);
nand UO_852 (O_852,N_14738,N_14864);
nor UO_853 (O_853,N_14939,N_14796);
nor UO_854 (O_854,N_14923,N_14985);
nand UO_855 (O_855,N_14781,N_14873);
or UO_856 (O_856,N_14851,N_14953);
nor UO_857 (O_857,N_14725,N_14850);
or UO_858 (O_858,N_14886,N_14843);
or UO_859 (O_859,N_14969,N_14739);
xor UO_860 (O_860,N_14943,N_14789);
or UO_861 (O_861,N_14843,N_14928);
or UO_862 (O_862,N_14895,N_14813);
or UO_863 (O_863,N_14815,N_14821);
or UO_864 (O_864,N_14706,N_14791);
and UO_865 (O_865,N_14701,N_14955);
and UO_866 (O_866,N_14881,N_14837);
xnor UO_867 (O_867,N_14726,N_14872);
nand UO_868 (O_868,N_14903,N_14891);
nor UO_869 (O_869,N_14729,N_14896);
or UO_870 (O_870,N_14914,N_14935);
xnor UO_871 (O_871,N_14782,N_14737);
and UO_872 (O_872,N_14974,N_14837);
nor UO_873 (O_873,N_14876,N_14775);
or UO_874 (O_874,N_14869,N_14762);
and UO_875 (O_875,N_14952,N_14950);
nor UO_876 (O_876,N_14724,N_14904);
xnor UO_877 (O_877,N_14728,N_14826);
nand UO_878 (O_878,N_14940,N_14718);
and UO_879 (O_879,N_14718,N_14798);
nand UO_880 (O_880,N_14830,N_14700);
nand UO_881 (O_881,N_14716,N_14700);
or UO_882 (O_882,N_14933,N_14849);
and UO_883 (O_883,N_14708,N_14787);
or UO_884 (O_884,N_14929,N_14977);
nor UO_885 (O_885,N_14805,N_14933);
or UO_886 (O_886,N_14877,N_14985);
nand UO_887 (O_887,N_14778,N_14722);
or UO_888 (O_888,N_14708,N_14756);
nor UO_889 (O_889,N_14822,N_14872);
and UO_890 (O_890,N_14799,N_14708);
nand UO_891 (O_891,N_14957,N_14955);
nand UO_892 (O_892,N_14889,N_14948);
nand UO_893 (O_893,N_14872,N_14818);
or UO_894 (O_894,N_14799,N_14721);
and UO_895 (O_895,N_14771,N_14800);
and UO_896 (O_896,N_14785,N_14726);
nand UO_897 (O_897,N_14938,N_14791);
nor UO_898 (O_898,N_14747,N_14714);
nor UO_899 (O_899,N_14981,N_14990);
and UO_900 (O_900,N_14996,N_14846);
xnor UO_901 (O_901,N_14785,N_14891);
nor UO_902 (O_902,N_14941,N_14818);
and UO_903 (O_903,N_14974,N_14897);
nand UO_904 (O_904,N_14936,N_14849);
or UO_905 (O_905,N_14810,N_14987);
or UO_906 (O_906,N_14746,N_14977);
or UO_907 (O_907,N_14723,N_14933);
xnor UO_908 (O_908,N_14977,N_14764);
and UO_909 (O_909,N_14806,N_14953);
and UO_910 (O_910,N_14727,N_14702);
nand UO_911 (O_911,N_14768,N_14720);
xnor UO_912 (O_912,N_14809,N_14846);
xnor UO_913 (O_913,N_14941,N_14861);
and UO_914 (O_914,N_14909,N_14947);
xnor UO_915 (O_915,N_14747,N_14775);
xnor UO_916 (O_916,N_14762,N_14884);
nand UO_917 (O_917,N_14990,N_14929);
and UO_918 (O_918,N_14862,N_14781);
nand UO_919 (O_919,N_14943,N_14990);
nor UO_920 (O_920,N_14958,N_14927);
nor UO_921 (O_921,N_14833,N_14823);
nand UO_922 (O_922,N_14797,N_14801);
nand UO_923 (O_923,N_14856,N_14940);
xor UO_924 (O_924,N_14858,N_14820);
nor UO_925 (O_925,N_14804,N_14753);
nand UO_926 (O_926,N_14756,N_14705);
nand UO_927 (O_927,N_14838,N_14793);
xor UO_928 (O_928,N_14876,N_14847);
xnor UO_929 (O_929,N_14715,N_14786);
or UO_930 (O_930,N_14865,N_14917);
and UO_931 (O_931,N_14972,N_14971);
and UO_932 (O_932,N_14897,N_14910);
nor UO_933 (O_933,N_14727,N_14817);
and UO_934 (O_934,N_14889,N_14863);
and UO_935 (O_935,N_14810,N_14970);
or UO_936 (O_936,N_14902,N_14930);
and UO_937 (O_937,N_14871,N_14753);
or UO_938 (O_938,N_14955,N_14900);
or UO_939 (O_939,N_14715,N_14935);
or UO_940 (O_940,N_14889,N_14866);
or UO_941 (O_941,N_14714,N_14884);
nor UO_942 (O_942,N_14714,N_14934);
and UO_943 (O_943,N_14794,N_14971);
nor UO_944 (O_944,N_14700,N_14818);
or UO_945 (O_945,N_14897,N_14759);
nor UO_946 (O_946,N_14703,N_14717);
xnor UO_947 (O_947,N_14764,N_14991);
and UO_948 (O_948,N_14913,N_14837);
or UO_949 (O_949,N_14894,N_14956);
nand UO_950 (O_950,N_14897,N_14885);
or UO_951 (O_951,N_14949,N_14927);
or UO_952 (O_952,N_14873,N_14787);
nand UO_953 (O_953,N_14960,N_14803);
nor UO_954 (O_954,N_14801,N_14936);
or UO_955 (O_955,N_14926,N_14950);
nor UO_956 (O_956,N_14954,N_14975);
nand UO_957 (O_957,N_14925,N_14932);
nand UO_958 (O_958,N_14740,N_14791);
xor UO_959 (O_959,N_14789,N_14858);
or UO_960 (O_960,N_14796,N_14714);
xor UO_961 (O_961,N_14814,N_14851);
xnor UO_962 (O_962,N_14726,N_14736);
and UO_963 (O_963,N_14746,N_14876);
and UO_964 (O_964,N_14908,N_14812);
or UO_965 (O_965,N_14955,N_14938);
xnor UO_966 (O_966,N_14831,N_14971);
nand UO_967 (O_967,N_14904,N_14831);
or UO_968 (O_968,N_14932,N_14999);
nand UO_969 (O_969,N_14879,N_14958);
or UO_970 (O_970,N_14750,N_14941);
and UO_971 (O_971,N_14701,N_14957);
nor UO_972 (O_972,N_14791,N_14767);
or UO_973 (O_973,N_14854,N_14857);
nand UO_974 (O_974,N_14986,N_14892);
or UO_975 (O_975,N_14839,N_14916);
nor UO_976 (O_976,N_14821,N_14795);
nor UO_977 (O_977,N_14716,N_14913);
nand UO_978 (O_978,N_14986,N_14941);
or UO_979 (O_979,N_14827,N_14826);
or UO_980 (O_980,N_14769,N_14947);
or UO_981 (O_981,N_14860,N_14857);
nor UO_982 (O_982,N_14728,N_14879);
nor UO_983 (O_983,N_14861,N_14970);
and UO_984 (O_984,N_14903,N_14893);
xnor UO_985 (O_985,N_14842,N_14874);
and UO_986 (O_986,N_14708,N_14823);
nand UO_987 (O_987,N_14928,N_14893);
nand UO_988 (O_988,N_14930,N_14734);
xnor UO_989 (O_989,N_14932,N_14990);
nor UO_990 (O_990,N_14768,N_14786);
xor UO_991 (O_991,N_14701,N_14869);
and UO_992 (O_992,N_14773,N_14912);
and UO_993 (O_993,N_14793,N_14990);
nor UO_994 (O_994,N_14746,N_14988);
and UO_995 (O_995,N_14806,N_14708);
xnor UO_996 (O_996,N_14776,N_14963);
xnor UO_997 (O_997,N_14785,N_14788);
and UO_998 (O_998,N_14854,N_14984);
nand UO_999 (O_999,N_14764,N_14897);
nor UO_1000 (O_1000,N_14825,N_14851);
xnor UO_1001 (O_1001,N_14723,N_14811);
xnor UO_1002 (O_1002,N_14765,N_14914);
and UO_1003 (O_1003,N_14938,N_14852);
and UO_1004 (O_1004,N_14989,N_14816);
and UO_1005 (O_1005,N_14999,N_14856);
or UO_1006 (O_1006,N_14981,N_14978);
xnor UO_1007 (O_1007,N_14837,N_14789);
nand UO_1008 (O_1008,N_14851,N_14842);
and UO_1009 (O_1009,N_14850,N_14790);
xnor UO_1010 (O_1010,N_14893,N_14981);
and UO_1011 (O_1011,N_14797,N_14878);
xnor UO_1012 (O_1012,N_14752,N_14976);
xnor UO_1013 (O_1013,N_14942,N_14831);
xor UO_1014 (O_1014,N_14967,N_14944);
nand UO_1015 (O_1015,N_14740,N_14836);
nand UO_1016 (O_1016,N_14976,N_14788);
and UO_1017 (O_1017,N_14716,N_14907);
nor UO_1018 (O_1018,N_14793,N_14810);
nand UO_1019 (O_1019,N_14911,N_14709);
and UO_1020 (O_1020,N_14985,N_14880);
or UO_1021 (O_1021,N_14794,N_14779);
xor UO_1022 (O_1022,N_14892,N_14724);
nand UO_1023 (O_1023,N_14917,N_14730);
xor UO_1024 (O_1024,N_14879,N_14771);
nor UO_1025 (O_1025,N_14728,N_14953);
and UO_1026 (O_1026,N_14739,N_14931);
nand UO_1027 (O_1027,N_14855,N_14829);
and UO_1028 (O_1028,N_14723,N_14908);
nor UO_1029 (O_1029,N_14742,N_14762);
and UO_1030 (O_1030,N_14976,N_14975);
nand UO_1031 (O_1031,N_14840,N_14975);
or UO_1032 (O_1032,N_14811,N_14905);
nor UO_1033 (O_1033,N_14882,N_14945);
and UO_1034 (O_1034,N_14873,N_14716);
xnor UO_1035 (O_1035,N_14877,N_14732);
and UO_1036 (O_1036,N_14865,N_14751);
and UO_1037 (O_1037,N_14879,N_14929);
nor UO_1038 (O_1038,N_14731,N_14814);
nand UO_1039 (O_1039,N_14703,N_14823);
nor UO_1040 (O_1040,N_14704,N_14758);
or UO_1041 (O_1041,N_14782,N_14859);
xnor UO_1042 (O_1042,N_14896,N_14758);
nor UO_1043 (O_1043,N_14758,N_14891);
xnor UO_1044 (O_1044,N_14900,N_14920);
nand UO_1045 (O_1045,N_14701,N_14728);
nor UO_1046 (O_1046,N_14905,N_14802);
xor UO_1047 (O_1047,N_14903,N_14984);
xnor UO_1048 (O_1048,N_14856,N_14837);
or UO_1049 (O_1049,N_14775,N_14713);
or UO_1050 (O_1050,N_14951,N_14807);
and UO_1051 (O_1051,N_14950,N_14846);
xnor UO_1052 (O_1052,N_14898,N_14802);
and UO_1053 (O_1053,N_14981,N_14878);
or UO_1054 (O_1054,N_14914,N_14807);
nor UO_1055 (O_1055,N_14904,N_14910);
nor UO_1056 (O_1056,N_14827,N_14872);
xor UO_1057 (O_1057,N_14973,N_14966);
or UO_1058 (O_1058,N_14996,N_14973);
and UO_1059 (O_1059,N_14915,N_14968);
and UO_1060 (O_1060,N_14832,N_14724);
and UO_1061 (O_1061,N_14995,N_14759);
or UO_1062 (O_1062,N_14912,N_14847);
nand UO_1063 (O_1063,N_14789,N_14781);
xnor UO_1064 (O_1064,N_14737,N_14833);
or UO_1065 (O_1065,N_14837,N_14728);
and UO_1066 (O_1066,N_14733,N_14730);
and UO_1067 (O_1067,N_14804,N_14733);
nand UO_1068 (O_1068,N_14737,N_14756);
nand UO_1069 (O_1069,N_14759,N_14936);
nand UO_1070 (O_1070,N_14898,N_14817);
nand UO_1071 (O_1071,N_14798,N_14912);
xor UO_1072 (O_1072,N_14922,N_14726);
nor UO_1073 (O_1073,N_14971,N_14726);
and UO_1074 (O_1074,N_14796,N_14956);
nor UO_1075 (O_1075,N_14875,N_14801);
nand UO_1076 (O_1076,N_14779,N_14836);
nor UO_1077 (O_1077,N_14806,N_14744);
xnor UO_1078 (O_1078,N_14845,N_14800);
and UO_1079 (O_1079,N_14726,N_14777);
nor UO_1080 (O_1080,N_14985,N_14870);
nand UO_1081 (O_1081,N_14821,N_14709);
xnor UO_1082 (O_1082,N_14843,N_14726);
xor UO_1083 (O_1083,N_14890,N_14831);
nor UO_1084 (O_1084,N_14867,N_14755);
nor UO_1085 (O_1085,N_14810,N_14835);
nor UO_1086 (O_1086,N_14932,N_14840);
nand UO_1087 (O_1087,N_14727,N_14833);
or UO_1088 (O_1088,N_14723,N_14769);
nor UO_1089 (O_1089,N_14908,N_14785);
nor UO_1090 (O_1090,N_14862,N_14891);
xor UO_1091 (O_1091,N_14785,N_14916);
or UO_1092 (O_1092,N_14986,N_14751);
nand UO_1093 (O_1093,N_14913,N_14743);
nor UO_1094 (O_1094,N_14768,N_14838);
xor UO_1095 (O_1095,N_14760,N_14892);
or UO_1096 (O_1096,N_14990,N_14885);
nor UO_1097 (O_1097,N_14948,N_14800);
or UO_1098 (O_1098,N_14701,N_14830);
and UO_1099 (O_1099,N_14754,N_14839);
or UO_1100 (O_1100,N_14966,N_14724);
or UO_1101 (O_1101,N_14899,N_14807);
nor UO_1102 (O_1102,N_14862,N_14775);
and UO_1103 (O_1103,N_14955,N_14821);
nor UO_1104 (O_1104,N_14747,N_14930);
nand UO_1105 (O_1105,N_14951,N_14928);
nor UO_1106 (O_1106,N_14845,N_14911);
and UO_1107 (O_1107,N_14709,N_14885);
xor UO_1108 (O_1108,N_14878,N_14798);
nor UO_1109 (O_1109,N_14934,N_14905);
or UO_1110 (O_1110,N_14921,N_14779);
nand UO_1111 (O_1111,N_14794,N_14936);
or UO_1112 (O_1112,N_14996,N_14741);
xnor UO_1113 (O_1113,N_14976,N_14751);
and UO_1114 (O_1114,N_14933,N_14774);
nor UO_1115 (O_1115,N_14742,N_14861);
and UO_1116 (O_1116,N_14957,N_14981);
xnor UO_1117 (O_1117,N_14948,N_14750);
nand UO_1118 (O_1118,N_14712,N_14857);
or UO_1119 (O_1119,N_14939,N_14824);
nor UO_1120 (O_1120,N_14818,N_14946);
or UO_1121 (O_1121,N_14716,N_14813);
xnor UO_1122 (O_1122,N_14943,N_14796);
nor UO_1123 (O_1123,N_14730,N_14826);
xor UO_1124 (O_1124,N_14900,N_14740);
nand UO_1125 (O_1125,N_14938,N_14815);
nand UO_1126 (O_1126,N_14731,N_14802);
xor UO_1127 (O_1127,N_14870,N_14806);
and UO_1128 (O_1128,N_14912,N_14991);
or UO_1129 (O_1129,N_14849,N_14963);
or UO_1130 (O_1130,N_14794,N_14860);
and UO_1131 (O_1131,N_14786,N_14718);
xor UO_1132 (O_1132,N_14953,N_14776);
nand UO_1133 (O_1133,N_14751,N_14918);
xor UO_1134 (O_1134,N_14786,N_14939);
xnor UO_1135 (O_1135,N_14924,N_14961);
xnor UO_1136 (O_1136,N_14906,N_14721);
xnor UO_1137 (O_1137,N_14910,N_14746);
xnor UO_1138 (O_1138,N_14860,N_14728);
nor UO_1139 (O_1139,N_14863,N_14784);
xnor UO_1140 (O_1140,N_14982,N_14768);
nand UO_1141 (O_1141,N_14973,N_14817);
xor UO_1142 (O_1142,N_14798,N_14704);
or UO_1143 (O_1143,N_14977,N_14962);
nand UO_1144 (O_1144,N_14982,N_14918);
nand UO_1145 (O_1145,N_14801,N_14842);
nor UO_1146 (O_1146,N_14976,N_14861);
xor UO_1147 (O_1147,N_14747,N_14954);
or UO_1148 (O_1148,N_14998,N_14855);
nand UO_1149 (O_1149,N_14974,N_14960);
nand UO_1150 (O_1150,N_14740,N_14824);
nor UO_1151 (O_1151,N_14940,N_14803);
xor UO_1152 (O_1152,N_14813,N_14971);
or UO_1153 (O_1153,N_14899,N_14784);
nor UO_1154 (O_1154,N_14844,N_14776);
or UO_1155 (O_1155,N_14734,N_14809);
nor UO_1156 (O_1156,N_14857,N_14778);
xnor UO_1157 (O_1157,N_14936,N_14910);
and UO_1158 (O_1158,N_14876,N_14731);
nand UO_1159 (O_1159,N_14744,N_14921);
nor UO_1160 (O_1160,N_14710,N_14901);
xor UO_1161 (O_1161,N_14860,N_14757);
nand UO_1162 (O_1162,N_14868,N_14971);
nor UO_1163 (O_1163,N_14799,N_14828);
and UO_1164 (O_1164,N_14809,N_14747);
xnor UO_1165 (O_1165,N_14879,N_14880);
nor UO_1166 (O_1166,N_14833,N_14783);
xor UO_1167 (O_1167,N_14746,N_14952);
or UO_1168 (O_1168,N_14869,N_14934);
nor UO_1169 (O_1169,N_14704,N_14943);
xnor UO_1170 (O_1170,N_14815,N_14801);
or UO_1171 (O_1171,N_14800,N_14702);
xor UO_1172 (O_1172,N_14954,N_14722);
nand UO_1173 (O_1173,N_14814,N_14736);
nand UO_1174 (O_1174,N_14719,N_14826);
nor UO_1175 (O_1175,N_14920,N_14730);
nand UO_1176 (O_1176,N_14866,N_14788);
xnor UO_1177 (O_1177,N_14929,N_14740);
or UO_1178 (O_1178,N_14942,N_14835);
and UO_1179 (O_1179,N_14978,N_14739);
nor UO_1180 (O_1180,N_14772,N_14784);
nor UO_1181 (O_1181,N_14723,N_14887);
or UO_1182 (O_1182,N_14893,N_14768);
nand UO_1183 (O_1183,N_14869,N_14831);
nand UO_1184 (O_1184,N_14754,N_14989);
nor UO_1185 (O_1185,N_14990,N_14776);
xnor UO_1186 (O_1186,N_14933,N_14877);
nand UO_1187 (O_1187,N_14779,N_14839);
nand UO_1188 (O_1188,N_14977,N_14774);
nand UO_1189 (O_1189,N_14771,N_14956);
nor UO_1190 (O_1190,N_14910,N_14802);
nand UO_1191 (O_1191,N_14773,N_14810);
nor UO_1192 (O_1192,N_14913,N_14965);
nor UO_1193 (O_1193,N_14870,N_14711);
or UO_1194 (O_1194,N_14810,N_14823);
xor UO_1195 (O_1195,N_14716,N_14901);
nand UO_1196 (O_1196,N_14826,N_14757);
xnor UO_1197 (O_1197,N_14763,N_14789);
or UO_1198 (O_1198,N_14724,N_14991);
xor UO_1199 (O_1199,N_14940,N_14967);
or UO_1200 (O_1200,N_14716,N_14893);
or UO_1201 (O_1201,N_14808,N_14777);
nand UO_1202 (O_1202,N_14849,N_14857);
nor UO_1203 (O_1203,N_14803,N_14841);
nor UO_1204 (O_1204,N_14801,N_14758);
nand UO_1205 (O_1205,N_14924,N_14778);
xor UO_1206 (O_1206,N_14826,N_14894);
nand UO_1207 (O_1207,N_14761,N_14841);
nor UO_1208 (O_1208,N_14811,N_14840);
and UO_1209 (O_1209,N_14790,N_14829);
xor UO_1210 (O_1210,N_14776,N_14840);
or UO_1211 (O_1211,N_14863,N_14966);
nor UO_1212 (O_1212,N_14736,N_14769);
xnor UO_1213 (O_1213,N_14944,N_14708);
nor UO_1214 (O_1214,N_14896,N_14837);
or UO_1215 (O_1215,N_14952,N_14912);
and UO_1216 (O_1216,N_14812,N_14920);
or UO_1217 (O_1217,N_14912,N_14705);
and UO_1218 (O_1218,N_14856,N_14708);
nor UO_1219 (O_1219,N_14748,N_14788);
nand UO_1220 (O_1220,N_14747,N_14771);
nand UO_1221 (O_1221,N_14973,N_14745);
and UO_1222 (O_1222,N_14782,N_14838);
nor UO_1223 (O_1223,N_14946,N_14805);
nand UO_1224 (O_1224,N_14748,N_14972);
nand UO_1225 (O_1225,N_14761,N_14780);
or UO_1226 (O_1226,N_14708,N_14988);
xnor UO_1227 (O_1227,N_14994,N_14740);
and UO_1228 (O_1228,N_14982,N_14872);
and UO_1229 (O_1229,N_14858,N_14841);
or UO_1230 (O_1230,N_14997,N_14764);
nor UO_1231 (O_1231,N_14999,N_14841);
and UO_1232 (O_1232,N_14703,N_14869);
nor UO_1233 (O_1233,N_14835,N_14960);
xnor UO_1234 (O_1234,N_14779,N_14708);
nand UO_1235 (O_1235,N_14866,N_14932);
nor UO_1236 (O_1236,N_14762,N_14711);
xnor UO_1237 (O_1237,N_14722,N_14818);
xnor UO_1238 (O_1238,N_14995,N_14732);
or UO_1239 (O_1239,N_14865,N_14960);
or UO_1240 (O_1240,N_14749,N_14765);
nor UO_1241 (O_1241,N_14744,N_14931);
and UO_1242 (O_1242,N_14769,N_14750);
or UO_1243 (O_1243,N_14980,N_14757);
or UO_1244 (O_1244,N_14759,N_14710);
nand UO_1245 (O_1245,N_14853,N_14854);
xor UO_1246 (O_1246,N_14779,N_14890);
and UO_1247 (O_1247,N_14926,N_14822);
nand UO_1248 (O_1248,N_14816,N_14821);
or UO_1249 (O_1249,N_14885,N_14964);
and UO_1250 (O_1250,N_14897,N_14925);
nor UO_1251 (O_1251,N_14918,N_14826);
nor UO_1252 (O_1252,N_14863,N_14953);
nand UO_1253 (O_1253,N_14736,N_14900);
nor UO_1254 (O_1254,N_14890,N_14906);
nand UO_1255 (O_1255,N_14856,N_14761);
and UO_1256 (O_1256,N_14723,N_14783);
or UO_1257 (O_1257,N_14980,N_14817);
or UO_1258 (O_1258,N_14705,N_14852);
nand UO_1259 (O_1259,N_14831,N_14754);
nand UO_1260 (O_1260,N_14786,N_14719);
and UO_1261 (O_1261,N_14851,N_14950);
xor UO_1262 (O_1262,N_14945,N_14858);
xor UO_1263 (O_1263,N_14942,N_14872);
or UO_1264 (O_1264,N_14885,N_14779);
and UO_1265 (O_1265,N_14740,N_14760);
nand UO_1266 (O_1266,N_14828,N_14970);
xor UO_1267 (O_1267,N_14954,N_14755);
nor UO_1268 (O_1268,N_14781,N_14941);
or UO_1269 (O_1269,N_14789,N_14775);
or UO_1270 (O_1270,N_14870,N_14846);
xor UO_1271 (O_1271,N_14712,N_14771);
or UO_1272 (O_1272,N_14856,N_14871);
nand UO_1273 (O_1273,N_14835,N_14907);
xnor UO_1274 (O_1274,N_14710,N_14920);
nand UO_1275 (O_1275,N_14823,N_14996);
and UO_1276 (O_1276,N_14798,N_14706);
nand UO_1277 (O_1277,N_14981,N_14858);
xnor UO_1278 (O_1278,N_14993,N_14840);
and UO_1279 (O_1279,N_14878,N_14725);
or UO_1280 (O_1280,N_14722,N_14856);
nand UO_1281 (O_1281,N_14704,N_14796);
nor UO_1282 (O_1282,N_14822,N_14773);
nor UO_1283 (O_1283,N_14965,N_14807);
or UO_1284 (O_1284,N_14919,N_14787);
nand UO_1285 (O_1285,N_14785,N_14714);
xor UO_1286 (O_1286,N_14883,N_14841);
and UO_1287 (O_1287,N_14969,N_14877);
and UO_1288 (O_1288,N_14810,N_14761);
nor UO_1289 (O_1289,N_14910,N_14826);
xnor UO_1290 (O_1290,N_14777,N_14877);
nor UO_1291 (O_1291,N_14943,N_14724);
and UO_1292 (O_1292,N_14886,N_14824);
nor UO_1293 (O_1293,N_14781,N_14738);
nor UO_1294 (O_1294,N_14871,N_14989);
and UO_1295 (O_1295,N_14716,N_14843);
or UO_1296 (O_1296,N_14700,N_14720);
and UO_1297 (O_1297,N_14703,N_14769);
nand UO_1298 (O_1298,N_14960,N_14973);
and UO_1299 (O_1299,N_14991,N_14825);
or UO_1300 (O_1300,N_14981,N_14808);
nand UO_1301 (O_1301,N_14839,N_14960);
nand UO_1302 (O_1302,N_14725,N_14998);
nor UO_1303 (O_1303,N_14744,N_14822);
nor UO_1304 (O_1304,N_14827,N_14770);
nor UO_1305 (O_1305,N_14951,N_14995);
nand UO_1306 (O_1306,N_14771,N_14819);
and UO_1307 (O_1307,N_14963,N_14910);
and UO_1308 (O_1308,N_14857,N_14706);
or UO_1309 (O_1309,N_14838,N_14858);
xor UO_1310 (O_1310,N_14749,N_14746);
xnor UO_1311 (O_1311,N_14713,N_14793);
nor UO_1312 (O_1312,N_14733,N_14921);
or UO_1313 (O_1313,N_14808,N_14908);
xor UO_1314 (O_1314,N_14998,N_14958);
xnor UO_1315 (O_1315,N_14861,N_14858);
or UO_1316 (O_1316,N_14827,N_14803);
xor UO_1317 (O_1317,N_14906,N_14727);
xnor UO_1318 (O_1318,N_14743,N_14802);
nor UO_1319 (O_1319,N_14835,N_14818);
and UO_1320 (O_1320,N_14897,N_14743);
xor UO_1321 (O_1321,N_14752,N_14953);
or UO_1322 (O_1322,N_14825,N_14845);
nor UO_1323 (O_1323,N_14835,N_14933);
nor UO_1324 (O_1324,N_14985,N_14775);
and UO_1325 (O_1325,N_14738,N_14855);
xor UO_1326 (O_1326,N_14884,N_14965);
nor UO_1327 (O_1327,N_14949,N_14734);
and UO_1328 (O_1328,N_14921,N_14761);
nand UO_1329 (O_1329,N_14761,N_14762);
xor UO_1330 (O_1330,N_14912,N_14954);
xor UO_1331 (O_1331,N_14810,N_14894);
and UO_1332 (O_1332,N_14816,N_14859);
nand UO_1333 (O_1333,N_14825,N_14708);
and UO_1334 (O_1334,N_14708,N_14800);
and UO_1335 (O_1335,N_14756,N_14931);
or UO_1336 (O_1336,N_14762,N_14947);
nand UO_1337 (O_1337,N_14849,N_14987);
and UO_1338 (O_1338,N_14832,N_14788);
nand UO_1339 (O_1339,N_14807,N_14872);
nor UO_1340 (O_1340,N_14909,N_14813);
nor UO_1341 (O_1341,N_14983,N_14887);
xnor UO_1342 (O_1342,N_14957,N_14885);
and UO_1343 (O_1343,N_14938,N_14718);
nor UO_1344 (O_1344,N_14938,N_14894);
and UO_1345 (O_1345,N_14960,N_14815);
and UO_1346 (O_1346,N_14740,N_14703);
nand UO_1347 (O_1347,N_14912,N_14996);
nand UO_1348 (O_1348,N_14801,N_14840);
and UO_1349 (O_1349,N_14861,N_14820);
xnor UO_1350 (O_1350,N_14926,N_14923);
and UO_1351 (O_1351,N_14739,N_14945);
or UO_1352 (O_1352,N_14719,N_14727);
nor UO_1353 (O_1353,N_14954,N_14740);
nand UO_1354 (O_1354,N_14804,N_14990);
nor UO_1355 (O_1355,N_14788,N_14781);
xor UO_1356 (O_1356,N_14975,N_14854);
nor UO_1357 (O_1357,N_14960,N_14762);
nor UO_1358 (O_1358,N_14848,N_14753);
or UO_1359 (O_1359,N_14982,N_14875);
xor UO_1360 (O_1360,N_14925,N_14788);
and UO_1361 (O_1361,N_14731,N_14950);
nand UO_1362 (O_1362,N_14831,N_14779);
and UO_1363 (O_1363,N_14826,N_14927);
xnor UO_1364 (O_1364,N_14746,N_14941);
nor UO_1365 (O_1365,N_14938,N_14826);
or UO_1366 (O_1366,N_14916,N_14901);
nor UO_1367 (O_1367,N_14915,N_14887);
and UO_1368 (O_1368,N_14812,N_14856);
or UO_1369 (O_1369,N_14816,N_14892);
or UO_1370 (O_1370,N_14942,N_14714);
and UO_1371 (O_1371,N_14760,N_14786);
nor UO_1372 (O_1372,N_14760,N_14737);
xnor UO_1373 (O_1373,N_14856,N_14781);
nor UO_1374 (O_1374,N_14909,N_14750);
or UO_1375 (O_1375,N_14895,N_14771);
nand UO_1376 (O_1376,N_14749,N_14995);
or UO_1377 (O_1377,N_14746,N_14859);
and UO_1378 (O_1378,N_14780,N_14813);
nand UO_1379 (O_1379,N_14736,N_14756);
or UO_1380 (O_1380,N_14724,N_14992);
or UO_1381 (O_1381,N_14917,N_14720);
or UO_1382 (O_1382,N_14744,N_14788);
nor UO_1383 (O_1383,N_14707,N_14762);
xor UO_1384 (O_1384,N_14702,N_14900);
nor UO_1385 (O_1385,N_14869,N_14860);
or UO_1386 (O_1386,N_14845,N_14892);
and UO_1387 (O_1387,N_14825,N_14903);
nor UO_1388 (O_1388,N_14903,N_14962);
or UO_1389 (O_1389,N_14936,N_14722);
and UO_1390 (O_1390,N_14763,N_14881);
nand UO_1391 (O_1391,N_14726,N_14821);
and UO_1392 (O_1392,N_14937,N_14921);
xor UO_1393 (O_1393,N_14817,N_14729);
nor UO_1394 (O_1394,N_14709,N_14829);
and UO_1395 (O_1395,N_14873,N_14841);
nand UO_1396 (O_1396,N_14738,N_14919);
nand UO_1397 (O_1397,N_14836,N_14948);
and UO_1398 (O_1398,N_14740,N_14958);
nand UO_1399 (O_1399,N_14762,N_14808);
and UO_1400 (O_1400,N_14802,N_14988);
nor UO_1401 (O_1401,N_14953,N_14909);
nand UO_1402 (O_1402,N_14819,N_14817);
xnor UO_1403 (O_1403,N_14980,N_14831);
and UO_1404 (O_1404,N_14740,N_14721);
or UO_1405 (O_1405,N_14768,N_14742);
xnor UO_1406 (O_1406,N_14726,N_14999);
or UO_1407 (O_1407,N_14836,N_14982);
nor UO_1408 (O_1408,N_14942,N_14832);
and UO_1409 (O_1409,N_14985,N_14786);
and UO_1410 (O_1410,N_14765,N_14886);
and UO_1411 (O_1411,N_14987,N_14884);
or UO_1412 (O_1412,N_14794,N_14762);
and UO_1413 (O_1413,N_14819,N_14958);
nand UO_1414 (O_1414,N_14828,N_14703);
nor UO_1415 (O_1415,N_14988,N_14730);
nor UO_1416 (O_1416,N_14941,N_14994);
xnor UO_1417 (O_1417,N_14885,N_14867);
and UO_1418 (O_1418,N_14858,N_14750);
and UO_1419 (O_1419,N_14708,N_14795);
nor UO_1420 (O_1420,N_14923,N_14876);
nand UO_1421 (O_1421,N_14778,N_14773);
xnor UO_1422 (O_1422,N_14953,N_14841);
or UO_1423 (O_1423,N_14755,N_14836);
nand UO_1424 (O_1424,N_14829,N_14901);
and UO_1425 (O_1425,N_14802,N_14724);
nand UO_1426 (O_1426,N_14753,N_14925);
nand UO_1427 (O_1427,N_14946,N_14963);
xnor UO_1428 (O_1428,N_14797,N_14782);
xor UO_1429 (O_1429,N_14988,N_14889);
nor UO_1430 (O_1430,N_14816,N_14844);
xor UO_1431 (O_1431,N_14788,N_14821);
nand UO_1432 (O_1432,N_14976,N_14954);
or UO_1433 (O_1433,N_14945,N_14981);
xor UO_1434 (O_1434,N_14899,N_14730);
and UO_1435 (O_1435,N_14700,N_14903);
nand UO_1436 (O_1436,N_14793,N_14930);
or UO_1437 (O_1437,N_14873,N_14863);
nand UO_1438 (O_1438,N_14768,N_14883);
nand UO_1439 (O_1439,N_14830,N_14886);
xor UO_1440 (O_1440,N_14776,N_14800);
and UO_1441 (O_1441,N_14848,N_14817);
xnor UO_1442 (O_1442,N_14745,N_14736);
nand UO_1443 (O_1443,N_14867,N_14717);
and UO_1444 (O_1444,N_14735,N_14817);
xor UO_1445 (O_1445,N_14769,N_14714);
and UO_1446 (O_1446,N_14940,N_14930);
nand UO_1447 (O_1447,N_14857,N_14773);
and UO_1448 (O_1448,N_14726,N_14797);
nand UO_1449 (O_1449,N_14780,N_14716);
and UO_1450 (O_1450,N_14927,N_14871);
and UO_1451 (O_1451,N_14756,N_14893);
xnor UO_1452 (O_1452,N_14827,N_14787);
and UO_1453 (O_1453,N_14829,N_14835);
nor UO_1454 (O_1454,N_14975,N_14734);
nand UO_1455 (O_1455,N_14770,N_14714);
or UO_1456 (O_1456,N_14958,N_14704);
xnor UO_1457 (O_1457,N_14788,N_14782);
nand UO_1458 (O_1458,N_14826,N_14940);
and UO_1459 (O_1459,N_14747,N_14950);
nand UO_1460 (O_1460,N_14795,N_14774);
nand UO_1461 (O_1461,N_14701,N_14866);
nand UO_1462 (O_1462,N_14743,N_14900);
or UO_1463 (O_1463,N_14747,N_14874);
and UO_1464 (O_1464,N_14974,N_14834);
nor UO_1465 (O_1465,N_14933,N_14907);
and UO_1466 (O_1466,N_14858,N_14881);
nand UO_1467 (O_1467,N_14893,N_14770);
nor UO_1468 (O_1468,N_14729,N_14814);
xor UO_1469 (O_1469,N_14753,N_14810);
or UO_1470 (O_1470,N_14941,N_14724);
nor UO_1471 (O_1471,N_14927,N_14919);
or UO_1472 (O_1472,N_14804,N_14981);
xor UO_1473 (O_1473,N_14983,N_14866);
xnor UO_1474 (O_1474,N_14741,N_14978);
or UO_1475 (O_1475,N_14705,N_14869);
nand UO_1476 (O_1476,N_14755,N_14935);
and UO_1477 (O_1477,N_14977,N_14897);
nand UO_1478 (O_1478,N_14806,N_14755);
or UO_1479 (O_1479,N_14829,N_14844);
and UO_1480 (O_1480,N_14941,N_14989);
nor UO_1481 (O_1481,N_14908,N_14787);
xor UO_1482 (O_1482,N_14925,N_14850);
or UO_1483 (O_1483,N_14818,N_14857);
nor UO_1484 (O_1484,N_14948,N_14965);
nand UO_1485 (O_1485,N_14977,N_14917);
and UO_1486 (O_1486,N_14923,N_14892);
and UO_1487 (O_1487,N_14802,N_14858);
nor UO_1488 (O_1488,N_14925,N_14968);
and UO_1489 (O_1489,N_14863,N_14752);
nor UO_1490 (O_1490,N_14884,N_14738);
or UO_1491 (O_1491,N_14716,N_14806);
xnor UO_1492 (O_1492,N_14944,N_14960);
nand UO_1493 (O_1493,N_14706,N_14813);
nand UO_1494 (O_1494,N_14927,N_14843);
or UO_1495 (O_1495,N_14854,N_14840);
nand UO_1496 (O_1496,N_14973,N_14989);
nor UO_1497 (O_1497,N_14837,N_14933);
xnor UO_1498 (O_1498,N_14909,N_14954);
or UO_1499 (O_1499,N_14736,N_14781);
nand UO_1500 (O_1500,N_14897,N_14737);
xnor UO_1501 (O_1501,N_14953,N_14720);
xor UO_1502 (O_1502,N_14962,N_14772);
and UO_1503 (O_1503,N_14915,N_14749);
xnor UO_1504 (O_1504,N_14801,N_14813);
xor UO_1505 (O_1505,N_14795,N_14980);
nor UO_1506 (O_1506,N_14840,N_14906);
or UO_1507 (O_1507,N_14750,N_14731);
and UO_1508 (O_1508,N_14881,N_14745);
and UO_1509 (O_1509,N_14822,N_14766);
nand UO_1510 (O_1510,N_14721,N_14980);
nor UO_1511 (O_1511,N_14969,N_14703);
nor UO_1512 (O_1512,N_14738,N_14826);
or UO_1513 (O_1513,N_14850,N_14707);
nand UO_1514 (O_1514,N_14962,N_14935);
xor UO_1515 (O_1515,N_14975,N_14960);
nand UO_1516 (O_1516,N_14753,N_14806);
and UO_1517 (O_1517,N_14927,N_14778);
nor UO_1518 (O_1518,N_14744,N_14897);
nor UO_1519 (O_1519,N_14735,N_14824);
nor UO_1520 (O_1520,N_14823,N_14740);
xnor UO_1521 (O_1521,N_14826,N_14743);
or UO_1522 (O_1522,N_14793,N_14939);
nand UO_1523 (O_1523,N_14768,N_14764);
and UO_1524 (O_1524,N_14878,N_14967);
nand UO_1525 (O_1525,N_14849,N_14926);
and UO_1526 (O_1526,N_14757,N_14906);
nor UO_1527 (O_1527,N_14760,N_14819);
nand UO_1528 (O_1528,N_14766,N_14879);
or UO_1529 (O_1529,N_14743,N_14715);
nor UO_1530 (O_1530,N_14806,N_14884);
nor UO_1531 (O_1531,N_14872,N_14837);
and UO_1532 (O_1532,N_14965,N_14789);
nor UO_1533 (O_1533,N_14718,N_14945);
and UO_1534 (O_1534,N_14950,N_14857);
nand UO_1535 (O_1535,N_14708,N_14744);
and UO_1536 (O_1536,N_14814,N_14728);
nand UO_1537 (O_1537,N_14787,N_14732);
and UO_1538 (O_1538,N_14711,N_14712);
nand UO_1539 (O_1539,N_14869,N_14804);
and UO_1540 (O_1540,N_14796,N_14781);
xnor UO_1541 (O_1541,N_14878,N_14857);
nand UO_1542 (O_1542,N_14998,N_14719);
nand UO_1543 (O_1543,N_14940,N_14860);
nand UO_1544 (O_1544,N_14804,N_14717);
or UO_1545 (O_1545,N_14713,N_14817);
nor UO_1546 (O_1546,N_14985,N_14959);
xnor UO_1547 (O_1547,N_14733,N_14747);
nand UO_1548 (O_1548,N_14860,N_14739);
xnor UO_1549 (O_1549,N_14757,N_14895);
nand UO_1550 (O_1550,N_14978,N_14865);
or UO_1551 (O_1551,N_14855,N_14859);
xnor UO_1552 (O_1552,N_14744,N_14790);
and UO_1553 (O_1553,N_14751,N_14701);
xor UO_1554 (O_1554,N_14854,N_14961);
nor UO_1555 (O_1555,N_14920,N_14902);
and UO_1556 (O_1556,N_14900,N_14766);
and UO_1557 (O_1557,N_14845,N_14812);
nand UO_1558 (O_1558,N_14981,N_14726);
nor UO_1559 (O_1559,N_14731,N_14907);
or UO_1560 (O_1560,N_14832,N_14888);
nand UO_1561 (O_1561,N_14869,N_14700);
nor UO_1562 (O_1562,N_14755,N_14819);
nand UO_1563 (O_1563,N_14979,N_14780);
or UO_1564 (O_1564,N_14995,N_14742);
and UO_1565 (O_1565,N_14903,N_14898);
nand UO_1566 (O_1566,N_14731,N_14875);
xor UO_1567 (O_1567,N_14943,N_14995);
and UO_1568 (O_1568,N_14931,N_14757);
or UO_1569 (O_1569,N_14881,N_14988);
or UO_1570 (O_1570,N_14753,N_14997);
and UO_1571 (O_1571,N_14986,N_14934);
or UO_1572 (O_1572,N_14770,N_14752);
xnor UO_1573 (O_1573,N_14719,N_14751);
xor UO_1574 (O_1574,N_14920,N_14962);
and UO_1575 (O_1575,N_14728,N_14863);
or UO_1576 (O_1576,N_14747,N_14729);
xor UO_1577 (O_1577,N_14717,N_14963);
or UO_1578 (O_1578,N_14945,N_14979);
or UO_1579 (O_1579,N_14996,N_14895);
nand UO_1580 (O_1580,N_14770,N_14947);
xnor UO_1581 (O_1581,N_14788,N_14809);
and UO_1582 (O_1582,N_14928,N_14855);
or UO_1583 (O_1583,N_14889,N_14943);
and UO_1584 (O_1584,N_14830,N_14871);
nand UO_1585 (O_1585,N_14744,N_14941);
and UO_1586 (O_1586,N_14970,N_14800);
nor UO_1587 (O_1587,N_14859,N_14927);
xnor UO_1588 (O_1588,N_14806,N_14728);
or UO_1589 (O_1589,N_14751,N_14724);
xnor UO_1590 (O_1590,N_14831,N_14738);
nor UO_1591 (O_1591,N_14832,N_14983);
nor UO_1592 (O_1592,N_14932,N_14935);
nand UO_1593 (O_1593,N_14931,N_14789);
and UO_1594 (O_1594,N_14987,N_14877);
xor UO_1595 (O_1595,N_14790,N_14799);
or UO_1596 (O_1596,N_14982,N_14929);
nand UO_1597 (O_1597,N_14781,N_14729);
nand UO_1598 (O_1598,N_14797,N_14764);
nor UO_1599 (O_1599,N_14798,N_14963);
nand UO_1600 (O_1600,N_14940,N_14858);
nor UO_1601 (O_1601,N_14980,N_14876);
nor UO_1602 (O_1602,N_14835,N_14975);
nor UO_1603 (O_1603,N_14965,N_14717);
xnor UO_1604 (O_1604,N_14743,N_14906);
and UO_1605 (O_1605,N_14768,N_14959);
or UO_1606 (O_1606,N_14760,N_14830);
xor UO_1607 (O_1607,N_14923,N_14860);
nor UO_1608 (O_1608,N_14718,N_14811);
nand UO_1609 (O_1609,N_14795,N_14966);
xnor UO_1610 (O_1610,N_14915,N_14723);
and UO_1611 (O_1611,N_14748,N_14881);
or UO_1612 (O_1612,N_14723,N_14968);
xnor UO_1613 (O_1613,N_14867,N_14915);
xnor UO_1614 (O_1614,N_14938,N_14879);
and UO_1615 (O_1615,N_14884,N_14721);
nor UO_1616 (O_1616,N_14961,N_14737);
and UO_1617 (O_1617,N_14937,N_14823);
or UO_1618 (O_1618,N_14827,N_14713);
nor UO_1619 (O_1619,N_14824,N_14880);
or UO_1620 (O_1620,N_14967,N_14759);
and UO_1621 (O_1621,N_14804,N_14789);
and UO_1622 (O_1622,N_14776,N_14966);
nand UO_1623 (O_1623,N_14896,N_14734);
nor UO_1624 (O_1624,N_14966,N_14880);
nand UO_1625 (O_1625,N_14950,N_14874);
or UO_1626 (O_1626,N_14880,N_14954);
nand UO_1627 (O_1627,N_14901,N_14800);
nand UO_1628 (O_1628,N_14862,N_14721);
xnor UO_1629 (O_1629,N_14936,N_14976);
xnor UO_1630 (O_1630,N_14956,N_14712);
xnor UO_1631 (O_1631,N_14866,N_14834);
or UO_1632 (O_1632,N_14961,N_14985);
or UO_1633 (O_1633,N_14793,N_14943);
xnor UO_1634 (O_1634,N_14730,N_14774);
nor UO_1635 (O_1635,N_14779,N_14705);
and UO_1636 (O_1636,N_14909,N_14748);
nand UO_1637 (O_1637,N_14807,N_14794);
nand UO_1638 (O_1638,N_14898,N_14942);
nand UO_1639 (O_1639,N_14892,N_14793);
xnor UO_1640 (O_1640,N_14771,N_14718);
nand UO_1641 (O_1641,N_14857,N_14915);
and UO_1642 (O_1642,N_14955,N_14898);
or UO_1643 (O_1643,N_14775,N_14829);
and UO_1644 (O_1644,N_14883,N_14720);
and UO_1645 (O_1645,N_14996,N_14850);
and UO_1646 (O_1646,N_14863,N_14853);
and UO_1647 (O_1647,N_14820,N_14940);
and UO_1648 (O_1648,N_14838,N_14824);
xnor UO_1649 (O_1649,N_14735,N_14898);
nor UO_1650 (O_1650,N_14834,N_14806);
nand UO_1651 (O_1651,N_14933,N_14897);
and UO_1652 (O_1652,N_14765,N_14995);
and UO_1653 (O_1653,N_14945,N_14800);
or UO_1654 (O_1654,N_14755,N_14882);
nand UO_1655 (O_1655,N_14800,N_14829);
nand UO_1656 (O_1656,N_14953,N_14906);
and UO_1657 (O_1657,N_14851,N_14948);
xor UO_1658 (O_1658,N_14844,N_14925);
nand UO_1659 (O_1659,N_14915,N_14833);
nor UO_1660 (O_1660,N_14991,N_14946);
xor UO_1661 (O_1661,N_14908,N_14736);
and UO_1662 (O_1662,N_14879,N_14844);
xor UO_1663 (O_1663,N_14977,N_14939);
nor UO_1664 (O_1664,N_14733,N_14744);
nor UO_1665 (O_1665,N_14785,N_14971);
nor UO_1666 (O_1666,N_14800,N_14937);
nor UO_1667 (O_1667,N_14848,N_14993);
xor UO_1668 (O_1668,N_14956,N_14871);
xnor UO_1669 (O_1669,N_14718,N_14716);
nor UO_1670 (O_1670,N_14795,N_14927);
and UO_1671 (O_1671,N_14907,N_14828);
or UO_1672 (O_1672,N_14944,N_14801);
nor UO_1673 (O_1673,N_14847,N_14996);
xor UO_1674 (O_1674,N_14811,N_14716);
or UO_1675 (O_1675,N_14722,N_14804);
and UO_1676 (O_1676,N_14857,N_14941);
or UO_1677 (O_1677,N_14835,N_14789);
nand UO_1678 (O_1678,N_14777,N_14875);
nand UO_1679 (O_1679,N_14741,N_14830);
or UO_1680 (O_1680,N_14815,N_14711);
nor UO_1681 (O_1681,N_14999,N_14739);
nand UO_1682 (O_1682,N_14755,N_14723);
and UO_1683 (O_1683,N_14864,N_14806);
nor UO_1684 (O_1684,N_14816,N_14933);
or UO_1685 (O_1685,N_14888,N_14752);
xor UO_1686 (O_1686,N_14872,N_14884);
xor UO_1687 (O_1687,N_14712,N_14960);
xor UO_1688 (O_1688,N_14837,N_14784);
and UO_1689 (O_1689,N_14876,N_14941);
nor UO_1690 (O_1690,N_14891,N_14850);
nand UO_1691 (O_1691,N_14982,N_14951);
xnor UO_1692 (O_1692,N_14868,N_14934);
and UO_1693 (O_1693,N_14861,N_14880);
or UO_1694 (O_1694,N_14758,N_14942);
and UO_1695 (O_1695,N_14880,N_14899);
and UO_1696 (O_1696,N_14968,N_14955);
nand UO_1697 (O_1697,N_14796,N_14903);
nor UO_1698 (O_1698,N_14932,N_14781);
or UO_1699 (O_1699,N_14919,N_14709);
xor UO_1700 (O_1700,N_14866,N_14999);
nor UO_1701 (O_1701,N_14802,N_14804);
and UO_1702 (O_1702,N_14816,N_14915);
or UO_1703 (O_1703,N_14899,N_14700);
or UO_1704 (O_1704,N_14950,N_14816);
nor UO_1705 (O_1705,N_14917,N_14712);
or UO_1706 (O_1706,N_14899,N_14913);
and UO_1707 (O_1707,N_14751,N_14768);
xnor UO_1708 (O_1708,N_14976,N_14881);
or UO_1709 (O_1709,N_14782,N_14789);
and UO_1710 (O_1710,N_14845,N_14923);
nand UO_1711 (O_1711,N_14764,N_14861);
or UO_1712 (O_1712,N_14796,N_14968);
nor UO_1713 (O_1713,N_14846,N_14864);
and UO_1714 (O_1714,N_14846,N_14944);
and UO_1715 (O_1715,N_14785,N_14959);
nor UO_1716 (O_1716,N_14962,N_14879);
xnor UO_1717 (O_1717,N_14937,N_14977);
xnor UO_1718 (O_1718,N_14898,N_14808);
nand UO_1719 (O_1719,N_14742,N_14793);
nor UO_1720 (O_1720,N_14870,N_14733);
nand UO_1721 (O_1721,N_14778,N_14851);
or UO_1722 (O_1722,N_14915,N_14714);
nand UO_1723 (O_1723,N_14893,N_14818);
or UO_1724 (O_1724,N_14852,N_14995);
xor UO_1725 (O_1725,N_14965,N_14809);
and UO_1726 (O_1726,N_14918,N_14915);
and UO_1727 (O_1727,N_14954,N_14999);
or UO_1728 (O_1728,N_14889,N_14939);
nand UO_1729 (O_1729,N_14989,N_14726);
nand UO_1730 (O_1730,N_14999,N_14754);
nor UO_1731 (O_1731,N_14831,N_14789);
nor UO_1732 (O_1732,N_14919,N_14768);
and UO_1733 (O_1733,N_14703,N_14719);
or UO_1734 (O_1734,N_14847,N_14831);
nand UO_1735 (O_1735,N_14901,N_14939);
nand UO_1736 (O_1736,N_14768,N_14779);
nand UO_1737 (O_1737,N_14795,N_14965);
and UO_1738 (O_1738,N_14732,N_14770);
or UO_1739 (O_1739,N_14998,N_14759);
nand UO_1740 (O_1740,N_14765,N_14984);
nor UO_1741 (O_1741,N_14873,N_14724);
nor UO_1742 (O_1742,N_14741,N_14761);
or UO_1743 (O_1743,N_14852,N_14975);
xor UO_1744 (O_1744,N_14987,N_14956);
nand UO_1745 (O_1745,N_14836,N_14745);
and UO_1746 (O_1746,N_14826,N_14987);
xor UO_1747 (O_1747,N_14958,N_14972);
or UO_1748 (O_1748,N_14785,N_14995);
nor UO_1749 (O_1749,N_14744,N_14729);
or UO_1750 (O_1750,N_14995,N_14783);
or UO_1751 (O_1751,N_14782,N_14815);
nor UO_1752 (O_1752,N_14791,N_14766);
nand UO_1753 (O_1753,N_14954,N_14883);
or UO_1754 (O_1754,N_14821,N_14910);
and UO_1755 (O_1755,N_14976,N_14915);
xnor UO_1756 (O_1756,N_14960,N_14896);
nand UO_1757 (O_1757,N_14985,N_14832);
nor UO_1758 (O_1758,N_14734,N_14748);
nor UO_1759 (O_1759,N_14819,N_14887);
or UO_1760 (O_1760,N_14903,N_14860);
nor UO_1761 (O_1761,N_14952,N_14974);
or UO_1762 (O_1762,N_14941,N_14962);
nand UO_1763 (O_1763,N_14748,N_14926);
nor UO_1764 (O_1764,N_14780,N_14762);
and UO_1765 (O_1765,N_14716,N_14914);
xor UO_1766 (O_1766,N_14974,N_14840);
or UO_1767 (O_1767,N_14787,N_14999);
or UO_1768 (O_1768,N_14742,N_14814);
and UO_1769 (O_1769,N_14944,N_14994);
nor UO_1770 (O_1770,N_14889,N_14953);
xor UO_1771 (O_1771,N_14996,N_14884);
nor UO_1772 (O_1772,N_14889,N_14903);
nand UO_1773 (O_1773,N_14777,N_14949);
and UO_1774 (O_1774,N_14822,N_14952);
nor UO_1775 (O_1775,N_14817,N_14895);
nand UO_1776 (O_1776,N_14823,N_14965);
or UO_1777 (O_1777,N_14982,N_14924);
xor UO_1778 (O_1778,N_14901,N_14922);
xor UO_1779 (O_1779,N_14811,N_14983);
nand UO_1780 (O_1780,N_14908,N_14967);
nand UO_1781 (O_1781,N_14849,N_14906);
or UO_1782 (O_1782,N_14882,N_14730);
nor UO_1783 (O_1783,N_14845,N_14909);
and UO_1784 (O_1784,N_14941,N_14881);
and UO_1785 (O_1785,N_14805,N_14847);
nor UO_1786 (O_1786,N_14792,N_14955);
xor UO_1787 (O_1787,N_14938,N_14800);
xnor UO_1788 (O_1788,N_14812,N_14712);
nand UO_1789 (O_1789,N_14799,N_14804);
or UO_1790 (O_1790,N_14801,N_14762);
and UO_1791 (O_1791,N_14718,N_14888);
xnor UO_1792 (O_1792,N_14950,N_14791);
or UO_1793 (O_1793,N_14993,N_14793);
nor UO_1794 (O_1794,N_14883,N_14973);
and UO_1795 (O_1795,N_14971,N_14847);
or UO_1796 (O_1796,N_14969,N_14818);
or UO_1797 (O_1797,N_14751,N_14814);
nor UO_1798 (O_1798,N_14873,N_14915);
or UO_1799 (O_1799,N_14776,N_14832);
and UO_1800 (O_1800,N_14750,N_14907);
xor UO_1801 (O_1801,N_14969,N_14708);
nand UO_1802 (O_1802,N_14913,N_14990);
nor UO_1803 (O_1803,N_14739,N_14962);
nand UO_1804 (O_1804,N_14963,N_14869);
nand UO_1805 (O_1805,N_14751,N_14885);
or UO_1806 (O_1806,N_14845,N_14798);
and UO_1807 (O_1807,N_14951,N_14964);
xor UO_1808 (O_1808,N_14866,N_14918);
or UO_1809 (O_1809,N_14758,N_14849);
xnor UO_1810 (O_1810,N_14905,N_14986);
and UO_1811 (O_1811,N_14904,N_14987);
or UO_1812 (O_1812,N_14747,N_14973);
nand UO_1813 (O_1813,N_14869,N_14764);
nor UO_1814 (O_1814,N_14704,N_14783);
nand UO_1815 (O_1815,N_14911,N_14875);
xor UO_1816 (O_1816,N_14866,N_14716);
nand UO_1817 (O_1817,N_14842,N_14831);
and UO_1818 (O_1818,N_14873,N_14785);
and UO_1819 (O_1819,N_14864,N_14760);
nor UO_1820 (O_1820,N_14886,N_14742);
nand UO_1821 (O_1821,N_14949,N_14980);
or UO_1822 (O_1822,N_14711,N_14919);
nand UO_1823 (O_1823,N_14847,N_14846);
or UO_1824 (O_1824,N_14713,N_14937);
or UO_1825 (O_1825,N_14909,N_14859);
xor UO_1826 (O_1826,N_14988,N_14965);
nand UO_1827 (O_1827,N_14764,N_14716);
xor UO_1828 (O_1828,N_14887,N_14841);
or UO_1829 (O_1829,N_14995,N_14987);
xor UO_1830 (O_1830,N_14797,N_14825);
xor UO_1831 (O_1831,N_14940,N_14948);
nand UO_1832 (O_1832,N_14937,N_14859);
xnor UO_1833 (O_1833,N_14796,N_14805);
or UO_1834 (O_1834,N_14943,N_14736);
xnor UO_1835 (O_1835,N_14723,N_14799);
xnor UO_1836 (O_1836,N_14957,N_14710);
and UO_1837 (O_1837,N_14909,N_14858);
or UO_1838 (O_1838,N_14929,N_14912);
nor UO_1839 (O_1839,N_14929,N_14913);
and UO_1840 (O_1840,N_14819,N_14823);
nand UO_1841 (O_1841,N_14845,N_14721);
nor UO_1842 (O_1842,N_14743,N_14851);
and UO_1843 (O_1843,N_14987,N_14878);
and UO_1844 (O_1844,N_14720,N_14967);
or UO_1845 (O_1845,N_14861,N_14881);
nand UO_1846 (O_1846,N_14977,N_14726);
or UO_1847 (O_1847,N_14888,N_14757);
xor UO_1848 (O_1848,N_14823,N_14741);
or UO_1849 (O_1849,N_14770,N_14795);
nand UO_1850 (O_1850,N_14755,N_14889);
and UO_1851 (O_1851,N_14775,N_14835);
nor UO_1852 (O_1852,N_14949,N_14935);
or UO_1853 (O_1853,N_14987,N_14707);
and UO_1854 (O_1854,N_14943,N_14875);
nor UO_1855 (O_1855,N_14704,N_14984);
nor UO_1856 (O_1856,N_14976,N_14731);
nor UO_1857 (O_1857,N_14913,N_14769);
and UO_1858 (O_1858,N_14780,N_14970);
and UO_1859 (O_1859,N_14947,N_14970);
or UO_1860 (O_1860,N_14707,N_14774);
and UO_1861 (O_1861,N_14912,N_14863);
nand UO_1862 (O_1862,N_14999,N_14946);
or UO_1863 (O_1863,N_14827,N_14707);
nand UO_1864 (O_1864,N_14961,N_14794);
or UO_1865 (O_1865,N_14829,N_14846);
nor UO_1866 (O_1866,N_14779,N_14981);
and UO_1867 (O_1867,N_14920,N_14860);
xor UO_1868 (O_1868,N_14824,N_14801);
xnor UO_1869 (O_1869,N_14709,N_14833);
nor UO_1870 (O_1870,N_14771,N_14973);
xor UO_1871 (O_1871,N_14829,N_14861);
nor UO_1872 (O_1872,N_14787,N_14853);
and UO_1873 (O_1873,N_14832,N_14923);
xnor UO_1874 (O_1874,N_14917,N_14705);
xnor UO_1875 (O_1875,N_14961,N_14990);
nor UO_1876 (O_1876,N_14974,N_14816);
or UO_1877 (O_1877,N_14927,N_14733);
nor UO_1878 (O_1878,N_14853,N_14999);
nand UO_1879 (O_1879,N_14747,N_14999);
nor UO_1880 (O_1880,N_14734,N_14915);
nor UO_1881 (O_1881,N_14899,N_14870);
xnor UO_1882 (O_1882,N_14803,N_14752);
nand UO_1883 (O_1883,N_14996,N_14878);
nand UO_1884 (O_1884,N_14970,N_14805);
and UO_1885 (O_1885,N_14738,N_14770);
or UO_1886 (O_1886,N_14786,N_14866);
nor UO_1887 (O_1887,N_14753,N_14929);
xor UO_1888 (O_1888,N_14916,N_14962);
xor UO_1889 (O_1889,N_14933,N_14873);
nand UO_1890 (O_1890,N_14793,N_14933);
nand UO_1891 (O_1891,N_14991,N_14784);
nand UO_1892 (O_1892,N_14983,N_14726);
nand UO_1893 (O_1893,N_14756,N_14733);
or UO_1894 (O_1894,N_14944,N_14763);
or UO_1895 (O_1895,N_14820,N_14980);
or UO_1896 (O_1896,N_14957,N_14887);
and UO_1897 (O_1897,N_14848,N_14743);
nand UO_1898 (O_1898,N_14894,N_14965);
nand UO_1899 (O_1899,N_14828,N_14976);
nand UO_1900 (O_1900,N_14971,N_14750);
nand UO_1901 (O_1901,N_14957,N_14830);
nor UO_1902 (O_1902,N_14753,N_14712);
xor UO_1903 (O_1903,N_14719,N_14974);
or UO_1904 (O_1904,N_14711,N_14845);
xnor UO_1905 (O_1905,N_14889,N_14893);
nor UO_1906 (O_1906,N_14816,N_14964);
nor UO_1907 (O_1907,N_14795,N_14877);
xnor UO_1908 (O_1908,N_14752,N_14827);
nand UO_1909 (O_1909,N_14956,N_14916);
and UO_1910 (O_1910,N_14913,N_14982);
nand UO_1911 (O_1911,N_14945,N_14707);
xor UO_1912 (O_1912,N_14782,N_14915);
nand UO_1913 (O_1913,N_14926,N_14914);
nor UO_1914 (O_1914,N_14937,N_14730);
or UO_1915 (O_1915,N_14819,N_14889);
and UO_1916 (O_1916,N_14951,N_14730);
or UO_1917 (O_1917,N_14835,N_14908);
nor UO_1918 (O_1918,N_14831,N_14936);
or UO_1919 (O_1919,N_14760,N_14795);
or UO_1920 (O_1920,N_14745,N_14780);
and UO_1921 (O_1921,N_14730,N_14791);
and UO_1922 (O_1922,N_14912,N_14729);
and UO_1923 (O_1923,N_14716,N_14849);
nand UO_1924 (O_1924,N_14818,N_14780);
or UO_1925 (O_1925,N_14913,N_14866);
nor UO_1926 (O_1926,N_14923,N_14764);
and UO_1927 (O_1927,N_14775,N_14898);
nand UO_1928 (O_1928,N_14797,N_14996);
or UO_1929 (O_1929,N_14960,N_14945);
and UO_1930 (O_1930,N_14719,N_14724);
and UO_1931 (O_1931,N_14868,N_14851);
nor UO_1932 (O_1932,N_14749,N_14860);
or UO_1933 (O_1933,N_14900,N_14892);
nand UO_1934 (O_1934,N_14911,N_14877);
xor UO_1935 (O_1935,N_14814,N_14971);
or UO_1936 (O_1936,N_14877,N_14910);
xor UO_1937 (O_1937,N_14939,N_14757);
xor UO_1938 (O_1938,N_14786,N_14779);
and UO_1939 (O_1939,N_14706,N_14731);
or UO_1940 (O_1940,N_14952,N_14768);
nor UO_1941 (O_1941,N_14843,N_14913);
or UO_1942 (O_1942,N_14810,N_14962);
xor UO_1943 (O_1943,N_14725,N_14767);
xor UO_1944 (O_1944,N_14831,N_14998);
nor UO_1945 (O_1945,N_14808,N_14886);
and UO_1946 (O_1946,N_14994,N_14884);
xor UO_1947 (O_1947,N_14706,N_14827);
nand UO_1948 (O_1948,N_14874,N_14983);
and UO_1949 (O_1949,N_14823,N_14755);
nor UO_1950 (O_1950,N_14892,N_14759);
or UO_1951 (O_1951,N_14896,N_14709);
and UO_1952 (O_1952,N_14859,N_14885);
nor UO_1953 (O_1953,N_14868,N_14821);
nor UO_1954 (O_1954,N_14967,N_14921);
nor UO_1955 (O_1955,N_14711,N_14739);
nor UO_1956 (O_1956,N_14918,N_14774);
or UO_1957 (O_1957,N_14731,N_14958);
and UO_1958 (O_1958,N_14731,N_14774);
and UO_1959 (O_1959,N_14894,N_14911);
or UO_1960 (O_1960,N_14706,N_14893);
nand UO_1961 (O_1961,N_14705,N_14771);
xnor UO_1962 (O_1962,N_14887,N_14803);
or UO_1963 (O_1963,N_14816,N_14759);
and UO_1964 (O_1964,N_14816,N_14873);
or UO_1965 (O_1965,N_14757,N_14915);
nand UO_1966 (O_1966,N_14728,N_14791);
or UO_1967 (O_1967,N_14868,N_14914);
nand UO_1968 (O_1968,N_14986,N_14865);
or UO_1969 (O_1969,N_14889,N_14833);
nand UO_1970 (O_1970,N_14762,N_14827);
nor UO_1971 (O_1971,N_14746,N_14863);
nor UO_1972 (O_1972,N_14974,N_14726);
or UO_1973 (O_1973,N_14854,N_14936);
nor UO_1974 (O_1974,N_14802,N_14822);
xor UO_1975 (O_1975,N_14933,N_14815);
nand UO_1976 (O_1976,N_14933,N_14900);
and UO_1977 (O_1977,N_14863,N_14807);
xor UO_1978 (O_1978,N_14820,N_14950);
and UO_1979 (O_1979,N_14945,N_14829);
nor UO_1980 (O_1980,N_14727,N_14865);
xnor UO_1981 (O_1981,N_14945,N_14751);
xor UO_1982 (O_1982,N_14748,N_14791);
and UO_1983 (O_1983,N_14770,N_14957);
nor UO_1984 (O_1984,N_14944,N_14864);
nand UO_1985 (O_1985,N_14898,N_14912);
xnor UO_1986 (O_1986,N_14836,N_14996);
and UO_1987 (O_1987,N_14825,N_14717);
nor UO_1988 (O_1988,N_14845,N_14829);
nand UO_1989 (O_1989,N_14859,N_14993);
or UO_1990 (O_1990,N_14762,N_14785);
nor UO_1991 (O_1991,N_14833,N_14959);
and UO_1992 (O_1992,N_14918,N_14993);
and UO_1993 (O_1993,N_14733,N_14803);
or UO_1994 (O_1994,N_14775,N_14889);
xor UO_1995 (O_1995,N_14924,N_14946);
or UO_1996 (O_1996,N_14719,N_14981);
or UO_1997 (O_1997,N_14792,N_14943);
xor UO_1998 (O_1998,N_14979,N_14718);
and UO_1999 (O_1999,N_14722,N_14758);
endmodule