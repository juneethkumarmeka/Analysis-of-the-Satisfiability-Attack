module basic_2500_25000_3000_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_2031,In_1931);
xnor U1 (N_1,In_1763,In_1366);
and U2 (N_2,In_1077,In_1694);
xor U3 (N_3,In_2465,In_2230);
and U4 (N_4,In_258,In_114);
or U5 (N_5,In_1497,In_2406);
and U6 (N_6,In_814,In_905);
nor U7 (N_7,In_1258,In_43);
xor U8 (N_8,In_578,In_1253);
or U9 (N_9,In_61,In_1805);
or U10 (N_10,In_348,In_416);
nor U11 (N_11,In_2264,In_443);
nand U12 (N_12,In_1057,In_609);
nand U13 (N_13,In_1768,In_1575);
nor U14 (N_14,In_132,In_699);
or U15 (N_15,In_627,In_1091);
and U16 (N_16,In_1908,In_694);
nor U17 (N_17,In_1483,In_2302);
or U18 (N_18,In_1667,In_1549);
nand U19 (N_19,In_1059,In_1925);
or U20 (N_20,In_1417,In_292);
nor U21 (N_21,In_1254,In_2038);
and U22 (N_22,In_1699,In_2351);
nor U23 (N_23,In_169,In_1580);
nand U24 (N_24,In_2016,In_1875);
and U25 (N_25,In_1297,In_150);
or U26 (N_26,In_639,In_123);
or U27 (N_27,In_1240,In_726);
or U28 (N_28,In_1716,In_580);
xor U29 (N_29,In_712,In_17);
nor U30 (N_30,In_1161,In_642);
and U31 (N_31,In_834,In_1036);
nor U32 (N_32,In_1100,In_2262);
xnor U33 (N_33,In_852,In_915);
and U34 (N_34,In_2483,In_1191);
or U35 (N_35,In_1939,In_2396);
xnor U36 (N_36,In_817,In_504);
and U37 (N_37,In_1396,In_374);
and U38 (N_38,In_619,In_953);
xor U39 (N_39,In_718,In_1369);
and U40 (N_40,In_1419,In_1511);
xnor U41 (N_41,In_1291,In_1724);
and U42 (N_42,In_349,In_1565);
nand U43 (N_43,In_1532,In_1139);
and U44 (N_44,In_955,In_625);
nor U45 (N_45,In_484,In_1268);
nand U46 (N_46,In_530,In_2208);
nand U47 (N_47,In_2300,In_1971);
and U48 (N_48,In_1202,In_154);
or U49 (N_49,In_645,In_1435);
xnor U50 (N_50,In_1309,In_2414);
nor U51 (N_51,In_2149,In_1491);
xor U52 (N_52,In_2137,In_192);
nor U53 (N_53,In_462,In_822);
nand U54 (N_54,In_1034,In_1692);
nand U55 (N_55,In_2372,In_575);
xnor U56 (N_56,In_1840,In_2460);
xnor U57 (N_57,In_554,In_856);
xnor U58 (N_58,In_785,In_1416);
nor U59 (N_59,In_350,In_1665);
nand U60 (N_60,In_608,In_2180);
and U61 (N_61,In_1022,In_1543);
or U62 (N_62,In_2075,In_1027);
xor U63 (N_63,In_1870,In_850);
or U64 (N_64,In_1195,In_2443);
nand U65 (N_65,In_1718,In_242);
nand U66 (N_66,In_1962,In_786);
and U67 (N_67,In_537,In_2403);
or U68 (N_68,In_1337,In_1661);
nand U69 (N_69,In_1074,In_1437);
nor U70 (N_70,In_2340,In_1358);
nand U71 (N_71,In_1278,In_903);
or U72 (N_72,In_1539,In_1212);
xnor U73 (N_73,In_30,In_1097);
xor U74 (N_74,In_1898,In_2266);
xor U75 (N_75,In_1720,In_2172);
nor U76 (N_76,In_1111,In_138);
xnor U77 (N_77,In_509,In_764);
nand U78 (N_78,In_859,In_2417);
or U79 (N_79,In_130,In_1573);
nand U80 (N_80,In_2468,In_1929);
xor U81 (N_81,In_961,In_2193);
nand U82 (N_82,In_2148,In_2320);
nand U83 (N_83,In_1192,In_266);
and U84 (N_84,In_1176,In_1484);
nor U85 (N_85,In_2487,In_2413);
xnor U86 (N_86,In_815,In_288);
nand U87 (N_87,In_2476,In_2190);
or U88 (N_88,In_2184,In_686);
or U89 (N_89,In_628,In_1657);
or U90 (N_90,In_1713,In_897);
nand U91 (N_91,In_2462,In_2187);
nand U92 (N_92,In_2138,In_1299);
nand U93 (N_93,In_73,In_835);
and U94 (N_94,In_552,In_2448);
xnor U95 (N_95,In_520,In_2174);
nand U96 (N_96,In_315,In_579);
or U97 (N_97,In_365,In_872);
and U98 (N_98,In_1521,In_1125);
xnor U99 (N_99,In_1852,In_26);
nor U100 (N_100,In_1408,In_665);
or U101 (N_101,In_818,In_1544);
nand U102 (N_102,In_1024,In_2065);
nor U103 (N_103,In_1385,In_2318);
or U104 (N_104,In_187,In_1230);
xor U105 (N_105,In_811,In_1554);
nor U106 (N_106,In_1640,In_2191);
nor U107 (N_107,In_803,In_260);
and U108 (N_108,In_1783,In_143);
nand U109 (N_109,In_1981,In_1888);
nand U110 (N_110,In_1514,In_1480);
and U111 (N_111,In_1945,In_1364);
nand U112 (N_112,In_377,In_368);
and U113 (N_113,In_1209,In_1885);
or U114 (N_114,In_1287,In_773);
xnor U115 (N_115,In_1179,In_1612);
nand U116 (N_116,In_2154,In_2244);
xnor U117 (N_117,In_213,In_1406);
and U118 (N_118,In_2360,In_857);
and U119 (N_119,In_866,In_1663);
or U120 (N_120,In_257,In_81);
nand U121 (N_121,In_1155,In_165);
nor U122 (N_122,In_469,In_2077);
nand U123 (N_123,In_1576,In_1819);
xnor U124 (N_124,In_152,In_1616);
xor U125 (N_125,In_201,In_538);
nor U126 (N_126,In_1154,In_740);
nand U127 (N_127,In_236,In_965);
and U128 (N_128,In_225,In_88);
or U129 (N_129,In_743,In_1158);
nor U130 (N_130,In_2247,In_1001);
and U131 (N_131,In_1114,In_2299);
or U132 (N_132,In_1577,In_1910);
or U133 (N_133,In_2181,In_1513);
nand U134 (N_134,In_1828,In_177);
nor U135 (N_135,In_505,In_1051);
nand U136 (N_136,In_1376,In_503);
nand U137 (N_137,In_1141,In_2357);
or U138 (N_138,In_1150,In_757);
xor U139 (N_139,In_1993,In_735);
nor U140 (N_140,In_2020,In_995);
xnor U141 (N_141,In_767,In_209);
nor U142 (N_142,In_780,In_2245);
xnor U143 (N_143,In_1460,In_429);
nor U144 (N_144,In_1711,In_46);
nand U145 (N_145,In_188,In_2072);
and U146 (N_146,In_704,In_2324);
or U147 (N_147,In_21,In_2341);
nand U148 (N_148,In_1181,In_1171);
or U149 (N_149,In_1293,In_620);
or U150 (N_150,In_1648,In_1106);
xnor U151 (N_151,In_1917,In_2177);
nand U152 (N_152,In_2197,In_1918);
or U153 (N_153,In_148,In_1433);
or U154 (N_154,In_1854,In_1975);
or U155 (N_155,In_705,In_147);
nand U156 (N_156,In_2293,In_697);
and U157 (N_157,In_1065,In_1619);
and U158 (N_158,In_876,In_1053);
and U159 (N_159,In_990,In_998);
or U160 (N_160,In_247,In_615);
nand U161 (N_161,In_1956,In_2046);
or U162 (N_162,In_1994,In_2285);
or U163 (N_163,In_865,In_1545);
and U164 (N_164,In_836,In_1316);
nand U165 (N_165,In_2375,In_2039);
xor U166 (N_166,In_415,In_2253);
and U167 (N_167,In_1887,In_216);
nor U168 (N_168,In_1178,In_140);
or U169 (N_169,In_2382,In_572);
xor U170 (N_170,In_1928,In_1219);
or U171 (N_171,In_1164,In_2227);
nand U172 (N_172,In_1301,In_2116);
and U173 (N_173,In_1757,In_2364);
nor U174 (N_174,In_2298,In_2472);
xor U175 (N_175,In_1121,In_729);
or U176 (N_176,In_2120,In_1120);
xnor U177 (N_177,In_1463,In_1349);
and U178 (N_178,In_1361,In_643);
or U179 (N_179,In_1478,In_2006);
nand U180 (N_180,In_1581,In_1658);
nor U181 (N_181,In_1893,In_2394);
nor U182 (N_182,In_1826,In_1168);
nand U183 (N_183,In_1441,In_1210);
xnor U184 (N_184,In_491,In_1409);
and U185 (N_185,In_678,In_2307);
xor U186 (N_186,In_119,In_1030);
and U187 (N_187,In_1182,In_2325);
nand U188 (N_188,In_2223,In_2135);
nand U189 (N_189,In_1827,In_45);
xor U190 (N_190,In_1221,In_1515);
or U191 (N_191,In_2366,In_1501);
xor U192 (N_192,In_692,In_2007);
nand U193 (N_193,In_914,In_2226);
xor U194 (N_194,In_1541,In_2454);
and U195 (N_195,In_1217,In_2453);
nor U196 (N_196,In_610,In_2117);
nand U197 (N_197,In_709,In_211);
xor U198 (N_198,In_483,In_1901);
and U199 (N_199,In_18,In_1330);
nor U200 (N_200,In_1608,In_302);
nand U201 (N_201,In_1076,In_2000);
nand U202 (N_202,In_1818,In_2150);
and U203 (N_203,In_1319,In_991);
and U204 (N_204,In_105,In_917);
or U205 (N_205,In_1339,In_2335);
nor U206 (N_206,In_1225,In_278);
nand U207 (N_207,In_796,In_1535);
and U208 (N_208,In_1811,In_561);
nand U209 (N_209,In_1353,In_2311);
nand U210 (N_210,In_2017,In_375);
nor U211 (N_211,In_1397,In_1820);
and U212 (N_212,In_373,In_1402);
and U213 (N_213,In_878,In_634);
and U214 (N_214,In_1932,In_2368);
and U215 (N_215,In_2122,In_978);
xnor U216 (N_216,In_1600,In_189);
nand U217 (N_217,In_1180,In_1428);
xnor U218 (N_218,In_284,In_401);
xnor U219 (N_219,In_751,In_376);
xnor U220 (N_220,In_184,In_1979);
and U221 (N_221,In_389,In_782);
xor U222 (N_222,In_331,In_1902);
nand U223 (N_223,In_2133,In_1907);
xor U224 (N_224,In_551,In_2012);
nor U225 (N_225,In_1427,In_1738);
and U226 (N_226,In_337,In_1183);
xnor U227 (N_227,In_6,In_765);
xor U228 (N_228,In_471,In_355);
and U229 (N_229,In_741,In_285);
xnor U230 (N_230,In_999,In_1872);
xor U231 (N_231,In_1346,In_1031);
or U232 (N_232,In_1654,In_2027);
or U233 (N_233,In_1504,In_378);
nand U234 (N_234,In_1064,In_2260);
and U235 (N_235,In_1571,In_1160);
and U236 (N_236,In_414,In_1933);
nand U237 (N_237,In_1630,In_598);
nor U238 (N_238,In_2370,In_84);
or U239 (N_239,In_1715,In_393);
and U240 (N_240,In_1609,In_958);
nand U241 (N_241,In_1567,In_771);
and U242 (N_242,In_2447,In_1257);
and U243 (N_243,In_316,In_1126);
nor U244 (N_244,In_988,In_1794);
or U245 (N_245,In_1598,In_1578);
and U246 (N_246,In_333,In_403);
nand U247 (N_247,In_759,In_997);
nor U248 (N_248,In_2048,In_727);
nor U249 (N_249,In_425,In_809);
nor U250 (N_250,In_534,In_638);
nor U251 (N_251,In_219,In_166);
xor U252 (N_252,In_508,In_117);
nand U253 (N_253,In_1216,In_2319);
nor U254 (N_254,In_1863,In_755);
and U255 (N_255,In_203,In_1599);
nand U256 (N_256,In_1015,In_0);
nor U257 (N_257,In_1333,In_2182);
xnor U258 (N_258,In_2478,In_480);
xor U259 (N_259,In_77,In_1508);
or U260 (N_260,In_1582,In_227);
nand U261 (N_261,In_833,In_523);
nor U262 (N_262,In_2052,In_879);
nand U263 (N_263,In_394,In_684);
nand U264 (N_264,In_200,In_89);
and U265 (N_265,In_2222,In_1320);
nand U266 (N_266,In_870,In_1823);
xor U267 (N_267,In_513,In_2159);
or U268 (N_268,In_338,In_2346);
xor U269 (N_269,In_2390,In_1285);
or U270 (N_270,In_1815,In_2189);
xnor U271 (N_271,In_1006,In_2466);
or U272 (N_272,In_1991,In_1013);
or U273 (N_273,In_664,In_1996);
nor U274 (N_274,In_1373,In_1528);
and U275 (N_275,In_395,In_369);
or U276 (N_276,In_2369,In_234);
nor U277 (N_277,In_701,In_1213);
or U278 (N_278,In_889,In_2494);
or U279 (N_279,In_439,In_1947);
nand U280 (N_280,In_1453,In_1270);
nor U281 (N_281,In_2326,In_2014);
nor U282 (N_282,In_823,In_456);
nand U283 (N_283,In_1159,In_1882);
nor U284 (N_284,In_44,In_929);
nand U285 (N_285,In_969,In_734);
nor U286 (N_286,In_599,In_992);
and U287 (N_287,In_2332,In_1223);
nand U288 (N_288,In_1686,In_1042);
xor U289 (N_289,In_2336,In_1703);
xnor U290 (N_290,In_1843,In_2037);
or U291 (N_291,In_1556,In_2115);
xnor U292 (N_292,In_2240,In_58);
nor U293 (N_293,In_565,In_1890);
nor U294 (N_294,In_685,In_1915);
or U295 (N_295,In_550,In_1835);
or U296 (N_296,In_498,In_840);
xnor U297 (N_297,In_248,In_1510);
nand U298 (N_298,In_2458,In_1211);
nor U299 (N_299,In_194,In_595);
nor U300 (N_300,In_2395,In_968);
xor U301 (N_301,In_1551,In_637);
xnor U302 (N_302,In_967,In_566);
nor U303 (N_303,In_2186,In_175);
nor U304 (N_304,In_526,In_1698);
nand U305 (N_305,In_2282,In_1842);
and U306 (N_306,In_1856,In_475);
nand U307 (N_307,In_1967,In_93);
and U308 (N_308,In_1802,In_2459);
xor U309 (N_309,In_1526,In_358);
nand U310 (N_310,In_490,In_1533);
nand U311 (N_311,In_1371,In_111);
nor U312 (N_312,In_2444,In_1186);
and U313 (N_313,In_753,In_2078);
xor U314 (N_314,In_1680,In_576);
nor U315 (N_315,In_2477,In_482);
or U316 (N_316,In_654,In_2042);
and U317 (N_317,In_1531,In_1924);
and U318 (N_318,In_1520,In_67);
nand U319 (N_319,In_1712,In_2207);
and U320 (N_320,In_533,In_1267);
or U321 (N_321,In_214,In_1974);
nand U322 (N_322,In_1555,In_1804);
and U323 (N_323,In_212,In_819);
nand U324 (N_324,In_2463,In_182);
and U325 (N_325,In_80,In_2158);
and U326 (N_326,In_1462,In_923);
and U327 (N_327,In_1756,In_162);
nor U328 (N_328,In_2358,In_445);
and U329 (N_329,In_1392,In_1662);
and U330 (N_330,In_2473,In_2424);
nor U331 (N_331,In_1399,In_145);
or U332 (N_332,In_1099,In_2092);
xnor U333 (N_333,In_1790,In_2131);
and U334 (N_334,In_1771,In_573);
and U335 (N_335,In_336,In_1821);
and U336 (N_336,In_1921,In_2114);
nand U337 (N_337,In_1930,In_2126);
xnor U338 (N_338,In_459,In_1318);
nand U339 (N_339,In_1518,In_2391);
xnor U340 (N_340,In_1973,In_1629);
nand U341 (N_341,In_56,In_1425);
and U342 (N_342,In_524,In_1559);
nand U343 (N_343,In_806,In_742);
xor U344 (N_344,In_632,In_1023);
or U345 (N_345,In_408,In_2152);
and U346 (N_346,In_66,In_1475);
or U347 (N_347,In_1454,In_2350);
xnor U348 (N_348,In_2015,In_564);
xnor U349 (N_349,In_2164,In_1675);
xnor U350 (N_350,In_2231,In_2429);
nand U351 (N_351,In_205,In_1553);
xnor U352 (N_352,In_1199,In_2384);
and U353 (N_353,In_1292,In_398);
xnor U354 (N_354,In_2322,In_962);
nor U355 (N_355,In_920,In_2328);
xnor U356 (N_356,In_825,In_1999);
xnor U357 (N_357,In_185,In_412);
nor U358 (N_358,In_563,In_805);
nor U359 (N_359,In_949,In_1156);
nor U360 (N_360,In_2291,In_1748);
nor U361 (N_361,In_1701,In_1853);
or U362 (N_362,In_659,In_1761);
nand U363 (N_363,In_1540,In_1274);
or U364 (N_364,In_383,In_529);
nor U365 (N_365,In_243,In_458);
nand U366 (N_366,In_1688,In_1446);
or U367 (N_367,In_52,In_324);
nor U368 (N_368,In_1145,In_783);
xor U369 (N_369,In_1208,In_1807);
and U370 (N_370,In_1415,In_474);
and U371 (N_371,In_1868,In_190);
nor U372 (N_372,In_2030,In_2107);
nor U373 (N_373,In_1537,In_467);
or U374 (N_374,In_586,In_1205);
nor U375 (N_375,In_1775,In_364);
and U376 (N_376,In_594,In_1758);
nand U377 (N_377,In_2044,In_1218);
nand U378 (N_378,In_669,In_255);
nand U379 (N_379,In_952,In_226);
and U380 (N_380,In_1886,In_1423);
and U381 (N_381,In_1911,In_1836);
and U382 (N_382,In_1940,In_1388);
or U383 (N_383,In_2228,In_1845);
and U384 (N_384,In_347,In_356);
nor U385 (N_385,In_1079,In_1259);
xor U386 (N_386,In_286,In_821);
nor U387 (N_387,In_340,In_2130);
and U388 (N_388,In_2229,In_275);
nor U389 (N_389,In_882,In_1017);
and U390 (N_390,In_2067,In_1639);
xnor U391 (N_391,In_1604,In_1379);
nor U392 (N_392,In_845,In_1594);
and U393 (N_393,In_1770,In_2495);
nand U394 (N_394,In_984,In_1652);
xnor U395 (N_395,In_1586,In_1904);
nand U396 (N_396,In_134,In_940);
or U397 (N_397,In_2111,In_623);
nand U398 (N_398,In_1755,In_362);
nor U399 (N_399,In_1774,In_671);
nand U400 (N_400,In_1874,In_2216);
nand U401 (N_401,In_2345,In_388);
xnor U402 (N_402,In_320,In_1547);
or U403 (N_403,In_1951,In_109);
and U404 (N_404,In_1260,In_2026);
or U405 (N_405,In_1982,In_100);
nand U406 (N_406,In_2296,In_1903);
nor U407 (N_407,In_37,In_2087);
xor U408 (N_408,In_1054,In_676);
xor U409 (N_409,In_1892,In_313);
xor U410 (N_410,In_933,In_1632);
xnor U411 (N_411,In_5,In_3);
or U412 (N_412,In_271,In_1250);
or U413 (N_413,In_2308,In_883);
xor U414 (N_414,In_1328,In_1080);
or U415 (N_415,In_353,In_94);
or U416 (N_416,In_1193,In_1283);
nor U417 (N_417,In_1793,In_1081);
xor U418 (N_418,In_402,In_863);
or U419 (N_419,In_2125,In_2110);
nand U420 (N_420,In_82,In_2408);
xor U421 (N_421,In_979,In_256);
or U422 (N_422,In_312,In_1039);
and U423 (N_423,In_157,In_848);
nor U424 (N_424,In_1009,In_2010);
or U425 (N_425,In_1372,In_107);
xnor U426 (N_426,In_1447,In_179);
xnor U427 (N_427,In_249,In_380);
or U428 (N_428,In_1461,In_946);
and U429 (N_429,In_435,In_1367);
or U430 (N_430,In_1857,In_1083);
nor U431 (N_431,In_1127,In_1782);
nand U432 (N_432,In_1044,In_1912);
nor U433 (N_433,In_1666,In_2023);
xnor U434 (N_434,In_716,In_2410);
and U435 (N_435,In_1313,In_1627);
nand U436 (N_436,In_1336,In_2456);
nor U437 (N_437,In_1374,In_2201);
xnor U438 (N_438,In_1492,In_1509);
or U439 (N_439,In_749,In_1846);
nor U440 (N_440,In_2002,In_877);
and U441 (N_441,In_862,In_1233);
nor U442 (N_442,In_421,In_2203);
and U443 (N_443,In_2101,In_2198);
xnor U444 (N_444,In_2062,In_1140);
xnor U445 (N_445,In_2166,In_1273);
nand U446 (N_446,In_2086,In_1272);
and U447 (N_447,In_706,In_2090);
nor U448 (N_448,In_1220,In_1781);
and U449 (N_449,In_163,In_2081);
nand U450 (N_450,In_2128,In_1421);
xor U451 (N_451,In_1759,In_186);
or U452 (N_452,In_486,In_305);
nand U453 (N_453,In_2428,In_1558);
or U454 (N_454,In_1844,In_2430);
or U455 (N_455,In_541,In_924);
nor U456 (N_456,In_481,In_1832);
xor U457 (N_457,In_2259,In_1308);
nand U458 (N_458,In_2267,In_2276);
or U459 (N_459,In_1245,In_2373);
or U460 (N_460,In_2132,In_277);
and U461 (N_461,In_1621,In_1574);
and U462 (N_462,In_2224,In_1198);
xor U463 (N_463,In_858,In_1611);
and U464 (N_464,In_789,In_2277);
or U465 (N_465,In_352,In_1082);
and U466 (N_466,In_4,In_2013);
xor U467 (N_467,In_521,In_2338);
or U468 (N_468,In_2292,In_1296);
nor U469 (N_469,In_1187,In_233);
xnor U470 (N_470,In_1517,In_2035);
and U471 (N_471,In_2297,In_174);
xor U472 (N_472,In_14,In_2251);
xor U473 (N_473,In_15,In_1597);
xor U474 (N_474,In_567,In_1305);
xnor U475 (N_475,In_571,In_1086);
or U476 (N_476,In_1167,In_1038);
xnor U477 (N_477,In_2422,In_2210);
nor U478 (N_478,In_793,In_1847);
nor U479 (N_479,In_2213,In_631);
nand U480 (N_480,In_1324,In_2426);
nor U481 (N_481,In_1734,In_2496);
nand U482 (N_482,In_2236,In_2353);
and U483 (N_483,In_1949,In_569);
or U484 (N_484,In_149,In_230);
and U485 (N_485,In_2237,In_1656);
nor U486 (N_486,In_1375,In_1331);
or U487 (N_487,In_2365,In_74);
and U488 (N_488,In_2275,In_500);
xor U489 (N_489,In_193,In_2082);
and U490 (N_490,In_1746,In_522);
and U491 (N_491,In_1413,In_2470);
nor U492 (N_492,In_2220,In_2356);
nand U493 (N_493,In_2480,In_54);
nand U494 (N_494,In_50,In_2045);
xnor U495 (N_495,In_423,In_1527);
and U496 (N_496,In_853,In_2270);
xnor U497 (N_497,In_540,In_1112);
and U498 (N_498,In_510,In_1380);
nand U499 (N_499,In_1426,In_994);
nor U500 (N_500,In_1060,In_2219);
xor U501 (N_501,In_1306,In_913);
or U502 (N_502,In_1116,N_98);
and U503 (N_503,N_385,In_2074);
nand U504 (N_504,In_115,In_38);
or U505 (N_505,In_2112,In_2310);
and U506 (N_506,In_1063,In_495);
nor U507 (N_507,In_2339,In_23);
nor U508 (N_508,In_159,In_1614);
and U509 (N_509,In_535,In_2446);
and U510 (N_510,In_1118,In_1286);
and U511 (N_511,In_1624,In_974);
or U512 (N_512,In_2147,In_795);
and U513 (N_513,In_34,In_907);
xnor U514 (N_514,N_196,In_1153);
or U515 (N_515,In_1977,In_2412);
or U516 (N_516,In_2175,In_732);
and U517 (N_517,N_253,In_2151);
and U518 (N_518,In_1025,In_553);
nand U519 (N_519,N_244,In_2497);
xor U520 (N_520,N_313,In_860);
nand U521 (N_521,In_1449,In_947);
and U522 (N_522,In_900,In_744);
xnor U523 (N_523,N_458,In_2162);
or U524 (N_524,In_601,In_1310);
nor U525 (N_525,In_2136,In_2153);
and U526 (N_526,N_318,In_2441);
nor U527 (N_527,In_1980,In_600);
nor U528 (N_528,In_750,In_2008);
and U529 (N_529,In_261,In_2286);
and U530 (N_530,In_2314,In_1148);
nand U531 (N_531,In_407,In_826);
xor U532 (N_532,In_2032,N_406);
xor U533 (N_533,In_1839,In_202);
or U534 (N_534,In_1429,In_1834);
nor U535 (N_535,In_2239,In_1669);
or U536 (N_536,In_392,N_413);
and U537 (N_537,In_1288,In_1860);
nor U538 (N_538,In_1569,N_420);
nand U539 (N_539,In_762,In_1329);
or U540 (N_540,N_287,In_1867);
or U541 (N_541,In_2387,N_445);
and U542 (N_542,In_1020,In_1725);
nor U543 (N_543,In_1264,In_720);
and U544 (N_544,In_1452,In_930);
nand U545 (N_545,In_2232,In_1029);
xor U546 (N_546,In_2071,In_335);
nor U547 (N_547,In_1239,In_2388);
nand U548 (N_548,N_147,In_367);
or U549 (N_549,In_956,In_2057);
nand U550 (N_550,In_1709,In_327);
xnor U551 (N_551,N_278,In_164);
xnor U552 (N_552,In_779,In_919);
xnor U553 (N_553,In_1056,N_250);
and U554 (N_554,In_2011,N_47);
or U555 (N_555,In_2344,In_178);
or U556 (N_556,In_454,In_2452);
nand U557 (N_557,N_210,N_56);
xor U558 (N_558,N_324,In_950);
xor U559 (N_559,In_1978,In_1613);
nand U560 (N_560,In_584,In_1678);
xnor U561 (N_561,In_1953,In_746);
nor U562 (N_562,N_399,N_32);
xor U563 (N_563,In_2022,In_1849);
and U564 (N_564,In_1344,In_1937);
xnor U565 (N_565,In_1637,In_1157);
nor U566 (N_566,In_1078,In_1377);
and U567 (N_567,In_363,In_299);
xnor U568 (N_568,In_422,In_1055);
nand U569 (N_569,In_1494,In_791);
nand U570 (N_570,In_1105,N_100);
xor U571 (N_571,In_1585,N_168);
nand U572 (N_572,In_1728,In_1830);
nor U573 (N_573,N_251,In_518);
xnor U574 (N_574,N_184,In_1398);
or U575 (N_575,In_1457,In_804);
nand U576 (N_576,In_989,In_1049);
xnor U577 (N_577,In_1583,In_2156);
or U578 (N_578,In_724,In_568);
nand U579 (N_579,In_1045,N_54);
xnor U580 (N_580,In_1751,N_224);
or U581 (N_581,N_109,N_165);
and U582 (N_582,In_1298,In_1866);
and U583 (N_583,In_1184,N_188);
nor U584 (N_584,In_411,In_515);
xor U585 (N_585,N_6,N_421);
or U586 (N_586,N_134,In_675);
nor U587 (N_587,In_64,N_387);
nand U588 (N_588,In_1073,N_59);
xnor U589 (N_589,In_91,N_190);
xnor U590 (N_590,In_1891,In_2363);
nor U591 (N_591,N_396,In_797);
or U592 (N_592,N_308,In_1797);
or U593 (N_593,N_229,N_16);
or U594 (N_594,In_1955,In_1691);
nand U595 (N_595,N_439,In_270);
nor U596 (N_596,In_2157,In_379);
nand U597 (N_597,N_246,In_673);
nand U598 (N_598,In_2437,N_279);
and U599 (N_599,N_178,In_1177);
nor U600 (N_600,N_414,In_1618);
or U601 (N_601,N_207,In_1880);
or U602 (N_602,In_1922,In_936);
or U603 (N_603,N_271,In_813);
nor U604 (N_604,In_916,In_2254);
or U605 (N_605,In_2398,N_444);
or U606 (N_606,In_2315,In_559);
nand U607 (N_607,In_2405,In_1222);
nor U608 (N_608,In_941,In_1169);
nor U609 (N_609,In_776,N_35);
nor U610 (N_610,In_622,N_434);
and U611 (N_611,In_381,In_733);
nand U612 (N_612,In_1799,N_284);
nor U613 (N_613,In_1143,In_1207);
or U614 (N_614,In_1767,In_2379);
xnor U615 (N_615,In_1269,In_1473);
nand U616 (N_616,In_1271,N_494);
and U617 (N_617,N_297,In_2376);
xnor U618 (N_618,In_2273,N_163);
xor U619 (N_619,In_2475,In_330);
nand U620 (N_620,N_50,In_1448);
nor U621 (N_621,In_2290,In_650);
xor U622 (N_622,In_2389,N_53);
or U623 (N_623,In_36,In_1058);
xor U624 (N_624,In_2248,In_1312);
xnor U625 (N_625,N_101,In_1393);
and U626 (N_626,N_368,In_618);
xor U627 (N_627,N_311,N_298);
xnor U628 (N_628,N_227,In_1280);
and U629 (N_629,In_332,In_1670);
nand U630 (N_630,In_868,In_106);
and U631 (N_631,In_648,In_1684);
xnor U632 (N_632,In_1228,N_67);
nand U633 (N_633,N_152,In_1390);
nor U634 (N_634,N_180,In_293);
xor U635 (N_635,In_1395,In_204);
nand U636 (N_636,N_3,In_721);
xnor U637 (N_637,N_263,N_283);
xor U638 (N_638,N_148,In_167);
and U639 (N_639,N_247,In_1693);
xnor U640 (N_640,N_202,N_374);
xnor U641 (N_641,In_644,In_766);
or U642 (N_642,In_1340,In_925);
xnor U643 (N_643,In_306,N_329);
or U644 (N_644,N_348,In_1455);
nand U645 (N_645,In_62,In_69);
nor U646 (N_646,In_772,In_1307);
and U647 (N_647,N_415,In_1474);
and U648 (N_648,In_2,In_1162);
and U649 (N_649,In_1704,In_1719);
nor U650 (N_650,In_492,N_17);
and U651 (N_651,In_139,In_2185);
and U652 (N_652,In_661,In_31);
nand U653 (N_653,In_715,In_1944);
or U654 (N_654,In_314,In_1489);
and U655 (N_655,N_293,In_1387);
or U656 (N_656,In_611,In_1403);
and U657 (N_657,In_1562,In_581);
nor U658 (N_658,In_450,In_1735);
or U659 (N_659,In_341,In_273);
nor U660 (N_660,In_2421,In_343);
nand U661 (N_661,In_1708,N_309);
xor U662 (N_662,N_235,N_462);
nor U663 (N_663,In_251,In_898);
or U664 (N_664,In_1424,In_235);
nand U665 (N_665,In_2295,In_1351);
and U666 (N_666,In_2342,In_1072);
xnor U667 (N_667,N_485,In_2113);
and U668 (N_668,In_1859,In_1314);
and U669 (N_669,N_409,In_397);
xnor U670 (N_670,In_2402,In_2305);
xnor U671 (N_671,In_1443,N_482);
nand U672 (N_672,N_392,N_496);
xor U673 (N_673,In_1035,In_210);
or U674 (N_674,N_424,In_406);
and U675 (N_675,In_263,N_130);
and U676 (N_676,In_191,In_635);
nor U677 (N_677,In_63,In_1899);
and U678 (N_678,In_1721,N_110);
nor U679 (N_679,In_1765,In_1163);
nand U680 (N_680,In_1342,In_479);
or U681 (N_681,In_339,In_921);
and U682 (N_682,N_52,In_507);
nand U683 (N_683,In_501,In_1108);
nand U684 (N_684,In_2055,In_2347);
xor U685 (N_685,In_60,N_355);
xnor U686 (N_686,In_1092,In_1479);
and U687 (N_687,N_39,In_1332);
xor U688 (N_688,In_1381,In_2274);
nor U689 (N_689,In_16,In_301);
nor U690 (N_690,N_144,In_2461);
nand U691 (N_691,In_1838,In_1414);
xor U692 (N_692,In_1696,In_1625);
nor U693 (N_693,N_490,N_177);
nand U694 (N_694,N_401,In_1095);
xor U695 (N_695,In_2019,In_1589);
or U696 (N_696,In_497,In_156);
or U697 (N_697,N_218,N_89);
and U698 (N_698,In_1606,In_792);
nand U699 (N_699,N_254,In_1946);
nand U700 (N_700,In_624,In_334);
nand U701 (N_701,In_1800,In_1777);
and U702 (N_702,In_1041,N_143);
and U703 (N_703,N_149,In_1747);
xor U704 (N_704,N_95,In_1175);
nor U705 (N_705,In_574,In_2214);
or U706 (N_706,N_469,In_778);
or U707 (N_707,In_1674,In_2140);
xor U708 (N_708,In_254,In_931);
nand U709 (N_709,In_874,In_72);
nor U710 (N_710,In_2058,N_172);
nand U711 (N_711,In_660,In_1502);
and U712 (N_712,In_980,N_212);
and U713 (N_713,In_472,In_1523);
nand U714 (N_714,N_70,In_1740);
xor U715 (N_715,N_301,N_214);
nand U716 (N_716,In_2047,In_2380);
or U717 (N_717,In_707,In_649);
nand U718 (N_718,In_1593,In_1394);
nor U719 (N_719,In_2036,In_2362);
and U720 (N_720,In_71,In_1026);
nor U721 (N_721,N_103,In_433);
or U722 (N_722,In_2085,N_226);
nor U723 (N_723,N_60,In_926);
nor U724 (N_724,In_1007,N_383);
nand U725 (N_725,In_1610,In_99);
xnor U726 (N_726,N_363,N_450);
or U727 (N_727,N_8,N_335);
nand U728 (N_728,In_1516,In_1004);
or U729 (N_729,In_2105,In_641);
nor U730 (N_730,N_398,In_2123);
and U731 (N_731,N_466,N_461);
xnor U732 (N_732,N_68,In_1697);
nor U733 (N_733,In_1304,In_1788);
and U734 (N_734,In_1507,In_2221);
nand U735 (N_735,In_1655,In_688);
xor U736 (N_736,N_146,N_82);
xnor U737 (N_737,In_222,In_1386);
xnor U738 (N_738,N_18,In_1472);
and U739 (N_739,In_437,N_225);
and U740 (N_740,In_674,N_2);
nand U741 (N_741,N_171,In_40);
xnor U742 (N_742,In_713,N_328);
nand U743 (N_743,In_837,In_652);
nand U744 (N_744,In_430,In_180);
and U745 (N_745,In_1634,In_1347);
xnor U746 (N_746,In_2200,In_2076);
xor U747 (N_747,In_512,N_314);
nand U748 (N_748,In_1151,In_1110);
and U749 (N_749,N_487,In_1215);
nor U750 (N_750,In_2215,N_416);
nand U751 (N_751,In_2194,N_12);
nand U752 (N_752,In_323,N_258);
or U753 (N_753,In_1732,In_442);
nor U754 (N_754,In_945,In_1101);
or U755 (N_755,In_1934,In_1439);
nor U756 (N_756,In_1241,In_2225);
nor U757 (N_757,In_1871,In_722);
nand U758 (N_758,N_372,In_1354);
xnor U759 (N_759,In_1753,In_973);
and U760 (N_760,N_169,In_228);
nand U761 (N_761,N_333,In_28);
xor U762 (N_762,In_1075,In_122);
xor U763 (N_763,In_2033,In_2066);
or U764 (N_764,In_446,In_1672);
or U765 (N_765,In_557,N_274);
xnor U766 (N_766,In_1173,N_288);
nor U767 (N_767,N_23,In_2009);
nand U768 (N_768,N_366,N_265);
and U769 (N_769,N_200,N_0);
nor U770 (N_770,N_108,In_2018);
nand U771 (N_771,N_24,In_2329);
and U772 (N_772,In_1764,In_2060);
and U773 (N_773,In_128,In_399);
nand U774 (N_774,In_1277,N_339);
and U775 (N_775,In_1679,In_27);
or U776 (N_776,In_2409,In_1986);
and U777 (N_777,In_268,In_626);
or U778 (N_778,In_1477,In_1348);
or U779 (N_779,In_1128,In_1563);
xnor U780 (N_780,N_262,In_413);
nor U781 (N_781,In_2281,In_1522);
and U782 (N_782,In_2348,In_1923);
nand U783 (N_783,N_121,In_39);
and U784 (N_784,In_1229,In_820);
xor U785 (N_785,In_975,N_97);
xnor U786 (N_786,In_2284,In_146);
nand U787 (N_787,In_2261,In_1206);
xor U788 (N_788,N_491,In_1458);
and U789 (N_789,In_2349,N_369);
and U790 (N_790,In_274,In_781);
or U791 (N_791,In_830,In_2196);
or U792 (N_792,N_111,In_514);
and U793 (N_793,N_493,In_1459);
or U794 (N_794,In_2257,In_220);
nor U795 (N_795,In_96,In_2474);
nor U796 (N_796,In_253,In_2059);
xnor U797 (N_797,N_437,In_1638);
or U798 (N_798,In_400,N_158);
nor U799 (N_799,In_463,In_1360);
xor U800 (N_800,In_259,In_1984);
nand U801 (N_801,In_2491,In_2490);
nor U802 (N_802,In_280,N_189);
nand U803 (N_803,In_1247,In_1102);
nor U804 (N_804,In_2371,In_802);
xnor U805 (N_805,N_456,In_1650);
and U806 (N_806,In_125,In_2435);
and U807 (N_807,In_1295,In_1189);
and U808 (N_808,In_1043,In_1005);
nand U809 (N_809,N_78,In_11);
and U810 (N_810,In_92,In_502);
nand U811 (N_811,In_1776,In_1248);
nand U812 (N_812,In_583,In_307);
and U813 (N_813,In_1300,In_887);
nor U814 (N_814,N_371,In_1113);
and U815 (N_815,In_354,N_483);
nand U816 (N_816,In_893,In_544);
xor U817 (N_817,In_668,In_1190);
or U818 (N_818,N_411,In_1);
nand U819 (N_819,N_80,N_62);
and U820 (N_820,In_1862,In_777);
nand U821 (N_821,N_484,In_517);
nor U822 (N_822,In_176,In_2381);
or U823 (N_823,In_95,In_1519);
nor U824 (N_824,In_97,In_1837);
and U825 (N_825,In_310,In_1263);
nand U826 (N_826,In_799,In_2094);
or U827 (N_827,In_1410,In_131);
or U828 (N_828,In_1290,In_703);
xnor U829 (N_829,In_1542,In_1687);
nand U830 (N_830,In_417,In_181);
nor U831 (N_831,In_2004,In_141);
xnor U832 (N_832,In_912,In_1950);
and U833 (N_833,In_2212,N_248);
and U834 (N_834,In_1482,In_1965);
or U835 (N_835,In_221,N_216);
and U836 (N_836,In_922,In_1959);
xnor U837 (N_837,In_647,N_129);
xnor U838 (N_838,In_151,N_289);
nor U839 (N_839,In_2420,N_429);
or U840 (N_840,In_1016,In_2051);
nor U841 (N_841,In_590,In_1032);
and U842 (N_842,In_1972,In_1564);
or U843 (N_843,N_266,In_465);
nor U844 (N_844,In_754,In_1942);
xnor U845 (N_845,N_362,N_359);
and U846 (N_846,In_1677,In_404);
and U847 (N_847,In_1400,In_1165);
nor U848 (N_848,In_1752,N_19);
nor U849 (N_849,In_985,In_2183);
and U850 (N_850,In_1588,In_133);
nand U851 (N_851,In_2139,In_577);
nand U852 (N_852,In_2165,In_880);
nand U853 (N_853,In_982,In_1014);
xor U854 (N_854,In_1881,In_1570);
or U855 (N_855,In_1355,In_1235);
nand U856 (N_856,In_102,In_525);
xor U857 (N_857,In_1084,In_1960);
and U858 (N_858,In_869,In_851);
nand U859 (N_859,N_305,In_2492);
xor U860 (N_860,In_670,In_981);
nand U861 (N_861,In_1913,In_2049);
or U862 (N_862,In_431,N_454);
or U863 (N_863,In_485,N_164);
and U864 (N_864,N_125,In_432);
nand U865 (N_865,N_81,In_562);
xor U866 (N_866,N_22,In_2097);
nor U867 (N_867,In_1089,In_1315);
or U868 (N_868,In_774,N_217);
xor U869 (N_869,In_2287,N_455);
or U870 (N_870,In_1450,In_1591);
or U871 (N_871,In_1200,In_1172);
nand U872 (N_872,In_1098,In_195);
nand U873 (N_873,In_901,In_2054);
xnor U874 (N_874,N_33,In_424);
xnor U875 (N_875,In_1958,In_127);
and U876 (N_876,In_2029,N_418);
nand U877 (N_877,In_2499,In_2471);
or U878 (N_878,In_731,In_2070);
nand U879 (N_879,In_1546,In_2401);
nor U880 (N_880,In_1040,N_84);
and U881 (N_881,In_1048,In_2238);
nand U882 (N_882,In_2312,In_745);
xnor U883 (N_883,In_2258,In_1088);
nor U884 (N_884,In_1008,In_229);
and U885 (N_885,N_426,In_1345);
nand U886 (N_886,In_885,In_75);
nor U887 (N_887,N_28,In_738);
xor U888 (N_888,N_476,N_221);
and U889 (N_889,In_2204,In_1281);
nor U890 (N_890,In_112,In_325);
nor U891 (N_891,N_187,N_112);
xnor U892 (N_892,In_1916,In_1552);
nor U893 (N_893,In_1762,In_290);
xnor U894 (N_894,N_365,In_1493);
nor U895 (N_895,In_653,In_2205);
xnor U896 (N_896,In_1096,In_928);
xor U897 (N_897,In_2093,In_2330);
xor U898 (N_898,In_2278,In_1906);
or U899 (N_899,In_279,In_683);
and U900 (N_900,N_243,N_162);
and U901 (N_901,In_1249,In_291);
nor U902 (N_902,N_393,In_1224);
or U903 (N_903,In_344,N_435);
and U904 (N_904,In_51,In_309);
xnor U905 (N_905,In_1188,In_1969);
xor U906 (N_906,N_277,N_304);
nand U907 (N_907,N_38,N_478);
and U908 (N_908,In_328,N_122);
nand U909 (N_909,N_272,In_2028);
nor U910 (N_910,In_1276,N_459);
nor U911 (N_911,In_593,In_262);
or U912 (N_912,In_1990,N_432);
nor U913 (N_913,In_1261,N_131);
and U914 (N_914,In_633,In_451);
nand U915 (N_915,In_1237,In_2451);
nand U916 (N_916,In_2146,N_477);
nor U917 (N_917,In_847,N_428);
or U918 (N_918,In_1119,In_2119);
and U919 (N_919,In_493,In_2053);
or U920 (N_920,In_614,N_181);
or U921 (N_921,In_2343,In_1723);
and U922 (N_922,In_2450,In_1359);
xor U923 (N_923,In_2241,N_449);
xnor U924 (N_924,In_1796,In_1592);
and U925 (N_925,N_140,In_1370);
nand U926 (N_926,N_9,N_440);
nor U927 (N_927,N_15,N_102);
nor U928 (N_928,N_238,In_828);
or U929 (N_929,In_596,In_1737);
xnor U930 (N_930,In_1935,In_494);
or U931 (N_931,In_937,In_2327);
xor U932 (N_932,In_680,In_1879);
xor U933 (N_933,N_280,In_2352);
and U934 (N_934,In_1850,In_768);
or U935 (N_935,In_2378,In_536);
nor U936 (N_936,In_1742,In_1470);
nand U937 (N_937,In_265,In_1232);
nor U938 (N_938,N_72,N_473);
nand U939 (N_939,In_658,In_1702);
xnor U940 (N_940,In_758,In_1787);
nand U941 (N_941,In_473,N_452);
or U942 (N_942,In_1631,In_2404);
xor U943 (N_943,In_1196,In_1087);
xor U944 (N_944,In_1919,In_208);
and U945 (N_945,N_380,In_1144);
nor U946 (N_946,N_256,N_317);
or U947 (N_947,In_440,In_2337);
or U948 (N_948,N_475,In_543);
or U949 (N_949,In_2289,In_104);
and U950 (N_950,In_390,In_2323);
or U951 (N_951,In_2355,In_1524);
or U952 (N_952,In_1068,In_886);
nor U953 (N_953,In_1660,In_2168);
nand U954 (N_954,In_2280,In_1129);
and U955 (N_955,In_304,In_906);
xor U956 (N_956,In_405,N_378);
nand U957 (N_957,In_2025,In_32);
and U958 (N_958,In_651,In_1561);
xnor U959 (N_959,N_124,In_250);
and U960 (N_960,In_155,In_1590);
xnor U961 (N_961,In_1214,In_1486);
nor U962 (N_962,In_2098,In_47);
nand U963 (N_963,N_457,In_531);
and U964 (N_964,In_2061,In_996);
xor U965 (N_965,In_1047,In_2269);
and U966 (N_966,In_963,In_2109);
xnor U967 (N_967,In_844,In_2195);
nor U968 (N_968,In_656,N_352);
or U969 (N_969,In_1676,In_1343);
xor U970 (N_970,In_873,N_211);
nor U971 (N_971,In_849,In_2246);
or U972 (N_972,In_1322,In_370);
or U973 (N_973,In_1383,In_391);
xor U974 (N_974,N_106,In_1896);
nand U975 (N_975,In_2317,In_2173);
xnor U976 (N_976,In_1467,In_1998);
xnor U977 (N_977,N_389,In_496);
and U978 (N_978,In_532,In_558);
and U979 (N_979,In_1779,N_268);
and U980 (N_980,In_951,N_240);
xor U981 (N_981,N_45,N_360);
xor U982 (N_982,In_1107,N_36);
xnor U983 (N_983,In_1620,In_719);
nand U984 (N_984,In_1773,In_1873);
and U985 (N_985,N_282,In_1130);
and U986 (N_986,In_827,In_1067);
nor U987 (N_987,In_161,In_282);
xnor U988 (N_988,In_824,N_322);
or U989 (N_989,In_747,In_841);
nand U990 (N_990,N_136,In_1341);
nand U991 (N_991,In_1861,In_2043);
xnor U992 (N_992,N_74,In_1431);
nand U993 (N_993,In_1989,In_477);
or U994 (N_994,N_57,In_1816);
xor U995 (N_995,In_570,N_296);
and U996 (N_996,In_918,In_603);
and U997 (N_997,In_1943,N_257);
nor U998 (N_998,In_2235,In_606);
and U999 (N_999,In_2118,In_2488);
and U1000 (N_1000,In_65,In_1530);
and U1001 (N_1001,N_443,N_940);
xor U1002 (N_1002,N_123,N_572);
xor U1003 (N_1003,N_744,N_321);
and U1004 (N_1004,In_2439,N_818);
nand U1005 (N_1005,N_793,In_1936);
xor U1006 (N_1006,In_2445,N_633);
xor U1007 (N_1007,In_217,In_1066);
nand U1008 (N_1008,N_986,In_1749);
and U1009 (N_1009,N_590,N_132);
xnor U1010 (N_1010,N_319,N_906);
xnor U1011 (N_1011,N_453,N_777);
xor U1012 (N_1012,In_1695,In_1895);
or U1013 (N_1013,In_1649,In_434);
and U1014 (N_1014,In_13,In_787);
or U1015 (N_1015,In_2464,N_233);
or U1016 (N_1016,N_542,In_281);
nand U1017 (N_1017,In_1142,N_290);
nand U1018 (N_1018,N_521,In_585);
and U1019 (N_1019,In_1568,In_136);
and U1020 (N_1020,In_2419,In_287);
or U1021 (N_1021,In_1302,In_206);
and U1022 (N_1022,In_1325,N_630);
or U1023 (N_1023,In_2169,N_730);
nand U1024 (N_1024,In_1825,In_864);
nor U1025 (N_1025,N_627,N_610);
nand U1026 (N_1026,N_959,N_341);
nand U1027 (N_1027,N_524,In_1405);
and U1028 (N_1028,N_900,N_950);
nor U1029 (N_1029,In_2192,N_622);
nor U1030 (N_1030,In_1471,N_989);
xnor U1031 (N_1031,In_1123,In_1335);
nand U1032 (N_1032,In_2455,N_847);
and U1033 (N_1033,In_2423,N_670);
or U1034 (N_1034,In_1238,In_927);
nand U1035 (N_1035,N_699,N_861);
nand U1036 (N_1036,In_2301,In_587);
nand U1037 (N_1037,In_240,In_2265);
xnor U1038 (N_1038,N_909,N_876);
or U1039 (N_1039,In_1814,N_894);
or U1040 (N_1040,N_245,N_974);
nand U1041 (N_1041,In_2306,N_557);
nand U1042 (N_1042,N_814,N_617);
xor U1043 (N_1043,In_1668,N_660);
and U1044 (N_1044,N_750,N_51);
and U1045 (N_1045,In_1689,In_447);
xor U1046 (N_1046,N_948,N_871);
xor U1047 (N_1047,In_158,N_715);
or U1048 (N_1048,N_835,N_802);
nor U1049 (N_1049,N_767,N_76);
nand U1050 (N_1050,In_1789,N_673);
xnor U1051 (N_1051,N_628,N_994);
or U1052 (N_1052,In_1432,N_527);
xor U1053 (N_1053,In_361,N_307);
nor U1054 (N_1054,N_127,In_801);
and U1055 (N_1055,N_504,In_2392);
nand U1056 (N_1056,N_862,N_969);
nand U1057 (N_1057,In_2108,In_2243);
or U1058 (N_1058,N_94,N_911);
and U1059 (N_1059,N_798,N_817);
or U1060 (N_1060,In_241,N_201);
nand U1061 (N_1061,N_778,In_2099);
xnor U1062 (N_1062,In_1864,N_96);
nor U1063 (N_1063,In_2250,N_513);
or U1064 (N_1064,N_377,In_1003);
or U1065 (N_1065,N_942,In_1548);
or U1066 (N_1066,In_2171,In_1829);
xor U1067 (N_1067,N_907,In_2486);
nand U1068 (N_1068,In_842,N_713);
or U1069 (N_1069,In_1234,In_196);
nor U1070 (N_1070,In_1033,In_2167);
xor U1071 (N_1071,N_634,N_554);
and U1072 (N_1072,N_874,N_43);
xnor U1073 (N_1073,N_463,In_2124);
xor U1074 (N_1074,In_41,In_519);
nand U1075 (N_1075,In_2096,In_2001);
and U1076 (N_1076,In_932,N_779);
nand U1077 (N_1077,In_875,In_1534);
and U1078 (N_1078,In_957,N_239);
xor U1079 (N_1079,In_2041,In_591);
and U1080 (N_1080,In_1813,In_22);
or U1081 (N_1081,In_1926,In_790);
nor U1082 (N_1082,N_705,N_815);
and U1083 (N_1083,In_322,In_1997);
nand U1084 (N_1084,N_376,In_1659);
xor U1085 (N_1085,N_532,In_428);
xnor U1086 (N_1086,In_2218,In_1784);
nor U1087 (N_1087,N_467,In_1920);
nor U1088 (N_1088,In_351,N_505);
or U1089 (N_1089,N_919,In_153);
and U1090 (N_1090,N_11,N_533);
and U1091 (N_1091,N_883,In_2449);
nand U1092 (N_1092,N_796,In_1792);
xnor U1093 (N_1093,In_2288,In_2209);
nand U1094 (N_1094,In_871,N_357);
nor U1095 (N_1095,In_2479,In_1707);
or U1096 (N_1096,In_1878,In_20);
xor U1097 (N_1097,In_1769,N_192);
nand U1098 (N_1098,In_909,N_441);
or U1099 (N_1099,N_537,In_1384);
and U1100 (N_1100,In_85,N_742);
nand U1101 (N_1101,In_1134,N_829);
xnor U1102 (N_1102,In_1733,In_617);
xnor U1103 (N_1103,N_843,In_2073);
nand U1104 (N_1104,N_680,N_936);
xor U1105 (N_1105,N_142,In_2068);
nand U1106 (N_1106,In_2163,In_418);
xor U1107 (N_1107,In_329,In_441);
or U1108 (N_1108,N_966,In_2482);
nand U1109 (N_1109,In_386,N_497);
and U1110 (N_1110,N_830,In_798);
nor U1111 (N_1111,N_841,N_840);
or U1112 (N_1112,In_987,N_998);
nand U1113 (N_1113,N_185,N_338);
nor U1114 (N_1114,In_763,N_529);
or U1115 (N_1115,N_115,N_388);
or U1116 (N_1116,In_1201,In_2436);
xnor U1117 (N_1117,N_553,N_816);
xor U1118 (N_1118,In_964,In_2399);
nand U1119 (N_1119,In_224,N_737);
nand U1120 (N_1120,In_1062,In_110);
nor U1121 (N_1121,N_552,N_327);
or U1122 (N_1122,N_315,In_2134);
nand U1123 (N_1123,In_1085,N_592);
and U1124 (N_1124,N_972,In_1124);
or U1125 (N_1125,In_231,In_1061);
xnor U1126 (N_1126,N_695,N_926);
nor U1127 (N_1127,N_783,In_2416);
nor U1128 (N_1128,N_770,N_786);
or U1129 (N_1129,In_667,In_296);
and U1130 (N_1130,N_589,In_366);
xnor U1131 (N_1131,N_203,In_438);
and U1132 (N_1132,In_1617,In_1244);
xnor U1133 (N_1133,N_120,N_932);
or U1134 (N_1134,N_935,N_656);
nor U1135 (N_1135,N_870,In_679);
or U1136 (N_1136,N_611,N_25);
and U1137 (N_1137,In_1894,N_822);
xor U1138 (N_1138,In_2386,N_87);
nand U1139 (N_1139,In_1817,N_10);
or U1140 (N_1140,N_860,N_973);
and U1141 (N_1141,In_794,N_800);
nand U1142 (N_1142,N_550,N_735);
xor U1143 (N_1143,N_775,In_1538);
or U1144 (N_1144,N_41,N_930);
xnor U1145 (N_1145,N_358,In_1938);
nand U1146 (N_1146,N_600,N_568);
and U1147 (N_1147,In_938,N_27);
nor U1148 (N_1148,In_2374,N_733);
xnor U1149 (N_1149,In_1745,N_342);
nor U1150 (N_1150,In_839,N_689);
xnor U1151 (N_1151,In_1572,In_881);
xnor U1152 (N_1152,N_291,N_510);
or U1153 (N_1153,N_649,N_166);
nand U1154 (N_1154,In_711,N_37);
xnor U1155 (N_1155,N_788,In_1905);
or U1156 (N_1156,N_754,N_752);
nand U1157 (N_1157,In_2433,In_2069);
xnor U1158 (N_1158,In_33,In_1731);
and U1159 (N_1159,In_867,In_2064);
nand U1160 (N_1160,In_687,In_1282);
or U1161 (N_1161,N_325,In_1002);
and U1162 (N_1162,N_390,N_769);
nor U1163 (N_1163,In_1927,In_487);
or U1164 (N_1164,N_851,In_761);
xor U1165 (N_1165,N_751,N_213);
or U1166 (N_1166,N_294,In_49);
nand U1167 (N_1167,N_639,In_173);
nand U1168 (N_1168,N_13,In_1798);
xnor U1169 (N_1169,In_1603,N_337);
or U1170 (N_1170,In_605,N_780);
xor U1171 (N_1171,In_1810,In_555);
or U1172 (N_1172,In_1265,N_464);
and U1173 (N_1173,N_782,In_911);
nor U1174 (N_1174,N_113,In_10);
xor U1175 (N_1175,N_5,In_545);
or U1176 (N_1176,N_956,N_606);
nor U1177 (N_1177,In_1587,In_1651);
or U1178 (N_1178,N_269,In_1137);
xnor U1179 (N_1179,N_888,In_690);
nor U1180 (N_1180,N_629,N_316);
nor U1181 (N_1181,In_1362,In_657);
xnor U1182 (N_1182,N_562,In_2397);
xor U1183 (N_1183,In_2354,In_1809);
xor U1184 (N_1184,In_698,N_356);
nand U1185 (N_1185,N_583,In_384);
or U1186 (N_1186,In_2176,N_465);
nand U1187 (N_1187,In_121,In_90);
nor U1188 (N_1188,N_619,In_890);
or U1189 (N_1189,N_150,N_724);
nand U1190 (N_1190,In_2418,In_223);
xnor U1191 (N_1191,N_241,N_503);
and U1192 (N_1192,N_336,In_1995);
nor U1193 (N_1193,N_762,N_765);
or U1194 (N_1194,N_612,N_479);
nor U1195 (N_1195,In_1203,N_624);
xnor U1196 (N_1196,In_1466,N_997);
xor U1197 (N_1197,N_107,N_616);
or U1198 (N_1198,In_993,In_460);
nand U1199 (N_1199,In_455,In_689);
or U1200 (N_1200,N_747,N_349);
nor U1201 (N_1201,In_1070,N_182);
or U1202 (N_1202,In_2121,In_775);
nand U1203 (N_1203,In_2427,N_66);
xor U1204 (N_1204,N_999,In_2100);
xnor U1205 (N_1205,In_183,In_636);
xnor U1206 (N_1206,N_884,In_326);
nand U1207 (N_1207,N_249,In_892);
nor U1208 (N_1208,N_489,N_787);
or U1209 (N_1209,In_2242,In_1671);
or U1210 (N_1210,In_2102,In_1052);
or U1211 (N_1211,N_460,In_342);
xnor U1212 (N_1212,N_712,In_1204);
nor U1213 (N_1213,In_2481,In_1876);
and U1214 (N_1214,In_466,In_1744);
or U1215 (N_1215,N_952,N_99);
and U1216 (N_1216,N_979,In_2129);
nand U1217 (N_1217,N_885,In_1506);
xor U1218 (N_1218,In_986,N_607);
nor U1219 (N_1219,N_519,In_359);
nor U1220 (N_1220,N_842,In_1808);
xor U1221 (N_1221,N_555,N_61);
nor U1222 (N_1222,N_945,N_636);
nand U1223 (N_1223,In_1831,In_1246);
and U1224 (N_1224,N_507,In_1434);
nor U1225 (N_1225,In_1090,In_829);
xnor U1226 (N_1226,In_1726,In_420);
xnor U1227 (N_1227,In_1976,In_1174);
nand U1228 (N_1228,N_785,N_173);
or U1229 (N_1229,N_873,N_716);
nor U1230 (N_1230,N_685,In_602);
xnor U1231 (N_1231,In_630,In_1812);
and U1232 (N_1232,In_1714,N_668);
or U1233 (N_1233,N_598,N_637);
and U1234 (N_1234,N_846,N_197);
and U1235 (N_1235,N_193,N_495);
xor U1236 (N_1236,N_613,In_2040);
xnor U1237 (N_1237,N_824,N_364);
or U1238 (N_1238,N_531,In_468);
nand U1239 (N_1239,In_2457,In_1010);
xor U1240 (N_1240,N_647,In_1255);
nand U1241 (N_1241,N_849,N_659);
xnor U1242 (N_1242,In_1011,In_1485);
or U1243 (N_1243,N_520,N_206);
nor U1244 (N_1244,In_9,N_625);
xor U1245 (N_1245,N_955,N_255);
or U1246 (N_1246,In_1550,In_2255);
nor U1247 (N_1247,N_155,In_710);
nand U1248 (N_1248,In_910,In_1700);
nor U1249 (N_1249,In_1275,N_350);
and U1250 (N_1250,In_943,N_658);
nor U1251 (N_1251,N_323,N_544);
nand U1252 (N_1252,N_615,N_881);
or U1253 (N_1253,In_1754,In_1987);
nor U1254 (N_1254,In_1231,In_464);
nor U1255 (N_1255,N_64,N_571);
nand U1256 (N_1256,In_1422,N_967);
nor U1257 (N_1257,N_407,In_297);
nand U1258 (N_1258,N_734,In_2106);
xnor U1259 (N_1259,N_897,N_516);
or U1260 (N_1260,N_204,In_756);
and U1261 (N_1261,N_771,N_561);
and U1262 (N_1262,N_430,N_991);
xnor U1263 (N_1263,In_527,N_116);
nor U1264 (N_1264,In_1456,N_438);
and U1265 (N_1265,N_650,In_1050);
or U1266 (N_1266,In_646,In_2440);
nand U1267 (N_1267,In_1251,N_844);
nor U1268 (N_1268,N_913,N_492);
nand U1269 (N_1269,N_215,N_139);
nor U1270 (N_1270,N_603,In_838);
or U1271 (N_1271,In_1103,In_548);
nand U1272 (N_1272,In_1884,N_962);
or U1273 (N_1273,N_586,N_135);
nor U1274 (N_1274,N_681,In_1496);
nor U1275 (N_1275,In_1536,N_331);
xnor U1276 (N_1276,N_470,N_488);
nand U1277 (N_1277,In_556,In_142);
nor U1278 (N_1278,N_604,In_730);
and U1279 (N_1279,N_865,In_1012);
nor U1280 (N_1280,In_2050,N_757);
nor U1281 (N_1281,N_963,N_914);
or U1282 (N_1282,In_700,N_958);
nand U1283 (N_1283,In_1529,In_1653);
or U1284 (N_1284,N_941,N_801);
xnor U1285 (N_1285,In_2127,In_79);
nor U1286 (N_1286,N_764,N_867);
nand U1287 (N_1287,In_1628,N_400);
or U1288 (N_1288,In_238,In_983);
xor U1289 (N_1289,N_792,In_666);
or U1290 (N_1290,N_183,In_2313);
nand U1291 (N_1291,N_21,N_593);
nand U1292 (N_1292,N_838,In_1323);
nand U1293 (N_1293,N_644,N_664);
nor U1294 (N_1294,N_632,In_1685);
and U1295 (N_1295,N_698,N_799);
nor U1296 (N_1296,N_361,N_853);
or U1297 (N_1297,N_534,In_2333);
and U1298 (N_1298,In_616,In_1401);
nand U1299 (N_1299,In_1411,N_635);
or U1300 (N_1300,In_1566,N_347);
xnor U1301 (N_1301,N_573,In_1279);
or U1302 (N_1302,In_197,In_419);
xor U1303 (N_1303,In_1104,N_875);
nor U1304 (N_1304,N_275,N_813);
and U1305 (N_1305,N_30,N_731);
or U1306 (N_1306,In_2432,In_387);
nand U1307 (N_1307,N_806,In_2088);
and U1308 (N_1308,In_1877,N_790);
nand U1309 (N_1309,N_923,In_448);
xor U1310 (N_1310,N_205,N_784);
and U1311 (N_1311,N_386,In_2206);
nand U1312 (N_1312,In_116,N_903);
or U1313 (N_1313,In_453,N_672);
or U1314 (N_1314,In_1136,N_345);
nand U1315 (N_1315,N_602,In_98);
xor U1316 (N_1316,In_2411,In_944);
xnor U1317 (N_1317,N_69,In_2234);
and U1318 (N_1318,N_745,N_714);
nand U1319 (N_1319,In_1626,In_607);
nand U1320 (N_1320,N_167,In_808);
and U1321 (N_1321,In_1505,N_270);
and U1322 (N_1322,N_285,N_599);
or U1323 (N_1323,In_1488,In_1512);
nor U1324 (N_1324,N_721,In_1605);
or U1325 (N_1325,N_117,N_905);
nor U1326 (N_1326,N_812,In_582);
or U1327 (N_1327,In_1262,In_2485);
xnor U1328 (N_1328,In_1636,In_549);
and U1329 (N_1329,N_49,In_207);
nand U1330 (N_1330,N_833,N_86);
nand U1331 (N_1331,N_153,N_920);
or U1332 (N_1332,N_423,In_542);
xor U1333 (N_1333,In_2303,In_118);
xor U1334 (N_1334,In_1465,In_2271);
nand U1335 (N_1335,In_1500,N_576);
nand U1336 (N_1336,In_1503,In_861);
or U1337 (N_1337,N_901,N_702);
nor U1338 (N_1338,In_2142,In_1028);
xnor U1339 (N_1339,In_171,N_587);
nor U1340 (N_1340,N_605,In_1641);
and U1341 (N_1341,In_1848,In_1018);
and U1342 (N_1342,In_457,N_403);
and U1343 (N_1343,N_209,N_312);
xor U1344 (N_1344,N_866,In_1801);
or U1345 (N_1345,N_645,In_1115);
xnor U1346 (N_1346,N_597,In_1149);
nor U1347 (N_1347,In_2103,In_1803);
nor U1348 (N_1348,In_1858,N_302);
and U1349 (N_1349,N_230,In_237);
nand U1350 (N_1350,In_2489,N_776);
nor U1351 (N_1351,In_2309,N_404);
nand U1352 (N_1352,In_7,N_882);
or U1353 (N_1353,N_228,In_2400);
nand U1354 (N_1354,N_191,N_330);
or U1355 (N_1355,In_816,N_559);
nor U1356 (N_1356,In_1730,In_1941);
or U1357 (N_1357,N_692,In_2056);
xor U1358 (N_1358,N_982,N_448);
and U1359 (N_1359,N_276,In_2316);
or U1360 (N_1360,N_219,In_101);
xor U1361 (N_1361,In_1964,In_2145);
nand U1362 (N_1362,In_311,N_688);
and U1363 (N_1363,N_71,In_2084);
nand U1364 (N_1364,In_1952,N_917);
nand U1365 (N_1365,N_697,In_1741);
nor U1366 (N_1366,In_410,N_976);
or U1367 (N_1367,In_1152,In_2438);
nand U1368 (N_1368,In_2498,In_1495);
and U1369 (N_1369,In_908,In_103);
xor U1370 (N_1370,In_276,In_1786);
and U1371 (N_1371,N_367,In_29);
and U1372 (N_1372,In_87,In_1690);
nor U1373 (N_1373,In_1855,N_581);
and U1374 (N_1374,In_1365,In_1378);
and U1375 (N_1375,In_2294,N_156);
nand U1376 (N_1376,N_77,N_981);
nor U1377 (N_1377,In_1961,N_320);
nor U1378 (N_1378,N_717,In_1750);
nor U1379 (N_1379,In_267,In_1743);
xnor U1380 (N_1380,N_575,N_988);
nor U1381 (N_1381,In_1350,In_935);
or U1382 (N_1382,In_1739,In_1883);
xor U1383 (N_1383,In_1481,In_1122);
xnor U1384 (N_1384,N_195,N_937);
xor U1385 (N_1385,N_468,N_236);
xor U1386 (N_1386,In_592,In_895);
nor U1387 (N_1387,In_86,In_1094);
and U1388 (N_1388,In_1389,In_1418);
and U1389 (N_1389,N_582,In_1736);
and U1390 (N_1390,In_1442,In_409);
and U1391 (N_1391,In_1407,In_662);
nand U1392 (N_1392,N_427,N_655);
nand U1393 (N_1393,In_1311,N_995);
nand U1394 (N_1394,N_585,N_351);
nor U1395 (N_1395,In_300,In_1266);
nand U1396 (N_1396,In_137,In_2331);
nor U1397 (N_1397,In_739,N_946);
and U1398 (N_1398,N_886,N_700);
and U1399 (N_1399,N_300,In_528);
nor U1400 (N_1400,In_894,In_1132);
nand U1401 (N_1401,In_2141,N_662);
nand U1402 (N_1402,In_372,In_1791);
nand U1403 (N_1403,N_79,In_888);
nor U1404 (N_1404,N_151,In_2425);
or U1405 (N_1405,N_703,In_831);
nor U1406 (N_1406,In_1069,N_910);
nand U1407 (N_1407,In_1468,In_2079);
nand U1408 (N_1408,In_613,In_1760);
nor U1409 (N_1409,N_346,In_629);
nand U1410 (N_1410,In_2484,N_237);
or U1411 (N_1411,In_2083,N_382);
nand U1412 (N_1412,N_683,N_992);
or U1413 (N_1413,In_289,In_1469);
nand U1414 (N_1414,N_498,N_591);
or U1415 (N_1415,N_539,In_1046);
xor U1416 (N_1416,N_412,In_1772);
nand U1417 (N_1417,N_543,N_727);
xor U1418 (N_1418,N_310,In_977);
nor U1419 (N_1419,N_522,In_124);
nand U1420 (N_1420,N_933,N_83);
xnor U1421 (N_1421,In_1131,In_264);
nand U1422 (N_1422,N_433,N_915);
or U1423 (N_1423,N_964,N_854);
nand U1424 (N_1424,In_1957,In_489);
nor U1425 (N_1425,In_385,N_898);
nor U1426 (N_1426,N_766,In_588);
and U1427 (N_1427,N_729,N_810);
and U1428 (N_1428,N_523,In_1226);
xnor U1429 (N_1429,N_686,N_160);
nor U1430 (N_1430,N_922,In_1135);
nand U1431 (N_1431,N_565,In_788);
xnor U1432 (N_1432,In_2143,In_770);
nor U1433 (N_1433,In_1642,N_384);
nand U1434 (N_1434,N_748,In_135);
nand U1435 (N_1435,N_88,N_749);
xor U1436 (N_1436,N_934,In_2091);
nor U1437 (N_1437,In_360,In_1037);
xor U1438 (N_1438,N_643,In_246);
nor U1439 (N_1439,In_1490,In_2021);
nor U1440 (N_1440,In_506,In_1806);
nor U1441 (N_1441,In_846,In_318);
xor U1442 (N_1442,N_985,N_711);
nor U1443 (N_1443,N_267,In_702);
and U1444 (N_1444,N_137,N_809);
nand U1445 (N_1445,In_1985,N_640);
nor U1446 (N_1446,N_987,N_34);
or U1447 (N_1447,N_878,N_558);
nand U1448 (N_1448,N_677,In_126);
nand U1449 (N_1449,In_1623,N_512);
or U1450 (N_1450,In_2003,In_748);
xnor U1451 (N_1451,N_506,In_1970);
and U1452 (N_1452,In_1851,N_128);
xor U1453 (N_1453,In_371,In_476);
xnor U1454 (N_1454,N_578,In_298);
and U1455 (N_1455,N_667,In_1236);
or U1456 (N_1456,N_912,N_208);
nand U1457 (N_1457,N_514,In_1185);
nor U1458 (N_1458,N_231,N_526);
nor U1459 (N_1459,N_344,In_295);
nor U1460 (N_1460,N_722,N_805);
nand U1461 (N_1461,In_2442,N_560);
nor U1462 (N_1462,N_904,In_1356);
nor U1463 (N_1463,N_743,In_655);
xnor U1464 (N_1464,In_1584,N_718);
nor U1465 (N_1465,In_2334,N_676);
xnor U1466 (N_1466,In_2179,N_857);
nor U1467 (N_1467,In_1197,N_704);
and U1468 (N_1468,N_7,N_696);
nor U1469 (N_1469,In_478,N_395);
and U1470 (N_1470,N_652,In_42);
and U1471 (N_1471,N_104,In_2170);
and U1472 (N_1472,In_1596,N_405);
or U1473 (N_1473,In_2256,N_73);
nand U1474 (N_1474,N_868,N_620);
nand U1475 (N_1475,In_1303,N_665);
xnor U1476 (N_1476,N_85,In_2431);
xor U1477 (N_1477,N_161,In_2188);
and U1478 (N_1478,In_1643,N_789);
xor U1479 (N_1479,N_674,In_2233);
or U1480 (N_1480,In_2415,N_965);
xor U1481 (N_1481,In_2383,N_863);
and U1482 (N_1482,In_1710,N_756);
or U1483 (N_1483,In_2393,In_83);
nand U1484 (N_1484,In_1909,N_446);
or U1485 (N_1485,In_1615,In_218);
nand U1486 (N_1486,N_687,N_951);
or U1487 (N_1487,N_157,N_855);
and U1488 (N_1488,N_623,N_194);
nor U1489 (N_1489,In_640,N_471);
xor U1490 (N_1490,N_682,N_306);
or U1491 (N_1491,In_539,In_1607);
and U1492 (N_1492,N_199,In_2104);
xor U1493 (N_1493,In_1897,N_826);
or U1494 (N_1494,N_141,N_540);
or U1495 (N_1495,In_1438,In_168);
nand U1496 (N_1496,N_299,N_601);
nor U1497 (N_1497,In_1729,In_2199);
or U1498 (N_1498,In_855,In_1444);
nor U1499 (N_1499,N_899,In_1147);
or U1500 (N_1500,N_1093,N_1468);
or U1501 (N_1501,N_397,N_819);
and U1502 (N_1502,N_1097,N_1246);
or U1503 (N_1503,In_1464,N_1298);
or U1504 (N_1504,In_1404,N_924);
xor U1505 (N_1505,N_1132,N_621);
or U1506 (N_1506,N_1213,N_1477);
nand U1507 (N_1507,N_694,In_57);
xnor U1508 (N_1508,N_1170,In_55);
nor U1509 (N_1509,N_1163,N_1304);
xor U1510 (N_1510,N_370,N_1455);
xor U1511 (N_1511,N_1055,N_1159);
xor U1512 (N_1512,In_891,N_1343);
or U1513 (N_1513,N_1098,N_410);
nor U1514 (N_1514,N_1281,N_1374);
or U1515 (N_1515,In_244,N_1221);
xnor U1516 (N_1516,N_1422,N_978);
xor U1517 (N_1517,N_1239,N_690);
or U1518 (N_1518,In_896,N_1369);
nor U1519 (N_1519,N_1035,N_1331);
nand U1520 (N_1520,N_1418,N_872);
nand U1521 (N_1521,N_1259,N_1146);
xnor U1522 (N_1522,N_1424,N_710);
xor U1523 (N_1523,In_470,N_334);
xor U1524 (N_1524,N_1140,N_1006);
and U1525 (N_1525,In_1242,N_1332);
nand U1526 (N_1526,N_1254,In_2321);
xor U1527 (N_1527,In_2263,N_580);
nor U1528 (N_1528,N_706,N_1349);
nor U1529 (N_1529,N_175,N_1032);
nand U1530 (N_1530,N_1184,N_93);
and U1531 (N_1531,N_827,N_1393);
or U1532 (N_1532,In_696,N_1172);
nand U1533 (N_1533,In_1645,In_2367);
xor U1534 (N_1534,In_160,N_1101);
nand U1535 (N_1535,N_159,N_1021);
nor U1536 (N_1536,N_1287,N_1256);
xnor U1537 (N_1537,In_2252,N_738);
and U1538 (N_1538,N_1451,In_108);
and U1539 (N_1539,N_1014,N_1071);
and U1540 (N_1540,N_502,In_2160);
and U1541 (N_1541,In_1557,In_2268);
nand U1542 (N_1542,N_222,In_1019);
nor U1543 (N_1543,N_1201,N_530);
nand U1544 (N_1544,N_1472,N_1397);
nor U1545 (N_1545,N_823,In_621);
and U1546 (N_1546,N_1316,N_474);
nand U1547 (N_1547,N_1238,In_1727);
xnor U1548 (N_1548,N_1350,N_303);
nor U1549 (N_1549,N_259,N_1203);
xor U1550 (N_1550,N_1497,N_1387);
nor U1551 (N_1551,In_2377,N_1122);
nand U1552 (N_1552,N_1312,N_1094);
or U1553 (N_1553,N_145,N_1233);
xor U1554 (N_1554,N_1300,N_1029);
and U1555 (N_1555,N_1416,N_1430);
nor U1556 (N_1556,N_1116,N_1037);
or U1557 (N_1557,N_1191,In_725);
or U1558 (N_1558,N_1067,In_1646);
nand U1559 (N_1559,N_1443,In_547);
and U1560 (N_1560,N_1268,N_1200);
xor U1561 (N_1561,N_1381,In_346);
xnor U1562 (N_1562,N_1015,N_1235);
and U1563 (N_1563,In_1436,In_1766);
or U1564 (N_1564,N_741,N_511);
or U1565 (N_1565,N_1118,N_1127);
nor U1566 (N_1566,N_286,N_1216);
and U1567 (N_1567,N_726,In_1622);
nand U1568 (N_1568,N_891,N_1417);
and U1569 (N_1569,N_1475,In_1451);
and U1570 (N_1570,N_1237,N_1411);
or U1571 (N_1571,N_869,In_976);
or U1572 (N_1572,N_1117,N_1380);
nor U1573 (N_1573,N_1234,N_1026);
nor U1574 (N_1574,In_1252,N_1103);
and U1575 (N_1575,N_55,In_199);
nor U1576 (N_1576,N_1107,N_1222);
or U1577 (N_1577,N_508,N_58);
or U1578 (N_1578,N_1211,In_2385);
nand U1579 (N_1579,In_2361,N_535);
xor U1580 (N_1580,N_1473,N_893);
and U1581 (N_1581,In_1822,N_556);
or U1582 (N_1582,N_648,N_1167);
nor U1583 (N_1583,In_1579,N_1210);
nand U1584 (N_1584,N_1013,In_2089);
or U1585 (N_1585,N_1450,In_682);
xor U1586 (N_1586,In_1412,N_1);
or U1587 (N_1587,N_1306,N_1370);
nor U1588 (N_1588,N_1137,N_1408);
and U1589 (N_1589,In_1146,In_1683);
xor U1590 (N_1590,N_772,N_1485);
nand U1591 (N_1591,N_1181,N_1358);
nand U1592 (N_1592,N_1257,In_1644);
or U1593 (N_1593,In_2178,N_1039);
nor U1594 (N_1594,N_1145,N_31);
nor U1595 (N_1595,N_1012,In_812);
and U1596 (N_1596,N_1175,In_1357);
nand U1597 (N_1597,In_2063,N_1119);
nor U1598 (N_1598,N_566,In_1778);
nor U1599 (N_1599,N_968,N_931);
nor U1600 (N_1600,In_589,N_1056);
nor U1601 (N_1601,N_1025,N_1484);
and U1602 (N_1602,N_1034,N_1396);
nand U1603 (N_1603,N_1091,N_14);
and U1604 (N_1604,N_480,N_1465);
xor U1605 (N_1605,In_427,N_551);
nand U1606 (N_1606,N_927,N_1173);
nand U1607 (N_1607,In_35,N_1318);
nand U1608 (N_1608,N_1290,N_1206);
xor U1609 (N_1609,In_426,N_1368);
and U1610 (N_1610,N_990,N_1125);
nand U1611 (N_1611,In_1326,In_695);
nor U1612 (N_1612,N_638,N_1470);
nand U1613 (N_1613,N_114,N_154);
nor U1614 (N_1614,N_1187,In_810);
or U1615 (N_1615,In_1000,N_1390);
or U1616 (N_1616,N_641,N_1134);
nor U1617 (N_1617,N_1018,N_661);
nor U1618 (N_1618,N_746,N_1412);
nand U1619 (N_1619,N_326,N_1453);
nor U1620 (N_1620,N_1068,N_1362);
nand U1621 (N_1621,In_1681,N_1218);
and U1622 (N_1622,N_1344,N_1367);
and U1623 (N_1623,N_1142,In_1833);
xnor U1624 (N_1624,In_597,N_1440);
nor U1625 (N_1625,N_720,N_1309);
xnor U1626 (N_1626,N_563,In_1289);
nand U1627 (N_1627,N_579,N_1208);
nor U1628 (N_1628,N_1372,N_1478);
nor U1629 (N_1629,In_884,N_1249);
nor U1630 (N_1630,N_354,In_1602);
nor U1631 (N_1631,In_449,N_1214);
nor U1632 (N_1632,N_186,N_791);
xor U1633 (N_1633,N_693,N_654);
nand U1634 (N_1634,N_1169,In_1785);
xnor U1635 (N_1635,N_675,N_1467);
xnor U1636 (N_1636,N_119,N_1041);
and U1637 (N_1637,In_8,N_850);
xnor U1638 (N_1638,N_1064,In_800);
nand U1639 (N_1639,N_1202,N_1204);
xor U1640 (N_1640,N_1051,In_321);
and U1641 (N_1641,N_1148,N_758);
nand U1642 (N_1642,N_1095,In_2202);
and U1643 (N_1643,N_1199,N_755);
or U1644 (N_1644,N_975,N_1436);
and U1645 (N_1645,In_1138,N_1087);
xnor U1646 (N_1646,N_1313,N_340);
or U1647 (N_1647,N_1420,In_1914);
nor U1648 (N_1648,N_1152,N_1247);
and U1649 (N_1649,N_577,N_1019);
nand U1650 (N_1650,N_1174,N_1225);
or U1651 (N_1651,N_1263,N_1435);
nor U1652 (N_1652,N_1385,N_618);
or U1653 (N_1653,N_1048,N_1124);
xnor U1654 (N_1654,N_1295,N_1399);
nor U1655 (N_1655,N_1166,In_1706);
nor U1656 (N_1656,N_1339,N_1441);
and U1657 (N_1657,N_1150,N_1275);
nand U1658 (N_1658,N_408,N_273);
nor U1659 (N_1659,N_1000,N_1498);
and U1660 (N_1660,N_1409,N_1315);
nor U1661 (N_1661,N_1302,N_1022);
nor U1662 (N_1662,N_908,N_797);
and U1663 (N_1663,N_75,N_820);
or U1664 (N_1664,In_1021,N_1400);
nand U1665 (N_1665,N_832,In_714);
nand U1666 (N_1666,N_1059,N_1293);
nor U1667 (N_1667,In_1722,N_1311);
nor U1668 (N_1668,N_1080,N_781);
nor U1669 (N_1669,N_1156,N_1286);
nand U1670 (N_1670,N_1189,In_2407);
xor U1671 (N_1671,N_1359,N_1317);
and U1672 (N_1672,In_1963,N_1490);
nor U1673 (N_1673,N_1326,N_993);
nand U1674 (N_1674,N_1027,N_1002);
nor U1675 (N_1675,N_1182,N_1147);
nor U1676 (N_1676,N_133,In_1633);
or U1677 (N_1677,N_1066,In_1440);
nand U1678 (N_1678,N_1195,N_1266);
and U1679 (N_1679,N_1277,N_373);
or U1680 (N_1680,N_1158,N_657);
xnor U1681 (N_1681,N_1232,In_1109);
and U1682 (N_1682,N_1354,N_1310);
or U1683 (N_1683,In_53,N_1045);
nand U1684 (N_1684,N_92,N_118);
and U1685 (N_1685,In_1673,N_1459);
nor U1686 (N_1686,N_1105,N_845);
and U1687 (N_1687,N_1325,N_1267);
xor U1688 (N_1688,N_1043,N_921);
or U1689 (N_1689,N_1322,N_422);
nor U1690 (N_1690,N_759,N_1241);
or U1691 (N_1691,N_232,N_379);
or U1692 (N_1692,N_1391,N_1229);
or U1693 (N_1693,N_1480,N_1328);
and U1694 (N_1694,N_1243,In_345);
nor U1695 (N_1695,N_1437,N_1338);
nand U1696 (N_1696,In_902,N_1086);
nor U1697 (N_1697,N_821,In_1430);
nor U1698 (N_1698,N_1128,N_1272);
xnor U1699 (N_1699,N_774,N_1255);
nand U1700 (N_1700,N_1405,N_1378);
nor U1701 (N_1701,N_536,N_1323);
xor U1702 (N_1702,N_1461,N_1296);
and U1703 (N_1703,N_1346,N_1428);
and U1704 (N_1704,In_396,In_48);
nand U1705 (N_1705,N_1355,N_1162);
or U1706 (N_1706,N_1361,N_1090);
nand U1707 (N_1707,N_1143,N_925);
nor U1708 (N_1708,N_517,N_486);
or U1709 (N_1709,In_239,In_444);
xor U1710 (N_1710,N_1220,N_1395);
or U1711 (N_1711,N_723,N_808);
and U1712 (N_1712,N_1016,N_44);
or U1713 (N_1713,N_1274,N_1321);
nor U1714 (N_1714,N_1177,N_1429);
nor U1715 (N_1715,In_499,N_1212);
nor U1716 (N_1716,In_1647,N_499);
or U1717 (N_1717,N_996,N_939);
nand U1718 (N_1718,N_1042,N_431);
and U1719 (N_1719,N_1058,In_1869);
xnor U1720 (N_1720,N_1262,In_939);
xnor U1721 (N_1721,In_245,N_1379);
nor U1722 (N_1722,N_892,In_317);
xor U1723 (N_1723,N_1063,N_1138);
nor U1724 (N_1724,N_1342,N_1144);
or U1725 (N_1725,N_402,N_760);
nor U1726 (N_1726,N_1193,N_839);
nor U1727 (N_1727,N_1226,In_1635);
nor U1728 (N_1728,N_1444,In_1560);
xnor U1729 (N_1729,In_843,N_834);
nand U1730 (N_1730,N_916,N_1336);
nand U1731 (N_1731,N_1129,In_769);
nor U1732 (N_1732,N_1340,In_19);
xor U1733 (N_1733,N_1327,N_1010);
and U1734 (N_1734,N_1419,In_2249);
and U1735 (N_1735,In_2469,N_1375);
xor U1736 (N_1736,In_2283,N_1130);
xnor U1737 (N_1737,N_1265,In_784);
and U1738 (N_1738,N_1194,N_666);
nor U1739 (N_1739,N_509,N_42);
nand U1740 (N_1740,In_1705,N_1463);
nand U1741 (N_1741,N_1292,N_1100);
and U1742 (N_1742,N_1111,In_1294);
or U1743 (N_1743,In_708,In_1420);
nand U1744 (N_1744,N_1062,N_1383);
xnor U1745 (N_1745,In_461,In_1363);
or U1746 (N_1746,In_272,N_1269);
and U1747 (N_1747,N_1495,N_547);
nand U1748 (N_1748,N_1242,N_252);
nor U1749 (N_1749,N_1464,N_859);
or U1750 (N_1750,In_269,In_959);
xnor U1751 (N_1751,N_170,In_1525);
nor U1752 (N_1752,In_283,N_1324);
nor U1753 (N_1753,N_970,N_918);
or U1754 (N_1754,In_172,N_1357);
nand U1755 (N_1755,N_1054,N_887);
or U1756 (N_1756,N_1394,In_1368);
nand U1757 (N_1757,N_1230,N_980);
nand U1758 (N_1758,N_1421,N_736);
nor U1759 (N_1759,N_1431,N_1044);
nand U1760 (N_1760,In_604,In_723);
and U1761 (N_1761,N_1060,N_295);
xor U1762 (N_1762,N_1228,N_1007);
and U1763 (N_1763,In_736,N_1223);
and U1764 (N_1764,N_1365,N_481);
nand U1765 (N_1765,N_451,N_1449);
or U1766 (N_1766,In_232,N_126);
xnor U1767 (N_1767,N_1489,N_837);
or U1768 (N_1768,In_971,In_970);
or U1769 (N_1769,N_1192,N_332);
nor U1770 (N_1770,N_1001,N_375);
and U1771 (N_1771,N_1154,N_1433);
nor U1772 (N_1772,N_1377,N_1329);
and U1773 (N_1773,N_1360,N_1185);
nand U1774 (N_1774,N_1320,N_1407);
or U1775 (N_1775,N_260,N_1479);
and U1776 (N_1776,N_983,N_763);
nand U1777 (N_1777,In_120,N_1115);
or U1778 (N_1778,N_1289,N_1109);
nand U1779 (N_1779,In_1487,N_1186);
or U1780 (N_1780,N_1305,N_1283);
nand U1781 (N_1781,N_1009,N_1386);
xor U1782 (N_1782,In_2272,N_425);
nor U1783 (N_1783,In_854,N_631);
nand U1784 (N_1784,N_1448,In_24);
or U1785 (N_1785,N_1057,N_1426);
and U1786 (N_1786,N_902,N_541);
and U1787 (N_1787,N_570,In_1595);
or U1788 (N_1788,N_1047,N_1217);
and U1789 (N_1789,N_1072,In_1992);
xnor U1790 (N_1790,In_954,N_381);
or U1791 (N_1791,In_1824,N_1423);
nand U1792 (N_1792,In_760,N_179);
xor U1793 (N_1793,N_1089,In_560);
and U1794 (N_1794,N_856,N_1053);
nor U1795 (N_1795,N_1092,N_773);
and U1796 (N_1796,N_1425,N_1088);
and U1797 (N_1797,N_548,N_176);
nand U1798 (N_1798,N_1341,N_1384);
nor U1799 (N_1799,N_564,N_957);
nor U1800 (N_1800,N_954,In_2467);
or U1801 (N_1801,N_1176,N_1307);
nor U1802 (N_1802,N_472,N_707);
and U1803 (N_1803,In_1717,N_4);
nand U1804 (N_1804,In_76,N_1356);
nand U1805 (N_1805,N_663,In_717);
and U1806 (N_1806,N_1197,In_319);
or U1807 (N_1807,N_1040,N_595);
or U1808 (N_1808,In_1352,N_1398);
xnor U1809 (N_1809,N_1165,N_220);
nand U1810 (N_1810,N_1347,N_1244);
nor U1811 (N_1811,N_1149,N_1337);
or U1812 (N_1812,N_1081,In_546);
nand U1813 (N_1813,N_1078,N_614);
and U1814 (N_1814,N_1496,N_174);
nor U1815 (N_1815,N_1073,N_1270);
and U1816 (N_1816,N_1294,N_1382);
and U1817 (N_1817,In_1954,N_1434);
and U1818 (N_1818,In_1391,N_1446);
nor U1819 (N_1819,N_811,N_1258);
and U1820 (N_1820,N_1108,N_1179);
and U1821 (N_1821,In_129,N_1401);
nor U1822 (N_1822,In_1499,N_1288);
nand U1823 (N_1823,N_971,N_588);
xor U1824 (N_1824,N_65,In_1256);
and U1825 (N_1825,N_669,N_889);
xor U1826 (N_1826,N_1126,In_1317);
xor U1827 (N_1827,In_612,N_895);
nand U1828 (N_1828,N_1297,N_1084);
nor U1829 (N_1829,N_1215,N_1240);
and U1830 (N_1830,N_1178,N_1028);
or U1831 (N_1831,N_1075,In_972);
nand U1832 (N_1832,N_1456,N_1279);
xnor U1833 (N_1833,N_1236,N_1348);
xnor U1834 (N_1834,N_1276,In_832);
nand U1835 (N_1835,In_12,In_1865);
nand U1836 (N_1836,N_1363,N_1492);
or U1837 (N_1837,N_609,In_1889);
nand U1838 (N_1838,N_1494,N_1427);
nand U1839 (N_1839,N_626,In_170);
xnor U1840 (N_1840,N_725,N_234);
and U1841 (N_1841,N_1131,N_1314);
or U1842 (N_1842,N_1432,N_1458);
xor U1843 (N_1843,N_292,N_1392);
xor U1844 (N_1844,N_1261,N_1333);
nor U1845 (N_1845,N_836,N_1413);
nor U1846 (N_1846,In_1117,N_1036);
xor U1847 (N_1847,N_1488,N_198);
nor U1848 (N_1848,N_419,In_1988);
and U1849 (N_1849,N_1038,N_1112);
nand U1850 (N_1850,N_46,In_2005);
or U1851 (N_1851,In_1795,N_768);
nor U1852 (N_1852,N_1011,In_904);
nor U1853 (N_1853,In_2304,N_1457);
nand U1854 (N_1854,N_679,N_1005);
nand U1855 (N_1855,N_596,N_739);
xor U1856 (N_1856,In_215,N_794);
nand U1857 (N_1857,In_677,N_223);
xor U1858 (N_1858,In_2279,N_1250);
nand U1859 (N_1859,In_1780,N_1133);
nand U1860 (N_1860,N_938,N_29);
xnor U1861 (N_1861,N_1023,In_663);
xor U1862 (N_1862,N_1121,N_1123);
nor U1863 (N_1863,N_105,In_681);
nor U1864 (N_1864,N_1079,N_761);
xor U1865 (N_1865,N_1491,N_26);
and U1866 (N_1866,In_452,N_653);
and U1867 (N_1867,N_1224,In_59);
and U1868 (N_1868,N_1319,In_1948);
and U1869 (N_1869,N_343,N_807);
and U1870 (N_1870,N_91,In_1093);
or U1871 (N_1871,N_1403,N_1070);
xnor U1872 (N_1872,N_691,N_1110);
and U1873 (N_1873,N_1483,N_928);
nand U1874 (N_1874,N_1280,N_1164);
nor U1875 (N_1875,N_594,N_1003);
nand U1876 (N_1876,N_929,N_1077);
or U1877 (N_1877,N_1106,In_2024);
nor U1878 (N_1878,N_1161,In_960);
or U1879 (N_1879,N_753,In_1166);
nand U1880 (N_1880,N_1445,N_1482);
xor U1881 (N_1881,N_528,In_2211);
xor U1882 (N_1882,N_1373,N_1352);
xor U1883 (N_1883,In_511,In_1841);
and U1884 (N_1884,In_752,N_1487);
nor U1885 (N_1885,In_1338,In_357);
nor U1886 (N_1886,N_890,N_1168);
nor U1887 (N_1887,N_1260,In_2493);
nand U1888 (N_1888,N_1499,N_40);
nor U1889 (N_1889,N_447,N_1160);
or U1890 (N_1890,In_1966,N_1020);
nor U1891 (N_1891,N_671,N_880);
xor U1892 (N_1892,N_1096,N_977);
or U1893 (N_1893,In_899,N_709);
xnor U1894 (N_1894,N_684,N_1330);
nand U1895 (N_1895,In_2161,In_942);
xor U1896 (N_1896,N_1139,N_701);
nand U1897 (N_1897,In_1170,In_252);
nand U1898 (N_1898,In_672,N_1209);
and U1899 (N_1899,N_1008,N_545);
nor U1900 (N_1900,N_574,In_2144);
nor U1901 (N_1901,N_1273,N_1061);
or U1902 (N_1902,In_2095,N_242);
nor U1903 (N_1903,N_1151,N_1345);
and U1904 (N_1904,N_825,N_567);
or U1905 (N_1905,N_1046,N_1402);
nand U1906 (N_1906,N_1180,N_1074);
xor U1907 (N_1907,N_1389,N_719);
nand U1908 (N_1908,In_1321,N_1406);
nand U1909 (N_1909,In_807,N_1452);
and U1910 (N_1910,N_264,N_708);
nor U1911 (N_1911,N_1410,In_1194);
xnor U1912 (N_1912,In_1664,N_584);
xor U1913 (N_1913,In_728,In_934);
or U1914 (N_1914,N_1114,N_1371);
nor U1915 (N_1915,In_294,N_1207);
nand U1916 (N_1916,N_394,N_1469);
and U1917 (N_1917,In_198,N_1155);
nor U1918 (N_1918,N_261,In_1476);
xnor U1919 (N_1919,N_90,N_1474);
nand U1920 (N_1920,In_2155,N_984);
and U1921 (N_1921,N_1454,In_1900);
and U1922 (N_1922,In_2034,N_1284);
and U1923 (N_1923,In_303,N_1017);
and U1924 (N_1924,In_25,In_68);
nand U1925 (N_1925,N_1415,In_1682);
or U1926 (N_1926,N_740,N_1198);
and U1927 (N_1927,N_1076,N_1353);
nand U1928 (N_1928,N_546,N_1291);
xor U1929 (N_1929,N_1136,N_442);
nand U1930 (N_1930,In_966,N_1219);
xnor U1931 (N_1931,N_1285,In_691);
nand U1932 (N_1932,In_1227,In_2080);
nor U1933 (N_1933,N_947,N_953);
xnor U1934 (N_1934,N_20,N_1252);
xor U1935 (N_1935,N_1486,In_70);
and U1936 (N_1936,In_948,N_642);
nor U1937 (N_1937,N_1334,In_1968);
and U1938 (N_1938,N_1171,N_549);
xnor U1939 (N_1939,N_943,In_516);
xnor U1940 (N_1940,N_1050,N_1231);
nor U1941 (N_1941,N_436,In_1334);
xor U1942 (N_1942,N_1083,N_1466);
nand U1943 (N_1943,In_1445,N_1351);
xnor U1944 (N_1944,N_864,N_353);
or U1945 (N_1945,In_436,N_515);
nand U1946 (N_1946,N_1376,In_1983);
nand U1947 (N_1947,N_831,N_1030);
or U1948 (N_1948,N_501,N_1082);
nand U1949 (N_1949,N_1301,N_944);
and U1950 (N_1950,N_1065,N_828);
nand U1951 (N_1951,N_1481,In_78);
nand U1952 (N_1952,N_1282,N_608);
and U1953 (N_1953,N_1205,N_1366);
nor U1954 (N_1954,In_308,N_1476);
or U1955 (N_1955,N_949,N_1404);
or U1956 (N_1956,N_1253,N_1335);
nor U1957 (N_1957,N_1153,In_1382);
nand U1958 (N_1958,N_1157,N_732);
or U1959 (N_1959,N_852,N_1190);
or U1960 (N_1960,N_1099,N_1113);
xnor U1961 (N_1961,N_1188,N_1245);
or U1962 (N_1962,N_1299,N_896);
xnor U1963 (N_1963,In_488,N_1493);
nor U1964 (N_1964,In_1133,N_1183);
or U1965 (N_1965,N_877,In_1071);
or U1966 (N_1966,N_1271,N_500);
nand U1967 (N_1967,N_961,In_2217);
or U1968 (N_1968,N_1031,In_382);
and U1969 (N_1969,N_858,N_1264);
nand U1970 (N_1970,N_1308,N_1460);
or U1971 (N_1971,In_2359,N_391);
and U1972 (N_1972,N_1248,N_1414);
xor U1973 (N_1973,N_569,N_1104);
and U1974 (N_1974,N_1462,N_803);
or U1975 (N_1975,N_678,In_737);
nand U1976 (N_1976,In_2434,N_138);
or U1977 (N_1977,N_1052,N_848);
and U1978 (N_1978,N_1388,N_1227);
nor U1979 (N_1979,In_1601,N_417);
xnor U1980 (N_1980,In_1284,N_804);
nand U1981 (N_1981,N_1364,N_1438);
xnor U1982 (N_1982,N_1303,In_693);
or U1983 (N_1983,N_1049,N_1196);
nand U1984 (N_1984,N_728,N_1439);
xnor U1985 (N_1985,N_646,N_1135);
nand U1986 (N_1986,N_63,N_1141);
or U1987 (N_1987,In_113,N_651);
or U1988 (N_1988,In_1498,N_281);
nand U1989 (N_1989,N_1471,N_48);
nor U1990 (N_1990,N_518,In_1243);
nor U1991 (N_1991,N_1004,N_1442);
nor U1992 (N_1992,N_1024,N_1069);
nor U1993 (N_1993,N_960,N_879);
nor U1994 (N_1994,N_1033,N_795);
or U1995 (N_1995,N_1102,N_1278);
xor U1996 (N_1996,In_144,N_538);
and U1997 (N_1997,In_1327,N_1251);
or U1998 (N_1998,N_525,N_1085);
xnor U1999 (N_1999,N_1447,N_1120);
nor U2000 (N_2000,N_1808,N_1549);
and U2001 (N_2001,N_1690,N_1575);
and U2002 (N_2002,N_1835,N_1977);
nor U2003 (N_2003,N_1743,N_1833);
or U2004 (N_2004,N_1726,N_1681);
and U2005 (N_2005,N_1997,N_1898);
nand U2006 (N_2006,N_1752,N_1962);
nand U2007 (N_2007,N_1713,N_1518);
nand U2008 (N_2008,N_1841,N_1736);
nand U2009 (N_2009,N_1846,N_1951);
nand U2010 (N_2010,N_1674,N_1954);
nor U2011 (N_2011,N_1545,N_1702);
xnor U2012 (N_2012,N_1783,N_1552);
nor U2013 (N_2013,N_1916,N_1853);
or U2014 (N_2014,N_1899,N_1836);
xor U2015 (N_2015,N_1934,N_1999);
and U2016 (N_2016,N_1857,N_1687);
nor U2017 (N_2017,N_1647,N_1597);
nor U2018 (N_2018,N_1861,N_1521);
and U2019 (N_2019,N_1500,N_1598);
nand U2020 (N_2020,N_1580,N_1856);
xnor U2021 (N_2021,N_1508,N_1721);
xnor U2022 (N_2022,N_1538,N_1534);
xor U2023 (N_2023,N_1769,N_1745);
or U2024 (N_2024,N_1582,N_1682);
nand U2025 (N_2025,N_1666,N_1848);
or U2026 (N_2026,N_1523,N_1659);
nand U2027 (N_2027,N_1531,N_1603);
nand U2028 (N_2028,N_1730,N_1617);
and U2029 (N_2029,N_1878,N_1512);
xor U2030 (N_2030,N_1821,N_1592);
and U2031 (N_2031,N_1505,N_1688);
nor U2032 (N_2032,N_1635,N_1664);
and U2033 (N_2033,N_1616,N_1636);
and U2034 (N_2034,N_1615,N_1718);
and U2035 (N_2035,N_1980,N_1527);
nand U2036 (N_2036,N_1988,N_1648);
and U2037 (N_2037,N_1594,N_1696);
xnor U2038 (N_2038,N_1849,N_1858);
xnor U2039 (N_2039,N_1969,N_1548);
xnor U2040 (N_2040,N_1756,N_1754);
xnor U2041 (N_2041,N_1517,N_1959);
or U2042 (N_2042,N_1778,N_1697);
xor U2043 (N_2043,N_1797,N_1850);
or U2044 (N_2044,N_1581,N_1896);
nand U2045 (N_2045,N_1680,N_1908);
and U2046 (N_2046,N_1672,N_1707);
nor U2047 (N_2047,N_1657,N_1873);
nor U2048 (N_2048,N_1976,N_1689);
nand U2049 (N_2049,N_1609,N_1871);
nand U2050 (N_2050,N_1734,N_1803);
nand U2051 (N_2051,N_1719,N_1723);
and U2052 (N_2052,N_1784,N_1795);
and U2053 (N_2053,N_1562,N_1760);
xor U2054 (N_2054,N_1619,N_1930);
xnor U2055 (N_2055,N_1968,N_1608);
nand U2056 (N_2056,N_1663,N_1600);
or U2057 (N_2057,N_1839,N_1502);
and U2058 (N_2058,N_1940,N_1987);
nor U2059 (N_2059,N_1771,N_1535);
or U2060 (N_2060,N_1879,N_1842);
or U2061 (N_2061,N_1624,N_1532);
or U2062 (N_2062,N_1605,N_1550);
or U2063 (N_2063,N_1679,N_1554);
or U2064 (N_2064,N_1904,N_1601);
and U2065 (N_2065,N_1780,N_1546);
xnor U2066 (N_2066,N_1553,N_1963);
nor U2067 (N_2067,N_1982,N_1642);
nand U2068 (N_2068,N_1639,N_1812);
xor U2069 (N_2069,N_1923,N_1995);
xor U2070 (N_2070,N_1870,N_1889);
or U2071 (N_2071,N_1887,N_1801);
nor U2072 (N_2072,N_1654,N_1753);
nor U2073 (N_2073,N_1641,N_1746);
or U2074 (N_2074,N_1526,N_1590);
nor U2075 (N_2075,N_1569,N_1727);
and U2076 (N_2076,N_1906,N_1935);
or U2077 (N_2077,N_1606,N_1573);
nor U2078 (N_2078,N_1984,N_1578);
xor U2079 (N_2079,N_1875,N_1970);
nor U2080 (N_2080,N_1832,N_1519);
nand U2081 (N_2081,N_1708,N_1911);
and U2082 (N_2082,N_1541,N_1621);
nor U2083 (N_2083,N_1514,N_1834);
and U2084 (N_2084,N_1540,N_1503);
and U2085 (N_2085,N_1924,N_1943);
nor U2086 (N_2086,N_1710,N_1890);
or U2087 (N_2087,N_1975,N_1577);
nand U2088 (N_2088,N_1670,N_1576);
or U2089 (N_2089,N_1915,N_1998);
nor U2090 (N_2090,N_1640,N_1974);
and U2091 (N_2091,N_1626,N_1838);
or U2092 (N_2092,N_1809,N_1757);
nor U2093 (N_2093,N_1794,N_1902);
nand U2094 (N_2094,N_1990,N_1806);
and U2095 (N_2095,N_1993,N_1955);
nand U2096 (N_2096,N_1564,N_1637);
nand U2097 (N_2097,N_1869,N_1933);
nor U2098 (N_2098,N_1817,N_1586);
and U2099 (N_2099,N_1884,N_1814);
xnor U2100 (N_2100,N_1767,N_1900);
or U2101 (N_2101,N_1936,N_1775);
and U2102 (N_2102,N_1633,N_1671);
and U2103 (N_2103,N_1630,N_1925);
nand U2104 (N_2104,N_1777,N_1952);
nor U2105 (N_2105,N_1851,N_1660);
or U2106 (N_2106,N_1650,N_1910);
xor U2107 (N_2107,N_1661,N_1766);
and U2108 (N_2108,N_1551,N_1728);
or U2109 (N_2109,N_1542,N_1927);
xor U2110 (N_2110,N_1613,N_1725);
and U2111 (N_2111,N_1826,N_1705);
or U2112 (N_2112,N_1986,N_1949);
and U2113 (N_2113,N_1882,N_1758);
nor U2114 (N_2114,N_1863,N_1926);
or U2115 (N_2115,N_1789,N_1932);
or U2116 (N_2116,N_1589,N_1942);
and U2117 (N_2117,N_1507,N_1610);
or U2118 (N_2118,N_1867,N_1764);
xor U2119 (N_2119,N_1894,N_1805);
nor U2120 (N_2120,N_1897,N_1929);
nor U2121 (N_2121,N_1845,N_1827);
or U2122 (N_2122,N_1628,N_1792);
nand U2123 (N_2123,N_1620,N_1691);
nor U2124 (N_2124,N_1996,N_1810);
nor U2125 (N_2125,N_1668,N_1669);
xor U2126 (N_2126,N_1945,N_1744);
or U2127 (N_2127,N_1825,N_1618);
xnor U2128 (N_2128,N_1868,N_1565);
or U2129 (N_2129,N_1732,N_1622);
nand U2130 (N_2130,N_1957,N_1556);
nand U2131 (N_2131,N_1676,N_1561);
xnor U2132 (N_2132,N_1574,N_1828);
xnor U2133 (N_2133,N_1706,N_1655);
or U2134 (N_2134,N_1729,N_1872);
nor U2135 (N_2135,N_1651,N_1599);
or U2136 (N_2136,N_1874,N_1847);
nor U2137 (N_2137,N_1860,N_1536);
or U2138 (N_2138,N_1678,N_1509);
xnor U2139 (N_2139,N_1749,N_1774);
or U2140 (N_2140,N_1737,N_1917);
nor U2141 (N_2141,N_1511,N_1765);
xnor U2142 (N_2142,N_1885,N_1629);
and U2143 (N_2143,N_1510,N_1716);
nand U2144 (N_2144,N_1859,N_1614);
and U2145 (N_2145,N_1739,N_1938);
xnor U2146 (N_2146,N_1520,N_1742);
xnor U2147 (N_2147,N_1722,N_1750);
nand U2148 (N_2148,N_1931,N_1593);
nor U2149 (N_2149,N_1584,N_1596);
nand U2150 (N_2150,N_1568,N_1971);
nor U2151 (N_2151,N_1829,N_1567);
xor U2152 (N_2152,N_1703,N_1903);
or U2153 (N_2153,N_1761,N_1956);
and U2154 (N_2154,N_1587,N_1816);
xnor U2155 (N_2155,N_1704,N_1886);
and U2156 (N_2156,N_1559,N_1768);
or U2157 (N_2157,N_1770,N_1937);
nor U2158 (N_2158,N_1570,N_1649);
nand U2159 (N_2159,N_1796,N_1607);
nor U2160 (N_2160,N_1572,N_1819);
xor U2161 (N_2161,N_1720,N_1985);
or U2162 (N_2162,N_1733,N_1524);
xor U2163 (N_2163,N_1731,N_1709);
nand U2164 (N_2164,N_1920,N_1843);
and U2165 (N_2165,N_1665,N_1790);
xnor U2166 (N_2166,N_1991,N_1791);
or U2167 (N_2167,N_1822,N_1960);
nor U2168 (N_2168,N_1712,N_1634);
and U2169 (N_2169,N_1529,N_1948);
nor U2170 (N_2170,N_1966,N_1675);
xor U2171 (N_2171,N_1504,N_1513);
and U2172 (N_2172,N_1862,N_1905);
or U2173 (N_2173,N_1939,N_1788);
xnor U2174 (N_2174,N_1714,N_1544);
xnor U2175 (N_2175,N_1683,N_1785);
nor U2176 (N_2176,N_1979,N_1588);
nor U2177 (N_2177,N_1953,N_1909);
nand U2178 (N_2178,N_1692,N_1965);
xor U2179 (N_2179,N_1646,N_1748);
and U2180 (N_2180,N_1698,N_1662);
or U2181 (N_2181,N_1560,N_1741);
xnor U2182 (N_2182,N_1891,N_1981);
xor U2183 (N_2183,N_1543,N_1928);
xor U2184 (N_2184,N_1611,N_1811);
xnor U2185 (N_2185,N_1978,N_1781);
xnor U2186 (N_2186,N_1989,N_1579);
nand U2187 (N_2187,N_1528,N_1824);
xnor U2188 (N_2188,N_1837,N_1912);
xor U2189 (N_2189,N_1667,N_1530);
xnor U2190 (N_2190,N_1763,N_1612);
or U2191 (N_2191,N_1913,N_1652);
nand U2192 (N_2192,N_1632,N_1844);
nor U2193 (N_2193,N_1516,N_1602);
xor U2194 (N_2194,N_1918,N_1786);
or U2195 (N_2195,N_1677,N_1604);
nor U2196 (N_2196,N_1645,N_1711);
xor U2197 (N_2197,N_1625,N_1571);
xor U2198 (N_2198,N_1525,N_1585);
and U2199 (N_2199,N_1701,N_1694);
and U2200 (N_2200,N_1595,N_1946);
nor U2201 (N_2201,N_1563,N_1653);
or U2202 (N_2202,N_1880,N_1643);
or U2203 (N_2203,N_1755,N_1695);
and U2204 (N_2204,N_1907,N_1967);
or U2205 (N_2205,N_1798,N_1501);
nand U2206 (N_2206,N_1994,N_1950);
and U2207 (N_2207,N_1804,N_1892);
xor U2208 (N_2208,N_1921,N_1793);
or U2209 (N_2209,N_1964,N_1762);
nand U2210 (N_2210,N_1877,N_1947);
xor U2211 (N_2211,N_1644,N_1865);
nor U2212 (N_2212,N_1591,N_1883);
nand U2213 (N_2213,N_1773,N_1700);
and U2214 (N_2214,N_1854,N_1866);
and U2215 (N_2215,N_1547,N_1972);
nor U2216 (N_2216,N_1717,N_1776);
xnor U2217 (N_2217,N_1914,N_1693);
and U2218 (N_2218,N_1901,N_1747);
nand U2219 (N_2219,N_1627,N_1631);
and U2220 (N_2220,N_1557,N_1855);
and U2221 (N_2221,N_1919,N_1961);
and U2222 (N_2222,N_1818,N_1506);
or U2223 (N_2223,N_1623,N_1735);
xnor U2224 (N_2224,N_1715,N_1782);
and U2225 (N_2225,N_1876,N_1815);
and U2226 (N_2226,N_1799,N_1992);
or U2227 (N_2227,N_1656,N_1820);
xor U2228 (N_2228,N_1537,N_1922);
xnor U2229 (N_2229,N_1759,N_1673);
nor U2230 (N_2230,N_1881,N_1888);
xor U2231 (N_2231,N_1539,N_1638);
nand U2232 (N_2232,N_1779,N_1558);
nand U2233 (N_2233,N_1852,N_1566);
nor U2234 (N_2234,N_1864,N_1813);
nor U2235 (N_2235,N_1807,N_1802);
or U2236 (N_2236,N_1973,N_1941);
xnor U2237 (N_2237,N_1555,N_1831);
and U2238 (N_2238,N_1515,N_1684);
or U2239 (N_2239,N_1583,N_1830);
nand U2240 (N_2240,N_1686,N_1800);
and U2241 (N_2241,N_1958,N_1944);
and U2242 (N_2242,N_1533,N_1738);
xnor U2243 (N_2243,N_1772,N_1840);
nand U2244 (N_2244,N_1751,N_1893);
or U2245 (N_2245,N_1522,N_1895);
nand U2246 (N_2246,N_1699,N_1823);
xnor U2247 (N_2247,N_1658,N_1983);
nand U2248 (N_2248,N_1787,N_1724);
xnor U2249 (N_2249,N_1740,N_1685);
and U2250 (N_2250,N_1619,N_1600);
and U2251 (N_2251,N_1503,N_1927);
or U2252 (N_2252,N_1503,N_1550);
nor U2253 (N_2253,N_1777,N_1681);
xnor U2254 (N_2254,N_1954,N_1725);
nor U2255 (N_2255,N_1939,N_1734);
and U2256 (N_2256,N_1837,N_1961);
or U2257 (N_2257,N_1687,N_1604);
nand U2258 (N_2258,N_1689,N_1595);
xnor U2259 (N_2259,N_1616,N_1554);
or U2260 (N_2260,N_1631,N_1910);
or U2261 (N_2261,N_1682,N_1867);
nor U2262 (N_2262,N_1762,N_1757);
or U2263 (N_2263,N_1971,N_1518);
nand U2264 (N_2264,N_1593,N_1554);
and U2265 (N_2265,N_1686,N_1949);
xor U2266 (N_2266,N_1659,N_1936);
and U2267 (N_2267,N_1508,N_1774);
xor U2268 (N_2268,N_1843,N_1553);
and U2269 (N_2269,N_1802,N_1862);
or U2270 (N_2270,N_1880,N_1915);
xnor U2271 (N_2271,N_1888,N_1603);
and U2272 (N_2272,N_1647,N_1782);
nor U2273 (N_2273,N_1947,N_1567);
and U2274 (N_2274,N_1647,N_1798);
nand U2275 (N_2275,N_1999,N_1575);
nand U2276 (N_2276,N_1565,N_1712);
or U2277 (N_2277,N_1564,N_1726);
or U2278 (N_2278,N_1548,N_1584);
and U2279 (N_2279,N_1607,N_1857);
nor U2280 (N_2280,N_1937,N_1724);
nand U2281 (N_2281,N_1945,N_1704);
or U2282 (N_2282,N_1906,N_1736);
xnor U2283 (N_2283,N_1940,N_1787);
nand U2284 (N_2284,N_1539,N_1744);
or U2285 (N_2285,N_1609,N_1652);
nor U2286 (N_2286,N_1961,N_1584);
xnor U2287 (N_2287,N_1517,N_1821);
xnor U2288 (N_2288,N_1942,N_1698);
or U2289 (N_2289,N_1915,N_1740);
or U2290 (N_2290,N_1551,N_1970);
nand U2291 (N_2291,N_1762,N_1989);
nor U2292 (N_2292,N_1539,N_1684);
and U2293 (N_2293,N_1901,N_1762);
or U2294 (N_2294,N_1911,N_1795);
xor U2295 (N_2295,N_1838,N_1565);
nor U2296 (N_2296,N_1999,N_1606);
nand U2297 (N_2297,N_1802,N_1546);
xor U2298 (N_2298,N_1845,N_1551);
or U2299 (N_2299,N_1798,N_1863);
or U2300 (N_2300,N_1855,N_1937);
or U2301 (N_2301,N_1850,N_1781);
and U2302 (N_2302,N_1880,N_1635);
or U2303 (N_2303,N_1840,N_1966);
xnor U2304 (N_2304,N_1563,N_1559);
nor U2305 (N_2305,N_1575,N_1508);
or U2306 (N_2306,N_1777,N_1707);
or U2307 (N_2307,N_1655,N_1578);
or U2308 (N_2308,N_1545,N_1874);
xor U2309 (N_2309,N_1573,N_1545);
xnor U2310 (N_2310,N_1859,N_1646);
nand U2311 (N_2311,N_1876,N_1854);
nand U2312 (N_2312,N_1731,N_1930);
xor U2313 (N_2313,N_1555,N_1563);
nand U2314 (N_2314,N_1674,N_1807);
or U2315 (N_2315,N_1858,N_1769);
nor U2316 (N_2316,N_1873,N_1807);
nand U2317 (N_2317,N_1614,N_1919);
nor U2318 (N_2318,N_1587,N_1537);
or U2319 (N_2319,N_1647,N_1964);
and U2320 (N_2320,N_1812,N_1553);
or U2321 (N_2321,N_1858,N_1915);
or U2322 (N_2322,N_1820,N_1934);
nor U2323 (N_2323,N_1522,N_1935);
nand U2324 (N_2324,N_1841,N_1681);
or U2325 (N_2325,N_1984,N_1847);
nand U2326 (N_2326,N_1934,N_1654);
xor U2327 (N_2327,N_1941,N_1883);
nand U2328 (N_2328,N_1747,N_1705);
xnor U2329 (N_2329,N_1605,N_1787);
nor U2330 (N_2330,N_1785,N_1950);
and U2331 (N_2331,N_1500,N_1652);
nor U2332 (N_2332,N_1640,N_1711);
and U2333 (N_2333,N_1745,N_1913);
xnor U2334 (N_2334,N_1742,N_1675);
nor U2335 (N_2335,N_1819,N_1504);
and U2336 (N_2336,N_1673,N_1940);
nand U2337 (N_2337,N_1787,N_1817);
nor U2338 (N_2338,N_1665,N_1514);
nand U2339 (N_2339,N_1874,N_1975);
nor U2340 (N_2340,N_1595,N_1724);
xor U2341 (N_2341,N_1841,N_1633);
xor U2342 (N_2342,N_1689,N_1985);
and U2343 (N_2343,N_1786,N_1916);
xnor U2344 (N_2344,N_1618,N_1753);
nand U2345 (N_2345,N_1583,N_1738);
nand U2346 (N_2346,N_1738,N_1893);
and U2347 (N_2347,N_1562,N_1973);
xnor U2348 (N_2348,N_1665,N_1809);
or U2349 (N_2349,N_1942,N_1947);
nor U2350 (N_2350,N_1793,N_1890);
nand U2351 (N_2351,N_1872,N_1967);
nor U2352 (N_2352,N_1572,N_1713);
nand U2353 (N_2353,N_1985,N_1916);
xor U2354 (N_2354,N_1937,N_1760);
nand U2355 (N_2355,N_1610,N_1901);
xnor U2356 (N_2356,N_1655,N_1798);
nand U2357 (N_2357,N_1864,N_1700);
and U2358 (N_2358,N_1883,N_1933);
and U2359 (N_2359,N_1543,N_1766);
nand U2360 (N_2360,N_1968,N_1785);
or U2361 (N_2361,N_1645,N_1740);
and U2362 (N_2362,N_1899,N_1733);
or U2363 (N_2363,N_1536,N_1730);
and U2364 (N_2364,N_1858,N_1563);
and U2365 (N_2365,N_1528,N_1501);
nand U2366 (N_2366,N_1628,N_1713);
nor U2367 (N_2367,N_1906,N_1516);
or U2368 (N_2368,N_1544,N_1831);
nor U2369 (N_2369,N_1535,N_1916);
xor U2370 (N_2370,N_1925,N_1930);
or U2371 (N_2371,N_1886,N_1601);
or U2372 (N_2372,N_1607,N_1653);
and U2373 (N_2373,N_1518,N_1863);
or U2374 (N_2374,N_1731,N_1572);
xnor U2375 (N_2375,N_1545,N_1994);
nor U2376 (N_2376,N_1768,N_1503);
or U2377 (N_2377,N_1718,N_1797);
nand U2378 (N_2378,N_1529,N_1838);
or U2379 (N_2379,N_1500,N_1924);
xor U2380 (N_2380,N_1600,N_1612);
and U2381 (N_2381,N_1750,N_1810);
and U2382 (N_2382,N_1873,N_1633);
xnor U2383 (N_2383,N_1918,N_1835);
and U2384 (N_2384,N_1589,N_1601);
xor U2385 (N_2385,N_1833,N_1816);
nor U2386 (N_2386,N_1588,N_1621);
or U2387 (N_2387,N_1683,N_1751);
xnor U2388 (N_2388,N_1538,N_1612);
xor U2389 (N_2389,N_1702,N_1806);
xor U2390 (N_2390,N_1568,N_1923);
or U2391 (N_2391,N_1532,N_1812);
nand U2392 (N_2392,N_1508,N_1683);
nand U2393 (N_2393,N_1886,N_1664);
and U2394 (N_2394,N_1624,N_1719);
nor U2395 (N_2395,N_1686,N_1805);
nor U2396 (N_2396,N_1508,N_1896);
and U2397 (N_2397,N_1523,N_1956);
nand U2398 (N_2398,N_1628,N_1730);
nor U2399 (N_2399,N_1810,N_1500);
or U2400 (N_2400,N_1929,N_1971);
nand U2401 (N_2401,N_1638,N_1555);
nor U2402 (N_2402,N_1799,N_1741);
nand U2403 (N_2403,N_1942,N_1814);
and U2404 (N_2404,N_1869,N_1891);
nand U2405 (N_2405,N_1806,N_1507);
and U2406 (N_2406,N_1992,N_1964);
nor U2407 (N_2407,N_1806,N_1794);
xnor U2408 (N_2408,N_1899,N_1734);
or U2409 (N_2409,N_1637,N_1532);
xnor U2410 (N_2410,N_1879,N_1503);
xor U2411 (N_2411,N_1990,N_1985);
or U2412 (N_2412,N_1936,N_1538);
nor U2413 (N_2413,N_1776,N_1730);
nand U2414 (N_2414,N_1658,N_1668);
nand U2415 (N_2415,N_1801,N_1947);
xor U2416 (N_2416,N_1955,N_1829);
xor U2417 (N_2417,N_1953,N_1558);
or U2418 (N_2418,N_1765,N_1801);
nor U2419 (N_2419,N_1794,N_1787);
or U2420 (N_2420,N_1673,N_1898);
or U2421 (N_2421,N_1731,N_1509);
xnor U2422 (N_2422,N_1670,N_1667);
nand U2423 (N_2423,N_1844,N_1583);
and U2424 (N_2424,N_1757,N_1947);
nor U2425 (N_2425,N_1763,N_1520);
xnor U2426 (N_2426,N_1876,N_1829);
nand U2427 (N_2427,N_1788,N_1770);
nor U2428 (N_2428,N_1631,N_1883);
or U2429 (N_2429,N_1985,N_1511);
nand U2430 (N_2430,N_1735,N_1507);
or U2431 (N_2431,N_1823,N_1781);
and U2432 (N_2432,N_1755,N_1661);
nand U2433 (N_2433,N_1654,N_1798);
nand U2434 (N_2434,N_1705,N_1827);
nand U2435 (N_2435,N_1585,N_1714);
and U2436 (N_2436,N_1999,N_1859);
xor U2437 (N_2437,N_1847,N_1543);
or U2438 (N_2438,N_1760,N_1658);
nor U2439 (N_2439,N_1850,N_1958);
or U2440 (N_2440,N_1670,N_1580);
or U2441 (N_2441,N_1891,N_1944);
and U2442 (N_2442,N_1627,N_1700);
xnor U2443 (N_2443,N_1955,N_1956);
xor U2444 (N_2444,N_1986,N_1889);
nand U2445 (N_2445,N_1643,N_1877);
and U2446 (N_2446,N_1530,N_1816);
or U2447 (N_2447,N_1906,N_1653);
and U2448 (N_2448,N_1662,N_1919);
nand U2449 (N_2449,N_1848,N_1654);
and U2450 (N_2450,N_1968,N_1584);
or U2451 (N_2451,N_1703,N_1924);
nor U2452 (N_2452,N_1947,N_1772);
or U2453 (N_2453,N_1687,N_1931);
nor U2454 (N_2454,N_1800,N_1963);
xor U2455 (N_2455,N_1922,N_1628);
and U2456 (N_2456,N_1999,N_1598);
nand U2457 (N_2457,N_1864,N_1830);
or U2458 (N_2458,N_1668,N_1506);
or U2459 (N_2459,N_1804,N_1690);
xnor U2460 (N_2460,N_1686,N_1542);
or U2461 (N_2461,N_1675,N_1567);
or U2462 (N_2462,N_1808,N_1708);
xnor U2463 (N_2463,N_1502,N_1844);
and U2464 (N_2464,N_1718,N_1990);
nor U2465 (N_2465,N_1688,N_1778);
xor U2466 (N_2466,N_1592,N_1621);
nor U2467 (N_2467,N_1772,N_1742);
nand U2468 (N_2468,N_1698,N_1877);
and U2469 (N_2469,N_1760,N_1762);
xnor U2470 (N_2470,N_1750,N_1964);
xnor U2471 (N_2471,N_1827,N_1895);
nand U2472 (N_2472,N_1856,N_1548);
nor U2473 (N_2473,N_1752,N_1519);
nand U2474 (N_2474,N_1614,N_1567);
or U2475 (N_2475,N_1835,N_1931);
and U2476 (N_2476,N_1622,N_1730);
xor U2477 (N_2477,N_1883,N_1836);
or U2478 (N_2478,N_1948,N_1532);
xor U2479 (N_2479,N_1561,N_1821);
or U2480 (N_2480,N_1596,N_1706);
or U2481 (N_2481,N_1897,N_1985);
nor U2482 (N_2482,N_1630,N_1565);
xnor U2483 (N_2483,N_1642,N_1637);
nand U2484 (N_2484,N_1585,N_1514);
and U2485 (N_2485,N_1838,N_1730);
xor U2486 (N_2486,N_1600,N_1884);
nand U2487 (N_2487,N_1903,N_1900);
xor U2488 (N_2488,N_1515,N_1524);
or U2489 (N_2489,N_1841,N_1973);
xor U2490 (N_2490,N_1516,N_1691);
nor U2491 (N_2491,N_1659,N_1571);
nand U2492 (N_2492,N_1988,N_1622);
nand U2493 (N_2493,N_1885,N_1735);
and U2494 (N_2494,N_1888,N_1773);
nand U2495 (N_2495,N_1604,N_1606);
nor U2496 (N_2496,N_1959,N_1894);
nor U2497 (N_2497,N_1964,N_1546);
nand U2498 (N_2498,N_1821,N_1853);
nand U2499 (N_2499,N_1505,N_1603);
nand U2500 (N_2500,N_2207,N_2223);
and U2501 (N_2501,N_2079,N_2123);
nor U2502 (N_2502,N_2346,N_2382);
nand U2503 (N_2503,N_2366,N_2029);
nor U2504 (N_2504,N_2217,N_2280);
nor U2505 (N_2505,N_2352,N_2497);
nor U2506 (N_2506,N_2394,N_2047);
nor U2507 (N_2507,N_2290,N_2025);
xnor U2508 (N_2508,N_2036,N_2057);
nand U2509 (N_2509,N_2181,N_2289);
nand U2510 (N_2510,N_2337,N_2372);
or U2511 (N_2511,N_2271,N_2420);
nor U2512 (N_2512,N_2315,N_2134);
xnor U2513 (N_2513,N_2208,N_2215);
nor U2514 (N_2514,N_2474,N_2451);
and U2515 (N_2515,N_2182,N_2388);
nor U2516 (N_2516,N_2068,N_2204);
and U2517 (N_2517,N_2026,N_2233);
xor U2518 (N_2518,N_2450,N_2375);
or U2519 (N_2519,N_2058,N_2359);
and U2520 (N_2520,N_2381,N_2065);
nor U2521 (N_2521,N_2228,N_2463);
or U2522 (N_2522,N_2019,N_2066);
xnor U2523 (N_2523,N_2370,N_2010);
nor U2524 (N_2524,N_2041,N_2246);
nor U2525 (N_2525,N_2301,N_2384);
nand U2526 (N_2526,N_2368,N_2465);
or U2527 (N_2527,N_2303,N_2383);
or U2528 (N_2528,N_2177,N_2356);
nand U2529 (N_2529,N_2224,N_2109);
and U2530 (N_2530,N_2250,N_2050);
or U2531 (N_2531,N_2415,N_2358);
nor U2532 (N_2532,N_2138,N_2434);
and U2533 (N_2533,N_2159,N_2401);
nor U2534 (N_2534,N_2333,N_2400);
xor U2535 (N_2535,N_2437,N_2328);
and U2536 (N_2536,N_2425,N_2034);
xor U2537 (N_2537,N_2214,N_2476);
or U2538 (N_2538,N_2110,N_2202);
nand U2539 (N_2539,N_2220,N_2410);
and U2540 (N_2540,N_2418,N_2431);
and U2541 (N_2541,N_2113,N_2348);
xor U2542 (N_2542,N_2236,N_2162);
or U2543 (N_2543,N_2049,N_2374);
xor U2544 (N_2544,N_2169,N_2242);
nor U2545 (N_2545,N_2335,N_2069);
xnor U2546 (N_2546,N_2496,N_2260);
nor U2547 (N_2547,N_2408,N_2080);
nor U2548 (N_2548,N_2402,N_2037);
and U2549 (N_2549,N_2287,N_2184);
nand U2550 (N_2550,N_2227,N_2221);
nor U2551 (N_2551,N_2145,N_2442);
xor U2552 (N_2552,N_2435,N_2413);
nand U2553 (N_2553,N_2040,N_2320);
nand U2554 (N_2554,N_2340,N_2059);
xnor U2555 (N_2555,N_2300,N_2281);
and U2556 (N_2556,N_2183,N_2063);
and U2557 (N_2557,N_2179,N_2457);
nand U2558 (N_2558,N_2210,N_2475);
xnor U2559 (N_2559,N_2255,N_2393);
nand U2560 (N_2560,N_2441,N_2129);
xor U2561 (N_2561,N_2015,N_2114);
xnor U2562 (N_2562,N_2060,N_2193);
xnor U2563 (N_2563,N_2272,N_2211);
nand U2564 (N_2564,N_2254,N_2445);
and U2565 (N_2565,N_2455,N_2460);
xor U2566 (N_2566,N_2318,N_2095);
or U2567 (N_2567,N_2051,N_2013);
xnor U2568 (N_2568,N_2175,N_2288);
nand U2569 (N_2569,N_2354,N_2226);
or U2570 (N_2570,N_2365,N_2351);
nor U2571 (N_2571,N_2297,N_2155);
nand U2572 (N_2572,N_2122,N_2126);
nand U2573 (N_2573,N_2212,N_2489);
nor U2574 (N_2574,N_2192,N_2453);
and U2575 (N_2575,N_2104,N_2349);
and U2576 (N_2576,N_2077,N_2235);
and U2577 (N_2577,N_2367,N_2230);
xor U2578 (N_2578,N_2231,N_2148);
xor U2579 (N_2579,N_2412,N_2006);
and U2580 (N_2580,N_2485,N_2433);
nand U2581 (N_2581,N_2152,N_2108);
and U2582 (N_2582,N_2482,N_2062);
xnor U2583 (N_2583,N_2116,N_2296);
nor U2584 (N_2584,N_2054,N_2088);
and U2585 (N_2585,N_2491,N_2127);
or U2586 (N_2586,N_2244,N_2343);
and U2587 (N_2587,N_2106,N_2407);
and U2588 (N_2588,N_2285,N_2310);
or U2589 (N_2589,N_2423,N_2143);
nor U2590 (N_2590,N_2461,N_2339);
or U2591 (N_2591,N_2016,N_2298);
nor U2592 (N_2592,N_2200,N_2133);
and U2593 (N_2593,N_2456,N_2305);
and U2594 (N_2594,N_2174,N_2444);
or U2595 (N_2595,N_2330,N_2416);
and U2596 (N_2596,N_2336,N_2101);
xnor U2597 (N_2597,N_2389,N_2279);
or U2598 (N_2598,N_2257,N_2486);
xor U2599 (N_2599,N_2203,N_2046);
and U2600 (N_2600,N_2276,N_2021);
nand U2601 (N_2601,N_2259,N_2308);
or U2602 (N_2602,N_2171,N_2406);
or U2603 (N_2603,N_2331,N_2076);
nor U2604 (N_2604,N_2136,N_2239);
nand U2605 (N_2605,N_2099,N_2332);
or U2606 (N_2606,N_2341,N_2316);
nand U2607 (N_2607,N_2107,N_2100);
nand U2608 (N_2608,N_2125,N_2170);
and U2609 (N_2609,N_2355,N_2185);
xnor U2610 (N_2610,N_2091,N_2199);
or U2611 (N_2611,N_2386,N_2467);
xor U2612 (N_2612,N_2197,N_2005);
and U2613 (N_2613,N_2111,N_2481);
or U2614 (N_2614,N_2168,N_2414);
xor U2615 (N_2615,N_2306,N_2253);
nand U2616 (N_2616,N_2241,N_2090);
nor U2617 (N_2617,N_2072,N_2020);
and U2618 (N_2618,N_2292,N_2395);
nor U2619 (N_2619,N_2422,N_2493);
nand U2620 (N_2620,N_2269,N_2478);
nand U2621 (N_2621,N_2030,N_2409);
nand U2622 (N_2622,N_2345,N_2466);
and U2623 (N_2623,N_2428,N_2229);
nand U2624 (N_2624,N_2373,N_2014);
xor U2625 (N_2625,N_2284,N_2448);
or U2626 (N_2626,N_2258,N_2377);
and U2627 (N_2627,N_2309,N_2243);
and U2628 (N_2628,N_2319,N_2151);
or U2629 (N_2629,N_2085,N_2167);
nand U2630 (N_2630,N_2024,N_2156);
or U2631 (N_2631,N_2130,N_2299);
nand U2632 (N_2632,N_2083,N_2484);
nand U2633 (N_2633,N_2446,N_2237);
or U2634 (N_2634,N_2492,N_2487);
nor U2635 (N_2635,N_2018,N_2342);
xor U2636 (N_2636,N_2454,N_2031);
nand U2637 (N_2637,N_2061,N_2124);
or U2638 (N_2638,N_2118,N_2096);
nand U2639 (N_2639,N_2247,N_2173);
and U2640 (N_2640,N_2273,N_2004);
xor U2641 (N_2641,N_2186,N_2153);
nor U2642 (N_2642,N_2261,N_2039);
nor U2643 (N_2643,N_2089,N_2398);
nor U2644 (N_2644,N_2424,N_2074);
and U2645 (N_2645,N_2141,N_2033);
or U2646 (N_2646,N_2321,N_2283);
xnor U2647 (N_2647,N_2387,N_2234);
nor U2648 (N_2648,N_2105,N_2043);
nand U2649 (N_2649,N_2144,N_2286);
and U2650 (N_2650,N_2135,N_2295);
xnor U2651 (N_2651,N_2147,N_2201);
nor U2652 (N_2652,N_2225,N_2073);
nor U2653 (N_2653,N_2396,N_2098);
nand U2654 (N_2654,N_2190,N_2092);
xor U2655 (N_2655,N_2007,N_2205);
or U2656 (N_2656,N_2371,N_2364);
or U2657 (N_2657,N_2084,N_2291);
xor U2658 (N_2658,N_2275,N_2160);
and U2659 (N_2659,N_2322,N_2178);
nor U2660 (N_2660,N_2274,N_2003);
nand U2661 (N_2661,N_2112,N_2344);
xnor U2662 (N_2662,N_2302,N_2067);
and U2663 (N_2663,N_2154,N_2468);
and U2664 (N_2664,N_2120,N_2103);
xnor U2665 (N_2665,N_2480,N_2458);
and U2666 (N_2666,N_2464,N_2027);
nor U2667 (N_2667,N_2002,N_2044);
nor U2668 (N_2668,N_2232,N_2093);
and U2669 (N_2669,N_2188,N_2449);
nor U2670 (N_2670,N_2000,N_2161);
xor U2671 (N_2671,N_2042,N_2350);
or U2672 (N_2672,N_2035,N_2140);
nand U2673 (N_2673,N_2198,N_2459);
nand U2674 (N_2674,N_2439,N_2317);
nor U2675 (N_2675,N_2334,N_2128);
nor U2676 (N_2676,N_2209,N_2150);
xor U2677 (N_2677,N_2252,N_2157);
and U2678 (N_2678,N_2379,N_2189);
nand U2679 (N_2679,N_2432,N_2472);
nand U2680 (N_2680,N_2477,N_2495);
xnor U2681 (N_2681,N_2078,N_2429);
nor U2682 (N_2682,N_2360,N_2403);
xnor U2683 (N_2683,N_2086,N_2045);
and U2684 (N_2684,N_2251,N_2264);
or U2685 (N_2685,N_2294,N_2277);
xnor U2686 (N_2686,N_2163,N_2430);
and U2687 (N_2687,N_2385,N_2158);
and U2688 (N_2688,N_2440,N_2146);
nand U2689 (N_2689,N_2070,N_2488);
nor U2690 (N_2690,N_2421,N_2325);
or U2691 (N_2691,N_2195,N_2038);
nor U2692 (N_2692,N_2053,N_2329);
and U2693 (N_2693,N_2139,N_2048);
nand U2694 (N_2694,N_2056,N_2149);
and U2695 (N_2695,N_2075,N_2378);
or U2696 (N_2696,N_2001,N_2417);
and U2697 (N_2697,N_2304,N_2311);
nand U2698 (N_2698,N_2165,N_2017);
or U2699 (N_2699,N_2248,N_2249);
nor U2700 (N_2700,N_2405,N_2240);
nand U2701 (N_2701,N_2119,N_2102);
xor U2702 (N_2702,N_2347,N_2052);
xor U2703 (N_2703,N_2397,N_2473);
xor U2704 (N_2704,N_2266,N_2022);
xnor U2705 (N_2705,N_2121,N_2191);
nand U2706 (N_2706,N_2187,N_2363);
nand U2707 (N_2707,N_2282,N_2064);
and U2708 (N_2708,N_2267,N_2082);
nand U2709 (N_2709,N_2314,N_2219);
xnor U2710 (N_2710,N_2426,N_2452);
and U2711 (N_2711,N_2206,N_2362);
and U2712 (N_2712,N_2357,N_2399);
and U2713 (N_2713,N_2131,N_2307);
xor U2714 (N_2714,N_2238,N_2443);
nor U2715 (N_2715,N_2256,N_2166);
xnor U2716 (N_2716,N_2479,N_2419);
xnor U2717 (N_2717,N_2216,N_2380);
xnor U2718 (N_2718,N_2268,N_2471);
or U2719 (N_2719,N_2499,N_2222);
nand U2720 (N_2720,N_2012,N_2218);
nor U2721 (N_2721,N_2494,N_2115);
nand U2722 (N_2722,N_2498,N_2097);
or U2723 (N_2723,N_2245,N_2194);
nor U2724 (N_2724,N_2390,N_2132);
and U2725 (N_2725,N_2324,N_2376);
nor U2726 (N_2726,N_2353,N_2263);
nor U2727 (N_2727,N_2023,N_2081);
nor U2728 (N_2728,N_2213,N_2164);
and U2729 (N_2729,N_2447,N_2176);
nand U2730 (N_2730,N_2323,N_2071);
and U2731 (N_2731,N_2262,N_2436);
nand U2732 (N_2732,N_2327,N_2338);
nor U2733 (N_2733,N_2391,N_2427);
xor U2734 (N_2734,N_2392,N_2404);
and U2735 (N_2735,N_2278,N_2438);
nor U2736 (N_2736,N_2313,N_2326);
and U2737 (N_2737,N_2369,N_2172);
and U2738 (N_2738,N_2411,N_2483);
xnor U2739 (N_2739,N_2055,N_2469);
xor U2740 (N_2740,N_2490,N_2462);
nor U2741 (N_2741,N_2270,N_2137);
or U2742 (N_2742,N_2011,N_2094);
and U2743 (N_2743,N_2032,N_2180);
or U2744 (N_2744,N_2142,N_2361);
xnor U2745 (N_2745,N_2087,N_2312);
nor U2746 (N_2746,N_2196,N_2008);
and U2747 (N_2747,N_2028,N_2293);
and U2748 (N_2748,N_2470,N_2265);
nor U2749 (N_2749,N_2009,N_2117);
xor U2750 (N_2750,N_2013,N_2466);
and U2751 (N_2751,N_2028,N_2143);
xnor U2752 (N_2752,N_2399,N_2320);
and U2753 (N_2753,N_2360,N_2213);
and U2754 (N_2754,N_2014,N_2257);
or U2755 (N_2755,N_2182,N_2330);
and U2756 (N_2756,N_2096,N_2240);
nor U2757 (N_2757,N_2404,N_2039);
and U2758 (N_2758,N_2048,N_2065);
or U2759 (N_2759,N_2377,N_2065);
or U2760 (N_2760,N_2154,N_2447);
nor U2761 (N_2761,N_2129,N_2256);
xor U2762 (N_2762,N_2111,N_2325);
or U2763 (N_2763,N_2082,N_2400);
nand U2764 (N_2764,N_2181,N_2478);
or U2765 (N_2765,N_2357,N_2457);
or U2766 (N_2766,N_2177,N_2209);
nor U2767 (N_2767,N_2178,N_2436);
xnor U2768 (N_2768,N_2429,N_2064);
xor U2769 (N_2769,N_2290,N_2263);
nand U2770 (N_2770,N_2192,N_2327);
xor U2771 (N_2771,N_2441,N_2377);
xnor U2772 (N_2772,N_2060,N_2353);
xnor U2773 (N_2773,N_2446,N_2480);
and U2774 (N_2774,N_2488,N_2076);
or U2775 (N_2775,N_2425,N_2339);
xor U2776 (N_2776,N_2100,N_2315);
or U2777 (N_2777,N_2289,N_2303);
and U2778 (N_2778,N_2086,N_2020);
and U2779 (N_2779,N_2385,N_2005);
nor U2780 (N_2780,N_2360,N_2382);
and U2781 (N_2781,N_2064,N_2483);
nor U2782 (N_2782,N_2055,N_2260);
nand U2783 (N_2783,N_2380,N_2147);
nand U2784 (N_2784,N_2191,N_2145);
and U2785 (N_2785,N_2038,N_2406);
xnor U2786 (N_2786,N_2246,N_2471);
nor U2787 (N_2787,N_2313,N_2474);
xnor U2788 (N_2788,N_2293,N_2436);
xnor U2789 (N_2789,N_2337,N_2102);
xor U2790 (N_2790,N_2282,N_2469);
xor U2791 (N_2791,N_2030,N_2285);
and U2792 (N_2792,N_2121,N_2188);
or U2793 (N_2793,N_2127,N_2023);
xor U2794 (N_2794,N_2232,N_2285);
or U2795 (N_2795,N_2369,N_2435);
and U2796 (N_2796,N_2388,N_2059);
nor U2797 (N_2797,N_2434,N_2191);
nand U2798 (N_2798,N_2296,N_2096);
and U2799 (N_2799,N_2216,N_2381);
nor U2800 (N_2800,N_2036,N_2206);
nand U2801 (N_2801,N_2391,N_2422);
nand U2802 (N_2802,N_2016,N_2418);
nor U2803 (N_2803,N_2419,N_2262);
and U2804 (N_2804,N_2089,N_2024);
nor U2805 (N_2805,N_2067,N_2322);
xnor U2806 (N_2806,N_2409,N_2391);
or U2807 (N_2807,N_2144,N_2238);
and U2808 (N_2808,N_2227,N_2356);
and U2809 (N_2809,N_2142,N_2482);
or U2810 (N_2810,N_2268,N_2151);
nor U2811 (N_2811,N_2051,N_2169);
nor U2812 (N_2812,N_2236,N_2361);
or U2813 (N_2813,N_2348,N_2457);
xor U2814 (N_2814,N_2205,N_2321);
or U2815 (N_2815,N_2184,N_2109);
and U2816 (N_2816,N_2221,N_2351);
or U2817 (N_2817,N_2395,N_2242);
and U2818 (N_2818,N_2350,N_2060);
or U2819 (N_2819,N_2209,N_2074);
nand U2820 (N_2820,N_2066,N_2102);
xnor U2821 (N_2821,N_2268,N_2266);
nor U2822 (N_2822,N_2304,N_2209);
and U2823 (N_2823,N_2370,N_2020);
xor U2824 (N_2824,N_2248,N_2350);
or U2825 (N_2825,N_2095,N_2039);
nand U2826 (N_2826,N_2046,N_2072);
or U2827 (N_2827,N_2288,N_2436);
nand U2828 (N_2828,N_2112,N_2441);
nor U2829 (N_2829,N_2204,N_2198);
or U2830 (N_2830,N_2321,N_2231);
xnor U2831 (N_2831,N_2410,N_2390);
xor U2832 (N_2832,N_2376,N_2430);
xor U2833 (N_2833,N_2357,N_2028);
nand U2834 (N_2834,N_2301,N_2349);
nand U2835 (N_2835,N_2359,N_2029);
nand U2836 (N_2836,N_2377,N_2411);
or U2837 (N_2837,N_2484,N_2164);
xor U2838 (N_2838,N_2115,N_2112);
xnor U2839 (N_2839,N_2467,N_2097);
nand U2840 (N_2840,N_2497,N_2418);
and U2841 (N_2841,N_2299,N_2037);
nor U2842 (N_2842,N_2366,N_2484);
or U2843 (N_2843,N_2326,N_2232);
or U2844 (N_2844,N_2154,N_2183);
xor U2845 (N_2845,N_2484,N_2234);
nand U2846 (N_2846,N_2476,N_2088);
nor U2847 (N_2847,N_2151,N_2489);
and U2848 (N_2848,N_2389,N_2139);
or U2849 (N_2849,N_2178,N_2392);
nand U2850 (N_2850,N_2240,N_2327);
xnor U2851 (N_2851,N_2336,N_2003);
and U2852 (N_2852,N_2008,N_2422);
nor U2853 (N_2853,N_2101,N_2255);
or U2854 (N_2854,N_2202,N_2077);
nand U2855 (N_2855,N_2188,N_2158);
and U2856 (N_2856,N_2237,N_2449);
and U2857 (N_2857,N_2209,N_2171);
or U2858 (N_2858,N_2112,N_2085);
nand U2859 (N_2859,N_2230,N_2100);
or U2860 (N_2860,N_2470,N_2131);
or U2861 (N_2861,N_2248,N_2348);
nor U2862 (N_2862,N_2488,N_2485);
xor U2863 (N_2863,N_2115,N_2026);
nor U2864 (N_2864,N_2177,N_2384);
nor U2865 (N_2865,N_2136,N_2032);
or U2866 (N_2866,N_2476,N_2042);
nor U2867 (N_2867,N_2295,N_2364);
nor U2868 (N_2868,N_2381,N_2446);
xnor U2869 (N_2869,N_2053,N_2398);
and U2870 (N_2870,N_2465,N_2041);
and U2871 (N_2871,N_2486,N_2262);
nor U2872 (N_2872,N_2335,N_2113);
nand U2873 (N_2873,N_2232,N_2177);
or U2874 (N_2874,N_2259,N_2495);
and U2875 (N_2875,N_2190,N_2363);
nand U2876 (N_2876,N_2402,N_2490);
xnor U2877 (N_2877,N_2469,N_2121);
or U2878 (N_2878,N_2394,N_2122);
or U2879 (N_2879,N_2196,N_2028);
nor U2880 (N_2880,N_2136,N_2195);
or U2881 (N_2881,N_2378,N_2076);
and U2882 (N_2882,N_2133,N_2390);
xor U2883 (N_2883,N_2085,N_2065);
nor U2884 (N_2884,N_2256,N_2435);
nand U2885 (N_2885,N_2422,N_2299);
xnor U2886 (N_2886,N_2238,N_2339);
xor U2887 (N_2887,N_2317,N_2142);
xor U2888 (N_2888,N_2019,N_2098);
xnor U2889 (N_2889,N_2210,N_2428);
or U2890 (N_2890,N_2239,N_2213);
or U2891 (N_2891,N_2287,N_2122);
xnor U2892 (N_2892,N_2177,N_2343);
or U2893 (N_2893,N_2131,N_2431);
xnor U2894 (N_2894,N_2106,N_2499);
nor U2895 (N_2895,N_2128,N_2189);
xnor U2896 (N_2896,N_2309,N_2017);
nor U2897 (N_2897,N_2379,N_2162);
nor U2898 (N_2898,N_2004,N_2475);
xor U2899 (N_2899,N_2179,N_2095);
and U2900 (N_2900,N_2184,N_2416);
and U2901 (N_2901,N_2445,N_2207);
and U2902 (N_2902,N_2173,N_2378);
and U2903 (N_2903,N_2379,N_2448);
nand U2904 (N_2904,N_2090,N_2405);
xor U2905 (N_2905,N_2278,N_2174);
xnor U2906 (N_2906,N_2131,N_2493);
or U2907 (N_2907,N_2114,N_2085);
nor U2908 (N_2908,N_2064,N_2216);
xor U2909 (N_2909,N_2088,N_2052);
nand U2910 (N_2910,N_2069,N_2353);
and U2911 (N_2911,N_2192,N_2109);
nand U2912 (N_2912,N_2496,N_2429);
xor U2913 (N_2913,N_2244,N_2088);
xnor U2914 (N_2914,N_2389,N_2186);
xnor U2915 (N_2915,N_2016,N_2165);
nor U2916 (N_2916,N_2358,N_2418);
xnor U2917 (N_2917,N_2087,N_2008);
xnor U2918 (N_2918,N_2277,N_2479);
and U2919 (N_2919,N_2342,N_2068);
nor U2920 (N_2920,N_2103,N_2383);
and U2921 (N_2921,N_2318,N_2199);
xnor U2922 (N_2922,N_2161,N_2404);
or U2923 (N_2923,N_2147,N_2362);
nand U2924 (N_2924,N_2161,N_2135);
nor U2925 (N_2925,N_2440,N_2367);
or U2926 (N_2926,N_2321,N_2461);
or U2927 (N_2927,N_2026,N_2495);
and U2928 (N_2928,N_2208,N_2495);
and U2929 (N_2929,N_2191,N_2182);
nor U2930 (N_2930,N_2192,N_2039);
nand U2931 (N_2931,N_2332,N_2246);
or U2932 (N_2932,N_2160,N_2068);
xor U2933 (N_2933,N_2429,N_2010);
xnor U2934 (N_2934,N_2199,N_2377);
and U2935 (N_2935,N_2382,N_2494);
nand U2936 (N_2936,N_2438,N_2325);
and U2937 (N_2937,N_2344,N_2393);
and U2938 (N_2938,N_2050,N_2219);
xor U2939 (N_2939,N_2266,N_2498);
and U2940 (N_2940,N_2324,N_2066);
and U2941 (N_2941,N_2220,N_2218);
nand U2942 (N_2942,N_2216,N_2279);
nor U2943 (N_2943,N_2116,N_2312);
xnor U2944 (N_2944,N_2097,N_2480);
nand U2945 (N_2945,N_2267,N_2174);
or U2946 (N_2946,N_2343,N_2438);
nand U2947 (N_2947,N_2434,N_2301);
or U2948 (N_2948,N_2209,N_2323);
xor U2949 (N_2949,N_2049,N_2250);
xnor U2950 (N_2950,N_2144,N_2156);
xnor U2951 (N_2951,N_2239,N_2267);
nand U2952 (N_2952,N_2099,N_2404);
and U2953 (N_2953,N_2111,N_2368);
nor U2954 (N_2954,N_2063,N_2341);
nand U2955 (N_2955,N_2244,N_2380);
or U2956 (N_2956,N_2402,N_2175);
xor U2957 (N_2957,N_2384,N_2368);
nor U2958 (N_2958,N_2343,N_2368);
or U2959 (N_2959,N_2339,N_2195);
or U2960 (N_2960,N_2475,N_2449);
xnor U2961 (N_2961,N_2490,N_2103);
nand U2962 (N_2962,N_2159,N_2151);
or U2963 (N_2963,N_2262,N_2337);
xnor U2964 (N_2964,N_2180,N_2006);
or U2965 (N_2965,N_2042,N_2388);
nand U2966 (N_2966,N_2482,N_2139);
nand U2967 (N_2967,N_2434,N_2335);
xnor U2968 (N_2968,N_2163,N_2205);
nor U2969 (N_2969,N_2064,N_2495);
nor U2970 (N_2970,N_2369,N_2181);
xor U2971 (N_2971,N_2347,N_2305);
nand U2972 (N_2972,N_2110,N_2134);
nor U2973 (N_2973,N_2335,N_2094);
and U2974 (N_2974,N_2452,N_2149);
nand U2975 (N_2975,N_2024,N_2495);
xor U2976 (N_2976,N_2296,N_2143);
and U2977 (N_2977,N_2448,N_2033);
or U2978 (N_2978,N_2178,N_2267);
and U2979 (N_2979,N_2158,N_2321);
and U2980 (N_2980,N_2499,N_2298);
nand U2981 (N_2981,N_2396,N_2275);
and U2982 (N_2982,N_2083,N_2064);
nand U2983 (N_2983,N_2178,N_2062);
xnor U2984 (N_2984,N_2080,N_2417);
nor U2985 (N_2985,N_2191,N_2106);
or U2986 (N_2986,N_2061,N_2446);
nand U2987 (N_2987,N_2187,N_2412);
nand U2988 (N_2988,N_2130,N_2223);
or U2989 (N_2989,N_2279,N_2199);
or U2990 (N_2990,N_2127,N_2148);
or U2991 (N_2991,N_2032,N_2443);
xnor U2992 (N_2992,N_2211,N_2013);
nor U2993 (N_2993,N_2176,N_2470);
or U2994 (N_2994,N_2177,N_2485);
xnor U2995 (N_2995,N_2363,N_2430);
or U2996 (N_2996,N_2455,N_2312);
nor U2997 (N_2997,N_2340,N_2226);
nand U2998 (N_2998,N_2382,N_2161);
and U2999 (N_2999,N_2067,N_2107);
or U3000 (N_3000,N_2552,N_2565);
and U3001 (N_3001,N_2627,N_2912);
xor U3002 (N_3002,N_2982,N_2761);
nand U3003 (N_3003,N_2558,N_2839);
xnor U3004 (N_3004,N_2603,N_2866);
nor U3005 (N_3005,N_2891,N_2846);
nor U3006 (N_3006,N_2831,N_2769);
nand U3007 (N_3007,N_2788,N_2832);
nor U3008 (N_3008,N_2680,N_2529);
nor U3009 (N_3009,N_2981,N_2507);
nand U3010 (N_3010,N_2521,N_2734);
nand U3011 (N_3011,N_2554,N_2805);
nand U3012 (N_3012,N_2931,N_2724);
or U3013 (N_3013,N_2581,N_2870);
nand U3014 (N_3014,N_2617,N_2753);
or U3015 (N_3015,N_2726,N_2875);
nor U3016 (N_3016,N_2571,N_2932);
xor U3017 (N_3017,N_2557,N_2975);
nor U3018 (N_3018,N_2503,N_2682);
or U3019 (N_3019,N_2798,N_2822);
nor U3020 (N_3020,N_2711,N_2659);
xnor U3021 (N_3021,N_2989,N_2671);
and U3022 (N_3022,N_2934,N_2770);
or U3023 (N_3023,N_2904,N_2656);
xnor U3024 (N_3024,N_2625,N_2840);
xnor U3025 (N_3025,N_2909,N_2930);
nor U3026 (N_3026,N_2698,N_2675);
and U3027 (N_3027,N_2823,N_2559);
nand U3028 (N_3028,N_2983,N_2512);
and U3029 (N_3029,N_2588,N_2797);
or U3030 (N_3030,N_2876,N_2593);
nand U3031 (N_3031,N_2774,N_2985);
nor U3032 (N_3032,N_2735,N_2632);
xnor U3033 (N_3033,N_2778,N_2764);
nand U3034 (N_3034,N_2949,N_2992);
nand U3035 (N_3035,N_2629,N_2514);
or U3036 (N_3036,N_2825,N_2852);
or U3037 (N_3037,N_2886,N_2964);
nor U3038 (N_3038,N_2663,N_2515);
nor U3039 (N_3039,N_2619,N_2841);
nor U3040 (N_3040,N_2705,N_2993);
and U3041 (N_3041,N_2898,N_2725);
or U3042 (N_3042,N_2795,N_2543);
and U3043 (N_3043,N_2796,N_2945);
nor U3044 (N_3044,N_2635,N_2608);
or U3045 (N_3045,N_2649,N_2513);
nor U3046 (N_3046,N_2793,N_2707);
nand U3047 (N_3047,N_2908,N_2598);
or U3048 (N_3048,N_2921,N_2884);
or U3049 (N_3049,N_2845,N_2570);
nor U3050 (N_3050,N_2673,N_2703);
xor U3051 (N_3051,N_2509,N_2561);
nor U3052 (N_3052,N_2547,N_2991);
or U3053 (N_3053,N_2887,N_2601);
or U3054 (N_3054,N_2791,N_2551);
xor U3055 (N_3055,N_2502,N_2938);
nand U3056 (N_3056,N_2639,N_2879);
xnor U3057 (N_3057,N_2910,N_2718);
nand U3058 (N_3058,N_2616,N_2668);
and U3059 (N_3059,N_2689,N_2584);
xor U3060 (N_3060,N_2928,N_2759);
and U3061 (N_3061,N_2751,N_2944);
nor U3062 (N_3062,N_2654,N_2517);
nor U3063 (N_3063,N_2924,N_2585);
nand U3064 (N_3064,N_2860,N_2942);
nand U3065 (N_3065,N_2569,N_2713);
or U3066 (N_3066,N_2524,N_2536);
xnor U3067 (N_3067,N_2665,N_2741);
xor U3068 (N_3068,N_2747,N_2806);
or U3069 (N_3069,N_2669,N_2922);
or U3070 (N_3070,N_2530,N_2987);
nor U3071 (N_3071,N_2553,N_2997);
nor U3072 (N_3072,N_2549,N_2775);
nand U3073 (N_3073,N_2780,N_2920);
nor U3074 (N_3074,N_2810,N_2939);
and U3075 (N_3075,N_2790,N_2526);
nand U3076 (N_3076,N_2963,N_2564);
or U3077 (N_3077,N_2956,N_2664);
nand U3078 (N_3078,N_2693,N_2697);
nand U3079 (N_3079,N_2749,N_2511);
and U3080 (N_3080,N_2737,N_2978);
and U3081 (N_3081,N_2634,N_2960);
xor U3082 (N_3082,N_2732,N_2900);
xor U3083 (N_3083,N_2733,N_2504);
xnor U3084 (N_3084,N_2510,N_2731);
xnor U3085 (N_3085,N_2946,N_2618);
nand U3086 (N_3086,N_2636,N_2519);
and U3087 (N_3087,N_2973,N_2817);
xnor U3088 (N_3088,N_2804,N_2915);
xnor U3089 (N_3089,N_2869,N_2853);
and U3090 (N_3090,N_2525,N_2701);
nand U3091 (N_3091,N_2534,N_2962);
xor U3092 (N_3092,N_2905,N_2811);
or U3093 (N_3093,N_2678,N_2913);
xor U3094 (N_3094,N_2628,N_2615);
and U3095 (N_3095,N_2843,N_2833);
or U3096 (N_3096,N_2799,N_2899);
and U3097 (N_3097,N_2646,N_2858);
and U3098 (N_3098,N_2901,N_2609);
nor U3099 (N_3099,N_2683,N_2859);
nor U3100 (N_3100,N_2624,N_2835);
and U3101 (N_3101,N_2729,N_2847);
and U3102 (N_3102,N_2578,N_2856);
nor U3103 (N_3103,N_2610,N_2850);
nor U3104 (N_3104,N_2638,N_2730);
and U3105 (N_3105,N_2955,N_2763);
nand U3106 (N_3106,N_2590,N_2935);
or U3107 (N_3107,N_2816,N_2986);
nand U3108 (N_3108,N_2728,N_2613);
and U3109 (N_3109,N_2976,N_2980);
or U3110 (N_3110,N_2849,N_2742);
xor U3111 (N_3111,N_2819,N_2685);
or U3112 (N_3112,N_2988,N_2784);
or U3113 (N_3113,N_2661,N_2563);
or U3114 (N_3114,N_2885,N_2881);
or U3115 (N_3115,N_2597,N_2918);
or U3116 (N_3116,N_2889,N_2739);
and U3117 (N_3117,N_2560,N_2936);
nor U3118 (N_3118,N_2933,N_2827);
and U3119 (N_3119,N_2854,N_2523);
nand U3120 (N_3120,N_2604,N_2888);
and U3121 (N_3121,N_2974,N_2925);
xnor U3122 (N_3122,N_2591,N_2865);
or U3123 (N_3123,N_2868,N_2872);
or U3124 (N_3124,N_2723,N_2752);
and U3125 (N_3125,N_2531,N_2600);
or U3126 (N_3126,N_2917,N_2815);
or U3127 (N_3127,N_2861,N_2776);
xnor U3128 (N_3128,N_2951,N_2999);
and U3129 (N_3129,N_2589,N_2582);
and U3130 (N_3130,N_2710,N_2684);
or U3131 (N_3131,N_2950,N_2695);
or U3132 (N_3132,N_2568,N_2929);
or U3133 (N_3133,N_2644,N_2677);
or U3134 (N_3134,N_2690,N_2620);
nor U3135 (N_3135,N_2508,N_2660);
nand U3136 (N_3136,N_2757,N_2637);
xnor U3137 (N_3137,N_2541,N_2748);
nor U3138 (N_3138,N_2522,N_2567);
or U3139 (N_3139,N_2878,N_2969);
and U3140 (N_3140,N_2914,N_2652);
xor U3141 (N_3141,N_2653,N_2662);
and U3142 (N_3142,N_2679,N_2961);
or U3143 (N_3143,N_2532,N_2670);
nand U3144 (N_3144,N_2623,N_2607);
and U3145 (N_3145,N_2545,N_2834);
and U3146 (N_3146,N_2970,N_2655);
nor U3147 (N_3147,N_2583,N_2650);
xor U3148 (N_3148,N_2897,N_2765);
nor U3149 (N_3149,N_2596,N_2575);
and U3150 (N_3150,N_2855,N_2786);
or U3151 (N_3151,N_2605,N_2782);
nor U3152 (N_3152,N_2544,N_2681);
or U3153 (N_3153,N_2667,N_2626);
nor U3154 (N_3154,N_2996,N_2916);
or U3155 (N_3155,N_2645,N_2666);
nand U3156 (N_3156,N_2579,N_2779);
nor U3157 (N_3157,N_2621,N_2520);
nor U3158 (N_3158,N_2857,N_2802);
xnor U3159 (N_3159,N_2756,N_2768);
xor U3160 (N_3160,N_2577,N_2702);
or U3161 (N_3161,N_2893,N_2586);
nand U3162 (N_3162,N_2794,N_2592);
nor U3163 (N_3163,N_2995,N_2801);
or U3164 (N_3164,N_2630,N_2821);
xor U3165 (N_3165,N_2754,N_2542);
nand U3166 (N_3166,N_2674,N_2830);
and U3167 (N_3167,N_2880,N_2844);
nor U3168 (N_3168,N_2550,N_2708);
xor U3169 (N_3169,N_2574,N_2506);
or U3170 (N_3170,N_2959,N_2750);
nor U3171 (N_3171,N_2952,N_2744);
nand U3172 (N_3172,N_2958,N_2984);
nor U3173 (N_3173,N_2657,N_2937);
nor U3174 (N_3174,N_2712,N_2813);
nand U3175 (N_3175,N_2940,N_2760);
nor U3176 (N_3176,N_2562,N_2838);
nor U3177 (N_3177,N_2533,N_2687);
xnor U3178 (N_3178,N_2692,N_2848);
nand U3179 (N_3179,N_2783,N_2717);
or U3180 (N_3180,N_2647,N_2941);
xnor U3181 (N_3181,N_2537,N_2501);
xnor U3182 (N_3182,N_2863,N_2643);
nor U3183 (N_3183,N_2998,N_2926);
nor U3184 (N_3184,N_2923,N_2709);
or U3185 (N_3185,N_2965,N_2871);
nor U3186 (N_3186,N_2640,N_2594);
xor U3187 (N_3187,N_2696,N_2967);
and U3188 (N_3188,N_2648,N_2612);
nor U3189 (N_3189,N_2927,N_2867);
nand U3190 (N_3190,N_2611,N_2546);
nor U3191 (N_3191,N_2785,N_2676);
nand U3192 (N_3192,N_2743,N_2721);
and U3193 (N_3193,N_2505,N_2540);
or U3194 (N_3194,N_2812,N_2957);
and U3195 (N_3195,N_2826,N_2953);
xnor U3196 (N_3196,N_2755,N_2716);
and U3197 (N_3197,N_2527,N_2758);
and U3198 (N_3198,N_2633,N_2727);
nand U3199 (N_3199,N_2837,N_2792);
xor U3200 (N_3200,N_2902,N_2736);
and U3201 (N_3201,N_2738,N_2836);
nor U3202 (N_3202,N_2943,N_2911);
nand U3203 (N_3203,N_2704,N_2548);
and U3204 (N_3204,N_2714,N_2641);
and U3205 (N_3205,N_2528,N_2971);
or U3206 (N_3206,N_2882,N_2691);
and U3207 (N_3207,N_2566,N_2556);
nor U3208 (N_3208,N_2800,N_2948);
and U3209 (N_3209,N_2658,N_2972);
nor U3210 (N_3210,N_2614,N_2602);
nand U3211 (N_3211,N_2947,N_2883);
nand U3212 (N_3212,N_2890,N_2580);
xnor U3213 (N_3213,N_2873,N_2535);
nor U3214 (N_3214,N_2771,N_2672);
xnor U3215 (N_3215,N_2824,N_2722);
nand U3216 (N_3216,N_2954,N_2777);
nor U3217 (N_3217,N_2894,N_2700);
xnor U3218 (N_3218,N_2500,N_2818);
xnor U3219 (N_3219,N_2706,N_2968);
and U3220 (N_3220,N_2595,N_2694);
or U3221 (N_3221,N_2572,N_2599);
nand U3222 (N_3222,N_2979,N_2809);
and U3223 (N_3223,N_2587,N_2686);
xnor U3224 (N_3224,N_2745,N_2919);
or U3225 (N_3225,N_2842,N_2896);
nand U3226 (N_3226,N_2977,N_2906);
and U3227 (N_3227,N_2720,N_2767);
and U3228 (N_3228,N_2808,N_2781);
and U3229 (N_3229,N_2994,N_2576);
nor U3230 (N_3230,N_2789,N_2766);
nand U3231 (N_3231,N_2688,N_2719);
nand U3232 (N_3232,N_2555,N_2803);
and U3233 (N_3233,N_2762,N_2990);
nor U3234 (N_3234,N_2622,N_2787);
nor U3235 (N_3235,N_2606,N_2877);
or U3236 (N_3236,N_2746,N_2966);
nor U3237 (N_3237,N_2773,N_2772);
and U3238 (N_3238,N_2740,N_2642);
and U3239 (N_3239,N_2631,N_2715);
xor U3240 (N_3240,N_2828,N_2895);
and U3241 (N_3241,N_2864,N_2807);
xor U3242 (N_3242,N_2814,N_2699);
and U3243 (N_3243,N_2573,N_2538);
nor U3244 (N_3244,N_2651,N_2862);
and U3245 (N_3245,N_2539,N_2907);
nand U3246 (N_3246,N_2820,N_2851);
xor U3247 (N_3247,N_2892,N_2829);
and U3248 (N_3248,N_2874,N_2518);
xnor U3249 (N_3249,N_2903,N_2516);
or U3250 (N_3250,N_2929,N_2977);
or U3251 (N_3251,N_2733,N_2829);
or U3252 (N_3252,N_2712,N_2697);
or U3253 (N_3253,N_2984,N_2888);
nand U3254 (N_3254,N_2639,N_2758);
and U3255 (N_3255,N_2670,N_2969);
and U3256 (N_3256,N_2629,N_2764);
nor U3257 (N_3257,N_2822,N_2953);
and U3258 (N_3258,N_2602,N_2848);
nor U3259 (N_3259,N_2851,N_2679);
nand U3260 (N_3260,N_2707,N_2536);
nor U3261 (N_3261,N_2578,N_2950);
nor U3262 (N_3262,N_2994,N_2744);
or U3263 (N_3263,N_2965,N_2731);
nor U3264 (N_3264,N_2711,N_2710);
and U3265 (N_3265,N_2730,N_2994);
xnor U3266 (N_3266,N_2901,N_2770);
xor U3267 (N_3267,N_2755,N_2839);
nor U3268 (N_3268,N_2505,N_2783);
xor U3269 (N_3269,N_2954,N_2966);
and U3270 (N_3270,N_2727,N_2524);
xnor U3271 (N_3271,N_2933,N_2669);
or U3272 (N_3272,N_2889,N_2641);
nor U3273 (N_3273,N_2995,N_2563);
nor U3274 (N_3274,N_2820,N_2840);
xor U3275 (N_3275,N_2680,N_2546);
nand U3276 (N_3276,N_2903,N_2931);
or U3277 (N_3277,N_2522,N_2717);
and U3278 (N_3278,N_2642,N_2717);
xnor U3279 (N_3279,N_2928,N_2556);
or U3280 (N_3280,N_2785,N_2729);
or U3281 (N_3281,N_2522,N_2679);
nor U3282 (N_3282,N_2604,N_2856);
nand U3283 (N_3283,N_2780,N_2584);
xor U3284 (N_3284,N_2642,N_2731);
nor U3285 (N_3285,N_2554,N_2772);
xnor U3286 (N_3286,N_2536,N_2874);
and U3287 (N_3287,N_2869,N_2756);
or U3288 (N_3288,N_2956,N_2866);
nand U3289 (N_3289,N_2877,N_2966);
or U3290 (N_3290,N_2709,N_2662);
nor U3291 (N_3291,N_2868,N_2867);
or U3292 (N_3292,N_2700,N_2994);
and U3293 (N_3293,N_2987,N_2515);
nand U3294 (N_3294,N_2676,N_2842);
or U3295 (N_3295,N_2728,N_2881);
nand U3296 (N_3296,N_2890,N_2884);
nor U3297 (N_3297,N_2667,N_2589);
xnor U3298 (N_3298,N_2842,N_2915);
and U3299 (N_3299,N_2725,N_2792);
nand U3300 (N_3300,N_2527,N_2645);
or U3301 (N_3301,N_2929,N_2751);
xnor U3302 (N_3302,N_2808,N_2769);
xor U3303 (N_3303,N_2991,N_2735);
or U3304 (N_3304,N_2962,N_2723);
nand U3305 (N_3305,N_2876,N_2788);
or U3306 (N_3306,N_2862,N_2989);
xor U3307 (N_3307,N_2894,N_2996);
nor U3308 (N_3308,N_2536,N_2617);
nand U3309 (N_3309,N_2567,N_2840);
and U3310 (N_3310,N_2920,N_2519);
or U3311 (N_3311,N_2527,N_2842);
nand U3312 (N_3312,N_2534,N_2825);
nand U3313 (N_3313,N_2860,N_2804);
nor U3314 (N_3314,N_2620,N_2681);
and U3315 (N_3315,N_2575,N_2781);
or U3316 (N_3316,N_2908,N_2696);
nor U3317 (N_3317,N_2671,N_2813);
and U3318 (N_3318,N_2745,N_2620);
and U3319 (N_3319,N_2746,N_2656);
nand U3320 (N_3320,N_2929,N_2746);
or U3321 (N_3321,N_2591,N_2661);
nor U3322 (N_3322,N_2582,N_2940);
nor U3323 (N_3323,N_2909,N_2775);
and U3324 (N_3324,N_2724,N_2599);
nor U3325 (N_3325,N_2783,N_2830);
nor U3326 (N_3326,N_2583,N_2565);
and U3327 (N_3327,N_2690,N_2604);
xnor U3328 (N_3328,N_2752,N_2671);
xnor U3329 (N_3329,N_2748,N_2515);
or U3330 (N_3330,N_2901,N_2920);
xor U3331 (N_3331,N_2986,N_2778);
nand U3332 (N_3332,N_2969,N_2675);
and U3333 (N_3333,N_2685,N_2593);
xor U3334 (N_3334,N_2874,N_2509);
nor U3335 (N_3335,N_2808,N_2723);
xnor U3336 (N_3336,N_2909,N_2536);
nand U3337 (N_3337,N_2986,N_2607);
nor U3338 (N_3338,N_2649,N_2693);
and U3339 (N_3339,N_2708,N_2979);
or U3340 (N_3340,N_2971,N_2871);
and U3341 (N_3341,N_2718,N_2825);
or U3342 (N_3342,N_2606,N_2953);
and U3343 (N_3343,N_2626,N_2508);
and U3344 (N_3344,N_2562,N_2964);
and U3345 (N_3345,N_2716,N_2641);
or U3346 (N_3346,N_2815,N_2942);
and U3347 (N_3347,N_2688,N_2558);
or U3348 (N_3348,N_2533,N_2880);
or U3349 (N_3349,N_2589,N_2556);
xnor U3350 (N_3350,N_2682,N_2727);
nor U3351 (N_3351,N_2691,N_2873);
nor U3352 (N_3352,N_2700,N_2726);
nor U3353 (N_3353,N_2958,N_2688);
nor U3354 (N_3354,N_2801,N_2724);
nand U3355 (N_3355,N_2984,N_2764);
or U3356 (N_3356,N_2786,N_2640);
or U3357 (N_3357,N_2898,N_2890);
or U3358 (N_3358,N_2975,N_2540);
and U3359 (N_3359,N_2553,N_2659);
nand U3360 (N_3360,N_2988,N_2697);
or U3361 (N_3361,N_2846,N_2511);
xor U3362 (N_3362,N_2632,N_2796);
and U3363 (N_3363,N_2944,N_2578);
and U3364 (N_3364,N_2999,N_2642);
and U3365 (N_3365,N_2789,N_2937);
nand U3366 (N_3366,N_2932,N_2634);
nor U3367 (N_3367,N_2799,N_2653);
nand U3368 (N_3368,N_2661,N_2911);
nor U3369 (N_3369,N_2948,N_2792);
nor U3370 (N_3370,N_2993,N_2640);
xor U3371 (N_3371,N_2650,N_2579);
or U3372 (N_3372,N_2927,N_2793);
nor U3373 (N_3373,N_2821,N_2883);
nor U3374 (N_3374,N_2619,N_2802);
or U3375 (N_3375,N_2601,N_2714);
nand U3376 (N_3376,N_2533,N_2580);
xnor U3377 (N_3377,N_2886,N_2579);
or U3378 (N_3378,N_2918,N_2851);
and U3379 (N_3379,N_2907,N_2632);
nand U3380 (N_3380,N_2798,N_2882);
nand U3381 (N_3381,N_2566,N_2847);
xor U3382 (N_3382,N_2914,N_2593);
or U3383 (N_3383,N_2568,N_2803);
nand U3384 (N_3384,N_2848,N_2690);
and U3385 (N_3385,N_2777,N_2696);
xnor U3386 (N_3386,N_2704,N_2715);
or U3387 (N_3387,N_2857,N_2524);
or U3388 (N_3388,N_2641,N_2554);
xnor U3389 (N_3389,N_2871,N_2862);
nor U3390 (N_3390,N_2683,N_2679);
and U3391 (N_3391,N_2890,N_2685);
nor U3392 (N_3392,N_2646,N_2621);
nor U3393 (N_3393,N_2667,N_2755);
nand U3394 (N_3394,N_2679,N_2787);
and U3395 (N_3395,N_2892,N_2817);
or U3396 (N_3396,N_2999,N_2716);
nand U3397 (N_3397,N_2966,N_2691);
nor U3398 (N_3398,N_2999,N_2558);
xor U3399 (N_3399,N_2968,N_2851);
nor U3400 (N_3400,N_2945,N_2628);
nor U3401 (N_3401,N_2712,N_2819);
xnor U3402 (N_3402,N_2977,N_2841);
nand U3403 (N_3403,N_2893,N_2722);
or U3404 (N_3404,N_2608,N_2792);
nor U3405 (N_3405,N_2907,N_2874);
nor U3406 (N_3406,N_2851,N_2771);
and U3407 (N_3407,N_2650,N_2611);
nor U3408 (N_3408,N_2744,N_2793);
xnor U3409 (N_3409,N_2578,N_2924);
or U3410 (N_3410,N_2934,N_2929);
nor U3411 (N_3411,N_2970,N_2832);
xor U3412 (N_3412,N_2836,N_2653);
and U3413 (N_3413,N_2642,N_2562);
and U3414 (N_3414,N_2904,N_2852);
and U3415 (N_3415,N_2836,N_2857);
xnor U3416 (N_3416,N_2683,N_2792);
nand U3417 (N_3417,N_2633,N_2778);
xnor U3418 (N_3418,N_2573,N_2755);
nor U3419 (N_3419,N_2719,N_2810);
xnor U3420 (N_3420,N_2607,N_2879);
nor U3421 (N_3421,N_2551,N_2680);
nor U3422 (N_3422,N_2909,N_2512);
nor U3423 (N_3423,N_2983,N_2563);
xor U3424 (N_3424,N_2871,N_2516);
xor U3425 (N_3425,N_2974,N_2940);
nor U3426 (N_3426,N_2523,N_2605);
nand U3427 (N_3427,N_2768,N_2915);
or U3428 (N_3428,N_2870,N_2631);
and U3429 (N_3429,N_2524,N_2911);
nor U3430 (N_3430,N_2985,N_2520);
nor U3431 (N_3431,N_2510,N_2911);
or U3432 (N_3432,N_2801,N_2657);
and U3433 (N_3433,N_2851,N_2852);
or U3434 (N_3434,N_2815,N_2622);
nor U3435 (N_3435,N_2775,N_2816);
nand U3436 (N_3436,N_2972,N_2866);
nor U3437 (N_3437,N_2672,N_2675);
xnor U3438 (N_3438,N_2786,N_2646);
xor U3439 (N_3439,N_2928,N_2515);
nand U3440 (N_3440,N_2757,N_2725);
nand U3441 (N_3441,N_2846,N_2719);
nor U3442 (N_3442,N_2870,N_2780);
nor U3443 (N_3443,N_2619,N_2891);
and U3444 (N_3444,N_2932,N_2880);
nor U3445 (N_3445,N_2665,N_2623);
nand U3446 (N_3446,N_2956,N_2847);
xor U3447 (N_3447,N_2774,N_2673);
xnor U3448 (N_3448,N_2574,N_2541);
nand U3449 (N_3449,N_2548,N_2902);
and U3450 (N_3450,N_2610,N_2836);
and U3451 (N_3451,N_2722,N_2515);
nor U3452 (N_3452,N_2837,N_2629);
or U3453 (N_3453,N_2506,N_2748);
nor U3454 (N_3454,N_2821,N_2571);
nand U3455 (N_3455,N_2577,N_2933);
nand U3456 (N_3456,N_2876,N_2501);
or U3457 (N_3457,N_2987,N_2773);
nand U3458 (N_3458,N_2840,N_2915);
and U3459 (N_3459,N_2533,N_2903);
or U3460 (N_3460,N_2793,N_2752);
nand U3461 (N_3461,N_2888,N_2511);
and U3462 (N_3462,N_2621,N_2917);
nor U3463 (N_3463,N_2683,N_2530);
and U3464 (N_3464,N_2540,N_2745);
nor U3465 (N_3465,N_2851,N_2788);
or U3466 (N_3466,N_2958,N_2710);
nand U3467 (N_3467,N_2762,N_2880);
or U3468 (N_3468,N_2755,N_2916);
and U3469 (N_3469,N_2799,N_2771);
xnor U3470 (N_3470,N_2557,N_2708);
xor U3471 (N_3471,N_2977,N_2541);
xor U3472 (N_3472,N_2913,N_2599);
nand U3473 (N_3473,N_2919,N_2952);
or U3474 (N_3474,N_2834,N_2533);
nand U3475 (N_3475,N_2844,N_2513);
and U3476 (N_3476,N_2957,N_2659);
and U3477 (N_3477,N_2900,N_2787);
nor U3478 (N_3478,N_2708,N_2792);
nand U3479 (N_3479,N_2855,N_2897);
or U3480 (N_3480,N_2569,N_2502);
or U3481 (N_3481,N_2559,N_2987);
nor U3482 (N_3482,N_2923,N_2753);
nand U3483 (N_3483,N_2604,N_2723);
and U3484 (N_3484,N_2958,N_2693);
nor U3485 (N_3485,N_2571,N_2804);
and U3486 (N_3486,N_2918,N_2669);
nand U3487 (N_3487,N_2698,N_2619);
nor U3488 (N_3488,N_2665,N_2941);
nand U3489 (N_3489,N_2838,N_2790);
nor U3490 (N_3490,N_2580,N_2601);
or U3491 (N_3491,N_2713,N_2642);
or U3492 (N_3492,N_2512,N_2896);
or U3493 (N_3493,N_2917,N_2969);
or U3494 (N_3494,N_2842,N_2727);
xor U3495 (N_3495,N_2831,N_2656);
nor U3496 (N_3496,N_2816,N_2625);
and U3497 (N_3497,N_2816,N_2771);
and U3498 (N_3498,N_2976,N_2760);
xor U3499 (N_3499,N_2788,N_2737);
or U3500 (N_3500,N_3419,N_3464);
nor U3501 (N_3501,N_3346,N_3083);
or U3502 (N_3502,N_3459,N_3022);
and U3503 (N_3503,N_3390,N_3029);
and U3504 (N_3504,N_3077,N_3063);
xnor U3505 (N_3505,N_3446,N_3236);
xor U3506 (N_3506,N_3131,N_3408);
nand U3507 (N_3507,N_3074,N_3386);
xnor U3508 (N_3508,N_3358,N_3240);
nor U3509 (N_3509,N_3338,N_3052);
or U3510 (N_3510,N_3411,N_3364);
xor U3511 (N_3511,N_3001,N_3102);
and U3512 (N_3512,N_3277,N_3324);
nand U3513 (N_3513,N_3002,N_3312);
or U3514 (N_3514,N_3397,N_3153);
xor U3515 (N_3515,N_3202,N_3165);
nor U3516 (N_3516,N_3299,N_3495);
and U3517 (N_3517,N_3264,N_3439);
nand U3518 (N_3518,N_3460,N_3339);
and U3519 (N_3519,N_3210,N_3492);
nor U3520 (N_3520,N_3127,N_3059);
or U3521 (N_3521,N_3219,N_3391);
or U3522 (N_3522,N_3200,N_3152);
and U3523 (N_3523,N_3173,N_3204);
or U3524 (N_3524,N_3344,N_3413);
xor U3525 (N_3525,N_3349,N_3020);
nor U3526 (N_3526,N_3087,N_3129);
nand U3527 (N_3527,N_3280,N_3222);
xor U3528 (N_3528,N_3073,N_3212);
nor U3529 (N_3529,N_3137,N_3490);
xor U3530 (N_3530,N_3148,N_3021);
nand U3531 (N_3531,N_3337,N_3448);
nor U3532 (N_3532,N_3079,N_3463);
nor U3533 (N_3533,N_3076,N_3314);
xnor U3534 (N_3534,N_3479,N_3383);
xnor U3535 (N_3535,N_3011,N_3159);
and U3536 (N_3536,N_3010,N_3190);
nor U3537 (N_3537,N_3350,N_3288);
nor U3538 (N_3538,N_3496,N_3354);
and U3539 (N_3539,N_3427,N_3160);
and U3540 (N_3540,N_3032,N_3154);
and U3541 (N_3541,N_3453,N_3370);
or U3542 (N_3542,N_3319,N_3326);
nor U3543 (N_3543,N_3357,N_3382);
or U3544 (N_3544,N_3385,N_3488);
or U3545 (N_3545,N_3053,N_3051);
and U3546 (N_3546,N_3150,N_3341);
and U3547 (N_3547,N_3351,N_3374);
xnor U3548 (N_3548,N_3449,N_3207);
nand U3549 (N_3549,N_3033,N_3213);
nor U3550 (N_3550,N_3230,N_3362);
nand U3551 (N_3551,N_3157,N_3273);
xnor U3552 (N_3552,N_3293,N_3115);
xor U3553 (N_3553,N_3205,N_3146);
xnor U3554 (N_3554,N_3166,N_3430);
xnor U3555 (N_3555,N_3256,N_3260);
and U3556 (N_3556,N_3468,N_3109);
xnor U3557 (N_3557,N_3359,N_3356);
or U3558 (N_3558,N_3306,N_3461);
xnor U3559 (N_3559,N_3130,N_3257);
xor U3560 (N_3560,N_3151,N_3423);
or U3561 (N_3561,N_3380,N_3315);
nand U3562 (N_3562,N_3226,N_3353);
and U3563 (N_3563,N_3434,N_3469);
nor U3564 (N_3564,N_3118,N_3367);
and U3565 (N_3565,N_3497,N_3333);
nand U3566 (N_3566,N_3307,N_3134);
or U3567 (N_3567,N_3193,N_3223);
and U3568 (N_3568,N_3061,N_3431);
and U3569 (N_3569,N_3041,N_3366);
or U3570 (N_3570,N_3106,N_3238);
and U3571 (N_3571,N_3388,N_3111);
nor U3572 (N_3572,N_3368,N_3247);
and U3573 (N_3573,N_3283,N_3140);
or U3574 (N_3574,N_3278,N_3178);
and U3575 (N_3575,N_3142,N_3425);
or U3576 (N_3576,N_3286,N_3440);
or U3577 (N_3577,N_3327,N_3062);
xnor U3578 (N_3578,N_3476,N_3398);
and U3579 (N_3579,N_3184,N_3169);
xnor U3580 (N_3580,N_3114,N_3034);
or U3581 (N_3581,N_3329,N_3447);
xnor U3582 (N_3582,N_3285,N_3217);
xnor U3583 (N_3583,N_3484,N_3234);
xor U3584 (N_3584,N_3451,N_3465);
or U3585 (N_3585,N_3231,N_3404);
nor U3586 (N_3586,N_3069,N_3158);
xor U3587 (N_3587,N_3136,N_3008);
xnor U3588 (N_3588,N_3026,N_3214);
nor U3589 (N_3589,N_3443,N_3117);
and U3590 (N_3590,N_3271,N_3313);
or U3591 (N_3591,N_3302,N_3135);
or U3592 (N_3592,N_3420,N_3120);
nor U3593 (N_3593,N_3099,N_3013);
and U3594 (N_3594,N_3429,N_3263);
or U3595 (N_3595,N_3177,N_3309);
or U3596 (N_3596,N_3037,N_3252);
nand U3597 (N_3597,N_3057,N_3025);
nor U3598 (N_3598,N_3220,N_3477);
and U3599 (N_3599,N_3227,N_3458);
and U3600 (N_3600,N_3405,N_3147);
or U3601 (N_3601,N_3498,N_3108);
xnor U3602 (N_3602,N_3412,N_3239);
or U3603 (N_3603,N_3081,N_3416);
or U3604 (N_3604,N_3325,N_3332);
and U3605 (N_3605,N_3144,N_3308);
xor U3606 (N_3606,N_3028,N_3279);
nor U3607 (N_3607,N_3094,N_3375);
nand U3608 (N_3608,N_3365,N_3065);
xnor U3609 (N_3609,N_3191,N_3133);
nand U3610 (N_3610,N_3066,N_3348);
xnor U3611 (N_3611,N_3345,N_3276);
or U3612 (N_3612,N_3267,N_3244);
and U3613 (N_3613,N_3067,N_3036);
and U3614 (N_3614,N_3304,N_3005);
nand U3615 (N_3615,N_3107,N_3183);
nand U3616 (N_3616,N_3038,N_3249);
nor U3617 (N_3617,N_3141,N_3409);
xor U3618 (N_3618,N_3282,N_3289);
nor U3619 (N_3619,N_3387,N_3172);
nand U3620 (N_3620,N_3377,N_3229);
nor U3621 (N_3621,N_3410,N_3424);
and U3622 (N_3622,N_3342,N_3018);
nor U3623 (N_3623,N_3167,N_3196);
nor U3624 (N_3624,N_3188,N_3078);
xor U3625 (N_3625,N_3072,N_3093);
xor U3626 (N_3626,N_3044,N_3487);
or U3627 (N_3627,N_3369,N_3334);
xnor U3628 (N_3628,N_3261,N_3444);
nor U3629 (N_3629,N_3352,N_3281);
or U3630 (N_3630,N_3189,N_3291);
xor U3631 (N_3631,N_3015,N_3457);
nor U3632 (N_3632,N_3237,N_3486);
nor U3633 (N_3633,N_3262,N_3201);
nor U3634 (N_3634,N_3401,N_3268);
and U3635 (N_3635,N_3456,N_3426);
nand U3636 (N_3636,N_3270,N_3128);
or U3637 (N_3637,N_3432,N_3499);
xor U3638 (N_3638,N_3428,N_3030);
and U3639 (N_3639,N_3480,N_3121);
and U3640 (N_3640,N_3211,N_3295);
xnor U3641 (N_3641,N_3320,N_3472);
nor U3642 (N_3642,N_3489,N_3376);
or U3643 (N_3643,N_3441,N_3049);
nand U3644 (N_3644,N_3355,N_3467);
or U3645 (N_3645,N_3481,N_3347);
xnor U3646 (N_3646,N_3216,N_3475);
and U3647 (N_3647,N_3290,N_3360);
nand U3648 (N_3648,N_3292,N_3126);
nand U3649 (N_3649,N_3174,N_3123);
or U3650 (N_3650,N_3048,N_3180);
xnor U3651 (N_3651,N_3040,N_3361);
nand U3652 (N_3652,N_3050,N_3009);
nand U3653 (N_3653,N_3155,N_3395);
nand U3654 (N_3654,N_3466,N_3023);
nand U3655 (N_3655,N_3266,N_3328);
nand U3656 (N_3656,N_3491,N_3101);
and U3657 (N_3657,N_3161,N_3179);
and U3658 (N_3658,N_3149,N_3493);
or U3659 (N_3659,N_3483,N_3272);
or U3660 (N_3660,N_3006,N_3335);
or U3661 (N_3661,N_3317,N_3163);
nor U3662 (N_3662,N_3417,N_3071);
nor U3663 (N_3663,N_3372,N_3233);
and U3664 (N_3664,N_3402,N_3445);
nand U3665 (N_3665,N_3186,N_3340);
or U3666 (N_3666,N_3403,N_3259);
and U3667 (N_3667,N_3242,N_3470);
nand U3668 (N_3668,N_3406,N_3321);
nand U3669 (N_3669,N_3045,N_3436);
xor U3670 (N_3670,N_3132,N_3474);
or U3671 (N_3671,N_3092,N_3396);
nor U3672 (N_3672,N_3206,N_3039);
nand U3673 (N_3673,N_3343,N_3287);
nand U3674 (N_3674,N_3225,N_3415);
nand U3675 (N_3675,N_3203,N_3000);
and U3676 (N_3676,N_3450,N_3215);
xor U3677 (N_3677,N_3125,N_3455);
or U3678 (N_3678,N_3218,N_3494);
nand U3679 (N_3679,N_3182,N_3209);
or U3680 (N_3680,N_3012,N_3122);
or U3681 (N_3681,N_3085,N_3265);
nor U3682 (N_3682,N_3473,N_3228);
nand U3683 (N_3683,N_3454,N_3197);
or U3684 (N_3684,N_3103,N_3086);
or U3685 (N_3685,N_3322,N_3331);
xor U3686 (N_3686,N_3414,N_3298);
xor U3687 (N_3687,N_3068,N_3407);
nor U3688 (N_3688,N_3003,N_3082);
nand U3689 (N_3689,N_3399,N_3323);
xor U3690 (N_3690,N_3296,N_3185);
xnor U3691 (N_3691,N_3090,N_3379);
or U3692 (N_3692,N_3007,N_3031);
xor U3693 (N_3693,N_3253,N_3139);
nand U3694 (N_3694,N_3100,N_3042);
or U3695 (N_3695,N_3330,N_3088);
xor U3696 (N_3696,N_3187,N_3195);
nand U3697 (N_3697,N_3274,N_3112);
or U3698 (N_3698,N_3363,N_3097);
xnor U3699 (N_3699,N_3438,N_3176);
or U3700 (N_3700,N_3208,N_3046);
xnor U3701 (N_3701,N_3194,N_3171);
nor U3702 (N_3702,N_3232,N_3269);
and U3703 (N_3703,N_3113,N_3170);
and U3704 (N_3704,N_3110,N_3175);
xor U3705 (N_3705,N_3145,N_3224);
nor U3706 (N_3706,N_3014,N_3243);
nand U3707 (N_3707,N_3381,N_3373);
or U3708 (N_3708,N_3442,N_3254);
and U3709 (N_3709,N_3394,N_3084);
nand U3710 (N_3710,N_3258,N_3168);
or U3711 (N_3711,N_3162,N_3422);
nor U3712 (N_3712,N_3482,N_3452);
nor U3713 (N_3713,N_3004,N_3384);
and U3714 (N_3714,N_3433,N_3080);
and U3715 (N_3715,N_3310,N_3156);
xor U3716 (N_3716,N_3393,N_3116);
nor U3717 (N_3717,N_3305,N_3070);
and U3718 (N_3718,N_3301,N_3318);
xor U3719 (N_3719,N_3297,N_3019);
nor U3720 (N_3720,N_3462,N_3392);
or U3721 (N_3721,N_3058,N_3248);
and U3722 (N_3722,N_3199,N_3075);
nor U3723 (N_3723,N_3047,N_3437);
or U3724 (N_3724,N_3035,N_3192);
and U3725 (N_3725,N_3246,N_3303);
or U3726 (N_3726,N_3284,N_3138);
and U3727 (N_3727,N_3471,N_3378);
nor U3728 (N_3728,N_3435,N_3235);
or U3729 (N_3729,N_3024,N_3245);
or U3730 (N_3730,N_3198,N_3275);
nor U3731 (N_3731,N_3095,N_3478);
and U3732 (N_3732,N_3060,N_3089);
and U3733 (N_3733,N_3124,N_3294);
or U3734 (N_3734,N_3389,N_3221);
and U3735 (N_3735,N_3421,N_3311);
and U3736 (N_3736,N_3250,N_3300);
or U3737 (N_3737,N_3336,N_3017);
xnor U3738 (N_3738,N_3043,N_3485);
nand U3739 (N_3739,N_3143,N_3371);
nand U3740 (N_3740,N_3251,N_3418);
nand U3741 (N_3741,N_3255,N_3164);
and U3742 (N_3742,N_3055,N_3105);
nor U3743 (N_3743,N_3119,N_3056);
nand U3744 (N_3744,N_3400,N_3241);
xor U3745 (N_3745,N_3064,N_3098);
nor U3746 (N_3746,N_3096,N_3091);
and U3747 (N_3747,N_3054,N_3181);
and U3748 (N_3748,N_3104,N_3316);
and U3749 (N_3749,N_3016,N_3027);
nor U3750 (N_3750,N_3240,N_3146);
or U3751 (N_3751,N_3484,N_3250);
or U3752 (N_3752,N_3433,N_3364);
xnor U3753 (N_3753,N_3303,N_3420);
or U3754 (N_3754,N_3288,N_3127);
nor U3755 (N_3755,N_3449,N_3293);
nand U3756 (N_3756,N_3378,N_3288);
and U3757 (N_3757,N_3303,N_3142);
or U3758 (N_3758,N_3243,N_3125);
xor U3759 (N_3759,N_3179,N_3455);
xnor U3760 (N_3760,N_3407,N_3051);
nand U3761 (N_3761,N_3123,N_3248);
and U3762 (N_3762,N_3037,N_3154);
and U3763 (N_3763,N_3474,N_3349);
and U3764 (N_3764,N_3347,N_3393);
or U3765 (N_3765,N_3471,N_3400);
xor U3766 (N_3766,N_3015,N_3045);
and U3767 (N_3767,N_3071,N_3241);
and U3768 (N_3768,N_3180,N_3271);
and U3769 (N_3769,N_3000,N_3139);
nand U3770 (N_3770,N_3235,N_3451);
or U3771 (N_3771,N_3467,N_3052);
nor U3772 (N_3772,N_3248,N_3060);
nor U3773 (N_3773,N_3261,N_3388);
nand U3774 (N_3774,N_3033,N_3160);
or U3775 (N_3775,N_3384,N_3247);
nand U3776 (N_3776,N_3127,N_3066);
xor U3777 (N_3777,N_3065,N_3418);
xnor U3778 (N_3778,N_3195,N_3227);
and U3779 (N_3779,N_3416,N_3000);
nand U3780 (N_3780,N_3461,N_3010);
and U3781 (N_3781,N_3007,N_3418);
or U3782 (N_3782,N_3193,N_3374);
nor U3783 (N_3783,N_3409,N_3219);
and U3784 (N_3784,N_3178,N_3390);
nand U3785 (N_3785,N_3098,N_3232);
nor U3786 (N_3786,N_3219,N_3462);
nand U3787 (N_3787,N_3492,N_3457);
or U3788 (N_3788,N_3366,N_3069);
nand U3789 (N_3789,N_3155,N_3020);
nand U3790 (N_3790,N_3167,N_3464);
nand U3791 (N_3791,N_3174,N_3284);
or U3792 (N_3792,N_3213,N_3266);
xor U3793 (N_3793,N_3403,N_3124);
or U3794 (N_3794,N_3173,N_3008);
nand U3795 (N_3795,N_3386,N_3469);
and U3796 (N_3796,N_3100,N_3398);
or U3797 (N_3797,N_3232,N_3195);
nand U3798 (N_3798,N_3013,N_3372);
and U3799 (N_3799,N_3232,N_3497);
nor U3800 (N_3800,N_3406,N_3122);
nand U3801 (N_3801,N_3348,N_3154);
xnor U3802 (N_3802,N_3225,N_3272);
nor U3803 (N_3803,N_3293,N_3048);
or U3804 (N_3804,N_3466,N_3360);
nor U3805 (N_3805,N_3127,N_3403);
nor U3806 (N_3806,N_3445,N_3497);
and U3807 (N_3807,N_3324,N_3310);
or U3808 (N_3808,N_3336,N_3248);
xor U3809 (N_3809,N_3109,N_3201);
xnor U3810 (N_3810,N_3223,N_3493);
xor U3811 (N_3811,N_3052,N_3013);
nor U3812 (N_3812,N_3487,N_3050);
xnor U3813 (N_3813,N_3496,N_3165);
xor U3814 (N_3814,N_3236,N_3173);
nor U3815 (N_3815,N_3339,N_3396);
xnor U3816 (N_3816,N_3220,N_3469);
nor U3817 (N_3817,N_3059,N_3324);
nor U3818 (N_3818,N_3342,N_3238);
nor U3819 (N_3819,N_3140,N_3088);
xor U3820 (N_3820,N_3226,N_3330);
or U3821 (N_3821,N_3300,N_3273);
or U3822 (N_3822,N_3188,N_3169);
xor U3823 (N_3823,N_3042,N_3064);
nand U3824 (N_3824,N_3199,N_3231);
nor U3825 (N_3825,N_3357,N_3373);
and U3826 (N_3826,N_3281,N_3061);
nand U3827 (N_3827,N_3358,N_3131);
or U3828 (N_3828,N_3386,N_3104);
nor U3829 (N_3829,N_3247,N_3275);
nand U3830 (N_3830,N_3023,N_3060);
nor U3831 (N_3831,N_3209,N_3294);
xnor U3832 (N_3832,N_3049,N_3487);
and U3833 (N_3833,N_3096,N_3286);
nand U3834 (N_3834,N_3073,N_3088);
and U3835 (N_3835,N_3052,N_3039);
xor U3836 (N_3836,N_3466,N_3470);
and U3837 (N_3837,N_3318,N_3349);
nor U3838 (N_3838,N_3443,N_3063);
nand U3839 (N_3839,N_3460,N_3480);
nor U3840 (N_3840,N_3049,N_3212);
and U3841 (N_3841,N_3260,N_3031);
or U3842 (N_3842,N_3064,N_3253);
and U3843 (N_3843,N_3071,N_3253);
nor U3844 (N_3844,N_3237,N_3134);
and U3845 (N_3845,N_3324,N_3015);
or U3846 (N_3846,N_3072,N_3193);
xnor U3847 (N_3847,N_3446,N_3100);
and U3848 (N_3848,N_3113,N_3361);
and U3849 (N_3849,N_3290,N_3365);
and U3850 (N_3850,N_3478,N_3375);
nor U3851 (N_3851,N_3002,N_3297);
and U3852 (N_3852,N_3214,N_3346);
and U3853 (N_3853,N_3343,N_3219);
nand U3854 (N_3854,N_3333,N_3479);
xnor U3855 (N_3855,N_3431,N_3364);
xnor U3856 (N_3856,N_3301,N_3234);
and U3857 (N_3857,N_3468,N_3117);
xor U3858 (N_3858,N_3151,N_3122);
xnor U3859 (N_3859,N_3185,N_3475);
and U3860 (N_3860,N_3134,N_3123);
xor U3861 (N_3861,N_3448,N_3477);
nand U3862 (N_3862,N_3392,N_3295);
nand U3863 (N_3863,N_3067,N_3016);
or U3864 (N_3864,N_3444,N_3404);
nor U3865 (N_3865,N_3113,N_3490);
xor U3866 (N_3866,N_3268,N_3433);
and U3867 (N_3867,N_3483,N_3205);
nor U3868 (N_3868,N_3293,N_3019);
and U3869 (N_3869,N_3387,N_3041);
nor U3870 (N_3870,N_3306,N_3250);
or U3871 (N_3871,N_3082,N_3455);
nor U3872 (N_3872,N_3148,N_3212);
nor U3873 (N_3873,N_3304,N_3118);
nor U3874 (N_3874,N_3027,N_3423);
or U3875 (N_3875,N_3427,N_3273);
and U3876 (N_3876,N_3111,N_3185);
nor U3877 (N_3877,N_3334,N_3286);
or U3878 (N_3878,N_3015,N_3366);
nand U3879 (N_3879,N_3280,N_3478);
xnor U3880 (N_3880,N_3131,N_3421);
and U3881 (N_3881,N_3460,N_3304);
nor U3882 (N_3882,N_3150,N_3098);
xnor U3883 (N_3883,N_3392,N_3283);
nor U3884 (N_3884,N_3449,N_3006);
and U3885 (N_3885,N_3254,N_3136);
nand U3886 (N_3886,N_3215,N_3046);
xnor U3887 (N_3887,N_3154,N_3295);
xnor U3888 (N_3888,N_3191,N_3039);
nor U3889 (N_3889,N_3491,N_3290);
nand U3890 (N_3890,N_3297,N_3192);
xnor U3891 (N_3891,N_3176,N_3224);
nor U3892 (N_3892,N_3447,N_3175);
or U3893 (N_3893,N_3309,N_3137);
xnor U3894 (N_3894,N_3165,N_3075);
xnor U3895 (N_3895,N_3120,N_3204);
xor U3896 (N_3896,N_3324,N_3037);
nand U3897 (N_3897,N_3150,N_3329);
xor U3898 (N_3898,N_3114,N_3130);
xnor U3899 (N_3899,N_3196,N_3405);
nand U3900 (N_3900,N_3425,N_3463);
and U3901 (N_3901,N_3180,N_3372);
and U3902 (N_3902,N_3198,N_3143);
xnor U3903 (N_3903,N_3390,N_3019);
or U3904 (N_3904,N_3237,N_3263);
nand U3905 (N_3905,N_3144,N_3301);
or U3906 (N_3906,N_3194,N_3319);
or U3907 (N_3907,N_3353,N_3411);
nor U3908 (N_3908,N_3203,N_3348);
nand U3909 (N_3909,N_3228,N_3181);
and U3910 (N_3910,N_3155,N_3032);
or U3911 (N_3911,N_3497,N_3260);
nor U3912 (N_3912,N_3231,N_3019);
nand U3913 (N_3913,N_3303,N_3006);
or U3914 (N_3914,N_3151,N_3228);
nand U3915 (N_3915,N_3326,N_3286);
nand U3916 (N_3916,N_3493,N_3459);
xor U3917 (N_3917,N_3441,N_3199);
and U3918 (N_3918,N_3396,N_3342);
nor U3919 (N_3919,N_3366,N_3379);
nor U3920 (N_3920,N_3032,N_3450);
nor U3921 (N_3921,N_3416,N_3053);
xnor U3922 (N_3922,N_3363,N_3105);
xnor U3923 (N_3923,N_3367,N_3199);
nand U3924 (N_3924,N_3025,N_3194);
and U3925 (N_3925,N_3209,N_3091);
xor U3926 (N_3926,N_3386,N_3109);
nand U3927 (N_3927,N_3239,N_3012);
nor U3928 (N_3928,N_3413,N_3024);
nand U3929 (N_3929,N_3027,N_3108);
or U3930 (N_3930,N_3116,N_3205);
nor U3931 (N_3931,N_3359,N_3341);
nor U3932 (N_3932,N_3441,N_3205);
xnor U3933 (N_3933,N_3040,N_3285);
xnor U3934 (N_3934,N_3233,N_3145);
and U3935 (N_3935,N_3177,N_3379);
nand U3936 (N_3936,N_3453,N_3021);
nor U3937 (N_3937,N_3461,N_3057);
or U3938 (N_3938,N_3450,N_3070);
nor U3939 (N_3939,N_3406,N_3043);
nor U3940 (N_3940,N_3195,N_3496);
xor U3941 (N_3941,N_3279,N_3466);
or U3942 (N_3942,N_3024,N_3305);
nand U3943 (N_3943,N_3495,N_3187);
or U3944 (N_3944,N_3038,N_3077);
xnor U3945 (N_3945,N_3447,N_3400);
or U3946 (N_3946,N_3266,N_3412);
and U3947 (N_3947,N_3247,N_3150);
xnor U3948 (N_3948,N_3252,N_3230);
nand U3949 (N_3949,N_3172,N_3004);
and U3950 (N_3950,N_3173,N_3348);
nand U3951 (N_3951,N_3433,N_3220);
nand U3952 (N_3952,N_3137,N_3349);
nand U3953 (N_3953,N_3056,N_3001);
xnor U3954 (N_3954,N_3411,N_3164);
nor U3955 (N_3955,N_3448,N_3153);
nor U3956 (N_3956,N_3310,N_3475);
or U3957 (N_3957,N_3011,N_3138);
nand U3958 (N_3958,N_3029,N_3409);
xnor U3959 (N_3959,N_3178,N_3288);
and U3960 (N_3960,N_3179,N_3089);
nor U3961 (N_3961,N_3467,N_3333);
nand U3962 (N_3962,N_3130,N_3032);
xor U3963 (N_3963,N_3006,N_3387);
or U3964 (N_3964,N_3128,N_3044);
or U3965 (N_3965,N_3020,N_3129);
nand U3966 (N_3966,N_3442,N_3032);
and U3967 (N_3967,N_3286,N_3175);
and U3968 (N_3968,N_3097,N_3017);
nor U3969 (N_3969,N_3489,N_3206);
nor U3970 (N_3970,N_3032,N_3288);
and U3971 (N_3971,N_3473,N_3421);
nor U3972 (N_3972,N_3322,N_3193);
nor U3973 (N_3973,N_3462,N_3051);
or U3974 (N_3974,N_3054,N_3339);
nor U3975 (N_3975,N_3208,N_3049);
xor U3976 (N_3976,N_3210,N_3305);
and U3977 (N_3977,N_3454,N_3270);
and U3978 (N_3978,N_3278,N_3001);
or U3979 (N_3979,N_3235,N_3401);
xnor U3980 (N_3980,N_3340,N_3314);
or U3981 (N_3981,N_3402,N_3413);
nor U3982 (N_3982,N_3349,N_3018);
xor U3983 (N_3983,N_3410,N_3206);
nor U3984 (N_3984,N_3457,N_3253);
xor U3985 (N_3985,N_3021,N_3435);
nand U3986 (N_3986,N_3263,N_3079);
and U3987 (N_3987,N_3352,N_3493);
xor U3988 (N_3988,N_3292,N_3407);
or U3989 (N_3989,N_3266,N_3439);
xnor U3990 (N_3990,N_3159,N_3180);
xor U3991 (N_3991,N_3241,N_3404);
and U3992 (N_3992,N_3087,N_3469);
nor U3993 (N_3993,N_3073,N_3490);
xor U3994 (N_3994,N_3494,N_3496);
xor U3995 (N_3995,N_3102,N_3018);
and U3996 (N_3996,N_3236,N_3461);
and U3997 (N_3997,N_3377,N_3352);
xnor U3998 (N_3998,N_3074,N_3314);
xnor U3999 (N_3999,N_3246,N_3394);
or U4000 (N_4000,N_3610,N_3948);
nor U4001 (N_4001,N_3826,N_3972);
xnor U4002 (N_4002,N_3821,N_3785);
xor U4003 (N_4003,N_3879,N_3678);
nand U4004 (N_4004,N_3900,N_3712);
xor U4005 (N_4005,N_3582,N_3630);
xnor U4006 (N_4006,N_3771,N_3860);
or U4007 (N_4007,N_3650,N_3578);
xnor U4008 (N_4008,N_3933,N_3534);
nand U4009 (N_4009,N_3721,N_3543);
nand U4010 (N_4010,N_3736,N_3985);
xnor U4011 (N_4011,N_3554,N_3802);
xnor U4012 (N_4012,N_3844,N_3761);
or U4013 (N_4013,N_3926,N_3586);
nor U4014 (N_4014,N_3507,N_3853);
or U4015 (N_4015,N_3648,N_3904);
and U4016 (N_4016,N_3697,N_3838);
or U4017 (N_4017,N_3791,N_3541);
or U4018 (N_4018,N_3855,N_3835);
nand U4019 (N_4019,N_3868,N_3684);
and U4020 (N_4020,N_3703,N_3544);
and U4021 (N_4021,N_3576,N_3790);
nand U4022 (N_4022,N_3639,N_3929);
xor U4023 (N_4023,N_3606,N_3612);
or U4024 (N_4024,N_3695,N_3661);
nor U4025 (N_4025,N_3741,N_3865);
nand U4026 (N_4026,N_3866,N_3622);
xnor U4027 (N_4027,N_3524,N_3694);
and U4028 (N_4028,N_3573,N_3773);
and U4029 (N_4029,N_3980,N_3881);
nor U4030 (N_4030,N_3581,N_3618);
and U4031 (N_4031,N_3979,N_3729);
nor U4032 (N_4032,N_3696,N_3869);
nand U4033 (N_4033,N_3583,N_3940);
xor U4034 (N_4034,N_3803,N_3861);
and U4035 (N_4035,N_3913,N_3911);
or U4036 (N_4036,N_3997,N_3545);
xnor U4037 (N_4037,N_3594,N_3934);
xor U4038 (N_4038,N_3845,N_3537);
xnor U4039 (N_4039,N_3525,N_3782);
nand U4040 (N_4040,N_3636,N_3956);
nor U4041 (N_4041,N_3964,N_3723);
or U4042 (N_4042,N_3863,N_3779);
and U4043 (N_4043,N_3688,N_3804);
nand U4044 (N_4044,N_3704,N_3888);
xor U4045 (N_4045,N_3994,N_3500);
xnor U4046 (N_4046,N_3579,N_3658);
and U4047 (N_4047,N_3664,N_3959);
or U4048 (N_4048,N_3936,N_3671);
nor U4049 (N_4049,N_3722,N_3589);
nor U4050 (N_4050,N_3814,N_3669);
or U4051 (N_4051,N_3825,N_3757);
nor U4052 (N_4052,N_3982,N_3841);
xnor U4053 (N_4053,N_3530,N_3725);
nand U4054 (N_4054,N_3760,N_3724);
nand U4055 (N_4055,N_3914,N_3574);
nor U4056 (N_4056,N_3572,N_3735);
and U4057 (N_4057,N_3717,N_3990);
xnor U4058 (N_4058,N_3986,N_3877);
nor U4059 (N_4059,N_3522,N_3852);
xor U4060 (N_4060,N_3727,N_3607);
nor U4061 (N_4061,N_3854,N_3520);
or U4062 (N_4062,N_3691,N_3508);
nand U4063 (N_4063,N_3649,N_3905);
and U4064 (N_4064,N_3859,N_3943);
nand U4065 (N_4065,N_3617,N_3796);
nand U4066 (N_4066,N_3909,N_3818);
nand U4067 (N_4067,N_3620,N_3693);
nor U4068 (N_4068,N_3864,N_3876);
xnor U4069 (N_4069,N_3756,N_3856);
nand U4070 (N_4070,N_3798,N_3754);
nand U4071 (N_4071,N_3631,N_3599);
or U4072 (N_4072,N_3647,N_3532);
and U4073 (N_4073,N_3941,N_3939);
and U4074 (N_4074,N_3775,N_3849);
nand U4075 (N_4075,N_3553,N_3969);
xor U4076 (N_4076,N_3840,N_3682);
nor U4077 (N_4077,N_3999,N_3906);
nand U4078 (N_4078,N_3820,N_3621);
nor U4079 (N_4079,N_3638,N_3983);
and U4080 (N_4080,N_3752,N_3800);
or U4081 (N_4081,N_3517,N_3958);
nand U4082 (N_4082,N_3737,N_3656);
or U4083 (N_4083,N_3659,N_3512);
nor U4084 (N_4084,N_3566,N_3733);
and U4085 (N_4085,N_3758,N_3787);
nand U4086 (N_4086,N_3542,N_3984);
xnor U4087 (N_4087,N_3673,N_3963);
or U4088 (N_4088,N_3885,N_3968);
or U4089 (N_4089,N_3720,N_3558);
xnor U4090 (N_4090,N_3884,N_3609);
nand U4091 (N_4091,N_3588,N_3768);
xor U4092 (N_4092,N_3946,N_3922);
xor U4093 (N_4093,N_3872,N_3942);
or U4094 (N_4094,N_3827,N_3731);
or U4095 (N_4095,N_3992,N_3732);
or U4096 (N_4096,N_3742,N_3960);
xor U4097 (N_4097,N_3966,N_3891);
nor U4098 (N_4098,N_3931,N_3910);
xnor U4099 (N_4099,N_3561,N_3812);
and U4100 (N_4100,N_3944,N_3570);
or U4101 (N_4101,N_3778,N_3847);
and U4102 (N_4102,N_3924,N_3726);
xor U4103 (N_4103,N_3753,N_3679);
or U4104 (N_4104,N_3952,N_3998);
nor U4105 (N_4105,N_3886,N_3614);
nand U4106 (N_4106,N_3837,N_3632);
or U4107 (N_4107,N_3672,N_3975);
nor U4108 (N_4108,N_3625,N_3894);
and U4109 (N_4109,N_3813,N_3692);
nand U4110 (N_4110,N_3832,N_3899);
or U4111 (N_4111,N_3681,N_3957);
nand U4112 (N_4112,N_3738,N_3591);
and U4113 (N_4113,N_3509,N_3575);
nor U4114 (N_4114,N_3751,N_3815);
nand U4115 (N_4115,N_3536,N_3836);
nand U4116 (N_4116,N_3858,N_3557);
nor U4117 (N_4117,N_3862,N_3605);
and U4118 (N_4118,N_3502,N_3590);
and U4119 (N_4119,N_3700,N_3627);
nand U4120 (N_4120,N_3764,N_3531);
xor U4121 (N_4121,N_3555,N_3674);
or U4122 (N_4122,N_3623,N_3817);
nand U4123 (N_4123,N_3938,N_3521);
nand U4124 (N_4124,N_3792,N_3846);
nand U4125 (N_4125,N_3719,N_3547);
nand U4126 (N_4126,N_3867,N_3597);
or U4127 (N_4127,N_3875,N_3784);
xnor U4128 (N_4128,N_3641,N_3970);
nor U4129 (N_4129,N_3670,N_3713);
xnor U4130 (N_4130,N_3564,N_3908);
nand U4131 (N_4131,N_3585,N_3923);
nor U4132 (N_4132,N_3925,N_3795);
nor U4133 (N_4133,N_3645,N_3539);
or U4134 (N_4134,N_3513,N_3907);
nand U4135 (N_4135,N_3893,N_3897);
or U4136 (N_4136,N_3635,N_3668);
nor U4137 (N_4137,N_3971,N_3708);
nand U4138 (N_4138,N_3552,N_3637);
nand U4139 (N_4139,N_3951,N_3828);
and U4140 (N_4140,N_3538,N_3823);
nand U4141 (N_4141,N_3608,N_3560);
nor U4142 (N_4142,N_3950,N_3976);
xnor U4143 (N_4143,N_3546,N_3794);
nand U4144 (N_4144,N_3715,N_3967);
and U4145 (N_4145,N_3718,N_3780);
and U4146 (N_4146,N_3662,N_3519);
and U4147 (N_4147,N_3624,N_3710);
xnor U4148 (N_4148,N_3776,N_3699);
nand U4149 (N_4149,N_3805,N_3932);
or U4150 (N_4150,N_3686,N_3523);
nor U4151 (N_4151,N_3902,N_3880);
or U4152 (N_4152,N_3857,N_3730);
nor U4153 (N_4153,N_3947,N_3748);
xor U4154 (N_4154,N_3680,N_3501);
nor U4155 (N_4155,N_3954,N_3824);
or U4156 (N_4156,N_3653,N_3604);
and U4157 (N_4157,N_3766,N_3991);
nor U4158 (N_4158,N_3919,N_3706);
or U4159 (N_4159,N_3799,N_3830);
or U4160 (N_4160,N_3548,N_3615);
and U4161 (N_4161,N_3831,N_3644);
and U4162 (N_4162,N_3961,N_3642);
nand U4163 (N_4163,N_3613,N_3709);
and U4164 (N_4164,N_3598,N_3660);
xor U4165 (N_4165,N_3556,N_3666);
nor U4166 (N_4166,N_3981,N_3810);
nor U4167 (N_4167,N_3774,N_3870);
nand U4168 (N_4168,N_3740,N_3759);
or U4169 (N_4169,N_3626,N_3750);
xnor U4170 (N_4170,N_3928,N_3901);
nand U4171 (N_4171,N_3667,N_3807);
or U4172 (N_4172,N_3628,N_3993);
or U4173 (N_4173,N_3788,N_3716);
or U4174 (N_4174,N_3734,N_3611);
and U4175 (N_4175,N_3580,N_3739);
or U4176 (N_4176,N_3744,N_3707);
nand U4177 (N_4177,N_3789,N_3749);
nor U4178 (N_4178,N_3685,N_3781);
nand U4179 (N_4179,N_3510,N_3930);
or U4180 (N_4180,N_3777,N_3848);
nor U4181 (N_4181,N_3833,N_3883);
nor U4182 (N_4182,N_3569,N_3786);
xor U4183 (N_4183,N_3746,N_3801);
xor U4184 (N_4184,N_3915,N_3701);
xnor U4185 (N_4185,N_3955,N_3743);
nor U4186 (N_4186,N_3528,N_3829);
nand U4187 (N_4187,N_3714,N_3987);
or U4188 (N_4188,N_3651,N_3895);
nor U4189 (N_4189,N_3655,N_3903);
or U4190 (N_4190,N_3505,N_3745);
and U4191 (N_4191,N_3677,N_3962);
nand U4192 (N_4192,N_3878,N_3965);
nand U4193 (N_4193,N_3596,N_3917);
nor U4194 (N_4194,N_3765,N_3973);
and U4195 (N_4195,N_3592,N_3887);
xnor U4196 (N_4196,N_3978,N_3629);
nand U4197 (N_4197,N_3595,N_3996);
nor U4198 (N_4198,N_3518,N_3563);
nand U4199 (N_4199,N_3584,N_3698);
nor U4200 (N_4200,N_3702,N_3892);
nand U4201 (N_4201,N_3526,N_3806);
xor U4202 (N_4202,N_3770,N_3811);
nor U4203 (N_4203,N_3889,N_3550);
nor U4204 (N_4204,N_3603,N_3945);
or U4205 (N_4205,N_3949,N_3977);
xor U4206 (N_4206,N_3654,N_3797);
and U4207 (N_4207,N_3504,N_3874);
and U4208 (N_4208,N_3772,N_3747);
or U4209 (N_4209,N_3690,N_3587);
nor U4210 (N_4210,N_3600,N_3871);
nor U4211 (N_4211,N_3619,N_3640);
or U4212 (N_4212,N_3665,N_3882);
nand U4213 (N_4213,N_3646,N_3529);
nand U4214 (N_4214,N_3562,N_3515);
or U4215 (N_4215,N_3809,N_3514);
nor U4216 (N_4216,N_3974,N_3593);
nand U4217 (N_4217,N_3602,N_3989);
nand U4218 (N_4218,N_3559,N_3676);
or U4219 (N_4219,N_3793,N_3808);
or U4220 (N_4220,N_3988,N_3912);
nor U4221 (N_4221,N_3898,N_3937);
xor U4222 (N_4222,N_3920,N_3540);
xor U4223 (N_4223,N_3896,N_3567);
nor U4224 (N_4224,N_3842,N_3839);
or U4225 (N_4225,N_3767,N_3571);
xnor U4226 (N_4226,N_3850,N_3675);
nor U4227 (N_4227,N_3728,N_3873);
nor U4228 (N_4228,N_3890,N_3551);
nand U4229 (N_4229,N_3601,N_3783);
or U4230 (N_4230,N_3511,N_3921);
nor U4231 (N_4231,N_3843,N_3916);
or U4232 (N_4232,N_3687,N_3834);
or U4233 (N_4233,N_3927,N_3516);
or U4234 (N_4234,N_3643,N_3527);
nor U4235 (N_4235,N_3816,N_3663);
nand U4236 (N_4236,N_3769,N_3577);
nor U4237 (N_4237,N_3918,N_3705);
nor U4238 (N_4238,N_3535,N_3689);
nand U4239 (N_4239,N_3633,N_3763);
nor U4240 (N_4240,N_3533,N_3683);
nand U4241 (N_4241,N_3616,N_3953);
xor U4242 (N_4242,N_3819,N_3506);
and U4243 (N_4243,N_3755,N_3634);
and U4244 (N_4244,N_3822,N_3503);
nor U4245 (N_4245,N_3549,N_3995);
or U4246 (N_4246,N_3568,N_3711);
nand U4247 (N_4247,N_3565,N_3935);
xor U4248 (N_4248,N_3657,N_3762);
or U4249 (N_4249,N_3851,N_3652);
xnor U4250 (N_4250,N_3658,N_3664);
nand U4251 (N_4251,N_3672,N_3831);
xor U4252 (N_4252,N_3686,N_3803);
nand U4253 (N_4253,N_3886,N_3916);
and U4254 (N_4254,N_3760,N_3755);
or U4255 (N_4255,N_3609,N_3973);
xor U4256 (N_4256,N_3577,N_3569);
nand U4257 (N_4257,N_3726,N_3526);
nor U4258 (N_4258,N_3912,N_3552);
or U4259 (N_4259,N_3932,N_3508);
nand U4260 (N_4260,N_3902,N_3761);
nand U4261 (N_4261,N_3975,N_3569);
nor U4262 (N_4262,N_3674,N_3917);
nand U4263 (N_4263,N_3964,N_3678);
nand U4264 (N_4264,N_3803,N_3611);
xnor U4265 (N_4265,N_3731,N_3793);
or U4266 (N_4266,N_3837,N_3939);
and U4267 (N_4267,N_3780,N_3880);
nand U4268 (N_4268,N_3780,N_3928);
or U4269 (N_4269,N_3891,N_3548);
xor U4270 (N_4270,N_3776,N_3545);
or U4271 (N_4271,N_3775,N_3966);
and U4272 (N_4272,N_3714,N_3527);
nand U4273 (N_4273,N_3941,N_3753);
xor U4274 (N_4274,N_3768,N_3650);
nand U4275 (N_4275,N_3682,N_3632);
nand U4276 (N_4276,N_3610,N_3978);
or U4277 (N_4277,N_3718,N_3877);
and U4278 (N_4278,N_3639,N_3936);
xnor U4279 (N_4279,N_3514,N_3561);
xnor U4280 (N_4280,N_3555,N_3516);
nand U4281 (N_4281,N_3854,N_3506);
xor U4282 (N_4282,N_3701,N_3907);
or U4283 (N_4283,N_3847,N_3696);
nand U4284 (N_4284,N_3917,N_3741);
nand U4285 (N_4285,N_3786,N_3863);
nor U4286 (N_4286,N_3979,N_3529);
nor U4287 (N_4287,N_3697,N_3814);
or U4288 (N_4288,N_3650,N_3534);
and U4289 (N_4289,N_3656,N_3654);
and U4290 (N_4290,N_3745,N_3870);
xnor U4291 (N_4291,N_3696,N_3824);
and U4292 (N_4292,N_3976,N_3734);
nand U4293 (N_4293,N_3689,N_3874);
or U4294 (N_4294,N_3622,N_3927);
nor U4295 (N_4295,N_3856,N_3843);
or U4296 (N_4296,N_3597,N_3935);
xnor U4297 (N_4297,N_3829,N_3519);
xor U4298 (N_4298,N_3543,N_3517);
nand U4299 (N_4299,N_3640,N_3904);
nand U4300 (N_4300,N_3553,N_3745);
and U4301 (N_4301,N_3834,N_3555);
and U4302 (N_4302,N_3781,N_3801);
nor U4303 (N_4303,N_3846,N_3834);
nor U4304 (N_4304,N_3996,N_3809);
xor U4305 (N_4305,N_3691,N_3966);
xnor U4306 (N_4306,N_3935,N_3555);
nand U4307 (N_4307,N_3936,N_3564);
xnor U4308 (N_4308,N_3951,N_3745);
or U4309 (N_4309,N_3689,N_3606);
or U4310 (N_4310,N_3754,N_3976);
xor U4311 (N_4311,N_3700,N_3686);
xor U4312 (N_4312,N_3695,N_3868);
or U4313 (N_4313,N_3738,N_3950);
xor U4314 (N_4314,N_3615,N_3722);
nand U4315 (N_4315,N_3758,N_3921);
nand U4316 (N_4316,N_3842,N_3826);
xor U4317 (N_4317,N_3845,N_3751);
or U4318 (N_4318,N_3822,N_3732);
nor U4319 (N_4319,N_3765,N_3724);
and U4320 (N_4320,N_3732,N_3552);
nor U4321 (N_4321,N_3996,N_3721);
nand U4322 (N_4322,N_3562,N_3532);
nor U4323 (N_4323,N_3758,N_3929);
xnor U4324 (N_4324,N_3801,N_3760);
xor U4325 (N_4325,N_3556,N_3604);
nor U4326 (N_4326,N_3743,N_3935);
or U4327 (N_4327,N_3639,N_3598);
nand U4328 (N_4328,N_3663,N_3549);
nor U4329 (N_4329,N_3998,N_3862);
and U4330 (N_4330,N_3748,N_3527);
nor U4331 (N_4331,N_3934,N_3630);
and U4332 (N_4332,N_3657,N_3948);
or U4333 (N_4333,N_3718,N_3977);
nor U4334 (N_4334,N_3713,N_3705);
xor U4335 (N_4335,N_3898,N_3995);
and U4336 (N_4336,N_3506,N_3892);
nand U4337 (N_4337,N_3513,N_3923);
nor U4338 (N_4338,N_3598,N_3579);
nand U4339 (N_4339,N_3613,N_3714);
nor U4340 (N_4340,N_3792,N_3892);
xor U4341 (N_4341,N_3973,N_3510);
or U4342 (N_4342,N_3800,N_3990);
nand U4343 (N_4343,N_3976,N_3932);
nor U4344 (N_4344,N_3634,N_3850);
and U4345 (N_4345,N_3981,N_3761);
or U4346 (N_4346,N_3510,N_3922);
nand U4347 (N_4347,N_3651,N_3535);
nor U4348 (N_4348,N_3748,N_3741);
or U4349 (N_4349,N_3588,N_3543);
nor U4350 (N_4350,N_3510,N_3860);
or U4351 (N_4351,N_3738,N_3675);
or U4352 (N_4352,N_3588,N_3508);
or U4353 (N_4353,N_3869,N_3683);
or U4354 (N_4354,N_3969,N_3565);
xnor U4355 (N_4355,N_3517,N_3558);
nor U4356 (N_4356,N_3770,N_3949);
and U4357 (N_4357,N_3912,N_3904);
or U4358 (N_4358,N_3946,N_3729);
nand U4359 (N_4359,N_3549,N_3986);
nor U4360 (N_4360,N_3881,N_3910);
or U4361 (N_4361,N_3512,N_3572);
nor U4362 (N_4362,N_3708,N_3974);
and U4363 (N_4363,N_3511,N_3635);
xnor U4364 (N_4364,N_3896,N_3777);
nor U4365 (N_4365,N_3880,N_3982);
xnor U4366 (N_4366,N_3756,N_3892);
nand U4367 (N_4367,N_3579,N_3583);
nor U4368 (N_4368,N_3918,N_3685);
or U4369 (N_4369,N_3590,N_3914);
nor U4370 (N_4370,N_3846,N_3584);
and U4371 (N_4371,N_3803,N_3869);
nor U4372 (N_4372,N_3766,N_3736);
xnor U4373 (N_4373,N_3776,N_3973);
and U4374 (N_4374,N_3634,N_3992);
or U4375 (N_4375,N_3581,N_3998);
nor U4376 (N_4376,N_3877,N_3764);
xor U4377 (N_4377,N_3922,N_3758);
or U4378 (N_4378,N_3947,N_3848);
or U4379 (N_4379,N_3551,N_3950);
nand U4380 (N_4380,N_3821,N_3673);
xnor U4381 (N_4381,N_3913,N_3595);
xor U4382 (N_4382,N_3842,N_3877);
nor U4383 (N_4383,N_3768,N_3970);
and U4384 (N_4384,N_3710,N_3990);
nand U4385 (N_4385,N_3656,N_3713);
nand U4386 (N_4386,N_3725,N_3990);
nor U4387 (N_4387,N_3971,N_3729);
nand U4388 (N_4388,N_3762,N_3986);
nor U4389 (N_4389,N_3712,N_3902);
xnor U4390 (N_4390,N_3513,N_3618);
xnor U4391 (N_4391,N_3950,N_3864);
or U4392 (N_4392,N_3503,N_3601);
nor U4393 (N_4393,N_3830,N_3706);
and U4394 (N_4394,N_3722,N_3979);
xnor U4395 (N_4395,N_3901,N_3793);
or U4396 (N_4396,N_3856,N_3655);
nor U4397 (N_4397,N_3715,N_3794);
or U4398 (N_4398,N_3632,N_3907);
nand U4399 (N_4399,N_3585,N_3788);
and U4400 (N_4400,N_3527,N_3581);
or U4401 (N_4401,N_3882,N_3981);
nand U4402 (N_4402,N_3617,N_3702);
and U4403 (N_4403,N_3816,N_3951);
nor U4404 (N_4404,N_3930,N_3763);
or U4405 (N_4405,N_3551,N_3635);
xor U4406 (N_4406,N_3723,N_3724);
or U4407 (N_4407,N_3999,N_3929);
xnor U4408 (N_4408,N_3904,N_3983);
and U4409 (N_4409,N_3534,N_3802);
nand U4410 (N_4410,N_3688,N_3867);
xor U4411 (N_4411,N_3883,N_3706);
xor U4412 (N_4412,N_3856,N_3739);
or U4413 (N_4413,N_3535,N_3865);
or U4414 (N_4414,N_3973,N_3987);
or U4415 (N_4415,N_3732,N_3618);
or U4416 (N_4416,N_3713,N_3975);
nand U4417 (N_4417,N_3983,N_3933);
nor U4418 (N_4418,N_3921,N_3603);
xor U4419 (N_4419,N_3848,N_3632);
or U4420 (N_4420,N_3837,N_3605);
nand U4421 (N_4421,N_3656,N_3941);
or U4422 (N_4422,N_3569,N_3678);
xor U4423 (N_4423,N_3959,N_3814);
or U4424 (N_4424,N_3914,N_3836);
nor U4425 (N_4425,N_3899,N_3866);
xnor U4426 (N_4426,N_3714,N_3682);
nor U4427 (N_4427,N_3684,N_3544);
or U4428 (N_4428,N_3925,N_3743);
nand U4429 (N_4429,N_3741,N_3796);
xor U4430 (N_4430,N_3921,N_3683);
xor U4431 (N_4431,N_3741,N_3817);
nand U4432 (N_4432,N_3640,N_3502);
or U4433 (N_4433,N_3851,N_3758);
nor U4434 (N_4434,N_3702,N_3638);
nand U4435 (N_4435,N_3547,N_3988);
xnor U4436 (N_4436,N_3923,N_3582);
xnor U4437 (N_4437,N_3938,N_3820);
nor U4438 (N_4438,N_3550,N_3816);
nand U4439 (N_4439,N_3578,N_3814);
xor U4440 (N_4440,N_3705,N_3848);
nand U4441 (N_4441,N_3899,N_3810);
xnor U4442 (N_4442,N_3994,N_3884);
xnor U4443 (N_4443,N_3855,N_3838);
nor U4444 (N_4444,N_3773,N_3985);
and U4445 (N_4445,N_3790,N_3808);
xor U4446 (N_4446,N_3602,N_3926);
nand U4447 (N_4447,N_3741,N_3970);
and U4448 (N_4448,N_3955,N_3795);
and U4449 (N_4449,N_3543,N_3954);
and U4450 (N_4450,N_3875,N_3771);
nand U4451 (N_4451,N_3760,N_3878);
xnor U4452 (N_4452,N_3523,N_3534);
nor U4453 (N_4453,N_3526,N_3897);
and U4454 (N_4454,N_3573,N_3792);
nand U4455 (N_4455,N_3781,N_3802);
and U4456 (N_4456,N_3960,N_3696);
xor U4457 (N_4457,N_3579,N_3756);
nor U4458 (N_4458,N_3961,N_3635);
or U4459 (N_4459,N_3627,N_3694);
xor U4460 (N_4460,N_3847,N_3534);
xor U4461 (N_4461,N_3658,N_3599);
nand U4462 (N_4462,N_3634,N_3772);
xor U4463 (N_4463,N_3874,N_3611);
or U4464 (N_4464,N_3737,N_3707);
xor U4465 (N_4465,N_3720,N_3951);
or U4466 (N_4466,N_3548,N_3863);
nand U4467 (N_4467,N_3877,N_3901);
nand U4468 (N_4468,N_3868,N_3739);
nand U4469 (N_4469,N_3875,N_3566);
xnor U4470 (N_4470,N_3664,N_3513);
nand U4471 (N_4471,N_3858,N_3985);
xor U4472 (N_4472,N_3834,N_3849);
xor U4473 (N_4473,N_3823,N_3750);
and U4474 (N_4474,N_3938,N_3874);
nand U4475 (N_4475,N_3565,N_3658);
and U4476 (N_4476,N_3590,N_3980);
or U4477 (N_4477,N_3618,N_3701);
xnor U4478 (N_4478,N_3943,N_3927);
xnor U4479 (N_4479,N_3754,N_3995);
nand U4480 (N_4480,N_3885,N_3647);
or U4481 (N_4481,N_3788,N_3989);
xor U4482 (N_4482,N_3824,N_3798);
nand U4483 (N_4483,N_3881,N_3945);
nand U4484 (N_4484,N_3889,N_3775);
xnor U4485 (N_4485,N_3771,N_3507);
nand U4486 (N_4486,N_3898,N_3892);
or U4487 (N_4487,N_3637,N_3922);
and U4488 (N_4488,N_3571,N_3559);
and U4489 (N_4489,N_3934,N_3635);
or U4490 (N_4490,N_3717,N_3602);
or U4491 (N_4491,N_3940,N_3506);
and U4492 (N_4492,N_3735,N_3630);
and U4493 (N_4493,N_3928,N_3515);
or U4494 (N_4494,N_3698,N_3717);
nor U4495 (N_4495,N_3836,N_3919);
xnor U4496 (N_4496,N_3854,N_3789);
nand U4497 (N_4497,N_3847,N_3596);
nor U4498 (N_4498,N_3842,N_3574);
and U4499 (N_4499,N_3599,N_3815);
and U4500 (N_4500,N_4349,N_4207);
nor U4501 (N_4501,N_4430,N_4445);
and U4502 (N_4502,N_4378,N_4222);
or U4503 (N_4503,N_4201,N_4146);
or U4504 (N_4504,N_4015,N_4488);
and U4505 (N_4505,N_4240,N_4336);
xor U4506 (N_4506,N_4099,N_4475);
and U4507 (N_4507,N_4069,N_4265);
nand U4508 (N_4508,N_4022,N_4266);
nand U4509 (N_4509,N_4320,N_4221);
nand U4510 (N_4510,N_4354,N_4351);
and U4511 (N_4511,N_4389,N_4101);
nor U4512 (N_4512,N_4420,N_4193);
and U4513 (N_4513,N_4299,N_4048);
xnor U4514 (N_4514,N_4197,N_4142);
and U4515 (N_4515,N_4318,N_4186);
and U4516 (N_4516,N_4411,N_4128);
and U4517 (N_4517,N_4010,N_4412);
xor U4518 (N_4518,N_4074,N_4208);
nand U4519 (N_4519,N_4437,N_4084);
xor U4520 (N_4520,N_4245,N_4458);
nand U4521 (N_4521,N_4111,N_4493);
or U4522 (N_4522,N_4305,N_4310);
and U4523 (N_4523,N_4397,N_4108);
xor U4524 (N_4524,N_4243,N_4161);
xor U4525 (N_4525,N_4492,N_4017);
nor U4526 (N_4526,N_4147,N_4055);
and U4527 (N_4527,N_4306,N_4263);
xor U4528 (N_4528,N_4394,N_4052);
or U4529 (N_4529,N_4482,N_4477);
nand U4530 (N_4530,N_4214,N_4089);
xor U4531 (N_4531,N_4148,N_4220);
nand U4532 (N_4532,N_4296,N_4380);
xor U4533 (N_4533,N_4273,N_4041);
nand U4534 (N_4534,N_4433,N_4345);
or U4535 (N_4535,N_4171,N_4417);
nand U4536 (N_4536,N_4036,N_4016);
nand U4537 (N_4537,N_4153,N_4129);
xnor U4538 (N_4538,N_4331,N_4029);
and U4539 (N_4539,N_4086,N_4205);
nor U4540 (N_4540,N_4091,N_4409);
nand U4541 (N_4541,N_4377,N_4063);
xnor U4542 (N_4542,N_4313,N_4003);
nand U4543 (N_4543,N_4210,N_4230);
xor U4544 (N_4544,N_4044,N_4151);
xor U4545 (N_4545,N_4100,N_4189);
nor U4546 (N_4546,N_4032,N_4115);
or U4547 (N_4547,N_4013,N_4035);
or U4548 (N_4548,N_4157,N_4190);
nand U4549 (N_4549,N_4059,N_4117);
nor U4550 (N_4550,N_4355,N_4158);
nor U4551 (N_4551,N_4384,N_4172);
and U4552 (N_4552,N_4167,N_4046);
nor U4553 (N_4553,N_4049,N_4102);
xor U4554 (N_4554,N_4238,N_4322);
nor U4555 (N_4555,N_4133,N_4436);
nor U4556 (N_4556,N_4302,N_4196);
nand U4557 (N_4557,N_4116,N_4457);
nor U4558 (N_4558,N_4490,N_4034);
and U4559 (N_4559,N_4056,N_4346);
xor U4560 (N_4560,N_4070,N_4300);
xor U4561 (N_4561,N_4042,N_4427);
xor U4562 (N_4562,N_4379,N_4469);
nand U4563 (N_4563,N_4050,N_4082);
xor U4564 (N_4564,N_4043,N_4183);
nor U4565 (N_4565,N_4474,N_4261);
nor U4566 (N_4566,N_4260,N_4314);
nand U4567 (N_4567,N_4062,N_4339);
xnor U4568 (N_4568,N_4040,N_4264);
xnor U4569 (N_4569,N_4472,N_4159);
nand U4570 (N_4570,N_4256,N_4223);
and U4571 (N_4571,N_4288,N_4195);
xor U4572 (N_4572,N_4203,N_4291);
nor U4573 (N_4573,N_4149,N_4467);
nor U4574 (N_4574,N_4473,N_4415);
and U4575 (N_4575,N_4438,N_4136);
and U4576 (N_4576,N_4249,N_4143);
nor U4577 (N_4577,N_4400,N_4166);
xnor U4578 (N_4578,N_4145,N_4232);
or U4579 (N_4579,N_4225,N_4418);
or U4580 (N_4580,N_4200,N_4154);
xor U4581 (N_4581,N_4303,N_4247);
xnor U4582 (N_4582,N_4434,N_4293);
nand U4583 (N_4583,N_4138,N_4316);
or U4584 (N_4584,N_4294,N_4267);
or U4585 (N_4585,N_4104,N_4095);
nand U4586 (N_4586,N_4061,N_4374);
and U4587 (N_4587,N_4065,N_4463);
or U4588 (N_4588,N_4150,N_4485);
xor U4589 (N_4589,N_4376,N_4077);
xor U4590 (N_4590,N_4386,N_4276);
and U4591 (N_4591,N_4275,N_4290);
or U4592 (N_4592,N_4182,N_4404);
xor U4593 (N_4593,N_4323,N_4449);
xor U4594 (N_4594,N_4371,N_4068);
nor U4595 (N_4595,N_4370,N_4385);
xor U4596 (N_4596,N_4058,N_4357);
xor U4597 (N_4597,N_4093,N_4483);
or U4598 (N_4598,N_4399,N_4423);
or U4599 (N_4599,N_4484,N_4004);
nand U4600 (N_4600,N_4496,N_4144);
nand U4601 (N_4601,N_4164,N_4359);
xnor U4602 (N_4602,N_4448,N_4312);
or U4603 (N_4603,N_4461,N_4368);
nor U4604 (N_4604,N_4255,N_4227);
and U4605 (N_4605,N_4217,N_4254);
nor U4606 (N_4606,N_4421,N_4155);
nor U4607 (N_4607,N_4039,N_4373);
or U4608 (N_4608,N_4090,N_4343);
nor U4609 (N_4609,N_4206,N_4466);
or U4610 (N_4610,N_4465,N_4092);
or U4611 (N_4611,N_4011,N_4124);
xnor U4612 (N_4612,N_4076,N_4403);
nand U4613 (N_4613,N_4367,N_4067);
nor U4614 (N_4614,N_4361,N_4495);
xnor U4615 (N_4615,N_4080,N_4226);
nand U4616 (N_4616,N_4185,N_4350);
nand U4617 (N_4617,N_4248,N_4491);
nor U4618 (N_4618,N_4441,N_4381);
and U4619 (N_4619,N_4025,N_4277);
nor U4620 (N_4620,N_4447,N_4321);
nand U4621 (N_4621,N_4340,N_4204);
nand U4622 (N_4622,N_4066,N_4250);
nor U4623 (N_4623,N_4088,N_4324);
nand U4624 (N_4624,N_4252,N_4218);
or U4625 (N_4625,N_4352,N_4459);
nand U4626 (N_4626,N_4237,N_4301);
xor U4627 (N_4627,N_4216,N_4442);
or U4628 (N_4628,N_4008,N_4413);
xor U4629 (N_4629,N_4363,N_4118);
nand U4630 (N_4630,N_4338,N_4071);
and U4631 (N_4631,N_4372,N_4173);
nor U4632 (N_4632,N_4175,N_4045);
xnor U4633 (N_4633,N_4019,N_4060);
xor U4634 (N_4634,N_4038,N_4282);
nand U4635 (N_4635,N_4219,N_4356);
xor U4636 (N_4636,N_4298,N_4194);
xnor U4637 (N_4637,N_4396,N_4072);
xor U4638 (N_4638,N_4094,N_4083);
nor U4639 (N_4639,N_4137,N_4215);
xnor U4640 (N_4640,N_4271,N_4253);
or U4641 (N_4641,N_4439,N_4122);
xor U4642 (N_4642,N_4317,N_4168);
and U4643 (N_4643,N_4431,N_4358);
or U4644 (N_4644,N_4307,N_4410);
nand U4645 (N_4645,N_4191,N_4470);
or U4646 (N_4646,N_4342,N_4181);
xor U4647 (N_4647,N_4236,N_4366);
or U4648 (N_4648,N_4251,N_4486);
nand U4649 (N_4649,N_4494,N_4235);
nand U4650 (N_4650,N_4353,N_4177);
nand U4651 (N_4651,N_4462,N_4012);
or U4652 (N_4652,N_4234,N_4390);
xnor U4653 (N_4653,N_4244,N_4212);
xnor U4654 (N_4654,N_4114,N_4471);
nor U4655 (N_4655,N_4387,N_4304);
nor U4656 (N_4656,N_4454,N_4481);
or U4657 (N_4657,N_4174,N_4156);
and U4658 (N_4658,N_4416,N_4152);
nor U4659 (N_4659,N_4053,N_4364);
or U4660 (N_4660,N_4333,N_4269);
nor U4661 (N_4661,N_4229,N_4480);
nand U4662 (N_4662,N_4383,N_4451);
nand U4663 (N_4663,N_4281,N_4239);
or U4664 (N_4664,N_4362,N_4257);
or U4665 (N_4665,N_4435,N_4075);
and U4666 (N_4666,N_4308,N_4408);
nand U4667 (N_4667,N_4406,N_4393);
nor U4668 (N_4668,N_4369,N_4132);
xor U4669 (N_4669,N_4391,N_4130);
nand U4670 (N_4670,N_4401,N_4005);
or U4671 (N_4671,N_4107,N_4178);
nand U4672 (N_4672,N_4424,N_4279);
nor U4673 (N_4673,N_4024,N_4228);
xnor U4674 (N_4674,N_4453,N_4382);
nor U4675 (N_4675,N_4140,N_4329);
nor U4676 (N_4676,N_4468,N_4139);
and U4677 (N_4677,N_4425,N_4319);
or U4678 (N_4678,N_4037,N_4344);
nor U4679 (N_4679,N_4169,N_4162);
nand U4680 (N_4680,N_4028,N_4270);
or U4681 (N_4681,N_4452,N_4414);
xor U4682 (N_4682,N_4365,N_4007);
nand U4683 (N_4683,N_4078,N_4487);
nand U4684 (N_4684,N_4213,N_4478);
and U4685 (N_4685,N_4284,N_4341);
and U4686 (N_4686,N_4160,N_4297);
xor U4687 (N_4687,N_4476,N_4064);
xnor U4688 (N_4688,N_4426,N_4335);
xor U4689 (N_4689,N_4311,N_4163);
nor U4690 (N_4690,N_4272,N_4428);
or U4691 (N_4691,N_4443,N_4398);
nand U4692 (N_4692,N_4327,N_4405);
nor U4693 (N_4693,N_4006,N_4112);
and U4694 (N_4694,N_4199,N_4274);
and U4695 (N_4695,N_4258,N_4280);
and U4696 (N_4696,N_4106,N_4334);
or U4697 (N_4697,N_4202,N_4119);
xnor U4698 (N_4698,N_4109,N_4031);
or U4699 (N_4699,N_4096,N_4033);
xnor U4700 (N_4700,N_4192,N_4021);
nor U4701 (N_4701,N_4002,N_4315);
nor U4702 (N_4702,N_4141,N_4287);
nor U4703 (N_4703,N_4444,N_4464);
xnor U4704 (N_4704,N_4026,N_4054);
and U4705 (N_4705,N_4000,N_4268);
xor U4706 (N_4706,N_4120,N_4198);
nand U4707 (N_4707,N_4047,N_4392);
xnor U4708 (N_4708,N_4020,N_4081);
xor U4709 (N_4709,N_4499,N_4231);
nand U4710 (N_4710,N_4242,N_4450);
and U4711 (N_4711,N_4209,N_4233);
or U4712 (N_4712,N_4030,N_4347);
or U4713 (N_4713,N_4429,N_4224);
or U4714 (N_4714,N_4211,N_4460);
xnor U4715 (N_4715,N_4134,N_4422);
nand U4716 (N_4716,N_4079,N_4085);
xor U4717 (N_4717,N_4489,N_4184);
xor U4718 (N_4718,N_4375,N_4001);
or U4719 (N_4719,N_4326,N_4103);
and U4720 (N_4720,N_4023,N_4057);
nor U4721 (N_4721,N_4407,N_4246);
nor U4722 (N_4722,N_4395,N_4497);
xnor U4723 (N_4723,N_4309,N_4176);
xor U4724 (N_4724,N_4360,N_4170);
nor U4725 (N_4725,N_4498,N_4087);
and U4726 (N_4726,N_4330,N_4180);
nor U4727 (N_4727,N_4325,N_4123);
xor U4728 (N_4728,N_4337,N_4328);
and U4729 (N_4729,N_4440,N_4097);
and U4730 (N_4730,N_4121,N_4295);
or U4731 (N_4731,N_4456,N_4014);
nand U4732 (N_4732,N_4446,N_4127);
nand U4733 (N_4733,N_4388,N_4286);
and U4734 (N_4734,N_4126,N_4027);
and U4735 (N_4735,N_4283,N_4188);
or U4736 (N_4736,N_4131,N_4165);
nor U4737 (N_4737,N_4332,N_4073);
or U4738 (N_4738,N_4432,N_4113);
nand U4739 (N_4739,N_4018,N_4110);
or U4740 (N_4740,N_4292,N_4241);
xor U4741 (N_4741,N_4259,N_4402);
nor U4742 (N_4742,N_4098,N_4187);
nand U4743 (N_4743,N_4278,N_4179);
xor U4744 (N_4744,N_4285,N_4262);
or U4745 (N_4745,N_4125,N_4105);
xnor U4746 (N_4746,N_4135,N_4348);
and U4747 (N_4747,N_4419,N_4009);
nand U4748 (N_4748,N_4455,N_4051);
and U4749 (N_4749,N_4479,N_4289);
nor U4750 (N_4750,N_4079,N_4185);
or U4751 (N_4751,N_4008,N_4120);
xor U4752 (N_4752,N_4039,N_4471);
or U4753 (N_4753,N_4224,N_4072);
or U4754 (N_4754,N_4009,N_4474);
nand U4755 (N_4755,N_4302,N_4070);
and U4756 (N_4756,N_4020,N_4057);
xnor U4757 (N_4757,N_4029,N_4491);
nand U4758 (N_4758,N_4152,N_4304);
xnor U4759 (N_4759,N_4152,N_4316);
xnor U4760 (N_4760,N_4240,N_4322);
or U4761 (N_4761,N_4063,N_4285);
nand U4762 (N_4762,N_4335,N_4162);
and U4763 (N_4763,N_4146,N_4037);
xor U4764 (N_4764,N_4487,N_4322);
and U4765 (N_4765,N_4458,N_4173);
xor U4766 (N_4766,N_4283,N_4191);
or U4767 (N_4767,N_4482,N_4273);
nand U4768 (N_4768,N_4461,N_4005);
nand U4769 (N_4769,N_4042,N_4469);
and U4770 (N_4770,N_4366,N_4362);
nor U4771 (N_4771,N_4421,N_4469);
or U4772 (N_4772,N_4184,N_4402);
or U4773 (N_4773,N_4493,N_4057);
nor U4774 (N_4774,N_4167,N_4288);
or U4775 (N_4775,N_4390,N_4455);
xor U4776 (N_4776,N_4092,N_4073);
and U4777 (N_4777,N_4313,N_4291);
or U4778 (N_4778,N_4089,N_4294);
and U4779 (N_4779,N_4036,N_4240);
or U4780 (N_4780,N_4494,N_4492);
nand U4781 (N_4781,N_4047,N_4128);
and U4782 (N_4782,N_4161,N_4350);
or U4783 (N_4783,N_4151,N_4033);
nor U4784 (N_4784,N_4392,N_4198);
nor U4785 (N_4785,N_4473,N_4482);
and U4786 (N_4786,N_4027,N_4179);
xor U4787 (N_4787,N_4220,N_4370);
nor U4788 (N_4788,N_4295,N_4378);
and U4789 (N_4789,N_4070,N_4458);
nor U4790 (N_4790,N_4388,N_4391);
nor U4791 (N_4791,N_4183,N_4417);
and U4792 (N_4792,N_4399,N_4335);
nor U4793 (N_4793,N_4024,N_4464);
or U4794 (N_4794,N_4049,N_4261);
nor U4795 (N_4795,N_4163,N_4076);
or U4796 (N_4796,N_4196,N_4082);
or U4797 (N_4797,N_4487,N_4472);
nand U4798 (N_4798,N_4302,N_4354);
nand U4799 (N_4799,N_4089,N_4332);
nand U4800 (N_4800,N_4462,N_4245);
xnor U4801 (N_4801,N_4420,N_4135);
or U4802 (N_4802,N_4184,N_4412);
nor U4803 (N_4803,N_4284,N_4247);
and U4804 (N_4804,N_4463,N_4104);
and U4805 (N_4805,N_4128,N_4496);
nand U4806 (N_4806,N_4415,N_4489);
xnor U4807 (N_4807,N_4072,N_4469);
or U4808 (N_4808,N_4406,N_4160);
xor U4809 (N_4809,N_4228,N_4453);
and U4810 (N_4810,N_4177,N_4430);
nand U4811 (N_4811,N_4209,N_4383);
nand U4812 (N_4812,N_4237,N_4405);
nor U4813 (N_4813,N_4324,N_4338);
or U4814 (N_4814,N_4291,N_4135);
xor U4815 (N_4815,N_4392,N_4485);
or U4816 (N_4816,N_4053,N_4354);
nor U4817 (N_4817,N_4439,N_4127);
or U4818 (N_4818,N_4355,N_4005);
and U4819 (N_4819,N_4351,N_4424);
or U4820 (N_4820,N_4375,N_4023);
or U4821 (N_4821,N_4235,N_4398);
and U4822 (N_4822,N_4326,N_4131);
xor U4823 (N_4823,N_4179,N_4370);
nor U4824 (N_4824,N_4182,N_4348);
or U4825 (N_4825,N_4324,N_4490);
xor U4826 (N_4826,N_4147,N_4337);
nand U4827 (N_4827,N_4421,N_4094);
nor U4828 (N_4828,N_4076,N_4224);
nor U4829 (N_4829,N_4051,N_4399);
xnor U4830 (N_4830,N_4127,N_4487);
xor U4831 (N_4831,N_4079,N_4468);
nand U4832 (N_4832,N_4343,N_4345);
and U4833 (N_4833,N_4111,N_4426);
xnor U4834 (N_4834,N_4061,N_4262);
nand U4835 (N_4835,N_4211,N_4273);
nand U4836 (N_4836,N_4278,N_4470);
xnor U4837 (N_4837,N_4224,N_4354);
nor U4838 (N_4838,N_4491,N_4059);
and U4839 (N_4839,N_4045,N_4457);
xnor U4840 (N_4840,N_4210,N_4491);
xnor U4841 (N_4841,N_4380,N_4204);
nor U4842 (N_4842,N_4433,N_4273);
and U4843 (N_4843,N_4083,N_4061);
xnor U4844 (N_4844,N_4414,N_4430);
and U4845 (N_4845,N_4491,N_4207);
xor U4846 (N_4846,N_4494,N_4467);
or U4847 (N_4847,N_4362,N_4316);
and U4848 (N_4848,N_4291,N_4490);
and U4849 (N_4849,N_4330,N_4340);
nand U4850 (N_4850,N_4466,N_4452);
xor U4851 (N_4851,N_4428,N_4174);
xor U4852 (N_4852,N_4282,N_4073);
nor U4853 (N_4853,N_4487,N_4359);
and U4854 (N_4854,N_4430,N_4381);
nand U4855 (N_4855,N_4140,N_4199);
or U4856 (N_4856,N_4234,N_4213);
xnor U4857 (N_4857,N_4242,N_4184);
xor U4858 (N_4858,N_4295,N_4450);
nor U4859 (N_4859,N_4435,N_4019);
or U4860 (N_4860,N_4451,N_4107);
xor U4861 (N_4861,N_4310,N_4253);
xor U4862 (N_4862,N_4178,N_4462);
xnor U4863 (N_4863,N_4330,N_4112);
xnor U4864 (N_4864,N_4207,N_4377);
or U4865 (N_4865,N_4149,N_4250);
nor U4866 (N_4866,N_4138,N_4144);
and U4867 (N_4867,N_4112,N_4390);
or U4868 (N_4868,N_4189,N_4336);
or U4869 (N_4869,N_4182,N_4279);
nand U4870 (N_4870,N_4107,N_4201);
or U4871 (N_4871,N_4070,N_4160);
nand U4872 (N_4872,N_4383,N_4262);
xnor U4873 (N_4873,N_4164,N_4364);
or U4874 (N_4874,N_4313,N_4187);
xnor U4875 (N_4875,N_4316,N_4468);
nor U4876 (N_4876,N_4103,N_4020);
xor U4877 (N_4877,N_4179,N_4499);
nand U4878 (N_4878,N_4222,N_4009);
and U4879 (N_4879,N_4192,N_4027);
xnor U4880 (N_4880,N_4121,N_4240);
nand U4881 (N_4881,N_4111,N_4155);
or U4882 (N_4882,N_4242,N_4061);
nand U4883 (N_4883,N_4245,N_4351);
and U4884 (N_4884,N_4158,N_4265);
or U4885 (N_4885,N_4245,N_4170);
and U4886 (N_4886,N_4039,N_4263);
nor U4887 (N_4887,N_4376,N_4369);
or U4888 (N_4888,N_4232,N_4495);
or U4889 (N_4889,N_4385,N_4033);
xnor U4890 (N_4890,N_4268,N_4329);
or U4891 (N_4891,N_4298,N_4315);
and U4892 (N_4892,N_4151,N_4206);
nand U4893 (N_4893,N_4351,N_4294);
xor U4894 (N_4894,N_4308,N_4347);
or U4895 (N_4895,N_4227,N_4072);
nor U4896 (N_4896,N_4257,N_4103);
nor U4897 (N_4897,N_4203,N_4437);
nor U4898 (N_4898,N_4075,N_4253);
and U4899 (N_4899,N_4392,N_4237);
nand U4900 (N_4900,N_4058,N_4139);
xnor U4901 (N_4901,N_4283,N_4346);
nand U4902 (N_4902,N_4398,N_4306);
or U4903 (N_4903,N_4408,N_4030);
nand U4904 (N_4904,N_4233,N_4485);
nand U4905 (N_4905,N_4193,N_4023);
nor U4906 (N_4906,N_4088,N_4031);
xor U4907 (N_4907,N_4141,N_4201);
or U4908 (N_4908,N_4133,N_4325);
nor U4909 (N_4909,N_4317,N_4433);
nor U4910 (N_4910,N_4072,N_4037);
nor U4911 (N_4911,N_4355,N_4233);
nand U4912 (N_4912,N_4207,N_4459);
or U4913 (N_4913,N_4319,N_4288);
or U4914 (N_4914,N_4239,N_4296);
nand U4915 (N_4915,N_4110,N_4117);
xor U4916 (N_4916,N_4067,N_4290);
xnor U4917 (N_4917,N_4302,N_4007);
or U4918 (N_4918,N_4084,N_4435);
or U4919 (N_4919,N_4007,N_4169);
xnor U4920 (N_4920,N_4372,N_4352);
xor U4921 (N_4921,N_4319,N_4372);
or U4922 (N_4922,N_4352,N_4006);
or U4923 (N_4923,N_4468,N_4256);
and U4924 (N_4924,N_4286,N_4312);
nand U4925 (N_4925,N_4013,N_4072);
nand U4926 (N_4926,N_4419,N_4244);
xnor U4927 (N_4927,N_4019,N_4332);
and U4928 (N_4928,N_4450,N_4055);
nand U4929 (N_4929,N_4387,N_4375);
nand U4930 (N_4930,N_4423,N_4089);
and U4931 (N_4931,N_4078,N_4080);
and U4932 (N_4932,N_4135,N_4230);
and U4933 (N_4933,N_4395,N_4462);
nor U4934 (N_4934,N_4467,N_4453);
nor U4935 (N_4935,N_4085,N_4475);
and U4936 (N_4936,N_4329,N_4248);
xor U4937 (N_4937,N_4078,N_4290);
xor U4938 (N_4938,N_4498,N_4308);
nand U4939 (N_4939,N_4222,N_4284);
xnor U4940 (N_4940,N_4296,N_4394);
xnor U4941 (N_4941,N_4341,N_4051);
nand U4942 (N_4942,N_4391,N_4213);
nor U4943 (N_4943,N_4408,N_4084);
or U4944 (N_4944,N_4477,N_4215);
and U4945 (N_4945,N_4002,N_4231);
and U4946 (N_4946,N_4352,N_4351);
xnor U4947 (N_4947,N_4086,N_4165);
nor U4948 (N_4948,N_4389,N_4286);
and U4949 (N_4949,N_4037,N_4189);
nand U4950 (N_4950,N_4045,N_4453);
or U4951 (N_4951,N_4424,N_4220);
or U4952 (N_4952,N_4088,N_4438);
nor U4953 (N_4953,N_4435,N_4148);
nand U4954 (N_4954,N_4020,N_4226);
and U4955 (N_4955,N_4495,N_4157);
nor U4956 (N_4956,N_4484,N_4338);
nand U4957 (N_4957,N_4412,N_4066);
and U4958 (N_4958,N_4452,N_4036);
or U4959 (N_4959,N_4153,N_4274);
or U4960 (N_4960,N_4005,N_4378);
and U4961 (N_4961,N_4138,N_4082);
nand U4962 (N_4962,N_4140,N_4050);
xnor U4963 (N_4963,N_4290,N_4043);
xor U4964 (N_4964,N_4381,N_4245);
xnor U4965 (N_4965,N_4027,N_4483);
and U4966 (N_4966,N_4337,N_4448);
xor U4967 (N_4967,N_4206,N_4452);
xor U4968 (N_4968,N_4013,N_4194);
nand U4969 (N_4969,N_4000,N_4219);
and U4970 (N_4970,N_4119,N_4273);
xor U4971 (N_4971,N_4089,N_4102);
and U4972 (N_4972,N_4409,N_4104);
nor U4973 (N_4973,N_4332,N_4265);
nor U4974 (N_4974,N_4482,N_4347);
and U4975 (N_4975,N_4484,N_4082);
nand U4976 (N_4976,N_4127,N_4453);
nand U4977 (N_4977,N_4197,N_4410);
nor U4978 (N_4978,N_4332,N_4058);
nand U4979 (N_4979,N_4123,N_4408);
nand U4980 (N_4980,N_4011,N_4304);
nand U4981 (N_4981,N_4496,N_4184);
or U4982 (N_4982,N_4205,N_4124);
xnor U4983 (N_4983,N_4285,N_4060);
xor U4984 (N_4984,N_4053,N_4334);
or U4985 (N_4985,N_4302,N_4118);
nor U4986 (N_4986,N_4082,N_4389);
or U4987 (N_4987,N_4350,N_4466);
or U4988 (N_4988,N_4110,N_4242);
or U4989 (N_4989,N_4337,N_4462);
or U4990 (N_4990,N_4012,N_4030);
and U4991 (N_4991,N_4033,N_4421);
or U4992 (N_4992,N_4487,N_4148);
or U4993 (N_4993,N_4229,N_4465);
and U4994 (N_4994,N_4364,N_4252);
nand U4995 (N_4995,N_4386,N_4407);
xor U4996 (N_4996,N_4167,N_4051);
xnor U4997 (N_4997,N_4035,N_4342);
and U4998 (N_4998,N_4170,N_4451);
or U4999 (N_4999,N_4200,N_4350);
or U5000 (N_5000,N_4717,N_4906);
nand U5001 (N_5001,N_4968,N_4962);
nand U5002 (N_5002,N_4935,N_4514);
nor U5003 (N_5003,N_4722,N_4917);
nor U5004 (N_5004,N_4716,N_4829);
or U5005 (N_5005,N_4837,N_4539);
nand U5006 (N_5006,N_4546,N_4573);
or U5007 (N_5007,N_4768,N_4886);
or U5008 (N_5008,N_4934,N_4729);
or U5009 (N_5009,N_4859,N_4647);
xnor U5010 (N_5010,N_4506,N_4736);
or U5011 (N_5011,N_4614,N_4732);
nand U5012 (N_5012,N_4791,N_4952);
nand U5013 (N_5013,N_4684,N_4590);
nor U5014 (N_5014,N_4788,N_4845);
or U5015 (N_5015,N_4510,N_4844);
xnor U5016 (N_5016,N_4687,N_4712);
xor U5017 (N_5017,N_4621,N_4942);
or U5018 (N_5018,N_4867,N_4508);
nand U5019 (N_5019,N_4554,N_4578);
and U5020 (N_5020,N_4612,N_4737);
xnor U5021 (N_5021,N_4725,N_4946);
or U5022 (N_5022,N_4750,N_4600);
or U5023 (N_5023,N_4629,N_4957);
or U5024 (N_5024,N_4599,N_4607);
nand U5025 (N_5025,N_4511,N_4615);
or U5026 (N_5026,N_4792,N_4756);
xnor U5027 (N_5027,N_4985,N_4515);
and U5028 (N_5028,N_4727,N_4733);
or U5029 (N_5029,N_4770,N_4806);
nor U5030 (N_5030,N_4964,N_4709);
or U5031 (N_5031,N_4826,N_4929);
or U5032 (N_5032,N_4780,N_4742);
nand U5033 (N_5033,N_4537,N_4698);
xor U5034 (N_5034,N_4993,N_4778);
and U5035 (N_5035,N_4943,N_4601);
or U5036 (N_5036,N_4741,N_4526);
and U5037 (N_5037,N_4828,N_4821);
nand U5038 (N_5038,N_4623,N_4931);
nor U5039 (N_5039,N_4823,N_4719);
or U5040 (N_5040,N_4919,N_4730);
or U5041 (N_5041,N_4790,N_4670);
nor U5042 (N_5042,N_4852,N_4521);
nand U5043 (N_5043,N_4998,N_4914);
nor U5044 (N_5044,N_4881,N_4916);
nand U5045 (N_5045,N_4619,N_4793);
nand U5046 (N_5046,N_4992,N_4609);
xor U5047 (N_5047,N_4787,N_4691);
xor U5048 (N_5048,N_4873,N_4561);
xnor U5049 (N_5049,N_4635,N_4933);
xor U5050 (N_5050,N_4813,N_4830);
or U5051 (N_5051,N_4569,N_4882);
nand U5052 (N_5052,N_4827,N_4699);
xnor U5053 (N_5053,N_4755,N_4786);
and U5054 (N_5054,N_4901,N_4707);
and U5055 (N_5055,N_4804,N_4972);
nand U5056 (N_5056,N_4738,N_4944);
nand U5057 (N_5057,N_4721,N_4803);
and U5058 (N_5058,N_4883,N_4863);
and U5059 (N_5059,N_4949,N_4678);
xor U5060 (N_5060,N_4855,N_4524);
nor U5061 (N_5061,N_4613,N_4555);
and U5062 (N_5062,N_4660,N_4956);
nand U5063 (N_5063,N_4978,N_4587);
and U5064 (N_5064,N_4889,N_4961);
xnor U5065 (N_5065,N_4825,N_4564);
xor U5066 (N_5066,N_4584,N_4885);
or U5067 (N_5067,N_4645,N_4950);
or U5068 (N_5068,N_4891,N_4566);
or U5069 (N_5069,N_4834,N_4651);
xnor U5070 (N_5070,N_4870,N_4657);
nor U5071 (N_5071,N_4988,N_4631);
or U5072 (N_5072,N_4525,N_4986);
and U5073 (N_5073,N_4617,N_4689);
and U5074 (N_5074,N_4688,N_4577);
and U5075 (N_5075,N_4708,N_4533);
nor U5076 (N_5076,N_4954,N_4763);
nor U5077 (N_5077,N_4588,N_4802);
xnor U5078 (N_5078,N_4560,N_4766);
and U5079 (N_5079,N_4912,N_4849);
or U5080 (N_5080,N_4783,N_4580);
or U5081 (N_5081,N_4582,N_4746);
xnor U5082 (N_5082,N_4663,N_4749);
or U5083 (N_5083,N_4692,N_4853);
nand U5084 (N_5084,N_4936,N_4846);
xnor U5085 (N_5085,N_4734,N_4711);
and U5086 (N_5086,N_4974,N_4981);
nor U5087 (N_5087,N_4851,N_4715);
xor U5088 (N_5088,N_4996,N_4502);
xor U5089 (N_5089,N_4743,N_4926);
nand U5090 (N_5090,N_4810,N_4757);
nand U5091 (N_5091,N_4748,N_4864);
nor U5092 (N_5092,N_4579,N_4505);
xor U5093 (N_5093,N_4562,N_4527);
nand U5094 (N_5094,N_4809,N_4948);
nand U5095 (N_5095,N_4900,N_4928);
and U5096 (N_5096,N_4745,N_4841);
and U5097 (N_5097,N_4666,N_4685);
nand U5098 (N_5098,N_4634,N_4536);
nor U5099 (N_5099,N_4632,N_4983);
nor U5100 (N_5100,N_4905,N_4528);
and U5101 (N_5101,N_4747,N_4694);
or U5102 (N_5102,N_4547,N_4695);
xor U5103 (N_5103,N_4517,N_4927);
nand U5104 (N_5104,N_4907,N_4606);
xor U5105 (N_5105,N_4913,N_4989);
nor U5106 (N_5106,N_4626,N_4958);
and U5107 (N_5107,N_4642,N_4503);
and U5108 (N_5108,N_4611,N_4622);
or U5109 (N_5109,N_4690,N_4535);
or U5110 (N_5110,N_4581,N_4824);
nand U5111 (N_5111,N_4897,N_4960);
and U5112 (N_5112,N_4697,N_4764);
nand U5113 (N_5113,N_4625,N_4572);
and U5114 (N_5114,N_4909,N_4641);
or U5115 (N_5115,N_4673,N_4682);
nand U5116 (N_5116,N_4876,N_4610);
nor U5117 (N_5117,N_4710,N_4575);
or U5118 (N_5118,N_4973,N_4520);
nor U5119 (N_5119,N_4620,N_4676);
and U5120 (N_5120,N_4596,N_4571);
nand U5121 (N_5121,N_4899,N_4618);
xor U5122 (N_5122,N_4879,N_4649);
xnor U5123 (N_5123,N_4800,N_4661);
nor U5124 (N_5124,N_4924,N_4677);
and U5125 (N_5125,N_4822,N_4977);
or U5126 (N_5126,N_4723,N_4713);
nand U5127 (N_5127,N_4875,N_4898);
xnor U5128 (N_5128,N_4516,N_4656);
nor U5129 (N_5129,N_4781,N_4534);
xnor U5130 (N_5130,N_4593,N_4874);
nand U5131 (N_5131,N_4818,N_4541);
xor U5132 (N_5132,N_4976,N_4653);
xor U5133 (N_5133,N_4565,N_4808);
or U5134 (N_5134,N_4843,N_4947);
nor U5135 (N_5135,N_4967,N_4784);
nand U5136 (N_5136,N_4604,N_4718);
nand U5137 (N_5137,N_4728,N_4815);
or U5138 (N_5138,N_4671,N_4854);
nor U5139 (N_5139,N_4878,N_4807);
or U5140 (N_5140,N_4814,N_4598);
and U5141 (N_5141,N_4769,N_4938);
and U5142 (N_5142,N_4819,N_4595);
and U5143 (N_5143,N_4556,N_4568);
nand U5144 (N_5144,N_4777,N_4762);
xnor U5145 (N_5145,N_4731,N_4591);
nor U5146 (N_5146,N_4840,N_4911);
nor U5147 (N_5147,N_4668,N_4925);
nor U5148 (N_5148,N_4662,N_4820);
xor U5149 (N_5149,N_4785,N_4920);
xor U5150 (N_5150,N_4811,N_4500);
and U5151 (N_5151,N_4551,N_4754);
and U5152 (N_5152,N_4563,N_4842);
xnor U5153 (N_5153,N_4744,N_4979);
or U5154 (N_5154,N_4558,N_4872);
xor U5155 (N_5155,N_4548,N_4772);
nor U5156 (N_5156,N_4586,N_4639);
and U5157 (N_5157,N_4550,N_4965);
nand U5158 (N_5158,N_4616,N_4765);
nand U5159 (N_5159,N_4799,N_4549);
nand U5160 (N_5160,N_4894,N_4759);
nor U5161 (N_5161,N_4848,N_4890);
or U5162 (N_5162,N_4608,N_4805);
nor U5163 (N_5163,N_4969,N_4892);
nor U5164 (N_5164,N_4951,N_4628);
nand U5165 (N_5165,N_4760,N_4816);
or U5166 (N_5166,N_4739,N_4908);
nor U5167 (N_5167,N_4589,N_4839);
and U5168 (N_5168,N_4995,N_4970);
xor U5169 (N_5169,N_4726,N_4939);
and U5170 (N_5170,N_4831,N_4658);
and U5171 (N_5171,N_4518,N_4735);
or U5172 (N_5172,N_4774,N_4888);
xnor U5173 (N_5173,N_4833,N_4861);
xnor U5174 (N_5174,N_4513,N_4963);
or U5175 (N_5175,N_4990,N_4940);
or U5176 (N_5176,N_4838,N_4922);
nand U5177 (N_5177,N_4672,N_4585);
nor U5178 (N_5178,N_4771,N_4576);
or U5179 (N_5179,N_4686,N_4557);
nand U5180 (N_5180,N_4531,N_4674);
or U5181 (N_5181,N_4869,N_4504);
nor U5182 (N_5182,N_4812,N_4636);
nand U5183 (N_5183,N_4543,N_4782);
nor U5184 (N_5184,N_4923,N_4857);
or U5185 (N_5185,N_4984,N_4910);
nand U5186 (N_5186,N_4798,N_4835);
and U5187 (N_5187,N_4696,N_4862);
xnor U5188 (N_5188,N_4507,N_4523);
or U5189 (N_5189,N_4630,N_4982);
and U5190 (N_5190,N_4866,N_4650);
or U5191 (N_5191,N_4544,N_4602);
nand U5192 (N_5192,N_4501,N_4794);
and U5193 (N_5193,N_4884,N_4776);
nor U5194 (N_5194,N_4999,N_4779);
nor U5195 (N_5195,N_4637,N_4654);
xnor U5196 (N_5196,N_4603,N_4644);
nand U5197 (N_5197,N_4592,N_4624);
or U5198 (N_5198,N_4646,N_4966);
and U5199 (N_5199,N_4532,N_4529);
nand U5200 (N_5200,N_4887,N_4959);
and U5201 (N_5201,N_4720,N_4937);
or U5202 (N_5202,N_4903,N_4703);
or U5203 (N_5203,N_4594,N_4918);
nor U5204 (N_5204,N_4761,N_4640);
nor U5205 (N_5205,N_4597,N_4655);
nor U5206 (N_5206,N_4795,N_4895);
or U5207 (N_5207,N_4583,N_4509);
or U5208 (N_5208,N_4789,N_4932);
and U5209 (N_5209,N_4991,N_4545);
and U5210 (N_5210,N_4701,N_4871);
and U5211 (N_5211,N_4856,N_4904);
and U5212 (N_5212,N_4850,N_4994);
nor U5213 (N_5213,N_4652,N_4740);
and U5214 (N_5214,N_4955,N_4775);
and U5215 (N_5215,N_4512,N_4773);
nand U5216 (N_5216,N_4858,N_4706);
nor U5217 (N_5217,N_4753,N_4797);
and U5218 (N_5218,N_4633,N_4680);
nor U5219 (N_5219,N_4542,N_4605);
nor U5220 (N_5220,N_4700,N_4648);
or U5221 (N_5221,N_4559,N_4627);
or U5222 (N_5222,N_4847,N_4553);
xnor U5223 (N_5223,N_4987,N_4638);
nand U5224 (N_5224,N_4683,N_4679);
nor U5225 (N_5225,N_4540,N_4675);
nor U5226 (N_5226,N_4801,N_4941);
or U5227 (N_5227,N_4643,N_4915);
nor U5228 (N_5228,N_4665,N_4832);
xor U5229 (N_5229,N_4836,N_4705);
or U5230 (N_5230,N_4567,N_4758);
and U5231 (N_5231,N_4860,N_4538);
nand U5232 (N_5232,N_4877,N_4865);
or U5233 (N_5233,N_4880,N_4702);
nand U5234 (N_5234,N_4817,N_4519);
xor U5235 (N_5235,N_4664,N_4980);
nor U5236 (N_5236,N_4669,N_4570);
or U5237 (N_5237,N_4667,N_4704);
or U5238 (N_5238,N_4659,N_4724);
or U5239 (N_5239,N_4751,N_4522);
nor U5240 (N_5240,N_4945,N_4693);
nor U5241 (N_5241,N_4997,N_4971);
or U5242 (N_5242,N_4902,N_4953);
or U5243 (N_5243,N_4752,N_4921);
nand U5244 (N_5244,N_4530,N_4796);
nand U5245 (N_5245,N_4868,N_4681);
nor U5246 (N_5246,N_4930,N_4893);
nand U5247 (N_5247,N_4975,N_4896);
nor U5248 (N_5248,N_4574,N_4714);
and U5249 (N_5249,N_4767,N_4552);
xnor U5250 (N_5250,N_4525,N_4895);
xnor U5251 (N_5251,N_4771,N_4682);
and U5252 (N_5252,N_4869,N_4764);
xor U5253 (N_5253,N_4544,N_4931);
nor U5254 (N_5254,N_4560,N_4889);
xor U5255 (N_5255,N_4804,N_4745);
nor U5256 (N_5256,N_4641,N_4645);
and U5257 (N_5257,N_4843,N_4523);
nor U5258 (N_5258,N_4706,N_4519);
xnor U5259 (N_5259,N_4830,N_4572);
nor U5260 (N_5260,N_4872,N_4975);
and U5261 (N_5261,N_4505,N_4827);
nor U5262 (N_5262,N_4856,N_4591);
or U5263 (N_5263,N_4742,N_4743);
or U5264 (N_5264,N_4873,N_4946);
or U5265 (N_5265,N_4829,N_4544);
nand U5266 (N_5266,N_4520,N_4611);
nand U5267 (N_5267,N_4792,N_4981);
xor U5268 (N_5268,N_4523,N_4864);
xnor U5269 (N_5269,N_4661,N_4781);
or U5270 (N_5270,N_4662,N_4892);
or U5271 (N_5271,N_4711,N_4577);
nor U5272 (N_5272,N_4881,N_4773);
nand U5273 (N_5273,N_4924,N_4515);
xor U5274 (N_5274,N_4836,N_4958);
or U5275 (N_5275,N_4519,N_4636);
xor U5276 (N_5276,N_4562,N_4983);
nand U5277 (N_5277,N_4987,N_4577);
or U5278 (N_5278,N_4831,N_4877);
and U5279 (N_5279,N_4581,N_4542);
nand U5280 (N_5280,N_4511,N_4739);
and U5281 (N_5281,N_4571,N_4665);
xor U5282 (N_5282,N_4806,N_4969);
or U5283 (N_5283,N_4577,N_4878);
and U5284 (N_5284,N_4623,N_4876);
and U5285 (N_5285,N_4508,N_4705);
and U5286 (N_5286,N_4789,N_4903);
or U5287 (N_5287,N_4997,N_4517);
xor U5288 (N_5288,N_4536,N_4949);
xor U5289 (N_5289,N_4823,N_4972);
nor U5290 (N_5290,N_4972,N_4577);
xnor U5291 (N_5291,N_4618,N_4700);
nand U5292 (N_5292,N_4646,N_4559);
and U5293 (N_5293,N_4726,N_4895);
or U5294 (N_5294,N_4940,N_4816);
xnor U5295 (N_5295,N_4651,N_4589);
and U5296 (N_5296,N_4573,N_4717);
xor U5297 (N_5297,N_4538,N_4975);
nor U5298 (N_5298,N_4766,N_4713);
nor U5299 (N_5299,N_4809,N_4625);
and U5300 (N_5300,N_4921,N_4849);
xnor U5301 (N_5301,N_4866,N_4726);
nor U5302 (N_5302,N_4666,N_4550);
nand U5303 (N_5303,N_4968,N_4754);
and U5304 (N_5304,N_4595,N_4996);
nand U5305 (N_5305,N_4881,N_4920);
nor U5306 (N_5306,N_4843,N_4996);
nand U5307 (N_5307,N_4942,N_4553);
and U5308 (N_5308,N_4622,N_4873);
nor U5309 (N_5309,N_4639,N_4522);
nor U5310 (N_5310,N_4639,N_4971);
or U5311 (N_5311,N_4707,N_4598);
nand U5312 (N_5312,N_4677,N_4998);
nand U5313 (N_5313,N_4805,N_4725);
nor U5314 (N_5314,N_4809,N_4526);
nor U5315 (N_5315,N_4912,N_4537);
xor U5316 (N_5316,N_4874,N_4997);
or U5317 (N_5317,N_4732,N_4559);
and U5318 (N_5318,N_4504,N_4854);
or U5319 (N_5319,N_4815,N_4804);
and U5320 (N_5320,N_4935,N_4869);
nor U5321 (N_5321,N_4812,N_4985);
and U5322 (N_5322,N_4597,N_4694);
or U5323 (N_5323,N_4722,N_4632);
xnor U5324 (N_5324,N_4838,N_4821);
nor U5325 (N_5325,N_4875,N_4760);
nor U5326 (N_5326,N_4606,N_4773);
xor U5327 (N_5327,N_4894,N_4915);
xnor U5328 (N_5328,N_4978,N_4971);
nor U5329 (N_5329,N_4517,N_4852);
xnor U5330 (N_5330,N_4687,N_4844);
or U5331 (N_5331,N_4985,N_4611);
nor U5332 (N_5332,N_4767,N_4817);
or U5333 (N_5333,N_4776,N_4753);
nand U5334 (N_5334,N_4586,N_4737);
and U5335 (N_5335,N_4520,N_4939);
xor U5336 (N_5336,N_4799,N_4885);
or U5337 (N_5337,N_4573,N_4508);
nor U5338 (N_5338,N_4673,N_4985);
nor U5339 (N_5339,N_4615,N_4763);
xnor U5340 (N_5340,N_4787,N_4690);
xor U5341 (N_5341,N_4719,N_4609);
and U5342 (N_5342,N_4818,N_4699);
and U5343 (N_5343,N_4675,N_4720);
and U5344 (N_5344,N_4753,N_4932);
nor U5345 (N_5345,N_4689,N_4867);
nand U5346 (N_5346,N_4691,N_4588);
xor U5347 (N_5347,N_4977,N_4859);
xor U5348 (N_5348,N_4790,N_4869);
nand U5349 (N_5349,N_4949,N_4850);
nand U5350 (N_5350,N_4608,N_4758);
and U5351 (N_5351,N_4652,N_4842);
xnor U5352 (N_5352,N_4858,N_4882);
and U5353 (N_5353,N_4744,N_4779);
nor U5354 (N_5354,N_4617,N_4603);
nand U5355 (N_5355,N_4812,N_4920);
nand U5356 (N_5356,N_4743,N_4990);
nand U5357 (N_5357,N_4628,N_4794);
or U5358 (N_5358,N_4559,N_4553);
and U5359 (N_5359,N_4593,N_4940);
nor U5360 (N_5360,N_4526,N_4924);
nor U5361 (N_5361,N_4513,N_4817);
xor U5362 (N_5362,N_4939,N_4513);
nand U5363 (N_5363,N_4891,N_4902);
xor U5364 (N_5364,N_4832,N_4921);
xnor U5365 (N_5365,N_4975,N_4752);
nor U5366 (N_5366,N_4884,N_4544);
or U5367 (N_5367,N_4662,N_4503);
xor U5368 (N_5368,N_4999,N_4994);
xnor U5369 (N_5369,N_4549,N_4727);
nor U5370 (N_5370,N_4813,N_4976);
xnor U5371 (N_5371,N_4760,N_4759);
xor U5372 (N_5372,N_4841,N_4658);
nor U5373 (N_5373,N_4683,N_4612);
nand U5374 (N_5374,N_4739,N_4502);
nand U5375 (N_5375,N_4957,N_4792);
nor U5376 (N_5376,N_4594,N_4680);
and U5377 (N_5377,N_4689,N_4891);
or U5378 (N_5378,N_4578,N_4617);
nand U5379 (N_5379,N_4678,N_4926);
and U5380 (N_5380,N_4989,N_4697);
and U5381 (N_5381,N_4813,N_4965);
nor U5382 (N_5382,N_4914,N_4594);
xor U5383 (N_5383,N_4729,N_4906);
xnor U5384 (N_5384,N_4908,N_4645);
or U5385 (N_5385,N_4893,N_4883);
or U5386 (N_5386,N_4522,N_4879);
nand U5387 (N_5387,N_4573,N_4722);
and U5388 (N_5388,N_4771,N_4546);
xor U5389 (N_5389,N_4597,N_4715);
or U5390 (N_5390,N_4565,N_4904);
nand U5391 (N_5391,N_4621,N_4813);
xor U5392 (N_5392,N_4547,N_4655);
and U5393 (N_5393,N_4700,N_4727);
xor U5394 (N_5394,N_4840,N_4783);
and U5395 (N_5395,N_4675,N_4914);
nand U5396 (N_5396,N_4943,N_4550);
or U5397 (N_5397,N_4756,N_4610);
nor U5398 (N_5398,N_4949,N_4737);
xnor U5399 (N_5399,N_4991,N_4847);
or U5400 (N_5400,N_4700,N_4815);
nand U5401 (N_5401,N_4531,N_4669);
nor U5402 (N_5402,N_4509,N_4903);
nand U5403 (N_5403,N_4525,N_4958);
nor U5404 (N_5404,N_4603,N_4588);
nor U5405 (N_5405,N_4674,N_4830);
xor U5406 (N_5406,N_4768,N_4649);
xor U5407 (N_5407,N_4811,N_4620);
or U5408 (N_5408,N_4533,N_4853);
nand U5409 (N_5409,N_4549,N_4617);
and U5410 (N_5410,N_4971,N_4628);
or U5411 (N_5411,N_4784,N_4965);
nand U5412 (N_5412,N_4725,N_4859);
xnor U5413 (N_5413,N_4981,N_4810);
nand U5414 (N_5414,N_4705,N_4671);
and U5415 (N_5415,N_4955,N_4516);
or U5416 (N_5416,N_4706,N_4786);
nand U5417 (N_5417,N_4867,N_4545);
xor U5418 (N_5418,N_4916,N_4575);
or U5419 (N_5419,N_4801,N_4699);
and U5420 (N_5420,N_4950,N_4786);
nand U5421 (N_5421,N_4729,N_4797);
nor U5422 (N_5422,N_4733,N_4605);
nand U5423 (N_5423,N_4996,N_4692);
nand U5424 (N_5424,N_4928,N_4530);
nand U5425 (N_5425,N_4776,N_4981);
or U5426 (N_5426,N_4636,N_4723);
xor U5427 (N_5427,N_4981,N_4785);
or U5428 (N_5428,N_4603,N_4699);
nor U5429 (N_5429,N_4906,N_4867);
and U5430 (N_5430,N_4931,N_4872);
nand U5431 (N_5431,N_4752,N_4885);
or U5432 (N_5432,N_4606,N_4876);
nor U5433 (N_5433,N_4964,N_4801);
or U5434 (N_5434,N_4671,N_4862);
nand U5435 (N_5435,N_4516,N_4925);
xor U5436 (N_5436,N_4940,N_4658);
or U5437 (N_5437,N_4634,N_4943);
and U5438 (N_5438,N_4918,N_4667);
nand U5439 (N_5439,N_4856,N_4564);
or U5440 (N_5440,N_4699,N_4903);
or U5441 (N_5441,N_4700,N_4726);
xnor U5442 (N_5442,N_4891,N_4785);
nand U5443 (N_5443,N_4861,N_4694);
nand U5444 (N_5444,N_4800,N_4775);
or U5445 (N_5445,N_4639,N_4860);
xnor U5446 (N_5446,N_4999,N_4566);
and U5447 (N_5447,N_4517,N_4804);
and U5448 (N_5448,N_4900,N_4853);
or U5449 (N_5449,N_4625,N_4894);
nor U5450 (N_5450,N_4580,N_4954);
and U5451 (N_5451,N_4656,N_4609);
or U5452 (N_5452,N_4647,N_4887);
xor U5453 (N_5453,N_4601,N_4917);
nand U5454 (N_5454,N_4840,N_4951);
and U5455 (N_5455,N_4984,N_4594);
or U5456 (N_5456,N_4892,N_4968);
nor U5457 (N_5457,N_4798,N_4910);
nor U5458 (N_5458,N_4990,N_4693);
or U5459 (N_5459,N_4817,N_4524);
nor U5460 (N_5460,N_4644,N_4811);
and U5461 (N_5461,N_4517,N_4746);
and U5462 (N_5462,N_4814,N_4533);
or U5463 (N_5463,N_4945,N_4815);
and U5464 (N_5464,N_4926,N_4839);
or U5465 (N_5465,N_4853,N_4660);
nor U5466 (N_5466,N_4942,N_4997);
xor U5467 (N_5467,N_4774,N_4941);
and U5468 (N_5468,N_4572,N_4917);
nor U5469 (N_5469,N_4811,N_4506);
nor U5470 (N_5470,N_4583,N_4711);
xor U5471 (N_5471,N_4848,N_4635);
and U5472 (N_5472,N_4559,N_4607);
or U5473 (N_5473,N_4508,N_4658);
nand U5474 (N_5474,N_4921,N_4719);
nor U5475 (N_5475,N_4884,N_4811);
nand U5476 (N_5476,N_4724,N_4606);
and U5477 (N_5477,N_4625,N_4868);
xnor U5478 (N_5478,N_4799,N_4572);
and U5479 (N_5479,N_4794,N_4517);
nor U5480 (N_5480,N_4651,N_4836);
and U5481 (N_5481,N_4517,N_4757);
or U5482 (N_5482,N_4565,N_4785);
nand U5483 (N_5483,N_4981,N_4914);
or U5484 (N_5484,N_4645,N_4681);
nand U5485 (N_5485,N_4721,N_4645);
or U5486 (N_5486,N_4858,N_4960);
xnor U5487 (N_5487,N_4785,N_4743);
and U5488 (N_5488,N_4515,N_4990);
nand U5489 (N_5489,N_4763,N_4989);
xnor U5490 (N_5490,N_4657,N_4799);
or U5491 (N_5491,N_4550,N_4662);
or U5492 (N_5492,N_4777,N_4529);
xnor U5493 (N_5493,N_4611,N_4777);
and U5494 (N_5494,N_4868,N_4988);
or U5495 (N_5495,N_4628,N_4635);
or U5496 (N_5496,N_4608,N_4657);
or U5497 (N_5497,N_4749,N_4678);
nor U5498 (N_5498,N_4794,N_4589);
nand U5499 (N_5499,N_4618,N_4612);
nand U5500 (N_5500,N_5220,N_5376);
nand U5501 (N_5501,N_5452,N_5051);
nand U5502 (N_5502,N_5102,N_5407);
and U5503 (N_5503,N_5019,N_5396);
and U5504 (N_5504,N_5058,N_5101);
or U5505 (N_5505,N_5193,N_5275);
nand U5506 (N_5506,N_5115,N_5195);
nand U5507 (N_5507,N_5207,N_5171);
and U5508 (N_5508,N_5088,N_5347);
nand U5509 (N_5509,N_5394,N_5231);
and U5510 (N_5510,N_5449,N_5397);
and U5511 (N_5511,N_5338,N_5271);
nor U5512 (N_5512,N_5285,N_5146);
or U5513 (N_5513,N_5063,N_5162);
nor U5514 (N_5514,N_5110,N_5380);
or U5515 (N_5515,N_5147,N_5428);
and U5516 (N_5516,N_5348,N_5400);
xor U5517 (N_5517,N_5015,N_5364);
nor U5518 (N_5518,N_5450,N_5175);
xor U5519 (N_5519,N_5234,N_5490);
xor U5520 (N_5520,N_5496,N_5018);
nor U5521 (N_5521,N_5368,N_5025);
and U5522 (N_5522,N_5432,N_5411);
nand U5523 (N_5523,N_5337,N_5096);
xnor U5524 (N_5524,N_5196,N_5289);
nand U5525 (N_5525,N_5427,N_5090);
or U5526 (N_5526,N_5247,N_5483);
xnor U5527 (N_5527,N_5322,N_5164);
nor U5528 (N_5528,N_5371,N_5216);
nor U5529 (N_5529,N_5303,N_5445);
nor U5530 (N_5530,N_5441,N_5374);
nand U5531 (N_5531,N_5122,N_5140);
and U5532 (N_5532,N_5143,N_5073);
nor U5533 (N_5533,N_5237,N_5230);
nor U5534 (N_5534,N_5050,N_5240);
nor U5535 (N_5535,N_5480,N_5125);
or U5536 (N_5536,N_5165,N_5153);
nor U5537 (N_5537,N_5443,N_5304);
nor U5538 (N_5538,N_5270,N_5087);
xnor U5539 (N_5539,N_5023,N_5226);
or U5540 (N_5540,N_5020,N_5393);
nand U5541 (N_5541,N_5349,N_5273);
and U5542 (N_5542,N_5229,N_5280);
nor U5543 (N_5543,N_5069,N_5199);
xnor U5544 (N_5544,N_5384,N_5189);
or U5545 (N_5545,N_5053,N_5156);
or U5546 (N_5546,N_5013,N_5442);
or U5547 (N_5547,N_5404,N_5318);
or U5548 (N_5548,N_5116,N_5118);
xnor U5549 (N_5549,N_5106,N_5042);
nor U5550 (N_5550,N_5222,N_5287);
xnor U5551 (N_5551,N_5067,N_5484);
and U5552 (N_5552,N_5072,N_5361);
and U5553 (N_5553,N_5281,N_5401);
or U5554 (N_5554,N_5470,N_5472);
nor U5555 (N_5555,N_5149,N_5469);
nor U5556 (N_5556,N_5346,N_5468);
nand U5557 (N_5557,N_5012,N_5011);
or U5558 (N_5558,N_5100,N_5037);
xor U5559 (N_5559,N_5253,N_5258);
nor U5560 (N_5560,N_5099,N_5487);
and U5561 (N_5561,N_5276,N_5036);
xor U5562 (N_5562,N_5232,N_5137);
and U5563 (N_5563,N_5084,N_5028);
xnor U5564 (N_5564,N_5353,N_5499);
and U5565 (N_5565,N_5486,N_5462);
nor U5566 (N_5566,N_5208,N_5184);
nor U5567 (N_5567,N_5246,N_5182);
and U5568 (N_5568,N_5279,N_5370);
nor U5569 (N_5569,N_5154,N_5402);
nor U5570 (N_5570,N_5435,N_5382);
xor U5571 (N_5571,N_5215,N_5465);
and U5572 (N_5572,N_5075,N_5167);
or U5573 (N_5573,N_5004,N_5282);
xor U5574 (N_5574,N_5398,N_5214);
nor U5575 (N_5575,N_5498,N_5440);
or U5576 (N_5576,N_5326,N_5181);
nor U5577 (N_5577,N_5225,N_5277);
nand U5578 (N_5578,N_5212,N_5413);
xnor U5579 (N_5579,N_5485,N_5148);
or U5580 (N_5580,N_5309,N_5111);
nor U5581 (N_5581,N_5330,N_5333);
xor U5582 (N_5582,N_5160,N_5244);
or U5583 (N_5583,N_5478,N_5113);
xor U5584 (N_5584,N_5493,N_5410);
or U5585 (N_5585,N_5306,N_5366);
xor U5586 (N_5586,N_5161,N_5310);
nor U5587 (N_5587,N_5217,N_5286);
xnor U5588 (N_5588,N_5000,N_5201);
nor U5589 (N_5589,N_5121,N_5467);
and U5590 (N_5590,N_5060,N_5294);
and U5591 (N_5591,N_5205,N_5259);
nand U5592 (N_5592,N_5006,N_5040);
xnor U5593 (N_5593,N_5495,N_5352);
or U5594 (N_5594,N_5123,N_5224);
or U5595 (N_5595,N_5068,N_5412);
xor U5596 (N_5596,N_5250,N_5491);
nand U5597 (N_5597,N_5488,N_5359);
or U5598 (N_5598,N_5190,N_5301);
and U5599 (N_5599,N_5362,N_5200);
and U5600 (N_5600,N_5218,N_5245);
xnor U5601 (N_5601,N_5424,N_5097);
xnor U5602 (N_5602,N_5455,N_5134);
or U5603 (N_5603,N_5296,N_5071);
and U5604 (N_5604,N_5431,N_5320);
xor U5605 (N_5605,N_5249,N_5031);
nand U5606 (N_5606,N_5492,N_5355);
or U5607 (N_5607,N_5264,N_5083);
xnor U5608 (N_5608,N_5086,N_5065);
xnor U5609 (N_5609,N_5295,N_5336);
nand U5610 (N_5610,N_5016,N_5302);
nor U5611 (N_5611,N_5372,N_5290);
or U5612 (N_5612,N_5183,N_5079);
nor U5613 (N_5613,N_5390,N_5010);
nand U5614 (N_5614,N_5461,N_5415);
nor U5615 (N_5615,N_5152,N_5210);
and U5616 (N_5616,N_5057,N_5267);
or U5617 (N_5617,N_5409,N_5062);
xnor U5618 (N_5618,N_5239,N_5344);
nor U5619 (N_5619,N_5104,N_5003);
xnor U5620 (N_5620,N_5185,N_5339);
xor U5621 (N_5621,N_5414,N_5095);
nor U5622 (N_5622,N_5298,N_5064);
or U5623 (N_5623,N_5399,N_5489);
and U5624 (N_5624,N_5300,N_5261);
and U5625 (N_5625,N_5345,N_5022);
nand U5626 (N_5626,N_5177,N_5438);
xnor U5627 (N_5627,N_5299,N_5001);
and U5628 (N_5628,N_5466,N_5494);
and U5629 (N_5629,N_5363,N_5408);
xnor U5630 (N_5630,N_5248,N_5151);
nand U5631 (N_5631,N_5365,N_5029);
xnor U5632 (N_5632,N_5383,N_5213);
nor U5633 (N_5633,N_5454,N_5074);
xor U5634 (N_5634,N_5308,N_5117);
and U5635 (N_5635,N_5108,N_5091);
xor U5636 (N_5636,N_5098,N_5227);
xor U5637 (N_5637,N_5360,N_5136);
nor U5638 (N_5638,N_5233,N_5460);
nor U5639 (N_5639,N_5076,N_5288);
nand U5640 (N_5640,N_5420,N_5129);
nand U5641 (N_5641,N_5202,N_5292);
nor U5642 (N_5642,N_5186,N_5257);
nand U5643 (N_5643,N_5173,N_5479);
xnor U5644 (N_5644,N_5124,N_5406);
nor U5645 (N_5645,N_5446,N_5350);
nor U5646 (N_5646,N_5158,N_5203);
nor U5647 (N_5647,N_5238,N_5343);
or U5648 (N_5648,N_5451,N_5439);
nand U5649 (N_5649,N_5197,N_5473);
nand U5650 (N_5650,N_5033,N_5430);
nand U5651 (N_5651,N_5314,N_5317);
xnor U5652 (N_5652,N_5166,N_5260);
nor U5653 (N_5653,N_5005,N_5312);
or U5654 (N_5654,N_5319,N_5114);
or U5655 (N_5655,N_5180,N_5142);
or U5656 (N_5656,N_5170,N_5092);
and U5657 (N_5657,N_5313,N_5265);
nor U5658 (N_5658,N_5085,N_5423);
nand U5659 (N_5659,N_5219,N_5323);
nor U5660 (N_5660,N_5047,N_5437);
or U5661 (N_5661,N_5388,N_5112);
nand U5662 (N_5662,N_5444,N_5082);
and U5663 (N_5663,N_5351,N_5132);
xor U5664 (N_5664,N_5476,N_5387);
nand U5665 (N_5665,N_5297,N_5262);
nor U5666 (N_5666,N_5155,N_5236);
nand U5667 (N_5667,N_5059,N_5070);
nand U5668 (N_5668,N_5327,N_5335);
and U5669 (N_5669,N_5332,N_5284);
and U5670 (N_5670,N_5429,N_5135);
nor U5671 (N_5671,N_5139,N_5127);
nand U5672 (N_5672,N_5128,N_5223);
nor U5673 (N_5673,N_5375,N_5176);
or U5674 (N_5674,N_5268,N_5103);
nand U5675 (N_5675,N_5456,N_5340);
and U5676 (N_5676,N_5316,N_5341);
nand U5677 (N_5677,N_5477,N_5405);
nand U5678 (N_5678,N_5055,N_5174);
nand U5679 (N_5679,N_5369,N_5130);
nor U5680 (N_5680,N_5272,N_5089);
or U5681 (N_5681,N_5459,N_5081);
nand U5682 (N_5682,N_5315,N_5043);
nor U5683 (N_5683,N_5367,N_5169);
nand U5684 (N_5684,N_5354,N_5178);
and U5685 (N_5685,N_5386,N_5241);
xor U5686 (N_5686,N_5024,N_5044);
nand U5687 (N_5687,N_5187,N_5093);
and U5688 (N_5688,N_5311,N_5263);
nor U5689 (N_5689,N_5356,N_5426);
and U5690 (N_5690,N_5436,N_5391);
nor U5691 (N_5691,N_5358,N_5243);
nand U5692 (N_5692,N_5325,N_5209);
xnor U5693 (N_5693,N_5221,N_5283);
and U5694 (N_5694,N_5039,N_5418);
nand U5695 (N_5695,N_5256,N_5206);
and U5696 (N_5696,N_5389,N_5434);
or U5697 (N_5697,N_5497,N_5052);
or U5698 (N_5698,N_5464,N_5471);
nor U5699 (N_5699,N_5119,N_5048);
and U5700 (N_5700,N_5274,N_5379);
nand U5701 (N_5701,N_5251,N_5373);
and U5702 (N_5702,N_5255,N_5453);
nor U5703 (N_5703,N_5254,N_5378);
nor U5704 (N_5704,N_5080,N_5021);
and U5705 (N_5705,N_5192,N_5045);
nor U5706 (N_5706,N_5194,N_5094);
and U5707 (N_5707,N_5107,N_5009);
nor U5708 (N_5708,N_5321,N_5377);
nor U5709 (N_5709,N_5381,N_5026);
nand U5710 (N_5710,N_5120,N_5144);
and U5711 (N_5711,N_5046,N_5228);
and U5712 (N_5712,N_5007,N_5481);
or U5713 (N_5713,N_5331,N_5014);
nand U5714 (N_5714,N_5357,N_5416);
nor U5715 (N_5715,N_5054,N_5448);
and U5716 (N_5716,N_5403,N_5385);
xor U5717 (N_5717,N_5126,N_5041);
or U5718 (N_5718,N_5457,N_5235);
xnor U5719 (N_5719,N_5422,N_5002);
nor U5720 (N_5720,N_5293,N_5334);
nor U5721 (N_5721,N_5269,N_5038);
and U5722 (N_5722,N_5305,N_5474);
nand U5723 (N_5723,N_5105,N_5419);
nor U5724 (N_5724,N_5395,N_5168);
and U5725 (N_5725,N_5032,N_5463);
or U5726 (N_5726,N_5417,N_5066);
nor U5727 (N_5727,N_5035,N_5475);
or U5728 (N_5728,N_5278,N_5133);
nand U5729 (N_5729,N_5425,N_5077);
nand U5730 (N_5730,N_5008,N_5138);
nor U5731 (N_5731,N_5266,N_5163);
xnor U5732 (N_5732,N_5027,N_5307);
xnor U5733 (N_5733,N_5179,N_5482);
and U5734 (N_5734,N_5458,N_5291);
nand U5735 (N_5735,N_5141,N_5242);
xnor U5736 (N_5736,N_5328,N_5150);
nor U5737 (N_5737,N_5198,N_5324);
nor U5738 (N_5738,N_5211,N_5433);
xor U5739 (N_5739,N_5030,N_5017);
nand U5740 (N_5740,N_5034,N_5061);
nor U5741 (N_5741,N_5392,N_5188);
or U5742 (N_5742,N_5109,N_5252);
nor U5743 (N_5743,N_5172,N_5329);
or U5744 (N_5744,N_5421,N_5145);
and U5745 (N_5745,N_5447,N_5191);
and U5746 (N_5746,N_5078,N_5056);
and U5747 (N_5747,N_5049,N_5131);
or U5748 (N_5748,N_5157,N_5342);
nor U5749 (N_5749,N_5159,N_5204);
and U5750 (N_5750,N_5032,N_5438);
xor U5751 (N_5751,N_5369,N_5450);
xor U5752 (N_5752,N_5239,N_5110);
xnor U5753 (N_5753,N_5441,N_5194);
nor U5754 (N_5754,N_5476,N_5479);
xor U5755 (N_5755,N_5188,N_5307);
and U5756 (N_5756,N_5259,N_5098);
nand U5757 (N_5757,N_5348,N_5253);
xor U5758 (N_5758,N_5497,N_5430);
nor U5759 (N_5759,N_5472,N_5056);
nand U5760 (N_5760,N_5402,N_5462);
nor U5761 (N_5761,N_5180,N_5017);
or U5762 (N_5762,N_5478,N_5011);
and U5763 (N_5763,N_5430,N_5409);
and U5764 (N_5764,N_5435,N_5437);
and U5765 (N_5765,N_5426,N_5307);
nand U5766 (N_5766,N_5356,N_5407);
xor U5767 (N_5767,N_5202,N_5276);
nor U5768 (N_5768,N_5182,N_5317);
xor U5769 (N_5769,N_5403,N_5490);
and U5770 (N_5770,N_5089,N_5038);
and U5771 (N_5771,N_5196,N_5477);
nor U5772 (N_5772,N_5209,N_5135);
nand U5773 (N_5773,N_5211,N_5127);
nor U5774 (N_5774,N_5210,N_5260);
nand U5775 (N_5775,N_5131,N_5355);
xor U5776 (N_5776,N_5132,N_5251);
xnor U5777 (N_5777,N_5289,N_5432);
or U5778 (N_5778,N_5172,N_5043);
and U5779 (N_5779,N_5144,N_5301);
or U5780 (N_5780,N_5304,N_5362);
or U5781 (N_5781,N_5475,N_5179);
xor U5782 (N_5782,N_5446,N_5018);
xor U5783 (N_5783,N_5393,N_5358);
and U5784 (N_5784,N_5131,N_5000);
or U5785 (N_5785,N_5350,N_5433);
nor U5786 (N_5786,N_5474,N_5092);
or U5787 (N_5787,N_5294,N_5284);
and U5788 (N_5788,N_5144,N_5136);
xnor U5789 (N_5789,N_5080,N_5005);
xor U5790 (N_5790,N_5088,N_5459);
nor U5791 (N_5791,N_5171,N_5038);
or U5792 (N_5792,N_5098,N_5189);
and U5793 (N_5793,N_5144,N_5247);
or U5794 (N_5794,N_5112,N_5305);
nor U5795 (N_5795,N_5175,N_5014);
nor U5796 (N_5796,N_5404,N_5481);
and U5797 (N_5797,N_5384,N_5424);
and U5798 (N_5798,N_5499,N_5323);
xnor U5799 (N_5799,N_5319,N_5469);
xnor U5800 (N_5800,N_5484,N_5109);
and U5801 (N_5801,N_5324,N_5466);
or U5802 (N_5802,N_5054,N_5414);
nand U5803 (N_5803,N_5460,N_5353);
nand U5804 (N_5804,N_5168,N_5080);
or U5805 (N_5805,N_5389,N_5008);
xnor U5806 (N_5806,N_5063,N_5145);
nor U5807 (N_5807,N_5336,N_5226);
nand U5808 (N_5808,N_5398,N_5466);
nor U5809 (N_5809,N_5307,N_5263);
nand U5810 (N_5810,N_5398,N_5308);
nand U5811 (N_5811,N_5039,N_5316);
and U5812 (N_5812,N_5446,N_5335);
nand U5813 (N_5813,N_5415,N_5111);
nand U5814 (N_5814,N_5342,N_5427);
xnor U5815 (N_5815,N_5448,N_5161);
and U5816 (N_5816,N_5092,N_5383);
or U5817 (N_5817,N_5224,N_5276);
nor U5818 (N_5818,N_5499,N_5015);
nand U5819 (N_5819,N_5112,N_5308);
nor U5820 (N_5820,N_5415,N_5440);
nand U5821 (N_5821,N_5322,N_5058);
nand U5822 (N_5822,N_5063,N_5065);
xnor U5823 (N_5823,N_5016,N_5006);
or U5824 (N_5824,N_5349,N_5314);
nor U5825 (N_5825,N_5472,N_5337);
xnor U5826 (N_5826,N_5077,N_5267);
xor U5827 (N_5827,N_5366,N_5129);
nand U5828 (N_5828,N_5418,N_5077);
or U5829 (N_5829,N_5219,N_5252);
xor U5830 (N_5830,N_5156,N_5077);
xor U5831 (N_5831,N_5127,N_5192);
nand U5832 (N_5832,N_5316,N_5086);
and U5833 (N_5833,N_5425,N_5254);
or U5834 (N_5834,N_5423,N_5259);
nand U5835 (N_5835,N_5100,N_5301);
or U5836 (N_5836,N_5136,N_5449);
xnor U5837 (N_5837,N_5200,N_5305);
nand U5838 (N_5838,N_5117,N_5068);
and U5839 (N_5839,N_5228,N_5156);
and U5840 (N_5840,N_5275,N_5209);
nor U5841 (N_5841,N_5092,N_5070);
and U5842 (N_5842,N_5097,N_5111);
and U5843 (N_5843,N_5145,N_5111);
nor U5844 (N_5844,N_5380,N_5233);
or U5845 (N_5845,N_5392,N_5069);
and U5846 (N_5846,N_5449,N_5264);
and U5847 (N_5847,N_5312,N_5300);
or U5848 (N_5848,N_5401,N_5191);
xnor U5849 (N_5849,N_5328,N_5032);
or U5850 (N_5850,N_5044,N_5058);
and U5851 (N_5851,N_5458,N_5408);
nor U5852 (N_5852,N_5207,N_5235);
or U5853 (N_5853,N_5049,N_5194);
and U5854 (N_5854,N_5223,N_5209);
xor U5855 (N_5855,N_5468,N_5259);
and U5856 (N_5856,N_5240,N_5336);
or U5857 (N_5857,N_5295,N_5286);
xor U5858 (N_5858,N_5420,N_5272);
or U5859 (N_5859,N_5272,N_5207);
xnor U5860 (N_5860,N_5156,N_5495);
xor U5861 (N_5861,N_5106,N_5213);
nand U5862 (N_5862,N_5140,N_5358);
nor U5863 (N_5863,N_5463,N_5325);
nor U5864 (N_5864,N_5309,N_5304);
xor U5865 (N_5865,N_5471,N_5449);
nand U5866 (N_5866,N_5328,N_5492);
or U5867 (N_5867,N_5418,N_5215);
nand U5868 (N_5868,N_5095,N_5396);
nor U5869 (N_5869,N_5350,N_5246);
xnor U5870 (N_5870,N_5272,N_5376);
nor U5871 (N_5871,N_5405,N_5146);
xor U5872 (N_5872,N_5452,N_5036);
or U5873 (N_5873,N_5254,N_5407);
nor U5874 (N_5874,N_5496,N_5246);
xnor U5875 (N_5875,N_5333,N_5430);
nand U5876 (N_5876,N_5034,N_5317);
and U5877 (N_5877,N_5337,N_5095);
nor U5878 (N_5878,N_5041,N_5193);
and U5879 (N_5879,N_5096,N_5293);
nand U5880 (N_5880,N_5260,N_5071);
nand U5881 (N_5881,N_5186,N_5413);
xnor U5882 (N_5882,N_5443,N_5047);
nor U5883 (N_5883,N_5065,N_5209);
xor U5884 (N_5884,N_5271,N_5430);
or U5885 (N_5885,N_5263,N_5237);
xnor U5886 (N_5886,N_5359,N_5142);
xor U5887 (N_5887,N_5280,N_5117);
and U5888 (N_5888,N_5149,N_5311);
or U5889 (N_5889,N_5242,N_5409);
xnor U5890 (N_5890,N_5201,N_5047);
or U5891 (N_5891,N_5304,N_5122);
nand U5892 (N_5892,N_5204,N_5126);
and U5893 (N_5893,N_5357,N_5031);
and U5894 (N_5894,N_5121,N_5452);
nor U5895 (N_5895,N_5195,N_5160);
nand U5896 (N_5896,N_5446,N_5247);
xor U5897 (N_5897,N_5349,N_5194);
nor U5898 (N_5898,N_5162,N_5215);
or U5899 (N_5899,N_5250,N_5123);
and U5900 (N_5900,N_5464,N_5327);
or U5901 (N_5901,N_5467,N_5457);
or U5902 (N_5902,N_5261,N_5057);
nand U5903 (N_5903,N_5161,N_5023);
nand U5904 (N_5904,N_5411,N_5438);
or U5905 (N_5905,N_5195,N_5450);
nand U5906 (N_5906,N_5347,N_5206);
nand U5907 (N_5907,N_5382,N_5447);
and U5908 (N_5908,N_5118,N_5463);
or U5909 (N_5909,N_5176,N_5260);
xnor U5910 (N_5910,N_5493,N_5305);
xor U5911 (N_5911,N_5333,N_5382);
and U5912 (N_5912,N_5354,N_5068);
and U5913 (N_5913,N_5390,N_5444);
and U5914 (N_5914,N_5127,N_5370);
xnor U5915 (N_5915,N_5188,N_5295);
nand U5916 (N_5916,N_5206,N_5434);
and U5917 (N_5917,N_5140,N_5189);
xnor U5918 (N_5918,N_5497,N_5248);
or U5919 (N_5919,N_5403,N_5226);
or U5920 (N_5920,N_5272,N_5357);
and U5921 (N_5921,N_5081,N_5038);
xnor U5922 (N_5922,N_5427,N_5297);
xor U5923 (N_5923,N_5004,N_5189);
or U5924 (N_5924,N_5341,N_5260);
xnor U5925 (N_5925,N_5018,N_5443);
nand U5926 (N_5926,N_5494,N_5370);
xor U5927 (N_5927,N_5083,N_5027);
nor U5928 (N_5928,N_5266,N_5221);
xor U5929 (N_5929,N_5151,N_5240);
and U5930 (N_5930,N_5232,N_5283);
nand U5931 (N_5931,N_5090,N_5126);
nand U5932 (N_5932,N_5174,N_5475);
nor U5933 (N_5933,N_5013,N_5010);
nand U5934 (N_5934,N_5402,N_5388);
nor U5935 (N_5935,N_5189,N_5151);
and U5936 (N_5936,N_5450,N_5321);
and U5937 (N_5937,N_5030,N_5432);
or U5938 (N_5938,N_5214,N_5209);
nor U5939 (N_5939,N_5404,N_5115);
nor U5940 (N_5940,N_5285,N_5036);
nand U5941 (N_5941,N_5129,N_5163);
nor U5942 (N_5942,N_5081,N_5263);
and U5943 (N_5943,N_5293,N_5241);
xnor U5944 (N_5944,N_5453,N_5339);
nor U5945 (N_5945,N_5096,N_5239);
nand U5946 (N_5946,N_5046,N_5187);
nor U5947 (N_5947,N_5177,N_5020);
nor U5948 (N_5948,N_5452,N_5302);
or U5949 (N_5949,N_5431,N_5382);
and U5950 (N_5950,N_5007,N_5009);
nor U5951 (N_5951,N_5116,N_5495);
nand U5952 (N_5952,N_5230,N_5280);
nor U5953 (N_5953,N_5310,N_5043);
and U5954 (N_5954,N_5257,N_5465);
xnor U5955 (N_5955,N_5069,N_5093);
or U5956 (N_5956,N_5289,N_5409);
nor U5957 (N_5957,N_5203,N_5038);
and U5958 (N_5958,N_5490,N_5023);
or U5959 (N_5959,N_5254,N_5326);
xor U5960 (N_5960,N_5150,N_5261);
and U5961 (N_5961,N_5129,N_5067);
xor U5962 (N_5962,N_5252,N_5212);
nand U5963 (N_5963,N_5430,N_5015);
or U5964 (N_5964,N_5307,N_5479);
and U5965 (N_5965,N_5039,N_5237);
or U5966 (N_5966,N_5164,N_5199);
and U5967 (N_5967,N_5004,N_5109);
and U5968 (N_5968,N_5375,N_5155);
and U5969 (N_5969,N_5455,N_5200);
nand U5970 (N_5970,N_5242,N_5044);
and U5971 (N_5971,N_5136,N_5422);
or U5972 (N_5972,N_5167,N_5053);
xor U5973 (N_5973,N_5321,N_5368);
and U5974 (N_5974,N_5171,N_5358);
nand U5975 (N_5975,N_5031,N_5047);
and U5976 (N_5976,N_5413,N_5297);
or U5977 (N_5977,N_5137,N_5376);
nor U5978 (N_5978,N_5061,N_5214);
xnor U5979 (N_5979,N_5094,N_5492);
xor U5980 (N_5980,N_5127,N_5368);
nand U5981 (N_5981,N_5439,N_5358);
nor U5982 (N_5982,N_5096,N_5278);
nand U5983 (N_5983,N_5202,N_5141);
nand U5984 (N_5984,N_5102,N_5018);
and U5985 (N_5985,N_5280,N_5078);
nand U5986 (N_5986,N_5103,N_5469);
and U5987 (N_5987,N_5175,N_5253);
xnor U5988 (N_5988,N_5028,N_5049);
or U5989 (N_5989,N_5041,N_5322);
nand U5990 (N_5990,N_5061,N_5158);
xnor U5991 (N_5991,N_5160,N_5148);
xor U5992 (N_5992,N_5012,N_5056);
xor U5993 (N_5993,N_5365,N_5241);
nand U5994 (N_5994,N_5467,N_5472);
or U5995 (N_5995,N_5176,N_5383);
xnor U5996 (N_5996,N_5296,N_5141);
or U5997 (N_5997,N_5343,N_5419);
xnor U5998 (N_5998,N_5373,N_5479);
nand U5999 (N_5999,N_5145,N_5206);
xor U6000 (N_6000,N_5564,N_5893);
xor U6001 (N_6001,N_5825,N_5658);
xor U6002 (N_6002,N_5911,N_5934);
nand U6003 (N_6003,N_5515,N_5928);
and U6004 (N_6004,N_5545,N_5558);
and U6005 (N_6005,N_5628,N_5806);
xor U6006 (N_6006,N_5646,N_5524);
nor U6007 (N_6007,N_5981,N_5886);
nor U6008 (N_6008,N_5565,N_5706);
and U6009 (N_6009,N_5547,N_5789);
or U6010 (N_6010,N_5796,N_5895);
nor U6011 (N_6011,N_5742,N_5923);
or U6012 (N_6012,N_5899,N_5753);
nor U6013 (N_6013,N_5920,N_5766);
xnor U6014 (N_6014,N_5717,N_5639);
nand U6015 (N_6015,N_5657,N_5559);
and U6016 (N_6016,N_5687,N_5567);
xnor U6017 (N_6017,N_5666,N_5574);
and U6018 (N_6018,N_5816,N_5964);
and U6019 (N_6019,N_5521,N_5793);
or U6020 (N_6020,N_5865,N_5955);
or U6021 (N_6021,N_5780,N_5739);
or U6022 (N_6022,N_5936,N_5840);
nor U6023 (N_6023,N_5686,N_5677);
xor U6024 (N_6024,N_5670,N_5653);
or U6025 (N_6025,N_5831,N_5710);
xnor U6026 (N_6026,N_5975,N_5808);
and U6027 (N_6027,N_5872,N_5999);
and U6028 (N_6028,N_5509,N_5751);
or U6029 (N_6029,N_5650,N_5620);
nor U6030 (N_6030,N_5728,N_5544);
and U6031 (N_6031,N_5866,N_5944);
nand U6032 (N_6032,N_5605,N_5651);
and U6033 (N_6033,N_5730,N_5659);
nor U6034 (N_6034,N_5966,N_5504);
and U6035 (N_6035,N_5933,N_5756);
nand U6036 (N_6036,N_5578,N_5554);
xnor U6037 (N_6037,N_5665,N_5634);
nand U6038 (N_6038,N_5917,N_5705);
and U6039 (N_6039,N_5845,N_5542);
nor U6040 (N_6040,N_5852,N_5674);
and U6041 (N_6041,N_5778,N_5617);
xnor U6042 (N_6042,N_5838,N_5681);
nor U6043 (N_6043,N_5848,N_5703);
or U6044 (N_6044,N_5506,N_5969);
or U6045 (N_6045,N_5712,N_5675);
nor U6046 (N_6046,N_5827,N_5697);
nor U6047 (N_6047,N_5773,N_5948);
or U6048 (N_6048,N_5992,N_5925);
or U6049 (N_6049,N_5669,N_5957);
xor U6050 (N_6050,N_5580,N_5711);
and U6051 (N_6051,N_5997,N_5685);
nand U6052 (N_6052,N_5864,N_5759);
xnor U6053 (N_6053,N_5531,N_5926);
nor U6054 (N_6054,N_5914,N_5757);
and U6055 (N_6055,N_5995,N_5523);
xnor U6056 (N_6056,N_5549,N_5783);
and U6057 (N_6057,N_5704,N_5630);
and U6058 (N_6058,N_5671,N_5570);
nand U6059 (N_6059,N_5566,N_5998);
or U6060 (N_6060,N_5528,N_5551);
nand U6061 (N_6061,N_5777,N_5880);
and U6062 (N_6062,N_5735,N_5738);
xor U6063 (N_6063,N_5889,N_5861);
and U6064 (N_6064,N_5961,N_5633);
and U6065 (N_6065,N_5573,N_5682);
nor U6066 (N_6066,N_5737,N_5505);
nor U6067 (N_6067,N_5618,N_5799);
xor U6068 (N_6068,N_5863,N_5968);
nor U6069 (N_6069,N_5820,N_5534);
xor U6070 (N_6070,N_5600,N_5815);
xnor U6071 (N_6071,N_5514,N_5599);
nor U6072 (N_6072,N_5813,N_5832);
nor U6073 (N_6073,N_5589,N_5718);
or U6074 (N_6074,N_5994,N_5904);
nand U6075 (N_6075,N_5945,N_5621);
or U6076 (N_6076,N_5696,N_5731);
or U6077 (N_6077,N_5942,N_5977);
nor U6078 (N_6078,N_5823,N_5941);
xnor U6079 (N_6079,N_5930,N_5905);
and U6080 (N_6080,N_5846,N_5588);
nand U6081 (N_6081,N_5550,N_5656);
nor U6082 (N_6082,N_5841,N_5919);
xnor U6083 (N_6083,N_5980,N_5859);
and U6084 (N_6084,N_5702,N_5987);
or U6085 (N_6085,N_5835,N_5803);
xor U6086 (N_6086,N_5877,N_5894);
xnor U6087 (N_6087,N_5597,N_5976);
or U6088 (N_6088,N_5684,N_5918);
and U6089 (N_6089,N_5819,N_5720);
and U6090 (N_6090,N_5912,N_5698);
nor U6091 (N_6091,N_5722,N_5826);
nor U6092 (N_6092,N_5887,N_5715);
xnor U6093 (N_6093,N_5527,N_5518);
or U6094 (N_6094,N_5770,N_5609);
xnor U6095 (N_6095,N_5922,N_5908);
or U6096 (N_6096,N_5790,N_5641);
xnor U6097 (N_6097,N_5931,N_5736);
nand U6098 (N_6098,N_5842,N_5851);
nor U6099 (N_6099,N_5507,N_5985);
nor U6100 (N_6100,N_5700,N_5781);
nor U6101 (N_6101,N_5878,N_5741);
or U6102 (N_6102,N_5667,N_5583);
nand U6103 (N_6103,N_5631,N_5619);
nand U6104 (N_6104,N_5533,N_5868);
nand U6105 (N_6105,N_5869,N_5626);
xnor U6106 (N_6106,N_5636,N_5805);
and U6107 (N_6107,N_5910,N_5690);
or U6108 (N_6108,N_5602,N_5592);
nor U6109 (N_6109,N_5986,N_5654);
nor U6110 (N_6110,N_5956,N_5937);
or U6111 (N_6111,N_5817,N_5638);
xor U6112 (N_6112,N_5530,N_5959);
xor U6113 (N_6113,N_5673,N_5557);
and U6114 (N_6114,N_5661,N_5511);
and U6115 (N_6115,N_5951,N_5939);
nand U6116 (N_6116,N_5679,N_5774);
nor U6117 (N_6117,N_5579,N_5884);
nor U6118 (N_6118,N_5595,N_5516);
nor U6119 (N_6119,N_5900,N_5973);
xnor U6120 (N_6120,N_5811,N_5744);
nor U6121 (N_6121,N_5556,N_5940);
nand U6122 (N_6122,N_5629,N_5586);
nand U6123 (N_6123,N_5584,N_5585);
or U6124 (N_6124,N_5726,N_5541);
nor U6125 (N_6125,N_5536,N_5879);
nor U6126 (N_6126,N_5555,N_5818);
and U6127 (N_6127,N_5635,N_5890);
xor U6128 (N_6128,N_5582,N_5867);
nand U6129 (N_6129,N_5915,N_5517);
nor U6130 (N_6130,N_5611,N_5576);
xor U6131 (N_6131,N_5642,N_5873);
nand U6132 (N_6132,N_5571,N_5947);
nand U6133 (N_6133,N_5984,N_5699);
xnor U6134 (N_6134,N_5891,N_5608);
or U6135 (N_6135,N_5779,N_5577);
nand U6136 (N_6136,N_5860,N_5768);
nand U6137 (N_6137,N_5938,N_5694);
xor U6138 (N_6138,N_5752,N_5708);
nand U6139 (N_6139,N_5809,N_5593);
and U6140 (N_6140,N_5668,N_5971);
nor U6141 (N_6141,N_5624,N_5786);
or U6142 (N_6142,N_5807,N_5672);
or U6143 (N_6143,N_5615,N_5834);
or U6144 (N_6144,N_5965,N_5622);
nand U6145 (N_6145,N_5643,N_5647);
nor U6146 (N_6146,N_5746,N_5902);
and U6147 (N_6147,N_5553,N_5892);
nor U6148 (N_6148,N_5798,N_5810);
xnor U6149 (N_6149,N_5637,N_5591);
and U6150 (N_6150,N_5683,N_5707);
nor U6151 (N_6151,N_5797,N_5855);
nor U6152 (N_6152,N_5896,N_5952);
and U6153 (N_6153,N_5644,N_5713);
and U6154 (N_6154,N_5843,N_5725);
nor U6155 (N_6155,N_5740,N_5916);
nand U6156 (N_6156,N_5996,N_5970);
nor U6157 (N_6157,N_5603,N_5794);
or U6158 (N_6158,N_5857,N_5989);
nor U6159 (N_6159,N_5932,N_5754);
nor U6160 (N_6160,N_5979,N_5525);
xor U6161 (N_6161,N_5623,N_5695);
and U6162 (N_6162,N_5849,N_5663);
or U6163 (N_6163,N_5765,N_5734);
nand U6164 (N_6164,N_5552,N_5983);
and U6165 (N_6165,N_5724,N_5874);
xnor U6166 (N_6166,N_5732,N_5572);
nand U6167 (N_6167,N_5787,N_5512);
or U6168 (N_6168,N_5540,N_5885);
nand U6169 (N_6169,N_5804,N_5755);
or U6170 (N_6170,N_5733,N_5689);
or U6171 (N_6171,N_5822,N_5836);
nor U6172 (N_6172,N_5821,N_5680);
nor U6173 (N_6173,N_5888,N_5883);
nand U6174 (N_6174,N_5616,N_5691);
and U6175 (N_6175,N_5792,N_5814);
and U6176 (N_6176,N_5802,N_5824);
nand U6177 (N_6177,N_5692,N_5575);
or U6178 (N_6178,N_5972,N_5581);
or U6179 (N_6179,N_5612,N_5538);
nor U6180 (N_6180,N_5750,N_5501);
xnor U6181 (N_6181,N_5988,N_5993);
nand U6182 (N_6182,N_5795,N_5830);
nor U6183 (N_6183,N_5748,N_5784);
nand U6184 (N_6184,N_5664,N_5719);
and U6185 (N_6185,N_5924,N_5991);
xor U6186 (N_6186,N_5769,N_5562);
nand U6187 (N_6187,N_5847,N_5871);
or U6188 (N_6188,N_5652,N_5648);
nand U6189 (N_6189,N_5901,N_5882);
xor U6190 (N_6190,N_5950,N_5532);
xnor U6191 (N_6191,N_5747,N_5844);
nand U6192 (N_6192,N_5771,N_5856);
xnor U6193 (N_6193,N_5729,N_5662);
and U6194 (N_6194,N_5791,N_5716);
nand U6195 (N_6195,N_5913,N_5526);
nor U6196 (N_6196,N_5508,N_5721);
and U6197 (N_6197,N_5963,N_5610);
or U6198 (N_6198,N_5870,N_5862);
and U6199 (N_6199,N_5604,N_5606);
and U6200 (N_6200,N_5812,N_5529);
and U6201 (N_6201,N_5876,N_5974);
nand U6202 (N_6202,N_5763,N_5548);
and U6203 (N_6203,N_5500,N_5943);
and U6204 (N_6204,N_5676,N_5776);
or U6205 (N_6205,N_5858,N_5960);
nor U6206 (N_6206,N_5967,N_5839);
xnor U6207 (N_6207,N_5520,N_5645);
nand U6208 (N_6208,N_5801,N_5775);
nor U6209 (N_6209,N_5762,N_5563);
or U6210 (N_6210,N_5560,N_5788);
nor U6211 (N_6211,N_5627,N_5640);
or U6212 (N_6212,N_5828,N_5953);
nor U6213 (N_6213,N_5785,N_5598);
nand U6214 (N_6214,N_5569,N_5502);
xnor U6215 (N_6215,N_5510,N_5594);
nand U6216 (N_6216,N_5561,N_5782);
and U6217 (N_6217,N_5897,N_5546);
nor U6218 (N_6218,N_5709,N_5833);
xor U6219 (N_6219,N_5927,N_5761);
nor U6220 (N_6220,N_5958,N_5854);
and U6221 (N_6221,N_5929,N_5660);
xnor U6222 (N_6222,N_5535,N_5767);
nand U6223 (N_6223,N_5906,N_5760);
nor U6224 (N_6224,N_5519,N_5587);
or U6225 (N_6225,N_5758,N_5954);
nand U6226 (N_6226,N_5935,N_5898);
or U6227 (N_6227,N_5649,N_5655);
and U6228 (N_6228,N_5982,N_5837);
nand U6229 (N_6229,N_5596,N_5539);
nor U6230 (N_6230,N_5962,N_5881);
or U6231 (N_6231,N_5853,N_5921);
xor U6232 (N_6232,N_5625,N_5613);
xnor U6233 (N_6233,N_5909,N_5727);
and U6234 (N_6234,N_5678,N_5714);
nor U6235 (N_6235,N_5522,N_5632);
nor U6236 (N_6236,N_5688,N_5568);
xor U6237 (N_6237,N_5601,N_5978);
and U6238 (N_6238,N_5764,N_5503);
nand U6239 (N_6239,N_5850,N_5614);
nor U6240 (N_6240,N_5800,N_5990);
or U6241 (N_6241,N_5743,N_5607);
and U6242 (N_6242,N_5537,N_5772);
and U6243 (N_6243,N_5745,N_5543);
xnor U6244 (N_6244,N_5907,N_5723);
nor U6245 (N_6245,N_5829,N_5701);
xnor U6246 (N_6246,N_5949,N_5693);
nor U6247 (N_6247,N_5513,N_5903);
nand U6248 (N_6248,N_5875,N_5749);
or U6249 (N_6249,N_5590,N_5946);
nor U6250 (N_6250,N_5931,N_5857);
nand U6251 (N_6251,N_5674,N_5947);
xor U6252 (N_6252,N_5569,N_5768);
nand U6253 (N_6253,N_5967,N_5950);
or U6254 (N_6254,N_5850,N_5648);
or U6255 (N_6255,N_5906,N_5539);
and U6256 (N_6256,N_5792,N_5766);
nand U6257 (N_6257,N_5571,N_5834);
nand U6258 (N_6258,N_5730,N_5986);
xnor U6259 (N_6259,N_5675,N_5752);
xor U6260 (N_6260,N_5697,N_5980);
xnor U6261 (N_6261,N_5833,N_5921);
nand U6262 (N_6262,N_5539,N_5589);
nor U6263 (N_6263,N_5589,N_5593);
and U6264 (N_6264,N_5541,N_5646);
or U6265 (N_6265,N_5819,N_5757);
and U6266 (N_6266,N_5728,N_5502);
or U6267 (N_6267,N_5579,N_5901);
and U6268 (N_6268,N_5618,N_5718);
and U6269 (N_6269,N_5619,N_5882);
xor U6270 (N_6270,N_5638,N_5729);
xnor U6271 (N_6271,N_5750,N_5917);
or U6272 (N_6272,N_5894,N_5755);
nor U6273 (N_6273,N_5985,N_5506);
or U6274 (N_6274,N_5786,N_5553);
nor U6275 (N_6275,N_5547,N_5511);
and U6276 (N_6276,N_5869,N_5764);
xor U6277 (N_6277,N_5568,N_5557);
nor U6278 (N_6278,N_5881,N_5653);
nand U6279 (N_6279,N_5809,N_5606);
nand U6280 (N_6280,N_5809,N_5882);
or U6281 (N_6281,N_5630,N_5501);
nor U6282 (N_6282,N_5792,N_5590);
or U6283 (N_6283,N_5684,N_5952);
nand U6284 (N_6284,N_5507,N_5781);
xnor U6285 (N_6285,N_5612,N_5585);
or U6286 (N_6286,N_5929,N_5959);
nor U6287 (N_6287,N_5842,N_5669);
nor U6288 (N_6288,N_5624,N_5533);
nand U6289 (N_6289,N_5667,N_5602);
or U6290 (N_6290,N_5968,N_5948);
nand U6291 (N_6291,N_5510,N_5977);
nor U6292 (N_6292,N_5958,N_5967);
nor U6293 (N_6293,N_5806,N_5553);
and U6294 (N_6294,N_5575,N_5673);
and U6295 (N_6295,N_5568,N_5947);
or U6296 (N_6296,N_5792,N_5555);
xnor U6297 (N_6297,N_5691,N_5819);
and U6298 (N_6298,N_5785,N_5902);
nor U6299 (N_6299,N_5755,N_5943);
nand U6300 (N_6300,N_5557,N_5772);
and U6301 (N_6301,N_5575,N_5902);
or U6302 (N_6302,N_5897,N_5852);
nor U6303 (N_6303,N_5935,N_5941);
xnor U6304 (N_6304,N_5854,N_5759);
or U6305 (N_6305,N_5561,N_5889);
and U6306 (N_6306,N_5827,N_5730);
nand U6307 (N_6307,N_5718,N_5782);
nand U6308 (N_6308,N_5668,N_5597);
xor U6309 (N_6309,N_5614,N_5651);
nor U6310 (N_6310,N_5537,N_5504);
or U6311 (N_6311,N_5617,N_5601);
or U6312 (N_6312,N_5583,N_5820);
or U6313 (N_6313,N_5657,N_5752);
and U6314 (N_6314,N_5833,N_5530);
or U6315 (N_6315,N_5558,N_5711);
and U6316 (N_6316,N_5839,N_5657);
or U6317 (N_6317,N_5955,N_5583);
or U6318 (N_6318,N_5573,N_5536);
nor U6319 (N_6319,N_5849,N_5831);
or U6320 (N_6320,N_5992,N_5698);
nor U6321 (N_6321,N_5893,N_5615);
and U6322 (N_6322,N_5936,N_5928);
xor U6323 (N_6323,N_5648,N_5861);
and U6324 (N_6324,N_5894,N_5658);
xnor U6325 (N_6325,N_5740,N_5596);
nor U6326 (N_6326,N_5587,N_5512);
nor U6327 (N_6327,N_5627,N_5560);
xnor U6328 (N_6328,N_5836,N_5916);
nor U6329 (N_6329,N_5839,N_5728);
or U6330 (N_6330,N_5582,N_5828);
nand U6331 (N_6331,N_5519,N_5887);
xor U6332 (N_6332,N_5884,N_5576);
nand U6333 (N_6333,N_5643,N_5989);
and U6334 (N_6334,N_5677,N_5752);
xnor U6335 (N_6335,N_5844,N_5902);
xnor U6336 (N_6336,N_5611,N_5760);
nand U6337 (N_6337,N_5673,N_5748);
nand U6338 (N_6338,N_5606,N_5520);
nand U6339 (N_6339,N_5636,N_5544);
and U6340 (N_6340,N_5808,N_5622);
nand U6341 (N_6341,N_5866,N_5762);
nor U6342 (N_6342,N_5575,N_5807);
and U6343 (N_6343,N_5793,N_5819);
nand U6344 (N_6344,N_5857,N_5554);
xor U6345 (N_6345,N_5825,N_5802);
or U6346 (N_6346,N_5562,N_5983);
xnor U6347 (N_6347,N_5644,N_5960);
nor U6348 (N_6348,N_5572,N_5550);
nor U6349 (N_6349,N_5578,N_5748);
xnor U6350 (N_6350,N_5564,N_5831);
and U6351 (N_6351,N_5842,N_5650);
xor U6352 (N_6352,N_5866,N_5535);
nor U6353 (N_6353,N_5992,N_5748);
nor U6354 (N_6354,N_5925,N_5635);
or U6355 (N_6355,N_5896,N_5799);
nor U6356 (N_6356,N_5768,N_5761);
nor U6357 (N_6357,N_5988,N_5629);
nor U6358 (N_6358,N_5899,N_5960);
xor U6359 (N_6359,N_5592,N_5661);
nor U6360 (N_6360,N_5531,N_5966);
nand U6361 (N_6361,N_5824,N_5723);
and U6362 (N_6362,N_5506,N_5619);
or U6363 (N_6363,N_5522,N_5737);
nand U6364 (N_6364,N_5738,N_5638);
xnor U6365 (N_6365,N_5926,N_5611);
and U6366 (N_6366,N_5680,N_5712);
xnor U6367 (N_6367,N_5691,N_5867);
nor U6368 (N_6368,N_5678,N_5516);
xnor U6369 (N_6369,N_5761,N_5861);
xnor U6370 (N_6370,N_5930,N_5991);
nor U6371 (N_6371,N_5503,N_5933);
and U6372 (N_6372,N_5742,N_5759);
or U6373 (N_6373,N_5708,N_5997);
nand U6374 (N_6374,N_5682,N_5697);
nor U6375 (N_6375,N_5800,N_5962);
and U6376 (N_6376,N_5565,N_5553);
or U6377 (N_6377,N_5628,N_5803);
nand U6378 (N_6378,N_5787,N_5925);
xor U6379 (N_6379,N_5853,N_5525);
nand U6380 (N_6380,N_5817,N_5878);
or U6381 (N_6381,N_5875,N_5590);
nor U6382 (N_6382,N_5999,N_5599);
nand U6383 (N_6383,N_5760,N_5723);
or U6384 (N_6384,N_5858,N_5673);
xor U6385 (N_6385,N_5995,N_5798);
nor U6386 (N_6386,N_5542,N_5638);
xnor U6387 (N_6387,N_5828,N_5588);
or U6388 (N_6388,N_5866,N_5969);
and U6389 (N_6389,N_5757,N_5842);
or U6390 (N_6390,N_5953,N_5774);
or U6391 (N_6391,N_5909,N_5537);
nand U6392 (N_6392,N_5982,N_5692);
nor U6393 (N_6393,N_5658,N_5633);
nand U6394 (N_6394,N_5731,N_5919);
nor U6395 (N_6395,N_5990,N_5693);
nand U6396 (N_6396,N_5851,N_5957);
or U6397 (N_6397,N_5918,N_5535);
xor U6398 (N_6398,N_5526,N_5967);
and U6399 (N_6399,N_5900,N_5505);
and U6400 (N_6400,N_5577,N_5765);
nand U6401 (N_6401,N_5899,N_5835);
or U6402 (N_6402,N_5602,N_5985);
and U6403 (N_6403,N_5513,N_5500);
xor U6404 (N_6404,N_5599,N_5816);
and U6405 (N_6405,N_5811,N_5870);
nor U6406 (N_6406,N_5662,N_5647);
xnor U6407 (N_6407,N_5945,N_5979);
or U6408 (N_6408,N_5896,N_5894);
or U6409 (N_6409,N_5993,N_5969);
or U6410 (N_6410,N_5981,N_5562);
nor U6411 (N_6411,N_5762,N_5676);
nor U6412 (N_6412,N_5907,N_5519);
and U6413 (N_6413,N_5528,N_5954);
nand U6414 (N_6414,N_5683,N_5578);
xor U6415 (N_6415,N_5737,N_5682);
and U6416 (N_6416,N_5978,N_5994);
xor U6417 (N_6417,N_5580,N_5638);
or U6418 (N_6418,N_5983,N_5942);
nor U6419 (N_6419,N_5764,N_5728);
and U6420 (N_6420,N_5891,N_5714);
and U6421 (N_6421,N_5987,N_5661);
xor U6422 (N_6422,N_5569,N_5872);
and U6423 (N_6423,N_5517,N_5914);
nor U6424 (N_6424,N_5720,N_5557);
nor U6425 (N_6425,N_5877,N_5747);
nor U6426 (N_6426,N_5575,N_5562);
and U6427 (N_6427,N_5642,N_5900);
xnor U6428 (N_6428,N_5646,N_5619);
or U6429 (N_6429,N_5917,N_5856);
and U6430 (N_6430,N_5888,N_5624);
nand U6431 (N_6431,N_5938,N_5631);
xor U6432 (N_6432,N_5884,N_5764);
xor U6433 (N_6433,N_5580,N_5548);
and U6434 (N_6434,N_5852,N_5784);
or U6435 (N_6435,N_5810,N_5828);
and U6436 (N_6436,N_5554,N_5906);
and U6437 (N_6437,N_5748,N_5610);
nor U6438 (N_6438,N_5566,N_5767);
and U6439 (N_6439,N_5655,N_5702);
or U6440 (N_6440,N_5957,N_5963);
nor U6441 (N_6441,N_5805,N_5607);
or U6442 (N_6442,N_5654,N_5993);
nor U6443 (N_6443,N_5598,N_5935);
xnor U6444 (N_6444,N_5600,N_5630);
or U6445 (N_6445,N_5958,N_5988);
nor U6446 (N_6446,N_5576,N_5741);
and U6447 (N_6447,N_5744,N_5771);
and U6448 (N_6448,N_5780,N_5652);
and U6449 (N_6449,N_5884,N_5515);
or U6450 (N_6450,N_5710,N_5792);
and U6451 (N_6451,N_5856,N_5522);
nor U6452 (N_6452,N_5905,N_5529);
or U6453 (N_6453,N_5636,N_5961);
and U6454 (N_6454,N_5875,N_5743);
and U6455 (N_6455,N_5570,N_5929);
xnor U6456 (N_6456,N_5799,N_5565);
or U6457 (N_6457,N_5927,N_5821);
xnor U6458 (N_6458,N_5591,N_5653);
xnor U6459 (N_6459,N_5905,N_5894);
nor U6460 (N_6460,N_5525,N_5541);
nor U6461 (N_6461,N_5822,N_5929);
nor U6462 (N_6462,N_5606,N_5998);
nand U6463 (N_6463,N_5996,N_5760);
nor U6464 (N_6464,N_5513,N_5815);
or U6465 (N_6465,N_5668,N_5920);
and U6466 (N_6466,N_5967,N_5529);
xnor U6467 (N_6467,N_5503,N_5590);
or U6468 (N_6468,N_5625,N_5898);
nor U6469 (N_6469,N_5769,N_5501);
and U6470 (N_6470,N_5996,N_5849);
and U6471 (N_6471,N_5938,N_5596);
or U6472 (N_6472,N_5967,N_5632);
and U6473 (N_6473,N_5975,N_5719);
nand U6474 (N_6474,N_5576,N_5559);
and U6475 (N_6475,N_5983,N_5939);
and U6476 (N_6476,N_5622,N_5530);
nand U6477 (N_6477,N_5743,N_5715);
xnor U6478 (N_6478,N_5788,N_5618);
nor U6479 (N_6479,N_5674,N_5637);
or U6480 (N_6480,N_5697,N_5713);
xor U6481 (N_6481,N_5804,N_5958);
nor U6482 (N_6482,N_5663,N_5539);
nor U6483 (N_6483,N_5610,N_5934);
nand U6484 (N_6484,N_5880,N_5943);
nand U6485 (N_6485,N_5529,N_5703);
xor U6486 (N_6486,N_5869,N_5775);
nand U6487 (N_6487,N_5520,N_5803);
xnor U6488 (N_6488,N_5885,N_5898);
xor U6489 (N_6489,N_5717,N_5527);
xor U6490 (N_6490,N_5815,N_5931);
xor U6491 (N_6491,N_5908,N_5852);
xnor U6492 (N_6492,N_5802,N_5769);
nor U6493 (N_6493,N_5526,N_5677);
xor U6494 (N_6494,N_5789,N_5553);
xor U6495 (N_6495,N_5537,N_5678);
xnor U6496 (N_6496,N_5801,N_5558);
or U6497 (N_6497,N_5973,N_5694);
nor U6498 (N_6498,N_5937,N_5799);
or U6499 (N_6499,N_5768,N_5577);
xor U6500 (N_6500,N_6301,N_6389);
nor U6501 (N_6501,N_6163,N_6381);
nor U6502 (N_6502,N_6114,N_6006);
xor U6503 (N_6503,N_6052,N_6143);
and U6504 (N_6504,N_6383,N_6087);
xnor U6505 (N_6505,N_6149,N_6127);
xor U6506 (N_6506,N_6132,N_6429);
xnor U6507 (N_6507,N_6042,N_6252);
nor U6508 (N_6508,N_6217,N_6165);
nand U6509 (N_6509,N_6162,N_6161);
xnor U6510 (N_6510,N_6287,N_6446);
xor U6511 (N_6511,N_6088,N_6219);
or U6512 (N_6512,N_6308,N_6311);
nor U6513 (N_6513,N_6228,N_6014);
nor U6514 (N_6514,N_6040,N_6216);
or U6515 (N_6515,N_6071,N_6321);
xor U6516 (N_6516,N_6164,N_6491);
nor U6517 (N_6517,N_6109,N_6101);
xnor U6518 (N_6518,N_6176,N_6498);
and U6519 (N_6519,N_6343,N_6017);
and U6520 (N_6520,N_6210,N_6255);
and U6521 (N_6521,N_6273,N_6489);
nand U6522 (N_6522,N_6118,N_6348);
xnor U6523 (N_6523,N_6371,N_6421);
and U6524 (N_6524,N_6449,N_6327);
xor U6525 (N_6525,N_6077,N_6465);
xor U6526 (N_6526,N_6471,N_6079);
nand U6527 (N_6527,N_6395,N_6278);
nand U6528 (N_6528,N_6001,N_6058);
or U6529 (N_6529,N_6485,N_6199);
and U6530 (N_6530,N_6072,N_6410);
or U6531 (N_6531,N_6106,N_6032);
nand U6532 (N_6532,N_6276,N_6335);
and U6533 (N_6533,N_6415,N_6112);
xor U6534 (N_6534,N_6248,N_6070);
and U6535 (N_6535,N_6055,N_6476);
nor U6536 (N_6536,N_6444,N_6379);
or U6537 (N_6537,N_6090,N_6263);
nand U6538 (N_6538,N_6150,N_6302);
nor U6539 (N_6539,N_6191,N_6495);
nand U6540 (N_6540,N_6221,N_6073);
nor U6541 (N_6541,N_6245,N_6043);
and U6542 (N_6542,N_6093,N_6294);
nand U6543 (N_6543,N_6051,N_6084);
xor U6544 (N_6544,N_6286,N_6213);
or U6545 (N_6545,N_6459,N_6303);
xnor U6546 (N_6546,N_6387,N_6212);
or U6547 (N_6547,N_6367,N_6416);
or U6548 (N_6548,N_6225,N_6095);
xor U6549 (N_6549,N_6400,N_6105);
and U6550 (N_6550,N_6102,N_6433);
and U6551 (N_6551,N_6128,N_6174);
xnor U6552 (N_6552,N_6440,N_6258);
or U6553 (N_6553,N_6204,N_6244);
nor U6554 (N_6554,N_6469,N_6190);
and U6555 (N_6555,N_6185,N_6307);
and U6556 (N_6556,N_6412,N_6352);
or U6557 (N_6557,N_6078,N_6354);
or U6558 (N_6558,N_6470,N_6281);
or U6559 (N_6559,N_6062,N_6194);
nor U6560 (N_6560,N_6430,N_6178);
and U6561 (N_6561,N_6130,N_6135);
xnor U6562 (N_6562,N_6115,N_6394);
xor U6563 (N_6563,N_6202,N_6414);
or U6564 (N_6564,N_6406,N_6365);
or U6565 (N_6565,N_6025,N_6325);
xor U6566 (N_6566,N_6240,N_6376);
or U6567 (N_6567,N_6427,N_6003);
nor U6568 (N_6568,N_6363,N_6175);
nand U6569 (N_6569,N_6155,N_6265);
nor U6570 (N_6570,N_6119,N_6493);
xor U6571 (N_6571,N_6349,N_6207);
nand U6572 (N_6572,N_6047,N_6408);
nand U6573 (N_6573,N_6405,N_6012);
and U6574 (N_6574,N_6438,N_6442);
nor U6575 (N_6575,N_6283,N_6329);
and U6576 (N_6576,N_6209,N_6401);
xnor U6577 (N_6577,N_6439,N_6499);
nor U6578 (N_6578,N_6274,N_6299);
xnor U6579 (N_6579,N_6375,N_6377);
and U6580 (N_6580,N_6324,N_6141);
or U6581 (N_6581,N_6111,N_6231);
xor U6582 (N_6582,N_6152,N_6230);
nor U6583 (N_6583,N_6447,N_6309);
nand U6584 (N_6584,N_6145,N_6494);
nor U6585 (N_6585,N_6063,N_6484);
nor U6586 (N_6586,N_6069,N_6186);
nand U6587 (N_6587,N_6188,N_6388);
nor U6588 (N_6588,N_6319,N_6172);
or U6589 (N_6589,N_6411,N_6249);
xnor U6590 (N_6590,N_6133,N_6113);
and U6591 (N_6591,N_6125,N_6466);
and U6592 (N_6592,N_6100,N_6288);
xnor U6593 (N_6593,N_6261,N_6167);
or U6594 (N_6594,N_6038,N_6369);
nor U6595 (N_6595,N_6253,N_6397);
nand U6596 (N_6596,N_6477,N_6214);
nand U6597 (N_6597,N_6378,N_6260);
and U6598 (N_6598,N_6323,N_6293);
or U6599 (N_6599,N_6462,N_6290);
and U6600 (N_6600,N_6305,N_6318);
or U6601 (N_6601,N_6487,N_6103);
xor U6602 (N_6602,N_6177,N_6220);
nor U6603 (N_6603,N_6392,N_6456);
xnor U6604 (N_6604,N_6269,N_6005);
and U6605 (N_6605,N_6390,N_6314);
nand U6606 (N_6606,N_6328,N_6479);
or U6607 (N_6607,N_6341,N_6346);
and U6608 (N_6608,N_6413,N_6226);
and U6609 (N_6609,N_6157,N_6002);
or U6610 (N_6610,N_6366,N_6009);
and U6611 (N_6611,N_6061,N_6297);
nor U6612 (N_6612,N_6180,N_6336);
nand U6613 (N_6613,N_6056,N_6268);
nand U6614 (N_6614,N_6277,N_6344);
nor U6615 (N_6615,N_6107,N_6312);
xnor U6616 (N_6616,N_6022,N_6361);
or U6617 (N_6617,N_6486,N_6004);
xor U6618 (N_6618,N_6173,N_6033);
nor U6619 (N_6619,N_6227,N_6028);
nand U6620 (N_6620,N_6048,N_6223);
xnor U6621 (N_6621,N_6151,N_6393);
nand U6622 (N_6622,N_6385,N_6422);
or U6623 (N_6623,N_6399,N_6086);
or U6624 (N_6624,N_6490,N_6126);
nor U6625 (N_6625,N_6436,N_6295);
or U6626 (N_6626,N_6315,N_6036);
and U6627 (N_6627,N_6235,N_6338);
and U6628 (N_6628,N_6085,N_6067);
xnor U6629 (N_6629,N_6262,N_6452);
or U6630 (N_6630,N_6306,N_6200);
or U6631 (N_6631,N_6454,N_6275);
xor U6632 (N_6632,N_6121,N_6171);
and U6633 (N_6633,N_6147,N_6030);
nand U6634 (N_6634,N_6254,N_6074);
xor U6635 (N_6635,N_6234,N_6098);
and U6636 (N_6636,N_6488,N_6224);
nand U6637 (N_6637,N_6148,N_6013);
or U6638 (N_6638,N_6313,N_6250);
nand U6639 (N_6639,N_6027,N_6448);
and U6640 (N_6640,N_6039,N_6453);
or U6641 (N_6641,N_6020,N_6187);
nor U6642 (N_6642,N_6168,N_6142);
nor U6643 (N_6643,N_6347,N_6316);
and U6644 (N_6644,N_6322,N_6082);
nor U6645 (N_6645,N_6026,N_6332);
and U6646 (N_6646,N_6007,N_6317);
and U6647 (N_6647,N_6360,N_6373);
and U6648 (N_6648,N_6053,N_6023);
or U6649 (N_6649,N_6131,N_6034);
nor U6650 (N_6650,N_6358,N_6296);
xor U6651 (N_6651,N_6140,N_6463);
and U6652 (N_6652,N_6496,N_6189);
or U6653 (N_6653,N_6357,N_6215);
xnor U6654 (N_6654,N_6257,N_6382);
nor U6655 (N_6655,N_6037,N_6356);
and U6656 (N_6656,N_6205,N_6169);
nand U6657 (N_6657,N_6068,N_6458);
xnor U6658 (N_6658,N_6451,N_6110);
nand U6659 (N_6659,N_6206,N_6242);
nand U6660 (N_6660,N_6368,N_6289);
and U6661 (N_6661,N_6256,N_6251);
or U6662 (N_6662,N_6492,N_6195);
and U6663 (N_6663,N_6179,N_6183);
nor U6664 (N_6664,N_6182,N_6460);
xor U6665 (N_6665,N_6247,N_6280);
xor U6666 (N_6666,N_6292,N_6457);
and U6667 (N_6667,N_6472,N_6218);
and U6668 (N_6668,N_6271,N_6091);
nor U6669 (N_6669,N_6331,N_6116);
nor U6670 (N_6670,N_6334,N_6031);
or U6671 (N_6671,N_6236,N_6021);
nor U6672 (N_6672,N_6246,N_6122);
nor U6673 (N_6673,N_6159,N_6450);
or U6674 (N_6674,N_6238,N_6426);
or U6675 (N_6675,N_6049,N_6089);
nor U6676 (N_6676,N_6419,N_6391);
and U6677 (N_6677,N_6066,N_6409);
nor U6678 (N_6678,N_6138,N_6282);
nor U6679 (N_6679,N_6266,N_6144);
or U6680 (N_6680,N_6480,N_6403);
and U6681 (N_6681,N_6351,N_6374);
or U6682 (N_6682,N_6229,N_6108);
nor U6683 (N_6683,N_6181,N_6298);
nor U6684 (N_6684,N_6284,N_6075);
or U6685 (N_6685,N_6264,N_6482);
nand U6686 (N_6686,N_6232,N_6473);
and U6687 (N_6687,N_6340,N_6418);
or U6688 (N_6688,N_6044,N_6104);
xnor U6689 (N_6689,N_6076,N_6483);
xnor U6690 (N_6690,N_6050,N_6123);
nor U6691 (N_6691,N_6211,N_6468);
xor U6692 (N_6692,N_6443,N_6279);
nor U6693 (N_6693,N_6441,N_6160);
or U6694 (N_6694,N_6241,N_6057);
nor U6695 (N_6695,N_6124,N_6337);
nand U6696 (N_6696,N_6402,N_6461);
nand U6697 (N_6697,N_6330,N_6478);
nor U6698 (N_6698,N_6139,N_6364);
and U6699 (N_6699,N_6092,N_6222);
xor U6700 (N_6700,N_6342,N_6407);
and U6701 (N_6701,N_6384,N_6184);
or U6702 (N_6702,N_6355,N_6203);
and U6703 (N_6703,N_6041,N_6080);
nor U6704 (N_6704,N_6239,N_6054);
and U6705 (N_6705,N_6060,N_6136);
nand U6706 (N_6706,N_6024,N_6000);
or U6707 (N_6707,N_6304,N_6158);
nor U6708 (N_6708,N_6166,N_6193);
or U6709 (N_6709,N_6497,N_6398);
and U6710 (N_6710,N_6016,N_6350);
nand U6711 (N_6711,N_6011,N_6435);
and U6712 (N_6712,N_6154,N_6475);
nor U6713 (N_6713,N_6197,N_6064);
or U6714 (N_6714,N_6156,N_6170);
or U6715 (N_6715,N_6134,N_6417);
or U6716 (N_6716,N_6423,N_6081);
or U6717 (N_6717,N_6035,N_6201);
and U6718 (N_6718,N_6474,N_6285);
or U6719 (N_6719,N_6481,N_6270);
and U6720 (N_6720,N_6320,N_6353);
xnor U6721 (N_6721,N_6097,N_6065);
and U6722 (N_6722,N_6464,N_6196);
or U6723 (N_6723,N_6326,N_6420);
xnor U6724 (N_6724,N_6008,N_6428);
or U6725 (N_6725,N_6018,N_6386);
or U6726 (N_6726,N_6117,N_6431);
or U6727 (N_6727,N_6272,N_6345);
xor U6728 (N_6728,N_6120,N_6445);
xor U6729 (N_6729,N_6359,N_6059);
nor U6730 (N_6730,N_6424,N_6083);
nand U6731 (N_6731,N_6099,N_6362);
nand U6732 (N_6732,N_6146,N_6333);
nand U6733 (N_6733,N_6370,N_6396);
or U6734 (N_6734,N_6310,N_6094);
nand U6735 (N_6735,N_6243,N_6029);
and U6736 (N_6736,N_6208,N_6432);
nand U6737 (N_6737,N_6237,N_6434);
xnor U6738 (N_6738,N_6339,N_6019);
nor U6739 (N_6739,N_6137,N_6437);
and U6740 (N_6740,N_6425,N_6259);
or U6741 (N_6741,N_6372,N_6015);
nand U6742 (N_6742,N_6380,N_6455);
or U6743 (N_6743,N_6467,N_6291);
xor U6744 (N_6744,N_6233,N_6096);
or U6745 (N_6745,N_6046,N_6300);
nor U6746 (N_6746,N_6129,N_6267);
nand U6747 (N_6747,N_6404,N_6010);
nand U6748 (N_6748,N_6153,N_6045);
and U6749 (N_6749,N_6198,N_6192);
nand U6750 (N_6750,N_6278,N_6495);
nand U6751 (N_6751,N_6358,N_6436);
and U6752 (N_6752,N_6416,N_6101);
xnor U6753 (N_6753,N_6087,N_6361);
xnor U6754 (N_6754,N_6485,N_6073);
xnor U6755 (N_6755,N_6107,N_6390);
nand U6756 (N_6756,N_6283,N_6491);
xor U6757 (N_6757,N_6311,N_6460);
xnor U6758 (N_6758,N_6211,N_6359);
and U6759 (N_6759,N_6193,N_6333);
xnor U6760 (N_6760,N_6345,N_6273);
and U6761 (N_6761,N_6313,N_6055);
and U6762 (N_6762,N_6188,N_6042);
nor U6763 (N_6763,N_6001,N_6022);
nor U6764 (N_6764,N_6320,N_6162);
and U6765 (N_6765,N_6331,N_6319);
and U6766 (N_6766,N_6359,N_6013);
or U6767 (N_6767,N_6339,N_6343);
and U6768 (N_6768,N_6064,N_6416);
and U6769 (N_6769,N_6048,N_6481);
nor U6770 (N_6770,N_6289,N_6454);
or U6771 (N_6771,N_6496,N_6063);
nor U6772 (N_6772,N_6403,N_6319);
nand U6773 (N_6773,N_6167,N_6145);
nor U6774 (N_6774,N_6071,N_6448);
xor U6775 (N_6775,N_6473,N_6286);
nor U6776 (N_6776,N_6057,N_6110);
nor U6777 (N_6777,N_6019,N_6134);
xor U6778 (N_6778,N_6142,N_6198);
or U6779 (N_6779,N_6415,N_6079);
or U6780 (N_6780,N_6261,N_6486);
nand U6781 (N_6781,N_6415,N_6362);
nor U6782 (N_6782,N_6480,N_6455);
or U6783 (N_6783,N_6128,N_6442);
or U6784 (N_6784,N_6395,N_6029);
xor U6785 (N_6785,N_6335,N_6394);
xor U6786 (N_6786,N_6017,N_6493);
nand U6787 (N_6787,N_6100,N_6121);
nand U6788 (N_6788,N_6086,N_6059);
xor U6789 (N_6789,N_6071,N_6141);
nor U6790 (N_6790,N_6479,N_6421);
or U6791 (N_6791,N_6154,N_6111);
nor U6792 (N_6792,N_6000,N_6341);
nor U6793 (N_6793,N_6050,N_6061);
and U6794 (N_6794,N_6072,N_6436);
nand U6795 (N_6795,N_6188,N_6199);
and U6796 (N_6796,N_6093,N_6080);
nand U6797 (N_6797,N_6379,N_6243);
nand U6798 (N_6798,N_6255,N_6147);
and U6799 (N_6799,N_6284,N_6484);
xor U6800 (N_6800,N_6385,N_6206);
and U6801 (N_6801,N_6395,N_6092);
nand U6802 (N_6802,N_6398,N_6449);
nand U6803 (N_6803,N_6309,N_6279);
xnor U6804 (N_6804,N_6138,N_6328);
and U6805 (N_6805,N_6042,N_6183);
or U6806 (N_6806,N_6204,N_6455);
nor U6807 (N_6807,N_6498,N_6406);
xor U6808 (N_6808,N_6393,N_6236);
or U6809 (N_6809,N_6231,N_6205);
nor U6810 (N_6810,N_6216,N_6198);
and U6811 (N_6811,N_6252,N_6439);
and U6812 (N_6812,N_6041,N_6103);
xnor U6813 (N_6813,N_6341,N_6290);
xnor U6814 (N_6814,N_6271,N_6295);
and U6815 (N_6815,N_6217,N_6306);
xor U6816 (N_6816,N_6048,N_6255);
and U6817 (N_6817,N_6156,N_6254);
or U6818 (N_6818,N_6395,N_6301);
xnor U6819 (N_6819,N_6267,N_6331);
xnor U6820 (N_6820,N_6448,N_6097);
nor U6821 (N_6821,N_6117,N_6359);
xor U6822 (N_6822,N_6174,N_6344);
and U6823 (N_6823,N_6327,N_6069);
and U6824 (N_6824,N_6390,N_6152);
xor U6825 (N_6825,N_6498,N_6043);
and U6826 (N_6826,N_6113,N_6482);
nand U6827 (N_6827,N_6225,N_6258);
nand U6828 (N_6828,N_6365,N_6399);
or U6829 (N_6829,N_6386,N_6039);
xor U6830 (N_6830,N_6312,N_6207);
nor U6831 (N_6831,N_6448,N_6171);
or U6832 (N_6832,N_6069,N_6262);
and U6833 (N_6833,N_6121,N_6195);
xnor U6834 (N_6834,N_6364,N_6420);
or U6835 (N_6835,N_6439,N_6294);
or U6836 (N_6836,N_6185,N_6063);
or U6837 (N_6837,N_6067,N_6203);
nand U6838 (N_6838,N_6077,N_6417);
and U6839 (N_6839,N_6466,N_6010);
and U6840 (N_6840,N_6284,N_6316);
nor U6841 (N_6841,N_6396,N_6474);
nand U6842 (N_6842,N_6163,N_6226);
or U6843 (N_6843,N_6410,N_6277);
and U6844 (N_6844,N_6438,N_6416);
and U6845 (N_6845,N_6051,N_6286);
and U6846 (N_6846,N_6367,N_6209);
xnor U6847 (N_6847,N_6401,N_6178);
or U6848 (N_6848,N_6136,N_6296);
or U6849 (N_6849,N_6347,N_6379);
nor U6850 (N_6850,N_6220,N_6481);
or U6851 (N_6851,N_6182,N_6300);
xnor U6852 (N_6852,N_6378,N_6054);
nand U6853 (N_6853,N_6374,N_6330);
xnor U6854 (N_6854,N_6373,N_6044);
nand U6855 (N_6855,N_6165,N_6489);
xor U6856 (N_6856,N_6145,N_6085);
xnor U6857 (N_6857,N_6194,N_6196);
nand U6858 (N_6858,N_6448,N_6145);
or U6859 (N_6859,N_6189,N_6183);
and U6860 (N_6860,N_6235,N_6085);
nor U6861 (N_6861,N_6067,N_6275);
nand U6862 (N_6862,N_6201,N_6076);
xor U6863 (N_6863,N_6075,N_6058);
or U6864 (N_6864,N_6481,N_6072);
nor U6865 (N_6865,N_6452,N_6004);
or U6866 (N_6866,N_6441,N_6412);
xnor U6867 (N_6867,N_6051,N_6269);
and U6868 (N_6868,N_6379,N_6034);
and U6869 (N_6869,N_6420,N_6356);
nand U6870 (N_6870,N_6435,N_6241);
or U6871 (N_6871,N_6182,N_6063);
xnor U6872 (N_6872,N_6131,N_6457);
and U6873 (N_6873,N_6296,N_6337);
or U6874 (N_6874,N_6236,N_6470);
xor U6875 (N_6875,N_6329,N_6397);
nor U6876 (N_6876,N_6143,N_6225);
and U6877 (N_6877,N_6229,N_6469);
nor U6878 (N_6878,N_6176,N_6448);
xnor U6879 (N_6879,N_6151,N_6392);
nor U6880 (N_6880,N_6196,N_6371);
xor U6881 (N_6881,N_6397,N_6474);
xnor U6882 (N_6882,N_6280,N_6359);
and U6883 (N_6883,N_6243,N_6331);
or U6884 (N_6884,N_6081,N_6059);
xnor U6885 (N_6885,N_6284,N_6401);
nor U6886 (N_6886,N_6297,N_6067);
or U6887 (N_6887,N_6191,N_6027);
nand U6888 (N_6888,N_6032,N_6257);
xor U6889 (N_6889,N_6012,N_6155);
nand U6890 (N_6890,N_6443,N_6482);
xnor U6891 (N_6891,N_6148,N_6006);
xor U6892 (N_6892,N_6133,N_6356);
nand U6893 (N_6893,N_6402,N_6123);
nand U6894 (N_6894,N_6440,N_6080);
and U6895 (N_6895,N_6000,N_6284);
or U6896 (N_6896,N_6371,N_6404);
or U6897 (N_6897,N_6148,N_6272);
nand U6898 (N_6898,N_6372,N_6156);
nand U6899 (N_6899,N_6425,N_6022);
nor U6900 (N_6900,N_6455,N_6434);
xnor U6901 (N_6901,N_6099,N_6162);
and U6902 (N_6902,N_6027,N_6253);
xnor U6903 (N_6903,N_6214,N_6428);
nand U6904 (N_6904,N_6287,N_6133);
nand U6905 (N_6905,N_6485,N_6278);
xor U6906 (N_6906,N_6473,N_6061);
nor U6907 (N_6907,N_6342,N_6104);
xnor U6908 (N_6908,N_6144,N_6281);
nand U6909 (N_6909,N_6223,N_6350);
and U6910 (N_6910,N_6337,N_6317);
nand U6911 (N_6911,N_6186,N_6247);
or U6912 (N_6912,N_6338,N_6292);
and U6913 (N_6913,N_6315,N_6057);
xnor U6914 (N_6914,N_6312,N_6444);
xor U6915 (N_6915,N_6436,N_6207);
nand U6916 (N_6916,N_6070,N_6002);
and U6917 (N_6917,N_6082,N_6424);
or U6918 (N_6918,N_6494,N_6414);
or U6919 (N_6919,N_6439,N_6231);
and U6920 (N_6920,N_6101,N_6220);
xor U6921 (N_6921,N_6041,N_6016);
nand U6922 (N_6922,N_6065,N_6397);
or U6923 (N_6923,N_6041,N_6127);
or U6924 (N_6924,N_6491,N_6192);
nor U6925 (N_6925,N_6106,N_6382);
nand U6926 (N_6926,N_6142,N_6066);
nand U6927 (N_6927,N_6441,N_6341);
and U6928 (N_6928,N_6059,N_6076);
xor U6929 (N_6929,N_6038,N_6250);
xor U6930 (N_6930,N_6334,N_6262);
and U6931 (N_6931,N_6401,N_6223);
and U6932 (N_6932,N_6109,N_6313);
xnor U6933 (N_6933,N_6033,N_6199);
nand U6934 (N_6934,N_6339,N_6310);
and U6935 (N_6935,N_6339,N_6267);
nor U6936 (N_6936,N_6175,N_6005);
xor U6937 (N_6937,N_6407,N_6348);
nand U6938 (N_6938,N_6394,N_6289);
nand U6939 (N_6939,N_6176,N_6399);
or U6940 (N_6940,N_6378,N_6436);
nor U6941 (N_6941,N_6429,N_6410);
or U6942 (N_6942,N_6272,N_6241);
nor U6943 (N_6943,N_6240,N_6089);
nand U6944 (N_6944,N_6402,N_6437);
xor U6945 (N_6945,N_6314,N_6140);
xor U6946 (N_6946,N_6077,N_6253);
nor U6947 (N_6947,N_6035,N_6409);
nor U6948 (N_6948,N_6396,N_6058);
and U6949 (N_6949,N_6243,N_6466);
xor U6950 (N_6950,N_6246,N_6372);
or U6951 (N_6951,N_6042,N_6433);
nand U6952 (N_6952,N_6019,N_6241);
xnor U6953 (N_6953,N_6454,N_6282);
nor U6954 (N_6954,N_6002,N_6106);
and U6955 (N_6955,N_6223,N_6066);
and U6956 (N_6956,N_6046,N_6321);
nand U6957 (N_6957,N_6072,N_6077);
xnor U6958 (N_6958,N_6301,N_6317);
nor U6959 (N_6959,N_6072,N_6146);
xnor U6960 (N_6960,N_6108,N_6145);
and U6961 (N_6961,N_6065,N_6262);
and U6962 (N_6962,N_6451,N_6014);
xnor U6963 (N_6963,N_6375,N_6073);
and U6964 (N_6964,N_6150,N_6119);
xor U6965 (N_6965,N_6313,N_6107);
nor U6966 (N_6966,N_6457,N_6161);
nor U6967 (N_6967,N_6280,N_6487);
nor U6968 (N_6968,N_6005,N_6276);
nand U6969 (N_6969,N_6177,N_6386);
or U6970 (N_6970,N_6166,N_6230);
and U6971 (N_6971,N_6194,N_6070);
xor U6972 (N_6972,N_6280,N_6440);
xnor U6973 (N_6973,N_6095,N_6097);
nor U6974 (N_6974,N_6439,N_6395);
nand U6975 (N_6975,N_6293,N_6492);
nand U6976 (N_6976,N_6171,N_6287);
or U6977 (N_6977,N_6217,N_6366);
xor U6978 (N_6978,N_6142,N_6022);
nand U6979 (N_6979,N_6173,N_6280);
nor U6980 (N_6980,N_6360,N_6458);
xnor U6981 (N_6981,N_6289,N_6212);
xnor U6982 (N_6982,N_6056,N_6364);
xnor U6983 (N_6983,N_6167,N_6296);
nand U6984 (N_6984,N_6395,N_6169);
or U6985 (N_6985,N_6481,N_6160);
nor U6986 (N_6986,N_6289,N_6304);
nor U6987 (N_6987,N_6462,N_6054);
or U6988 (N_6988,N_6155,N_6166);
or U6989 (N_6989,N_6318,N_6097);
xnor U6990 (N_6990,N_6189,N_6455);
xor U6991 (N_6991,N_6430,N_6294);
xnor U6992 (N_6992,N_6396,N_6285);
xor U6993 (N_6993,N_6390,N_6467);
nor U6994 (N_6994,N_6001,N_6345);
and U6995 (N_6995,N_6329,N_6060);
or U6996 (N_6996,N_6325,N_6310);
nor U6997 (N_6997,N_6254,N_6203);
and U6998 (N_6998,N_6177,N_6323);
and U6999 (N_6999,N_6057,N_6355);
nand U7000 (N_7000,N_6568,N_6527);
and U7001 (N_7001,N_6944,N_6861);
and U7002 (N_7002,N_6851,N_6728);
nand U7003 (N_7003,N_6757,N_6597);
and U7004 (N_7004,N_6819,N_6781);
nand U7005 (N_7005,N_6760,N_6892);
nor U7006 (N_7006,N_6794,N_6839);
nand U7007 (N_7007,N_6906,N_6883);
nand U7008 (N_7008,N_6695,N_6809);
xnor U7009 (N_7009,N_6814,N_6535);
nor U7010 (N_7010,N_6684,N_6920);
nand U7011 (N_7011,N_6556,N_6987);
nand U7012 (N_7012,N_6507,N_6899);
nand U7013 (N_7013,N_6835,N_6855);
and U7014 (N_7014,N_6563,N_6617);
nand U7015 (N_7015,N_6529,N_6665);
nor U7016 (N_7016,N_6746,N_6661);
nor U7017 (N_7017,N_6744,N_6629);
and U7018 (N_7018,N_6618,N_6959);
xnor U7019 (N_7019,N_6748,N_6868);
nand U7020 (N_7020,N_6824,N_6612);
nor U7021 (N_7021,N_6997,N_6513);
nor U7022 (N_7022,N_6936,N_6631);
nand U7023 (N_7023,N_6880,N_6626);
nand U7024 (N_7024,N_6914,N_6860);
nand U7025 (N_7025,N_6820,N_6532);
nor U7026 (N_7026,N_6610,N_6589);
xnor U7027 (N_7027,N_6557,N_6667);
and U7028 (N_7028,N_6866,N_6601);
nand U7029 (N_7029,N_6831,N_6699);
nand U7030 (N_7030,N_6523,N_6521);
or U7031 (N_7031,N_6570,N_6700);
and U7032 (N_7032,N_6766,N_6600);
xnor U7033 (N_7033,N_6953,N_6594);
nand U7034 (N_7034,N_6782,N_6550);
xnor U7035 (N_7035,N_6873,N_6727);
xor U7036 (N_7036,N_6706,N_6984);
xor U7037 (N_7037,N_6951,N_6796);
nor U7038 (N_7038,N_6554,N_6526);
and U7039 (N_7039,N_6952,N_6965);
nand U7040 (N_7040,N_6547,N_6580);
nand U7041 (N_7041,N_6683,N_6714);
and U7042 (N_7042,N_6925,N_6614);
and U7043 (N_7043,N_6514,N_6697);
nor U7044 (N_7044,N_6886,N_6982);
xnor U7045 (N_7045,N_6551,N_6985);
xnor U7046 (N_7046,N_6719,N_6937);
nor U7047 (N_7047,N_6871,N_6756);
and U7048 (N_7048,N_6694,N_6623);
nand U7049 (N_7049,N_6518,N_6670);
or U7050 (N_7050,N_6804,N_6869);
nand U7051 (N_7051,N_6715,N_6764);
or U7052 (N_7052,N_6891,N_6639);
and U7053 (N_7053,N_6765,N_6912);
xor U7054 (N_7054,N_6864,N_6789);
or U7055 (N_7055,N_6785,N_6910);
xnor U7056 (N_7056,N_6818,N_6774);
nor U7057 (N_7057,N_6652,N_6896);
and U7058 (N_7058,N_6770,N_6988);
nand U7059 (N_7059,N_6561,N_6622);
xnor U7060 (N_7060,N_6674,N_6564);
nand U7061 (N_7061,N_6758,N_6691);
xor U7062 (N_7062,N_6917,N_6929);
nand U7063 (N_7063,N_6799,N_6608);
nand U7064 (N_7064,N_6994,N_6669);
xor U7065 (N_7065,N_6741,N_6558);
xor U7066 (N_7066,N_6957,N_6844);
nor U7067 (N_7067,N_6935,N_6897);
nor U7068 (N_7068,N_6907,N_6689);
and U7069 (N_7069,N_6771,N_6901);
xor U7070 (N_7070,N_6945,N_6606);
nand U7071 (N_7071,N_6878,N_6668);
nor U7072 (N_7072,N_6501,N_6811);
xor U7073 (N_7073,N_6792,N_6732);
or U7074 (N_7074,N_6575,N_6671);
nor U7075 (N_7075,N_6701,N_6979);
or U7076 (N_7076,N_6967,N_6643);
xor U7077 (N_7077,N_6676,N_6759);
nor U7078 (N_7078,N_6640,N_6660);
xor U7079 (N_7079,N_6578,N_6857);
xnor U7080 (N_7080,N_6881,N_6808);
or U7081 (N_7081,N_6533,N_6615);
and U7082 (N_7082,N_6971,N_6648);
xor U7083 (N_7083,N_6582,N_6711);
or U7084 (N_7084,N_6534,N_6609);
or U7085 (N_7085,N_6928,N_6562);
xnor U7086 (N_7086,N_6571,N_6955);
or U7087 (N_7087,N_6773,N_6963);
nor U7088 (N_7088,N_6680,N_6546);
xnor U7089 (N_7089,N_6520,N_6974);
or U7090 (N_7090,N_6877,N_6713);
or U7091 (N_7091,N_6583,N_6595);
and U7092 (N_7092,N_6560,N_6911);
or U7093 (N_7093,N_6704,N_6565);
xor U7094 (N_7094,N_6736,N_6509);
nor U7095 (N_7095,N_6502,N_6602);
xor U7096 (N_7096,N_6593,N_6823);
nand U7097 (N_7097,N_6947,N_6887);
nor U7098 (N_7098,N_6599,N_6613);
xor U7099 (N_7099,N_6553,N_6921);
and U7100 (N_7100,N_6948,N_6777);
and U7101 (N_7101,N_6707,N_6666);
nand U7102 (N_7102,N_6567,N_6503);
xor U7103 (N_7103,N_6751,N_6703);
nor U7104 (N_7104,N_6693,N_6651);
xnor U7105 (N_7105,N_6506,N_6934);
or U7106 (N_7106,N_6784,N_6552);
and U7107 (N_7107,N_6656,N_6510);
or U7108 (N_7108,N_6817,N_6747);
or U7109 (N_7109,N_6730,N_6650);
nor U7110 (N_7110,N_6950,N_6752);
nor U7111 (N_7111,N_6678,N_6696);
and U7112 (N_7112,N_6605,N_6592);
xnor U7113 (N_7113,N_6903,N_6685);
xnor U7114 (N_7114,N_6628,N_6588);
and U7115 (N_7115,N_6603,N_6902);
nor U7116 (N_7116,N_6939,N_6576);
xnor U7117 (N_7117,N_6976,N_6893);
and U7118 (N_7118,N_6772,N_6522);
xnor U7119 (N_7119,N_6989,N_6904);
nand U7120 (N_7120,N_6821,N_6972);
xor U7121 (N_7121,N_6806,N_6637);
nor U7122 (N_7122,N_6733,N_6717);
nor U7123 (N_7123,N_6649,N_6634);
xor U7124 (N_7124,N_6517,N_6739);
nand U7125 (N_7125,N_6702,N_6916);
xor U7126 (N_7126,N_6977,N_6919);
and U7127 (N_7127,N_6926,N_6783);
and U7128 (N_7128,N_6611,N_6810);
xnor U7129 (N_7129,N_6827,N_6712);
xnor U7130 (N_7130,N_6743,N_6981);
nor U7131 (N_7131,N_6826,N_6983);
nor U7132 (N_7132,N_6793,N_6538);
or U7133 (N_7133,N_6978,N_6800);
or U7134 (N_7134,N_6962,N_6731);
xor U7135 (N_7135,N_6973,N_6734);
nand U7136 (N_7136,N_6769,N_6627);
and U7137 (N_7137,N_6544,N_6812);
nand U7138 (N_7138,N_6745,N_6659);
or U7139 (N_7139,N_6579,N_6942);
nand U7140 (N_7140,N_6813,N_6585);
nor U7141 (N_7141,N_6619,N_6598);
or U7142 (N_7142,N_6716,N_6632);
nand U7143 (N_7143,N_6569,N_6581);
nand U7144 (N_7144,N_6710,N_6761);
xnor U7145 (N_7145,N_6616,N_6607);
or U7146 (N_7146,N_6923,N_6858);
nor U7147 (N_7147,N_6927,N_6688);
xor U7148 (N_7148,N_6961,N_6768);
xor U7149 (N_7149,N_6729,N_6918);
nand U7150 (N_7150,N_6762,N_6995);
and U7151 (N_7151,N_6508,N_6655);
nor U7152 (N_7152,N_6642,N_6980);
or U7153 (N_7153,N_6686,N_6735);
nor U7154 (N_7154,N_6644,N_6537);
nor U7155 (N_7155,N_6540,N_6624);
and U7156 (N_7156,N_6924,N_6549);
or U7157 (N_7157,N_6932,N_6663);
xor U7158 (N_7158,N_6991,N_6572);
or U7159 (N_7159,N_6705,N_6797);
or U7160 (N_7160,N_6675,N_6874);
or U7161 (N_7161,N_6949,N_6885);
nand U7162 (N_7162,N_6815,N_6836);
xor U7163 (N_7163,N_6516,N_6875);
and U7164 (N_7164,N_6723,N_6833);
or U7165 (N_7165,N_6838,N_6940);
nand U7166 (N_7166,N_6620,N_6519);
xnor U7167 (N_7167,N_6834,N_6867);
and U7168 (N_7168,N_6960,N_6573);
nor U7169 (N_7169,N_6725,N_6726);
nand U7170 (N_7170,N_6658,N_6905);
nand U7171 (N_7171,N_6722,N_6930);
nor U7172 (N_7172,N_6946,N_6798);
xor U7173 (N_7173,N_6841,N_6590);
xnor U7174 (N_7174,N_6890,N_6692);
and U7175 (N_7175,N_6788,N_6657);
and U7176 (N_7176,N_6763,N_6690);
xnor U7177 (N_7177,N_6536,N_6908);
and U7178 (N_7178,N_6641,N_6755);
nand U7179 (N_7179,N_6673,N_6913);
or U7180 (N_7180,N_6512,N_6698);
or U7181 (N_7181,N_6956,N_6721);
nor U7182 (N_7182,N_6970,N_6876);
or U7183 (N_7183,N_6966,N_6647);
and U7184 (N_7184,N_6822,N_6882);
nand U7185 (N_7185,N_6630,N_6559);
xor U7186 (N_7186,N_6879,N_6786);
nand U7187 (N_7187,N_6845,N_6504);
and U7188 (N_7188,N_6586,N_6825);
xnor U7189 (N_7189,N_6718,N_6847);
and U7190 (N_7190,N_6975,N_6574);
xnor U7191 (N_7191,N_6753,N_6832);
nand U7192 (N_7192,N_6709,N_6852);
or U7193 (N_7193,N_6587,N_6775);
nand U7194 (N_7194,N_6954,N_6604);
xor U7195 (N_7195,N_6635,N_6708);
and U7196 (N_7196,N_6802,N_6922);
nand U7197 (N_7197,N_6999,N_6993);
nor U7198 (N_7198,N_6941,N_6842);
xnor U7199 (N_7199,N_6500,N_6662);
nand U7200 (N_7200,N_6848,N_6870);
nor U7201 (N_7201,N_6515,N_6645);
xnor U7202 (N_7202,N_6646,N_6895);
or U7203 (N_7203,N_6633,N_6681);
nand U7204 (N_7204,N_6525,N_6889);
xnor U7205 (N_7205,N_6801,N_6779);
nand U7206 (N_7206,N_6542,N_6687);
nor U7207 (N_7207,N_6566,N_6964);
nand U7208 (N_7208,N_6530,N_6969);
xnor U7209 (N_7209,N_6539,N_6653);
and U7210 (N_7210,N_6767,N_6859);
and U7211 (N_7211,N_6545,N_6863);
xor U7212 (N_7212,N_6742,N_6780);
or U7213 (N_7213,N_6664,N_6931);
and U7214 (N_7214,N_6596,N_6720);
nor U7215 (N_7215,N_6998,N_6790);
nand U7216 (N_7216,N_6958,N_6738);
and U7217 (N_7217,N_6828,N_6840);
and U7218 (N_7218,N_6621,N_6791);
and U7219 (N_7219,N_6591,N_6778);
nor U7220 (N_7220,N_6843,N_6737);
xor U7221 (N_7221,N_6577,N_6830);
or U7222 (N_7222,N_6853,N_6943);
xor U7223 (N_7223,N_6541,N_6872);
xnor U7224 (N_7224,N_6584,N_6888);
or U7225 (N_7225,N_6865,N_6749);
and U7226 (N_7226,N_6636,N_6990);
xnor U7227 (N_7227,N_6900,N_6511);
or U7228 (N_7228,N_6807,N_6909);
or U7229 (N_7229,N_6654,N_6933);
xnor U7230 (N_7230,N_6805,N_6846);
and U7231 (N_7231,N_6795,N_6754);
and U7232 (N_7232,N_6531,N_6850);
nor U7233 (N_7233,N_6968,N_6740);
and U7234 (N_7234,N_6524,N_6682);
or U7235 (N_7235,N_6829,N_6862);
xnor U7236 (N_7236,N_6996,N_6816);
and U7237 (N_7237,N_6679,N_6837);
nor U7238 (N_7238,N_6787,N_6938);
and U7239 (N_7239,N_6677,N_6724);
nand U7240 (N_7240,N_6849,N_6638);
nand U7241 (N_7241,N_6894,N_6548);
or U7242 (N_7242,N_6992,N_6528);
or U7243 (N_7243,N_6750,N_6803);
or U7244 (N_7244,N_6915,N_6672);
xnor U7245 (N_7245,N_6555,N_6856);
nor U7246 (N_7246,N_6505,N_6543);
or U7247 (N_7247,N_6854,N_6898);
nand U7248 (N_7248,N_6884,N_6625);
nand U7249 (N_7249,N_6986,N_6776);
and U7250 (N_7250,N_6501,N_6968);
nand U7251 (N_7251,N_6647,N_6638);
nor U7252 (N_7252,N_6701,N_6727);
or U7253 (N_7253,N_6625,N_6768);
xor U7254 (N_7254,N_6958,N_6509);
xnor U7255 (N_7255,N_6611,N_6806);
nand U7256 (N_7256,N_6994,N_6813);
nor U7257 (N_7257,N_6592,N_6868);
nand U7258 (N_7258,N_6850,N_6734);
or U7259 (N_7259,N_6710,N_6847);
and U7260 (N_7260,N_6765,N_6916);
nand U7261 (N_7261,N_6758,N_6852);
xnor U7262 (N_7262,N_6625,N_6507);
xor U7263 (N_7263,N_6800,N_6581);
nand U7264 (N_7264,N_6683,N_6832);
nor U7265 (N_7265,N_6506,N_6542);
and U7266 (N_7266,N_6945,N_6808);
or U7267 (N_7267,N_6537,N_6650);
nand U7268 (N_7268,N_6658,N_6508);
and U7269 (N_7269,N_6671,N_6754);
nand U7270 (N_7270,N_6734,N_6510);
xnor U7271 (N_7271,N_6846,N_6908);
nor U7272 (N_7272,N_6877,N_6900);
xor U7273 (N_7273,N_6516,N_6938);
xor U7274 (N_7274,N_6566,N_6557);
nand U7275 (N_7275,N_6786,N_6657);
nor U7276 (N_7276,N_6582,N_6988);
nor U7277 (N_7277,N_6818,N_6832);
nand U7278 (N_7278,N_6653,N_6903);
xnor U7279 (N_7279,N_6823,N_6821);
or U7280 (N_7280,N_6951,N_6553);
nand U7281 (N_7281,N_6968,N_6570);
and U7282 (N_7282,N_6936,N_6730);
and U7283 (N_7283,N_6812,N_6682);
xor U7284 (N_7284,N_6861,N_6977);
and U7285 (N_7285,N_6670,N_6659);
or U7286 (N_7286,N_6921,N_6963);
nand U7287 (N_7287,N_6598,N_6509);
or U7288 (N_7288,N_6626,N_6777);
nor U7289 (N_7289,N_6649,N_6836);
or U7290 (N_7290,N_6575,N_6870);
and U7291 (N_7291,N_6660,N_6999);
or U7292 (N_7292,N_6652,N_6741);
and U7293 (N_7293,N_6748,N_6594);
nor U7294 (N_7294,N_6792,N_6864);
nor U7295 (N_7295,N_6557,N_6894);
and U7296 (N_7296,N_6868,N_6619);
or U7297 (N_7297,N_6942,N_6846);
nor U7298 (N_7298,N_6752,N_6534);
xor U7299 (N_7299,N_6656,N_6610);
nor U7300 (N_7300,N_6548,N_6639);
and U7301 (N_7301,N_6701,N_6999);
nor U7302 (N_7302,N_6507,N_6641);
or U7303 (N_7303,N_6650,N_6889);
or U7304 (N_7304,N_6864,N_6573);
or U7305 (N_7305,N_6917,N_6902);
or U7306 (N_7306,N_6876,N_6975);
nand U7307 (N_7307,N_6750,N_6701);
xnor U7308 (N_7308,N_6588,N_6599);
nand U7309 (N_7309,N_6786,N_6862);
xor U7310 (N_7310,N_6900,N_6888);
and U7311 (N_7311,N_6533,N_6804);
and U7312 (N_7312,N_6766,N_6617);
nor U7313 (N_7313,N_6777,N_6724);
nor U7314 (N_7314,N_6571,N_6608);
or U7315 (N_7315,N_6780,N_6826);
or U7316 (N_7316,N_6939,N_6927);
xor U7317 (N_7317,N_6908,N_6742);
or U7318 (N_7318,N_6747,N_6553);
and U7319 (N_7319,N_6556,N_6552);
nand U7320 (N_7320,N_6942,N_6511);
xor U7321 (N_7321,N_6865,N_6935);
nor U7322 (N_7322,N_6971,N_6856);
or U7323 (N_7323,N_6746,N_6906);
nor U7324 (N_7324,N_6587,N_6604);
nor U7325 (N_7325,N_6891,N_6562);
nand U7326 (N_7326,N_6873,N_6720);
nand U7327 (N_7327,N_6713,N_6702);
and U7328 (N_7328,N_6917,N_6703);
and U7329 (N_7329,N_6815,N_6510);
nor U7330 (N_7330,N_6554,N_6919);
or U7331 (N_7331,N_6573,N_6935);
xor U7332 (N_7332,N_6741,N_6855);
nand U7333 (N_7333,N_6615,N_6705);
nor U7334 (N_7334,N_6528,N_6553);
and U7335 (N_7335,N_6660,N_6537);
and U7336 (N_7336,N_6950,N_6867);
xor U7337 (N_7337,N_6721,N_6677);
xor U7338 (N_7338,N_6510,N_6782);
nor U7339 (N_7339,N_6722,N_6735);
xor U7340 (N_7340,N_6812,N_6610);
and U7341 (N_7341,N_6968,N_6768);
and U7342 (N_7342,N_6833,N_6770);
and U7343 (N_7343,N_6547,N_6788);
and U7344 (N_7344,N_6539,N_6925);
nand U7345 (N_7345,N_6966,N_6614);
or U7346 (N_7346,N_6864,N_6856);
nor U7347 (N_7347,N_6503,N_6518);
nor U7348 (N_7348,N_6737,N_6969);
and U7349 (N_7349,N_6826,N_6567);
or U7350 (N_7350,N_6985,N_6512);
nor U7351 (N_7351,N_6745,N_6548);
and U7352 (N_7352,N_6948,N_6790);
or U7353 (N_7353,N_6886,N_6639);
and U7354 (N_7354,N_6771,N_6602);
or U7355 (N_7355,N_6961,N_6626);
nand U7356 (N_7356,N_6591,N_6632);
and U7357 (N_7357,N_6944,N_6595);
nand U7358 (N_7358,N_6833,N_6976);
or U7359 (N_7359,N_6885,N_6878);
nand U7360 (N_7360,N_6646,N_6642);
or U7361 (N_7361,N_6981,N_6694);
and U7362 (N_7362,N_6683,N_6974);
nor U7363 (N_7363,N_6977,N_6596);
xnor U7364 (N_7364,N_6867,N_6602);
xor U7365 (N_7365,N_6791,N_6969);
nand U7366 (N_7366,N_6704,N_6984);
nor U7367 (N_7367,N_6690,N_6874);
nor U7368 (N_7368,N_6558,N_6771);
nor U7369 (N_7369,N_6718,N_6758);
xnor U7370 (N_7370,N_6515,N_6984);
nor U7371 (N_7371,N_6918,N_6662);
nor U7372 (N_7372,N_6704,N_6805);
or U7373 (N_7373,N_6927,N_6836);
or U7374 (N_7374,N_6690,N_6963);
nor U7375 (N_7375,N_6647,N_6590);
and U7376 (N_7376,N_6947,N_6529);
xor U7377 (N_7377,N_6950,N_6797);
nor U7378 (N_7378,N_6923,N_6927);
and U7379 (N_7379,N_6547,N_6693);
nand U7380 (N_7380,N_6782,N_6535);
and U7381 (N_7381,N_6500,N_6811);
or U7382 (N_7382,N_6604,N_6668);
and U7383 (N_7383,N_6976,N_6890);
nor U7384 (N_7384,N_6544,N_6637);
and U7385 (N_7385,N_6592,N_6539);
nand U7386 (N_7386,N_6814,N_6943);
nor U7387 (N_7387,N_6852,N_6984);
nor U7388 (N_7388,N_6767,N_6582);
or U7389 (N_7389,N_6606,N_6826);
nand U7390 (N_7390,N_6845,N_6707);
and U7391 (N_7391,N_6686,N_6714);
xnor U7392 (N_7392,N_6541,N_6833);
nor U7393 (N_7393,N_6757,N_6925);
xnor U7394 (N_7394,N_6601,N_6813);
xnor U7395 (N_7395,N_6548,N_6559);
nor U7396 (N_7396,N_6728,N_6971);
nand U7397 (N_7397,N_6762,N_6744);
nand U7398 (N_7398,N_6570,N_6975);
or U7399 (N_7399,N_6694,N_6978);
nand U7400 (N_7400,N_6846,N_6571);
nor U7401 (N_7401,N_6673,N_6509);
and U7402 (N_7402,N_6878,N_6859);
and U7403 (N_7403,N_6547,N_6958);
or U7404 (N_7404,N_6961,N_6923);
or U7405 (N_7405,N_6524,N_6546);
and U7406 (N_7406,N_6738,N_6804);
or U7407 (N_7407,N_6505,N_6941);
nand U7408 (N_7408,N_6973,N_6950);
nor U7409 (N_7409,N_6820,N_6548);
or U7410 (N_7410,N_6566,N_6885);
xnor U7411 (N_7411,N_6512,N_6796);
xor U7412 (N_7412,N_6956,N_6962);
nand U7413 (N_7413,N_6585,N_6665);
nor U7414 (N_7414,N_6873,N_6889);
xor U7415 (N_7415,N_6628,N_6964);
and U7416 (N_7416,N_6902,N_6888);
nand U7417 (N_7417,N_6569,N_6916);
xor U7418 (N_7418,N_6674,N_6841);
nor U7419 (N_7419,N_6557,N_6771);
nand U7420 (N_7420,N_6849,N_6740);
nand U7421 (N_7421,N_6509,N_6661);
and U7422 (N_7422,N_6963,N_6801);
nand U7423 (N_7423,N_6805,N_6946);
xnor U7424 (N_7424,N_6608,N_6640);
xnor U7425 (N_7425,N_6992,N_6998);
and U7426 (N_7426,N_6921,N_6923);
nor U7427 (N_7427,N_6551,N_6710);
nand U7428 (N_7428,N_6738,N_6571);
and U7429 (N_7429,N_6982,N_6520);
nor U7430 (N_7430,N_6805,N_6999);
nand U7431 (N_7431,N_6765,N_6612);
nor U7432 (N_7432,N_6971,N_6641);
xor U7433 (N_7433,N_6948,N_6859);
xor U7434 (N_7434,N_6914,N_6638);
nor U7435 (N_7435,N_6785,N_6517);
or U7436 (N_7436,N_6618,N_6586);
nor U7437 (N_7437,N_6649,N_6735);
nand U7438 (N_7438,N_6695,N_6550);
xnor U7439 (N_7439,N_6500,N_6982);
and U7440 (N_7440,N_6573,N_6703);
and U7441 (N_7441,N_6655,N_6789);
and U7442 (N_7442,N_6765,N_6760);
nand U7443 (N_7443,N_6542,N_6947);
and U7444 (N_7444,N_6519,N_6673);
or U7445 (N_7445,N_6904,N_6950);
xor U7446 (N_7446,N_6912,N_6858);
and U7447 (N_7447,N_6615,N_6546);
xnor U7448 (N_7448,N_6827,N_6996);
nand U7449 (N_7449,N_6608,N_6575);
xnor U7450 (N_7450,N_6969,N_6621);
nor U7451 (N_7451,N_6913,N_6650);
and U7452 (N_7452,N_6787,N_6523);
nand U7453 (N_7453,N_6913,N_6502);
and U7454 (N_7454,N_6537,N_6828);
xnor U7455 (N_7455,N_6832,N_6782);
or U7456 (N_7456,N_6976,N_6900);
and U7457 (N_7457,N_6561,N_6635);
and U7458 (N_7458,N_6985,N_6932);
nor U7459 (N_7459,N_6502,N_6936);
nand U7460 (N_7460,N_6693,N_6600);
xor U7461 (N_7461,N_6851,N_6989);
nor U7462 (N_7462,N_6598,N_6503);
xor U7463 (N_7463,N_6646,N_6686);
xor U7464 (N_7464,N_6583,N_6736);
xor U7465 (N_7465,N_6551,N_6574);
nor U7466 (N_7466,N_6593,N_6957);
or U7467 (N_7467,N_6509,N_6875);
and U7468 (N_7468,N_6781,N_6823);
nor U7469 (N_7469,N_6520,N_6685);
and U7470 (N_7470,N_6750,N_6759);
nor U7471 (N_7471,N_6715,N_6828);
xor U7472 (N_7472,N_6760,N_6520);
xor U7473 (N_7473,N_6978,N_6706);
and U7474 (N_7474,N_6799,N_6587);
nand U7475 (N_7475,N_6503,N_6696);
and U7476 (N_7476,N_6969,N_6806);
xor U7477 (N_7477,N_6649,N_6645);
nor U7478 (N_7478,N_6923,N_6566);
nor U7479 (N_7479,N_6681,N_6947);
nor U7480 (N_7480,N_6631,N_6870);
nor U7481 (N_7481,N_6960,N_6775);
xnor U7482 (N_7482,N_6928,N_6547);
or U7483 (N_7483,N_6706,N_6697);
and U7484 (N_7484,N_6810,N_6614);
and U7485 (N_7485,N_6954,N_6959);
and U7486 (N_7486,N_6911,N_6823);
and U7487 (N_7487,N_6782,N_6617);
or U7488 (N_7488,N_6647,N_6536);
nor U7489 (N_7489,N_6561,N_6944);
or U7490 (N_7490,N_6783,N_6930);
and U7491 (N_7491,N_6855,N_6886);
xor U7492 (N_7492,N_6564,N_6968);
nor U7493 (N_7493,N_6546,N_6668);
xnor U7494 (N_7494,N_6827,N_6980);
nand U7495 (N_7495,N_6737,N_6584);
xnor U7496 (N_7496,N_6677,N_6504);
nand U7497 (N_7497,N_6989,N_6604);
nor U7498 (N_7498,N_6834,N_6813);
nand U7499 (N_7499,N_6919,N_6982);
xnor U7500 (N_7500,N_7272,N_7122);
xnor U7501 (N_7501,N_7224,N_7025);
xnor U7502 (N_7502,N_7424,N_7046);
and U7503 (N_7503,N_7492,N_7363);
and U7504 (N_7504,N_7183,N_7069);
xnor U7505 (N_7505,N_7429,N_7368);
or U7506 (N_7506,N_7023,N_7418);
nor U7507 (N_7507,N_7433,N_7203);
or U7508 (N_7508,N_7177,N_7083);
or U7509 (N_7509,N_7485,N_7307);
nor U7510 (N_7510,N_7452,N_7048);
nor U7511 (N_7511,N_7073,N_7081);
nand U7512 (N_7512,N_7063,N_7490);
or U7513 (N_7513,N_7239,N_7487);
or U7514 (N_7514,N_7449,N_7134);
xnor U7515 (N_7515,N_7303,N_7341);
and U7516 (N_7516,N_7290,N_7060);
nor U7517 (N_7517,N_7446,N_7057);
or U7518 (N_7518,N_7343,N_7232);
nand U7519 (N_7519,N_7425,N_7310);
or U7520 (N_7520,N_7407,N_7188);
or U7521 (N_7521,N_7179,N_7067);
nor U7522 (N_7522,N_7215,N_7339);
and U7523 (N_7523,N_7037,N_7027);
nor U7524 (N_7524,N_7457,N_7047);
and U7525 (N_7525,N_7475,N_7022);
nor U7526 (N_7526,N_7344,N_7249);
or U7527 (N_7527,N_7152,N_7218);
nand U7528 (N_7528,N_7334,N_7128);
xor U7529 (N_7529,N_7171,N_7380);
xor U7530 (N_7530,N_7136,N_7143);
nor U7531 (N_7531,N_7039,N_7040);
and U7532 (N_7532,N_7328,N_7375);
and U7533 (N_7533,N_7358,N_7405);
xor U7534 (N_7534,N_7336,N_7021);
xor U7535 (N_7535,N_7116,N_7279);
and U7536 (N_7536,N_7453,N_7026);
nand U7537 (N_7537,N_7442,N_7350);
xnor U7538 (N_7538,N_7242,N_7496);
xnor U7539 (N_7539,N_7335,N_7052);
xnor U7540 (N_7540,N_7121,N_7056);
nor U7541 (N_7541,N_7031,N_7447);
and U7542 (N_7542,N_7379,N_7008);
nand U7543 (N_7543,N_7302,N_7278);
nor U7544 (N_7544,N_7337,N_7270);
xnor U7545 (N_7545,N_7119,N_7205);
or U7546 (N_7546,N_7109,N_7404);
nand U7547 (N_7547,N_7491,N_7186);
and U7548 (N_7548,N_7187,N_7062);
and U7549 (N_7549,N_7299,N_7364);
nand U7550 (N_7550,N_7480,N_7019);
xnor U7551 (N_7551,N_7080,N_7296);
xor U7552 (N_7552,N_7383,N_7311);
and U7553 (N_7553,N_7146,N_7172);
xor U7554 (N_7554,N_7414,N_7223);
nand U7555 (N_7555,N_7411,N_7243);
and U7556 (N_7556,N_7086,N_7118);
or U7557 (N_7557,N_7353,N_7458);
and U7558 (N_7558,N_7316,N_7061);
nand U7559 (N_7559,N_7427,N_7124);
or U7560 (N_7560,N_7200,N_7089);
and U7561 (N_7561,N_7402,N_7289);
nand U7562 (N_7562,N_7006,N_7182);
nand U7563 (N_7563,N_7126,N_7283);
or U7564 (N_7564,N_7013,N_7065);
xor U7565 (N_7565,N_7032,N_7180);
nand U7566 (N_7566,N_7245,N_7016);
nand U7567 (N_7567,N_7388,N_7276);
nand U7568 (N_7568,N_7269,N_7168);
nand U7569 (N_7569,N_7354,N_7413);
nor U7570 (N_7570,N_7438,N_7144);
nor U7571 (N_7571,N_7049,N_7162);
nor U7572 (N_7572,N_7390,N_7421);
and U7573 (N_7573,N_7064,N_7156);
nand U7574 (N_7574,N_7382,N_7036);
and U7575 (N_7575,N_7362,N_7185);
nand U7576 (N_7576,N_7478,N_7208);
xnor U7577 (N_7577,N_7415,N_7403);
xnor U7578 (N_7578,N_7422,N_7253);
or U7579 (N_7579,N_7158,N_7462);
and U7580 (N_7580,N_7135,N_7043);
and U7581 (N_7581,N_7288,N_7078);
nor U7582 (N_7582,N_7169,N_7197);
and U7583 (N_7583,N_7301,N_7266);
nor U7584 (N_7584,N_7199,N_7309);
and U7585 (N_7585,N_7014,N_7459);
nand U7586 (N_7586,N_7072,N_7314);
xnor U7587 (N_7587,N_7236,N_7366);
nor U7588 (N_7588,N_7099,N_7408);
or U7589 (N_7589,N_7294,N_7409);
xnor U7590 (N_7590,N_7356,N_7092);
nor U7591 (N_7591,N_7321,N_7317);
or U7592 (N_7592,N_7381,N_7389);
nor U7593 (N_7593,N_7258,N_7357);
and U7594 (N_7594,N_7004,N_7097);
and U7595 (N_7595,N_7175,N_7285);
or U7596 (N_7596,N_7167,N_7166);
nor U7597 (N_7597,N_7028,N_7035);
nand U7598 (N_7598,N_7011,N_7198);
nor U7599 (N_7599,N_7481,N_7050);
nand U7600 (N_7600,N_7479,N_7038);
xnor U7601 (N_7601,N_7472,N_7113);
nand U7602 (N_7602,N_7255,N_7140);
nand U7603 (N_7603,N_7160,N_7033);
and U7604 (N_7604,N_7306,N_7055);
or U7605 (N_7605,N_7385,N_7090);
or U7606 (N_7606,N_7286,N_7444);
or U7607 (N_7607,N_7318,N_7305);
or U7608 (N_7608,N_7466,N_7024);
and U7609 (N_7609,N_7178,N_7194);
or U7610 (N_7610,N_7149,N_7443);
nor U7611 (N_7611,N_7348,N_7018);
and U7612 (N_7612,N_7029,N_7320);
nand U7613 (N_7613,N_7088,N_7051);
nor U7614 (N_7614,N_7231,N_7191);
nor U7615 (N_7615,N_7387,N_7359);
nand U7616 (N_7616,N_7106,N_7114);
nand U7617 (N_7617,N_7094,N_7300);
xnor U7618 (N_7618,N_7132,N_7360);
xor U7619 (N_7619,N_7312,N_7184);
nor U7620 (N_7620,N_7399,N_7164);
and U7621 (N_7621,N_7133,N_7007);
and U7622 (N_7622,N_7082,N_7319);
nor U7623 (N_7623,N_7115,N_7495);
nand U7624 (N_7624,N_7228,N_7297);
or U7625 (N_7625,N_7325,N_7137);
and U7626 (N_7626,N_7391,N_7173);
xnor U7627 (N_7627,N_7202,N_7432);
or U7628 (N_7628,N_7315,N_7455);
nor U7629 (N_7629,N_7463,N_7304);
or U7630 (N_7630,N_7322,N_7281);
nor U7631 (N_7631,N_7210,N_7329);
nor U7632 (N_7632,N_7159,N_7298);
and U7633 (N_7633,N_7235,N_7079);
nand U7634 (N_7634,N_7486,N_7010);
nand U7635 (N_7635,N_7246,N_7112);
xor U7636 (N_7636,N_7476,N_7176);
nand U7637 (N_7637,N_7110,N_7257);
and U7638 (N_7638,N_7091,N_7274);
nor U7639 (N_7639,N_7410,N_7436);
nor U7640 (N_7640,N_7361,N_7423);
nand U7641 (N_7641,N_7141,N_7204);
nand U7642 (N_7642,N_7340,N_7251);
nor U7643 (N_7643,N_7244,N_7261);
or U7644 (N_7644,N_7398,N_7145);
nand U7645 (N_7645,N_7386,N_7372);
xnor U7646 (N_7646,N_7189,N_7003);
nor U7647 (N_7647,N_7001,N_7100);
nand U7648 (N_7648,N_7345,N_7127);
xnor U7649 (N_7649,N_7323,N_7488);
and U7650 (N_7650,N_7280,N_7397);
nor U7651 (N_7651,N_7256,N_7327);
nand U7652 (N_7652,N_7448,N_7005);
nor U7653 (N_7653,N_7221,N_7494);
nand U7654 (N_7654,N_7333,N_7434);
nor U7655 (N_7655,N_7464,N_7474);
xor U7656 (N_7656,N_7460,N_7170);
xor U7657 (N_7657,N_7401,N_7250);
xnor U7658 (N_7658,N_7222,N_7248);
or U7659 (N_7659,N_7220,N_7009);
or U7660 (N_7660,N_7017,N_7473);
nand U7661 (N_7661,N_7295,N_7234);
nand U7662 (N_7662,N_7441,N_7147);
nand U7663 (N_7663,N_7417,N_7428);
nand U7664 (N_7664,N_7497,N_7437);
nor U7665 (N_7665,N_7107,N_7431);
and U7666 (N_7666,N_7153,N_7493);
nand U7667 (N_7667,N_7015,N_7465);
nand U7668 (N_7668,N_7161,N_7454);
and U7669 (N_7669,N_7151,N_7045);
and U7670 (N_7670,N_7275,N_7111);
xor U7671 (N_7671,N_7267,N_7214);
nor U7672 (N_7672,N_7355,N_7277);
nand U7673 (N_7673,N_7477,N_7260);
nor U7674 (N_7674,N_7483,N_7207);
xor U7675 (N_7675,N_7247,N_7181);
xor U7676 (N_7676,N_7154,N_7347);
nor U7677 (N_7677,N_7393,N_7470);
and U7678 (N_7678,N_7456,N_7332);
and U7679 (N_7679,N_7252,N_7313);
nor U7680 (N_7680,N_7138,N_7211);
and U7681 (N_7681,N_7066,N_7201);
or U7682 (N_7682,N_7053,N_7482);
or U7683 (N_7683,N_7044,N_7209);
nor U7684 (N_7684,N_7471,N_7163);
nor U7685 (N_7685,N_7439,N_7042);
xnor U7686 (N_7686,N_7206,N_7440);
nor U7687 (N_7687,N_7216,N_7229);
nor U7688 (N_7688,N_7148,N_7367);
and U7689 (N_7689,N_7241,N_7058);
or U7690 (N_7690,N_7174,N_7030);
nor U7691 (N_7691,N_7284,N_7324);
and U7692 (N_7692,N_7461,N_7377);
nand U7693 (N_7693,N_7196,N_7219);
xor U7694 (N_7694,N_7282,N_7074);
or U7695 (N_7695,N_7095,N_7342);
and U7696 (N_7696,N_7416,N_7131);
or U7697 (N_7697,N_7371,N_7213);
or U7698 (N_7698,N_7435,N_7217);
nand U7699 (N_7699,N_7392,N_7394);
and U7700 (N_7700,N_7378,N_7130);
or U7701 (N_7701,N_7369,N_7263);
xor U7702 (N_7702,N_7426,N_7352);
nor U7703 (N_7703,N_7430,N_7308);
nor U7704 (N_7704,N_7139,N_7190);
or U7705 (N_7705,N_7000,N_7117);
and U7706 (N_7706,N_7268,N_7254);
xor U7707 (N_7707,N_7499,N_7212);
and U7708 (N_7708,N_7084,N_7076);
xor U7709 (N_7709,N_7230,N_7264);
nand U7710 (N_7710,N_7020,N_7104);
and U7711 (N_7711,N_7068,N_7384);
or U7712 (N_7712,N_7012,N_7075);
or U7713 (N_7713,N_7262,N_7396);
or U7714 (N_7714,N_7395,N_7225);
and U7715 (N_7715,N_7105,N_7484);
nand U7716 (N_7716,N_7059,N_7103);
nor U7717 (N_7717,N_7331,N_7259);
nand U7718 (N_7718,N_7098,N_7129);
and U7719 (N_7719,N_7101,N_7346);
xor U7720 (N_7720,N_7226,N_7293);
nand U7721 (N_7721,N_7291,N_7451);
nor U7722 (N_7722,N_7265,N_7227);
and U7723 (N_7723,N_7498,N_7338);
nand U7724 (N_7724,N_7237,N_7150);
or U7725 (N_7725,N_7412,N_7071);
and U7726 (N_7726,N_7108,N_7271);
xor U7727 (N_7727,N_7420,N_7193);
xor U7728 (N_7728,N_7374,N_7287);
xnor U7729 (N_7729,N_7400,N_7351);
or U7730 (N_7730,N_7233,N_7155);
and U7731 (N_7731,N_7165,N_7087);
and U7732 (N_7732,N_7467,N_7376);
nor U7733 (N_7733,N_7489,N_7370);
nor U7734 (N_7734,N_7034,N_7373);
nand U7735 (N_7735,N_7093,N_7273);
xnor U7736 (N_7736,N_7041,N_7330);
and U7737 (N_7737,N_7070,N_7102);
and U7738 (N_7738,N_7292,N_7468);
nor U7739 (N_7739,N_7419,N_7445);
or U7740 (N_7740,N_7406,N_7195);
and U7741 (N_7741,N_7142,N_7123);
and U7742 (N_7742,N_7469,N_7349);
or U7743 (N_7743,N_7002,N_7120);
xor U7744 (N_7744,N_7365,N_7096);
nor U7745 (N_7745,N_7192,N_7077);
or U7746 (N_7746,N_7326,N_7240);
nand U7747 (N_7747,N_7238,N_7125);
xnor U7748 (N_7748,N_7054,N_7450);
nand U7749 (N_7749,N_7157,N_7085);
nand U7750 (N_7750,N_7158,N_7145);
nor U7751 (N_7751,N_7337,N_7167);
xor U7752 (N_7752,N_7418,N_7260);
or U7753 (N_7753,N_7363,N_7431);
and U7754 (N_7754,N_7147,N_7436);
nor U7755 (N_7755,N_7370,N_7303);
nand U7756 (N_7756,N_7094,N_7439);
nand U7757 (N_7757,N_7073,N_7385);
nand U7758 (N_7758,N_7042,N_7172);
or U7759 (N_7759,N_7437,N_7106);
xnor U7760 (N_7760,N_7126,N_7350);
or U7761 (N_7761,N_7434,N_7170);
xor U7762 (N_7762,N_7132,N_7331);
nand U7763 (N_7763,N_7100,N_7053);
or U7764 (N_7764,N_7381,N_7476);
and U7765 (N_7765,N_7127,N_7280);
xor U7766 (N_7766,N_7155,N_7283);
xor U7767 (N_7767,N_7047,N_7195);
xnor U7768 (N_7768,N_7322,N_7050);
nand U7769 (N_7769,N_7349,N_7023);
nand U7770 (N_7770,N_7398,N_7140);
nor U7771 (N_7771,N_7157,N_7290);
and U7772 (N_7772,N_7468,N_7077);
nand U7773 (N_7773,N_7343,N_7060);
and U7774 (N_7774,N_7034,N_7412);
xnor U7775 (N_7775,N_7177,N_7188);
nor U7776 (N_7776,N_7371,N_7355);
nand U7777 (N_7777,N_7295,N_7035);
nand U7778 (N_7778,N_7341,N_7368);
and U7779 (N_7779,N_7364,N_7297);
or U7780 (N_7780,N_7089,N_7002);
xnor U7781 (N_7781,N_7428,N_7086);
or U7782 (N_7782,N_7154,N_7367);
xnor U7783 (N_7783,N_7028,N_7358);
nor U7784 (N_7784,N_7166,N_7233);
nor U7785 (N_7785,N_7414,N_7024);
and U7786 (N_7786,N_7004,N_7357);
nor U7787 (N_7787,N_7077,N_7080);
and U7788 (N_7788,N_7322,N_7300);
xnor U7789 (N_7789,N_7138,N_7278);
xnor U7790 (N_7790,N_7415,N_7360);
or U7791 (N_7791,N_7353,N_7130);
xnor U7792 (N_7792,N_7008,N_7479);
and U7793 (N_7793,N_7146,N_7413);
nor U7794 (N_7794,N_7150,N_7262);
and U7795 (N_7795,N_7071,N_7072);
or U7796 (N_7796,N_7077,N_7385);
or U7797 (N_7797,N_7459,N_7211);
nand U7798 (N_7798,N_7435,N_7133);
or U7799 (N_7799,N_7234,N_7182);
nor U7800 (N_7800,N_7374,N_7090);
and U7801 (N_7801,N_7424,N_7377);
nand U7802 (N_7802,N_7422,N_7202);
nand U7803 (N_7803,N_7255,N_7415);
nand U7804 (N_7804,N_7113,N_7420);
and U7805 (N_7805,N_7242,N_7362);
nand U7806 (N_7806,N_7164,N_7482);
nor U7807 (N_7807,N_7311,N_7357);
xnor U7808 (N_7808,N_7040,N_7265);
nand U7809 (N_7809,N_7324,N_7074);
xnor U7810 (N_7810,N_7223,N_7292);
nor U7811 (N_7811,N_7131,N_7346);
and U7812 (N_7812,N_7188,N_7467);
and U7813 (N_7813,N_7008,N_7320);
nor U7814 (N_7814,N_7180,N_7387);
nor U7815 (N_7815,N_7293,N_7232);
or U7816 (N_7816,N_7056,N_7301);
xor U7817 (N_7817,N_7454,N_7118);
and U7818 (N_7818,N_7168,N_7132);
nor U7819 (N_7819,N_7457,N_7482);
nor U7820 (N_7820,N_7052,N_7429);
nand U7821 (N_7821,N_7487,N_7201);
xor U7822 (N_7822,N_7046,N_7364);
nor U7823 (N_7823,N_7120,N_7315);
or U7824 (N_7824,N_7079,N_7041);
xor U7825 (N_7825,N_7072,N_7225);
nand U7826 (N_7826,N_7002,N_7118);
and U7827 (N_7827,N_7261,N_7164);
nor U7828 (N_7828,N_7180,N_7308);
and U7829 (N_7829,N_7087,N_7214);
or U7830 (N_7830,N_7213,N_7338);
or U7831 (N_7831,N_7279,N_7133);
xor U7832 (N_7832,N_7351,N_7158);
nand U7833 (N_7833,N_7342,N_7301);
or U7834 (N_7834,N_7443,N_7089);
nand U7835 (N_7835,N_7368,N_7391);
xnor U7836 (N_7836,N_7344,N_7276);
and U7837 (N_7837,N_7415,N_7389);
xnor U7838 (N_7838,N_7246,N_7277);
xor U7839 (N_7839,N_7455,N_7233);
xnor U7840 (N_7840,N_7291,N_7061);
or U7841 (N_7841,N_7371,N_7211);
or U7842 (N_7842,N_7098,N_7491);
and U7843 (N_7843,N_7196,N_7026);
or U7844 (N_7844,N_7442,N_7370);
and U7845 (N_7845,N_7035,N_7019);
and U7846 (N_7846,N_7215,N_7285);
nand U7847 (N_7847,N_7443,N_7420);
and U7848 (N_7848,N_7133,N_7205);
or U7849 (N_7849,N_7041,N_7142);
or U7850 (N_7850,N_7355,N_7489);
nor U7851 (N_7851,N_7214,N_7289);
nor U7852 (N_7852,N_7420,N_7038);
nand U7853 (N_7853,N_7372,N_7057);
nand U7854 (N_7854,N_7244,N_7328);
nor U7855 (N_7855,N_7040,N_7256);
nor U7856 (N_7856,N_7016,N_7344);
nand U7857 (N_7857,N_7035,N_7248);
xnor U7858 (N_7858,N_7340,N_7296);
and U7859 (N_7859,N_7417,N_7322);
nand U7860 (N_7860,N_7413,N_7322);
xnor U7861 (N_7861,N_7347,N_7355);
nand U7862 (N_7862,N_7332,N_7162);
nand U7863 (N_7863,N_7308,N_7314);
and U7864 (N_7864,N_7403,N_7480);
and U7865 (N_7865,N_7027,N_7474);
and U7866 (N_7866,N_7460,N_7426);
xor U7867 (N_7867,N_7000,N_7312);
and U7868 (N_7868,N_7411,N_7280);
nand U7869 (N_7869,N_7274,N_7033);
or U7870 (N_7870,N_7261,N_7369);
nor U7871 (N_7871,N_7008,N_7053);
xnor U7872 (N_7872,N_7262,N_7450);
nand U7873 (N_7873,N_7177,N_7131);
nand U7874 (N_7874,N_7473,N_7024);
or U7875 (N_7875,N_7093,N_7110);
nand U7876 (N_7876,N_7436,N_7418);
xor U7877 (N_7877,N_7389,N_7206);
nor U7878 (N_7878,N_7416,N_7173);
and U7879 (N_7879,N_7087,N_7251);
nand U7880 (N_7880,N_7087,N_7478);
nand U7881 (N_7881,N_7290,N_7224);
or U7882 (N_7882,N_7386,N_7037);
nand U7883 (N_7883,N_7404,N_7374);
and U7884 (N_7884,N_7477,N_7305);
nand U7885 (N_7885,N_7175,N_7274);
nand U7886 (N_7886,N_7377,N_7473);
xnor U7887 (N_7887,N_7166,N_7087);
xor U7888 (N_7888,N_7224,N_7483);
and U7889 (N_7889,N_7331,N_7151);
nor U7890 (N_7890,N_7432,N_7146);
or U7891 (N_7891,N_7261,N_7340);
or U7892 (N_7892,N_7328,N_7202);
xnor U7893 (N_7893,N_7406,N_7385);
nor U7894 (N_7894,N_7470,N_7336);
nor U7895 (N_7895,N_7488,N_7418);
and U7896 (N_7896,N_7123,N_7236);
xor U7897 (N_7897,N_7186,N_7158);
and U7898 (N_7898,N_7486,N_7122);
and U7899 (N_7899,N_7320,N_7083);
or U7900 (N_7900,N_7119,N_7424);
xnor U7901 (N_7901,N_7130,N_7305);
nand U7902 (N_7902,N_7398,N_7192);
nor U7903 (N_7903,N_7048,N_7360);
nor U7904 (N_7904,N_7243,N_7066);
nor U7905 (N_7905,N_7213,N_7392);
nand U7906 (N_7906,N_7259,N_7467);
xor U7907 (N_7907,N_7260,N_7144);
and U7908 (N_7908,N_7304,N_7174);
or U7909 (N_7909,N_7033,N_7043);
nor U7910 (N_7910,N_7302,N_7320);
xor U7911 (N_7911,N_7415,N_7449);
nor U7912 (N_7912,N_7160,N_7276);
nor U7913 (N_7913,N_7101,N_7416);
xnor U7914 (N_7914,N_7421,N_7366);
and U7915 (N_7915,N_7491,N_7358);
or U7916 (N_7916,N_7445,N_7015);
or U7917 (N_7917,N_7369,N_7052);
nand U7918 (N_7918,N_7369,N_7143);
nand U7919 (N_7919,N_7440,N_7460);
xor U7920 (N_7920,N_7358,N_7336);
and U7921 (N_7921,N_7369,N_7203);
nor U7922 (N_7922,N_7210,N_7295);
nor U7923 (N_7923,N_7400,N_7323);
or U7924 (N_7924,N_7075,N_7068);
and U7925 (N_7925,N_7481,N_7134);
or U7926 (N_7926,N_7325,N_7032);
or U7927 (N_7927,N_7427,N_7069);
or U7928 (N_7928,N_7030,N_7102);
and U7929 (N_7929,N_7136,N_7016);
nand U7930 (N_7930,N_7067,N_7071);
nor U7931 (N_7931,N_7070,N_7403);
xor U7932 (N_7932,N_7249,N_7037);
or U7933 (N_7933,N_7059,N_7372);
xnor U7934 (N_7934,N_7213,N_7287);
or U7935 (N_7935,N_7008,N_7036);
xor U7936 (N_7936,N_7239,N_7037);
nand U7937 (N_7937,N_7366,N_7275);
and U7938 (N_7938,N_7078,N_7264);
xor U7939 (N_7939,N_7245,N_7060);
nor U7940 (N_7940,N_7447,N_7197);
and U7941 (N_7941,N_7349,N_7336);
and U7942 (N_7942,N_7172,N_7350);
or U7943 (N_7943,N_7100,N_7196);
and U7944 (N_7944,N_7143,N_7444);
and U7945 (N_7945,N_7159,N_7474);
nor U7946 (N_7946,N_7030,N_7074);
or U7947 (N_7947,N_7144,N_7053);
nand U7948 (N_7948,N_7138,N_7075);
xor U7949 (N_7949,N_7486,N_7487);
nor U7950 (N_7950,N_7092,N_7334);
nand U7951 (N_7951,N_7065,N_7185);
or U7952 (N_7952,N_7012,N_7400);
xnor U7953 (N_7953,N_7172,N_7107);
xor U7954 (N_7954,N_7247,N_7332);
xnor U7955 (N_7955,N_7128,N_7001);
xor U7956 (N_7956,N_7423,N_7246);
xnor U7957 (N_7957,N_7375,N_7159);
and U7958 (N_7958,N_7466,N_7121);
nor U7959 (N_7959,N_7227,N_7448);
nand U7960 (N_7960,N_7458,N_7442);
and U7961 (N_7961,N_7193,N_7125);
nand U7962 (N_7962,N_7124,N_7077);
nand U7963 (N_7963,N_7387,N_7417);
xnor U7964 (N_7964,N_7446,N_7340);
nand U7965 (N_7965,N_7110,N_7441);
nor U7966 (N_7966,N_7205,N_7251);
and U7967 (N_7967,N_7189,N_7302);
and U7968 (N_7968,N_7377,N_7212);
nand U7969 (N_7969,N_7402,N_7133);
and U7970 (N_7970,N_7181,N_7251);
and U7971 (N_7971,N_7158,N_7405);
xor U7972 (N_7972,N_7289,N_7436);
or U7973 (N_7973,N_7098,N_7133);
nor U7974 (N_7974,N_7229,N_7414);
xnor U7975 (N_7975,N_7396,N_7146);
or U7976 (N_7976,N_7033,N_7161);
nor U7977 (N_7977,N_7304,N_7162);
nor U7978 (N_7978,N_7475,N_7028);
nor U7979 (N_7979,N_7436,N_7391);
nand U7980 (N_7980,N_7254,N_7485);
or U7981 (N_7981,N_7151,N_7473);
nand U7982 (N_7982,N_7111,N_7440);
xor U7983 (N_7983,N_7464,N_7092);
and U7984 (N_7984,N_7469,N_7299);
nor U7985 (N_7985,N_7193,N_7214);
xnor U7986 (N_7986,N_7078,N_7102);
nor U7987 (N_7987,N_7405,N_7283);
nor U7988 (N_7988,N_7191,N_7492);
or U7989 (N_7989,N_7077,N_7026);
nor U7990 (N_7990,N_7115,N_7153);
xor U7991 (N_7991,N_7402,N_7042);
xor U7992 (N_7992,N_7490,N_7268);
and U7993 (N_7993,N_7482,N_7121);
and U7994 (N_7994,N_7211,N_7486);
nor U7995 (N_7995,N_7328,N_7262);
and U7996 (N_7996,N_7259,N_7027);
or U7997 (N_7997,N_7029,N_7146);
nand U7998 (N_7998,N_7445,N_7498);
or U7999 (N_7999,N_7193,N_7286);
and U8000 (N_8000,N_7642,N_7895);
nand U8001 (N_8001,N_7953,N_7977);
nor U8002 (N_8002,N_7849,N_7587);
nand U8003 (N_8003,N_7767,N_7865);
nand U8004 (N_8004,N_7829,N_7777);
and U8005 (N_8005,N_7984,N_7721);
and U8006 (N_8006,N_7556,N_7923);
nand U8007 (N_8007,N_7745,N_7943);
xor U8008 (N_8008,N_7728,N_7706);
and U8009 (N_8009,N_7527,N_7627);
or U8010 (N_8010,N_7911,N_7744);
nand U8011 (N_8011,N_7680,N_7988);
nor U8012 (N_8012,N_7960,N_7586);
xnor U8013 (N_8013,N_7947,N_7872);
nor U8014 (N_8014,N_7776,N_7864);
nor U8015 (N_8015,N_7521,N_7726);
and U8016 (N_8016,N_7775,N_7717);
nor U8017 (N_8017,N_7814,N_7522);
nor U8018 (N_8018,N_7863,N_7945);
and U8019 (N_8019,N_7770,N_7533);
or U8020 (N_8020,N_7779,N_7672);
and U8021 (N_8021,N_7553,N_7557);
nand U8022 (N_8022,N_7646,N_7795);
nor U8023 (N_8023,N_7545,N_7564);
nand U8024 (N_8024,N_7641,N_7724);
or U8025 (N_8025,N_7520,N_7749);
xor U8026 (N_8026,N_7707,N_7825);
or U8027 (N_8027,N_7831,N_7824);
nor U8028 (N_8028,N_7759,N_7946);
xor U8029 (N_8029,N_7854,N_7568);
and U8030 (N_8030,N_7678,N_7720);
xor U8031 (N_8031,N_7866,N_7659);
nor U8032 (N_8032,N_7915,N_7789);
nand U8033 (N_8033,N_7700,N_7651);
or U8034 (N_8034,N_7692,N_7752);
or U8035 (N_8035,N_7772,N_7763);
xnor U8036 (N_8036,N_7559,N_7929);
or U8037 (N_8037,N_7903,N_7631);
nand U8038 (N_8038,N_7882,N_7912);
xor U8039 (N_8039,N_7990,N_7666);
xor U8040 (N_8040,N_7738,N_7755);
and U8041 (N_8041,N_7529,N_7561);
nor U8042 (N_8042,N_7937,N_7810);
nor U8043 (N_8043,N_7518,N_7832);
xnor U8044 (N_8044,N_7676,N_7590);
nor U8045 (N_8045,N_7602,N_7858);
or U8046 (N_8046,N_7699,N_7819);
nand U8047 (N_8047,N_7512,N_7917);
xnor U8048 (N_8048,N_7927,N_7565);
nand U8049 (N_8049,N_7563,N_7570);
or U8050 (N_8050,N_7743,N_7806);
nor U8051 (N_8051,N_7616,N_7993);
and U8052 (N_8052,N_7665,N_7804);
or U8053 (N_8053,N_7836,N_7941);
and U8054 (N_8054,N_7530,N_7841);
xor U8055 (N_8055,N_7628,N_7940);
or U8056 (N_8056,N_7867,N_7809);
xor U8057 (N_8057,N_7588,N_7820);
and U8058 (N_8058,N_7883,N_7515);
or U8059 (N_8059,N_7595,N_7732);
and U8060 (N_8060,N_7690,N_7861);
xor U8061 (N_8061,N_7753,N_7975);
nor U8062 (N_8062,N_7905,N_7794);
nand U8063 (N_8063,N_7509,N_7736);
xnor U8064 (N_8064,N_7837,N_7935);
and U8065 (N_8065,N_7904,N_7856);
nor U8066 (N_8066,N_7723,N_7902);
xor U8067 (N_8067,N_7609,N_7981);
and U8068 (N_8068,N_7955,N_7938);
nor U8069 (N_8069,N_7843,N_7514);
xnor U8070 (N_8070,N_7971,N_7839);
xor U8071 (N_8071,N_7624,N_7962);
nor U8072 (N_8072,N_7754,N_7765);
nor U8073 (N_8073,N_7661,N_7950);
nor U8074 (N_8074,N_7782,N_7932);
nand U8075 (N_8075,N_7899,N_7870);
xnor U8076 (N_8076,N_7722,N_7735);
xor U8077 (N_8077,N_7517,N_7614);
and U8078 (N_8078,N_7599,N_7606);
nand U8079 (N_8079,N_7705,N_7931);
and U8080 (N_8080,N_7584,N_7756);
and U8081 (N_8081,N_7890,N_7818);
nand U8082 (N_8082,N_7800,N_7604);
or U8083 (N_8083,N_7936,N_7897);
and U8084 (N_8084,N_7833,N_7539);
or U8085 (N_8085,N_7996,N_7970);
nand U8086 (N_8086,N_7852,N_7597);
or U8087 (N_8087,N_7558,N_7944);
or U8088 (N_8088,N_7611,N_7501);
nor U8089 (N_8089,N_7774,N_7876);
xnor U8090 (N_8090,N_7761,N_7875);
and U8091 (N_8091,N_7739,N_7859);
or U8092 (N_8092,N_7928,N_7808);
or U8093 (N_8093,N_7812,N_7516);
nand U8094 (N_8094,N_7693,N_7796);
xor U8095 (N_8095,N_7914,N_7788);
and U8096 (N_8096,N_7834,N_7653);
or U8097 (N_8097,N_7551,N_7654);
and U8098 (N_8098,N_7942,N_7815);
nand U8099 (N_8099,N_7908,N_7964);
nand U8100 (N_8100,N_7891,N_7910);
nor U8101 (N_8101,N_7510,N_7688);
nor U8102 (N_8102,N_7648,N_7827);
nor U8103 (N_8103,N_7741,N_7828);
nor U8104 (N_8104,N_7918,N_7650);
nor U8105 (N_8105,N_7538,N_7543);
nor U8106 (N_8106,N_7956,N_7781);
or U8107 (N_8107,N_7885,N_7888);
xor U8108 (N_8108,N_7546,N_7685);
nor U8109 (N_8109,N_7513,N_7746);
nand U8110 (N_8110,N_7764,N_7773);
or U8111 (N_8111,N_7845,N_7500);
nand U8112 (N_8112,N_7901,N_7507);
nand U8113 (N_8113,N_7686,N_7822);
or U8114 (N_8114,N_7673,N_7985);
and U8115 (N_8115,N_7725,N_7961);
xor U8116 (N_8116,N_7695,N_7647);
and U8117 (N_8117,N_7835,N_7670);
and U8118 (N_8118,N_7667,N_7934);
nand U8119 (N_8119,N_7634,N_7737);
xor U8120 (N_8120,N_7889,N_7992);
nand U8121 (N_8121,N_7589,N_7525);
xor U8122 (N_8122,N_7655,N_7807);
nand U8123 (N_8123,N_7535,N_7608);
nor U8124 (N_8124,N_7913,N_7892);
or U8125 (N_8125,N_7880,N_7508);
or U8126 (N_8126,N_7731,N_7592);
nand U8127 (N_8127,N_7537,N_7662);
or U8128 (N_8128,N_7848,N_7550);
or U8129 (N_8129,N_7689,N_7577);
xor U8130 (N_8130,N_7881,N_7817);
xnor U8131 (N_8131,N_7771,N_7768);
nand U8132 (N_8132,N_7747,N_7844);
nor U8133 (N_8133,N_7846,N_7930);
or U8134 (N_8134,N_7979,N_7709);
xnor U8135 (N_8135,N_7760,N_7573);
nor U8136 (N_8136,N_7734,N_7994);
and U8137 (N_8137,N_7612,N_7860);
or U8138 (N_8138,N_7886,N_7907);
nand U8139 (N_8139,N_7579,N_7694);
and U8140 (N_8140,N_7511,N_7583);
nand U8141 (N_8141,N_7951,N_7920);
and U8142 (N_8142,N_7571,N_7811);
nor U8143 (N_8143,N_7711,N_7610);
and U8144 (N_8144,N_7969,N_7791);
nor U8145 (N_8145,N_7790,N_7842);
nor U8146 (N_8146,N_7894,N_7963);
or U8147 (N_8147,N_7742,N_7576);
nand U8148 (N_8148,N_7900,N_7548);
nand U8149 (N_8149,N_7757,N_7851);
and U8150 (N_8150,N_7729,N_7593);
xor U8151 (N_8151,N_7585,N_7813);
or U8152 (N_8152,N_7504,N_7799);
or U8153 (N_8153,N_7919,N_7884);
nand U8154 (N_8154,N_7629,N_7893);
xnor U8155 (N_8155,N_7633,N_7823);
and U8156 (N_8156,N_7998,N_7959);
nor U8157 (N_8157,N_7600,N_7976);
nand U8158 (N_8158,N_7965,N_7869);
and U8159 (N_8159,N_7862,N_7974);
and U8160 (N_8160,N_7803,N_7784);
or U8161 (N_8161,N_7658,N_7640);
nor U8162 (N_8162,N_7802,N_7926);
or U8163 (N_8163,N_7536,N_7618);
nand U8164 (N_8164,N_7778,N_7555);
nor U8165 (N_8165,N_7544,N_7909);
xnor U8166 (N_8166,N_7523,N_7615);
nand U8167 (N_8167,N_7540,N_7704);
or U8168 (N_8168,N_7668,N_7581);
xnor U8169 (N_8169,N_7687,N_7838);
nor U8170 (N_8170,N_7531,N_7855);
nand U8171 (N_8171,N_7560,N_7986);
or U8172 (N_8172,N_7552,N_7991);
nor U8173 (N_8173,N_7797,N_7980);
xnor U8174 (N_8174,N_7780,N_7978);
or U8175 (N_8175,N_7503,N_7878);
xnor U8176 (N_8176,N_7574,N_7997);
nor U8177 (N_8177,N_7957,N_7715);
xor U8178 (N_8178,N_7973,N_7671);
nor U8179 (N_8179,N_7649,N_7566);
xnor U8180 (N_8180,N_7758,N_7830);
or U8181 (N_8181,N_7632,N_7983);
xor U8182 (N_8182,N_7675,N_7591);
nor U8183 (N_8183,N_7626,N_7684);
or U8184 (N_8184,N_7598,N_7718);
nor U8185 (N_8185,N_7657,N_7643);
xor U8186 (N_8186,N_7798,N_7816);
or U8187 (N_8187,N_7982,N_7625);
or U8188 (N_8188,N_7989,N_7948);
nand U8189 (N_8189,N_7664,N_7580);
or U8190 (N_8190,N_7748,N_7645);
nor U8191 (N_8191,N_7766,N_7644);
nand U8192 (N_8192,N_7541,N_7528);
and U8193 (N_8193,N_7638,N_7669);
nor U8194 (N_8194,N_7683,N_7871);
and U8195 (N_8195,N_7712,N_7605);
nand U8196 (N_8196,N_7787,N_7639);
or U8197 (N_8197,N_7708,N_7534);
or U8198 (N_8198,N_7792,N_7847);
nand U8199 (N_8199,N_7906,N_7575);
xor U8200 (N_8200,N_7542,N_7569);
and U8201 (N_8201,N_7702,N_7750);
nand U8202 (N_8202,N_7554,N_7594);
and U8203 (N_8203,N_7630,N_7506);
nand U8204 (N_8204,N_7623,N_7519);
or U8205 (N_8205,N_7727,N_7968);
xnor U8206 (N_8206,N_7660,N_7730);
and U8207 (N_8207,N_7873,N_7887);
and U8208 (N_8208,N_7691,N_7896);
nand U8209 (N_8209,N_7879,N_7572);
or U8210 (N_8210,N_7682,N_7696);
and U8211 (N_8211,N_7697,N_7769);
nor U8212 (N_8212,N_7898,N_7603);
xnor U8213 (N_8213,N_7698,N_7674);
xor U8214 (N_8214,N_7578,N_7958);
nor U8215 (N_8215,N_7621,N_7713);
xnor U8216 (N_8216,N_7617,N_7733);
or U8217 (N_8217,N_7762,N_7677);
and U8218 (N_8218,N_7567,N_7916);
nor U8219 (N_8219,N_7877,N_7656);
and U8220 (N_8220,N_7719,N_7853);
nor U8221 (N_8221,N_7972,N_7995);
xor U8222 (N_8222,N_7826,N_7987);
nand U8223 (N_8223,N_7922,N_7524);
or U8224 (N_8224,N_7714,N_7663);
or U8225 (N_8225,N_7954,N_7751);
nor U8226 (N_8226,N_7966,N_7549);
nand U8227 (N_8227,N_7786,N_7582);
nand U8228 (N_8228,N_7681,N_7939);
or U8229 (N_8229,N_7933,N_7840);
xor U8230 (N_8230,N_7636,N_7703);
and U8231 (N_8231,N_7793,N_7857);
or U8232 (N_8232,N_7679,N_7620);
nand U8233 (N_8233,N_7740,N_7925);
nand U8234 (N_8234,N_7502,N_7547);
or U8235 (N_8235,N_7783,N_7505);
xnor U8236 (N_8236,N_7924,N_7635);
nand U8237 (N_8237,N_7607,N_7601);
or U8238 (N_8238,N_7952,N_7949);
and U8239 (N_8239,N_7619,N_7868);
and U8240 (N_8240,N_7874,N_7562);
nor U8241 (N_8241,N_7532,N_7526);
xnor U8242 (N_8242,N_7967,N_7701);
nor U8243 (N_8243,N_7716,N_7785);
and U8244 (N_8244,N_7596,N_7622);
or U8245 (N_8245,N_7652,N_7999);
nor U8246 (N_8246,N_7850,N_7921);
and U8247 (N_8247,N_7805,N_7637);
nand U8248 (N_8248,N_7710,N_7821);
nand U8249 (N_8249,N_7801,N_7613);
or U8250 (N_8250,N_7804,N_7670);
and U8251 (N_8251,N_7916,N_7672);
nor U8252 (N_8252,N_7705,N_7792);
or U8253 (N_8253,N_7848,N_7796);
or U8254 (N_8254,N_7803,N_7507);
and U8255 (N_8255,N_7968,N_7588);
and U8256 (N_8256,N_7801,N_7920);
xnor U8257 (N_8257,N_7883,N_7526);
or U8258 (N_8258,N_7772,N_7592);
nand U8259 (N_8259,N_7831,N_7906);
xor U8260 (N_8260,N_7971,N_7855);
and U8261 (N_8261,N_7865,N_7884);
or U8262 (N_8262,N_7840,N_7946);
and U8263 (N_8263,N_7573,N_7506);
nand U8264 (N_8264,N_7936,N_7817);
or U8265 (N_8265,N_7938,N_7581);
and U8266 (N_8266,N_7851,N_7788);
or U8267 (N_8267,N_7774,N_7669);
nand U8268 (N_8268,N_7792,N_7584);
or U8269 (N_8269,N_7927,N_7617);
nand U8270 (N_8270,N_7806,N_7592);
nand U8271 (N_8271,N_7949,N_7790);
or U8272 (N_8272,N_7662,N_7569);
or U8273 (N_8273,N_7825,N_7720);
nand U8274 (N_8274,N_7897,N_7952);
nand U8275 (N_8275,N_7755,N_7914);
nor U8276 (N_8276,N_7887,N_7715);
and U8277 (N_8277,N_7888,N_7687);
and U8278 (N_8278,N_7894,N_7998);
nand U8279 (N_8279,N_7521,N_7612);
nand U8280 (N_8280,N_7901,N_7985);
xor U8281 (N_8281,N_7621,N_7946);
xnor U8282 (N_8282,N_7922,N_7727);
xnor U8283 (N_8283,N_7829,N_7611);
xor U8284 (N_8284,N_7874,N_7552);
and U8285 (N_8285,N_7733,N_7532);
nor U8286 (N_8286,N_7813,N_7982);
nand U8287 (N_8287,N_7912,N_7969);
nor U8288 (N_8288,N_7978,N_7598);
or U8289 (N_8289,N_7641,N_7924);
and U8290 (N_8290,N_7520,N_7615);
and U8291 (N_8291,N_7939,N_7782);
nor U8292 (N_8292,N_7664,N_7615);
or U8293 (N_8293,N_7942,N_7952);
and U8294 (N_8294,N_7651,N_7574);
nand U8295 (N_8295,N_7556,N_7930);
or U8296 (N_8296,N_7580,N_7525);
and U8297 (N_8297,N_7780,N_7938);
and U8298 (N_8298,N_7522,N_7947);
and U8299 (N_8299,N_7980,N_7650);
nand U8300 (N_8300,N_7913,N_7920);
xnor U8301 (N_8301,N_7900,N_7906);
nor U8302 (N_8302,N_7763,N_7875);
or U8303 (N_8303,N_7532,N_7903);
nand U8304 (N_8304,N_7814,N_7975);
xnor U8305 (N_8305,N_7805,N_7718);
nand U8306 (N_8306,N_7679,N_7851);
and U8307 (N_8307,N_7951,N_7730);
xnor U8308 (N_8308,N_7905,N_7670);
and U8309 (N_8309,N_7773,N_7668);
nor U8310 (N_8310,N_7620,N_7898);
and U8311 (N_8311,N_7510,N_7588);
or U8312 (N_8312,N_7676,N_7882);
xnor U8313 (N_8313,N_7825,N_7605);
nor U8314 (N_8314,N_7751,N_7710);
or U8315 (N_8315,N_7905,N_7518);
and U8316 (N_8316,N_7584,N_7668);
and U8317 (N_8317,N_7759,N_7587);
and U8318 (N_8318,N_7812,N_7994);
xor U8319 (N_8319,N_7988,N_7696);
or U8320 (N_8320,N_7723,N_7634);
nor U8321 (N_8321,N_7877,N_7903);
and U8322 (N_8322,N_7853,N_7637);
or U8323 (N_8323,N_7980,N_7603);
nand U8324 (N_8324,N_7579,N_7722);
nand U8325 (N_8325,N_7931,N_7963);
nor U8326 (N_8326,N_7872,N_7957);
or U8327 (N_8327,N_7686,N_7512);
and U8328 (N_8328,N_7919,N_7524);
nand U8329 (N_8329,N_7560,N_7859);
and U8330 (N_8330,N_7789,N_7853);
nand U8331 (N_8331,N_7637,N_7768);
xnor U8332 (N_8332,N_7984,N_7933);
nor U8333 (N_8333,N_7548,N_7726);
or U8334 (N_8334,N_7953,N_7955);
xor U8335 (N_8335,N_7615,N_7695);
nand U8336 (N_8336,N_7803,N_7903);
nor U8337 (N_8337,N_7719,N_7735);
nor U8338 (N_8338,N_7949,N_7992);
xor U8339 (N_8339,N_7749,N_7527);
or U8340 (N_8340,N_7691,N_7669);
and U8341 (N_8341,N_7590,N_7566);
nand U8342 (N_8342,N_7574,N_7569);
nand U8343 (N_8343,N_7613,N_7681);
or U8344 (N_8344,N_7528,N_7871);
nand U8345 (N_8345,N_7514,N_7556);
nand U8346 (N_8346,N_7639,N_7933);
nor U8347 (N_8347,N_7588,N_7596);
nor U8348 (N_8348,N_7562,N_7569);
nor U8349 (N_8349,N_7759,N_7858);
or U8350 (N_8350,N_7690,N_7862);
or U8351 (N_8351,N_7788,N_7545);
nor U8352 (N_8352,N_7664,N_7851);
nor U8353 (N_8353,N_7921,N_7893);
and U8354 (N_8354,N_7720,N_7874);
nor U8355 (N_8355,N_7859,N_7717);
or U8356 (N_8356,N_7658,N_7911);
and U8357 (N_8357,N_7929,N_7963);
xor U8358 (N_8358,N_7589,N_7950);
nor U8359 (N_8359,N_7849,N_7782);
xor U8360 (N_8360,N_7657,N_7644);
xnor U8361 (N_8361,N_7668,N_7508);
or U8362 (N_8362,N_7785,N_7764);
nand U8363 (N_8363,N_7953,N_7785);
and U8364 (N_8364,N_7509,N_7547);
xnor U8365 (N_8365,N_7954,N_7596);
nand U8366 (N_8366,N_7954,N_7896);
nand U8367 (N_8367,N_7793,N_7530);
and U8368 (N_8368,N_7736,N_7500);
nor U8369 (N_8369,N_7805,N_7862);
and U8370 (N_8370,N_7913,N_7815);
nand U8371 (N_8371,N_7513,N_7612);
and U8372 (N_8372,N_7553,N_7543);
or U8373 (N_8373,N_7739,N_7737);
and U8374 (N_8374,N_7898,N_7510);
xor U8375 (N_8375,N_7945,N_7705);
nor U8376 (N_8376,N_7877,N_7567);
nor U8377 (N_8377,N_7685,N_7509);
xor U8378 (N_8378,N_7923,N_7571);
and U8379 (N_8379,N_7887,N_7852);
nand U8380 (N_8380,N_7560,N_7960);
and U8381 (N_8381,N_7609,N_7840);
nand U8382 (N_8382,N_7817,N_7991);
or U8383 (N_8383,N_7838,N_7998);
and U8384 (N_8384,N_7812,N_7706);
or U8385 (N_8385,N_7714,N_7516);
or U8386 (N_8386,N_7791,N_7754);
nor U8387 (N_8387,N_7892,N_7768);
and U8388 (N_8388,N_7940,N_7989);
nand U8389 (N_8389,N_7959,N_7559);
and U8390 (N_8390,N_7622,N_7637);
nor U8391 (N_8391,N_7571,N_7501);
xnor U8392 (N_8392,N_7773,N_7884);
and U8393 (N_8393,N_7882,N_7593);
and U8394 (N_8394,N_7879,N_7795);
and U8395 (N_8395,N_7803,N_7853);
and U8396 (N_8396,N_7972,N_7834);
nand U8397 (N_8397,N_7768,N_7745);
and U8398 (N_8398,N_7777,N_7776);
nor U8399 (N_8399,N_7594,N_7656);
nor U8400 (N_8400,N_7770,N_7906);
nor U8401 (N_8401,N_7981,N_7675);
xor U8402 (N_8402,N_7735,N_7946);
nand U8403 (N_8403,N_7741,N_7711);
nor U8404 (N_8404,N_7854,N_7550);
nor U8405 (N_8405,N_7636,N_7587);
nand U8406 (N_8406,N_7540,N_7541);
nor U8407 (N_8407,N_7970,N_7750);
or U8408 (N_8408,N_7740,N_7750);
xor U8409 (N_8409,N_7579,N_7554);
nand U8410 (N_8410,N_7664,N_7984);
xnor U8411 (N_8411,N_7666,N_7517);
nand U8412 (N_8412,N_7967,N_7612);
nor U8413 (N_8413,N_7646,N_7534);
or U8414 (N_8414,N_7821,N_7637);
nand U8415 (N_8415,N_7632,N_7769);
xor U8416 (N_8416,N_7650,N_7712);
and U8417 (N_8417,N_7676,N_7880);
and U8418 (N_8418,N_7989,N_7606);
nor U8419 (N_8419,N_7754,N_7522);
nand U8420 (N_8420,N_7632,N_7516);
nand U8421 (N_8421,N_7783,N_7645);
and U8422 (N_8422,N_7659,N_7531);
and U8423 (N_8423,N_7620,N_7570);
or U8424 (N_8424,N_7671,N_7507);
xnor U8425 (N_8425,N_7699,N_7570);
and U8426 (N_8426,N_7980,N_7831);
xor U8427 (N_8427,N_7942,N_7544);
or U8428 (N_8428,N_7599,N_7967);
and U8429 (N_8429,N_7827,N_7966);
xnor U8430 (N_8430,N_7519,N_7575);
nor U8431 (N_8431,N_7758,N_7957);
nand U8432 (N_8432,N_7694,N_7905);
nor U8433 (N_8433,N_7870,N_7849);
or U8434 (N_8434,N_7712,N_7792);
nand U8435 (N_8435,N_7842,N_7784);
or U8436 (N_8436,N_7993,N_7763);
or U8437 (N_8437,N_7775,N_7547);
and U8438 (N_8438,N_7800,N_7754);
xor U8439 (N_8439,N_7690,N_7901);
or U8440 (N_8440,N_7744,N_7754);
xnor U8441 (N_8441,N_7808,N_7537);
and U8442 (N_8442,N_7522,N_7508);
xor U8443 (N_8443,N_7710,N_7869);
xor U8444 (N_8444,N_7659,N_7627);
nand U8445 (N_8445,N_7734,N_7811);
nand U8446 (N_8446,N_7783,N_7621);
and U8447 (N_8447,N_7610,N_7649);
xnor U8448 (N_8448,N_7512,N_7926);
and U8449 (N_8449,N_7696,N_7996);
or U8450 (N_8450,N_7824,N_7596);
or U8451 (N_8451,N_7953,N_7550);
xnor U8452 (N_8452,N_7528,N_7890);
nand U8453 (N_8453,N_7706,N_7591);
or U8454 (N_8454,N_7665,N_7904);
or U8455 (N_8455,N_7552,N_7877);
xor U8456 (N_8456,N_7604,N_7881);
and U8457 (N_8457,N_7526,N_7959);
xor U8458 (N_8458,N_7653,N_7580);
or U8459 (N_8459,N_7775,N_7576);
and U8460 (N_8460,N_7745,N_7551);
or U8461 (N_8461,N_7947,N_7760);
nor U8462 (N_8462,N_7608,N_7801);
xnor U8463 (N_8463,N_7995,N_7728);
and U8464 (N_8464,N_7930,N_7584);
and U8465 (N_8465,N_7513,N_7968);
and U8466 (N_8466,N_7940,N_7559);
nand U8467 (N_8467,N_7930,N_7845);
or U8468 (N_8468,N_7627,N_7529);
nand U8469 (N_8469,N_7824,N_7840);
nor U8470 (N_8470,N_7592,N_7991);
nand U8471 (N_8471,N_7649,N_7546);
nand U8472 (N_8472,N_7756,N_7612);
and U8473 (N_8473,N_7849,N_7506);
nand U8474 (N_8474,N_7846,N_7633);
nand U8475 (N_8475,N_7501,N_7570);
nor U8476 (N_8476,N_7820,N_7655);
or U8477 (N_8477,N_7682,N_7736);
xor U8478 (N_8478,N_7607,N_7931);
or U8479 (N_8479,N_7910,N_7780);
or U8480 (N_8480,N_7530,N_7649);
xnor U8481 (N_8481,N_7824,N_7701);
or U8482 (N_8482,N_7693,N_7696);
nor U8483 (N_8483,N_7682,N_7578);
xor U8484 (N_8484,N_7702,N_7955);
and U8485 (N_8485,N_7819,N_7604);
xnor U8486 (N_8486,N_7524,N_7964);
nor U8487 (N_8487,N_7762,N_7514);
or U8488 (N_8488,N_7950,N_7734);
xnor U8489 (N_8489,N_7757,N_7543);
or U8490 (N_8490,N_7702,N_7667);
or U8491 (N_8491,N_7791,N_7601);
or U8492 (N_8492,N_7872,N_7734);
nor U8493 (N_8493,N_7503,N_7509);
nor U8494 (N_8494,N_7702,N_7928);
xnor U8495 (N_8495,N_7905,N_7620);
and U8496 (N_8496,N_7796,N_7993);
nand U8497 (N_8497,N_7714,N_7995);
xor U8498 (N_8498,N_7600,N_7850);
or U8499 (N_8499,N_7726,N_7719);
or U8500 (N_8500,N_8283,N_8123);
and U8501 (N_8501,N_8164,N_8036);
xor U8502 (N_8502,N_8181,N_8020);
nand U8503 (N_8503,N_8156,N_8117);
nand U8504 (N_8504,N_8368,N_8197);
nor U8505 (N_8505,N_8246,N_8161);
and U8506 (N_8506,N_8370,N_8402);
or U8507 (N_8507,N_8353,N_8355);
xnor U8508 (N_8508,N_8139,N_8388);
and U8509 (N_8509,N_8339,N_8075);
nor U8510 (N_8510,N_8321,N_8147);
nand U8511 (N_8511,N_8333,N_8429);
or U8512 (N_8512,N_8041,N_8350);
xnor U8513 (N_8513,N_8016,N_8182);
nor U8514 (N_8514,N_8054,N_8057);
nor U8515 (N_8515,N_8132,N_8284);
nand U8516 (N_8516,N_8103,N_8486);
xor U8517 (N_8517,N_8449,N_8243);
and U8518 (N_8518,N_8496,N_8348);
nand U8519 (N_8519,N_8310,N_8296);
xor U8520 (N_8520,N_8395,N_8302);
or U8521 (N_8521,N_8211,N_8374);
or U8522 (N_8522,N_8437,N_8415);
or U8523 (N_8523,N_8300,N_8495);
nor U8524 (N_8524,N_8144,N_8462);
and U8525 (N_8525,N_8129,N_8116);
nor U8526 (N_8526,N_8479,N_8229);
and U8527 (N_8527,N_8095,N_8043);
and U8528 (N_8528,N_8155,N_8322);
xor U8529 (N_8529,N_8173,N_8040);
xor U8530 (N_8530,N_8491,N_8143);
nand U8531 (N_8531,N_8397,N_8213);
or U8532 (N_8532,N_8042,N_8039);
nand U8533 (N_8533,N_8024,N_8448);
nand U8534 (N_8534,N_8455,N_8193);
or U8535 (N_8535,N_8110,N_8025);
and U8536 (N_8536,N_8471,N_8192);
or U8537 (N_8537,N_8081,N_8417);
or U8538 (N_8538,N_8454,N_8240);
nor U8539 (N_8539,N_8421,N_8241);
nand U8540 (N_8540,N_8194,N_8021);
nand U8541 (N_8541,N_8049,N_8230);
nor U8542 (N_8542,N_8019,N_8320);
or U8543 (N_8543,N_8023,N_8003);
xnor U8544 (N_8544,N_8162,N_8314);
or U8545 (N_8545,N_8071,N_8382);
xor U8546 (N_8546,N_8094,N_8092);
nor U8547 (N_8547,N_8336,N_8074);
and U8548 (N_8548,N_8137,N_8485);
nand U8549 (N_8549,N_8121,N_8498);
nand U8550 (N_8550,N_8086,N_8221);
nand U8551 (N_8551,N_8004,N_8377);
and U8552 (N_8552,N_8325,N_8048);
nand U8553 (N_8553,N_8428,N_8233);
or U8554 (N_8554,N_8256,N_8465);
and U8555 (N_8555,N_8318,N_8247);
and U8556 (N_8556,N_8278,N_8038);
and U8557 (N_8557,N_8292,N_8072);
xnor U8558 (N_8558,N_8165,N_8286);
nand U8559 (N_8559,N_8150,N_8101);
and U8560 (N_8560,N_8207,N_8079);
xor U8561 (N_8561,N_8060,N_8487);
and U8562 (N_8562,N_8384,N_8196);
nor U8563 (N_8563,N_8249,N_8404);
and U8564 (N_8564,N_8359,N_8285);
nor U8565 (N_8565,N_8090,N_8408);
xnor U8566 (N_8566,N_8293,N_8070);
nand U8567 (N_8567,N_8442,N_8389);
nor U8568 (N_8568,N_8187,N_8309);
or U8569 (N_8569,N_8254,N_8223);
nand U8570 (N_8570,N_8112,N_8459);
nand U8571 (N_8571,N_8017,N_8064);
or U8572 (N_8572,N_8326,N_8014);
nand U8573 (N_8573,N_8306,N_8379);
nor U8574 (N_8574,N_8276,N_8030);
or U8575 (N_8575,N_8499,N_8251);
nor U8576 (N_8576,N_8138,N_8061);
nor U8577 (N_8577,N_8253,N_8401);
and U8578 (N_8578,N_8085,N_8105);
and U8579 (N_8579,N_8228,N_8218);
nand U8580 (N_8580,N_8472,N_8268);
nand U8581 (N_8581,N_8347,N_8441);
nor U8582 (N_8582,N_8266,N_8248);
nand U8583 (N_8583,N_8093,N_8447);
nand U8584 (N_8584,N_8476,N_8206);
xor U8585 (N_8585,N_8338,N_8494);
nand U8586 (N_8586,N_8290,N_8250);
or U8587 (N_8587,N_8035,N_8179);
xor U8588 (N_8588,N_8364,N_8420);
nand U8589 (N_8589,N_8443,N_8341);
and U8590 (N_8590,N_8015,N_8073);
or U8591 (N_8591,N_8434,N_8154);
and U8592 (N_8592,N_8099,N_8104);
nor U8593 (N_8593,N_8344,N_8198);
nand U8594 (N_8594,N_8470,N_8052);
nor U8595 (N_8595,N_8069,N_8467);
or U8596 (N_8596,N_8264,N_8331);
nand U8597 (N_8597,N_8190,N_8134);
nor U8598 (N_8598,N_8342,N_8340);
xor U8599 (N_8599,N_8189,N_8378);
nand U8600 (N_8600,N_8362,N_8214);
xor U8601 (N_8601,N_8390,N_8425);
and U8602 (N_8602,N_8363,N_8445);
nand U8603 (N_8603,N_8204,N_8169);
xor U8604 (N_8604,N_8352,N_8373);
nand U8605 (N_8605,N_8224,N_8080);
nand U8606 (N_8606,N_8232,N_8050);
nand U8607 (N_8607,N_8311,N_8385);
or U8608 (N_8608,N_8097,N_8063);
and U8609 (N_8609,N_8267,N_8012);
nor U8610 (N_8610,N_8131,N_8409);
and U8611 (N_8611,N_8394,N_8119);
xor U8612 (N_8612,N_8219,N_8062);
or U8613 (N_8613,N_8209,N_8469);
xor U8614 (N_8614,N_8010,N_8427);
xnor U8615 (N_8615,N_8055,N_8483);
or U8616 (N_8616,N_8089,N_8056);
or U8617 (N_8617,N_8399,N_8461);
nor U8618 (N_8618,N_8088,N_8332);
or U8619 (N_8619,N_8478,N_8002);
or U8620 (N_8620,N_8386,N_8177);
and U8621 (N_8621,N_8205,N_8130);
and U8622 (N_8622,N_8148,N_8013);
nand U8623 (N_8623,N_8414,N_8167);
and U8624 (N_8624,N_8203,N_8396);
nor U8625 (N_8625,N_8371,N_8329);
nand U8626 (N_8626,N_8185,N_8160);
nor U8627 (N_8627,N_8059,N_8031);
nand U8628 (N_8628,N_8210,N_8280);
nor U8629 (N_8629,N_8277,N_8127);
nand U8630 (N_8630,N_8453,N_8133);
xor U8631 (N_8631,N_8317,N_8343);
nand U8632 (N_8632,N_8180,N_8032);
xor U8633 (N_8633,N_8436,N_8078);
xor U8634 (N_8634,N_8307,N_8393);
nand U8635 (N_8635,N_8354,N_8327);
and U8636 (N_8636,N_8493,N_8297);
nor U8637 (N_8637,N_8000,N_8098);
and U8638 (N_8638,N_8466,N_8186);
or U8639 (N_8639,N_8323,N_8366);
xor U8640 (N_8640,N_8011,N_8313);
and U8641 (N_8641,N_8188,N_8225);
nand U8642 (N_8642,N_8083,N_8315);
xnor U8643 (N_8643,N_8244,N_8324);
or U8644 (N_8644,N_8065,N_8245);
or U8645 (N_8645,N_8199,N_8480);
and U8646 (N_8646,N_8022,N_8122);
nor U8647 (N_8647,N_8005,N_8145);
nand U8648 (N_8648,N_8450,N_8365);
and U8649 (N_8649,N_8482,N_8142);
and U8650 (N_8650,N_8236,N_8183);
xor U8651 (N_8651,N_8328,N_8158);
nor U8652 (N_8652,N_8288,N_8176);
xnor U8653 (N_8653,N_8360,N_8376);
xor U8654 (N_8654,N_8216,N_8195);
and U8655 (N_8655,N_8146,N_8361);
xor U8656 (N_8656,N_8452,N_8432);
and U8657 (N_8657,N_8303,N_8380);
nor U8658 (N_8658,N_8419,N_8231);
or U8659 (N_8659,N_8261,N_8044);
nor U8660 (N_8660,N_8426,N_8037);
xor U8661 (N_8661,N_8298,N_8416);
nand U8662 (N_8662,N_8367,N_8175);
and U8663 (N_8663,N_8460,N_8423);
nor U8664 (N_8664,N_8208,N_8227);
or U8665 (N_8665,N_8200,N_8084);
xnor U8666 (N_8666,N_8201,N_8438);
nand U8667 (N_8667,N_8001,N_8424);
nor U8668 (N_8668,N_8481,N_8212);
and U8669 (N_8669,N_8163,N_8255);
nor U8670 (N_8670,N_8058,N_8108);
nand U8671 (N_8671,N_8184,N_8444);
or U8672 (N_8672,N_8114,N_8281);
nor U8673 (N_8673,N_8463,N_8440);
nor U8674 (N_8674,N_8113,N_8222);
or U8675 (N_8675,N_8474,N_8008);
nor U8676 (N_8676,N_8140,N_8398);
or U8677 (N_8677,N_8282,N_8152);
or U8678 (N_8678,N_8490,N_8202);
and U8679 (N_8679,N_8330,N_8242);
nand U8680 (N_8680,N_8111,N_8118);
nand U8681 (N_8681,N_8149,N_8220);
nand U8682 (N_8682,N_8270,N_8489);
xor U8683 (N_8683,N_8392,N_8406);
nor U8684 (N_8684,N_8120,N_8067);
or U8685 (N_8685,N_8369,N_8431);
nor U8686 (N_8686,N_8435,N_8456);
nor U8687 (N_8687,N_8102,N_8274);
or U8688 (N_8688,N_8488,N_8279);
and U8689 (N_8689,N_8046,N_8115);
nand U8690 (N_8690,N_8295,N_8451);
or U8691 (N_8691,N_8226,N_8291);
nor U8692 (N_8692,N_8215,N_8430);
and U8693 (N_8693,N_8045,N_8172);
xnor U8694 (N_8694,N_8077,N_8497);
nand U8695 (N_8695,N_8034,N_8477);
or U8696 (N_8696,N_8337,N_8458);
xor U8697 (N_8697,N_8107,N_8334);
and U8698 (N_8698,N_8351,N_8076);
or U8699 (N_8699,N_8258,N_8252);
xor U8700 (N_8700,N_8109,N_8271);
and U8701 (N_8701,N_8407,N_8418);
and U8702 (N_8702,N_8457,N_8289);
or U8703 (N_8703,N_8126,N_8166);
xnor U8704 (N_8704,N_8287,N_8464);
xor U8705 (N_8705,N_8151,N_8217);
nand U8706 (N_8706,N_8124,N_8135);
nand U8707 (N_8707,N_8446,N_8141);
nand U8708 (N_8708,N_8433,N_8053);
or U8709 (N_8709,N_8191,N_8257);
nand U8710 (N_8710,N_8029,N_8128);
nor U8711 (N_8711,N_8492,N_8301);
and U8712 (N_8712,N_8082,N_8068);
or U8713 (N_8713,N_8051,N_8170);
or U8714 (N_8714,N_8412,N_8299);
nor U8715 (N_8715,N_8027,N_8066);
nand U8716 (N_8716,N_8304,N_8272);
nor U8717 (N_8717,N_8381,N_8273);
nand U8718 (N_8718,N_8007,N_8405);
nor U8719 (N_8719,N_8159,N_8346);
nand U8720 (N_8720,N_8157,N_8372);
or U8721 (N_8721,N_8391,N_8400);
xnor U8722 (N_8722,N_8403,N_8269);
nor U8723 (N_8723,N_8484,N_8383);
nor U8724 (N_8724,N_8375,N_8294);
and U8725 (N_8725,N_8239,N_8009);
and U8726 (N_8726,N_8262,N_8106);
nand U8727 (N_8727,N_8178,N_8305);
or U8728 (N_8728,N_8308,N_8234);
nor U8729 (N_8729,N_8263,N_8006);
and U8730 (N_8730,N_8475,N_8100);
nand U8731 (N_8731,N_8345,N_8357);
and U8732 (N_8732,N_8260,N_8473);
xor U8733 (N_8733,N_8335,N_8171);
nor U8734 (N_8734,N_8026,N_8358);
nor U8735 (N_8735,N_8387,N_8265);
and U8736 (N_8736,N_8168,N_8422);
nand U8737 (N_8737,N_8153,N_8439);
and U8738 (N_8738,N_8312,N_8047);
and U8739 (N_8739,N_8018,N_8468);
or U8740 (N_8740,N_8235,N_8033);
nor U8741 (N_8741,N_8096,N_8091);
and U8742 (N_8742,N_8410,N_8411);
nand U8743 (N_8743,N_8125,N_8319);
nor U8744 (N_8744,N_8316,N_8259);
and U8745 (N_8745,N_8238,N_8237);
or U8746 (N_8746,N_8136,N_8349);
and U8747 (N_8747,N_8028,N_8275);
xnor U8748 (N_8748,N_8356,N_8087);
or U8749 (N_8749,N_8413,N_8174);
nand U8750 (N_8750,N_8222,N_8008);
nor U8751 (N_8751,N_8185,N_8407);
xnor U8752 (N_8752,N_8436,N_8042);
nor U8753 (N_8753,N_8231,N_8150);
or U8754 (N_8754,N_8409,N_8159);
or U8755 (N_8755,N_8242,N_8320);
nand U8756 (N_8756,N_8196,N_8499);
xnor U8757 (N_8757,N_8418,N_8345);
or U8758 (N_8758,N_8483,N_8328);
xor U8759 (N_8759,N_8434,N_8453);
xnor U8760 (N_8760,N_8264,N_8431);
or U8761 (N_8761,N_8247,N_8014);
nor U8762 (N_8762,N_8038,N_8327);
xor U8763 (N_8763,N_8244,N_8122);
or U8764 (N_8764,N_8432,N_8244);
nand U8765 (N_8765,N_8282,N_8313);
or U8766 (N_8766,N_8043,N_8345);
nand U8767 (N_8767,N_8293,N_8121);
and U8768 (N_8768,N_8418,N_8406);
nand U8769 (N_8769,N_8163,N_8121);
and U8770 (N_8770,N_8143,N_8497);
nand U8771 (N_8771,N_8206,N_8173);
nor U8772 (N_8772,N_8125,N_8462);
or U8773 (N_8773,N_8190,N_8458);
nand U8774 (N_8774,N_8363,N_8345);
or U8775 (N_8775,N_8163,N_8193);
xor U8776 (N_8776,N_8286,N_8275);
nor U8777 (N_8777,N_8432,N_8316);
and U8778 (N_8778,N_8498,N_8328);
xnor U8779 (N_8779,N_8108,N_8354);
and U8780 (N_8780,N_8154,N_8017);
or U8781 (N_8781,N_8250,N_8295);
and U8782 (N_8782,N_8352,N_8307);
nand U8783 (N_8783,N_8247,N_8148);
nor U8784 (N_8784,N_8358,N_8022);
nor U8785 (N_8785,N_8371,N_8072);
nor U8786 (N_8786,N_8377,N_8416);
or U8787 (N_8787,N_8223,N_8397);
and U8788 (N_8788,N_8086,N_8237);
xor U8789 (N_8789,N_8489,N_8139);
nor U8790 (N_8790,N_8415,N_8373);
nand U8791 (N_8791,N_8095,N_8354);
xor U8792 (N_8792,N_8279,N_8030);
nand U8793 (N_8793,N_8158,N_8355);
or U8794 (N_8794,N_8141,N_8285);
xnor U8795 (N_8795,N_8152,N_8332);
nor U8796 (N_8796,N_8331,N_8393);
nand U8797 (N_8797,N_8288,N_8191);
nor U8798 (N_8798,N_8263,N_8009);
or U8799 (N_8799,N_8285,N_8139);
nand U8800 (N_8800,N_8441,N_8165);
nor U8801 (N_8801,N_8485,N_8161);
nor U8802 (N_8802,N_8230,N_8235);
nand U8803 (N_8803,N_8182,N_8054);
xnor U8804 (N_8804,N_8007,N_8344);
nand U8805 (N_8805,N_8059,N_8017);
nor U8806 (N_8806,N_8257,N_8420);
and U8807 (N_8807,N_8341,N_8170);
nor U8808 (N_8808,N_8271,N_8498);
nand U8809 (N_8809,N_8434,N_8323);
xor U8810 (N_8810,N_8346,N_8011);
xor U8811 (N_8811,N_8158,N_8475);
xor U8812 (N_8812,N_8442,N_8486);
nand U8813 (N_8813,N_8179,N_8372);
and U8814 (N_8814,N_8424,N_8106);
or U8815 (N_8815,N_8373,N_8200);
nand U8816 (N_8816,N_8387,N_8450);
nor U8817 (N_8817,N_8210,N_8106);
and U8818 (N_8818,N_8220,N_8347);
nand U8819 (N_8819,N_8251,N_8099);
and U8820 (N_8820,N_8126,N_8245);
nand U8821 (N_8821,N_8402,N_8385);
or U8822 (N_8822,N_8446,N_8486);
and U8823 (N_8823,N_8074,N_8484);
and U8824 (N_8824,N_8024,N_8019);
or U8825 (N_8825,N_8114,N_8371);
xor U8826 (N_8826,N_8194,N_8081);
or U8827 (N_8827,N_8219,N_8296);
nor U8828 (N_8828,N_8374,N_8244);
nor U8829 (N_8829,N_8211,N_8130);
and U8830 (N_8830,N_8131,N_8488);
nor U8831 (N_8831,N_8156,N_8412);
nor U8832 (N_8832,N_8483,N_8191);
nand U8833 (N_8833,N_8128,N_8095);
nand U8834 (N_8834,N_8028,N_8373);
or U8835 (N_8835,N_8118,N_8371);
and U8836 (N_8836,N_8101,N_8093);
xnor U8837 (N_8837,N_8404,N_8150);
nand U8838 (N_8838,N_8050,N_8369);
or U8839 (N_8839,N_8070,N_8381);
nor U8840 (N_8840,N_8273,N_8334);
nor U8841 (N_8841,N_8250,N_8352);
and U8842 (N_8842,N_8338,N_8478);
nor U8843 (N_8843,N_8324,N_8039);
nand U8844 (N_8844,N_8326,N_8203);
xnor U8845 (N_8845,N_8443,N_8417);
nand U8846 (N_8846,N_8329,N_8337);
nand U8847 (N_8847,N_8222,N_8456);
nand U8848 (N_8848,N_8435,N_8008);
nor U8849 (N_8849,N_8409,N_8438);
and U8850 (N_8850,N_8075,N_8363);
xor U8851 (N_8851,N_8126,N_8390);
xor U8852 (N_8852,N_8208,N_8262);
and U8853 (N_8853,N_8172,N_8237);
nor U8854 (N_8854,N_8349,N_8025);
xor U8855 (N_8855,N_8192,N_8293);
and U8856 (N_8856,N_8142,N_8018);
nand U8857 (N_8857,N_8430,N_8413);
nand U8858 (N_8858,N_8240,N_8183);
xor U8859 (N_8859,N_8497,N_8073);
nand U8860 (N_8860,N_8187,N_8282);
nand U8861 (N_8861,N_8079,N_8291);
nand U8862 (N_8862,N_8389,N_8192);
or U8863 (N_8863,N_8019,N_8082);
xnor U8864 (N_8864,N_8058,N_8156);
and U8865 (N_8865,N_8272,N_8088);
and U8866 (N_8866,N_8070,N_8184);
nor U8867 (N_8867,N_8091,N_8200);
nor U8868 (N_8868,N_8042,N_8295);
and U8869 (N_8869,N_8378,N_8266);
nor U8870 (N_8870,N_8061,N_8100);
and U8871 (N_8871,N_8313,N_8446);
or U8872 (N_8872,N_8190,N_8034);
and U8873 (N_8873,N_8091,N_8022);
xor U8874 (N_8874,N_8096,N_8371);
and U8875 (N_8875,N_8303,N_8478);
xnor U8876 (N_8876,N_8001,N_8291);
and U8877 (N_8877,N_8386,N_8037);
xnor U8878 (N_8878,N_8174,N_8143);
nand U8879 (N_8879,N_8171,N_8319);
nor U8880 (N_8880,N_8173,N_8015);
and U8881 (N_8881,N_8075,N_8069);
and U8882 (N_8882,N_8099,N_8465);
nor U8883 (N_8883,N_8144,N_8032);
and U8884 (N_8884,N_8305,N_8099);
and U8885 (N_8885,N_8165,N_8164);
nand U8886 (N_8886,N_8346,N_8233);
xor U8887 (N_8887,N_8093,N_8367);
nand U8888 (N_8888,N_8492,N_8274);
or U8889 (N_8889,N_8051,N_8401);
or U8890 (N_8890,N_8091,N_8426);
nand U8891 (N_8891,N_8409,N_8309);
nor U8892 (N_8892,N_8041,N_8182);
nand U8893 (N_8893,N_8351,N_8141);
nor U8894 (N_8894,N_8433,N_8421);
and U8895 (N_8895,N_8341,N_8330);
nand U8896 (N_8896,N_8259,N_8206);
nand U8897 (N_8897,N_8070,N_8384);
xnor U8898 (N_8898,N_8140,N_8450);
nor U8899 (N_8899,N_8096,N_8252);
or U8900 (N_8900,N_8207,N_8428);
and U8901 (N_8901,N_8077,N_8056);
nand U8902 (N_8902,N_8122,N_8478);
nor U8903 (N_8903,N_8498,N_8375);
xor U8904 (N_8904,N_8434,N_8192);
and U8905 (N_8905,N_8104,N_8011);
or U8906 (N_8906,N_8199,N_8087);
nand U8907 (N_8907,N_8265,N_8147);
xnor U8908 (N_8908,N_8176,N_8332);
nand U8909 (N_8909,N_8216,N_8077);
xor U8910 (N_8910,N_8365,N_8474);
or U8911 (N_8911,N_8152,N_8352);
and U8912 (N_8912,N_8362,N_8077);
nand U8913 (N_8913,N_8482,N_8422);
or U8914 (N_8914,N_8036,N_8210);
or U8915 (N_8915,N_8273,N_8175);
xor U8916 (N_8916,N_8434,N_8175);
and U8917 (N_8917,N_8467,N_8408);
nand U8918 (N_8918,N_8038,N_8317);
xnor U8919 (N_8919,N_8005,N_8105);
or U8920 (N_8920,N_8390,N_8216);
and U8921 (N_8921,N_8253,N_8027);
nor U8922 (N_8922,N_8037,N_8017);
and U8923 (N_8923,N_8154,N_8232);
nor U8924 (N_8924,N_8403,N_8143);
nor U8925 (N_8925,N_8489,N_8482);
xnor U8926 (N_8926,N_8380,N_8074);
nand U8927 (N_8927,N_8298,N_8214);
or U8928 (N_8928,N_8422,N_8480);
nand U8929 (N_8929,N_8421,N_8404);
nor U8930 (N_8930,N_8125,N_8470);
and U8931 (N_8931,N_8177,N_8392);
nor U8932 (N_8932,N_8070,N_8386);
and U8933 (N_8933,N_8080,N_8094);
or U8934 (N_8934,N_8275,N_8292);
and U8935 (N_8935,N_8265,N_8315);
or U8936 (N_8936,N_8426,N_8481);
nand U8937 (N_8937,N_8150,N_8211);
and U8938 (N_8938,N_8006,N_8016);
nor U8939 (N_8939,N_8108,N_8274);
nor U8940 (N_8940,N_8113,N_8083);
and U8941 (N_8941,N_8298,N_8174);
or U8942 (N_8942,N_8344,N_8419);
or U8943 (N_8943,N_8323,N_8149);
nand U8944 (N_8944,N_8465,N_8094);
nand U8945 (N_8945,N_8471,N_8285);
and U8946 (N_8946,N_8283,N_8446);
or U8947 (N_8947,N_8018,N_8369);
xnor U8948 (N_8948,N_8086,N_8163);
nor U8949 (N_8949,N_8343,N_8054);
or U8950 (N_8950,N_8415,N_8231);
xnor U8951 (N_8951,N_8081,N_8210);
nor U8952 (N_8952,N_8092,N_8364);
nor U8953 (N_8953,N_8146,N_8371);
xnor U8954 (N_8954,N_8131,N_8321);
xor U8955 (N_8955,N_8008,N_8460);
or U8956 (N_8956,N_8063,N_8079);
nor U8957 (N_8957,N_8082,N_8247);
and U8958 (N_8958,N_8162,N_8170);
xnor U8959 (N_8959,N_8097,N_8239);
nor U8960 (N_8960,N_8150,N_8487);
xor U8961 (N_8961,N_8079,N_8442);
or U8962 (N_8962,N_8070,N_8128);
nor U8963 (N_8963,N_8052,N_8150);
nand U8964 (N_8964,N_8499,N_8106);
nand U8965 (N_8965,N_8357,N_8111);
or U8966 (N_8966,N_8394,N_8380);
nand U8967 (N_8967,N_8197,N_8087);
xor U8968 (N_8968,N_8110,N_8393);
nand U8969 (N_8969,N_8392,N_8471);
nand U8970 (N_8970,N_8154,N_8480);
or U8971 (N_8971,N_8064,N_8114);
and U8972 (N_8972,N_8408,N_8379);
and U8973 (N_8973,N_8432,N_8229);
or U8974 (N_8974,N_8381,N_8245);
nand U8975 (N_8975,N_8014,N_8301);
xnor U8976 (N_8976,N_8410,N_8263);
and U8977 (N_8977,N_8251,N_8483);
or U8978 (N_8978,N_8384,N_8058);
xnor U8979 (N_8979,N_8454,N_8401);
xor U8980 (N_8980,N_8241,N_8320);
nand U8981 (N_8981,N_8085,N_8207);
xnor U8982 (N_8982,N_8271,N_8290);
xnor U8983 (N_8983,N_8000,N_8107);
nand U8984 (N_8984,N_8400,N_8231);
xnor U8985 (N_8985,N_8343,N_8256);
nand U8986 (N_8986,N_8016,N_8461);
nor U8987 (N_8987,N_8464,N_8278);
and U8988 (N_8988,N_8187,N_8466);
or U8989 (N_8989,N_8408,N_8175);
and U8990 (N_8990,N_8486,N_8025);
or U8991 (N_8991,N_8133,N_8340);
nor U8992 (N_8992,N_8160,N_8400);
and U8993 (N_8993,N_8229,N_8347);
nand U8994 (N_8994,N_8050,N_8019);
and U8995 (N_8995,N_8047,N_8040);
nand U8996 (N_8996,N_8357,N_8411);
or U8997 (N_8997,N_8487,N_8039);
and U8998 (N_8998,N_8150,N_8057);
or U8999 (N_8999,N_8009,N_8388);
nor U9000 (N_9000,N_8816,N_8612);
nor U9001 (N_9001,N_8616,N_8715);
nor U9002 (N_9002,N_8844,N_8855);
nand U9003 (N_9003,N_8961,N_8545);
and U9004 (N_9004,N_8898,N_8508);
xnor U9005 (N_9005,N_8851,N_8659);
xor U9006 (N_9006,N_8657,N_8569);
nand U9007 (N_9007,N_8686,N_8631);
nand U9008 (N_9008,N_8893,N_8877);
nand U9009 (N_9009,N_8978,N_8505);
and U9010 (N_9010,N_8741,N_8788);
nand U9011 (N_9011,N_8534,N_8941);
xor U9012 (N_9012,N_8624,N_8579);
or U9013 (N_9013,N_8949,N_8539);
xor U9014 (N_9014,N_8845,N_8738);
nor U9015 (N_9015,N_8967,N_8608);
or U9016 (N_9016,N_8792,N_8717);
xnor U9017 (N_9017,N_8630,N_8884);
nand U9018 (N_9018,N_8793,N_8536);
and U9019 (N_9019,N_8698,N_8916);
or U9020 (N_9020,N_8869,N_8618);
and U9021 (N_9021,N_8521,N_8511);
and U9022 (N_9022,N_8925,N_8981);
and U9023 (N_9023,N_8901,N_8871);
nand U9024 (N_9024,N_8693,N_8723);
or U9025 (N_9025,N_8522,N_8736);
nand U9026 (N_9026,N_8990,N_8950);
nor U9027 (N_9027,N_8640,N_8790);
nor U9028 (N_9028,N_8839,N_8734);
xor U9029 (N_9029,N_8840,N_8722);
nor U9030 (N_9030,N_8865,N_8553);
and U9031 (N_9031,N_8680,N_8627);
or U9032 (N_9032,N_8571,N_8720);
nor U9033 (N_9033,N_8746,N_8908);
xor U9034 (N_9034,N_8825,N_8555);
or U9035 (N_9035,N_8643,N_8711);
xnor U9036 (N_9036,N_8633,N_8668);
xor U9037 (N_9037,N_8853,N_8594);
or U9038 (N_9038,N_8994,N_8516);
and U9039 (N_9039,N_8795,N_8577);
xor U9040 (N_9040,N_8747,N_8502);
nor U9041 (N_9041,N_8581,N_8781);
and U9042 (N_9042,N_8929,N_8974);
and U9043 (N_9043,N_8847,N_8989);
nor U9044 (N_9044,N_8743,N_8751);
or U9045 (N_9045,N_8661,N_8507);
and U9046 (N_9046,N_8917,N_8862);
or U9047 (N_9047,N_8671,N_8824);
nor U9048 (N_9048,N_8922,N_8718);
nor U9049 (N_9049,N_8510,N_8591);
nand U9050 (N_9050,N_8762,N_8683);
nand U9051 (N_9051,N_8637,N_8979);
nand U9052 (N_9052,N_8911,N_8954);
or U9053 (N_9053,N_8632,N_8697);
and U9054 (N_9054,N_8613,N_8710);
nand U9055 (N_9055,N_8764,N_8660);
nand U9056 (N_9056,N_8966,N_8857);
and U9057 (N_9057,N_8943,N_8754);
or U9058 (N_9058,N_8912,N_8780);
nand U9059 (N_9059,N_8573,N_8810);
xor U9060 (N_9060,N_8776,N_8551);
nand U9061 (N_9061,N_8629,N_8712);
xor U9062 (N_9062,N_8956,N_8849);
and U9063 (N_9063,N_8604,N_8935);
nand U9064 (N_9064,N_8542,N_8533);
and U9065 (N_9065,N_8938,N_8889);
nor U9066 (N_9066,N_8888,N_8782);
and U9067 (N_9067,N_8834,N_8813);
or U9068 (N_9068,N_8999,N_8867);
or U9069 (N_9069,N_8891,N_8980);
xor U9070 (N_9070,N_8965,N_8662);
nor U9071 (N_9071,N_8984,N_8859);
and U9072 (N_9072,N_8778,N_8786);
xnor U9073 (N_9073,N_8763,N_8727);
nor U9074 (N_9074,N_8615,N_8596);
nand U9075 (N_9075,N_8652,N_8599);
and U9076 (N_9076,N_8572,N_8537);
xor U9077 (N_9077,N_8815,N_8692);
nand U9078 (N_9078,N_8945,N_8977);
xnor U9079 (N_9079,N_8735,N_8872);
and U9080 (N_9080,N_8863,N_8759);
nand U9081 (N_9081,N_8868,N_8923);
or U9082 (N_9082,N_8664,N_8873);
xnor U9083 (N_9083,N_8852,N_8899);
nor U9084 (N_9084,N_8948,N_8695);
nor U9085 (N_9085,N_8641,N_8988);
xor U9086 (N_9086,N_8798,N_8688);
nand U9087 (N_9087,N_8940,N_8523);
nor U9088 (N_9088,N_8674,N_8766);
or U9089 (N_9089,N_8924,N_8757);
nand U9090 (N_9090,N_8562,N_8670);
nor U9091 (N_9091,N_8517,N_8655);
nor U9092 (N_9092,N_8706,N_8713);
and U9093 (N_9093,N_8580,N_8983);
and U9094 (N_9094,N_8559,N_8827);
xnor U9095 (N_9095,N_8520,N_8907);
nand U9096 (N_9096,N_8957,N_8566);
nand U9097 (N_9097,N_8666,N_8783);
nor U9098 (N_9098,N_8601,N_8600);
nor U9099 (N_9099,N_8811,N_8973);
xnor U9100 (N_9100,N_8719,N_8684);
and U9101 (N_9101,N_8543,N_8906);
xor U9102 (N_9102,N_8787,N_8875);
xor U9103 (N_9103,N_8739,N_8856);
nor U9104 (N_9104,N_8634,N_8879);
xnor U9105 (N_9105,N_8583,N_8947);
and U9106 (N_9106,N_8703,N_8714);
or U9107 (N_9107,N_8742,N_8667);
and U9108 (N_9108,N_8676,N_8682);
or U9109 (N_9109,N_8858,N_8535);
nor U9110 (N_9110,N_8876,N_8942);
nor U9111 (N_9111,N_8673,N_8937);
xor U9112 (N_9112,N_8531,N_8821);
and U9113 (N_9113,N_8915,N_8595);
nand U9114 (N_9114,N_8642,N_8758);
nor U9115 (N_9115,N_8690,N_8568);
xor U9116 (N_9116,N_8982,N_8920);
nor U9117 (N_9117,N_8696,N_8773);
or U9118 (N_9118,N_8833,N_8576);
nand U9119 (N_9119,N_8809,N_8808);
nand U9120 (N_9120,N_8678,N_8733);
xnor U9121 (N_9121,N_8800,N_8694);
nand U9122 (N_9122,N_8584,N_8638);
nor U9123 (N_9123,N_8930,N_8802);
xnor U9124 (N_9124,N_8606,N_8585);
nor U9125 (N_9125,N_8646,N_8563);
and U9126 (N_9126,N_8928,N_8603);
nand U9127 (N_9127,N_8968,N_8570);
nor U9128 (N_9128,N_8895,N_8910);
and U9129 (N_9129,N_8902,N_8817);
xor U9130 (N_9130,N_8550,N_8650);
xnor U9131 (N_9131,N_8832,N_8748);
nor U9132 (N_9132,N_8512,N_8995);
nand U9133 (N_9133,N_8985,N_8900);
xnor U9134 (N_9134,N_8997,N_8665);
nor U9135 (N_9135,N_8610,N_8532);
nand U9136 (N_9136,N_8970,N_8677);
nand U9137 (N_9137,N_8565,N_8560);
xnor U9138 (N_9138,N_8654,N_8885);
xnor U9139 (N_9139,N_8614,N_8647);
or U9140 (N_9140,N_8896,N_8913);
or U9141 (N_9141,N_8503,N_8651);
nor U9142 (N_9142,N_8784,N_8644);
or U9143 (N_9143,N_8744,N_8737);
xor U9144 (N_9144,N_8575,N_8767);
xor U9145 (N_9145,N_8609,N_8500);
nor U9146 (N_9146,N_8826,N_8894);
nand U9147 (N_9147,N_8526,N_8904);
xor U9148 (N_9148,N_8883,N_8504);
xor U9149 (N_9149,N_8831,N_8953);
nor U9150 (N_9150,N_8679,N_8626);
or U9151 (N_9151,N_8952,N_8528);
nor U9152 (N_9152,N_8992,N_8963);
nor U9153 (N_9153,N_8552,N_8617);
nor U9154 (N_9154,N_8549,N_8556);
nor U9155 (N_9155,N_8636,N_8903);
or U9156 (N_9156,N_8529,N_8822);
or U9157 (N_9157,N_8774,N_8527);
nor U9158 (N_9158,N_8602,N_8509);
xnor U9159 (N_9159,N_8590,N_8777);
and U9160 (N_9160,N_8843,N_8672);
or U9161 (N_9161,N_8598,N_8707);
or U9162 (N_9162,N_8622,N_8881);
nand U9163 (N_9163,N_8880,N_8918);
and U9164 (N_9164,N_8854,N_8975);
or U9165 (N_9165,N_8892,N_8506);
and U9166 (N_9166,N_8998,N_8501);
and U9167 (N_9167,N_8791,N_8548);
and U9168 (N_9168,N_8753,N_8860);
nand U9169 (N_9169,N_8820,N_8905);
or U9170 (N_9170,N_8756,N_8789);
and U9171 (N_9171,N_8681,N_8926);
nor U9172 (N_9172,N_8530,N_8933);
nand U9173 (N_9173,N_8829,N_8619);
xor U9174 (N_9174,N_8897,N_8700);
nor U9175 (N_9175,N_8927,N_8721);
or U9176 (N_9176,N_8567,N_8732);
xnor U9177 (N_9177,N_8772,N_8882);
and U9178 (N_9178,N_8760,N_8823);
and U9179 (N_9179,N_8592,N_8709);
xor U9180 (N_9180,N_8675,N_8837);
xor U9181 (N_9181,N_8547,N_8639);
nor U9182 (N_9182,N_8538,N_8976);
xor U9183 (N_9183,N_8931,N_8705);
xor U9184 (N_9184,N_8574,N_8724);
xnor U9185 (N_9185,N_8991,N_8740);
or U9186 (N_9186,N_8969,N_8525);
nand U9187 (N_9187,N_8914,N_8519);
or U9188 (N_9188,N_8861,N_8761);
nand U9189 (N_9189,N_8835,N_8623);
nor U9190 (N_9190,N_8749,N_8804);
or U9191 (N_9191,N_8770,N_8801);
nand U9192 (N_9192,N_8663,N_8726);
and U9193 (N_9193,N_8771,N_8807);
xor U9194 (N_9194,N_8582,N_8846);
and U9195 (N_9195,N_8794,N_8611);
and U9196 (N_9196,N_8635,N_8814);
nor U9197 (N_9197,N_8716,N_8909);
nor U9198 (N_9198,N_8620,N_8605);
or U9199 (N_9199,N_8962,N_8944);
nand U9200 (N_9200,N_8725,N_8828);
nand U9201 (N_9201,N_8607,N_8993);
or U9202 (N_9202,N_8874,N_8838);
and U9203 (N_9203,N_8669,N_8730);
nand U9204 (N_9204,N_8701,N_8518);
nor U9205 (N_9205,N_8936,N_8964);
or U9206 (N_9206,N_8812,N_8752);
or U9207 (N_9207,N_8541,N_8951);
nand U9208 (N_9208,N_8587,N_8554);
nor U9209 (N_9209,N_8960,N_8546);
and U9210 (N_9210,N_8987,N_8887);
or U9211 (N_9211,N_8799,N_8775);
and U9212 (N_9212,N_8768,N_8524);
xnor U9213 (N_9213,N_8955,N_8658);
and U9214 (N_9214,N_8625,N_8919);
xor U9215 (N_9215,N_8557,N_8996);
nor U9216 (N_9216,N_8729,N_8842);
and U9217 (N_9217,N_8765,N_8586);
and U9218 (N_9218,N_8841,N_8769);
and U9219 (N_9219,N_8870,N_8731);
nor U9220 (N_9220,N_8685,N_8702);
or U9221 (N_9221,N_8797,N_8515);
nor U9222 (N_9222,N_8785,N_8745);
xor U9223 (N_9223,N_8621,N_8958);
xor U9224 (N_9224,N_8878,N_8818);
xnor U9225 (N_9225,N_8971,N_8934);
nand U9226 (N_9226,N_8819,N_8561);
or U9227 (N_9227,N_8972,N_8803);
xnor U9228 (N_9228,N_8558,N_8645);
nor U9229 (N_9229,N_8755,N_8848);
xor U9230 (N_9230,N_8513,N_8540);
nand U9231 (N_9231,N_8830,N_8564);
or U9232 (N_9232,N_8691,N_8589);
and U9233 (N_9233,N_8578,N_8656);
and U9234 (N_9234,N_8708,N_8514);
xor U9235 (N_9235,N_8836,N_8886);
xnor U9236 (N_9236,N_8728,N_8544);
and U9237 (N_9237,N_8704,N_8921);
or U9238 (N_9238,N_8959,N_8850);
nand U9239 (N_9239,N_8939,N_8628);
and U9240 (N_9240,N_8593,N_8653);
xor U9241 (N_9241,N_8796,N_8986);
nor U9242 (N_9242,N_8649,N_8648);
xnor U9243 (N_9243,N_8890,N_8588);
and U9244 (N_9244,N_8805,N_8687);
xor U9245 (N_9245,N_8689,N_8750);
nor U9246 (N_9246,N_8946,N_8699);
or U9247 (N_9247,N_8932,N_8779);
and U9248 (N_9248,N_8864,N_8597);
and U9249 (N_9249,N_8806,N_8866);
nor U9250 (N_9250,N_8777,N_8548);
or U9251 (N_9251,N_8643,N_8811);
xor U9252 (N_9252,N_8603,N_8574);
or U9253 (N_9253,N_8757,N_8901);
xnor U9254 (N_9254,N_8859,N_8720);
nand U9255 (N_9255,N_8793,N_8921);
nor U9256 (N_9256,N_8845,N_8754);
nor U9257 (N_9257,N_8916,N_8587);
or U9258 (N_9258,N_8686,N_8742);
nand U9259 (N_9259,N_8514,N_8725);
xor U9260 (N_9260,N_8732,N_8750);
nand U9261 (N_9261,N_8843,N_8795);
nor U9262 (N_9262,N_8963,N_8835);
and U9263 (N_9263,N_8951,N_8983);
and U9264 (N_9264,N_8635,N_8749);
and U9265 (N_9265,N_8956,N_8746);
xor U9266 (N_9266,N_8758,N_8715);
nor U9267 (N_9267,N_8545,N_8819);
or U9268 (N_9268,N_8698,N_8964);
or U9269 (N_9269,N_8568,N_8725);
or U9270 (N_9270,N_8973,N_8997);
nand U9271 (N_9271,N_8548,N_8772);
xor U9272 (N_9272,N_8581,N_8986);
and U9273 (N_9273,N_8841,N_8580);
and U9274 (N_9274,N_8965,N_8769);
or U9275 (N_9275,N_8867,N_8554);
xnor U9276 (N_9276,N_8865,N_8919);
and U9277 (N_9277,N_8904,N_8674);
xor U9278 (N_9278,N_8668,N_8546);
or U9279 (N_9279,N_8732,N_8766);
nand U9280 (N_9280,N_8612,N_8727);
and U9281 (N_9281,N_8908,N_8547);
nor U9282 (N_9282,N_8925,N_8619);
nand U9283 (N_9283,N_8625,N_8791);
xor U9284 (N_9284,N_8612,N_8836);
or U9285 (N_9285,N_8786,N_8794);
or U9286 (N_9286,N_8870,N_8983);
nand U9287 (N_9287,N_8931,N_8792);
nand U9288 (N_9288,N_8901,N_8728);
nand U9289 (N_9289,N_8912,N_8778);
nor U9290 (N_9290,N_8743,N_8670);
or U9291 (N_9291,N_8748,N_8780);
xor U9292 (N_9292,N_8650,N_8975);
or U9293 (N_9293,N_8908,N_8737);
and U9294 (N_9294,N_8647,N_8835);
nor U9295 (N_9295,N_8722,N_8981);
and U9296 (N_9296,N_8669,N_8554);
nor U9297 (N_9297,N_8836,N_8757);
and U9298 (N_9298,N_8968,N_8901);
xor U9299 (N_9299,N_8722,N_8864);
or U9300 (N_9300,N_8874,N_8933);
and U9301 (N_9301,N_8689,N_8695);
xor U9302 (N_9302,N_8889,N_8669);
xnor U9303 (N_9303,N_8868,N_8600);
xnor U9304 (N_9304,N_8743,N_8897);
xnor U9305 (N_9305,N_8967,N_8929);
and U9306 (N_9306,N_8903,N_8919);
nor U9307 (N_9307,N_8615,N_8907);
xnor U9308 (N_9308,N_8752,N_8764);
xnor U9309 (N_9309,N_8925,N_8747);
xnor U9310 (N_9310,N_8709,N_8858);
xnor U9311 (N_9311,N_8815,N_8513);
xor U9312 (N_9312,N_8703,N_8707);
and U9313 (N_9313,N_8978,N_8796);
and U9314 (N_9314,N_8745,N_8605);
xnor U9315 (N_9315,N_8889,N_8751);
or U9316 (N_9316,N_8536,N_8766);
xnor U9317 (N_9317,N_8773,N_8893);
xor U9318 (N_9318,N_8897,N_8960);
nand U9319 (N_9319,N_8866,N_8957);
and U9320 (N_9320,N_8672,N_8862);
nor U9321 (N_9321,N_8861,N_8909);
or U9322 (N_9322,N_8871,N_8744);
xor U9323 (N_9323,N_8969,N_8512);
nor U9324 (N_9324,N_8770,N_8755);
xor U9325 (N_9325,N_8987,N_8699);
xnor U9326 (N_9326,N_8972,N_8817);
xnor U9327 (N_9327,N_8841,N_8571);
or U9328 (N_9328,N_8581,N_8828);
nor U9329 (N_9329,N_8826,N_8949);
nor U9330 (N_9330,N_8745,N_8513);
nand U9331 (N_9331,N_8607,N_8520);
nand U9332 (N_9332,N_8762,N_8839);
nand U9333 (N_9333,N_8644,N_8533);
xor U9334 (N_9334,N_8885,N_8848);
nand U9335 (N_9335,N_8824,N_8582);
nor U9336 (N_9336,N_8683,N_8591);
xnor U9337 (N_9337,N_8686,N_8509);
and U9338 (N_9338,N_8932,N_8902);
or U9339 (N_9339,N_8873,N_8636);
or U9340 (N_9340,N_8528,N_8541);
and U9341 (N_9341,N_8701,N_8798);
and U9342 (N_9342,N_8777,N_8571);
and U9343 (N_9343,N_8656,N_8735);
nor U9344 (N_9344,N_8542,N_8826);
nor U9345 (N_9345,N_8648,N_8843);
or U9346 (N_9346,N_8506,N_8570);
nand U9347 (N_9347,N_8571,N_8675);
or U9348 (N_9348,N_8744,N_8617);
xnor U9349 (N_9349,N_8517,N_8789);
xnor U9350 (N_9350,N_8786,N_8881);
nor U9351 (N_9351,N_8995,N_8702);
xor U9352 (N_9352,N_8517,N_8524);
or U9353 (N_9353,N_8797,N_8689);
xor U9354 (N_9354,N_8716,N_8918);
nand U9355 (N_9355,N_8806,N_8545);
nor U9356 (N_9356,N_8929,N_8805);
nand U9357 (N_9357,N_8735,N_8650);
nand U9358 (N_9358,N_8512,N_8590);
nor U9359 (N_9359,N_8773,N_8755);
nor U9360 (N_9360,N_8822,N_8570);
nand U9361 (N_9361,N_8882,N_8785);
or U9362 (N_9362,N_8676,N_8559);
nor U9363 (N_9363,N_8723,N_8662);
nand U9364 (N_9364,N_8837,N_8509);
nor U9365 (N_9365,N_8951,N_8597);
or U9366 (N_9366,N_8835,N_8767);
xnor U9367 (N_9367,N_8714,N_8577);
and U9368 (N_9368,N_8573,N_8753);
and U9369 (N_9369,N_8779,N_8628);
and U9370 (N_9370,N_8651,N_8689);
and U9371 (N_9371,N_8990,N_8673);
nand U9372 (N_9372,N_8727,N_8554);
nor U9373 (N_9373,N_8711,N_8753);
and U9374 (N_9374,N_8773,N_8825);
and U9375 (N_9375,N_8661,N_8961);
and U9376 (N_9376,N_8676,N_8641);
and U9377 (N_9377,N_8794,N_8910);
xnor U9378 (N_9378,N_8979,N_8984);
or U9379 (N_9379,N_8630,N_8767);
xor U9380 (N_9380,N_8965,N_8847);
nand U9381 (N_9381,N_8660,N_8530);
nand U9382 (N_9382,N_8595,N_8884);
nor U9383 (N_9383,N_8741,N_8625);
xnor U9384 (N_9384,N_8996,N_8786);
xor U9385 (N_9385,N_8917,N_8951);
nor U9386 (N_9386,N_8991,N_8536);
nand U9387 (N_9387,N_8689,N_8640);
nand U9388 (N_9388,N_8731,N_8814);
and U9389 (N_9389,N_8740,N_8900);
xor U9390 (N_9390,N_8529,N_8874);
xnor U9391 (N_9391,N_8544,N_8644);
nor U9392 (N_9392,N_8820,N_8747);
and U9393 (N_9393,N_8531,N_8528);
nor U9394 (N_9394,N_8509,N_8680);
xnor U9395 (N_9395,N_8707,N_8848);
or U9396 (N_9396,N_8916,N_8807);
nor U9397 (N_9397,N_8665,N_8884);
or U9398 (N_9398,N_8896,N_8875);
xnor U9399 (N_9399,N_8661,N_8898);
and U9400 (N_9400,N_8791,N_8662);
and U9401 (N_9401,N_8798,N_8974);
nor U9402 (N_9402,N_8636,N_8814);
nor U9403 (N_9403,N_8704,N_8840);
and U9404 (N_9404,N_8632,N_8509);
nand U9405 (N_9405,N_8654,N_8827);
nor U9406 (N_9406,N_8740,N_8542);
nor U9407 (N_9407,N_8693,N_8590);
and U9408 (N_9408,N_8513,N_8811);
and U9409 (N_9409,N_8834,N_8974);
xor U9410 (N_9410,N_8735,N_8540);
xnor U9411 (N_9411,N_8808,N_8667);
nor U9412 (N_9412,N_8942,N_8609);
xor U9413 (N_9413,N_8987,N_8600);
and U9414 (N_9414,N_8818,N_8584);
and U9415 (N_9415,N_8615,N_8537);
xnor U9416 (N_9416,N_8938,N_8669);
nor U9417 (N_9417,N_8918,N_8839);
xor U9418 (N_9418,N_8635,N_8539);
nand U9419 (N_9419,N_8989,N_8710);
nor U9420 (N_9420,N_8907,N_8717);
nand U9421 (N_9421,N_8756,N_8992);
or U9422 (N_9422,N_8721,N_8993);
and U9423 (N_9423,N_8662,N_8581);
or U9424 (N_9424,N_8870,N_8880);
or U9425 (N_9425,N_8582,N_8901);
or U9426 (N_9426,N_8813,N_8769);
xor U9427 (N_9427,N_8549,N_8649);
xor U9428 (N_9428,N_8947,N_8767);
and U9429 (N_9429,N_8998,N_8885);
and U9430 (N_9430,N_8934,N_8902);
xor U9431 (N_9431,N_8914,N_8783);
and U9432 (N_9432,N_8951,N_8672);
xor U9433 (N_9433,N_8749,N_8656);
nor U9434 (N_9434,N_8674,N_8754);
nand U9435 (N_9435,N_8966,N_8808);
nand U9436 (N_9436,N_8592,N_8811);
xor U9437 (N_9437,N_8790,N_8828);
nand U9438 (N_9438,N_8637,N_8639);
nor U9439 (N_9439,N_8654,N_8547);
nor U9440 (N_9440,N_8663,N_8785);
and U9441 (N_9441,N_8535,N_8754);
nand U9442 (N_9442,N_8823,N_8815);
nor U9443 (N_9443,N_8951,N_8683);
xor U9444 (N_9444,N_8601,N_8836);
and U9445 (N_9445,N_8752,N_8953);
nor U9446 (N_9446,N_8680,N_8731);
nor U9447 (N_9447,N_8562,N_8826);
nor U9448 (N_9448,N_8876,N_8614);
nand U9449 (N_9449,N_8900,N_8625);
or U9450 (N_9450,N_8602,N_8823);
nand U9451 (N_9451,N_8523,N_8654);
xor U9452 (N_9452,N_8629,N_8522);
and U9453 (N_9453,N_8822,N_8651);
and U9454 (N_9454,N_8989,N_8824);
or U9455 (N_9455,N_8959,N_8867);
nor U9456 (N_9456,N_8978,N_8707);
or U9457 (N_9457,N_8601,N_8988);
nand U9458 (N_9458,N_8943,N_8599);
and U9459 (N_9459,N_8541,N_8821);
nand U9460 (N_9460,N_8505,N_8538);
nor U9461 (N_9461,N_8677,N_8693);
and U9462 (N_9462,N_8848,N_8612);
and U9463 (N_9463,N_8672,N_8757);
nand U9464 (N_9464,N_8553,N_8850);
nor U9465 (N_9465,N_8521,N_8709);
nand U9466 (N_9466,N_8534,N_8639);
nand U9467 (N_9467,N_8642,N_8655);
or U9468 (N_9468,N_8578,N_8755);
nand U9469 (N_9469,N_8528,N_8925);
nand U9470 (N_9470,N_8908,N_8566);
and U9471 (N_9471,N_8580,N_8981);
and U9472 (N_9472,N_8500,N_8613);
and U9473 (N_9473,N_8973,N_8660);
or U9474 (N_9474,N_8743,N_8668);
xor U9475 (N_9475,N_8798,N_8659);
and U9476 (N_9476,N_8965,N_8646);
nand U9477 (N_9477,N_8988,N_8757);
xnor U9478 (N_9478,N_8948,N_8954);
nor U9479 (N_9479,N_8517,N_8996);
or U9480 (N_9480,N_8548,N_8529);
xnor U9481 (N_9481,N_8993,N_8793);
nor U9482 (N_9482,N_8745,N_8750);
and U9483 (N_9483,N_8955,N_8712);
nand U9484 (N_9484,N_8748,N_8777);
and U9485 (N_9485,N_8805,N_8563);
and U9486 (N_9486,N_8790,N_8842);
nor U9487 (N_9487,N_8645,N_8862);
nand U9488 (N_9488,N_8792,N_8824);
nand U9489 (N_9489,N_8977,N_8782);
xor U9490 (N_9490,N_8828,N_8543);
and U9491 (N_9491,N_8797,N_8829);
or U9492 (N_9492,N_8681,N_8905);
nand U9493 (N_9493,N_8760,N_8615);
xnor U9494 (N_9494,N_8819,N_8803);
nand U9495 (N_9495,N_8899,N_8566);
and U9496 (N_9496,N_8582,N_8783);
nor U9497 (N_9497,N_8501,N_8559);
nor U9498 (N_9498,N_8557,N_8936);
nand U9499 (N_9499,N_8800,N_8537);
nor U9500 (N_9500,N_9144,N_9455);
or U9501 (N_9501,N_9261,N_9358);
and U9502 (N_9502,N_9330,N_9161);
or U9503 (N_9503,N_9339,N_9220);
and U9504 (N_9504,N_9327,N_9119);
or U9505 (N_9505,N_9242,N_9205);
or U9506 (N_9506,N_9170,N_9422);
and U9507 (N_9507,N_9465,N_9055);
and U9508 (N_9508,N_9185,N_9085);
and U9509 (N_9509,N_9115,N_9298);
nand U9510 (N_9510,N_9370,N_9253);
nand U9511 (N_9511,N_9005,N_9341);
xnor U9512 (N_9512,N_9346,N_9128);
nor U9513 (N_9513,N_9270,N_9223);
or U9514 (N_9514,N_9363,N_9497);
or U9515 (N_9515,N_9340,N_9389);
or U9516 (N_9516,N_9124,N_9351);
nor U9517 (N_9517,N_9458,N_9284);
nand U9518 (N_9518,N_9191,N_9490);
or U9519 (N_9519,N_9256,N_9024);
xor U9520 (N_9520,N_9499,N_9335);
nor U9521 (N_9521,N_9426,N_9186);
and U9522 (N_9522,N_9314,N_9307);
nor U9523 (N_9523,N_9082,N_9381);
or U9524 (N_9524,N_9414,N_9175);
xor U9525 (N_9525,N_9072,N_9084);
nor U9526 (N_9526,N_9195,N_9252);
xor U9527 (N_9527,N_9047,N_9219);
nor U9528 (N_9528,N_9008,N_9086);
nand U9529 (N_9529,N_9123,N_9495);
xor U9530 (N_9530,N_9313,N_9204);
or U9531 (N_9531,N_9125,N_9421);
nand U9532 (N_9532,N_9338,N_9059);
and U9533 (N_9533,N_9294,N_9353);
and U9534 (N_9534,N_9439,N_9143);
and U9535 (N_9535,N_9441,N_9403);
xor U9536 (N_9536,N_9420,N_9491);
and U9537 (N_9537,N_9364,N_9326);
xnor U9538 (N_9538,N_9227,N_9333);
xor U9539 (N_9539,N_9405,N_9266);
and U9540 (N_9540,N_9021,N_9437);
xnor U9541 (N_9541,N_9035,N_9262);
or U9542 (N_9542,N_9336,N_9022);
xnor U9543 (N_9543,N_9231,N_9029);
nor U9544 (N_9544,N_9279,N_9183);
nor U9545 (N_9545,N_9442,N_9129);
nor U9546 (N_9546,N_9423,N_9287);
and U9547 (N_9547,N_9203,N_9462);
and U9548 (N_9548,N_9187,N_9077);
and U9549 (N_9549,N_9352,N_9464);
or U9550 (N_9550,N_9080,N_9017);
and U9551 (N_9551,N_9199,N_9039);
nor U9552 (N_9552,N_9100,N_9359);
nand U9553 (N_9553,N_9131,N_9428);
nand U9554 (N_9554,N_9147,N_9184);
and U9555 (N_9555,N_9344,N_9461);
or U9556 (N_9556,N_9305,N_9165);
nand U9557 (N_9557,N_9474,N_9216);
or U9558 (N_9558,N_9002,N_9498);
nand U9559 (N_9559,N_9054,N_9412);
or U9560 (N_9560,N_9237,N_9214);
and U9561 (N_9561,N_9483,N_9382);
or U9562 (N_9562,N_9137,N_9049);
xnor U9563 (N_9563,N_9297,N_9150);
nand U9564 (N_9564,N_9482,N_9496);
nand U9565 (N_9565,N_9269,N_9056);
nor U9566 (N_9566,N_9471,N_9289);
nand U9567 (N_9567,N_9375,N_9408);
or U9568 (N_9568,N_9145,N_9087);
nor U9569 (N_9569,N_9210,N_9319);
and U9570 (N_9570,N_9361,N_9095);
nor U9571 (N_9571,N_9485,N_9198);
and U9572 (N_9572,N_9241,N_9494);
or U9573 (N_9573,N_9480,N_9406);
nand U9574 (N_9574,N_9309,N_9157);
or U9575 (N_9575,N_9016,N_9174);
and U9576 (N_9576,N_9384,N_9090);
nor U9577 (N_9577,N_9107,N_9043);
xnor U9578 (N_9578,N_9487,N_9169);
or U9579 (N_9579,N_9371,N_9000);
nand U9580 (N_9580,N_9432,N_9083);
nand U9581 (N_9581,N_9078,N_9097);
nor U9582 (N_9582,N_9334,N_9098);
nand U9583 (N_9583,N_9492,N_9250);
nor U9584 (N_9584,N_9099,N_9068);
nor U9585 (N_9585,N_9489,N_9271);
nor U9586 (N_9586,N_9259,N_9139);
and U9587 (N_9587,N_9456,N_9197);
xor U9588 (N_9588,N_9173,N_9444);
xnor U9589 (N_9589,N_9387,N_9181);
and U9590 (N_9590,N_9272,N_9479);
and U9591 (N_9591,N_9239,N_9301);
nor U9592 (N_9592,N_9166,N_9162);
and U9593 (N_9593,N_9019,N_9160);
nand U9594 (N_9594,N_9134,N_9067);
nand U9595 (N_9595,N_9232,N_9106);
xor U9596 (N_9596,N_9202,N_9036);
nand U9597 (N_9597,N_9449,N_9234);
nor U9598 (N_9598,N_9247,N_9006);
or U9599 (N_9599,N_9065,N_9407);
nand U9600 (N_9600,N_9238,N_9276);
and U9601 (N_9601,N_9424,N_9399);
xor U9602 (N_9602,N_9410,N_9188);
nand U9603 (N_9603,N_9329,N_9053);
nand U9604 (N_9604,N_9395,N_9308);
xnor U9605 (N_9605,N_9274,N_9427);
or U9606 (N_9606,N_9117,N_9027);
and U9607 (N_9607,N_9189,N_9208);
nand U9608 (N_9608,N_9240,N_9121);
and U9609 (N_9609,N_9225,N_9295);
or U9610 (N_9610,N_9304,N_9416);
or U9611 (N_9611,N_9419,N_9164);
nand U9612 (N_9612,N_9092,N_9140);
and U9613 (N_9613,N_9267,N_9020);
nor U9614 (N_9614,N_9222,N_9062);
and U9615 (N_9615,N_9322,N_9376);
nor U9616 (N_9616,N_9317,N_9470);
and U9617 (N_9617,N_9343,N_9118);
and U9618 (N_9618,N_9292,N_9218);
and U9619 (N_9619,N_9443,N_9264);
xnor U9620 (N_9620,N_9433,N_9221);
nor U9621 (N_9621,N_9349,N_9094);
nor U9622 (N_9622,N_9026,N_9200);
and U9623 (N_9623,N_9025,N_9023);
nor U9624 (N_9624,N_9152,N_9321);
nor U9625 (N_9625,N_9457,N_9466);
nand U9626 (N_9626,N_9409,N_9473);
nand U9627 (N_9627,N_9122,N_9453);
or U9628 (N_9628,N_9211,N_9101);
or U9629 (N_9629,N_9212,N_9451);
and U9630 (N_9630,N_9469,N_9070);
nand U9631 (N_9631,N_9445,N_9369);
and U9632 (N_9632,N_9088,N_9037);
or U9633 (N_9633,N_9396,N_9255);
or U9634 (N_9634,N_9004,N_9064);
nor U9635 (N_9635,N_9076,N_9235);
xnor U9636 (N_9636,N_9111,N_9277);
nand U9637 (N_9637,N_9293,N_9377);
or U9638 (N_9638,N_9034,N_9438);
and U9639 (N_9639,N_9324,N_9477);
xnor U9640 (N_9640,N_9285,N_9430);
nor U9641 (N_9641,N_9354,N_9296);
or U9642 (N_9642,N_9397,N_9440);
nand U9643 (N_9643,N_9112,N_9075);
or U9644 (N_9644,N_9215,N_9435);
nor U9645 (N_9645,N_9050,N_9394);
or U9646 (N_9646,N_9138,N_9400);
or U9647 (N_9647,N_9013,N_9282);
and U9648 (N_9648,N_9182,N_9290);
nand U9649 (N_9649,N_9081,N_9207);
or U9650 (N_9650,N_9052,N_9378);
and U9651 (N_9651,N_9233,N_9246);
or U9652 (N_9652,N_9116,N_9044);
nand U9653 (N_9653,N_9136,N_9429);
nor U9654 (N_9654,N_9383,N_9127);
nor U9655 (N_9655,N_9374,N_9318);
and U9656 (N_9656,N_9196,N_9133);
nor U9657 (N_9657,N_9245,N_9066);
nor U9658 (N_9658,N_9130,N_9177);
and U9659 (N_9659,N_9108,N_9488);
xor U9660 (N_9660,N_9385,N_9347);
or U9661 (N_9661,N_9051,N_9171);
or U9662 (N_9662,N_9091,N_9159);
xnor U9663 (N_9663,N_9254,N_9096);
and U9664 (N_9664,N_9060,N_9434);
xnor U9665 (N_9665,N_9209,N_9486);
nor U9666 (N_9666,N_9398,N_9142);
or U9667 (N_9667,N_9265,N_9342);
and U9668 (N_9668,N_9328,N_9413);
nor U9669 (N_9669,N_9467,N_9356);
xnor U9670 (N_9670,N_9459,N_9010);
nor U9671 (N_9671,N_9436,N_9217);
nand U9672 (N_9672,N_9153,N_9074);
nand U9673 (N_9673,N_9114,N_9190);
xnor U9674 (N_9674,N_9109,N_9493);
nor U9675 (N_9675,N_9236,N_9325);
or U9676 (N_9676,N_9275,N_9355);
and U9677 (N_9677,N_9368,N_9404);
xnor U9678 (N_9678,N_9448,N_9417);
and U9679 (N_9679,N_9316,N_9300);
or U9680 (N_9680,N_9367,N_9093);
and U9681 (N_9681,N_9001,N_9251);
nand U9682 (N_9682,N_9257,N_9155);
and U9683 (N_9683,N_9201,N_9156);
nor U9684 (N_9684,N_9167,N_9079);
xor U9685 (N_9685,N_9362,N_9149);
nand U9686 (N_9686,N_9393,N_9105);
and U9687 (N_9687,N_9281,N_9332);
nor U9688 (N_9688,N_9447,N_9380);
or U9689 (N_9689,N_9303,N_9391);
xor U9690 (N_9690,N_9452,N_9366);
and U9691 (N_9691,N_9402,N_9249);
xor U9692 (N_9692,N_9041,N_9230);
and U9693 (N_9693,N_9446,N_9348);
xnor U9694 (N_9694,N_9014,N_9280);
or U9695 (N_9695,N_9323,N_9315);
nand U9696 (N_9696,N_9045,N_9038);
nand U9697 (N_9697,N_9379,N_9450);
and U9698 (N_9698,N_9015,N_9168);
nand U9699 (N_9699,N_9286,N_9320);
xor U9700 (N_9700,N_9063,N_9089);
and U9701 (N_9701,N_9263,N_9350);
and U9702 (N_9702,N_9229,N_9312);
nand U9703 (N_9703,N_9331,N_9151);
xnor U9704 (N_9704,N_9360,N_9372);
nand U9705 (N_9705,N_9057,N_9146);
or U9706 (N_9706,N_9048,N_9302);
nand U9707 (N_9707,N_9418,N_9102);
nand U9708 (N_9708,N_9104,N_9386);
and U9709 (N_9709,N_9311,N_9390);
or U9710 (N_9710,N_9180,N_9031);
and U9711 (N_9711,N_9179,N_9030);
nand U9712 (N_9712,N_9268,N_9206);
nand U9713 (N_9713,N_9345,N_9365);
or U9714 (N_9714,N_9310,N_9283);
or U9715 (N_9715,N_9481,N_9042);
and U9716 (N_9716,N_9046,N_9357);
and U9717 (N_9717,N_9244,N_9454);
nor U9718 (N_9718,N_9463,N_9178);
nand U9719 (N_9719,N_9018,N_9103);
or U9720 (N_9720,N_9192,N_9172);
and U9721 (N_9721,N_9411,N_9132);
nand U9722 (N_9722,N_9032,N_9299);
or U9723 (N_9723,N_9478,N_9135);
nand U9724 (N_9724,N_9278,N_9388);
nor U9725 (N_9725,N_9069,N_9154);
or U9726 (N_9726,N_9392,N_9040);
nor U9727 (N_9727,N_9472,N_9260);
nor U9728 (N_9728,N_9071,N_9009);
or U9729 (N_9729,N_9415,N_9126);
and U9730 (N_9730,N_9163,N_9224);
or U9731 (N_9731,N_9373,N_9061);
or U9732 (N_9732,N_9003,N_9337);
nor U9733 (N_9733,N_9248,N_9158);
and U9734 (N_9734,N_9058,N_9228);
and U9735 (N_9735,N_9258,N_9007);
nand U9736 (N_9736,N_9193,N_9141);
xnor U9737 (N_9737,N_9468,N_9028);
or U9738 (N_9738,N_9012,N_9288);
or U9739 (N_9739,N_9033,N_9273);
or U9740 (N_9740,N_9425,N_9306);
or U9741 (N_9741,N_9291,N_9484);
nor U9742 (N_9742,N_9176,N_9460);
and U9743 (N_9743,N_9110,N_9148);
xor U9744 (N_9744,N_9073,N_9475);
and U9745 (N_9745,N_9401,N_9226);
or U9746 (N_9746,N_9243,N_9194);
nor U9747 (N_9747,N_9431,N_9120);
or U9748 (N_9748,N_9113,N_9213);
nor U9749 (N_9749,N_9011,N_9476);
and U9750 (N_9750,N_9223,N_9357);
and U9751 (N_9751,N_9064,N_9001);
nand U9752 (N_9752,N_9066,N_9132);
nor U9753 (N_9753,N_9452,N_9288);
nor U9754 (N_9754,N_9027,N_9026);
and U9755 (N_9755,N_9441,N_9443);
and U9756 (N_9756,N_9079,N_9188);
and U9757 (N_9757,N_9330,N_9416);
and U9758 (N_9758,N_9455,N_9200);
nor U9759 (N_9759,N_9253,N_9127);
nand U9760 (N_9760,N_9045,N_9452);
and U9761 (N_9761,N_9437,N_9010);
nor U9762 (N_9762,N_9499,N_9468);
nor U9763 (N_9763,N_9370,N_9115);
and U9764 (N_9764,N_9148,N_9218);
nor U9765 (N_9765,N_9117,N_9178);
and U9766 (N_9766,N_9483,N_9372);
xor U9767 (N_9767,N_9398,N_9299);
xor U9768 (N_9768,N_9199,N_9276);
nor U9769 (N_9769,N_9126,N_9296);
nor U9770 (N_9770,N_9263,N_9486);
nand U9771 (N_9771,N_9015,N_9472);
xnor U9772 (N_9772,N_9213,N_9479);
xor U9773 (N_9773,N_9130,N_9175);
or U9774 (N_9774,N_9142,N_9408);
xnor U9775 (N_9775,N_9003,N_9042);
or U9776 (N_9776,N_9050,N_9470);
or U9777 (N_9777,N_9448,N_9447);
and U9778 (N_9778,N_9496,N_9295);
or U9779 (N_9779,N_9282,N_9167);
nand U9780 (N_9780,N_9406,N_9098);
xor U9781 (N_9781,N_9117,N_9366);
and U9782 (N_9782,N_9441,N_9438);
nand U9783 (N_9783,N_9407,N_9071);
or U9784 (N_9784,N_9345,N_9287);
nor U9785 (N_9785,N_9052,N_9003);
or U9786 (N_9786,N_9351,N_9242);
xor U9787 (N_9787,N_9448,N_9222);
xor U9788 (N_9788,N_9407,N_9037);
or U9789 (N_9789,N_9106,N_9228);
and U9790 (N_9790,N_9214,N_9412);
or U9791 (N_9791,N_9203,N_9443);
nand U9792 (N_9792,N_9184,N_9376);
nand U9793 (N_9793,N_9017,N_9448);
xnor U9794 (N_9794,N_9482,N_9190);
xor U9795 (N_9795,N_9463,N_9110);
and U9796 (N_9796,N_9017,N_9465);
xor U9797 (N_9797,N_9094,N_9410);
nor U9798 (N_9798,N_9308,N_9209);
or U9799 (N_9799,N_9353,N_9158);
and U9800 (N_9800,N_9363,N_9139);
and U9801 (N_9801,N_9415,N_9041);
nand U9802 (N_9802,N_9273,N_9378);
or U9803 (N_9803,N_9077,N_9072);
nand U9804 (N_9804,N_9101,N_9047);
nor U9805 (N_9805,N_9483,N_9026);
or U9806 (N_9806,N_9099,N_9293);
xor U9807 (N_9807,N_9041,N_9383);
and U9808 (N_9808,N_9306,N_9360);
xnor U9809 (N_9809,N_9409,N_9120);
and U9810 (N_9810,N_9402,N_9371);
nand U9811 (N_9811,N_9488,N_9368);
nand U9812 (N_9812,N_9424,N_9395);
and U9813 (N_9813,N_9207,N_9396);
nor U9814 (N_9814,N_9193,N_9239);
and U9815 (N_9815,N_9495,N_9061);
nand U9816 (N_9816,N_9422,N_9205);
nand U9817 (N_9817,N_9084,N_9499);
or U9818 (N_9818,N_9370,N_9118);
and U9819 (N_9819,N_9473,N_9053);
and U9820 (N_9820,N_9040,N_9257);
xnor U9821 (N_9821,N_9226,N_9175);
and U9822 (N_9822,N_9121,N_9120);
and U9823 (N_9823,N_9429,N_9319);
or U9824 (N_9824,N_9338,N_9431);
xor U9825 (N_9825,N_9330,N_9455);
nand U9826 (N_9826,N_9325,N_9200);
nand U9827 (N_9827,N_9015,N_9005);
nand U9828 (N_9828,N_9262,N_9026);
nor U9829 (N_9829,N_9243,N_9199);
or U9830 (N_9830,N_9088,N_9392);
nand U9831 (N_9831,N_9305,N_9308);
and U9832 (N_9832,N_9013,N_9310);
nor U9833 (N_9833,N_9132,N_9069);
nor U9834 (N_9834,N_9159,N_9337);
nand U9835 (N_9835,N_9065,N_9234);
nor U9836 (N_9836,N_9100,N_9437);
and U9837 (N_9837,N_9487,N_9301);
nand U9838 (N_9838,N_9431,N_9091);
nor U9839 (N_9839,N_9122,N_9274);
xnor U9840 (N_9840,N_9149,N_9085);
nor U9841 (N_9841,N_9182,N_9189);
and U9842 (N_9842,N_9177,N_9384);
xor U9843 (N_9843,N_9179,N_9208);
nand U9844 (N_9844,N_9436,N_9259);
and U9845 (N_9845,N_9146,N_9121);
nand U9846 (N_9846,N_9254,N_9466);
nand U9847 (N_9847,N_9289,N_9031);
or U9848 (N_9848,N_9358,N_9214);
xnor U9849 (N_9849,N_9138,N_9447);
and U9850 (N_9850,N_9241,N_9132);
xor U9851 (N_9851,N_9040,N_9024);
and U9852 (N_9852,N_9147,N_9224);
nor U9853 (N_9853,N_9171,N_9435);
nand U9854 (N_9854,N_9327,N_9303);
xor U9855 (N_9855,N_9391,N_9163);
xor U9856 (N_9856,N_9304,N_9279);
nor U9857 (N_9857,N_9307,N_9320);
or U9858 (N_9858,N_9177,N_9036);
and U9859 (N_9859,N_9274,N_9347);
or U9860 (N_9860,N_9405,N_9156);
nor U9861 (N_9861,N_9484,N_9046);
nand U9862 (N_9862,N_9493,N_9265);
xnor U9863 (N_9863,N_9237,N_9092);
or U9864 (N_9864,N_9242,N_9342);
and U9865 (N_9865,N_9401,N_9024);
nor U9866 (N_9866,N_9032,N_9269);
xor U9867 (N_9867,N_9016,N_9361);
xnor U9868 (N_9868,N_9091,N_9350);
xor U9869 (N_9869,N_9059,N_9008);
and U9870 (N_9870,N_9028,N_9179);
nand U9871 (N_9871,N_9152,N_9085);
nor U9872 (N_9872,N_9026,N_9168);
nand U9873 (N_9873,N_9412,N_9233);
and U9874 (N_9874,N_9405,N_9182);
nand U9875 (N_9875,N_9276,N_9171);
or U9876 (N_9876,N_9193,N_9396);
or U9877 (N_9877,N_9475,N_9023);
nor U9878 (N_9878,N_9236,N_9091);
or U9879 (N_9879,N_9063,N_9033);
xor U9880 (N_9880,N_9239,N_9230);
nand U9881 (N_9881,N_9076,N_9381);
or U9882 (N_9882,N_9442,N_9464);
xnor U9883 (N_9883,N_9217,N_9450);
xor U9884 (N_9884,N_9004,N_9235);
nand U9885 (N_9885,N_9350,N_9430);
nor U9886 (N_9886,N_9132,N_9111);
nand U9887 (N_9887,N_9425,N_9287);
xnor U9888 (N_9888,N_9230,N_9148);
nand U9889 (N_9889,N_9133,N_9205);
nand U9890 (N_9890,N_9059,N_9158);
nor U9891 (N_9891,N_9069,N_9025);
and U9892 (N_9892,N_9309,N_9362);
nor U9893 (N_9893,N_9276,N_9390);
and U9894 (N_9894,N_9444,N_9079);
and U9895 (N_9895,N_9110,N_9006);
or U9896 (N_9896,N_9150,N_9134);
and U9897 (N_9897,N_9293,N_9170);
xor U9898 (N_9898,N_9448,N_9436);
nand U9899 (N_9899,N_9301,N_9037);
and U9900 (N_9900,N_9173,N_9419);
or U9901 (N_9901,N_9270,N_9235);
or U9902 (N_9902,N_9020,N_9493);
nor U9903 (N_9903,N_9488,N_9449);
nor U9904 (N_9904,N_9300,N_9083);
or U9905 (N_9905,N_9083,N_9177);
and U9906 (N_9906,N_9457,N_9186);
nand U9907 (N_9907,N_9233,N_9480);
nand U9908 (N_9908,N_9349,N_9097);
and U9909 (N_9909,N_9361,N_9346);
nand U9910 (N_9910,N_9195,N_9241);
nor U9911 (N_9911,N_9210,N_9185);
and U9912 (N_9912,N_9322,N_9065);
or U9913 (N_9913,N_9156,N_9080);
and U9914 (N_9914,N_9293,N_9265);
or U9915 (N_9915,N_9124,N_9289);
xor U9916 (N_9916,N_9308,N_9368);
nor U9917 (N_9917,N_9188,N_9475);
or U9918 (N_9918,N_9456,N_9173);
and U9919 (N_9919,N_9268,N_9117);
nand U9920 (N_9920,N_9486,N_9396);
xor U9921 (N_9921,N_9125,N_9299);
nor U9922 (N_9922,N_9464,N_9313);
and U9923 (N_9923,N_9463,N_9290);
nand U9924 (N_9924,N_9024,N_9389);
xor U9925 (N_9925,N_9330,N_9118);
nand U9926 (N_9926,N_9139,N_9434);
nor U9927 (N_9927,N_9125,N_9431);
xor U9928 (N_9928,N_9407,N_9095);
nand U9929 (N_9929,N_9136,N_9047);
and U9930 (N_9930,N_9150,N_9475);
and U9931 (N_9931,N_9331,N_9049);
xnor U9932 (N_9932,N_9177,N_9379);
nand U9933 (N_9933,N_9161,N_9203);
nor U9934 (N_9934,N_9369,N_9106);
or U9935 (N_9935,N_9162,N_9214);
nand U9936 (N_9936,N_9420,N_9463);
nor U9937 (N_9937,N_9041,N_9281);
xor U9938 (N_9938,N_9410,N_9065);
or U9939 (N_9939,N_9354,N_9037);
nor U9940 (N_9940,N_9350,N_9413);
and U9941 (N_9941,N_9225,N_9145);
or U9942 (N_9942,N_9028,N_9122);
nor U9943 (N_9943,N_9327,N_9417);
xnor U9944 (N_9944,N_9215,N_9090);
nor U9945 (N_9945,N_9175,N_9454);
xnor U9946 (N_9946,N_9440,N_9236);
nor U9947 (N_9947,N_9151,N_9247);
xor U9948 (N_9948,N_9007,N_9092);
nor U9949 (N_9949,N_9496,N_9301);
xnor U9950 (N_9950,N_9300,N_9261);
or U9951 (N_9951,N_9084,N_9429);
xnor U9952 (N_9952,N_9075,N_9209);
xor U9953 (N_9953,N_9213,N_9460);
nor U9954 (N_9954,N_9305,N_9137);
xnor U9955 (N_9955,N_9368,N_9455);
or U9956 (N_9956,N_9307,N_9388);
nor U9957 (N_9957,N_9008,N_9307);
nor U9958 (N_9958,N_9010,N_9300);
xor U9959 (N_9959,N_9383,N_9325);
xor U9960 (N_9960,N_9015,N_9021);
xnor U9961 (N_9961,N_9435,N_9244);
and U9962 (N_9962,N_9298,N_9294);
and U9963 (N_9963,N_9457,N_9242);
nor U9964 (N_9964,N_9497,N_9322);
nor U9965 (N_9965,N_9491,N_9164);
nand U9966 (N_9966,N_9096,N_9426);
nand U9967 (N_9967,N_9303,N_9395);
nor U9968 (N_9968,N_9095,N_9050);
or U9969 (N_9969,N_9200,N_9429);
nand U9970 (N_9970,N_9335,N_9407);
xor U9971 (N_9971,N_9312,N_9181);
and U9972 (N_9972,N_9231,N_9224);
nor U9973 (N_9973,N_9479,N_9296);
or U9974 (N_9974,N_9411,N_9338);
or U9975 (N_9975,N_9070,N_9388);
nor U9976 (N_9976,N_9456,N_9137);
nand U9977 (N_9977,N_9408,N_9002);
nor U9978 (N_9978,N_9393,N_9426);
xor U9979 (N_9979,N_9311,N_9249);
xor U9980 (N_9980,N_9066,N_9362);
and U9981 (N_9981,N_9107,N_9265);
xor U9982 (N_9982,N_9475,N_9435);
xnor U9983 (N_9983,N_9346,N_9375);
or U9984 (N_9984,N_9281,N_9304);
xor U9985 (N_9985,N_9064,N_9017);
xor U9986 (N_9986,N_9320,N_9204);
or U9987 (N_9987,N_9450,N_9406);
or U9988 (N_9988,N_9338,N_9361);
or U9989 (N_9989,N_9188,N_9132);
xor U9990 (N_9990,N_9403,N_9318);
or U9991 (N_9991,N_9126,N_9451);
or U9992 (N_9992,N_9142,N_9258);
nand U9993 (N_9993,N_9123,N_9141);
nor U9994 (N_9994,N_9420,N_9067);
and U9995 (N_9995,N_9147,N_9320);
nor U9996 (N_9996,N_9278,N_9404);
and U9997 (N_9997,N_9152,N_9197);
xnor U9998 (N_9998,N_9384,N_9168);
xnor U9999 (N_9999,N_9036,N_9290);
xor U10000 (N_10000,N_9892,N_9883);
and U10001 (N_10001,N_9730,N_9561);
nand U10002 (N_10002,N_9682,N_9620);
or U10003 (N_10003,N_9797,N_9528);
and U10004 (N_10004,N_9980,N_9676);
and U10005 (N_10005,N_9681,N_9816);
and U10006 (N_10006,N_9568,N_9867);
or U10007 (N_10007,N_9667,N_9661);
nand U10008 (N_10008,N_9593,N_9887);
nor U10009 (N_10009,N_9830,N_9984);
nand U10010 (N_10010,N_9594,N_9734);
xnor U10011 (N_10011,N_9741,N_9928);
xnor U10012 (N_10012,N_9759,N_9587);
nor U10013 (N_10013,N_9680,N_9601);
xor U10014 (N_10014,N_9709,N_9787);
nand U10015 (N_10015,N_9881,N_9904);
xnor U10016 (N_10016,N_9882,N_9855);
and U10017 (N_10017,N_9534,N_9965);
and U10018 (N_10018,N_9754,N_9813);
nand U10019 (N_10019,N_9505,N_9862);
nand U10020 (N_10020,N_9993,N_9599);
nand U10021 (N_10021,N_9654,N_9686);
and U10022 (N_10022,N_9523,N_9755);
nor U10023 (N_10023,N_9874,N_9857);
xnor U10024 (N_10024,N_9538,N_9610);
nor U10025 (N_10025,N_9588,N_9564);
nand U10026 (N_10026,N_9912,N_9600);
nor U10027 (N_10027,N_9578,N_9995);
xor U10028 (N_10028,N_9781,N_9604);
and U10029 (N_10029,N_9915,N_9548);
and U10030 (N_10030,N_9689,N_9591);
nand U10031 (N_10031,N_9553,N_9959);
nand U10032 (N_10032,N_9868,N_9585);
xor U10033 (N_10033,N_9770,N_9836);
or U10034 (N_10034,N_9865,N_9786);
or U10035 (N_10035,N_9590,N_9990);
xnor U10036 (N_10036,N_9618,N_9721);
xnor U10037 (N_10037,N_9640,N_9695);
nor U10038 (N_10038,N_9964,N_9562);
and U10039 (N_10039,N_9545,N_9525);
nand U10040 (N_10040,N_9806,N_9979);
and U10041 (N_10041,N_9827,N_9924);
nand U10042 (N_10042,N_9753,N_9624);
nand U10043 (N_10043,N_9670,N_9758);
or U10044 (N_10044,N_9611,N_9856);
nor U10045 (N_10045,N_9608,N_9744);
nand U10046 (N_10046,N_9947,N_9869);
nor U10047 (N_10047,N_9605,N_9782);
and U10048 (N_10048,N_9650,N_9555);
nor U10049 (N_10049,N_9972,N_9699);
nand U10050 (N_10050,N_9771,N_9537);
or U10051 (N_10051,N_9802,N_9898);
and U10052 (N_10052,N_9678,N_9655);
or U10053 (N_10053,N_9844,N_9981);
nand U10054 (N_10054,N_9825,N_9668);
nor U10055 (N_10055,N_9873,N_9596);
nand U10056 (N_10056,N_9834,N_9745);
or U10057 (N_10057,N_9509,N_9902);
or U10058 (N_10058,N_9589,N_9549);
xnor U10059 (N_10059,N_9581,N_9765);
nor U10060 (N_10060,N_9629,N_9570);
or U10061 (N_10061,N_9943,N_9824);
nor U10062 (N_10062,N_9942,N_9918);
nand U10063 (N_10063,N_9921,N_9798);
nor U10064 (N_10064,N_9733,N_9949);
xnor U10065 (N_10065,N_9841,N_9506);
nand U10066 (N_10066,N_9653,N_9615);
nand U10067 (N_10067,N_9876,N_9580);
and U10068 (N_10068,N_9514,N_9634);
or U10069 (N_10069,N_9630,N_9783);
nor U10070 (N_10070,N_9749,N_9905);
xor U10071 (N_10071,N_9829,N_9767);
xor U10072 (N_10072,N_9565,N_9930);
or U10073 (N_10073,N_9953,N_9810);
nand U10074 (N_10074,N_9792,N_9890);
xnor U10075 (N_10075,N_9598,N_9584);
and U10076 (N_10076,N_9974,N_9919);
xor U10077 (N_10077,N_9547,N_9609);
nand U10078 (N_10078,N_9888,N_9662);
nor U10079 (N_10079,N_9842,N_9831);
and U10080 (N_10080,N_9633,N_9835);
and U10081 (N_10081,N_9986,N_9795);
xor U10082 (N_10082,N_9780,N_9536);
xnor U10083 (N_10083,N_9860,N_9625);
nand U10084 (N_10084,N_9966,N_9760);
and U10085 (N_10085,N_9688,N_9567);
xnor U10086 (N_10086,N_9926,N_9501);
and U10087 (N_10087,N_9697,N_9871);
or U10088 (N_10088,N_9727,N_9948);
xnor U10089 (N_10089,N_9722,N_9804);
nand U10090 (N_10090,N_9794,N_9612);
nand U10091 (N_10091,N_9907,N_9576);
nor U10092 (N_10092,N_9788,N_9544);
and U10093 (N_10093,N_9910,N_9691);
nor U10094 (N_10094,N_9517,N_9546);
xnor U10095 (N_10095,N_9657,N_9763);
xor U10096 (N_10096,N_9955,N_9996);
nor U10097 (N_10097,N_9896,N_9616);
and U10098 (N_10098,N_9775,N_9673);
nand U10099 (N_10099,N_9789,N_9854);
nor U10100 (N_10100,N_9696,N_9558);
and U10101 (N_10101,N_9838,N_9597);
xnor U10102 (N_10102,N_9756,N_9706);
xnor U10103 (N_10103,N_9714,N_9790);
nor U10104 (N_10104,N_9694,N_9901);
and U10105 (N_10105,N_9863,N_9672);
nor U10106 (N_10106,N_9885,N_9840);
xor U10107 (N_10107,N_9539,N_9929);
xnor U10108 (N_10108,N_9791,N_9743);
or U10109 (N_10109,N_9807,N_9524);
nand U10110 (N_10110,N_9645,N_9847);
nand U10111 (N_10111,N_9951,N_9870);
or U10112 (N_10112,N_9939,N_9977);
nand U10113 (N_10113,N_9636,N_9535);
and U10114 (N_10114,N_9988,N_9732);
nor U10115 (N_10115,N_9515,N_9726);
and U10116 (N_10116,N_9805,N_9626);
xor U10117 (N_10117,N_9768,N_9849);
and U10118 (N_10118,N_9803,N_9531);
and U10119 (N_10119,N_9989,N_9675);
and U10120 (N_10120,N_9917,N_9851);
or U10121 (N_10121,N_9529,N_9652);
nor U10122 (N_10122,N_9913,N_9684);
nor U10123 (N_10123,N_9521,N_9583);
and U10124 (N_10124,N_9976,N_9693);
or U10125 (N_10125,N_9961,N_9925);
nor U10126 (N_10126,N_9957,N_9540);
nand U10127 (N_10127,N_9735,N_9648);
nand U10128 (N_10128,N_9837,N_9508);
nand U10129 (N_10129,N_9846,N_9718);
xnor U10130 (N_10130,N_9592,N_9542);
xnor U10131 (N_10131,N_9705,N_9513);
nor U10132 (N_10132,N_9731,N_9569);
and U10133 (N_10133,N_9516,N_9893);
nor U10134 (N_10134,N_9911,N_9701);
nor U10135 (N_10135,N_9659,N_9715);
nor U10136 (N_10136,N_9526,N_9503);
or U10137 (N_10137,N_9700,N_9663);
nand U10138 (N_10138,N_9574,N_9669);
xor U10139 (N_10139,N_9878,N_9941);
or U10140 (N_10140,N_9889,N_9757);
nor U10141 (N_10141,N_9761,N_9665);
nand U10142 (N_10142,N_9906,N_9845);
or U10143 (N_10143,N_9677,N_9541);
xnor U10144 (N_10144,N_9935,N_9774);
nand U10145 (N_10145,N_9982,N_9821);
nand U10146 (N_10146,N_9850,N_9692);
and U10147 (N_10147,N_9660,N_9817);
nor U10148 (N_10148,N_9704,N_9617);
and U10149 (N_10149,N_9968,N_9772);
and U10150 (N_10150,N_9656,N_9740);
nor U10151 (N_10151,N_9796,N_9738);
nand U10152 (N_10152,N_9960,N_9725);
or U10153 (N_10153,N_9713,N_9962);
or U10154 (N_10154,N_9751,N_9853);
xor U10155 (N_10155,N_9637,N_9970);
nor U10156 (N_10156,N_9776,N_9698);
xnor U10157 (N_10157,N_9666,N_9823);
nor U10158 (N_10158,N_9766,N_9644);
or U10159 (N_10159,N_9945,N_9720);
and U10160 (N_10160,N_9631,N_9595);
nor U10161 (N_10161,N_9500,N_9674);
and U10162 (N_10162,N_9658,N_9764);
nor U10163 (N_10163,N_9543,N_9784);
xor U10164 (N_10164,N_9808,N_9978);
xnor U10165 (N_10165,N_9512,N_9839);
xor U10166 (N_10166,N_9891,N_9724);
nand U10167 (N_10167,N_9762,N_9779);
or U10168 (N_10168,N_9914,N_9958);
xnor U10169 (N_10169,N_9967,N_9582);
and U10170 (N_10170,N_9622,N_9687);
and U10171 (N_10171,N_9572,N_9818);
and U10172 (N_10172,N_9703,N_9712);
or U10173 (N_10173,N_9502,N_9985);
and U10174 (N_10174,N_9785,N_9638);
nor U10175 (N_10175,N_9533,N_9559);
xor U10176 (N_10176,N_9899,N_9801);
nor U10177 (N_10177,N_9671,N_9998);
nor U10178 (N_10178,N_9932,N_9809);
nor U10179 (N_10179,N_9864,N_9510);
nand U10180 (N_10180,N_9866,N_9938);
nor U10181 (N_10181,N_9623,N_9822);
xnor U10182 (N_10182,N_9635,N_9552);
nand U10183 (N_10183,N_9799,N_9518);
and U10184 (N_10184,N_9550,N_9683);
and U10185 (N_10185,N_9628,N_9880);
or U10186 (N_10186,N_9936,N_9973);
nor U10187 (N_10187,N_9619,N_9646);
nand U10188 (N_10188,N_9532,N_9952);
nand U10189 (N_10189,N_9923,N_9828);
xnor U10190 (N_10190,N_9560,N_9520);
nand U10191 (N_10191,N_9852,N_9614);
xnor U10192 (N_10192,N_9997,N_9971);
nand U10193 (N_10193,N_9859,N_9641);
xor U10194 (N_10194,N_9969,N_9579);
and U10195 (N_10195,N_9750,N_9563);
and U10196 (N_10196,N_9833,N_9994);
or U10197 (N_10197,N_9729,N_9877);
and U10198 (N_10198,N_9607,N_9963);
or U10199 (N_10199,N_9651,N_9747);
xor U10200 (N_10200,N_9717,N_9946);
or U10201 (N_10201,N_9944,N_9664);
xor U10202 (N_10202,N_9507,N_9987);
xor U10203 (N_10203,N_9642,N_9602);
and U10204 (N_10204,N_9940,N_9800);
or U10205 (N_10205,N_9954,N_9778);
or U10206 (N_10206,N_9711,N_9530);
and U10207 (N_10207,N_9903,N_9793);
nor U10208 (N_10208,N_9922,N_9848);
and U10209 (N_10209,N_9649,N_9639);
nand U10210 (N_10210,N_9820,N_9557);
nor U10211 (N_10211,N_9769,N_9736);
or U10212 (N_10212,N_9685,N_9707);
nor U10213 (N_10213,N_9690,N_9723);
or U10214 (N_10214,N_9708,N_9937);
and U10215 (N_10215,N_9613,N_9647);
nand U10216 (N_10216,N_9934,N_9742);
nand U10217 (N_10217,N_9746,N_9702);
xnor U10218 (N_10218,N_9643,N_9737);
or U10219 (N_10219,N_9504,N_9527);
and U10220 (N_10220,N_9992,N_9861);
or U10221 (N_10221,N_9627,N_9843);
xor U10222 (N_10222,N_9522,N_9777);
nand U10223 (N_10223,N_9920,N_9511);
xnor U10224 (N_10224,N_9897,N_9900);
nand U10225 (N_10225,N_9950,N_9710);
nor U10226 (N_10226,N_9752,N_9975);
or U10227 (N_10227,N_9956,N_9815);
or U10228 (N_10228,N_9575,N_9916);
xor U10229 (N_10229,N_9748,N_9879);
nor U10230 (N_10230,N_9551,N_9983);
or U10231 (N_10231,N_9716,N_9773);
and U10232 (N_10232,N_9573,N_9875);
nand U10233 (N_10233,N_9933,N_9931);
nand U10234 (N_10234,N_9872,N_9719);
xor U10235 (N_10235,N_9999,N_9858);
and U10236 (N_10236,N_9577,N_9679);
nor U10237 (N_10237,N_9556,N_9908);
nand U10238 (N_10238,N_9991,N_9571);
nand U10239 (N_10239,N_9566,N_9621);
nor U10240 (N_10240,N_9909,N_9895);
xor U10241 (N_10241,N_9606,N_9927);
and U10242 (N_10242,N_9586,N_9812);
nand U10243 (N_10243,N_9894,N_9739);
or U10244 (N_10244,N_9884,N_9554);
nor U10245 (N_10245,N_9811,N_9603);
xor U10246 (N_10246,N_9814,N_9819);
nor U10247 (N_10247,N_9826,N_9832);
nand U10248 (N_10248,N_9632,N_9728);
or U10249 (N_10249,N_9519,N_9886);
or U10250 (N_10250,N_9812,N_9931);
nor U10251 (N_10251,N_9628,N_9770);
nor U10252 (N_10252,N_9626,N_9831);
nand U10253 (N_10253,N_9961,N_9544);
and U10254 (N_10254,N_9575,N_9542);
nor U10255 (N_10255,N_9944,N_9538);
and U10256 (N_10256,N_9576,N_9667);
nand U10257 (N_10257,N_9762,N_9711);
nor U10258 (N_10258,N_9988,N_9663);
or U10259 (N_10259,N_9579,N_9736);
nand U10260 (N_10260,N_9701,N_9609);
or U10261 (N_10261,N_9681,N_9926);
nor U10262 (N_10262,N_9647,N_9704);
nand U10263 (N_10263,N_9620,N_9554);
or U10264 (N_10264,N_9739,N_9727);
nand U10265 (N_10265,N_9929,N_9726);
and U10266 (N_10266,N_9991,N_9633);
nor U10267 (N_10267,N_9932,N_9997);
xor U10268 (N_10268,N_9619,N_9831);
or U10269 (N_10269,N_9977,N_9988);
xor U10270 (N_10270,N_9597,N_9734);
xnor U10271 (N_10271,N_9920,N_9625);
nand U10272 (N_10272,N_9868,N_9549);
nand U10273 (N_10273,N_9858,N_9586);
xor U10274 (N_10274,N_9692,N_9866);
and U10275 (N_10275,N_9975,N_9631);
nand U10276 (N_10276,N_9958,N_9919);
and U10277 (N_10277,N_9898,N_9812);
or U10278 (N_10278,N_9637,N_9965);
or U10279 (N_10279,N_9773,N_9634);
or U10280 (N_10280,N_9724,N_9794);
and U10281 (N_10281,N_9965,N_9570);
nand U10282 (N_10282,N_9729,N_9535);
nand U10283 (N_10283,N_9754,N_9881);
or U10284 (N_10284,N_9964,N_9904);
nand U10285 (N_10285,N_9738,N_9967);
or U10286 (N_10286,N_9595,N_9906);
nand U10287 (N_10287,N_9947,N_9649);
or U10288 (N_10288,N_9523,N_9628);
nor U10289 (N_10289,N_9536,N_9945);
nor U10290 (N_10290,N_9834,N_9821);
or U10291 (N_10291,N_9614,N_9891);
and U10292 (N_10292,N_9957,N_9680);
xor U10293 (N_10293,N_9952,N_9980);
nor U10294 (N_10294,N_9752,N_9882);
and U10295 (N_10295,N_9879,N_9706);
nand U10296 (N_10296,N_9806,N_9929);
nor U10297 (N_10297,N_9511,N_9753);
or U10298 (N_10298,N_9584,N_9569);
nand U10299 (N_10299,N_9897,N_9760);
or U10300 (N_10300,N_9933,N_9949);
xor U10301 (N_10301,N_9623,N_9897);
and U10302 (N_10302,N_9799,N_9678);
or U10303 (N_10303,N_9730,N_9525);
nand U10304 (N_10304,N_9653,N_9616);
nor U10305 (N_10305,N_9939,N_9732);
and U10306 (N_10306,N_9538,N_9892);
xnor U10307 (N_10307,N_9760,N_9538);
or U10308 (N_10308,N_9784,N_9571);
and U10309 (N_10309,N_9694,N_9555);
or U10310 (N_10310,N_9802,N_9584);
nor U10311 (N_10311,N_9753,N_9965);
and U10312 (N_10312,N_9533,N_9569);
and U10313 (N_10313,N_9721,N_9880);
nand U10314 (N_10314,N_9517,N_9753);
and U10315 (N_10315,N_9946,N_9540);
nor U10316 (N_10316,N_9567,N_9706);
and U10317 (N_10317,N_9758,N_9524);
nand U10318 (N_10318,N_9763,N_9987);
xor U10319 (N_10319,N_9811,N_9528);
nand U10320 (N_10320,N_9622,N_9710);
or U10321 (N_10321,N_9905,N_9867);
and U10322 (N_10322,N_9951,N_9915);
xor U10323 (N_10323,N_9779,N_9669);
and U10324 (N_10324,N_9974,N_9881);
nor U10325 (N_10325,N_9659,N_9790);
xor U10326 (N_10326,N_9531,N_9887);
or U10327 (N_10327,N_9571,N_9681);
or U10328 (N_10328,N_9922,N_9563);
and U10329 (N_10329,N_9870,N_9960);
nand U10330 (N_10330,N_9647,N_9707);
or U10331 (N_10331,N_9549,N_9817);
xor U10332 (N_10332,N_9800,N_9827);
or U10333 (N_10333,N_9534,N_9862);
and U10334 (N_10334,N_9558,N_9677);
nor U10335 (N_10335,N_9750,N_9617);
nand U10336 (N_10336,N_9977,N_9757);
and U10337 (N_10337,N_9744,N_9731);
and U10338 (N_10338,N_9909,N_9546);
nor U10339 (N_10339,N_9770,N_9832);
nand U10340 (N_10340,N_9905,N_9663);
xnor U10341 (N_10341,N_9584,N_9902);
or U10342 (N_10342,N_9674,N_9984);
or U10343 (N_10343,N_9788,N_9973);
nor U10344 (N_10344,N_9772,N_9921);
or U10345 (N_10345,N_9868,N_9845);
nand U10346 (N_10346,N_9987,N_9581);
xnor U10347 (N_10347,N_9974,N_9633);
nor U10348 (N_10348,N_9732,N_9516);
nand U10349 (N_10349,N_9702,N_9527);
and U10350 (N_10350,N_9813,N_9944);
or U10351 (N_10351,N_9611,N_9724);
xor U10352 (N_10352,N_9830,N_9804);
and U10353 (N_10353,N_9982,N_9581);
xnor U10354 (N_10354,N_9699,N_9738);
nor U10355 (N_10355,N_9822,N_9503);
xnor U10356 (N_10356,N_9503,N_9784);
nor U10357 (N_10357,N_9894,N_9923);
xnor U10358 (N_10358,N_9714,N_9718);
and U10359 (N_10359,N_9573,N_9983);
xnor U10360 (N_10360,N_9548,N_9754);
and U10361 (N_10361,N_9920,N_9658);
and U10362 (N_10362,N_9705,N_9762);
or U10363 (N_10363,N_9689,N_9837);
xnor U10364 (N_10364,N_9503,N_9840);
nor U10365 (N_10365,N_9576,N_9977);
or U10366 (N_10366,N_9847,N_9707);
and U10367 (N_10367,N_9725,N_9867);
and U10368 (N_10368,N_9625,N_9726);
and U10369 (N_10369,N_9899,N_9700);
xor U10370 (N_10370,N_9627,N_9585);
or U10371 (N_10371,N_9674,N_9933);
nor U10372 (N_10372,N_9967,N_9500);
nor U10373 (N_10373,N_9969,N_9526);
nand U10374 (N_10374,N_9952,N_9795);
or U10375 (N_10375,N_9861,N_9771);
xnor U10376 (N_10376,N_9927,N_9886);
xor U10377 (N_10377,N_9635,N_9917);
nand U10378 (N_10378,N_9616,N_9786);
nor U10379 (N_10379,N_9884,N_9927);
nand U10380 (N_10380,N_9899,N_9585);
xor U10381 (N_10381,N_9737,N_9644);
or U10382 (N_10382,N_9893,N_9890);
nand U10383 (N_10383,N_9848,N_9880);
xnor U10384 (N_10384,N_9877,N_9787);
xnor U10385 (N_10385,N_9557,N_9693);
and U10386 (N_10386,N_9916,N_9921);
and U10387 (N_10387,N_9629,N_9593);
nand U10388 (N_10388,N_9589,N_9636);
xor U10389 (N_10389,N_9792,N_9834);
and U10390 (N_10390,N_9889,N_9823);
nand U10391 (N_10391,N_9825,N_9834);
or U10392 (N_10392,N_9514,N_9613);
nand U10393 (N_10393,N_9590,N_9962);
or U10394 (N_10394,N_9540,N_9860);
and U10395 (N_10395,N_9641,N_9670);
and U10396 (N_10396,N_9573,N_9559);
and U10397 (N_10397,N_9852,N_9825);
or U10398 (N_10398,N_9724,N_9621);
nand U10399 (N_10399,N_9909,N_9870);
nor U10400 (N_10400,N_9650,N_9704);
xnor U10401 (N_10401,N_9967,N_9685);
nor U10402 (N_10402,N_9962,N_9837);
and U10403 (N_10403,N_9600,N_9816);
nor U10404 (N_10404,N_9811,N_9586);
nand U10405 (N_10405,N_9561,N_9963);
nand U10406 (N_10406,N_9997,N_9705);
xnor U10407 (N_10407,N_9574,N_9547);
or U10408 (N_10408,N_9536,N_9724);
nand U10409 (N_10409,N_9848,N_9996);
xnor U10410 (N_10410,N_9735,N_9517);
nor U10411 (N_10411,N_9844,N_9533);
nor U10412 (N_10412,N_9956,N_9948);
nand U10413 (N_10413,N_9545,N_9831);
or U10414 (N_10414,N_9896,N_9509);
or U10415 (N_10415,N_9606,N_9843);
xor U10416 (N_10416,N_9900,N_9945);
and U10417 (N_10417,N_9941,N_9935);
nand U10418 (N_10418,N_9520,N_9549);
nor U10419 (N_10419,N_9666,N_9898);
nand U10420 (N_10420,N_9511,N_9576);
or U10421 (N_10421,N_9634,N_9960);
nand U10422 (N_10422,N_9514,N_9820);
and U10423 (N_10423,N_9992,N_9925);
nor U10424 (N_10424,N_9648,N_9566);
nor U10425 (N_10425,N_9549,N_9593);
xnor U10426 (N_10426,N_9767,N_9827);
xnor U10427 (N_10427,N_9813,N_9677);
or U10428 (N_10428,N_9585,N_9826);
xor U10429 (N_10429,N_9600,N_9992);
nand U10430 (N_10430,N_9985,N_9748);
nand U10431 (N_10431,N_9592,N_9655);
and U10432 (N_10432,N_9573,N_9761);
nand U10433 (N_10433,N_9867,N_9509);
nor U10434 (N_10434,N_9500,N_9698);
nor U10435 (N_10435,N_9762,N_9538);
xor U10436 (N_10436,N_9560,N_9642);
xor U10437 (N_10437,N_9915,N_9901);
xor U10438 (N_10438,N_9598,N_9567);
nand U10439 (N_10439,N_9957,N_9677);
and U10440 (N_10440,N_9558,N_9963);
nand U10441 (N_10441,N_9778,N_9739);
or U10442 (N_10442,N_9768,N_9674);
nor U10443 (N_10443,N_9859,N_9505);
or U10444 (N_10444,N_9535,N_9510);
or U10445 (N_10445,N_9986,N_9996);
nand U10446 (N_10446,N_9668,N_9954);
and U10447 (N_10447,N_9713,N_9943);
nand U10448 (N_10448,N_9990,N_9595);
and U10449 (N_10449,N_9830,N_9652);
xnor U10450 (N_10450,N_9685,N_9536);
nor U10451 (N_10451,N_9763,N_9598);
or U10452 (N_10452,N_9886,N_9625);
xnor U10453 (N_10453,N_9937,N_9776);
nor U10454 (N_10454,N_9766,N_9680);
xnor U10455 (N_10455,N_9973,N_9956);
and U10456 (N_10456,N_9577,N_9521);
nor U10457 (N_10457,N_9894,N_9749);
xnor U10458 (N_10458,N_9666,N_9703);
xor U10459 (N_10459,N_9834,N_9703);
nor U10460 (N_10460,N_9778,N_9837);
xor U10461 (N_10461,N_9883,N_9833);
xnor U10462 (N_10462,N_9713,N_9822);
and U10463 (N_10463,N_9635,N_9925);
and U10464 (N_10464,N_9879,N_9709);
xor U10465 (N_10465,N_9716,N_9545);
nor U10466 (N_10466,N_9756,N_9650);
xnor U10467 (N_10467,N_9934,N_9702);
xor U10468 (N_10468,N_9655,N_9631);
nand U10469 (N_10469,N_9522,N_9841);
nand U10470 (N_10470,N_9866,N_9982);
and U10471 (N_10471,N_9834,N_9504);
or U10472 (N_10472,N_9707,N_9694);
and U10473 (N_10473,N_9660,N_9521);
and U10474 (N_10474,N_9991,N_9557);
or U10475 (N_10475,N_9833,N_9701);
or U10476 (N_10476,N_9937,N_9810);
nor U10477 (N_10477,N_9544,N_9841);
and U10478 (N_10478,N_9722,N_9641);
and U10479 (N_10479,N_9608,N_9724);
nor U10480 (N_10480,N_9598,N_9506);
or U10481 (N_10481,N_9929,N_9974);
or U10482 (N_10482,N_9511,N_9638);
nand U10483 (N_10483,N_9891,N_9608);
nor U10484 (N_10484,N_9504,N_9626);
or U10485 (N_10485,N_9542,N_9762);
xor U10486 (N_10486,N_9957,N_9813);
or U10487 (N_10487,N_9996,N_9906);
nand U10488 (N_10488,N_9863,N_9661);
and U10489 (N_10489,N_9759,N_9702);
or U10490 (N_10490,N_9541,N_9624);
nand U10491 (N_10491,N_9789,N_9935);
and U10492 (N_10492,N_9778,N_9501);
nor U10493 (N_10493,N_9878,N_9562);
or U10494 (N_10494,N_9740,N_9935);
and U10495 (N_10495,N_9771,N_9660);
and U10496 (N_10496,N_9934,N_9812);
and U10497 (N_10497,N_9887,N_9578);
nor U10498 (N_10498,N_9670,N_9505);
nor U10499 (N_10499,N_9975,N_9685);
and U10500 (N_10500,N_10456,N_10316);
nor U10501 (N_10501,N_10037,N_10004);
or U10502 (N_10502,N_10288,N_10060);
xor U10503 (N_10503,N_10098,N_10173);
nand U10504 (N_10504,N_10074,N_10244);
or U10505 (N_10505,N_10373,N_10106);
nor U10506 (N_10506,N_10372,N_10213);
xnor U10507 (N_10507,N_10387,N_10398);
or U10508 (N_10508,N_10204,N_10082);
nor U10509 (N_10509,N_10169,N_10237);
and U10510 (N_10510,N_10338,N_10374);
nand U10511 (N_10511,N_10426,N_10013);
xor U10512 (N_10512,N_10076,N_10136);
and U10513 (N_10513,N_10267,N_10181);
and U10514 (N_10514,N_10081,N_10469);
nand U10515 (N_10515,N_10070,N_10337);
or U10516 (N_10516,N_10485,N_10216);
and U10517 (N_10517,N_10444,N_10393);
and U10518 (N_10518,N_10443,N_10012);
or U10519 (N_10519,N_10091,N_10352);
or U10520 (N_10520,N_10332,N_10232);
xor U10521 (N_10521,N_10206,N_10363);
nor U10522 (N_10522,N_10360,N_10245);
nor U10523 (N_10523,N_10172,N_10318);
nand U10524 (N_10524,N_10005,N_10479);
or U10525 (N_10525,N_10410,N_10424);
nor U10526 (N_10526,N_10001,N_10336);
nor U10527 (N_10527,N_10429,N_10080);
nor U10528 (N_10528,N_10180,N_10068);
or U10529 (N_10529,N_10157,N_10043);
nand U10530 (N_10530,N_10063,N_10349);
xnor U10531 (N_10531,N_10484,N_10225);
nor U10532 (N_10532,N_10039,N_10481);
and U10533 (N_10533,N_10170,N_10141);
nor U10534 (N_10534,N_10190,N_10164);
nor U10535 (N_10535,N_10038,N_10112);
nand U10536 (N_10536,N_10249,N_10073);
nand U10537 (N_10537,N_10416,N_10467);
nor U10538 (N_10538,N_10470,N_10064);
or U10539 (N_10539,N_10368,N_10330);
nor U10540 (N_10540,N_10021,N_10389);
or U10541 (N_10541,N_10397,N_10411);
and U10542 (N_10542,N_10289,N_10111);
xor U10543 (N_10543,N_10491,N_10129);
nand U10544 (N_10544,N_10320,N_10108);
xnor U10545 (N_10545,N_10313,N_10487);
or U10546 (N_10546,N_10051,N_10420);
and U10547 (N_10547,N_10119,N_10104);
nand U10548 (N_10548,N_10034,N_10161);
nand U10549 (N_10549,N_10100,N_10083);
nand U10550 (N_10550,N_10270,N_10417);
nand U10551 (N_10551,N_10194,N_10322);
nand U10552 (N_10552,N_10125,N_10002);
and U10553 (N_10553,N_10048,N_10380);
nor U10554 (N_10554,N_10301,N_10113);
nand U10555 (N_10555,N_10009,N_10408);
nor U10556 (N_10556,N_10378,N_10055);
nor U10557 (N_10557,N_10238,N_10159);
xnor U10558 (N_10558,N_10310,N_10124);
nor U10559 (N_10559,N_10192,N_10453);
and U10560 (N_10560,N_10264,N_10077);
or U10561 (N_10561,N_10400,N_10427);
or U10562 (N_10562,N_10221,N_10341);
or U10563 (N_10563,N_10032,N_10230);
or U10564 (N_10564,N_10292,N_10193);
nor U10565 (N_10565,N_10153,N_10242);
nor U10566 (N_10566,N_10137,N_10053);
and U10567 (N_10567,N_10354,N_10144);
and U10568 (N_10568,N_10268,N_10234);
and U10569 (N_10569,N_10403,N_10086);
and U10570 (N_10570,N_10347,N_10448);
xor U10571 (N_10571,N_10201,N_10257);
or U10572 (N_10572,N_10383,N_10256);
xnor U10573 (N_10573,N_10088,N_10440);
xnor U10574 (N_10574,N_10454,N_10473);
nor U10575 (N_10575,N_10024,N_10371);
or U10576 (N_10576,N_10262,N_10482);
or U10577 (N_10577,N_10284,N_10406);
or U10578 (N_10578,N_10003,N_10016);
nor U10579 (N_10579,N_10187,N_10195);
nor U10580 (N_10580,N_10394,N_10110);
nand U10581 (N_10581,N_10303,N_10135);
and U10582 (N_10582,N_10029,N_10071);
or U10583 (N_10583,N_10353,N_10236);
and U10584 (N_10584,N_10033,N_10460);
nand U10585 (N_10585,N_10131,N_10140);
nand U10586 (N_10586,N_10247,N_10449);
or U10587 (N_10587,N_10049,N_10059);
nor U10588 (N_10588,N_10233,N_10185);
xnor U10589 (N_10589,N_10050,N_10497);
nand U10590 (N_10590,N_10329,N_10258);
and U10591 (N_10591,N_10286,N_10299);
and U10592 (N_10592,N_10189,N_10174);
nand U10593 (N_10593,N_10306,N_10413);
nor U10594 (N_10594,N_10327,N_10182);
nand U10595 (N_10595,N_10312,N_10437);
or U10596 (N_10596,N_10311,N_10228);
nor U10597 (N_10597,N_10023,N_10324);
and U10598 (N_10598,N_10415,N_10396);
xnor U10599 (N_10599,N_10027,N_10280);
or U10600 (N_10600,N_10197,N_10078);
nor U10601 (N_10601,N_10425,N_10483);
nand U10602 (N_10602,N_10490,N_10478);
and U10603 (N_10603,N_10328,N_10466);
or U10604 (N_10604,N_10399,N_10428);
xor U10605 (N_10605,N_10158,N_10227);
and U10606 (N_10606,N_10287,N_10447);
xnor U10607 (N_10607,N_10344,N_10395);
nand U10608 (N_10608,N_10465,N_10222);
and U10609 (N_10609,N_10127,N_10145);
and U10610 (N_10610,N_10441,N_10252);
xnor U10611 (N_10611,N_10155,N_10370);
or U10612 (N_10612,N_10178,N_10294);
xor U10613 (N_10613,N_10210,N_10331);
nor U10614 (N_10614,N_10496,N_10401);
or U10615 (N_10615,N_10134,N_10480);
and U10616 (N_10616,N_10279,N_10281);
xnor U10617 (N_10617,N_10323,N_10295);
or U10618 (N_10618,N_10462,N_10376);
nor U10619 (N_10619,N_10386,N_10022);
and U10620 (N_10620,N_10379,N_10253);
nand U10621 (N_10621,N_10163,N_10414);
xor U10622 (N_10622,N_10026,N_10066);
xor U10623 (N_10623,N_10435,N_10333);
nor U10624 (N_10624,N_10296,N_10203);
nand U10625 (N_10625,N_10058,N_10177);
nor U10626 (N_10626,N_10278,N_10260);
or U10627 (N_10627,N_10304,N_10167);
xor U10628 (N_10628,N_10459,N_10007);
nand U10629 (N_10629,N_10028,N_10404);
or U10630 (N_10630,N_10369,N_10486);
xnor U10631 (N_10631,N_10439,N_10087);
xor U10632 (N_10632,N_10208,N_10057);
xnor U10633 (N_10633,N_10432,N_10340);
and U10634 (N_10634,N_10402,N_10095);
and U10635 (N_10635,N_10277,N_10291);
nor U10636 (N_10636,N_10229,N_10302);
nor U10637 (N_10637,N_10079,N_10054);
and U10638 (N_10638,N_10419,N_10239);
xor U10639 (N_10639,N_10248,N_10308);
and U10640 (N_10640,N_10162,N_10412);
and U10641 (N_10641,N_10075,N_10243);
nand U10642 (N_10642,N_10364,N_10321);
or U10643 (N_10643,N_10207,N_10219);
xnor U10644 (N_10644,N_10315,N_10365);
xnor U10645 (N_10645,N_10384,N_10198);
and U10646 (N_10646,N_10138,N_10274);
nor U10647 (N_10647,N_10103,N_10405);
nand U10648 (N_10648,N_10122,N_10421);
or U10649 (N_10649,N_10133,N_10196);
and U10650 (N_10650,N_10130,N_10309);
xnor U10651 (N_10651,N_10094,N_10494);
or U10652 (N_10652,N_10014,N_10297);
and U10653 (N_10653,N_10492,N_10356);
and U10654 (N_10654,N_10090,N_10474);
nand U10655 (N_10655,N_10209,N_10409);
and U10656 (N_10656,N_10117,N_10151);
nand U10657 (N_10657,N_10290,N_10255);
nand U10658 (N_10658,N_10132,N_10160);
or U10659 (N_10659,N_10099,N_10214);
and U10660 (N_10660,N_10107,N_10121);
or U10661 (N_10661,N_10040,N_10362);
xnor U10662 (N_10662,N_10105,N_10150);
or U10663 (N_10663,N_10351,N_10346);
nand U10664 (N_10664,N_10250,N_10025);
or U10665 (N_10665,N_10283,N_10388);
nor U10666 (N_10666,N_10041,N_10461);
and U10667 (N_10667,N_10020,N_10114);
and U10668 (N_10668,N_10326,N_10065);
xor U10669 (N_10669,N_10045,N_10042);
and U10670 (N_10670,N_10457,N_10361);
and U10671 (N_10671,N_10477,N_10377);
nor U10672 (N_10672,N_10455,N_10407);
or U10673 (N_10673,N_10226,N_10089);
nand U10674 (N_10674,N_10282,N_10176);
or U10675 (N_10675,N_10061,N_10202);
or U10676 (N_10676,N_10231,N_10343);
xor U10677 (N_10677,N_10017,N_10438);
nor U10678 (N_10678,N_10285,N_10271);
nor U10679 (N_10679,N_10392,N_10251);
nand U10680 (N_10680,N_10350,N_10224);
nand U10681 (N_10681,N_10272,N_10056);
nand U10682 (N_10682,N_10254,N_10220);
or U10683 (N_10683,N_10463,N_10334);
and U10684 (N_10684,N_10434,N_10215);
nand U10685 (N_10685,N_10146,N_10442);
or U10686 (N_10686,N_10468,N_10367);
nor U10687 (N_10687,N_10339,N_10093);
and U10688 (N_10688,N_10265,N_10205);
nand U10689 (N_10689,N_10472,N_10390);
xnor U10690 (N_10690,N_10446,N_10010);
and U10691 (N_10691,N_10186,N_10019);
or U10692 (N_10692,N_10069,N_10342);
and U10693 (N_10693,N_10123,N_10325);
and U10694 (N_10694,N_10355,N_10188);
xnor U10695 (N_10695,N_10006,N_10148);
nand U10696 (N_10696,N_10235,N_10223);
and U10697 (N_10697,N_10348,N_10471);
nand U10698 (N_10698,N_10476,N_10200);
nand U10699 (N_10699,N_10120,N_10000);
xor U10700 (N_10700,N_10199,N_10431);
or U10701 (N_10701,N_10031,N_10097);
or U10702 (N_10702,N_10433,N_10092);
or U10703 (N_10703,N_10030,N_10418);
nand U10704 (N_10704,N_10035,N_10358);
nor U10705 (N_10705,N_10382,N_10317);
nor U10706 (N_10706,N_10183,N_10464);
or U10707 (N_10707,N_10430,N_10391);
and U10708 (N_10708,N_10475,N_10165);
nand U10709 (N_10709,N_10147,N_10015);
and U10710 (N_10710,N_10175,N_10126);
or U10711 (N_10711,N_10116,N_10168);
nor U10712 (N_10712,N_10044,N_10212);
or U10713 (N_10713,N_10067,N_10018);
nand U10714 (N_10714,N_10179,N_10085);
nand U10715 (N_10715,N_10381,N_10345);
xor U10716 (N_10716,N_10263,N_10241);
nand U10717 (N_10717,N_10084,N_10298);
nor U10718 (N_10718,N_10217,N_10240);
and U10719 (N_10719,N_10366,N_10008);
or U10720 (N_10720,N_10047,N_10266);
nand U10721 (N_10721,N_10359,N_10276);
and U10722 (N_10722,N_10458,N_10499);
xnor U10723 (N_10723,N_10246,N_10335);
or U10724 (N_10724,N_10218,N_10305);
and U10725 (N_10725,N_10314,N_10445);
xor U10726 (N_10726,N_10171,N_10422);
or U10727 (N_10727,N_10184,N_10357);
and U10728 (N_10728,N_10011,N_10436);
xor U10729 (N_10729,N_10300,N_10452);
and U10730 (N_10730,N_10096,N_10450);
xor U10731 (N_10731,N_10046,N_10101);
nand U10732 (N_10732,N_10062,N_10072);
nand U10733 (N_10733,N_10375,N_10102);
and U10734 (N_10734,N_10149,N_10261);
nand U10735 (N_10735,N_10166,N_10128);
nand U10736 (N_10736,N_10493,N_10152);
nor U10737 (N_10737,N_10109,N_10052);
xor U10738 (N_10738,N_10488,N_10259);
nor U10739 (N_10739,N_10385,N_10307);
or U10740 (N_10740,N_10319,N_10273);
or U10741 (N_10741,N_10156,N_10293);
nand U10742 (N_10742,N_10498,N_10154);
nor U10743 (N_10743,N_10211,N_10275);
nor U10744 (N_10744,N_10036,N_10143);
nor U10745 (N_10745,N_10142,N_10451);
and U10746 (N_10746,N_10495,N_10115);
and U10747 (N_10747,N_10118,N_10191);
nor U10748 (N_10748,N_10489,N_10139);
nor U10749 (N_10749,N_10269,N_10423);
or U10750 (N_10750,N_10154,N_10404);
xor U10751 (N_10751,N_10432,N_10118);
xor U10752 (N_10752,N_10262,N_10137);
and U10753 (N_10753,N_10485,N_10056);
xor U10754 (N_10754,N_10228,N_10326);
xor U10755 (N_10755,N_10057,N_10485);
nor U10756 (N_10756,N_10084,N_10246);
xnor U10757 (N_10757,N_10185,N_10482);
nor U10758 (N_10758,N_10074,N_10398);
and U10759 (N_10759,N_10025,N_10335);
nand U10760 (N_10760,N_10307,N_10333);
nand U10761 (N_10761,N_10022,N_10297);
or U10762 (N_10762,N_10331,N_10356);
nand U10763 (N_10763,N_10227,N_10283);
xor U10764 (N_10764,N_10103,N_10364);
and U10765 (N_10765,N_10194,N_10366);
or U10766 (N_10766,N_10314,N_10007);
nor U10767 (N_10767,N_10315,N_10276);
and U10768 (N_10768,N_10231,N_10342);
xnor U10769 (N_10769,N_10128,N_10459);
or U10770 (N_10770,N_10273,N_10381);
and U10771 (N_10771,N_10199,N_10223);
and U10772 (N_10772,N_10143,N_10149);
nand U10773 (N_10773,N_10420,N_10437);
nor U10774 (N_10774,N_10109,N_10134);
xnor U10775 (N_10775,N_10286,N_10012);
nor U10776 (N_10776,N_10184,N_10414);
xnor U10777 (N_10777,N_10349,N_10353);
nor U10778 (N_10778,N_10206,N_10372);
xnor U10779 (N_10779,N_10264,N_10148);
nand U10780 (N_10780,N_10340,N_10168);
nand U10781 (N_10781,N_10177,N_10357);
xor U10782 (N_10782,N_10098,N_10392);
nor U10783 (N_10783,N_10162,N_10133);
and U10784 (N_10784,N_10309,N_10377);
nand U10785 (N_10785,N_10137,N_10185);
and U10786 (N_10786,N_10094,N_10001);
nand U10787 (N_10787,N_10298,N_10455);
and U10788 (N_10788,N_10470,N_10368);
and U10789 (N_10789,N_10328,N_10496);
nor U10790 (N_10790,N_10053,N_10422);
and U10791 (N_10791,N_10025,N_10423);
or U10792 (N_10792,N_10372,N_10127);
nand U10793 (N_10793,N_10285,N_10305);
or U10794 (N_10794,N_10259,N_10373);
xor U10795 (N_10795,N_10299,N_10175);
xor U10796 (N_10796,N_10113,N_10326);
xor U10797 (N_10797,N_10143,N_10071);
xnor U10798 (N_10798,N_10084,N_10395);
or U10799 (N_10799,N_10424,N_10241);
nor U10800 (N_10800,N_10064,N_10424);
or U10801 (N_10801,N_10430,N_10400);
or U10802 (N_10802,N_10337,N_10263);
and U10803 (N_10803,N_10147,N_10220);
and U10804 (N_10804,N_10009,N_10167);
or U10805 (N_10805,N_10194,N_10185);
and U10806 (N_10806,N_10343,N_10207);
or U10807 (N_10807,N_10423,N_10429);
or U10808 (N_10808,N_10265,N_10441);
nor U10809 (N_10809,N_10438,N_10159);
and U10810 (N_10810,N_10287,N_10144);
nand U10811 (N_10811,N_10180,N_10341);
nor U10812 (N_10812,N_10153,N_10187);
and U10813 (N_10813,N_10078,N_10213);
xor U10814 (N_10814,N_10294,N_10414);
and U10815 (N_10815,N_10179,N_10299);
and U10816 (N_10816,N_10422,N_10444);
nand U10817 (N_10817,N_10208,N_10186);
xor U10818 (N_10818,N_10295,N_10202);
nand U10819 (N_10819,N_10303,N_10086);
nor U10820 (N_10820,N_10467,N_10465);
and U10821 (N_10821,N_10435,N_10203);
and U10822 (N_10822,N_10459,N_10410);
xor U10823 (N_10823,N_10294,N_10029);
xnor U10824 (N_10824,N_10080,N_10425);
xor U10825 (N_10825,N_10006,N_10223);
nor U10826 (N_10826,N_10234,N_10379);
or U10827 (N_10827,N_10328,N_10005);
xnor U10828 (N_10828,N_10328,N_10464);
nor U10829 (N_10829,N_10423,N_10375);
nand U10830 (N_10830,N_10240,N_10179);
xnor U10831 (N_10831,N_10435,N_10436);
nor U10832 (N_10832,N_10010,N_10157);
or U10833 (N_10833,N_10087,N_10035);
or U10834 (N_10834,N_10029,N_10210);
or U10835 (N_10835,N_10351,N_10222);
nor U10836 (N_10836,N_10408,N_10204);
xor U10837 (N_10837,N_10156,N_10233);
and U10838 (N_10838,N_10165,N_10234);
nand U10839 (N_10839,N_10409,N_10013);
xor U10840 (N_10840,N_10429,N_10350);
and U10841 (N_10841,N_10475,N_10484);
xnor U10842 (N_10842,N_10219,N_10318);
nand U10843 (N_10843,N_10341,N_10239);
nand U10844 (N_10844,N_10422,N_10448);
and U10845 (N_10845,N_10490,N_10059);
and U10846 (N_10846,N_10444,N_10401);
xor U10847 (N_10847,N_10046,N_10131);
nand U10848 (N_10848,N_10304,N_10279);
nor U10849 (N_10849,N_10469,N_10087);
or U10850 (N_10850,N_10032,N_10034);
or U10851 (N_10851,N_10467,N_10129);
and U10852 (N_10852,N_10438,N_10037);
nor U10853 (N_10853,N_10352,N_10176);
nand U10854 (N_10854,N_10233,N_10011);
xnor U10855 (N_10855,N_10376,N_10407);
and U10856 (N_10856,N_10235,N_10340);
xor U10857 (N_10857,N_10408,N_10316);
or U10858 (N_10858,N_10034,N_10465);
nand U10859 (N_10859,N_10131,N_10319);
or U10860 (N_10860,N_10015,N_10428);
nand U10861 (N_10861,N_10223,N_10491);
or U10862 (N_10862,N_10228,N_10399);
nor U10863 (N_10863,N_10393,N_10441);
and U10864 (N_10864,N_10330,N_10464);
xor U10865 (N_10865,N_10274,N_10170);
and U10866 (N_10866,N_10361,N_10292);
xor U10867 (N_10867,N_10239,N_10363);
nand U10868 (N_10868,N_10020,N_10415);
and U10869 (N_10869,N_10438,N_10155);
xor U10870 (N_10870,N_10312,N_10412);
nor U10871 (N_10871,N_10042,N_10077);
nand U10872 (N_10872,N_10311,N_10353);
xor U10873 (N_10873,N_10073,N_10463);
xnor U10874 (N_10874,N_10345,N_10327);
or U10875 (N_10875,N_10367,N_10194);
nand U10876 (N_10876,N_10105,N_10034);
nor U10877 (N_10877,N_10481,N_10199);
nor U10878 (N_10878,N_10458,N_10341);
nand U10879 (N_10879,N_10474,N_10000);
nor U10880 (N_10880,N_10007,N_10096);
xnor U10881 (N_10881,N_10106,N_10168);
nor U10882 (N_10882,N_10029,N_10282);
nor U10883 (N_10883,N_10342,N_10336);
and U10884 (N_10884,N_10181,N_10345);
nand U10885 (N_10885,N_10355,N_10455);
nand U10886 (N_10886,N_10388,N_10212);
or U10887 (N_10887,N_10362,N_10454);
xor U10888 (N_10888,N_10144,N_10101);
xor U10889 (N_10889,N_10183,N_10064);
nand U10890 (N_10890,N_10354,N_10010);
nor U10891 (N_10891,N_10450,N_10058);
nor U10892 (N_10892,N_10326,N_10210);
nand U10893 (N_10893,N_10190,N_10333);
and U10894 (N_10894,N_10408,N_10144);
and U10895 (N_10895,N_10407,N_10399);
and U10896 (N_10896,N_10137,N_10410);
nand U10897 (N_10897,N_10060,N_10179);
and U10898 (N_10898,N_10206,N_10480);
xor U10899 (N_10899,N_10378,N_10431);
xnor U10900 (N_10900,N_10347,N_10053);
and U10901 (N_10901,N_10497,N_10015);
nor U10902 (N_10902,N_10424,N_10147);
nor U10903 (N_10903,N_10152,N_10091);
or U10904 (N_10904,N_10026,N_10420);
nand U10905 (N_10905,N_10355,N_10024);
nor U10906 (N_10906,N_10308,N_10011);
xnor U10907 (N_10907,N_10252,N_10164);
or U10908 (N_10908,N_10432,N_10209);
or U10909 (N_10909,N_10081,N_10489);
nand U10910 (N_10910,N_10018,N_10063);
or U10911 (N_10911,N_10072,N_10071);
xnor U10912 (N_10912,N_10137,N_10349);
or U10913 (N_10913,N_10289,N_10003);
nor U10914 (N_10914,N_10173,N_10343);
and U10915 (N_10915,N_10256,N_10366);
nand U10916 (N_10916,N_10436,N_10272);
nor U10917 (N_10917,N_10275,N_10031);
nand U10918 (N_10918,N_10336,N_10386);
xnor U10919 (N_10919,N_10243,N_10091);
nand U10920 (N_10920,N_10123,N_10109);
nor U10921 (N_10921,N_10300,N_10015);
nor U10922 (N_10922,N_10360,N_10397);
xor U10923 (N_10923,N_10023,N_10394);
xor U10924 (N_10924,N_10465,N_10139);
xor U10925 (N_10925,N_10079,N_10334);
xor U10926 (N_10926,N_10016,N_10430);
nand U10927 (N_10927,N_10348,N_10312);
xnor U10928 (N_10928,N_10287,N_10097);
or U10929 (N_10929,N_10362,N_10155);
xnor U10930 (N_10930,N_10347,N_10418);
nand U10931 (N_10931,N_10093,N_10236);
nor U10932 (N_10932,N_10001,N_10180);
or U10933 (N_10933,N_10285,N_10241);
nor U10934 (N_10934,N_10107,N_10037);
xor U10935 (N_10935,N_10042,N_10112);
and U10936 (N_10936,N_10152,N_10344);
and U10937 (N_10937,N_10451,N_10219);
nand U10938 (N_10938,N_10201,N_10443);
or U10939 (N_10939,N_10372,N_10150);
or U10940 (N_10940,N_10098,N_10052);
xnor U10941 (N_10941,N_10472,N_10439);
nor U10942 (N_10942,N_10316,N_10380);
or U10943 (N_10943,N_10057,N_10185);
and U10944 (N_10944,N_10436,N_10015);
and U10945 (N_10945,N_10325,N_10032);
nand U10946 (N_10946,N_10309,N_10399);
nand U10947 (N_10947,N_10014,N_10388);
or U10948 (N_10948,N_10470,N_10138);
nand U10949 (N_10949,N_10080,N_10025);
nor U10950 (N_10950,N_10040,N_10343);
nor U10951 (N_10951,N_10486,N_10277);
xnor U10952 (N_10952,N_10430,N_10424);
or U10953 (N_10953,N_10488,N_10309);
nand U10954 (N_10954,N_10403,N_10031);
xnor U10955 (N_10955,N_10457,N_10070);
nand U10956 (N_10956,N_10237,N_10207);
nand U10957 (N_10957,N_10001,N_10327);
or U10958 (N_10958,N_10156,N_10459);
xnor U10959 (N_10959,N_10069,N_10002);
and U10960 (N_10960,N_10420,N_10135);
and U10961 (N_10961,N_10408,N_10018);
or U10962 (N_10962,N_10484,N_10173);
xor U10963 (N_10963,N_10469,N_10113);
nor U10964 (N_10964,N_10419,N_10171);
nand U10965 (N_10965,N_10023,N_10461);
xnor U10966 (N_10966,N_10280,N_10191);
nand U10967 (N_10967,N_10250,N_10461);
and U10968 (N_10968,N_10031,N_10178);
and U10969 (N_10969,N_10057,N_10064);
nand U10970 (N_10970,N_10004,N_10002);
or U10971 (N_10971,N_10163,N_10139);
and U10972 (N_10972,N_10030,N_10024);
nand U10973 (N_10973,N_10492,N_10393);
nand U10974 (N_10974,N_10156,N_10001);
or U10975 (N_10975,N_10354,N_10161);
nand U10976 (N_10976,N_10387,N_10324);
nor U10977 (N_10977,N_10403,N_10056);
and U10978 (N_10978,N_10364,N_10463);
and U10979 (N_10979,N_10475,N_10223);
or U10980 (N_10980,N_10217,N_10424);
and U10981 (N_10981,N_10196,N_10247);
or U10982 (N_10982,N_10136,N_10442);
or U10983 (N_10983,N_10051,N_10183);
nor U10984 (N_10984,N_10036,N_10115);
and U10985 (N_10985,N_10277,N_10274);
or U10986 (N_10986,N_10240,N_10087);
or U10987 (N_10987,N_10392,N_10266);
nand U10988 (N_10988,N_10131,N_10342);
xor U10989 (N_10989,N_10302,N_10355);
nand U10990 (N_10990,N_10148,N_10428);
xnor U10991 (N_10991,N_10139,N_10398);
xor U10992 (N_10992,N_10014,N_10003);
xnor U10993 (N_10993,N_10091,N_10024);
and U10994 (N_10994,N_10297,N_10403);
and U10995 (N_10995,N_10434,N_10048);
and U10996 (N_10996,N_10130,N_10484);
or U10997 (N_10997,N_10390,N_10153);
and U10998 (N_10998,N_10329,N_10304);
nand U10999 (N_10999,N_10430,N_10144);
xnor U11000 (N_11000,N_10555,N_10800);
xnor U11001 (N_11001,N_10567,N_10522);
xnor U11002 (N_11002,N_10955,N_10702);
nor U11003 (N_11003,N_10748,N_10991);
xnor U11004 (N_11004,N_10851,N_10858);
xnor U11005 (N_11005,N_10773,N_10712);
nand U11006 (N_11006,N_10525,N_10862);
or U11007 (N_11007,N_10917,N_10737);
or U11008 (N_11008,N_10837,N_10983);
xor U11009 (N_11009,N_10823,N_10880);
xnor U11010 (N_11010,N_10713,N_10740);
xnor U11011 (N_11011,N_10887,N_10946);
nor U11012 (N_11012,N_10523,N_10648);
nor U11013 (N_11013,N_10583,N_10581);
nand U11014 (N_11014,N_10844,N_10985);
nand U11015 (N_11015,N_10625,N_10565);
or U11016 (N_11016,N_10811,N_10757);
or U11017 (N_11017,N_10847,N_10626);
or U11018 (N_11018,N_10741,N_10743);
nor U11019 (N_11019,N_10520,N_10597);
xnor U11020 (N_11020,N_10898,N_10810);
and U11021 (N_11021,N_10832,N_10639);
or U11022 (N_11022,N_10872,N_10979);
and U11023 (N_11023,N_10723,N_10646);
nand U11024 (N_11024,N_10509,N_10751);
or U11025 (N_11025,N_10997,N_10641);
nor U11026 (N_11026,N_10848,N_10503);
and U11027 (N_11027,N_10782,N_10596);
nor U11028 (N_11028,N_10927,N_10553);
nor U11029 (N_11029,N_10933,N_10778);
and U11030 (N_11030,N_10765,N_10502);
nor U11031 (N_11031,N_10679,N_10547);
or U11032 (N_11032,N_10513,N_10952);
xor U11033 (N_11033,N_10856,N_10662);
and U11034 (N_11034,N_10876,N_10850);
nor U11035 (N_11035,N_10894,N_10651);
nor U11036 (N_11036,N_10841,N_10527);
nand U11037 (N_11037,N_10675,N_10661);
xor U11038 (N_11038,N_10653,N_10964);
and U11039 (N_11039,N_10584,N_10804);
xor U11040 (N_11040,N_10635,N_10775);
and U11041 (N_11041,N_10956,N_10730);
nor U11042 (N_11042,N_10993,N_10936);
xnor U11043 (N_11043,N_10899,N_10589);
xnor U11044 (N_11044,N_10693,N_10521);
xor U11045 (N_11045,N_10826,N_10557);
nand U11046 (N_11046,N_10754,N_10577);
and U11047 (N_11047,N_10629,N_10692);
xnor U11048 (N_11048,N_10652,N_10621);
nand U11049 (N_11049,N_10886,N_10822);
xor U11050 (N_11050,N_10888,N_10882);
xor U11051 (N_11051,N_10569,N_10682);
xor U11052 (N_11052,N_10963,N_10689);
or U11053 (N_11053,N_10901,N_10785);
and U11054 (N_11054,N_10877,N_10590);
nand U11055 (N_11055,N_10611,N_10815);
nand U11056 (N_11056,N_10637,N_10854);
nor U11057 (N_11057,N_10758,N_10632);
nor U11058 (N_11058,N_10756,N_10911);
or U11059 (N_11059,N_10966,N_10515);
nor U11060 (N_11060,N_10715,N_10514);
nand U11061 (N_11061,N_10643,N_10820);
nor U11062 (N_11062,N_10912,N_10697);
and U11063 (N_11063,N_10763,N_10551);
nor U11064 (N_11064,N_10501,N_10588);
and U11065 (N_11065,N_10871,N_10990);
nand U11066 (N_11066,N_10771,N_10510);
nand U11067 (N_11067,N_10972,N_10928);
or U11068 (N_11068,N_10708,N_10606);
nor U11069 (N_11069,N_10973,N_10591);
xor U11070 (N_11070,N_10792,N_10721);
xnor U11071 (N_11071,N_10812,N_10500);
xnor U11072 (N_11072,N_10825,N_10750);
or U11073 (N_11073,N_10705,N_10559);
or U11074 (N_11074,N_10633,N_10879);
or U11075 (N_11075,N_10587,N_10685);
nor U11076 (N_11076,N_10656,N_10563);
nor U11077 (N_11077,N_10746,N_10953);
xor U11078 (N_11078,N_10504,N_10951);
nand U11079 (N_11079,N_10529,N_10944);
nand U11080 (N_11080,N_10579,N_10842);
nor U11081 (N_11081,N_10707,N_10922);
nor U11082 (N_11082,N_10885,N_10824);
and U11083 (N_11083,N_10536,N_10895);
and U11084 (N_11084,N_10994,N_10564);
or U11085 (N_11085,N_10918,N_10650);
or U11086 (N_11086,N_10916,N_10586);
nand U11087 (N_11087,N_10897,N_10676);
and U11088 (N_11088,N_10505,N_10552);
nand U11089 (N_11089,N_10634,N_10699);
nor U11090 (N_11090,N_10869,N_10829);
nor U11091 (N_11091,N_10709,N_10821);
nand U11092 (N_11092,N_10600,N_10943);
and U11093 (N_11093,N_10747,N_10627);
or U11094 (N_11094,N_10870,N_10645);
xor U11095 (N_11095,N_10932,N_10580);
and U11096 (N_11096,N_10638,N_10941);
and U11097 (N_11097,N_10924,N_10961);
nor U11098 (N_11098,N_10843,N_10549);
and U11099 (N_11099,N_10772,N_10716);
and U11100 (N_11100,N_10992,N_10512);
or U11101 (N_11101,N_10873,N_10769);
and U11102 (N_11102,N_10957,N_10849);
nand U11103 (N_11103,N_10797,N_10686);
nand U11104 (N_11104,N_10840,N_10789);
nand U11105 (N_11105,N_10749,N_10831);
or U11106 (N_11106,N_10610,N_10779);
nor U11107 (N_11107,N_10808,N_10921);
nand U11108 (N_11108,N_10526,N_10636);
or U11109 (N_11109,N_10677,N_10718);
xor U11110 (N_11110,N_10574,N_10863);
nand U11111 (N_11111,N_10604,N_10742);
xnor U11112 (N_11112,N_10908,N_10934);
or U11113 (N_11113,N_10791,N_10962);
or U11114 (N_11114,N_10900,N_10836);
xnor U11115 (N_11115,N_10893,N_10706);
nand U11116 (N_11116,N_10524,N_10672);
nor U11117 (N_11117,N_10725,N_10560);
or U11118 (N_11118,N_10538,N_10942);
or U11119 (N_11119,N_10704,N_10561);
or U11120 (N_11120,N_10535,N_10919);
nor U11121 (N_11121,N_10981,N_10755);
nand U11122 (N_11122,N_10687,N_10976);
xor U11123 (N_11123,N_10915,N_10864);
and U11124 (N_11124,N_10805,N_10660);
or U11125 (N_11125,N_10620,N_10786);
and U11126 (N_11126,N_10603,N_10828);
and U11127 (N_11127,N_10582,N_10925);
nor U11128 (N_11128,N_10818,N_10999);
xor U11129 (N_11129,N_10809,N_10947);
nand U11130 (N_11130,N_10827,N_10539);
xor U11131 (N_11131,N_10914,N_10732);
and U11132 (N_11132,N_10562,N_10780);
nand U11133 (N_11133,N_10673,N_10619);
nand U11134 (N_11134,N_10930,N_10788);
or U11135 (N_11135,N_10507,N_10640);
nor U11136 (N_11136,N_10683,N_10913);
nand U11137 (N_11137,N_10982,N_10774);
or U11138 (N_11138,N_10855,N_10770);
and U11139 (N_11139,N_10960,N_10519);
or U11140 (N_11140,N_10950,N_10830);
or U11141 (N_11141,N_10680,N_10926);
or U11142 (N_11142,N_10859,N_10996);
or U11143 (N_11143,N_10534,N_10910);
nor U11144 (N_11144,N_10544,N_10806);
nand U11145 (N_11145,N_10546,N_10733);
nor U11146 (N_11146,N_10678,N_10846);
nand U11147 (N_11147,N_10543,N_10592);
or U11148 (N_11148,N_10695,N_10937);
and U11149 (N_11149,N_10753,N_10719);
nor U11150 (N_11150,N_10541,N_10696);
xor U11151 (N_11151,N_10784,N_10903);
and U11152 (N_11152,N_10764,N_10508);
or U11153 (N_11153,N_10967,N_10670);
xor U11154 (N_11154,N_10874,N_10613);
nand U11155 (N_11155,N_10988,N_10669);
and U11156 (N_11156,N_10608,N_10852);
nor U11157 (N_11157,N_10601,N_10690);
and U11158 (N_11158,N_10865,N_10684);
xor U11159 (N_11159,N_10572,N_10986);
nor U11160 (N_11160,N_10694,N_10896);
nor U11161 (N_11161,N_10954,N_10868);
or U11162 (N_11162,N_10935,N_10701);
xor U11163 (N_11163,N_10984,N_10623);
xnor U11164 (N_11164,N_10776,N_10722);
nor U11165 (N_11165,N_10731,N_10971);
nand U11166 (N_11166,N_10866,N_10803);
and U11167 (N_11167,N_10720,N_10599);
nand U11168 (N_11168,N_10940,N_10724);
nor U11169 (N_11169,N_10698,N_10816);
or U11170 (N_11170,N_10595,N_10931);
xnor U11171 (N_11171,N_10545,N_10867);
or U11172 (N_11172,N_10605,N_10542);
nor U11173 (N_11173,N_10736,N_10834);
nand U11174 (N_11174,N_10995,N_10594);
and U11175 (N_11175,N_10790,N_10745);
nand U11176 (N_11176,N_10884,N_10533);
or U11177 (N_11177,N_10568,N_10668);
xnor U11178 (N_11178,N_10795,N_10609);
xor U11179 (N_11179,N_10839,N_10977);
or U11180 (N_11180,N_10612,N_10875);
and U11181 (N_11181,N_10729,N_10614);
nor U11182 (N_11182,N_10615,N_10655);
and U11183 (N_11183,N_10618,N_10658);
xor U11184 (N_11184,N_10906,N_10923);
or U11185 (N_11185,N_10518,N_10783);
nand U11186 (N_11186,N_10891,N_10578);
nand U11187 (N_11187,N_10807,N_10970);
xnor U11188 (N_11188,N_10738,N_10835);
and U11189 (N_11189,N_10566,N_10674);
or U11190 (N_11190,N_10531,N_10762);
nand U11191 (N_11191,N_10728,N_10593);
nor U11192 (N_11192,N_10647,N_10796);
nand U11193 (N_11193,N_10691,N_10727);
and U11194 (N_11194,N_10550,N_10681);
or U11195 (N_11195,N_10516,N_10909);
and U11196 (N_11196,N_10793,N_10554);
xnor U11197 (N_11197,N_10573,N_10883);
and U11198 (N_11198,N_10703,N_10767);
nand U11199 (N_11199,N_10766,N_10665);
or U11200 (N_11200,N_10761,N_10642);
nand U11201 (N_11201,N_10714,N_10987);
and U11202 (N_11202,N_10735,N_10624);
xor U11203 (N_11203,N_10860,N_10532);
nand U11204 (N_11204,N_10777,N_10734);
nand U11205 (N_11205,N_10890,N_10958);
nand U11206 (N_11206,N_10833,N_10666);
nand U11207 (N_11207,N_10853,N_10585);
and U11208 (N_11208,N_10861,N_10945);
and U11209 (N_11209,N_10659,N_10688);
nand U11210 (N_11210,N_10664,N_10929);
nand U11211 (N_11211,N_10571,N_10628);
and U11212 (N_11212,N_10630,N_10904);
and U11213 (N_11213,N_10878,N_10781);
nor U11214 (N_11214,N_10576,N_10540);
and U11215 (N_11215,N_10857,N_10817);
xor U11216 (N_11216,N_10980,N_10889);
xnor U11217 (N_11217,N_10607,N_10975);
xor U11218 (N_11218,N_10710,N_10949);
nor U11219 (N_11219,N_10819,N_10989);
or U11220 (N_11220,N_10948,N_10787);
and U11221 (N_11221,N_10938,N_10517);
xor U11222 (N_11222,N_10907,N_10902);
xnor U11223 (N_11223,N_10798,N_10617);
nor U11224 (N_11224,N_10759,N_10570);
and U11225 (N_11225,N_10801,N_10700);
nand U11226 (N_11226,N_10506,N_10556);
xnor U11227 (N_11227,N_10598,N_10622);
and U11228 (N_11228,N_10978,N_10813);
and U11229 (N_11229,N_10537,N_10511);
nor U11230 (N_11230,N_10905,N_10845);
nand U11231 (N_11231,N_10711,N_10744);
and U11232 (N_11232,N_10760,N_10794);
xor U11233 (N_11233,N_10965,N_10838);
and U11234 (N_11234,N_10802,N_10998);
nor U11235 (N_11235,N_10663,N_10726);
xnor U11236 (N_11236,N_10969,N_10644);
and U11237 (N_11237,N_10920,N_10974);
nand U11238 (N_11238,N_10654,N_10739);
nor U11239 (N_11239,N_10616,N_10548);
xor U11240 (N_11240,N_10717,N_10649);
nand U11241 (N_11241,N_10602,N_10530);
xor U11242 (N_11242,N_10881,N_10575);
and U11243 (N_11243,N_10667,N_10671);
or U11244 (N_11244,N_10558,N_10799);
and U11245 (N_11245,N_10657,N_10892);
nor U11246 (N_11246,N_10528,N_10752);
nor U11247 (N_11247,N_10814,N_10968);
xnor U11248 (N_11248,N_10939,N_10959);
and U11249 (N_11249,N_10768,N_10631);
xor U11250 (N_11250,N_10733,N_10871);
nor U11251 (N_11251,N_10805,N_10995);
nor U11252 (N_11252,N_10513,N_10707);
xnor U11253 (N_11253,N_10909,N_10914);
nor U11254 (N_11254,N_10793,N_10786);
or U11255 (N_11255,N_10587,N_10747);
or U11256 (N_11256,N_10942,N_10643);
and U11257 (N_11257,N_10650,N_10952);
and U11258 (N_11258,N_10726,N_10948);
nand U11259 (N_11259,N_10781,N_10862);
or U11260 (N_11260,N_10656,N_10673);
and U11261 (N_11261,N_10772,N_10912);
xnor U11262 (N_11262,N_10885,N_10556);
nand U11263 (N_11263,N_10953,N_10815);
nor U11264 (N_11264,N_10928,N_10799);
nand U11265 (N_11265,N_10535,N_10840);
nor U11266 (N_11266,N_10501,N_10614);
or U11267 (N_11267,N_10931,N_10808);
or U11268 (N_11268,N_10798,N_10576);
and U11269 (N_11269,N_10970,N_10561);
nor U11270 (N_11270,N_10627,N_10615);
nor U11271 (N_11271,N_10503,N_10587);
and U11272 (N_11272,N_10559,N_10555);
nand U11273 (N_11273,N_10802,N_10642);
or U11274 (N_11274,N_10740,N_10915);
nand U11275 (N_11275,N_10807,N_10631);
or U11276 (N_11276,N_10851,N_10962);
nand U11277 (N_11277,N_10605,N_10560);
nand U11278 (N_11278,N_10907,N_10678);
or U11279 (N_11279,N_10727,N_10581);
xnor U11280 (N_11280,N_10894,N_10988);
nand U11281 (N_11281,N_10713,N_10642);
or U11282 (N_11282,N_10544,N_10734);
and U11283 (N_11283,N_10830,N_10560);
nor U11284 (N_11284,N_10883,N_10582);
and U11285 (N_11285,N_10593,N_10636);
xor U11286 (N_11286,N_10627,N_10994);
and U11287 (N_11287,N_10533,N_10789);
and U11288 (N_11288,N_10803,N_10794);
nand U11289 (N_11289,N_10631,N_10667);
and U11290 (N_11290,N_10509,N_10583);
or U11291 (N_11291,N_10819,N_10788);
nor U11292 (N_11292,N_10559,N_10507);
nand U11293 (N_11293,N_10770,N_10512);
or U11294 (N_11294,N_10552,N_10653);
nor U11295 (N_11295,N_10869,N_10915);
nor U11296 (N_11296,N_10518,N_10583);
xnor U11297 (N_11297,N_10979,N_10964);
xnor U11298 (N_11298,N_10744,N_10795);
nor U11299 (N_11299,N_10568,N_10873);
xor U11300 (N_11300,N_10712,N_10983);
xor U11301 (N_11301,N_10794,N_10570);
and U11302 (N_11302,N_10956,N_10766);
or U11303 (N_11303,N_10568,N_10800);
nor U11304 (N_11304,N_10842,N_10692);
or U11305 (N_11305,N_10666,N_10957);
and U11306 (N_11306,N_10587,N_10649);
nor U11307 (N_11307,N_10710,N_10952);
xor U11308 (N_11308,N_10905,N_10537);
nor U11309 (N_11309,N_10703,N_10686);
nand U11310 (N_11310,N_10592,N_10852);
nor U11311 (N_11311,N_10874,N_10789);
and U11312 (N_11312,N_10928,N_10966);
nor U11313 (N_11313,N_10889,N_10930);
and U11314 (N_11314,N_10648,N_10753);
nor U11315 (N_11315,N_10598,N_10674);
nand U11316 (N_11316,N_10721,N_10744);
nor U11317 (N_11317,N_10544,N_10507);
nor U11318 (N_11318,N_10757,N_10778);
and U11319 (N_11319,N_10970,N_10990);
and U11320 (N_11320,N_10558,N_10873);
and U11321 (N_11321,N_10922,N_10831);
nor U11322 (N_11322,N_10614,N_10677);
and U11323 (N_11323,N_10730,N_10780);
and U11324 (N_11324,N_10886,N_10924);
and U11325 (N_11325,N_10750,N_10934);
nand U11326 (N_11326,N_10919,N_10510);
or U11327 (N_11327,N_10774,N_10574);
nand U11328 (N_11328,N_10611,N_10850);
xnor U11329 (N_11329,N_10615,N_10819);
xnor U11330 (N_11330,N_10934,N_10674);
nor U11331 (N_11331,N_10812,N_10732);
nand U11332 (N_11332,N_10922,N_10892);
or U11333 (N_11333,N_10836,N_10603);
nor U11334 (N_11334,N_10973,N_10582);
nor U11335 (N_11335,N_10845,N_10898);
xnor U11336 (N_11336,N_10910,N_10649);
nand U11337 (N_11337,N_10991,N_10706);
nand U11338 (N_11338,N_10698,N_10841);
xor U11339 (N_11339,N_10687,N_10873);
nand U11340 (N_11340,N_10820,N_10654);
or U11341 (N_11341,N_10764,N_10528);
and U11342 (N_11342,N_10798,N_10589);
xor U11343 (N_11343,N_10592,N_10563);
xor U11344 (N_11344,N_10520,N_10851);
xor U11345 (N_11345,N_10807,N_10587);
and U11346 (N_11346,N_10517,N_10826);
xnor U11347 (N_11347,N_10841,N_10779);
nor U11348 (N_11348,N_10990,N_10580);
nor U11349 (N_11349,N_10515,N_10538);
nand U11350 (N_11350,N_10982,N_10925);
nor U11351 (N_11351,N_10898,N_10660);
and U11352 (N_11352,N_10767,N_10764);
nor U11353 (N_11353,N_10857,N_10697);
nand U11354 (N_11354,N_10796,N_10518);
and U11355 (N_11355,N_10922,N_10642);
nand U11356 (N_11356,N_10968,N_10844);
or U11357 (N_11357,N_10709,N_10637);
nand U11358 (N_11358,N_10671,N_10795);
and U11359 (N_11359,N_10692,N_10662);
and U11360 (N_11360,N_10853,N_10726);
or U11361 (N_11361,N_10750,N_10561);
nor U11362 (N_11362,N_10817,N_10618);
or U11363 (N_11363,N_10916,N_10753);
xor U11364 (N_11364,N_10571,N_10551);
nor U11365 (N_11365,N_10715,N_10544);
nor U11366 (N_11366,N_10725,N_10958);
nand U11367 (N_11367,N_10727,N_10531);
nand U11368 (N_11368,N_10841,N_10828);
and U11369 (N_11369,N_10814,N_10650);
xor U11370 (N_11370,N_10673,N_10843);
nor U11371 (N_11371,N_10720,N_10690);
nor U11372 (N_11372,N_10560,N_10527);
and U11373 (N_11373,N_10754,N_10654);
nor U11374 (N_11374,N_10791,N_10922);
nor U11375 (N_11375,N_10882,N_10645);
xor U11376 (N_11376,N_10635,N_10861);
nor U11377 (N_11377,N_10511,N_10871);
nand U11378 (N_11378,N_10733,N_10567);
xor U11379 (N_11379,N_10586,N_10528);
or U11380 (N_11380,N_10756,N_10544);
nand U11381 (N_11381,N_10678,N_10687);
nand U11382 (N_11382,N_10771,N_10584);
xor U11383 (N_11383,N_10867,N_10653);
or U11384 (N_11384,N_10513,N_10873);
and U11385 (N_11385,N_10854,N_10711);
xor U11386 (N_11386,N_10817,N_10521);
and U11387 (N_11387,N_10959,N_10812);
or U11388 (N_11388,N_10585,N_10947);
nor U11389 (N_11389,N_10511,N_10502);
or U11390 (N_11390,N_10571,N_10699);
nand U11391 (N_11391,N_10843,N_10539);
and U11392 (N_11392,N_10829,N_10585);
nor U11393 (N_11393,N_10667,N_10733);
nor U11394 (N_11394,N_10601,N_10780);
and U11395 (N_11395,N_10700,N_10722);
or U11396 (N_11396,N_10890,N_10986);
and U11397 (N_11397,N_10881,N_10860);
nor U11398 (N_11398,N_10640,N_10548);
nor U11399 (N_11399,N_10770,N_10919);
nor U11400 (N_11400,N_10961,N_10596);
nand U11401 (N_11401,N_10828,N_10821);
nor U11402 (N_11402,N_10733,N_10961);
or U11403 (N_11403,N_10944,N_10982);
nand U11404 (N_11404,N_10505,N_10524);
and U11405 (N_11405,N_10518,N_10825);
and U11406 (N_11406,N_10892,N_10783);
or U11407 (N_11407,N_10842,N_10650);
xnor U11408 (N_11408,N_10522,N_10716);
nand U11409 (N_11409,N_10732,N_10535);
nand U11410 (N_11410,N_10825,N_10953);
nand U11411 (N_11411,N_10993,N_10512);
nor U11412 (N_11412,N_10707,N_10644);
or U11413 (N_11413,N_10829,N_10996);
and U11414 (N_11414,N_10982,N_10743);
xnor U11415 (N_11415,N_10795,N_10696);
xnor U11416 (N_11416,N_10993,N_10519);
nor U11417 (N_11417,N_10904,N_10621);
nor U11418 (N_11418,N_10668,N_10708);
or U11419 (N_11419,N_10794,N_10737);
nor U11420 (N_11420,N_10567,N_10601);
nand U11421 (N_11421,N_10665,N_10743);
and U11422 (N_11422,N_10574,N_10795);
nand U11423 (N_11423,N_10615,N_10618);
nand U11424 (N_11424,N_10858,N_10797);
nand U11425 (N_11425,N_10783,N_10878);
and U11426 (N_11426,N_10862,N_10570);
xor U11427 (N_11427,N_10766,N_10781);
nor U11428 (N_11428,N_10790,N_10776);
nor U11429 (N_11429,N_10906,N_10614);
xor U11430 (N_11430,N_10998,N_10943);
nand U11431 (N_11431,N_10544,N_10980);
xor U11432 (N_11432,N_10728,N_10665);
and U11433 (N_11433,N_10992,N_10575);
nor U11434 (N_11434,N_10903,N_10991);
and U11435 (N_11435,N_10534,N_10933);
and U11436 (N_11436,N_10681,N_10899);
nand U11437 (N_11437,N_10614,N_10556);
nand U11438 (N_11438,N_10887,N_10706);
nand U11439 (N_11439,N_10746,N_10600);
nor U11440 (N_11440,N_10706,N_10995);
nor U11441 (N_11441,N_10556,N_10698);
xnor U11442 (N_11442,N_10593,N_10837);
nor U11443 (N_11443,N_10966,N_10755);
or U11444 (N_11444,N_10527,N_10839);
or U11445 (N_11445,N_10839,N_10622);
or U11446 (N_11446,N_10785,N_10531);
or U11447 (N_11447,N_10565,N_10721);
or U11448 (N_11448,N_10935,N_10785);
and U11449 (N_11449,N_10716,N_10864);
xnor U11450 (N_11450,N_10873,N_10986);
or U11451 (N_11451,N_10717,N_10612);
nand U11452 (N_11452,N_10698,N_10516);
nand U11453 (N_11453,N_10751,N_10970);
nor U11454 (N_11454,N_10947,N_10751);
or U11455 (N_11455,N_10784,N_10726);
nor U11456 (N_11456,N_10842,N_10720);
xnor U11457 (N_11457,N_10949,N_10966);
or U11458 (N_11458,N_10897,N_10627);
nor U11459 (N_11459,N_10657,N_10645);
nor U11460 (N_11460,N_10927,N_10843);
nor U11461 (N_11461,N_10522,N_10707);
and U11462 (N_11462,N_10536,N_10503);
nand U11463 (N_11463,N_10824,N_10986);
and U11464 (N_11464,N_10519,N_10922);
and U11465 (N_11465,N_10820,N_10639);
or U11466 (N_11466,N_10948,N_10778);
and U11467 (N_11467,N_10555,N_10503);
nor U11468 (N_11468,N_10859,N_10710);
or U11469 (N_11469,N_10969,N_10567);
nor U11470 (N_11470,N_10841,N_10717);
nand U11471 (N_11471,N_10839,N_10521);
nor U11472 (N_11472,N_10998,N_10579);
xnor U11473 (N_11473,N_10554,N_10691);
xnor U11474 (N_11474,N_10592,N_10715);
nand U11475 (N_11475,N_10960,N_10563);
nor U11476 (N_11476,N_10679,N_10674);
or U11477 (N_11477,N_10847,N_10592);
and U11478 (N_11478,N_10544,N_10699);
or U11479 (N_11479,N_10851,N_10860);
or U11480 (N_11480,N_10827,N_10623);
or U11481 (N_11481,N_10581,N_10730);
nor U11482 (N_11482,N_10567,N_10550);
nor U11483 (N_11483,N_10747,N_10599);
and U11484 (N_11484,N_10979,N_10789);
and U11485 (N_11485,N_10916,N_10585);
xnor U11486 (N_11486,N_10953,N_10566);
xor U11487 (N_11487,N_10930,N_10544);
and U11488 (N_11488,N_10758,N_10997);
xor U11489 (N_11489,N_10682,N_10875);
and U11490 (N_11490,N_10847,N_10785);
nor U11491 (N_11491,N_10758,N_10926);
xor U11492 (N_11492,N_10712,N_10768);
nand U11493 (N_11493,N_10868,N_10904);
nand U11494 (N_11494,N_10531,N_10713);
nand U11495 (N_11495,N_10918,N_10854);
nor U11496 (N_11496,N_10681,N_10679);
and U11497 (N_11497,N_10843,N_10782);
or U11498 (N_11498,N_10666,N_10722);
or U11499 (N_11499,N_10993,N_10576);
xor U11500 (N_11500,N_11157,N_11491);
or U11501 (N_11501,N_11356,N_11118);
nor U11502 (N_11502,N_11100,N_11163);
xnor U11503 (N_11503,N_11489,N_11360);
and U11504 (N_11504,N_11062,N_11239);
and U11505 (N_11505,N_11327,N_11098);
nor U11506 (N_11506,N_11396,N_11310);
nor U11507 (N_11507,N_11135,N_11374);
nand U11508 (N_11508,N_11150,N_11268);
nor U11509 (N_11509,N_11347,N_11463);
or U11510 (N_11510,N_11137,N_11017);
or U11511 (N_11511,N_11292,N_11229);
and U11512 (N_11512,N_11402,N_11476);
nor U11513 (N_11513,N_11086,N_11115);
or U11514 (N_11514,N_11355,N_11466);
and U11515 (N_11515,N_11465,N_11040);
or U11516 (N_11516,N_11461,N_11253);
and U11517 (N_11517,N_11131,N_11187);
nand U11518 (N_11518,N_11404,N_11249);
and U11519 (N_11519,N_11052,N_11318);
xor U11520 (N_11520,N_11497,N_11336);
or U11521 (N_11521,N_11431,N_11054);
and U11522 (N_11522,N_11194,N_11147);
and U11523 (N_11523,N_11428,N_11076);
or U11524 (N_11524,N_11285,N_11316);
nand U11525 (N_11525,N_11289,N_11270);
nor U11526 (N_11526,N_11486,N_11204);
xor U11527 (N_11527,N_11481,N_11004);
nand U11528 (N_11528,N_11357,N_11275);
xor U11529 (N_11529,N_11032,N_11277);
nand U11530 (N_11530,N_11291,N_11274);
xor U11531 (N_11531,N_11425,N_11203);
nor U11532 (N_11532,N_11283,N_11315);
xor U11533 (N_11533,N_11273,N_11156);
xnor U11534 (N_11534,N_11044,N_11440);
and U11535 (N_11535,N_11041,N_11256);
nand U11536 (N_11536,N_11499,N_11300);
and U11537 (N_11537,N_11021,N_11317);
or U11538 (N_11538,N_11457,N_11104);
or U11539 (N_11539,N_11170,N_11089);
or U11540 (N_11540,N_11234,N_11320);
xnor U11541 (N_11541,N_11332,N_11001);
or U11542 (N_11542,N_11127,N_11394);
xnor U11543 (N_11543,N_11324,N_11141);
or U11544 (N_11544,N_11297,N_11210);
nor U11545 (N_11545,N_11395,N_11353);
and U11546 (N_11546,N_11050,N_11047);
or U11547 (N_11547,N_11397,N_11306);
nor U11548 (N_11548,N_11252,N_11091);
or U11549 (N_11549,N_11458,N_11368);
xnor U11550 (N_11550,N_11443,N_11454);
xnor U11551 (N_11551,N_11337,N_11217);
xnor U11552 (N_11552,N_11364,N_11418);
and U11553 (N_11553,N_11212,N_11031);
nor U11554 (N_11554,N_11186,N_11305);
nor U11555 (N_11555,N_11095,N_11201);
xnor U11556 (N_11556,N_11023,N_11140);
and U11557 (N_11557,N_11061,N_11278);
nor U11558 (N_11558,N_11208,N_11171);
nand U11559 (N_11559,N_11109,N_11205);
nand U11560 (N_11560,N_11412,N_11175);
and U11561 (N_11561,N_11480,N_11120);
and U11562 (N_11562,N_11084,N_11366);
nor U11563 (N_11563,N_11319,N_11279);
nor U11564 (N_11564,N_11479,N_11482);
xnor U11565 (N_11565,N_11471,N_11290);
and U11566 (N_11566,N_11011,N_11019);
and U11567 (N_11567,N_11375,N_11301);
nor U11568 (N_11568,N_11348,N_11258);
or U11569 (N_11569,N_11447,N_11034);
nor U11570 (N_11570,N_11035,N_11003);
and U11571 (N_11571,N_11060,N_11436);
xnor U11572 (N_11572,N_11340,N_11166);
or U11573 (N_11573,N_11262,N_11071);
nor U11574 (N_11574,N_11048,N_11000);
nand U11575 (N_11575,N_11237,N_11331);
and U11576 (N_11576,N_11072,N_11329);
and U11577 (N_11577,N_11370,N_11460);
or U11578 (N_11578,N_11488,N_11129);
nand U11579 (N_11579,N_11422,N_11354);
nand U11580 (N_11580,N_11092,N_11213);
and U11581 (N_11581,N_11117,N_11420);
and U11582 (N_11582,N_11106,N_11393);
or U11583 (N_11583,N_11039,N_11198);
xor U11584 (N_11584,N_11132,N_11246);
nor U11585 (N_11585,N_11287,N_11361);
nand U11586 (N_11586,N_11018,N_11407);
xnor U11587 (N_11587,N_11371,N_11267);
and U11588 (N_11588,N_11437,N_11493);
xor U11589 (N_11589,N_11349,N_11495);
nor U11590 (N_11590,N_11028,N_11083);
or U11591 (N_11591,N_11142,N_11452);
xor U11592 (N_11592,N_11439,N_11259);
and U11593 (N_11593,N_11008,N_11073);
nand U11594 (N_11594,N_11230,N_11335);
or U11595 (N_11595,N_11146,N_11302);
and U11596 (N_11596,N_11191,N_11243);
nand U11597 (N_11597,N_11236,N_11222);
or U11598 (N_11598,N_11006,N_11051);
or U11599 (N_11599,N_11167,N_11231);
nand U11600 (N_11600,N_11449,N_11174);
or U11601 (N_11601,N_11079,N_11383);
or U11602 (N_11602,N_11328,N_11260);
xnor U11603 (N_11603,N_11215,N_11244);
nand U11604 (N_11604,N_11211,N_11413);
or U11605 (N_11605,N_11139,N_11264);
xnor U11606 (N_11606,N_11430,N_11379);
and U11607 (N_11607,N_11369,N_11433);
xnor U11608 (N_11608,N_11330,N_11446);
or U11609 (N_11609,N_11272,N_11414);
nand U11610 (N_11610,N_11380,N_11358);
and U11611 (N_11611,N_11046,N_11112);
and U11612 (N_11612,N_11322,N_11299);
nand U11613 (N_11613,N_11392,N_11250);
and U11614 (N_11614,N_11389,N_11126);
nor U11615 (N_11615,N_11136,N_11055);
nand U11616 (N_11616,N_11138,N_11159);
nor U11617 (N_11617,N_11056,N_11029);
or U11618 (N_11618,N_11228,N_11030);
nor U11619 (N_11619,N_11043,N_11288);
nor U11620 (N_11620,N_11189,N_11474);
or U11621 (N_11621,N_11386,N_11013);
nand U11622 (N_11622,N_11464,N_11063);
and U11623 (N_11623,N_11101,N_11227);
xor U11624 (N_11624,N_11042,N_11445);
nand U11625 (N_11625,N_11200,N_11107);
nor U11626 (N_11626,N_11294,N_11225);
nand U11627 (N_11627,N_11341,N_11359);
and U11628 (N_11628,N_11188,N_11235);
nor U11629 (N_11629,N_11027,N_11350);
nor U11630 (N_11630,N_11220,N_11085);
nor U11631 (N_11631,N_11475,N_11192);
or U11632 (N_11632,N_11382,N_11207);
xnor U11633 (N_11633,N_11090,N_11453);
and U11634 (N_11634,N_11065,N_11321);
and U11635 (N_11635,N_11459,N_11469);
nand U11636 (N_11636,N_11399,N_11058);
and U11637 (N_11637,N_11053,N_11206);
nor U11638 (N_11638,N_11345,N_11049);
nand U11639 (N_11639,N_11180,N_11160);
xnor U11640 (N_11640,N_11088,N_11143);
and U11641 (N_11641,N_11417,N_11097);
xor U11642 (N_11642,N_11276,N_11036);
nand U11643 (N_11643,N_11007,N_11074);
nor U11644 (N_11644,N_11066,N_11421);
xor U11645 (N_11645,N_11400,N_11339);
nand U11646 (N_11646,N_11247,N_11080);
or U11647 (N_11647,N_11401,N_11390);
nor U11648 (N_11648,N_11432,N_11026);
or U11649 (N_11649,N_11245,N_11221);
xor U11650 (N_11650,N_11408,N_11196);
or U11651 (N_11651,N_11271,N_11110);
nand U11652 (N_11652,N_11162,N_11450);
nand U11653 (N_11653,N_11151,N_11185);
or U11654 (N_11654,N_11014,N_11391);
nand U11655 (N_11655,N_11442,N_11233);
and U11656 (N_11656,N_11202,N_11059);
nor U11657 (N_11657,N_11311,N_11184);
nand U11658 (N_11658,N_11093,N_11016);
or U11659 (N_11659,N_11165,N_11387);
nand U11660 (N_11660,N_11284,N_11251);
xor U11661 (N_11661,N_11381,N_11045);
or U11662 (N_11662,N_11438,N_11248);
xor U11663 (N_11663,N_11190,N_11304);
nand U11664 (N_11664,N_11009,N_11424);
nand U11665 (N_11665,N_11241,N_11492);
xor U11666 (N_11666,N_11351,N_11012);
nand U11667 (N_11667,N_11022,N_11265);
nor U11668 (N_11668,N_11099,N_11002);
or U11669 (N_11669,N_11119,N_11467);
or U11670 (N_11670,N_11209,N_11455);
and U11671 (N_11671,N_11176,N_11333);
nor U11672 (N_11672,N_11087,N_11462);
nor U11673 (N_11673,N_11238,N_11114);
nand U11674 (N_11674,N_11193,N_11344);
xor U11675 (N_11675,N_11307,N_11406);
nor U11676 (N_11676,N_11161,N_11484);
xnor U11677 (N_11677,N_11216,N_11472);
or U11678 (N_11678,N_11286,N_11255);
or U11679 (N_11679,N_11309,N_11451);
xnor U11680 (N_11680,N_11338,N_11130);
nor U11681 (N_11681,N_11257,N_11195);
xnor U11682 (N_11682,N_11173,N_11411);
nor U11683 (N_11683,N_11434,N_11064);
and U11684 (N_11684,N_11281,N_11182);
xor U11685 (N_11685,N_11070,N_11082);
or U11686 (N_11686,N_11125,N_11025);
or U11687 (N_11687,N_11128,N_11367);
or U11688 (N_11688,N_11263,N_11199);
nor U11689 (N_11689,N_11197,N_11282);
and U11690 (N_11690,N_11183,N_11308);
and U11691 (N_11691,N_11024,N_11232);
xnor U11692 (N_11692,N_11154,N_11403);
or U11693 (N_11693,N_11015,N_11298);
and U11694 (N_11694,N_11470,N_11121);
nor U11695 (N_11695,N_11113,N_11485);
and U11696 (N_11696,N_11385,N_11346);
or U11697 (N_11697,N_11473,N_11269);
xor U11698 (N_11698,N_11133,N_11240);
or U11699 (N_11699,N_11498,N_11342);
nand U11700 (N_11700,N_11168,N_11122);
xnor U11701 (N_11701,N_11254,N_11094);
xor U11702 (N_11702,N_11158,N_11312);
nor U11703 (N_11703,N_11037,N_11123);
nand U11704 (N_11704,N_11377,N_11323);
nor U11705 (N_11705,N_11384,N_11423);
or U11706 (N_11706,N_11295,N_11010);
and U11707 (N_11707,N_11378,N_11296);
and U11708 (N_11708,N_11155,N_11398);
nand U11709 (N_11709,N_11429,N_11134);
nor U11710 (N_11710,N_11441,N_11172);
xor U11711 (N_11711,N_11124,N_11177);
xor U11712 (N_11712,N_11069,N_11153);
or U11713 (N_11713,N_11145,N_11116);
and U11714 (N_11714,N_11102,N_11111);
nor U11715 (N_11715,N_11219,N_11444);
nand U11716 (N_11716,N_11179,N_11410);
and U11717 (N_11717,N_11103,N_11020);
xnor U11718 (N_11718,N_11068,N_11435);
nand U11719 (N_11719,N_11148,N_11426);
and U11720 (N_11720,N_11181,N_11362);
nand U11721 (N_11721,N_11477,N_11376);
nor U11722 (N_11722,N_11415,N_11487);
and U11723 (N_11723,N_11077,N_11325);
nand U11724 (N_11724,N_11038,N_11496);
and U11725 (N_11725,N_11144,N_11448);
nor U11726 (N_11726,N_11078,N_11419);
xnor U11727 (N_11727,N_11352,N_11149);
nand U11728 (N_11728,N_11261,N_11164);
xor U11729 (N_11729,N_11313,N_11363);
nand U11730 (N_11730,N_11005,N_11075);
nand U11731 (N_11731,N_11326,N_11468);
xnor U11732 (N_11732,N_11293,N_11456);
xnor U11733 (N_11733,N_11427,N_11280);
xor U11734 (N_11734,N_11105,N_11314);
and U11735 (N_11735,N_11365,N_11081);
nor U11736 (N_11736,N_11214,N_11057);
nand U11737 (N_11737,N_11416,N_11409);
and U11738 (N_11738,N_11303,N_11266);
nand U11739 (N_11739,N_11169,N_11483);
nor U11740 (N_11740,N_11033,N_11478);
nand U11741 (N_11741,N_11334,N_11372);
nor U11742 (N_11742,N_11218,N_11152);
xnor U11743 (N_11743,N_11096,N_11226);
nor U11744 (N_11744,N_11108,N_11373);
and U11745 (N_11745,N_11388,N_11242);
xnor U11746 (N_11746,N_11223,N_11405);
and U11747 (N_11747,N_11494,N_11178);
nor U11748 (N_11748,N_11067,N_11490);
nor U11749 (N_11749,N_11224,N_11343);
nand U11750 (N_11750,N_11387,N_11159);
and U11751 (N_11751,N_11054,N_11400);
and U11752 (N_11752,N_11314,N_11218);
and U11753 (N_11753,N_11336,N_11393);
nor U11754 (N_11754,N_11132,N_11458);
nor U11755 (N_11755,N_11201,N_11493);
and U11756 (N_11756,N_11470,N_11418);
nand U11757 (N_11757,N_11455,N_11159);
or U11758 (N_11758,N_11011,N_11121);
or U11759 (N_11759,N_11171,N_11057);
nor U11760 (N_11760,N_11429,N_11016);
nor U11761 (N_11761,N_11030,N_11266);
nor U11762 (N_11762,N_11368,N_11471);
nand U11763 (N_11763,N_11206,N_11177);
xor U11764 (N_11764,N_11244,N_11025);
or U11765 (N_11765,N_11492,N_11118);
nand U11766 (N_11766,N_11133,N_11227);
xnor U11767 (N_11767,N_11087,N_11275);
or U11768 (N_11768,N_11185,N_11340);
or U11769 (N_11769,N_11476,N_11444);
nand U11770 (N_11770,N_11089,N_11481);
or U11771 (N_11771,N_11323,N_11003);
xnor U11772 (N_11772,N_11288,N_11064);
nor U11773 (N_11773,N_11433,N_11060);
and U11774 (N_11774,N_11410,N_11487);
xor U11775 (N_11775,N_11112,N_11404);
nand U11776 (N_11776,N_11237,N_11069);
nor U11777 (N_11777,N_11329,N_11461);
xnor U11778 (N_11778,N_11374,N_11077);
nor U11779 (N_11779,N_11461,N_11062);
nor U11780 (N_11780,N_11192,N_11440);
nand U11781 (N_11781,N_11229,N_11326);
nor U11782 (N_11782,N_11473,N_11017);
nor U11783 (N_11783,N_11117,N_11082);
and U11784 (N_11784,N_11239,N_11202);
nand U11785 (N_11785,N_11142,N_11260);
nand U11786 (N_11786,N_11223,N_11240);
and U11787 (N_11787,N_11394,N_11365);
and U11788 (N_11788,N_11128,N_11019);
or U11789 (N_11789,N_11005,N_11473);
nand U11790 (N_11790,N_11196,N_11433);
xnor U11791 (N_11791,N_11429,N_11235);
and U11792 (N_11792,N_11137,N_11429);
nand U11793 (N_11793,N_11397,N_11149);
xnor U11794 (N_11794,N_11356,N_11237);
nor U11795 (N_11795,N_11248,N_11000);
xnor U11796 (N_11796,N_11135,N_11072);
xnor U11797 (N_11797,N_11134,N_11367);
nor U11798 (N_11798,N_11099,N_11158);
nor U11799 (N_11799,N_11415,N_11257);
nor U11800 (N_11800,N_11406,N_11239);
nor U11801 (N_11801,N_11278,N_11140);
and U11802 (N_11802,N_11157,N_11035);
nand U11803 (N_11803,N_11357,N_11074);
or U11804 (N_11804,N_11302,N_11186);
nand U11805 (N_11805,N_11489,N_11289);
or U11806 (N_11806,N_11247,N_11352);
nand U11807 (N_11807,N_11384,N_11478);
nor U11808 (N_11808,N_11325,N_11214);
nor U11809 (N_11809,N_11297,N_11436);
nand U11810 (N_11810,N_11004,N_11247);
xor U11811 (N_11811,N_11048,N_11185);
nand U11812 (N_11812,N_11361,N_11074);
xor U11813 (N_11813,N_11064,N_11392);
xor U11814 (N_11814,N_11410,N_11279);
nor U11815 (N_11815,N_11265,N_11278);
and U11816 (N_11816,N_11473,N_11132);
nand U11817 (N_11817,N_11011,N_11492);
nand U11818 (N_11818,N_11398,N_11442);
or U11819 (N_11819,N_11259,N_11213);
nor U11820 (N_11820,N_11377,N_11258);
xnor U11821 (N_11821,N_11060,N_11091);
or U11822 (N_11822,N_11361,N_11338);
nor U11823 (N_11823,N_11474,N_11088);
and U11824 (N_11824,N_11129,N_11084);
xnor U11825 (N_11825,N_11055,N_11426);
or U11826 (N_11826,N_11024,N_11295);
or U11827 (N_11827,N_11335,N_11288);
xor U11828 (N_11828,N_11135,N_11423);
and U11829 (N_11829,N_11246,N_11342);
xor U11830 (N_11830,N_11058,N_11387);
xnor U11831 (N_11831,N_11206,N_11307);
nand U11832 (N_11832,N_11306,N_11005);
and U11833 (N_11833,N_11429,N_11348);
nor U11834 (N_11834,N_11229,N_11184);
and U11835 (N_11835,N_11305,N_11103);
xor U11836 (N_11836,N_11002,N_11260);
xor U11837 (N_11837,N_11006,N_11260);
and U11838 (N_11838,N_11346,N_11412);
nand U11839 (N_11839,N_11113,N_11046);
or U11840 (N_11840,N_11198,N_11414);
xor U11841 (N_11841,N_11398,N_11326);
xnor U11842 (N_11842,N_11236,N_11199);
xor U11843 (N_11843,N_11197,N_11247);
nand U11844 (N_11844,N_11443,N_11476);
and U11845 (N_11845,N_11317,N_11200);
xor U11846 (N_11846,N_11271,N_11022);
nand U11847 (N_11847,N_11015,N_11469);
or U11848 (N_11848,N_11458,N_11090);
and U11849 (N_11849,N_11350,N_11438);
nand U11850 (N_11850,N_11244,N_11447);
nor U11851 (N_11851,N_11082,N_11366);
nor U11852 (N_11852,N_11251,N_11262);
nand U11853 (N_11853,N_11480,N_11370);
and U11854 (N_11854,N_11480,N_11488);
or U11855 (N_11855,N_11492,N_11261);
or U11856 (N_11856,N_11156,N_11152);
xnor U11857 (N_11857,N_11314,N_11462);
nor U11858 (N_11858,N_11117,N_11195);
xor U11859 (N_11859,N_11285,N_11311);
nor U11860 (N_11860,N_11241,N_11051);
xnor U11861 (N_11861,N_11364,N_11380);
nand U11862 (N_11862,N_11132,N_11232);
and U11863 (N_11863,N_11368,N_11437);
and U11864 (N_11864,N_11428,N_11429);
xnor U11865 (N_11865,N_11390,N_11417);
nand U11866 (N_11866,N_11075,N_11345);
nor U11867 (N_11867,N_11481,N_11095);
and U11868 (N_11868,N_11264,N_11062);
nand U11869 (N_11869,N_11065,N_11333);
nor U11870 (N_11870,N_11423,N_11392);
nand U11871 (N_11871,N_11304,N_11164);
and U11872 (N_11872,N_11345,N_11351);
and U11873 (N_11873,N_11214,N_11130);
and U11874 (N_11874,N_11279,N_11091);
or U11875 (N_11875,N_11236,N_11248);
and U11876 (N_11876,N_11105,N_11384);
xnor U11877 (N_11877,N_11212,N_11166);
and U11878 (N_11878,N_11488,N_11036);
nand U11879 (N_11879,N_11171,N_11212);
or U11880 (N_11880,N_11208,N_11097);
xor U11881 (N_11881,N_11427,N_11403);
or U11882 (N_11882,N_11038,N_11493);
xnor U11883 (N_11883,N_11011,N_11389);
xor U11884 (N_11884,N_11343,N_11253);
or U11885 (N_11885,N_11118,N_11388);
xnor U11886 (N_11886,N_11179,N_11297);
nor U11887 (N_11887,N_11178,N_11300);
or U11888 (N_11888,N_11054,N_11484);
or U11889 (N_11889,N_11219,N_11357);
or U11890 (N_11890,N_11415,N_11079);
xnor U11891 (N_11891,N_11377,N_11421);
nand U11892 (N_11892,N_11110,N_11074);
and U11893 (N_11893,N_11268,N_11016);
nor U11894 (N_11894,N_11493,N_11417);
xor U11895 (N_11895,N_11023,N_11413);
nor U11896 (N_11896,N_11407,N_11077);
and U11897 (N_11897,N_11017,N_11144);
nand U11898 (N_11898,N_11111,N_11277);
nor U11899 (N_11899,N_11373,N_11353);
nor U11900 (N_11900,N_11394,N_11054);
nor U11901 (N_11901,N_11113,N_11012);
or U11902 (N_11902,N_11180,N_11305);
or U11903 (N_11903,N_11068,N_11443);
xnor U11904 (N_11904,N_11046,N_11416);
or U11905 (N_11905,N_11305,N_11265);
xor U11906 (N_11906,N_11308,N_11247);
or U11907 (N_11907,N_11188,N_11292);
nor U11908 (N_11908,N_11255,N_11002);
xor U11909 (N_11909,N_11298,N_11353);
nor U11910 (N_11910,N_11447,N_11492);
nand U11911 (N_11911,N_11099,N_11220);
nand U11912 (N_11912,N_11128,N_11240);
nor U11913 (N_11913,N_11199,N_11287);
nand U11914 (N_11914,N_11463,N_11151);
nand U11915 (N_11915,N_11123,N_11374);
xor U11916 (N_11916,N_11127,N_11002);
nand U11917 (N_11917,N_11497,N_11141);
xnor U11918 (N_11918,N_11046,N_11395);
and U11919 (N_11919,N_11367,N_11257);
and U11920 (N_11920,N_11417,N_11348);
and U11921 (N_11921,N_11098,N_11323);
nor U11922 (N_11922,N_11116,N_11275);
and U11923 (N_11923,N_11239,N_11473);
xor U11924 (N_11924,N_11202,N_11370);
nand U11925 (N_11925,N_11385,N_11465);
nor U11926 (N_11926,N_11072,N_11490);
nor U11927 (N_11927,N_11475,N_11016);
nand U11928 (N_11928,N_11092,N_11042);
or U11929 (N_11929,N_11376,N_11491);
or U11930 (N_11930,N_11026,N_11221);
and U11931 (N_11931,N_11092,N_11352);
nand U11932 (N_11932,N_11238,N_11243);
and U11933 (N_11933,N_11302,N_11416);
xnor U11934 (N_11934,N_11045,N_11138);
and U11935 (N_11935,N_11170,N_11244);
or U11936 (N_11936,N_11348,N_11145);
nand U11937 (N_11937,N_11088,N_11330);
or U11938 (N_11938,N_11063,N_11380);
and U11939 (N_11939,N_11341,N_11118);
and U11940 (N_11940,N_11431,N_11079);
or U11941 (N_11941,N_11261,N_11195);
or U11942 (N_11942,N_11173,N_11061);
nor U11943 (N_11943,N_11080,N_11453);
or U11944 (N_11944,N_11310,N_11389);
and U11945 (N_11945,N_11337,N_11065);
nor U11946 (N_11946,N_11410,N_11217);
or U11947 (N_11947,N_11190,N_11350);
nand U11948 (N_11948,N_11378,N_11209);
and U11949 (N_11949,N_11312,N_11369);
and U11950 (N_11950,N_11363,N_11090);
and U11951 (N_11951,N_11051,N_11137);
xor U11952 (N_11952,N_11086,N_11401);
nor U11953 (N_11953,N_11424,N_11076);
or U11954 (N_11954,N_11099,N_11180);
nand U11955 (N_11955,N_11292,N_11437);
or U11956 (N_11956,N_11017,N_11172);
nand U11957 (N_11957,N_11040,N_11086);
or U11958 (N_11958,N_11228,N_11411);
nor U11959 (N_11959,N_11181,N_11358);
or U11960 (N_11960,N_11169,N_11385);
and U11961 (N_11961,N_11180,N_11357);
nand U11962 (N_11962,N_11459,N_11440);
nand U11963 (N_11963,N_11027,N_11165);
and U11964 (N_11964,N_11291,N_11030);
or U11965 (N_11965,N_11190,N_11296);
nand U11966 (N_11966,N_11432,N_11174);
nand U11967 (N_11967,N_11403,N_11232);
nor U11968 (N_11968,N_11061,N_11002);
nor U11969 (N_11969,N_11348,N_11045);
and U11970 (N_11970,N_11336,N_11212);
and U11971 (N_11971,N_11426,N_11300);
or U11972 (N_11972,N_11084,N_11364);
and U11973 (N_11973,N_11478,N_11059);
nor U11974 (N_11974,N_11208,N_11360);
nor U11975 (N_11975,N_11464,N_11444);
or U11976 (N_11976,N_11050,N_11365);
nand U11977 (N_11977,N_11404,N_11256);
nor U11978 (N_11978,N_11359,N_11174);
or U11979 (N_11979,N_11244,N_11078);
and U11980 (N_11980,N_11137,N_11444);
nor U11981 (N_11981,N_11143,N_11236);
or U11982 (N_11982,N_11328,N_11387);
and U11983 (N_11983,N_11090,N_11472);
nor U11984 (N_11984,N_11244,N_11347);
and U11985 (N_11985,N_11188,N_11438);
nand U11986 (N_11986,N_11040,N_11167);
xor U11987 (N_11987,N_11096,N_11062);
nor U11988 (N_11988,N_11324,N_11100);
nand U11989 (N_11989,N_11085,N_11329);
xor U11990 (N_11990,N_11118,N_11276);
nor U11991 (N_11991,N_11150,N_11197);
or U11992 (N_11992,N_11329,N_11074);
or U11993 (N_11993,N_11122,N_11343);
nor U11994 (N_11994,N_11164,N_11166);
or U11995 (N_11995,N_11357,N_11028);
nor U11996 (N_11996,N_11059,N_11436);
nand U11997 (N_11997,N_11372,N_11326);
nor U11998 (N_11998,N_11105,N_11159);
nand U11999 (N_11999,N_11157,N_11200);
or U12000 (N_12000,N_11566,N_11712);
and U12001 (N_12001,N_11982,N_11599);
nand U12002 (N_12002,N_11502,N_11877);
nand U12003 (N_12003,N_11521,N_11578);
xnor U12004 (N_12004,N_11680,N_11682);
and U12005 (N_12005,N_11872,N_11823);
or U12006 (N_12006,N_11933,N_11814);
and U12007 (N_12007,N_11840,N_11978);
and U12008 (N_12008,N_11824,N_11544);
xor U12009 (N_12009,N_11861,N_11790);
nand U12010 (N_12010,N_11789,N_11985);
and U12011 (N_12011,N_11621,N_11703);
nor U12012 (N_12012,N_11768,N_11618);
nor U12013 (N_12013,N_11857,N_11896);
nand U12014 (N_12014,N_11555,N_11633);
or U12015 (N_12015,N_11788,N_11670);
xor U12016 (N_12016,N_11734,N_11523);
nor U12017 (N_12017,N_11837,N_11846);
nor U12018 (N_12018,N_11783,N_11802);
nand U12019 (N_12019,N_11809,N_11808);
or U12020 (N_12020,N_11679,N_11644);
or U12021 (N_12021,N_11554,N_11708);
and U12022 (N_12022,N_11606,N_11540);
nor U12023 (N_12023,N_11864,N_11818);
or U12024 (N_12024,N_11647,N_11649);
nand U12025 (N_12025,N_11795,N_11828);
or U12026 (N_12026,N_11505,N_11968);
or U12027 (N_12027,N_11582,N_11537);
nand U12028 (N_12028,N_11817,N_11662);
xnor U12029 (N_12029,N_11605,N_11929);
and U12030 (N_12030,N_11799,N_11671);
or U12031 (N_12031,N_11518,N_11743);
nand U12032 (N_12032,N_11683,N_11742);
or U12033 (N_12033,N_11884,N_11515);
nand U12034 (N_12034,N_11695,N_11794);
xor U12035 (N_12035,N_11776,N_11863);
nor U12036 (N_12036,N_11765,N_11520);
and U12037 (N_12037,N_11858,N_11890);
and U12038 (N_12038,N_11586,N_11673);
nand U12039 (N_12039,N_11563,N_11653);
nand U12040 (N_12040,N_11562,N_11851);
xor U12041 (N_12041,N_11980,N_11951);
or U12042 (N_12042,N_11592,N_11995);
nand U12043 (N_12043,N_11888,N_11661);
nor U12044 (N_12044,N_11845,N_11865);
xor U12045 (N_12045,N_11902,N_11559);
nor U12046 (N_12046,N_11767,N_11862);
nor U12047 (N_12047,N_11587,N_11882);
or U12048 (N_12048,N_11964,N_11732);
nand U12049 (N_12049,N_11741,N_11623);
nor U12050 (N_12050,N_11950,N_11906);
and U12051 (N_12051,N_11519,N_11651);
or U12052 (N_12052,N_11829,N_11745);
or U12053 (N_12053,N_11833,N_11836);
or U12054 (N_12054,N_11539,N_11739);
xnor U12055 (N_12055,N_11590,N_11760);
nor U12056 (N_12056,N_11634,N_11686);
and U12057 (N_12057,N_11860,N_11979);
nand U12058 (N_12058,N_11992,N_11855);
nand U12059 (N_12059,N_11900,N_11782);
and U12060 (N_12060,N_11927,N_11875);
nor U12061 (N_12061,N_11904,N_11804);
and U12062 (N_12062,N_11677,N_11800);
xor U12063 (N_12063,N_11674,N_11556);
xnor U12064 (N_12064,N_11735,N_11572);
xor U12065 (N_12065,N_11819,N_11645);
or U12066 (N_12066,N_11959,N_11758);
nand U12067 (N_12067,N_11666,N_11748);
nor U12068 (N_12068,N_11928,N_11763);
nand U12069 (N_12069,N_11567,N_11785);
xor U12070 (N_12070,N_11962,N_11723);
nand U12071 (N_12071,N_11963,N_11910);
nor U12072 (N_12072,N_11803,N_11919);
xor U12073 (N_12073,N_11898,N_11622);
xnor U12074 (N_12074,N_11917,N_11759);
nand U12075 (N_12075,N_11841,N_11847);
and U12076 (N_12076,N_11905,N_11697);
nand U12077 (N_12077,N_11895,N_11635);
nand U12078 (N_12078,N_11969,N_11557);
and U12079 (N_12079,N_11810,N_11603);
nor U12080 (N_12080,N_11775,N_11564);
or U12081 (N_12081,N_11757,N_11988);
xor U12082 (N_12082,N_11774,N_11692);
and U12083 (N_12083,N_11991,N_11584);
and U12084 (N_12084,N_11798,N_11663);
or U12085 (N_12085,N_11713,N_11528);
and U12086 (N_12086,N_11573,N_11656);
nand U12087 (N_12087,N_11601,N_11591);
nand U12088 (N_12088,N_11730,N_11630);
nor U12089 (N_12089,N_11721,N_11657);
xor U12090 (N_12090,N_11580,N_11533);
or U12091 (N_12091,N_11737,N_11812);
nor U12092 (N_12092,N_11999,N_11893);
xnor U12093 (N_12093,N_11655,N_11935);
nand U12094 (N_12094,N_11838,N_11733);
xnor U12095 (N_12095,N_11705,N_11638);
xnor U12096 (N_12096,N_11957,N_11827);
nor U12097 (N_12097,N_11853,N_11527);
nand U12098 (N_12098,N_11848,N_11772);
and U12099 (N_12099,N_11835,N_11507);
xor U12100 (N_12100,N_11652,N_11639);
xnor U12101 (N_12101,N_11522,N_11690);
xor U12102 (N_12102,N_11920,N_11922);
and U12103 (N_12103,N_11719,N_11553);
nand U12104 (N_12104,N_11543,N_11883);
nand U12105 (N_12105,N_11524,N_11706);
or U12106 (N_12106,N_11948,N_11820);
xor U12107 (N_12107,N_11725,N_11932);
nand U12108 (N_12108,N_11547,N_11628);
xor U12109 (N_12109,N_11854,N_11736);
or U12110 (N_12110,N_11984,N_11756);
xnor U12111 (N_12111,N_11546,N_11873);
nor U12112 (N_12112,N_11830,N_11576);
or U12113 (N_12113,N_11608,N_11811);
and U12114 (N_12114,N_11887,N_11921);
or U12115 (N_12115,N_11755,N_11541);
and U12116 (N_12116,N_11616,N_11512);
xor U12117 (N_12117,N_11629,N_11886);
and U12118 (N_12118,N_11668,N_11958);
or U12119 (N_12119,N_11869,N_11825);
nor U12120 (N_12120,N_11728,N_11571);
xnor U12121 (N_12121,N_11891,N_11570);
xnor U12122 (N_12122,N_11870,N_11624);
or U12123 (N_12123,N_11844,N_11826);
and U12124 (N_12124,N_11579,N_11642);
and U12125 (N_12125,N_11611,N_11952);
nor U12126 (N_12126,N_11807,N_11947);
xor U12127 (N_12127,N_11577,N_11646);
nor U12128 (N_12128,N_11698,N_11504);
nor U12129 (N_12129,N_11761,N_11640);
or U12130 (N_12130,N_11878,N_11913);
xor U12131 (N_12131,N_11797,N_11648);
nand U12132 (N_12132,N_11500,N_11583);
or U12133 (N_12133,N_11778,N_11724);
nor U12134 (N_12134,N_11977,N_11746);
nor U12135 (N_12135,N_11509,N_11970);
nor U12136 (N_12136,N_11720,N_11931);
nor U12137 (N_12137,N_11923,N_11604);
or U12138 (N_12138,N_11868,N_11822);
xnor U12139 (N_12139,N_11531,N_11702);
or U12140 (N_12140,N_11626,N_11912);
nor U12141 (N_12141,N_11770,N_11843);
xor U12142 (N_12142,N_11766,N_11994);
and U12143 (N_12143,N_11612,N_11687);
or U12144 (N_12144,N_11955,N_11976);
nor U12145 (N_12145,N_11796,N_11613);
nor U12146 (N_12146,N_11598,N_11967);
or U12147 (N_12147,N_11997,N_11946);
nor U12148 (N_12148,N_11525,N_11619);
nand U12149 (N_12149,N_11691,N_11609);
and U12150 (N_12150,N_11729,N_11777);
and U12151 (N_12151,N_11696,N_11986);
and U12152 (N_12152,N_11936,N_11529);
xnor U12153 (N_12153,N_11908,N_11918);
and U12154 (N_12154,N_11569,N_11753);
nor U12155 (N_12155,N_11784,N_11615);
and U12156 (N_12156,N_11676,N_11889);
or U12157 (N_12157,N_11538,N_11740);
nor U12158 (N_12158,N_11801,N_11542);
or U12159 (N_12159,N_11773,N_11602);
nand U12160 (N_12160,N_11975,N_11506);
xor U12161 (N_12161,N_11596,N_11954);
or U12162 (N_12162,N_11791,N_11575);
or U12163 (N_12163,N_11953,N_11530);
nand U12164 (N_12164,N_11534,N_11793);
nor U12165 (N_12165,N_11514,N_11727);
and U12166 (N_12166,N_11558,N_11924);
and U12167 (N_12167,N_11709,N_11658);
xnor U12168 (N_12168,N_11508,N_11595);
xor U12169 (N_12169,N_11659,N_11548);
xnor U12170 (N_12170,N_11942,N_11675);
or U12171 (N_12171,N_11714,N_11627);
nor U12172 (N_12172,N_11961,N_11956);
and U12173 (N_12173,N_11834,N_11589);
or U12174 (N_12174,N_11684,N_11832);
nor U12175 (N_12175,N_11806,N_11916);
nand U12176 (N_12176,N_11856,N_11867);
or U12177 (N_12177,N_11532,N_11925);
and U12178 (N_12178,N_11937,N_11664);
or U12179 (N_12179,N_11915,N_11701);
nor U12180 (N_12180,N_11744,N_11849);
xor U12181 (N_12181,N_11535,N_11940);
xnor U12182 (N_12182,N_11780,N_11769);
nor U12183 (N_12183,N_11501,N_11989);
xnor U12184 (N_12184,N_11551,N_11631);
and U12185 (N_12185,N_11694,N_11930);
nand U12186 (N_12186,N_11786,N_11568);
xor U12187 (N_12187,N_11839,N_11667);
and U12188 (N_12188,N_11688,N_11938);
and U12189 (N_12189,N_11711,N_11911);
and U12190 (N_12190,N_11901,N_11715);
xor U12191 (N_12191,N_11973,N_11718);
or U12192 (N_12192,N_11636,N_11998);
xor U12193 (N_12193,N_11749,N_11678);
nor U12194 (N_12194,N_11771,N_11850);
nand U12195 (N_12195,N_11752,N_11750);
nand U12196 (N_12196,N_11874,N_11876);
nand U12197 (N_12197,N_11960,N_11536);
xor U12198 (N_12198,N_11710,N_11892);
nor U12199 (N_12199,N_11972,N_11754);
nand U12200 (N_12200,N_11894,N_11821);
nor U12201 (N_12201,N_11641,N_11510);
xnor U12202 (N_12202,N_11614,N_11593);
or U12203 (N_12203,N_11731,N_11738);
nor U12204 (N_12204,N_11805,N_11944);
and U12205 (N_12205,N_11859,N_11909);
or U12206 (N_12206,N_11971,N_11665);
nor U12207 (N_12207,N_11585,N_11871);
or U12208 (N_12208,N_11966,N_11813);
nand U12209 (N_12209,N_11643,N_11654);
and U12210 (N_12210,N_11747,N_11685);
nand U12211 (N_12211,N_11594,N_11625);
and U12212 (N_12212,N_11517,N_11600);
xnor U12213 (N_12213,N_11897,N_11764);
nand U12214 (N_12214,N_11899,N_11693);
xor U12215 (N_12215,N_11751,N_11511);
and U12216 (N_12216,N_11607,N_11700);
and U12217 (N_12217,N_11545,N_11669);
and U12218 (N_12218,N_11974,N_11717);
nor U12219 (N_12219,N_11939,N_11610);
nand U12220 (N_12220,N_11852,N_11632);
xnor U12221 (N_12221,N_11581,N_11707);
nand U12222 (N_12222,N_11516,N_11549);
and U12223 (N_12223,N_11503,N_11983);
nand U12224 (N_12224,N_11949,N_11934);
and U12225 (N_12225,N_11866,N_11816);
or U12226 (N_12226,N_11704,N_11574);
nor U12227 (N_12227,N_11650,N_11617);
nor U12228 (N_12228,N_11981,N_11681);
nor U12229 (N_12229,N_11990,N_11565);
or U12230 (N_12230,N_11699,N_11987);
or U12231 (N_12231,N_11993,N_11660);
nor U12232 (N_12232,N_11880,N_11945);
xor U12233 (N_12233,N_11879,N_11965);
and U12234 (N_12234,N_11903,N_11513);
nor U12235 (N_12235,N_11842,N_11941);
nor U12236 (N_12236,N_11726,N_11637);
or U12237 (N_12237,N_11620,N_11526);
or U12238 (N_12238,N_11781,N_11792);
nand U12239 (N_12239,N_11779,N_11996);
or U12240 (N_12240,N_11907,N_11672);
xnor U12241 (N_12241,N_11716,N_11885);
and U12242 (N_12242,N_11943,N_11588);
nor U12243 (N_12243,N_11560,N_11914);
nor U12244 (N_12244,N_11815,N_11787);
or U12245 (N_12245,N_11550,N_11831);
nor U12246 (N_12246,N_11689,N_11881);
and U12247 (N_12247,N_11552,N_11597);
or U12248 (N_12248,N_11762,N_11926);
xnor U12249 (N_12249,N_11722,N_11561);
or U12250 (N_12250,N_11954,N_11676);
and U12251 (N_12251,N_11831,N_11952);
nand U12252 (N_12252,N_11716,N_11800);
nor U12253 (N_12253,N_11776,N_11535);
or U12254 (N_12254,N_11601,N_11731);
nor U12255 (N_12255,N_11570,N_11994);
nor U12256 (N_12256,N_11536,N_11513);
and U12257 (N_12257,N_11618,N_11685);
nand U12258 (N_12258,N_11688,N_11599);
and U12259 (N_12259,N_11569,N_11616);
nor U12260 (N_12260,N_11897,N_11520);
or U12261 (N_12261,N_11668,N_11992);
xnor U12262 (N_12262,N_11712,N_11990);
nor U12263 (N_12263,N_11908,N_11669);
nand U12264 (N_12264,N_11938,N_11611);
xnor U12265 (N_12265,N_11810,N_11858);
or U12266 (N_12266,N_11912,N_11669);
nor U12267 (N_12267,N_11754,N_11725);
and U12268 (N_12268,N_11755,N_11836);
xnor U12269 (N_12269,N_11760,N_11670);
nand U12270 (N_12270,N_11966,N_11649);
or U12271 (N_12271,N_11506,N_11909);
or U12272 (N_12272,N_11765,N_11525);
and U12273 (N_12273,N_11785,N_11789);
and U12274 (N_12274,N_11815,N_11838);
nand U12275 (N_12275,N_11931,N_11861);
nand U12276 (N_12276,N_11812,N_11934);
or U12277 (N_12277,N_11814,N_11593);
or U12278 (N_12278,N_11563,N_11646);
xnor U12279 (N_12279,N_11691,N_11571);
nor U12280 (N_12280,N_11783,N_11553);
and U12281 (N_12281,N_11906,N_11857);
nor U12282 (N_12282,N_11763,N_11824);
and U12283 (N_12283,N_11912,N_11676);
or U12284 (N_12284,N_11825,N_11748);
and U12285 (N_12285,N_11785,N_11984);
nor U12286 (N_12286,N_11753,N_11512);
xnor U12287 (N_12287,N_11950,N_11794);
nor U12288 (N_12288,N_11716,N_11824);
or U12289 (N_12289,N_11581,N_11738);
xnor U12290 (N_12290,N_11887,N_11504);
and U12291 (N_12291,N_11554,N_11657);
nor U12292 (N_12292,N_11750,N_11759);
or U12293 (N_12293,N_11606,N_11582);
or U12294 (N_12294,N_11540,N_11928);
nand U12295 (N_12295,N_11893,N_11675);
and U12296 (N_12296,N_11927,N_11527);
nor U12297 (N_12297,N_11683,N_11751);
nor U12298 (N_12298,N_11888,N_11932);
or U12299 (N_12299,N_11864,N_11638);
or U12300 (N_12300,N_11761,N_11501);
and U12301 (N_12301,N_11876,N_11907);
and U12302 (N_12302,N_11774,N_11799);
or U12303 (N_12303,N_11892,N_11871);
nand U12304 (N_12304,N_11733,N_11721);
or U12305 (N_12305,N_11571,N_11626);
xnor U12306 (N_12306,N_11524,N_11717);
and U12307 (N_12307,N_11963,N_11649);
nor U12308 (N_12308,N_11741,N_11931);
or U12309 (N_12309,N_11692,N_11899);
xor U12310 (N_12310,N_11702,N_11988);
xor U12311 (N_12311,N_11874,N_11828);
or U12312 (N_12312,N_11869,N_11543);
and U12313 (N_12313,N_11725,N_11638);
or U12314 (N_12314,N_11504,N_11670);
nor U12315 (N_12315,N_11933,N_11695);
or U12316 (N_12316,N_11592,N_11786);
nand U12317 (N_12317,N_11957,N_11653);
or U12318 (N_12318,N_11735,N_11505);
or U12319 (N_12319,N_11827,N_11578);
xor U12320 (N_12320,N_11833,N_11893);
nand U12321 (N_12321,N_11763,N_11663);
nand U12322 (N_12322,N_11700,N_11669);
or U12323 (N_12323,N_11660,N_11910);
or U12324 (N_12324,N_11534,N_11540);
xnor U12325 (N_12325,N_11973,N_11810);
xnor U12326 (N_12326,N_11912,N_11901);
and U12327 (N_12327,N_11879,N_11863);
or U12328 (N_12328,N_11791,N_11626);
or U12329 (N_12329,N_11712,N_11844);
xor U12330 (N_12330,N_11644,N_11670);
xnor U12331 (N_12331,N_11876,N_11656);
or U12332 (N_12332,N_11920,N_11569);
nand U12333 (N_12333,N_11686,N_11508);
nor U12334 (N_12334,N_11833,N_11581);
or U12335 (N_12335,N_11753,N_11970);
xor U12336 (N_12336,N_11640,N_11579);
and U12337 (N_12337,N_11651,N_11889);
xnor U12338 (N_12338,N_11583,N_11732);
nand U12339 (N_12339,N_11861,N_11694);
and U12340 (N_12340,N_11653,N_11970);
xnor U12341 (N_12341,N_11593,N_11961);
and U12342 (N_12342,N_11733,N_11822);
and U12343 (N_12343,N_11605,N_11798);
nor U12344 (N_12344,N_11884,N_11591);
or U12345 (N_12345,N_11677,N_11601);
nor U12346 (N_12346,N_11729,N_11595);
xnor U12347 (N_12347,N_11980,N_11956);
nor U12348 (N_12348,N_11505,N_11687);
or U12349 (N_12349,N_11898,N_11787);
nor U12350 (N_12350,N_11587,N_11822);
or U12351 (N_12351,N_11795,N_11805);
nor U12352 (N_12352,N_11810,N_11996);
or U12353 (N_12353,N_11987,N_11998);
xor U12354 (N_12354,N_11601,N_11740);
or U12355 (N_12355,N_11565,N_11665);
nor U12356 (N_12356,N_11785,N_11688);
or U12357 (N_12357,N_11504,N_11968);
and U12358 (N_12358,N_11789,N_11819);
nor U12359 (N_12359,N_11728,N_11538);
nand U12360 (N_12360,N_11813,N_11861);
or U12361 (N_12361,N_11717,N_11744);
and U12362 (N_12362,N_11660,N_11519);
xnor U12363 (N_12363,N_11970,N_11973);
or U12364 (N_12364,N_11760,N_11604);
nor U12365 (N_12365,N_11935,N_11931);
nand U12366 (N_12366,N_11772,N_11618);
or U12367 (N_12367,N_11799,N_11900);
nand U12368 (N_12368,N_11730,N_11980);
xor U12369 (N_12369,N_11885,N_11503);
and U12370 (N_12370,N_11549,N_11712);
or U12371 (N_12371,N_11697,N_11629);
xor U12372 (N_12372,N_11833,N_11689);
nand U12373 (N_12373,N_11885,N_11822);
or U12374 (N_12374,N_11951,N_11634);
or U12375 (N_12375,N_11970,N_11729);
and U12376 (N_12376,N_11656,N_11747);
nand U12377 (N_12377,N_11829,N_11896);
xnor U12378 (N_12378,N_11653,N_11601);
and U12379 (N_12379,N_11942,N_11810);
and U12380 (N_12380,N_11727,N_11899);
and U12381 (N_12381,N_11587,N_11573);
xor U12382 (N_12382,N_11945,N_11778);
nand U12383 (N_12383,N_11967,N_11926);
xnor U12384 (N_12384,N_11833,N_11845);
or U12385 (N_12385,N_11854,N_11812);
and U12386 (N_12386,N_11529,N_11747);
xnor U12387 (N_12387,N_11995,N_11967);
xor U12388 (N_12388,N_11746,N_11654);
nand U12389 (N_12389,N_11846,N_11657);
nand U12390 (N_12390,N_11712,N_11841);
and U12391 (N_12391,N_11774,N_11902);
xor U12392 (N_12392,N_11909,N_11918);
or U12393 (N_12393,N_11954,N_11915);
nor U12394 (N_12394,N_11847,N_11538);
xor U12395 (N_12395,N_11773,N_11524);
xor U12396 (N_12396,N_11950,N_11902);
or U12397 (N_12397,N_11576,N_11875);
or U12398 (N_12398,N_11597,N_11728);
and U12399 (N_12399,N_11592,N_11740);
nor U12400 (N_12400,N_11903,N_11522);
or U12401 (N_12401,N_11854,N_11920);
xor U12402 (N_12402,N_11848,N_11598);
and U12403 (N_12403,N_11950,N_11604);
xor U12404 (N_12404,N_11723,N_11933);
and U12405 (N_12405,N_11533,N_11966);
or U12406 (N_12406,N_11778,N_11942);
xnor U12407 (N_12407,N_11988,N_11981);
and U12408 (N_12408,N_11981,N_11943);
and U12409 (N_12409,N_11601,N_11645);
xor U12410 (N_12410,N_11527,N_11713);
nand U12411 (N_12411,N_11589,N_11705);
nand U12412 (N_12412,N_11638,N_11966);
or U12413 (N_12413,N_11953,N_11763);
xnor U12414 (N_12414,N_11923,N_11883);
nor U12415 (N_12415,N_11526,N_11978);
nand U12416 (N_12416,N_11773,N_11803);
and U12417 (N_12417,N_11670,N_11520);
and U12418 (N_12418,N_11590,N_11688);
nor U12419 (N_12419,N_11819,N_11513);
and U12420 (N_12420,N_11531,N_11890);
or U12421 (N_12421,N_11624,N_11556);
nand U12422 (N_12422,N_11854,N_11869);
or U12423 (N_12423,N_11600,N_11551);
nor U12424 (N_12424,N_11948,N_11622);
or U12425 (N_12425,N_11952,N_11599);
nand U12426 (N_12426,N_11852,N_11768);
or U12427 (N_12427,N_11814,N_11611);
and U12428 (N_12428,N_11771,N_11547);
xnor U12429 (N_12429,N_11840,N_11678);
nor U12430 (N_12430,N_11863,N_11604);
and U12431 (N_12431,N_11581,N_11514);
nor U12432 (N_12432,N_11941,N_11872);
nor U12433 (N_12433,N_11657,N_11896);
xnor U12434 (N_12434,N_11981,N_11709);
or U12435 (N_12435,N_11617,N_11972);
nor U12436 (N_12436,N_11543,N_11729);
nand U12437 (N_12437,N_11876,N_11598);
nand U12438 (N_12438,N_11542,N_11939);
nor U12439 (N_12439,N_11612,N_11696);
nor U12440 (N_12440,N_11513,N_11586);
and U12441 (N_12441,N_11939,N_11538);
xor U12442 (N_12442,N_11811,N_11990);
nand U12443 (N_12443,N_11586,N_11767);
or U12444 (N_12444,N_11879,N_11615);
nand U12445 (N_12445,N_11971,N_11735);
xor U12446 (N_12446,N_11572,N_11555);
or U12447 (N_12447,N_11944,N_11632);
and U12448 (N_12448,N_11963,N_11555);
nand U12449 (N_12449,N_11630,N_11576);
xnor U12450 (N_12450,N_11648,N_11684);
or U12451 (N_12451,N_11875,N_11526);
and U12452 (N_12452,N_11915,N_11508);
nor U12453 (N_12453,N_11687,N_11726);
or U12454 (N_12454,N_11781,N_11718);
nor U12455 (N_12455,N_11725,N_11504);
nand U12456 (N_12456,N_11616,N_11570);
nand U12457 (N_12457,N_11800,N_11951);
xor U12458 (N_12458,N_11977,N_11568);
nand U12459 (N_12459,N_11527,N_11613);
and U12460 (N_12460,N_11992,N_11645);
and U12461 (N_12461,N_11532,N_11759);
or U12462 (N_12462,N_11811,N_11552);
nand U12463 (N_12463,N_11580,N_11648);
nor U12464 (N_12464,N_11842,N_11699);
nand U12465 (N_12465,N_11502,N_11579);
and U12466 (N_12466,N_11767,N_11802);
xnor U12467 (N_12467,N_11785,N_11962);
nor U12468 (N_12468,N_11809,N_11802);
nor U12469 (N_12469,N_11975,N_11543);
nor U12470 (N_12470,N_11613,N_11560);
xnor U12471 (N_12471,N_11996,N_11532);
nor U12472 (N_12472,N_11765,N_11831);
and U12473 (N_12473,N_11832,N_11517);
or U12474 (N_12474,N_11698,N_11558);
and U12475 (N_12475,N_11696,N_11870);
nand U12476 (N_12476,N_11517,N_11712);
nor U12477 (N_12477,N_11990,N_11739);
or U12478 (N_12478,N_11680,N_11637);
nor U12479 (N_12479,N_11851,N_11518);
xnor U12480 (N_12480,N_11655,N_11982);
xor U12481 (N_12481,N_11818,N_11674);
and U12482 (N_12482,N_11694,N_11692);
nor U12483 (N_12483,N_11977,N_11959);
xor U12484 (N_12484,N_11658,N_11572);
or U12485 (N_12485,N_11649,N_11678);
or U12486 (N_12486,N_11860,N_11938);
nor U12487 (N_12487,N_11983,N_11834);
or U12488 (N_12488,N_11676,N_11858);
and U12489 (N_12489,N_11809,N_11507);
xor U12490 (N_12490,N_11694,N_11590);
nand U12491 (N_12491,N_11747,N_11689);
nor U12492 (N_12492,N_11674,N_11732);
or U12493 (N_12493,N_11949,N_11530);
nand U12494 (N_12494,N_11658,N_11541);
nor U12495 (N_12495,N_11518,N_11991);
or U12496 (N_12496,N_11931,N_11638);
nand U12497 (N_12497,N_11643,N_11858);
or U12498 (N_12498,N_11602,N_11507);
or U12499 (N_12499,N_11533,N_11654);
xor U12500 (N_12500,N_12468,N_12314);
nand U12501 (N_12501,N_12404,N_12021);
or U12502 (N_12502,N_12206,N_12480);
nor U12503 (N_12503,N_12348,N_12492);
xnor U12504 (N_12504,N_12462,N_12042);
nand U12505 (N_12505,N_12169,N_12176);
nand U12506 (N_12506,N_12472,N_12394);
xor U12507 (N_12507,N_12094,N_12450);
and U12508 (N_12508,N_12105,N_12174);
and U12509 (N_12509,N_12123,N_12217);
nor U12510 (N_12510,N_12451,N_12327);
or U12511 (N_12511,N_12034,N_12434);
nor U12512 (N_12512,N_12355,N_12049);
or U12513 (N_12513,N_12280,N_12099);
nor U12514 (N_12514,N_12183,N_12456);
nand U12515 (N_12515,N_12448,N_12320);
or U12516 (N_12516,N_12415,N_12358);
nand U12517 (N_12517,N_12454,N_12214);
and U12518 (N_12518,N_12211,N_12391);
xor U12519 (N_12519,N_12417,N_12184);
nor U12520 (N_12520,N_12427,N_12166);
and U12521 (N_12521,N_12283,N_12015);
xor U12522 (N_12522,N_12264,N_12317);
nand U12523 (N_12523,N_12298,N_12288);
xnor U12524 (N_12524,N_12428,N_12088);
and U12525 (N_12525,N_12224,N_12238);
nor U12526 (N_12526,N_12380,N_12086);
and U12527 (N_12527,N_12323,N_12261);
nor U12528 (N_12528,N_12340,N_12068);
xnor U12529 (N_12529,N_12381,N_12360);
or U12530 (N_12530,N_12148,N_12017);
and U12531 (N_12531,N_12396,N_12278);
nand U12532 (N_12532,N_12466,N_12220);
nand U12533 (N_12533,N_12406,N_12202);
and U12534 (N_12534,N_12098,N_12163);
or U12535 (N_12535,N_12442,N_12299);
nor U12536 (N_12536,N_12292,N_12044);
xnor U12537 (N_12537,N_12078,N_12012);
and U12538 (N_12538,N_12172,N_12002);
xor U12539 (N_12539,N_12197,N_12402);
nor U12540 (N_12540,N_12354,N_12065);
and U12541 (N_12541,N_12104,N_12305);
nor U12542 (N_12542,N_12365,N_12128);
nand U12543 (N_12543,N_12173,N_12095);
or U12544 (N_12544,N_12039,N_12331);
or U12545 (N_12545,N_12222,N_12393);
and U12546 (N_12546,N_12367,N_12204);
nand U12547 (N_12547,N_12066,N_12389);
nor U12548 (N_12548,N_12246,N_12435);
nand U12549 (N_12549,N_12338,N_12257);
nor U12550 (N_12550,N_12499,N_12439);
or U12551 (N_12551,N_12227,N_12410);
nand U12552 (N_12552,N_12158,N_12168);
nand U12553 (N_12553,N_12140,N_12014);
xor U12554 (N_12554,N_12420,N_12240);
and U12555 (N_12555,N_12187,N_12010);
xnor U12556 (N_12556,N_12141,N_12269);
or U12557 (N_12557,N_12271,N_12199);
or U12558 (N_12558,N_12255,N_12416);
and U12559 (N_12559,N_12074,N_12061);
nand U12560 (N_12560,N_12316,N_12216);
nor U12561 (N_12561,N_12397,N_12008);
nand U12562 (N_12562,N_12164,N_12481);
nor U12563 (N_12563,N_12102,N_12474);
and U12564 (N_12564,N_12242,N_12352);
or U12565 (N_12565,N_12342,N_12207);
and U12566 (N_12566,N_12115,N_12137);
or U12567 (N_12567,N_12073,N_12398);
and U12568 (N_12568,N_12134,N_12063);
nand U12569 (N_12569,N_12445,N_12009);
or U12570 (N_12570,N_12441,N_12362);
and U12571 (N_12571,N_12020,N_12223);
and U12572 (N_12572,N_12096,N_12013);
nor U12573 (N_12573,N_12248,N_12161);
nand U12574 (N_12574,N_12198,N_12000);
nand U12575 (N_12575,N_12275,N_12181);
or U12576 (N_12576,N_12180,N_12436);
xor U12577 (N_12577,N_12249,N_12325);
nand U12578 (N_12578,N_12090,N_12301);
or U12579 (N_12579,N_12465,N_12256);
nor U12580 (N_12580,N_12165,N_12023);
nor U12581 (N_12581,N_12471,N_12368);
nor U12582 (N_12582,N_12284,N_12219);
and U12583 (N_12583,N_12476,N_12313);
nand U12584 (N_12584,N_12228,N_12482);
nand U12585 (N_12585,N_12153,N_12453);
nand U12586 (N_12586,N_12421,N_12108);
nand U12587 (N_12587,N_12229,N_12159);
and U12588 (N_12588,N_12133,N_12233);
or U12589 (N_12589,N_12083,N_12405);
xor U12590 (N_12590,N_12241,N_12113);
and U12591 (N_12591,N_12029,N_12028);
nand U12592 (N_12592,N_12413,N_12375);
nor U12593 (N_12593,N_12129,N_12311);
and U12594 (N_12594,N_12024,N_12026);
nand U12595 (N_12595,N_12343,N_12419);
or U12596 (N_12596,N_12353,N_12359);
or U12597 (N_12597,N_12473,N_12139);
nand U12598 (N_12598,N_12218,N_12392);
or U12599 (N_12599,N_12213,N_12387);
and U12600 (N_12600,N_12265,N_12085);
nor U12601 (N_12601,N_12291,N_12370);
nand U12602 (N_12602,N_12205,N_12339);
nor U12603 (N_12603,N_12036,N_12443);
nand U12604 (N_12604,N_12127,N_12069);
and U12605 (N_12605,N_12433,N_12209);
xor U12606 (N_12606,N_12483,N_12383);
and U12607 (N_12607,N_12497,N_12003);
xnor U12608 (N_12608,N_12124,N_12236);
xor U12609 (N_12609,N_12109,N_12485);
nor U12610 (N_12610,N_12160,N_12239);
and U12611 (N_12611,N_12070,N_12270);
or U12612 (N_12612,N_12135,N_12328);
nor U12613 (N_12613,N_12189,N_12230);
nor U12614 (N_12614,N_12048,N_12486);
and U12615 (N_12615,N_12432,N_12458);
and U12616 (N_12616,N_12440,N_12136);
nand U12617 (N_12617,N_12156,N_12091);
nand U12618 (N_12618,N_12112,N_12491);
or U12619 (N_12619,N_12084,N_12245);
and U12620 (N_12620,N_12321,N_12379);
xor U12621 (N_12621,N_12201,N_12300);
or U12622 (N_12622,N_12175,N_12459);
nor U12623 (N_12623,N_12337,N_12011);
nor U12624 (N_12624,N_12424,N_12144);
nor U12625 (N_12625,N_12463,N_12267);
or U12626 (N_12626,N_12268,N_12312);
nor U12627 (N_12627,N_12341,N_12146);
or U12628 (N_12628,N_12422,N_12407);
nor U12629 (N_12629,N_12046,N_12281);
or U12630 (N_12630,N_12119,N_12460);
or U12631 (N_12631,N_12185,N_12263);
nor U12632 (N_12632,N_12058,N_12221);
or U12633 (N_12633,N_12496,N_12408);
nand U12634 (N_12634,N_12259,N_12147);
or U12635 (N_12635,N_12120,N_12452);
or U12636 (N_12636,N_12329,N_12056);
or U12637 (N_12637,N_12155,N_12005);
nand U12638 (N_12638,N_12082,N_12414);
or U12639 (N_12639,N_12194,N_12322);
nand U12640 (N_12640,N_12079,N_12423);
or U12641 (N_12641,N_12052,N_12431);
nand U12642 (N_12642,N_12346,N_12335);
nor U12643 (N_12643,N_12306,N_12045);
or U12644 (N_12644,N_12274,N_12131);
or U12645 (N_12645,N_12143,N_12234);
and U12646 (N_12646,N_12470,N_12032);
and U12647 (N_12647,N_12054,N_12333);
nand U12648 (N_12648,N_12294,N_12493);
nand U12649 (N_12649,N_12035,N_12072);
nor U12650 (N_12650,N_12179,N_12369);
or U12651 (N_12651,N_12336,N_12016);
and U12652 (N_12652,N_12019,N_12411);
or U12653 (N_12653,N_12494,N_12361);
and U12654 (N_12654,N_12177,N_12117);
xor U12655 (N_12655,N_12093,N_12097);
xor U12656 (N_12656,N_12378,N_12290);
nor U12657 (N_12657,N_12276,N_12412);
nor U12658 (N_12658,N_12043,N_12272);
nor U12659 (N_12659,N_12303,N_12089);
or U12660 (N_12660,N_12309,N_12430);
or U12661 (N_12661,N_12092,N_12488);
or U12662 (N_12662,N_12154,N_12372);
nand U12663 (N_12663,N_12193,N_12145);
nand U12664 (N_12664,N_12018,N_12081);
or U12665 (N_12665,N_12296,N_12373);
xnor U12666 (N_12666,N_12122,N_12118);
nand U12667 (N_12667,N_12385,N_12444);
or U12668 (N_12668,N_12364,N_12477);
xnor U12669 (N_12669,N_12231,N_12495);
xnor U12670 (N_12670,N_12399,N_12345);
nand U12671 (N_12671,N_12293,N_12196);
and U12672 (N_12672,N_12101,N_12064);
and U12673 (N_12673,N_12132,N_12210);
nand U12674 (N_12674,N_12006,N_12277);
nor U12675 (N_12675,N_12285,N_12304);
or U12676 (N_12676,N_12357,N_12076);
or U12677 (N_12677,N_12170,N_12171);
nor U12678 (N_12678,N_12429,N_12279);
xnor U12679 (N_12679,N_12350,N_12446);
xnor U12680 (N_12680,N_12190,N_12254);
xor U12681 (N_12681,N_12266,N_12212);
and U12682 (N_12682,N_12286,N_12038);
xor U12683 (N_12683,N_12426,N_12152);
nor U12684 (N_12684,N_12126,N_12116);
and U12685 (N_12685,N_12308,N_12386);
or U12686 (N_12686,N_12334,N_12403);
or U12687 (N_12687,N_12059,N_12363);
nand U12688 (N_12688,N_12037,N_12027);
xnor U12689 (N_12689,N_12282,N_12047);
and U12690 (N_12690,N_12077,N_12289);
and U12691 (N_12691,N_12247,N_12326);
or U12692 (N_12692,N_12244,N_12203);
and U12693 (N_12693,N_12178,N_12374);
or U12694 (N_12694,N_12191,N_12121);
xor U12695 (N_12695,N_12192,N_12400);
or U12696 (N_12696,N_12253,N_12041);
xnor U12697 (N_12697,N_12489,N_12457);
nor U12698 (N_12698,N_12251,N_12449);
nand U12699 (N_12699,N_12371,N_12087);
nor U12700 (N_12700,N_12273,N_12425);
and U12701 (N_12701,N_12467,N_12478);
xnor U12702 (N_12702,N_12200,N_12237);
nor U12703 (N_12703,N_12384,N_12100);
and U12704 (N_12704,N_12388,N_12111);
or U12705 (N_12705,N_12071,N_12366);
nand U12706 (N_12706,N_12031,N_12250);
nor U12707 (N_12707,N_12315,N_12344);
or U12708 (N_12708,N_12075,N_12001);
or U12709 (N_12709,N_12418,N_12258);
or U12710 (N_12710,N_12057,N_12347);
and U12711 (N_12711,N_12151,N_12060);
nand U12712 (N_12712,N_12150,N_12050);
nor U12713 (N_12713,N_12490,N_12007);
xor U12714 (N_12714,N_12208,N_12260);
and U12715 (N_12715,N_12356,N_12243);
nor U12716 (N_12716,N_12455,N_12464);
nand U12717 (N_12717,N_12390,N_12186);
or U12718 (N_12718,N_12142,N_12395);
nand U12719 (N_12719,N_12004,N_12226);
nor U12720 (N_12720,N_12461,N_12235);
and U12721 (N_12721,N_12484,N_12080);
or U12722 (N_12722,N_12324,N_12302);
or U12723 (N_12723,N_12103,N_12167);
or U12724 (N_12724,N_12157,N_12487);
xnor U12725 (N_12725,N_12188,N_12195);
nand U12726 (N_12726,N_12149,N_12040);
or U12727 (N_12727,N_12182,N_12215);
xor U12728 (N_12728,N_12138,N_12106);
and U12729 (N_12729,N_12025,N_12319);
or U12730 (N_12730,N_12107,N_12318);
or U12731 (N_12731,N_12162,N_12225);
and U12732 (N_12732,N_12401,N_12110);
and U12733 (N_12733,N_12232,N_12262);
and U12734 (N_12734,N_12051,N_12033);
xnor U12735 (N_12735,N_12022,N_12351);
nor U12736 (N_12736,N_12114,N_12332);
nor U12737 (N_12737,N_12030,N_12062);
nand U12738 (N_12738,N_12295,N_12252);
nand U12739 (N_12739,N_12055,N_12067);
nand U12740 (N_12740,N_12125,N_12447);
or U12741 (N_12741,N_12437,N_12310);
nor U12742 (N_12742,N_12377,N_12475);
and U12743 (N_12743,N_12479,N_12349);
nand U12744 (N_12744,N_12469,N_12376);
xnor U12745 (N_12745,N_12297,N_12053);
nand U12746 (N_12746,N_12438,N_12307);
nand U12747 (N_12747,N_12409,N_12130);
and U12748 (N_12748,N_12330,N_12498);
and U12749 (N_12749,N_12382,N_12287);
nand U12750 (N_12750,N_12055,N_12295);
or U12751 (N_12751,N_12420,N_12418);
xnor U12752 (N_12752,N_12428,N_12252);
or U12753 (N_12753,N_12329,N_12352);
and U12754 (N_12754,N_12173,N_12172);
or U12755 (N_12755,N_12388,N_12278);
xnor U12756 (N_12756,N_12427,N_12460);
or U12757 (N_12757,N_12448,N_12070);
nand U12758 (N_12758,N_12363,N_12356);
or U12759 (N_12759,N_12310,N_12290);
nor U12760 (N_12760,N_12326,N_12036);
or U12761 (N_12761,N_12292,N_12146);
nand U12762 (N_12762,N_12084,N_12324);
and U12763 (N_12763,N_12471,N_12011);
xnor U12764 (N_12764,N_12212,N_12431);
xor U12765 (N_12765,N_12385,N_12441);
and U12766 (N_12766,N_12332,N_12450);
and U12767 (N_12767,N_12461,N_12030);
nand U12768 (N_12768,N_12183,N_12443);
nor U12769 (N_12769,N_12167,N_12019);
and U12770 (N_12770,N_12290,N_12139);
nand U12771 (N_12771,N_12056,N_12453);
nand U12772 (N_12772,N_12379,N_12103);
nor U12773 (N_12773,N_12304,N_12422);
nor U12774 (N_12774,N_12001,N_12077);
nor U12775 (N_12775,N_12100,N_12424);
and U12776 (N_12776,N_12481,N_12052);
nor U12777 (N_12777,N_12173,N_12276);
nand U12778 (N_12778,N_12429,N_12233);
or U12779 (N_12779,N_12498,N_12255);
xor U12780 (N_12780,N_12392,N_12348);
or U12781 (N_12781,N_12284,N_12427);
and U12782 (N_12782,N_12235,N_12484);
and U12783 (N_12783,N_12427,N_12403);
nor U12784 (N_12784,N_12166,N_12403);
and U12785 (N_12785,N_12194,N_12242);
nand U12786 (N_12786,N_12232,N_12213);
nor U12787 (N_12787,N_12220,N_12373);
and U12788 (N_12788,N_12269,N_12220);
nor U12789 (N_12789,N_12247,N_12439);
or U12790 (N_12790,N_12408,N_12106);
nor U12791 (N_12791,N_12409,N_12162);
xnor U12792 (N_12792,N_12174,N_12339);
or U12793 (N_12793,N_12073,N_12057);
nor U12794 (N_12794,N_12471,N_12071);
xor U12795 (N_12795,N_12100,N_12082);
or U12796 (N_12796,N_12442,N_12334);
nor U12797 (N_12797,N_12372,N_12062);
nand U12798 (N_12798,N_12417,N_12497);
nand U12799 (N_12799,N_12476,N_12135);
xor U12800 (N_12800,N_12366,N_12181);
or U12801 (N_12801,N_12137,N_12314);
nand U12802 (N_12802,N_12266,N_12415);
or U12803 (N_12803,N_12061,N_12425);
and U12804 (N_12804,N_12384,N_12475);
and U12805 (N_12805,N_12074,N_12332);
nand U12806 (N_12806,N_12250,N_12025);
nand U12807 (N_12807,N_12206,N_12039);
or U12808 (N_12808,N_12338,N_12445);
xor U12809 (N_12809,N_12307,N_12309);
nor U12810 (N_12810,N_12153,N_12242);
xor U12811 (N_12811,N_12436,N_12245);
nor U12812 (N_12812,N_12389,N_12019);
xor U12813 (N_12813,N_12391,N_12006);
xor U12814 (N_12814,N_12010,N_12391);
or U12815 (N_12815,N_12491,N_12080);
and U12816 (N_12816,N_12174,N_12496);
and U12817 (N_12817,N_12316,N_12094);
and U12818 (N_12818,N_12332,N_12466);
or U12819 (N_12819,N_12434,N_12129);
nand U12820 (N_12820,N_12164,N_12361);
nand U12821 (N_12821,N_12046,N_12412);
or U12822 (N_12822,N_12256,N_12401);
nor U12823 (N_12823,N_12127,N_12032);
or U12824 (N_12824,N_12390,N_12350);
nor U12825 (N_12825,N_12181,N_12049);
nor U12826 (N_12826,N_12155,N_12052);
and U12827 (N_12827,N_12001,N_12264);
nor U12828 (N_12828,N_12086,N_12486);
or U12829 (N_12829,N_12273,N_12193);
xnor U12830 (N_12830,N_12120,N_12302);
xnor U12831 (N_12831,N_12195,N_12458);
or U12832 (N_12832,N_12383,N_12079);
or U12833 (N_12833,N_12340,N_12434);
xnor U12834 (N_12834,N_12198,N_12286);
and U12835 (N_12835,N_12094,N_12091);
xor U12836 (N_12836,N_12261,N_12193);
and U12837 (N_12837,N_12373,N_12309);
nand U12838 (N_12838,N_12307,N_12005);
and U12839 (N_12839,N_12334,N_12007);
xnor U12840 (N_12840,N_12227,N_12231);
nor U12841 (N_12841,N_12030,N_12452);
nand U12842 (N_12842,N_12496,N_12454);
nor U12843 (N_12843,N_12076,N_12061);
nor U12844 (N_12844,N_12158,N_12365);
or U12845 (N_12845,N_12239,N_12403);
or U12846 (N_12846,N_12101,N_12211);
nor U12847 (N_12847,N_12171,N_12053);
or U12848 (N_12848,N_12321,N_12160);
and U12849 (N_12849,N_12369,N_12217);
and U12850 (N_12850,N_12289,N_12165);
nor U12851 (N_12851,N_12333,N_12111);
and U12852 (N_12852,N_12357,N_12483);
xnor U12853 (N_12853,N_12391,N_12245);
xnor U12854 (N_12854,N_12170,N_12016);
nand U12855 (N_12855,N_12143,N_12317);
nor U12856 (N_12856,N_12443,N_12499);
nand U12857 (N_12857,N_12234,N_12400);
or U12858 (N_12858,N_12166,N_12153);
nor U12859 (N_12859,N_12491,N_12301);
or U12860 (N_12860,N_12346,N_12247);
xor U12861 (N_12861,N_12324,N_12135);
and U12862 (N_12862,N_12306,N_12268);
nor U12863 (N_12863,N_12378,N_12174);
or U12864 (N_12864,N_12064,N_12171);
nor U12865 (N_12865,N_12296,N_12197);
nand U12866 (N_12866,N_12168,N_12237);
nor U12867 (N_12867,N_12076,N_12100);
xor U12868 (N_12868,N_12192,N_12166);
nor U12869 (N_12869,N_12129,N_12112);
nor U12870 (N_12870,N_12295,N_12250);
nand U12871 (N_12871,N_12214,N_12156);
xor U12872 (N_12872,N_12137,N_12291);
nand U12873 (N_12873,N_12068,N_12426);
xnor U12874 (N_12874,N_12332,N_12083);
or U12875 (N_12875,N_12203,N_12263);
xor U12876 (N_12876,N_12124,N_12129);
xor U12877 (N_12877,N_12002,N_12420);
and U12878 (N_12878,N_12111,N_12183);
nand U12879 (N_12879,N_12144,N_12150);
nor U12880 (N_12880,N_12139,N_12384);
and U12881 (N_12881,N_12006,N_12176);
xor U12882 (N_12882,N_12305,N_12145);
and U12883 (N_12883,N_12375,N_12383);
and U12884 (N_12884,N_12042,N_12378);
and U12885 (N_12885,N_12201,N_12237);
and U12886 (N_12886,N_12401,N_12136);
nor U12887 (N_12887,N_12191,N_12232);
nand U12888 (N_12888,N_12014,N_12358);
xnor U12889 (N_12889,N_12170,N_12002);
xnor U12890 (N_12890,N_12301,N_12039);
or U12891 (N_12891,N_12432,N_12368);
xor U12892 (N_12892,N_12085,N_12430);
and U12893 (N_12893,N_12086,N_12217);
xnor U12894 (N_12894,N_12347,N_12126);
nor U12895 (N_12895,N_12122,N_12116);
or U12896 (N_12896,N_12408,N_12340);
and U12897 (N_12897,N_12155,N_12338);
and U12898 (N_12898,N_12092,N_12322);
nand U12899 (N_12899,N_12339,N_12269);
nand U12900 (N_12900,N_12316,N_12418);
and U12901 (N_12901,N_12095,N_12073);
and U12902 (N_12902,N_12348,N_12127);
or U12903 (N_12903,N_12468,N_12111);
xnor U12904 (N_12904,N_12190,N_12185);
nor U12905 (N_12905,N_12162,N_12304);
xor U12906 (N_12906,N_12072,N_12048);
xnor U12907 (N_12907,N_12482,N_12057);
nand U12908 (N_12908,N_12216,N_12254);
nor U12909 (N_12909,N_12407,N_12433);
nand U12910 (N_12910,N_12038,N_12252);
or U12911 (N_12911,N_12133,N_12286);
nor U12912 (N_12912,N_12243,N_12083);
nor U12913 (N_12913,N_12046,N_12469);
and U12914 (N_12914,N_12071,N_12430);
or U12915 (N_12915,N_12183,N_12474);
xor U12916 (N_12916,N_12027,N_12036);
xnor U12917 (N_12917,N_12290,N_12208);
and U12918 (N_12918,N_12387,N_12431);
and U12919 (N_12919,N_12085,N_12465);
nand U12920 (N_12920,N_12069,N_12481);
and U12921 (N_12921,N_12424,N_12050);
nand U12922 (N_12922,N_12265,N_12172);
xor U12923 (N_12923,N_12205,N_12254);
nand U12924 (N_12924,N_12443,N_12402);
nor U12925 (N_12925,N_12328,N_12118);
xor U12926 (N_12926,N_12196,N_12045);
or U12927 (N_12927,N_12257,N_12169);
and U12928 (N_12928,N_12354,N_12010);
xor U12929 (N_12929,N_12153,N_12193);
or U12930 (N_12930,N_12106,N_12411);
and U12931 (N_12931,N_12078,N_12479);
or U12932 (N_12932,N_12386,N_12150);
or U12933 (N_12933,N_12094,N_12048);
nor U12934 (N_12934,N_12187,N_12445);
and U12935 (N_12935,N_12095,N_12367);
and U12936 (N_12936,N_12026,N_12125);
xor U12937 (N_12937,N_12105,N_12068);
nor U12938 (N_12938,N_12465,N_12106);
and U12939 (N_12939,N_12116,N_12164);
or U12940 (N_12940,N_12078,N_12357);
and U12941 (N_12941,N_12280,N_12489);
nor U12942 (N_12942,N_12361,N_12316);
nor U12943 (N_12943,N_12224,N_12492);
xnor U12944 (N_12944,N_12029,N_12264);
or U12945 (N_12945,N_12005,N_12418);
xnor U12946 (N_12946,N_12041,N_12368);
nor U12947 (N_12947,N_12338,N_12478);
xor U12948 (N_12948,N_12384,N_12424);
and U12949 (N_12949,N_12446,N_12196);
xor U12950 (N_12950,N_12389,N_12381);
nand U12951 (N_12951,N_12343,N_12003);
and U12952 (N_12952,N_12181,N_12307);
nand U12953 (N_12953,N_12164,N_12268);
xor U12954 (N_12954,N_12179,N_12159);
nor U12955 (N_12955,N_12098,N_12006);
nand U12956 (N_12956,N_12391,N_12436);
nor U12957 (N_12957,N_12390,N_12319);
or U12958 (N_12958,N_12051,N_12473);
nand U12959 (N_12959,N_12272,N_12438);
xnor U12960 (N_12960,N_12447,N_12463);
xor U12961 (N_12961,N_12067,N_12046);
or U12962 (N_12962,N_12269,N_12379);
or U12963 (N_12963,N_12249,N_12417);
nor U12964 (N_12964,N_12284,N_12178);
nand U12965 (N_12965,N_12345,N_12045);
and U12966 (N_12966,N_12120,N_12242);
nor U12967 (N_12967,N_12428,N_12345);
xor U12968 (N_12968,N_12295,N_12289);
and U12969 (N_12969,N_12314,N_12246);
nor U12970 (N_12970,N_12233,N_12187);
xnor U12971 (N_12971,N_12453,N_12148);
and U12972 (N_12972,N_12014,N_12357);
nand U12973 (N_12973,N_12061,N_12001);
xnor U12974 (N_12974,N_12016,N_12246);
xnor U12975 (N_12975,N_12026,N_12113);
nor U12976 (N_12976,N_12244,N_12103);
nor U12977 (N_12977,N_12313,N_12049);
or U12978 (N_12978,N_12235,N_12266);
or U12979 (N_12979,N_12460,N_12324);
and U12980 (N_12980,N_12014,N_12336);
and U12981 (N_12981,N_12136,N_12190);
nor U12982 (N_12982,N_12329,N_12408);
and U12983 (N_12983,N_12309,N_12489);
xor U12984 (N_12984,N_12047,N_12127);
or U12985 (N_12985,N_12478,N_12140);
nor U12986 (N_12986,N_12384,N_12226);
and U12987 (N_12987,N_12341,N_12058);
nor U12988 (N_12988,N_12005,N_12450);
and U12989 (N_12989,N_12076,N_12145);
nor U12990 (N_12990,N_12346,N_12343);
and U12991 (N_12991,N_12141,N_12122);
nor U12992 (N_12992,N_12208,N_12241);
or U12993 (N_12993,N_12056,N_12177);
nand U12994 (N_12994,N_12167,N_12282);
xnor U12995 (N_12995,N_12112,N_12418);
nand U12996 (N_12996,N_12240,N_12371);
xor U12997 (N_12997,N_12379,N_12335);
and U12998 (N_12998,N_12390,N_12496);
xnor U12999 (N_12999,N_12467,N_12055);
nand U13000 (N_13000,N_12874,N_12611);
nor U13001 (N_13001,N_12884,N_12873);
nand U13002 (N_13002,N_12737,N_12607);
nand U13003 (N_13003,N_12672,N_12775);
and U13004 (N_13004,N_12533,N_12590);
or U13005 (N_13005,N_12870,N_12599);
xnor U13006 (N_13006,N_12595,N_12524);
xor U13007 (N_13007,N_12633,N_12805);
nor U13008 (N_13008,N_12876,N_12732);
nor U13009 (N_13009,N_12634,N_12703);
and U13010 (N_13010,N_12937,N_12632);
and U13011 (N_13011,N_12807,N_12908);
nor U13012 (N_13012,N_12577,N_12548);
nand U13013 (N_13013,N_12646,N_12973);
and U13014 (N_13014,N_12912,N_12994);
xor U13015 (N_13015,N_12858,N_12628);
or U13016 (N_13016,N_12835,N_12917);
xnor U13017 (N_13017,N_12772,N_12883);
nand U13018 (N_13018,N_12934,N_12783);
xnor U13019 (N_13019,N_12663,N_12981);
nand U13020 (N_13020,N_12790,N_12527);
or U13021 (N_13021,N_12508,N_12654);
nand U13022 (N_13022,N_12955,N_12553);
xnor U13023 (N_13023,N_12601,N_12780);
nor U13024 (N_13024,N_12963,N_12603);
nand U13025 (N_13025,N_12920,N_12926);
nor U13026 (N_13026,N_12704,N_12869);
nand U13027 (N_13027,N_12614,N_12759);
or U13028 (N_13028,N_12636,N_12593);
or U13029 (N_13029,N_12960,N_12733);
xnor U13030 (N_13030,N_12850,N_12653);
nor U13031 (N_13031,N_12962,N_12546);
xnor U13032 (N_13032,N_12512,N_12640);
xor U13033 (N_13033,N_12610,N_12896);
nor U13034 (N_13034,N_12735,N_12801);
and U13035 (N_13035,N_12972,N_12958);
xnor U13036 (N_13036,N_12530,N_12575);
nor U13037 (N_13037,N_12868,N_12929);
nand U13038 (N_13038,N_12826,N_12815);
nand U13039 (N_13039,N_12657,N_12539);
nor U13040 (N_13040,N_12674,N_12901);
xor U13041 (N_13041,N_12856,N_12931);
or U13042 (N_13042,N_12616,N_12596);
xor U13043 (N_13043,N_12866,N_12648);
nand U13044 (N_13044,N_12836,N_12786);
nand U13045 (N_13045,N_12589,N_12720);
or U13046 (N_13046,N_12693,N_12797);
nand U13047 (N_13047,N_12859,N_12882);
and U13048 (N_13048,N_12989,N_12935);
and U13049 (N_13049,N_12681,N_12839);
nand U13050 (N_13050,N_12840,N_12777);
xnor U13051 (N_13051,N_12586,N_12846);
nor U13052 (N_13052,N_12705,N_12682);
nand U13053 (N_13053,N_12650,N_12619);
xnor U13054 (N_13054,N_12608,N_12739);
and U13055 (N_13055,N_12965,N_12665);
nand U13056 (N_13056,N_12924,N_12905);
xor U13057 (N_13057,N_12979,N_12565);
or U13058 (N_13058,N_12558,N_12879);
or U13059 (N_13059,N_12848,N_12789);
nor U13060 (N_13060,N_12925,N_12729);
xor U13061 (N_13061,N_12605,N_12860);
nand U13062 (N_13062,N_12769,N_12932);
nor U13063 (N_13063,N_12871,N_12550);
and U13064 (N_13064,N_12571,N_12515);
nor U13065 (N_13065,N_12742,N_12773);
nand U13066 (N_13066,N_12712,N_12738);
or U13067 (N_13067,N_12624,N_12606);
xnor U13068 (N_13068,N_12647,N_12660);
and U13069 (N_13069,N_12950,N_12594);
nor U13070 (N_13070,N_12516,N_12952);
or U13071 (N_13071,N_12756,N_12602);
nor U13072 (N_13072,N_12991,N_12584);
nand U13073 (N_13073,N_12655,N_12670);
and U13074 (N_13074,N_12652,N_12863);
and U13075 (N_13075,N_12538,N_12851);
nor U13076 (N_13076,N_12552,N_12699);
nand U13077 (N_13077,N_12872,N_12715);
nand U13078 (N_13078,N_12765,N_12881);
nor U13079 (N_13079,N_12502,N_12617);
and U13080 (N_13080,N_12734,N_12942);
nand U13081 (N_13081,N_12829,N_12580);
nand U13082 (N_13082,N_12814,N_12597);
nor U13083 (N_13083,N_12921,N_12907);
and U13084 (N_13084,N_12673,N_12878);
xnor U13085 (N_13085,N_12534,N_12697);
and U13086 (N_13086,N_12642,N_12669);
and U13087 (N_13087,N_12744,N_12659);
xor U13088 (N_13088,N_12853,N_12988);
or U13089 (N_13089,N_12944,N_12880);
nand U13090 (N_13090,N_12827,N_12845);
nand U13091 (N_13091,N_12658,N_12549);
xor U13092 (N_13092,N_12844,N_12510);
or U13093 (N_13093,N_12837,N_12638);
nor U13094 (N_13094,N_12518,N_12700);
and U13095 (N_13095,N_12841,N_12581);
nand U13096 (N_13096,N_12587,N_12536);
nor U13097 (N_13097,N_12644,N_12849);
xor U13098 (N_13098,N_12909,N_12519);
nand U13099 (N_13099,N_12762,N_12875);
and U13100 (N_13100,N_12526,N_12641);
nand U13101 (N_13101,N_12517,N_12834);
nand U13102 (N_13102,N_12854,N_12645);
xor U13103 (N_13103,N_12522,N_12977);
or U13104 (N_13104,N_12885,N_12656);
or U13105 (N_13105,N_12600,N_12592);
or U13106 (N_13106,N_12781,N_12941);
nor U13107 (N_13107,N_12877,N_12887);
or U13108 (N_13108,N_12598,N_12916);
or U13109 (N_13109,N_12511,N_12588);
nor U13110 (N_13110,N_12802,N_12643);
nand U13111 (N_13111,N_12545,N_12778);
nor U13112 (N_13112,N_12514,N_12821);
nand U13113 (N_13113,N_12551,N_12583);
nand U13114 (N_13114,N_12813,N_12639);
and U13115 (N_13115,N_12831,N_12900);
nor U13116 (N_13116,N_12864,N_12919);
nand U13117 (N_13117,N_12531,N_12749);
xor U13118 (N_13118,N_12637,N_12609);
nor U13119 (N_13119,N_12707,N_12776);
or U13120 (N_13120,N_12902,N_12579);
or U13121 (N_13121,N_12661,N_12787);
or U13122 (N_13122,N_12562,N_12892);
nor U13123 (N_13123,N_12984,N_12573);
or U13124 (N_13124,N_12582,N_12623);
and U13125 (N_13125,N_12626,N_12535);
nand U13126 (N_13126,N_12555,N_12822);
or U13127 (N_13127,N_12891,N_12560);
xnor U13128 (N_13128,N_12709,N_12564);
nor U13129 (N_13129,N_12622,N_12847);
or U13130 (N_13130,N_12529,N_12940);
and U13131 (N_13131,N_12970,N_12615);
nand U13132 (N_13132,N_12855,N_12572);
xor U13133 (N_13133,N_12691,N_12726);
xor U13134 (N_13134,N_12898,N_12559);
and U13135 (N_13135,N_12861,N_12629);
nand U13136 (N_13136,N_12793,N_12904);
xor U13137 (N_13137,N_12723,N_12746);
nand U13138 (N_13138,N_12993,N_12507);
and U13139 (N_13139,N_12743,N_12753);
nor U13140 (N_13140,N_12927,N_12692);
and U13141 (N_13141,N_12574,N_12711);
xnor U13142 (N_13142,N_12544,N_12968);
nor U13143 (N_13143,N_12649,N_12812);
and U13144 (N_13144,N_12701,N_12949);
xor U13145 (N_13145,N_12690,N_12625);
nor U13146 (N_13146,N_12911,N_12717);
or U13147 (N_13147,N_12757,N_12532);
nand U13148 (N_13148,N_12718,N_12567);
or U13149 (N_13149,N_12767,N_12666);
and U13150 (N_13150,N_12967,N_12750);
nand U13151 (N_13151,N_12591,N_12945);
and U13152 (N_13152,N_12684,N_12943);
and U13153 (N_13153,N_12721,N_12930);
xor U13154 (N_13154,N_12928,N_12696);
or U13155 (N_13155,N_12999,N_12992);
nor U13156 (N_13156,N_12631,N_12811);
or U13157 (N_13157,N_12852,N_12630);
or U13158 (N_13158,N_12897,N_12953);
or U13159 (N_13159,N_12740,N_12620);
or U13160 (N_13160,N_12543,N_12865);
or U13161 (N_13161,N_12923,N_12635);
or U13162 (N_13162,N_12763,N_12713);
nor U13163 (N_13163,N_12770,N_12667);
xor U13164 (N_13164,N_12751,N_12677);
or U13165 (N_13165,N_12830,N_12889);
xnor U13166 (N_13166,N_12585,N_12725);
and U13167 (N_13167,N_12843,N_12817);
or U13168 (N_13168,N_12758,N_12987);
xor U13169 (N_13169,N_12795,N_12810);
and U13170 (N_13170,N_12986,N_12969);
nand U13171 (N_13171,N_12695,N_12966);
and U13172 (N_13172,N_12689,N_12686);
nor U13173 (N_13173,N_12706,N_12819);
nor U13174 (N_13174,N_12521,N_12974);
nand U13175 (N_13175,N_12996,N_12708);
and U13176 (N_13176,N_12867,N_12651);
or U13177 (N_13177,N_12833,N_12857);
and U13178 (N_13178,N_12792,N_12785);
or U13179 (N_13179,N_12683,N_12959);
xor U13180 (N_13180,N_12520,N_12687);
or U13181 (N_13181,N_12752,N_12886);
xnor U13182 (N_13182,N_12724,N_12755);
nand U13183 (N_13183,N_12728,N_12675);
or U13184 (N_13184,N_12782,N_12668);
and U13185 (N_13185,N_12557,N_12760);
and U13186 (N_13186,N_12664,N_12731);
and U13187 (N_13187,N_12980,N_12745);
or U13188 (N_13188,N_12922,N_12771);
or U13189 (N_13189,N_12806,N_12754);
or U13190 (N_13190,N_12774,N_12766);
and U13191 (N_13191,N_12768,N_12824);
nor U13192 (N_13192,N_12621,N_12976);
and U13193 (N_13193,N_12803,N_12933);
xor U13194 (N_13194,N_12505,N_12915);
or U13195 (N_13195,N_12890,N_12948);
nor U13196 (N_13196,N_12722,N_12820);
nand U13197 (N_13197,N_12685,N_12501);
nand U13198 (N_13198,N_12716,N_12936);
nand U13199 (N_13199,N_12513,N_12995);
or U13200 (N_13200,N_12804,N_12888);
or U13201 (N_13201,N_12719,N_12540);
nor U13202 (N_13202,N_12500,N_12828);
nand U13203 (N_13203,N_12971,N_12561);
nor U13204 (N_13204,N_12893,N_12694);
nand U13205 (N_13205,N_12947,N_12823);
xor U13206 (N_13206,N_12627,N_12764);
nor U13207 (N_13207,N_12906,N_12523);
nor U13208 (N_13208,N_12914,N_12506);
or U13209 (N_13209,N_12799,N_12983);
nand U13210 (N_13210,N_12570,N_12800);
or U13211 (N_13211,N_12556,N_12702);
xnor U13212 (N_13212,N_12714,N_12997);
and U13213 (N_13213,N_12794,N_12961);
or U13214 (N_13214,N_12939,N_12680);
nand U13215 (N_13215,N_12748,N_12618);
nand U13216 (N_13216,N_12964,N_12832);
and U13217 (N_13217,N_12862,N_12796);
or U13218 (N_13218,N_12537,N_12761);
xnor U13219 (N_13219,N_12842,N_12678);
xor U13220 (N_13220,N_12985,N_12688);
or U13221 (N_13221,N_12982,N_12747);
xnor U13222 (N_13222,N_12569,N_12808);
or U13223 (N_13223,N_12791,N_12809);
nand U13224 (N_13224,N_12838,N_12698);
nand U13225 (N_13225,N_12727,N_12509);
or U13226 (N_13226,N_12613,N_12525);
and U13227 (N_13227,N_12563,N_12676);
nand U13228 (N_13228,N_12504,N_12566);
nand U13229 (N_13229,N_12741,N_12503);
xnor U13230 (N_13230,N_12576,N_12541);
or U13231 (N_13231,N_12779,N_12918);
xnor U13232 (N_13232,N_12604,N_12825);
nor U13233 (N_13233,N_12730,N_12679);
or U13234 (N_13234,N_12956,N_12894);
or U13235 (N_13235,N_12612,N_12736);
nor U13236 (N_13236,N_12903,N_12816);
nand U13237 (N_13237,N_12990,N_12938);
or U13238 (N_13238,N_12975,N_12954);
or U13239 (N_13239,N_12710,N_12662);
xnor U13240 (N_13240,N_12899,N_12946);
nand U13241 (N_13241,N_12913,N_12568);
or U13242 (N_13242,N_12788,N_12542);
xnor U13243 (N_13243,N_12951,N_12910);
nand U13244 (N_13244,N_12784,N_12554);
or U13245 (N_13245,N_12957,N_12671);
nand U13246 (N_13246,N_12998,N_12578);
xor U13247 (N_13247,N_12528,N_12895);
nand U13248 (N_13248,N_12818,N_12547);
and U13249 (N_13249,N_12798,N_12978);
and U13250 (N_13250,N_12853,N_12944);
and U13251 (N_13251,N_12993,N_12786);
nand U13252 (N_13252,N_12734,N_12627);
xor U13253 (N_13253,N_12532,N_12558);
and U13254 (N_13254,N_12502,N_12546);
and U13255 (N_13255,N_12806,N_12838);
xor U13256 (N_13256,N_12993,N_12760);
or U13257 (N_13257,N_12690,N_12723);
and U13258 (N_13258,N_12975,N_12681);
xor U13259 (N_13259,N_12945,N_12967);
and U13260 (N_13260,N_12562,N_12547);
and U13261 (N_13261,N_12704,N_12985);
nand U13262 (N_13262,N_12594,N_12858);
or U13263 (N_13263,N_12746,N_12554);
nor U13264 (N_13264,N_12597,N_12896);
nand U13265 (N_13265,N_12537,N_12721);
or U13266 (N_13266,N_12637,N_12874);
nor U13267 (N_13267,N_12722,N_12603);
or U13268 (N_13268,N_12519,N_12819);
or U13269 (N_13269,N_12798,N_12647);
xor U13270 (N_13270,N_12880,N_12896);
nand U13271 (N_13271,N_12867,N_12703);
nand U13272 (N_13272,N_12805,N_12759);
or U13273 (N_13273,N_12945,N_12803);
nor U13274 (N_13274,N_12572,N_12644);
nor U13275 (N_13275,N_12667,N_12779);
and U13276 (N_13276,N_12533,N_12904);
nor U13277 (N_13277,N_12739,N_12899);
nand U13278 (N_13278,N_12707,N_12858);
and U13279 (N_13279,N_12873,N_12703);
nand U13280 (N_13280,N_12733,N_12626);
xor U13281 (N_13281,N_12599,N_12834);
and U13282 (N_13282,N_12699,N_12713);
or U13283 (N_13283,N_12910,N_12702);
nor U13284 (N_13284,N_12682,N_12530);
xnor U13285 (N_13285,N_12843,N_12925);
xnor U13286 (N_13286,N_12756,N_12743);
or U13287 (N_13287,N_12829,N_12645);
or U13288 (N_13288,N_12594,N_12815);
nand U13289 (N_13289,N_12534,N_12783);
nand U13290 (N_13290,N_12733,N_12630);
xor U13291 (N_13291,N_12790,N_12540);
or U13292 (N_13292,N_12534,N_12905);
nand U13293 (N_13293,N_12551,N_12714);
and U13294 (N_13294,N_12948,N_12901);
or U13295 (N_13295,N_12790,N_12998);
xor U13296 (N_13296,N_12756,N_12671);
nor U13297 (N_13297,N_12886,N_12616);
nor U13298 (N_13298,N_12544,N_12599);
nor U13299 (N_13299,N_12820,N_12558);
xor U13300 (N_13300,N_12958,N_12973);
xnor U13301 (N_13301,N_12913,N_12952);
nand U13302 (N_13302,N_12623,N_12521);
nand U13303 (N_13303,N_12928,N_12689);
and U13304 (N_13304,N_12751,N_12769);
and U13305 (N_13305,N_12561,N_12552);
nand U13306 (N_13306,N_12566,N_12849);
nand U13307 (N_13307,N_12941,N_12835);
nand U13308 (N_13308,N_12531,N_12756);
nand U13309 (N_13309,N_12888,N_12836);
nor U13310 (N_13310,N_12690,N_12630);
or U13311 (N_13311,N_12549,N_12518);
nand U13312 (N_13312,N_12624,N_12792);
or U13313 (N_13313,N_12553,N_12767);
and U13314 (N_13314,N_12982,N_12557);
nand U13315 (N_13315,N_12521,N_12629);
and U13316 (N_13316,N_12587,N_12543);
nor U13317 (N_13317,N_12735,N_12517);
or U13318 (N_13318,N_12837,N_12785);
nor U13319 (N_13319,N_12743,N_12724);
and U13320 (N_13320,N_12757,N_12746);
and U13321 (N_13321,N_12836,N_12821);
or U13322 (N_13322,N_12782,N_12968);
or U13323 (N_13323,N_12844,N_12531);
and U13324 (N_13324,N_12575,N_12742);
or U13325 (N_13325,N_12929,N_12662);
xor U13326 (N_13326,N_12770,N_12624);
nand U13327 (N_13327,N_12818,N_12868);
or U13328 (N_13328,N_12920,N_12973);
or U13329 (N_13329,N_12712,N_12642);
nor U13330 (N_13330,N_12729,N_12555);
xnor U13331 (N_13331,N_12557,N_12637);
nor U13332 (N_13332,N_12904,N_12937);
or U13333 (N_13333,N_12845,N_12516);
and U13334 (N_13334,N_12724,N_12578);
or U13335 (N_13335,N_12855,N_12763);
xor U13336 (N_13336,N_12834,N_12657);
and U13337 (N_13337,N_12985,N_12696);
or U13338 (N_13338,N_12964,N_12903);
nor U13339 (N_13339,N_12551,N_12565);
or U13340 (N_13340,N_12662,N_12604);
nor U13341 (N_13341,N_12793,N_12778);
nand U13342 (N_13342,N_12829,N_12883);
nand U13343 (N_13343,N_12825,N_12612);
or U13344 (N_13344,N_12788,N_12648);
or U13345 (N_13345,N_12692,N_12559);
xor U13346 (N_13346,N_12512,N_12696);
nor U13347 (N_13347,N_12957,N_12658);
or U13348 (N_13348,N_12560,N_12818);
xnor U13349 (N_13349,N_12517,N_12564);
nand U13350 (N_13350,N_12650,N_12823);
xor U13351 (N_13351,N_12527,N_12504);
or U13352 (N_13352,N_12959,N_12824);
nand U13353 (N_13353,N_12981,N_12887);
xnor U13354 (N_13354,N_12708,N_12690);
nand U13355 (N_13355,N_12974,N_12626);
nand U13356 (N_13356,N_12586,N_12572);
nor U13357 (N_13357,N_12649,N_12826);
or U13358 (N_13358,N_12670,N_12628);
xor U13359 (N_13359,N_12809,N_12613);
and U13360 (N_13360,N_12910,N_12986);
or U13361 (N_13361,N_12702,N_12784);
or U13362 (N_13362,N_12798,N_12893);
nand U13363 (N_13363,N_12835,N_12925);
nor U13364 (N_13364,N_12757,N_12881);
or U13365 (N_13365,N_12926,N_12553);
nor U13366 (N_13366,N_12837,N_12812);
nand U13367 (N_13367,N_12699,N_12821);
nand U13368 (N_13368,N_12866,N_12548);
xnor U13369 (N_13369,N_12932,N_12875);
or U13370 (N_13370,N_12650,N_12675);
nor U13371 (N_13371,N_12744,N_12949);
nor U13372 (N_13372,N_12880,N_12860);
nor U13373 (N_13373,N_12767,N_12606);
nor U13374 (N_13374,N_12714,N_12926);
nand U13375 (N_13375,N_12846,N_12738);
nor U13376 (N_13376,N_12819,N_12978);
xnor U13377 (N_13377,N_12562,N_12723);
and U13378 (N_13378,N_12515,N_12757);
and U13379 (N_13379,N_12858,N_12643);
nand U13380 (N_13380,N_12872,N_12707);
xnor U13381 (N_13381,N_12799,N_12736);
and U13382 (N_13382,N_12863,N_12557);
and U13383 (N_13383,N_12906,N_12609);
nor U13384 (N_13384,N_12865,N_12563);
and U13385 (N_13385,N_12622,N_12706);
nor U13386 (N_13386,N_12526,N_12505);
or U13387 (N_13387,N_12571,N_12639);
and U13388 (N_13388,N_12686,N_12627);
or U13389 (N_13389,N_12597,N_12685);
nor U13390 (N_13390,N_12722,N_12941);
nor U13391 (N_13391,N_12623,N_12921);
nand U13392 (N_13392,N_12930,N_12987);
xor U13393 (N_13393,N_12840,N_12723);
nand U13394 (N_13394,N_12709,N_12862);
nand U13395 (N_13395,N_12808,N_12846);
or U13396 (N_13396,N_12737,N_12708);
nor U13397 (N_13397,N_12656,N_12842);
or U13398 (N_13398,N_12628,N_12699);
and U13399 (N_13399,N_12861,N_12890);
and U13400 (N_13400,N_12680,N_12656);
nand U13401 (N_13401,N_12794,N_12690);
nand U13402 (N_13402,N_12877,N_12656);
xnor U13403 (N_13403,N_12574,N_12764);
nor U13404 (N_13404,N_12876,N_12784);
or U13405 (N_13405,N_12629,N_12695);
nor U13406 (N_13406,N_12787,N_12705);
and U13407 (N_13407,N_12882,N_12922);
xnor U13408 (N_13408,N_12630,N_12911);
nand U13409 (N_13409,N_12907,N_12549);
nor U13410 (N_13410,N_12755,N_12855);
nor U13411 (N_13411,N_12742,N_12831);
or U13412 (N_13412,N_12602,N_12935);
or U13413 (N_13413,N_12815,N_12578);
and U13414 (N_13414,N_12538,N_12718);
nand U13415 (N_13415,N_12702,N_12807);
xnor U13416 (N_13416,N_12660,N_12587);
nand U13417 (N_13417,N_12719,N_12599);
and U13418 (N_13418,N_12587,N_12759);
and U13419 (N_13419,N_12612,N_12587);
or U13420 (N_13420,N_12615,N_12911);
and U13421 (N_13421,N_12549,N_12704);
nand U13422 (N_13422,N_12605,N_12716);
and U13423 (N_13423,N_12681,N_12676);
and U13424 (N_13424,N_12654,N_12555);
or U13425 (N_13425,N_12516,N_12659);
nand U13426 (N_13426,N_12818,N_12564);
nor U13427 (N_13427,N_12714,N_12957);
xnor U13428 (N_13428,N_12990,N_12710);
xor U13429 (N_13429,N_12733,N_12608);
nand U13430 (N_13430,N_12669,N_12714);
or U13431 (N_13431,N_12870,N_12990);
nor U13432 (N_13432,N_12604,N_12959);
xnor U13433 (N_13433,N_12557,N_12980);
nor U13434 (N_13434,N_12962,N_12690);
or U13435 (N_13435,N_12821,N_12967);
or U13436 (N_13436,N_12582,N_12878);
or U13437 (N_13437,N_12564,N_12587);
nor U13438 (N_13438,N_12727,N_12695);
xnor U13439 (N_13439,N_12626,N_12896);
xnor U13440 (N_13440,N_12774,N_12967);
and U13441 (N_13441,N_12631,N_12686);
and U13442 (N_13442,N_12935,N_12796);
nand U13443 (N_13443,N_12795,N_12900);
nand U13444 (N_13444,N_12579,N_12896);
nand U13445 (N_13445,N_12943,N_12502);
or U13446 (N_13446,N_12770,N_12660);
and U13447 (N_13447,N_12787,N_12877);
or U13448 (N_13448,N_12568,N_12653);
xor U13449 (N_13449,N_12975,N_12880);
xnor U13450 (N_13450,N_12624,N_12816);
nand U13451 (N_13451,N_12547,N_12833);
xor U13452 (N_13452,N_12604,N_12824);
and U13453 (N_13453,N_12577,N_12763);
and U13454 (N_13454,N_12670,N_12806);
or U13455 (N_13455,N_12580,N_12919);
or U13456 (N_13456,N_12598,N_12807);
xor U13457 (N_13457,N_12897,N_12841);
nor U13458 (N_13458,N_12575,N_12804);
nor U13459 (N_13459,N_12963,N_12916);
nor U13460 (N_13460,N_12636,N_12662);
and U13461 (N_13461,N_12593,N_12822);
xnor U13462 (N_13462,N_12748,N_12860);
and U13463 (N_13463,N_12988,N_12733);
nand U13464 (N_13464,N_12808,N_12898);
or U13465 (N_13465,N_12675,N_12871);
nor U13466 (N_13466,N_12837,N_12943);
xor U13467 (N_13467,N_12695,N_12801);
nand U13468 (N_13468,N_12992,N_12678);
or U13469 (N_13469,N_12984,N_12854);
or U13470 (N_13470,N_12508,N_12755);
nand U13471 (N_13471,N_12910,N_12516);
xnor U13472 (N_13472,N_12686,N_12533);
or U13473 (N_13473,N_12645,N_12991);
xnor U13474 (N_13474,N_12996,N_12561);
nor U13475 (N_13475,N_12970,N_12707);
nor U13476 (N_13476,N_12500,N_12835);
xnor U13477 (N_13477,N_12606,N_12832);
xor U13478 (N_13478,N_12803,N_12843);
nand U13479 (N_13479,N_12733,N_12597);
and U13480 (N_13480,N_12861,N_12713);
xnor U13481 (N_13481,N_12598,N_12627);
and U13482 (N_13482,N_12532,N_12650);
xor U13483 (N_13483,N_12894,N_12938);
xnor U13484 (N_13484,N_12984,N_12554);
xor U13485 (N_13485,N_12901,N_12737);
and U13486 (N_13486,N_12894,N_12939);
or U13487 (N_13487,N_12527,N_12696);
nor U13488 (N_13488,N_12800,N_12643);
nor U13489 (N_13489,N_12692,N_12882);
and U13490 (N_13490,N_12607,N_12624);
xnor U13491 (N_13491,N_12570,N_12737);
nor U13492 (N_13492,N_12760,N_12562);
and U13493 (N_13493,N_12773,N_12945);
nor U13494 (N_13494,N_12531,N_12677);
or U13495 (N_13495,N_12735,N_12638);
nand U13496 (N_13496,N_12648,N_12726);
or U13497 (N_13497,N_12562,N_12512);
nand U13498 (N_13498,N_12571,N_12791);
nor U13499 (N_13499,N_12653,N_12860);
nor U13500 (N_13500,N_13014,N_13038);
xnor U13501 (N_13501,N_13159,N_13221);
nand U13502 (N_13502,N_13424,N_13392);
nor U13503 (N_13503,N_13396,N_13316);
and U13504 (N_13504,N_13262,N_13184);
xnor U13505 (N_13505,N_13348,N_13107);
nor U13506 (N_13506,N_13052,N_13298);
nand U13507 (N_13507,N_13323,N_13376);
and U13508 (N_13508,N_13279,N_13450);
or U13509 (N_13509,N_13039,N_13409);
or U13510 (N_13510,N_13374,N_13005);
or U13511 (N_13511,N_13166,N_13010);
nand U13512 (N_13512,N_13434,N_13017);
xor U13513 (N_13513,N_13433,N_13125);
nand U13514 (N_13514,N_13321,N_13296);
xor U13515 (N_13515,N_13241,N_13410);
nand U13516 (N_13516,N_13143,N_13269);
and U13517 (N_13517,N_13160,N_13464);
nand U13518 (N_13518,N_13310,N_13180);
and U13519 (N_13519,N_13449,N_13480);
nand U13520 (N_13520,N_13277,N_13233);
nor U13521 (N_13521,N_13360,N_13476);
nor U13522 (N_13522,N_13225,N_13103);
xnor U13523 (N_13523,N_13220,N_13185);
and U13524 (N_13524,N_13147,N_13398);
and U13525 (N_13525,N_13174,N_13055);
or U13526 (N_13526,N_13265,N_13164);
or U13527 (N_13527,N_13264,N_13253);
and U13528 (N_13528,N_13155,N_13413);
xnor U13529 (N_13529,N_13071,N_13249);
or U13530 (N_13530,N_13332,N_13420);
nand U13531 (N_13531,N_13140,N_13223);
or U13532 (N_13532,N_13157,N_13109);
xor U13533 (N_13533,N_13236,N_13491);
nor U13534 (N_13534,N_13317,N_13407);
nand U13535 (N_13535,N_13423,N_13377);
nor U13536 (N_13536,N_13445,N_13097);
and U13537 (N_13537,N_13403,N_13153);
or U13538 (N_13538,N_13192,N_13475);
nand U13539 (N_13539,N_13059,N_13282);
xnor U13540 (N_13540,N_13176,N_13066);
nand U13541 (N_13541,N_13268,N_13419);
xor U13542 (N_13542,N_13278,N_13337);
xor U13543 (N_13543,N_13388,N_13152);
nand U13544 (N_13544,N_13401,N_13128);
or U13545 (N_13545,N_13026,N_13124);
or U13546 (N_13546,N_13260,N_13254);
and U13547 (N_13547,N_13205,N_13255);
nor U13548 (N_13548,N_13045,N_13297);
and U13549 (N_13549,N_13108,N_13405);
nor U13550 (N_13550,N_13250,N_13497);
or U13551 (N_13551,N_13345,N_13161);
xnor U13552 (N_13552,N_13091,N_13092);
or U13553 (N_13553,N_13436,N_13472);
or U13554 (N_13554,N_13451,N_13425);
nor U13555 (N_13555,N_13415,N_13408);
nor U13556 (N_13556,N_13101,N_13313);
xnor U13557 (N_13557,N_13169,N_13359);
nand U13558 (N_13558,N_13293,N_13439);
and U13559 (N_13559,N_13366,N_13473);
nor U13560 (N_13560,N_13189,N_13181);
or U13561 (N_13561,N_13088,N_13304);
nand U13562 (N_13562,N_13435,N_13341);
or U13563 (N_13563,N_13458,N_13355);
nand U13564 (N_13564,N_13106,N_13467);
nor U13565 (N_13565,N_13358,N_13393);
xnor U13566 (N_13566,N_13133,N_13037);
and U13567 (N_13567,N_13432,N_13117);
nand U13568 (N_13568,N_13163,N_13488);
xor U13569 (N_13569,N_13004,N_13149);
nand U13570 (N_13570,N_13426,N_13350);
nor U13571 (N_13571,N_13102,N_13111);
nor U13572 (N_13572,N_13320,N_13493);
and U13573 (N_13573,N_13110,N_13459);
and U13574 (N_13574,N_13474,N_13251);
nand U13575 (N_13575,N_13150,N_13079);
xor U13576 (N_13576,N_13031,N_13170);
nand U13577 (N_13577,N_13058,N_13072);
or U13578 (N_13578,N_13272,N_13437);
nor U13579 (N_13579,N_13033,N_13077);
xor U13580 (N_13580,N_13378,N_13214);
and U13581 (N_13581,N_13383,N_13146);
and U13582 (N_13582,N_13196,N_13239);
nand U13583 (N_13583,N_13466,N_13482);
xor U13584 (N_13584,N_13200,N_13498);
nor U13585 (N_13585,N_13499,N_13123);
or U13586 (N_13586,N_13002,N_13258);
nor U13587 (N_13587,N_13489,N_13479);
or U13588 (N_13588,N_13369,N_13195);
xor U13589 (N_13589,N_13252,N_13283);
nand U13590 (N_13590,N_13120,N_13063);
xnor U13591 (N_13591,N_13019,N_13447);
nand U13592 (N_13592,N_13421,N_13346);
xor U13593 (N_13593,N_13271,N_13448);
nand U13594 (N_13594,N_13006,N_13070);
or U13595 (N_13595,N_13301,N_13230);
or U13596 (N_13596,N_13391,N_13386);
or U13597 (N_13597,N_13179,N_13216);
nand U13598 (N_13598,N_13406,N_13084);
or U13599 (N_13599,N_13087,N_13057);
or U13600 (N_13600,N_13414,N_13244);
or U13601 (N_13601,N_13203,N_13194);
and U13602 (N_13602,N_13395,N_13330);
nor U13603 (N_13603,N_13371,N_13368);
nor U13604 (N_13604,N_13046,N_13036);
or U13605 (N_13605,N_13427,N_13148);
nand U13606 (N_13606,N_13093,N_13197);
or U13607 (N_13607,N_13324,N_13144);
nor U13608 (N_13608,N_13051,N_13485);
nor U13609 (N_13609,N_13100,N_13023);
nor U13610 (N_13610,N_13053,N_13440);
and U13611 (N_13611,N_13064,N_13370);
xnor U13612 (N_13612,N_13462,N_13336);
nand U13613 (N_13613,N_13168,N_13129);
xnor U13614 (N_13614,N_13471,N_13372);
nor U13615 (N_13615,N_13118,N_13198);
or U13616 (N_13616,N_13492,N_13454);
nor U13617 (N_13617,N_13035,N_13013);
and U13618 (N_13618,N_13135,N_13154);
nor U13619 (N_13619,N_13257,N_13076);
nor U13620 (N_13620,N_13333,N_13380);
or U13621 (N_13621,N_13438,N_13231);
and U13622 (N_13622,N_13204,N_13020);
xor U13623 (N_13623,N_13429,N_13417);
or U13624 (N_13624,N_13306,N_13481);
nand U13625 (N_13625,N_13389,N_13385);
and U13626 (N_13626,N_13151,N_13465);
xor U13627 (N_13627,N_13291,N_13142);
nor U13628 (N_13628,N_13382,N_13238);
xor U13629 (N_13629,N_13276,N_13030);
nand U13630 (N_13630,N_13222,N_13027);
and U13631 (N_13631,N_13218,N_13127);
and U13632 (N_13632,N_13188,N_13325);
nor U13633 (N_13633,N_13281,N_13343);
nand U13634 (N_13634,N_13041,N_13299);
or U13635 (N_13635,N_13114,N_13259);
or U13636 (N_13636,N_13138,N_13029);
nor U13637 (N_13637,N_13182,N_13213);
or U13638 (N_13638,N_13165,N_13217);
nor U13639 (N_13639,N_13040,N_13215);
or U13640 (N_13640,N_13470,N_13292);
nor U13641 (N_13641,N_13080,N_13190);
nand U13642 (N_13642,N_13186,N_13352);
xnor U13643 (N_13643,N_13390,N_13009);
nor U13644 (N_13644,N_13351,N_13096);
nand U13645 (N_13645,N_13422,N_13248);
nor U13646 (N_13646,N_13339,N_13028);
nor U13647 (N_13647,N_13246,N_13043);
nand U13648 (N_13648,N_13210,N_13270);
and U13649 (N_13649,N_13363,N_13089);
nand U13650 (N_13650,N_13418,N_13441);
and U13651 (N_13651,N_13121,N_13209);
nor U13652 (N_13652,N_13007,N_13073);
or U13653 (N_13653,N_13453,N_13444);
xor U13654 (N_13654,N_13496,N_13050);
and U13655 (N_13655,N_13468,N_13187);
xnor U13656 (N_13656,N_13307,N_13086);
xor U13657 (N_13657,N_13237,N_13312);
and U13658 (N_13658,N_13021,N_13347);
nor U13659 (N_13659,N_13075,N_13099);
nand U13660 (N_13660,N_13286,N_13326);
and U13661 (N_13661,N_13314,N_13201);
nand U13662 (N_13662,N_13240,N_13308);
xor U13663 (N_13663,N_13340,N_13290);
or U13664 (N_13664,N_13012,N_13469);
or U13665 (N_13665,N_13207,N_13381);
xnor U13666 (N_13666,N_13139,N_13315);
or U13667 (N_13667,N_13208,N_13126);
nor U13668 (N_13668,N_13305,N_13478);
and U13669 (N_13669,N_13263,N_13494);
xor U13670 (N_13670,N_13047,N_13284);
and U13671 (N_13671,N_13094,N_13361);
or U13672 (N_13672,N_13397,N_13289);
and U13673 (N_13673,N_13056,N_13162);
nor U13674 (N_13674,N_13404,N_13261);
or U13675 (N_13675,N_13384,N_13115);
nand U13676 (N_13676,N_13234,N_13018);
xor U13677 (N_13677,N_13011,N_13034);
or U13678 (N_13678,N_13334,N_13048);
nor U13679 (N_13679,N_13116,N_13078);
and U13680 (N_13680,N_13068,N_13362);
or U13681 (N_13681,N_13191,N_13074);
nand U13682 (N_13682,N_13061,N_13338);
or U13683 (N_13683,N_13367,N_13156);
nor U13684 (N_13684,N_13373,N_13356);
nand U13685 (N_13685,N_13484,N_13311);
xnor U13686 (N_13686,N_13069,N_13394);
or U13687 (N_13687,N_13015,N_13416);
and U13688 (N_13688,N_13461,N_13145);
or U13689 (N_13689,N_13243,N_13452);
or U13690 (N_13690,N_13353,N_13235);
nor U13691 (N_13691,N_13486,N_13122);
or U13692 (N_13692,N_13460,N_13199);
nor U13693 (N_13693,N_13295,N_13067);
nor U13694 (N_13694,N_13227,N_13228);
nor U13695 (N_13695,N_13379,N_13387);
or U13696 (N_13696,N_13167,N_13016);
nand U13697 (N_13697,N_13065,N_13132);
and U13698 (N_13698,N_13171,N_13082);
nor U13699 (N_13699,N_13322,N_13273);
and U13700 (N_13700,N_13364,N_13411);
xnor U13701 (N_13701,N_13266,N_13224);
xor U13702 (N_13702,N_13219,N_13172);
nand U13703 (N_13703,N_13206,N_13232);
or U13704 (N_13704,N_13365,N_13487);
and U13705 (N_13705,N_13247,N_13490);
xor U13706 (N_13706,N_13226,N_13309);
xor U13707 (N_13707,N_13062,N_13303);
xnor U13708 (N_13708,N_13025,N_13455);
or U13709 (N_13709,N_13287,N_13173);
nor U13710 (N_13710,N_13331,N_13022);
or U13711 (N_13711,N_13141,N_13457);
or U13712 (N_13712,N_13104,N_13344);
nand U13713 (N_13713,N_13044,N_13175);
xor U13714 (N_13714,N_13008,N_13335);
or U13715 (N_13715,N_13098,N_13158);
nand U13716 (N_13716,N_13112,N_13267);
xnor U13717 (N_13717,N_13463,N_13329);
nor U13718 (N_13718,N_13177,N_13357);
nand U13719 (N_13719,N_13105,N_13202);
or U13720 (N_13720,N_13412,N_13137);
and U13721 (N_13721,N_13402,N_13285);
nand U13722 (N_13722,N_13245,N_13274);
xnor U13723 (N_13723,N_13083,N_13446);
nor U13724 (N_13724,N_13131,N_13300);
nor U13725 (N_13725,N_13183,N_13193);
nand U13726 (N_13726,N_13483,N_13477);
nor U13727 (N_13727,N_13042,N_13054);
and U13728 (N_13728,N_13456,N_13212);
nor U13729 (N_13729,N_13294,N_13134);
nor U13730 (N_13730,N_13001,N_13319);
xor U13731 (N_13731,N_13328,N_13229);
nand U13732 (N_13732,N_13211,N_13242);
nand U13733 (N_13733,N_13431,N_13318);
and U13734 (N_13734,N_13085,N_13400);
nand U13735 (N_13735,N_13302,N_13442);
or U13736 (N_13736,N_13399,N_13049);
xnor U13737 (N_13737,N_13081,N_13095);
or U13738 (N_13738,N_13113,N_13342);
and U13739 (N_13739,N_13136,N_13119);
and U13740 (N_13740,N_13430,N_13060);
nor U13741 (N_13741,N_13090,N_13428);
nor U13742 (N_13742,N_13443,N_13275);
xnor U13743 (N_13743,N_13327,N_13032);
nor U13744 (N_13744,N_13288,N_13024);
xnor U13745 (N_13745,N_13130,N_13178);
nor U13746 (N_13746,N_13280,N_13256);
nor U13747 (N_13747,N_13349,N_13000);
xnor U13748 (N_13748,N_13495,N_13003);
nor U13749 (N_13749,N_13375,N_13354);
nand U13750 (N_13750,N_13457,N_13035);
nand U13751 (N_13751,N_13086,N_13043);
or U13752 (N_13752,N_13407,N_13354);
xnor U13753 (N_13753,N_13096,N_13291);
or U13754 (N_13754,N_13368,N_13319);
and U13755 (N_13755,N_13301,N_13198);
nand U13756 (N_13756,N_13015,N_13421);
xnor U13757 (N_13757,N_13007,N_13391);
nand U13758 (N_13758,N_13005,N_13178);
xnor U13759 (N_13759,N_13394,N_13074);
or U13760 (N_13760,N_13109,N_13219);
nor U13761 (N_13761,N_13209,N_13157);
nor U13762 (N_13762,N_13285,N_13193);
nand U13763 (N_13763,N_13417,N_13416);
and U13764 (N_13764,N_13220,N_13177);
or U13765 (N_13765,N_13228,N_13498);
and U13766 (N_13766,N_13478,N_13237);
nand U13767 (N_13767,N_13158,N_13336);
or U13768 (N_13768,N_13376,N_13120);
nand U13769 (N_13769,N_13035,N_13348);
or U13770 (N_13770,N_13092,N_13417);
nand U13771 (N_13771,N_13336,N_13432);
nand U13772 (N_13772,N_13129,N_13347);
or U13773 (N_13773,N_13192,N_13365);
and U13774 (N_13774,N_13367,N_13256);
or U13775 (N_13775,N_13438,N_13306);
or U13776 (N_13776,N_13041,N_13386);
xnor U13777 (N_13777,N_13372,N_13263);
and U13778 (N_13778,N_13320,N_13434);
and U13779 (N_13779,N_13082,N_13061);
nand U13780 (N_13780,N_13084,N_13148);
nor U13781 (N_13781,N_13343,N_13475);
nor U13782 (N_13782,N_13448,N_13214);
xor U13783 (N_13783,N_13330,N_13448);
or U13784 (N_13784,N_13315,N_13234);
or U13785 (N_13785,N_13040,N_13138);
or U13786 (N_13786,N_13049,N_13289);
or U13787 (N_13787,N_13188,N_13454);
or U13788 (N_13788,N_13490,N_13340);
and U13789 (N_13789,N_13439,N_13011);
nor U13790 (N_13790,N_13493,N_13331);
or U13791 (N_13791,N_13397,N_13154);
nor U13792 (N_13792,N_13450,N_13066);
or U13793 (N_13793,N_13240,N_13403);
and U13794 (N_13794,N_13441,N_13415);
xnor U13795 (N_13795,N_13004,N_13476);
and U13796 (N_13796,N_13408,N_13292);
xor U13797 (N_13797,N_13370,N_13404);
nand U13798 (N_13798,N_13411,N_13023);
xnor U13799 (N_13799,N_13367,N_13253);
nor U13800 (N_13800,N_13428,N_13180);
xnor U13801 (N_13801,N_13488,N_13254);
nor U13802 (N_13802,N_13425,N_13243);
or U13803 (N_13803,N_13187,N_13024);
nor U13804 (N_13804,N_13025,N_13208);
xor U13805 (N_13805,N_13438,N_13358);
xor U13806 (N_13806,N_13265,N_13314);
nor U13807 (N_13807,N_13035,N_13024);
nand U13808 (N_13808,N_13437,N_13299);
and U13809 (N_13809,N_13016,N_13100);
or U13810 (N_13810,N_13101,N_13042);
nand U13811 (N_13811,N_13148,N_13196);
and U13812 (N_13812,N_13462,N_13467);
and U13813 (N_13813,N_13165,N_13302);
nor U13814 (N_13814,N_13302,N_13071);
xor U13815 (N_13815,N_13157,N_13207);
and U13816 (N_13816,N_13311,N_13200);
nand U13817 (N_13817,N_13435,N_13187);
or U13818 (N_13818,N_13300,N_13390);
nor U13819 (N_13819,N_13028,N_13285);
xnor U13820 (N_13820,N_13023,N_13477);
nor U13821 (N_13821,N_13214,N_13075);
and U13822 (N_13822,N_13284,N_13292);
xor U13823 (N_13823,N_13110,N_13116);
nand U13824 (N_13824,N_13278,N_13285);
nor U13825 (N_13825,N_13117,N_13490);
xor U13826 (N_13826,N_13145,N_13081);
xor U13827 (N_13827,N_13102,N_13170);
xnor U13828 (N_13828,N_13491,N_13030);
nand U13829 (N_13829,N_13070,N_13055);
xnor U13830 (N_13830,N_13447,N_13195);
nand U13831 (N_13831,N_13349,N_13189);
or U13832 (N_13832,N_13057,N_13488);
nor U13833 (N_13833,N_13243,N_13090);
nor U13834 (N_13834,N_13360,N_13291);
and U13835 (N_13835,N_13466,N_13159);
and U13836 (N_13836,N_13364,N_13431);
nand U13837 (N_13837,N_13355,N_13105);
xnor U13838 (N_13838,N_13469,N_13054);
and U13839 (N_13839,N_13186,N_13222);
and U13840 (N_13840,N_13181,N_13456);
or U13841 (N_13841,N_13146,N_13070);
nand U13842 (N_13842,N_13440,N_13081);
nor U13843 (N_13843,N_13470,N_13455);
nand U13844 (N_13844,N_13387,N_13190);
and U13845 (N_13845,N_13415,N_13341);
or U13846 (N_13846,N_13299,N_13311);
and U13847 (N_13847,N_13413,N_13184);
nor U13848 (N_13848,N_13430,N_13262);
xor U13849 (N_13849,N_13422,N_13012);
or U13850 (N_13850,N_13378,N_13225);
xnor U13851 (N_13851,N_13341,N_13087);
nor U13852 (N_13852,N_13208,N_13458);
nor U13853 (N_13853,N_13466,N_13434);
nand U13854 (N_13854,N_13162,N_13151);
and U13855 (N_13855,N_13176,N_13406);
or U13856 (N_13856,N_13066,N_13112);
or U13857 (N_13857,N_13246,N_13008);
xnor U13858 (N_13858,N_13465,N_13273);
xnor U13859 (N_13859,N_13222,N_13390);
xnor U13860 (N_13860,N_13454,N_13212);
nand U13861 (N_13861,N_13070,N_13497);
nor U13862 (N_13862,N_13206,N_13116);
and U13863 (N_13863,N_13055,N_13456);
or U13864 (N_13864,N_13080,N_13004);
or U13865 (N_13865,N_13232,N_13408);
nand U13866 (N_13866,N_13498,N_13224);
xnor U13867 (N_13867,N_13113,N_13161);
nand U13868 (N_13868,N_13445,N_13344);
or U13869 (N_13869,N_13053,N_13354);
or U13870 (N_13870,N_13321,N_13269);
nor U13871 (N_13871,N_13059,N_13411);
nor U13872 (N_13872,N_13460,N_13067);
xnor U13873 (N_13873,N_13400,N_13009);
nand U13874 (N_13874,N_13423,N_13142);
nand U13875 (N_13875,N_13203,N_13318);
nor U13876 (N_13876,N_13488,N_13470);
and U13877 (N_13877,N_13361,N_13179);
or U13878 (N_13878,N_13268,N_13381);
and U13879 (N_13879,N_13181,N_13137);
nor U13880 (N_13880,N_13034,N_13094);
and U13881 (N_13881,N_13344,N_13198);
or U13882 (N_13882,N_13349,N_13060);
nand U13883 (N_13883,N_13217,N_13329);
nand U13884 (N_13884,N_13473,N_13254);
and U13885 (N_13885,N_13236,N_13248);
xnor U13886 (N_13886,N_13478,N_13115);
and U13887 (N_13887,N_13261,N_13313);
nor U13888 (N_13888,N_13074,N_13197);
nand U13889 (N_13889,N_13295,N_13001);
nand U13890 (N_13890,N_13227,N_13198);
xor U13891 (N_13891,N_13468,N_13414);
xnor U13892 (N_13892,N_13094,N_13183);
or U13893 (N_13893,N_13448,N_13398);
or U13894 (N_13894,N_13012,N_13001);
nor U13895 (N_13895,N_13043,N_13163);
xor U13896 (N_13896,N_13204,N_13246);
or U13897 (N_13897,N_13152,N_13130);
nand U13898 (N_13898,N_13065,N_13000);
or U13899 (N_13899,N_13208,N_13388);
or U13900 (N_13900,N_13286,N_13006);
or U13901 (N_13901,N_13197,N_13309);
nand U13902 (N_13902,N_13244,N_13465);
and U13903 (N_13903,N_13385,N_13203);
nor U13904 (N_13904,N_13206,N_13211);
and U13905 (N_13905,N_13301,N_13411);
nor U13906 (N_13906,N_13290,N_13377);
or U13907 (N_13907,N_13342,N_13101);
and U13908 (N_13908,N_13095,N_13488);
nor U13909 (N_13909,N_13069,N_13363);
nand U13910 (N_13910,N_13276,N_13384);
and U13911 (N_13911,N_13336,N_13118);
nand U13912 (N_13912,N_13060,N_13311);
nand U13913 (N_13913,N_13294,N_13495);
xor U13914 (N_13914,N_13341,N_13166);
nor U13915 (N_13915,N_13380,N_13319);
and U13916 (N_13916,N_13260,N_13104);
nand U13917 (N_13917,N_13092,N_13313);
and U13918 (N_13918,N_13407,N_13167);
or U13919 (N_13919,N_13215,N_13283);
and U13920 (N_13920,N_13252,N_13091);
xor U13921 (N_13921,N_13421,N_13475);
xor U13922 (N_13922,N_13241,N_13395);
or U13923 (N_13923,N_13382,N_13208);
xnor U13924 (N_13924,N_13300,N_13428);
nor U13925 (N_13925,N_13017,N_13159);
or U13926 (N_13926,N_13406,N_13183);
and U13927 (N_13927,N_13425,N_13268);
or U13928 (N_13928,N_13052,N_13408);
xnor U13929 (N_13929,N_13272,N_13315);
and U13930 (N_13930,N_13387,N_13022);
nand U13931 (N_13931,N_13025,N_13412);
nand U13932 (N_13932,N_13368,N_13266);
nand U13933 (N_13933,N_13158,N_13084);
xnor U13934 (N_13934,N_13129,N_13029);
nor U13935 (N_13935,N_13129,N_13412);
and U13936 (N_13936,N_13395,N_13391);
nor U13937 (N_13937,N_13176,N_13230);
and U13938 (N_13938,N_13137,N_13491);
nor U13939 (N_13939,N_13257,N_13434);
and U13940 (N_13940,N_13195,N_13327);
or U13941 (N_13941,N_13048,N_13267);
nand U13942 (N_13942,N_13377,N_13076);
or U13943 (N_13943,N_13169,N_13185);
nand U13944 (N_13944,N_13002,N_13389);
or U13945 (N_13945,N_13312,N_13241);
nand U13946 (N_13946,N_13035,N_13071);
and U13947 (N_13947,N_13087,N_13196);
nor U13948 (N_13948,N_13344,N_13238);
and U13949 (N_13949,N_13133,N_13280);
nand U13950 (N_13950,N_13152,N_13208);
and U13951 (N_13951,N_13186,N_13212);
or U13952 (N_13952,N_13470,N_13157);
xnor U13953 (N_13953,N_13452,N_13359);
nand U13954 (N_13954,N_13372,N_13196);
nor U13955 (N_13955,N_13266,N_13115);
or U13956 (N_13956,N_13143,N_13074);
nor U13957 (N_13957,N_13368,N_13223);
or U13958 (N_13958,N_13296,N_13020);
nand U13959 (N_13959,N_13410,N_13283);
and U13960 (N_13960,N_13489,N_13374);
and U13961 (N_13961,N_13073,N_13303);
nand U13962 (N_13962,N_13222,N_13375);
nor U13963 (N_13963,N_13385,N_13182);
nor U13964 (N_13964,N_13396,N_13137);
and U13965 (N_13965,N_13209,N_13341);
xnor U13966 (N_13966,N_13066,N_13181);
xor U13967 (N_13967,N_13477,N_13137);
nor U13968 (N_13968,N_13256,N_13305);
and U13969 (N_13969,N_13455,N_13281);
or U13970 (N_13970,N_13478,N_13160);
and U13971 (N_13971,N_13272,N_13434);
or U13972 (N_13972,N_13248,N_13436);
and U13973 (N_13973,N_13188,N_13344);
and U13974 (N_13974,N_13491,N_13364);
or U13975 (N_13975,N_13210,N_13023);
and U13976 (N_13976,N_13119,N_13189);
and U13977 (N_13977,N_13202,N_13252);
nor U13978 (N_13978,N_13343,N_13161);
or U13979 (N_13979,N_13449,N_13132);
nor U13980 (N_13980,N_13099,N_13005);
nand U13981 (N_13981,N_13084,N_13432);
and U13982 (N_13982,N_13091,N_13488);
xor U13983 (N_13983,N_13163,N_13477);
or U13984 (N_13984,N_13014,N_13098);
and U13985 (N_13985,N_13256,N_13431);
nor U13986 (N_13986,N_13148,N_13377);
nor U13987 (N_13987,N_13166,N_13373);
and U13988 (N_13988,N_13324,N_13071);
or U13989 (N_13989,N_13470,N_13189);
nand U13990 (N_13990,N_13379,N_13238);
and U13991 (N_13991,N_13244,N_13427);
xnor U13992 (N_13992,N_13319,N_13307);
nor U13993 (N_13993,N_13297,N_13427);
nand U13994 (N_13994,N_13401,N_13499);
and U13995 (N_13995,N_13153,N_13004);
nand U13996 (N_13996,N_13363,N_13044);
xnor U13997 (N_13997,N_13321,N_13383);
nor U13998 (N_13998,N_13298,N_13051);
and U13999 (N_13999,N_13182,N_13369);
or U14000 (N_14000,N_13692,N_13915);
nor U14001 (N_14001,N_13694,N_13548);
and U14002 (N_14002,N_13547,N_13695);
nor U14003 (N_14003,N_13881,N_13959);
nand U14004 (N_14004,N_13968,N_13823);
nor U14005 (N_14005,N_13771,N_13923);
nor U14006 (N_14006,N_13888,N_13976);
xor U14007 (N_14007,N_13697,N_13797);
or U14008 (N_14008,N_13861,N_13805);
or U14009 (N_14009,N_13729,N_13570);
nor U14010 (N_14010,N_13782,N_13524);
nor U14011 (N_14011,N_13739,N_13641);
and U14012 (N_14012,N_13618,N_13855);
nor U14013 (N_14013,N_13671,N_13848);
nand U14014 (N_14014,N_13665,N_13687);
nand U14015 (N_14015,N_13520,N_13889);
xnor U14016 (N_14016,N_13660,N_13741);
xor U14017 (N_14017,N_13877,N_13972);
xnor U14018 (N_14018,N_13914,N_13519);
and U14019 (N_14019,N_13643,N_13640);
xor U14020 (N_14020,N_13613,N_13755);
or U14021 (N_14021,N_13700,N_13509);
nand U14022 (N_14022,N_13929,N_13963);
or U14023 (N_14023,N_13569,N_13607);
and U14024 (N_14024,N_13874,N_13710);
and U14025 (N_14025,N_13666,N_13880);
nand U14026 (N_14026,N_13870,N_13605);
nand U14027 (N_14027,N_13875,N_13730);
nor U14028 (N_14028,N_13985,N_13557);
and U14029 (N_14029,N_13952,N_13884);
and U14030 (N_14030,N_13562,N_13693);
and U14031 (N_14031,N_13736,N_13718);
nand U14032 (N_14032,N_13908,N_13811);
nor U14033 (N_14033,N_13876,N_13529);
xnor U14034 (N_14034,N_13933,N_13603);
nand U14035 (N_14035,N_13712,N_13584);
xnor U14036 (N_14036,N_13611,N_13826);
nor U14037 (N_14037,N_13589,N_13924);
nand U14038 (N_14038,N_13955,N_13792);
xnor U14039 (N_14039,N_13789,N_13659);
xnor U14040 (N_14040,N_13954,N_13673);
xor U14041 (N_14041,N_13701,N_13973);
nor U14042 (N_14042,N_13614,N_13636);
xor U14043 (N_14043,N_13910,N_13651);
xor U14044 (N_14044,N_13871,N_13819);
or U14045 (N_14045,N_13745,N_13844);
nand U14046 (N_14046,N_13662,N_13537);
and U14047 (N_14047,N_13765,N_13859);
nor U14048 (N_14048,N_13803,N_13586);
nand U14049 (N_14049,N_13783,N_13582);
nand U14050 (N_14050,N_13732,N_13540);
nand U14051 (N_14051,N_13912,N_13681);
nor U14052 (N_14052,N_13837,N_13958);
and U14053 (N_14053,N_13802,N_13523);
xnor U14054 (N_14054,N_13709,N_13772);
xnor U14055 (N_14055,N_13527,N_13901);
xor U14056 (N_14056,N_13868,N_13719);
and U14057 (N_14057,N_13935,N_13501);
or U14058 (N_14058,N_13720,N_13886);
or U14059 (N_14059,N_13946,N_13940);
nor U14060 (N_14060,N_13781,N_13635);
nand U14061 (N_14061,N_13865,N_13936);
nand U14062 (N_14062,N_13647,N_13894);
and U14063 (N_14063,N_13559,N_13835);
nor U14064 (N_14064,N_13810,N_13853);
nor U14065 (N_14065,N_13577,N_13734);
nor U14066 (N_14066,N_13911,N_13749);
or U14067 (N_14067,N_13552,N_13674);
nand U14068 (N_14068,N_13907,N_13689);
and U14069 (N_14069,N_13816,N_13573);
xnor U14070 (N_14070,N_13752,N_13615);
nand U14071 (N_14071,N_13938,N_13746);
or U14072 (N_14072,N_13794,N_13669);
xor U14073 (N_14073,N_13798,N_13622);
or U14074 (N_14074,N_13795,N_13944);
nor U14075 (N_14075,N_13599,N_13546);
and U14076 (N_14076,N_13895,N_13767);
xnor U14077 (N_14077,N_13808,N_13536);
or U14078 (N_14078,N_13762,N_13948);
or U14079 (N_14079,N_13813,N_13740);
and U14080 (N_14080,N_13517,N_13956);
nand U14081 (N_14081,N_13977,N_13757);
and U14082 (N_14082,N_13637,N_13715);
nand U14083 (N_14083,N_13723,N_13898);
nor U14084 (N_14084,N_13631,N_13626);
xnor U14085 (N_14085,N_13587,N_13549);
nand U14086 (N_14086,N_13775,N_13983);
or U14087 (N_14087,N_13576,N_13686);
nand U14088 (N_14088,N_13790,N_13706);
xnor U14089 (N_14089,N_13885,N_13621);
and U14090 (N_14090,N_13508,N_13610);
and U14091 (N_14091,N_13761,N_13512);
nor U14092 (N_14092,N_13581,N_13604);
xor U14093 (N_14093,N_13539,N_13769);
xnor U14094 (N_14094,N_13860,N_13751);
nand U14095 (N_14095,N_13941,N_13590);
and U14096 (N_14096,N_13992,N_13830);
nand U14097 (N_14097,N_13677,N_13937);
xnor U14098 (N_14098,N_13831,N_13784);
nor U14099 (N_14099,N_13690,N_13661);
xnor U14100 (N_14100,N_13550,N_13787);
nor U14101 (N_14101,N_13991,N_13617);
or U14102 (N_14102,N_13595,N_13768);
or U14103 (N_14103,N_13841,N_13777);
nor U14104 (N_14104,N_13864,N_13747);
xor U14105 (N_14105,N_13542,N_13834);
nand U14106 (N_14106,N_13516,N_13619);
or U14107 (N_14107,N_13644,N_13845);
nand U14108 (N_14108,N_13857,N_13571);
nand U14109 (N_14109,N_13737,N_13818);
xor U14110 (N_14110,N_13657,N_13564);
xor U14111 (N_14111,N_13869,N_13926);
xnor U14112 (N_14112,N_13708,N_13971);
xnor U14113 (N_14113,N_13591,N_13713);
nand U14114 (N_14114,N_13598,N_13817);
nand U14115 (N_14115,N_13957,N_13993);
or U14116 (N_14116,N_13629,N_13634);
xor U14117 (N_14117,N_13764,N_13535);
or U14118 (N_14118,N_13832,N_13851);
xnor U14119 (N_14119,N_13989,N_13939);
xnor U14120 (N_14120,N_13878,N_13879);
xor U14121 (N_14121,N_13648,N_13525);
nand U14122 (N_14122,N_13545,N_13703);
or U14123 (N_14123,N_13685,N_13829);
nand U14124 (N_14124,N_13670,N_13563);
nor U14125 (N_14125,N_13846,N_13932);
and U14126 (N_14126,N_13724,N_13779);
xor U14127 (N_14127,N_13986,N_13773);
or U14128 (N_14128,N_13696,N_13902);
xnor U14129 (N_14129,N_13825,N_13903);
or U14130 (N_14130,N_13791,N_13551);
and U14131 (N_14131,N_13975,N_13822);
nand U14132 (N_14132,N_13873,N_13632);
xnor U14133 (N_14133,N_13616,N_13961);
or U14134 (N_14134,N_13728,N_13964);
nand U14135 (N_14135,N_13801,N_13583);
xor U14136 (N_14136,N_13754,N_13649);
and U14137 (N_14137,N_13530,N_13565);
or U14138 (N_14138,N_13814,N_13854);
nand U14139 (N_14139,N_13566,N_13962);
nand U14140 (N_14140,N_13609,N_13942);
or U14141 (N_14141,N_13763,N_13554);
and U14142 (N_14142,N_13842,N_13639);
and U14143 (N_14143,N_13890,N_13684);
xnor U14144 (N_14144,N_13664,N_13620);
nand U14145 (N_14145,N_13922,N_13707);
or U14146 (N_14146,N_13691,N_13653);
nor U14147 (N_14147,N_13522,N_13780);
or U14148 (N_14148,N_13996,N_13553);
and U14149 (N_14149,N_13588,N_13978);
xnor U14150 (N_14150,N_13507,N_13678);
or U14151 (N_14151,N_13579,N_13943);
or U14152 (N_14152,N_13995,N_13960);
or U14153 (N_14153,N_13731,N_13518);
nand U14154 (N_14154,N_13514,N_13897);
xor U14155 (N_14155,N_13919,N_13920);
xor U14156 (N_14156,N_13774,N_13600);
nor U14157 (N_14157,N_13863,N_13558);
nand U14158 (N_14158,N_13916,N_13756);
or U14159 (N_14159,N_13680,N_13984);
and U14160 (N_14160,N_13650,N_13727);
xor U14161 (N_14161,N_13716,N_13623);
and U14162 (N_14162,N_13904,N_13882);
or U14163 (N_14163,N_13836,N_13658);
nand U14164 (N_14164,N_13887,N_13528);
and U14165 (N_14165,N_13750,N_13997);
nor U14166 (N_14166,N_13627,N_13821);
xor U14167 (N_14167,N_13606,N_13913);
xnor U14168 (N_14168,N_13515,N_13820);
nor U14169 (N_14169,N_13990,N_13796);
or U14170 (N_14170,N_13505,N_13556);
xor U14171 (N_14171,N_13891,N_13656);
nor U14172 (N_14172,N_13711,N_13793);
nor U14173 (N_14173,N_13714,N_13905);
nand U14174 (N_14174,N_13947,N_13642);
or U14175 (N_14175,N_13645,N_13506);
and U14176 (N_14176,N_13892,N_13800);
or U14177 (N_14177,N_13743,N_13951);
xnor U14178 (N_14178,N_13828,N_13578);
nor U14179 (N_14179,N_13511,N_13998);
and U14180 (N_14180,N_13928,N_13510);
or U14181 (N_14181,N_13602,N_13738);
or U14182 (N_14182,N_13799,N_13502);
xor U14183 (N_14183,N_13766,N_13717);
nor U14184 (N_14184,N_13572,N_13807);
xnor U14185 (N_14185,N_13945,N_13596);
nand U14186 (N_14186,N_13663,N_13900);
or U14187 (N_14187,N_13883,N_13654);
nand U14188 (N_14188,N_13698,N_13624);
and U14189 (N_14189,N_13840,N_13534);
nand U14190 (N_14190,N_13909,N_13679);
or U14191 (N_14191,N_13833,N_13504);
or U14192 (N_14192,N_13950,N_13965);
or U14193 (N_14193,N_13533,N_13594);
xor U14194 (N_14194,N_13560,N_13981);
nor U14195 (N_14195,N_13608,N_13721);
xor U14196 (N_14196,N_13704,N_13858);
nand U14197 (N_14197,N_13896,N_13770);
xnor U14198 (N_14198,N_13850,N_13899);
or U14199 (N_14199,N_13849,N_13521);
and U14200 (N_14200,N_13675,N_13702);
or U14201 (N_14201,N_13628,N_13967);
nand U14202 (N_14202,N_13760,N_13531);
nand U14203 (N_14203,N_13815,N_13742);
and U14204 (N_14204,N_13776,N_13974);
nor U14205 (N_14205,N_13544,N_13970);
or U14206 (N_14206,N_13538,N_13748);
xor U14207 (N_14207,N_13580,N_13682);
nor U14208 (N_14208,N_13667,N_13918);
or U14209 (N_14209,N_13931,N_13778);
xor U14210 (N_14210,N_13526,N_13574);
and U14211 (N_14211,N_13838,N_13966);
nand U14212 (N_14212,N_13585,N_13812);
and U14213 (N_14213,N_13735,N_13809);
xnor U14214 (N_14214,N_13655,N_13575);
xor U14215 (N_14215,N_13788,N_13930);
or U14216 (N_14216,N_13867,N_13688);
nor U14217 (N_14217,N_13969,N_13839);
or U14218 (N_14218,N_13543,N_13872);
nand U14219 (N_14219,N_13668,N_13733);
and U14220 (N_14220,N_13555,N_13906);
nand U14221 (N_14221,N_13567,N_13725);
xor U14222 (N_14222,N_13541,N_13722);
nand U14223 (N_14223,N_13758,N_13979);
xnor U14224 (N_14224,N_13921,N_13699);
or U14225 (N_14225,N_13852,N_13994);
nor U14226 (N_14226,N_13532,N_13638);
nor U14227 (N_14227,N_13987,N_13568);
xor U14228 (N_14228,N_13843,N_13705);
nand U14229 (N_14229,N_13934,N_13917);
xnor U14230 (N_14230,N_13601,N_13785);
and U14231 (N_14231,N_13726,N_13625);
xnor U14232 (N_14232,N_13856,N_13988);
or U14233 (N_14233,N_13949,N_13753);
nor U14234 (N_14234,N_13683,N_13513);
or U14235 (N_14235,N_13806,N_13927);
or U14236 (N_14236,N_13866,N_13503);
nand U14237 (N_14237,N_13804,N_13982);
nor U14238 (N_14238,N_13744,N_13633);
xnor U14239 (N_14239,N_13652,N_13862);
xnor U14240 (N_14240,N_13893,N_13847);
or U14241 (N_14241,N_13925,N_13786);
nor U14242 (N_14242,N_13672,N_13597);
or U14243 (N_14243,N_13759,N_13500);
and U14244 (N_14244,N_13630,N_13612);
nor U14245 (N_14245,N_13824,N_13646);
nor U14246 (N_14246,N_13561,N_13676);
or U14247 (N_14247,N_13592,N_13827);
xor U14248 (N_14248,N_13593,N_13999);
nand U14249 (N_14249,N_13953,N_13980);
nand U14250 (N_14250,N_13568,N_13559);
xnor U14251 (N_14251,N_13857,N_13636);
nor U14252 (N_14252,N_13763,N_13701);
or U14253 (N_14253,N_13526,N_13643);
xnor U14254 (N_14254,N_13531,N_13685);
nand U14255 (N_14255,N_13874,N_13924);
or U14256 (N_14256,N_13985,N_13704);
and U14257 (N_14257,N_13796,N_13526);
nand U14258 (N_14258,N_13578,N_13798);
or U14259 (N_14259,N_13863,N_13643);
and U14260 (N_14260,N_13627,N_13840);
nand U14261 (N_14261,N_13737,N_13947);
nor U14262 (N_14262,N_13969,N_13797);
nand U14263 (N_14263,N_13646,N_13826);
xor U14264 (N_14264,N_13549,N_13778);
and U14265 (N_14265,N_13629,N_13597);
nor U14266 (N_14266,N_13648,N_13969);
xor U14267 (N_14267,N_13965,N_13952);
nor U14268 (N_14268,N_13630,N_13650);
xnor U14269 (N_14269,N_13550,N_13894);
or U14270 (N_14270,N_13818,N_13849);
nand U14271 (N_14271,N_13557,N_13536);
nor U14272 (N_14272,N_13879,N_13584);
nand U14273 (N_14273,N_13857,N_13668);
xnor U14274 (N_14274,N_13995,N_13700);
and U14275 (N_14275,N_13693,N_13549);
or U14276 (N_14276,N_13526,N_13571);
and U14277 (N_14277,N_13689,N_13526);
nor U14278 (N_14278,N_13677,N_13745);
or U14279 (N_14279,N_13844,N_13807);
or U14280 (N_14280,N_13963,N_13752);
and U14281 (N_14281,N_13647,N_13733);
nor U14282 (N_14282,N_13796,N_13646);
xor U14283 (N_14283,N_13954,N_13883);
nor U14284 (N_14284,N_13936,N_13990);
or U14285 (N_14285,N_13906,N_13859);
or U14286 (N_14286,N_13798,N_13695);
or U14287 (N_14287,N_13702,N_13998);
nand U14288 (N_14288,N_13535,N_13826);
xnor U14289 (N_14289,N_13516,N_13505);
xnor U14290 (N_14290,N_13796,N_13589);
and U14291 (N_14291,N_13581,N_13729);
xnor U14292 (N_14292,N_13937,N_13880);
nor U14293 (N_14293,N_13907,N_13739);
and U14294 (N_14294,N_13763,N_13711);
or U14295 (N_14295,N_13522,N_13914);
nor U14296 (N_14296,N_13517,N_13806);
and U14297 (N_14297,N_13540,N_13726);
nand U14298 (N_14298,N_13967,N_13940);
or U14299 (N_14299,N_13923,N_13837);
and U14300 (N_14300,N_13533,N_13506);
xnor U14301 (N_14301,N_13515,N_13678);
nor U14302 (N_14302,N_13905,N_13804);
xor U14303 (N_14303,N_13701,N_13710);
nand U14304 (N_14304,N_13972,N_13563);
nor U14305 (N_14305,N_13668,N_13968);
or U14306 (N_14306,N_13880,N_13908);
xor U14307 (N_14307,N_13894,N_13907);
nand U14308 (N_14308,N_13629,N_13756);
and U14309 (N_14309,N_13848,N_13766);
or U14310 (N_14310,N_13788,N_13940);
and U14311 (N_14311,N_13535,N_13850);
and U14312 (N_14312,N_13990,N_13921);
or U14313 (N_14313,N_13977,N_13767);
xnor U14314 (N_14314,N_13832,N_13934);
and U14315 (N_14315,N_13585,N_13877);
nand U14316 (N_14316,N_13952,N_13861);
and U14317 (N_14317,N_13772,N_13742);
nor U14318 (N_14318,N_13773,N_13910);
or U14319 (N_14319,N_13942,N_13824);
nand U14320 (N_14320,N_13791,N_13522);
nor U14321 (N_14321,N_13588,N_13695);
or U14322 (N_14322,N_13888,N_13882);
nand U14323 (N_14323,N_13644,N_13917);
or U14324 (N_14324,N_13785,N_13797);
and U14325 (N_14325,N_13643,N_13825);
nand U14326 (N_14326,N_13939,N_13947);
and U14327 (N_14327,N_13786,N_13996);
nand U14328 (N_14328,N_13908,N_13527);
and U14329 (N_14329,N_13872,N_13859);
nand U14330 (N_14330,N_13805,N_13844);
xor U14331 (N_14331,N_13521,N_13971);
nand U14332 (N_14332,N_13862,N_13924);
nor U14333 (N_14333,N_13635,N_13790);
or U14334 (N_14334,N_13677,N_13692);
xnor U14335 (N_14335,N_13566,N_13693);
or U14336 (N_14336,N_13996,N_13531);
nor U14337 (N_14337,N_13622,N_13700);
or U14338 (N_14338,N_13750,N_13673);
nand U14339 (N_14339,N_13927,N_13723);
nor U14340 (N_14340,N_13527,N_13754);
nor U14341 (N_14341,N_13593,N_13885);
and U14342 (N_14342,N_13934,N_13529);
nand U14343 (N_14343,N_13678,N_13505);
xnor U14344 (N_14344,N_13811,N_13518);
or U14345 (N_14345,N_13707,N_13591);
xnor U14346 (N_14346,N_13657,N_13635);
and U14347 (N_14347,N_13956,N_13548);
nand U14348 (N_14348,N_13713,N_13916);
xnor U14349 (N_14349,N_13532,N_13941);
nand U14350 (N_14350,N_13557,N_13559);
or U14351 (N_14351,N_13915,N_13840);
or U14352 (N_14352,N_13824,N_13787);
or U14353 (N_14353,N_13875,N_13593);
nor U14354 (N_14354,N_13909,N_13786);
nand U14355 (N_14355,N_13837,N_13724);
xor U14356 (N_14356,N_13682,N_13503);
or U14357 (N_14357,N_13609,N_13764);
nand U14358 (N_14358,N_13725,N_13519);
xor U14359 (N_14359,N_13798,N_13955);
xor U14360 (N_14360,N_13830,N_13677);
nor U14361 (N_14361,N_13635,N_13893);
or U14362 (N_14362,N_13900,N_13822);
nand U14363 (N_14363,N_13955,N_13770);
xor U14364 (N_14364,N_13908,N_13863);
xor U14365 (N_14365,N_13859,N_13587);
nor U14366 (N_14366,N_13625,N_13638);
or U14367 (N_14367,N_13907,N_13766);
or U14368 (N_14368,N_13997,N_13987);
and U14369 (N_14369,N_13930,N_13722);
or U14370 (N_14370,N_13640,N_13611);
or U14371 (N_14371,N_13923,N_13691);
and U14372 (N_14372,N_13510,N_13815);
nor U14373 (N_14373,N_13844,N_13526);
and U14374 (N_14374,N_13594,N_13916);
xnor U14375 (N_14375,N_13835,N_13945);
nand U14376 (N_14376,N_13887,N_13854);
xnor U14377 (N_14377,N_13630,N_13806);
nor U14378 (N_14378,N_13820,N_13544);
and U14379 (N_14379,N_13711,N_13599);
nand U14380 (N_14380,N_13992,N_13858);
or U14381 (N_14381,N_13728,N_13789);
or U14382 (N_14382,N_13670,N_13655);
and U14383 (N_14383,N_13896,N_13607);
or U14384 (N_14384,N_13580,N_13881);
and U14385 (N_14385,N_13503,N_13799);
or U14386 (N_14386,N_13623,N_13677);
and U14387 (N_14387,N_13675,N_13549);
and U14388 (N_14388,N_13529,N_13697);
nand U14389 (N_14389,N_13543,N_13676);
and U14390 (N_14390,N_13874,N_13723);
and U14391 (N_14391,N_13789,N_13947);
or U14392 (N_14392,N_13652,N_13584);
nand U14393 (N_14393,N_13810,N_13844);
or U14394 (N_14394,N_13724,N_13540);
nor U14395 (N_14395,N_13669,N_13619);
xor U14396 (N_14396,N_13718,N_13576);
nor U14397 (N_14397,N_13975,N_13559);
nand U14398 (N_14398,N_13574,N_13692);
or U14399 (N_14399,N_13780,N_13801);
or U14400 (N_14400,N_13524,N_13754);
nand U14401 (N_14401,N_13942,N_13805);
nor U14402 (N_14402,N_13608,N_13977);
xnor U14403 (N_14403,N_13586,N_13841);
nor U14404 (N_14404,N_13745,N_13819);
nand U14405 (N_14405,N_13691,N_13804);
nand U14406 (N_14406,N_13500,N_13851);
nor U14407 (N_14407,N_13604,N_13612);
and U14408 (N_14408,N_13952,N_13781);
nor U14409 (N_14409,N_13554,N_13549);
nor U14410 (N_14410,N_13723,N_13847);
xnor U14411 (N_14411,N_13715,N_13733);
xnor U14412 (N_14412,N_13629,N_13859);
nor U14413 (N_14413,N_13643,N_13806);
or U14414 (N_14414,N_13529,N_13765);
and U14415 (N_14415,N_13976,N_13949);
nand U14416 (N_14416,N_13599,N_13591);
nor U14417 (N_14417,N_13647,N_13563);
and U14418 (N_14418,N_13872,N_13696);
nand U14419 (N_14419,N_13924,N_13628);
or U14420 (N_14420,N_13752,N_13920);
or U14421 (N_14421,N_13659,N_13837);
xor U14422 (N_14422,N_13769,N_13988);
nor U14423 (N_14423,N_13678,N_13613);
xnor U14424 (N_14424,N_13667,N_13772);
nor U14425 (N_14425,N_13985,N_13818);
and U14426 (N_14426,N_13956,N_13994);
or U14427 (N_14427,N_13810,N_13802);
nand U14428 (N_14428,N_13749,N_13816);
and U14429 (N_14429,N_13872,N_13734);
nand U14430 (N_14430,N_13589,N_13853);
nor U14431 (N_14431,N_13815,N_13746);
nand U14432 (N_14432,N_13725,N_13784);
or U14433 (N_14433,N_13808,N_13829);
xor U14434 (N_14434,N_13918,N_13759);
xnor U14435 (N_14435,N_13514,N_13850);
nor U14436 (N_14436,N_13555,N_13520);
nor U14437 (N_14437,N_13543,N_13920);
nor U14438 (N_14438,N_13576,N_13564);
and U14439 (N_14439,N_13852,N_13924);
and U14440 (N_14440,N_13690,N_13868);
nand U14441 (N_14441,N_13510,N_13514);
nor U14442 (N_14442,N_13937,N_13512);
nor U14443 (N_14443,N_13545,N_13916);
and U14444 (N_14444,N_13828,N_13730);
xnor U14445 (N_14445,N_13657,N_13998);
nor U14446 (N_14446,N_13797,N_13632);
nand U14447 (N_14447,N_13597,N_13902);
xnor U14448 (N_14448,N_13995,N_13981);
or U14449 (N_14449,N_13646,N_13510);
and U14450 (N_14450,N_13758,N_13701);
nand U14451 (N_14451,N_13662,N_13978);
nor U14452 (N_14452,N_13822,N_13767);
and U14453 (N_14453,N_13846,N_13623);
or U14454 (N_14454,N_13849,N_13957);
xnor U14455 (N_14455,N_13550,N_13526);
and U14456 (N_14456,N_13744,N_13878);
or U14457 (N_14457,N_13741,N_13687);
nor U14458 (N_14458,N_13651,N_13766);
xnor U14459 (N_14459,N_13594,N_13842);
nand U14460 (N_14460,N_13862,N_13883);
nand U14461 (N_14461,N_13704,N_13559);
nor U14462 (N_14462,N_13709,N_13683);
or U14463 (N_14463,N_13734,N_13893);
and U14464 (N_14464,N_13995,N_13950);
nor U14465 (N_14465,N_13850,N_13935);
and U14466 (N_14466,N_13539,N_13736);
or U14467 (N_14467,N_13509,N_13934);
nor U14468 (N_14468,N_13579,N_13620);
nand U14469 (N_14469,N_13736,N_13762);
xnor U14470 (N_14470,N_13593,N_13530);
nand U14471 (N_14471,N_13931,N_13663);
and U14472 (N_14472,N_13684,N_13662);
or U14473 (N_14473,N_13867,N_13896);
xnor U14474 (N_14474,N_13850,N_13642);
nand U14475 (N_14475,N_13701,N_13820);
nor U14476 (N_14476,N_13752,N_13930);
nor U14477 (N_14477,N_13997,N_13971);
or U14478 (N_14478,N_13720,N_13965);
xor U14479 (N_14479,N_13751,N_13818);
and U14480 (N_14480,N_13940,N_13930);
and U14481 (N_14481,N_13755,N_13690);
and U14482 (N_14482,N_13567,N_13930);
nor U14483 (N_14483,N_13587,N_13925);
and U14484 (N_14484,N_13787,N_13652);
or U14485 (N_14485,N_13632,N_13789);
nor U14486 (N_14486,N_13642,N_13857);
xor U14487 (N_14487,N_13591,N_13569);
nand U14488 (N_14488,N_13870,N_13844);
nor U14489 (N_14489,N_13510,N_13572);
xnor U14490 (N_14490,N_13759,N_13537);
nand U14491 (N_14491,N_13521,N_13512);
nand U14492 (N_14492,N_13752,N_13545);
nor U14493 (N_14493,N_13781,N_13861);
nor U14494 (N_14494,N_13668,N_13862);
or U14495 (N_14495,N_13678,N_13533);
nor U14496 (N_14496,N_13676,N_13738);
nor U14497 (N_14497,N_13802,N_13731);
xnor U14498 (N_14498,N_13977,N_13905);
nand U14499 (N_14499,N_13569,N_13848);
xnor U14500 (N_14500,N_14219,N_14413);
and U14501 (N_14501,N_14152,N_14007);
nand U14502 (N_14502,N_14010,N_14227);
nand U14503 (N_14503,N_14398,N_14352);
nor U14504 (N_14504,N_14367,N_14351);
nand U14505 (N_14505,N_14267,N_14162);
and U14506 (N_14506,N_14478,N_14487);
and U14507 (N_14507,N_14097,N_14276);
nand U14508 (N_14508,N_14042,N_14106);
nor U14509 (N_14509,N_14446,N_14239);
nor U14510 (N_14510,N_14386,N_14279);
and U14511 (N_14511,N_14455,N_14223);
nand U14512 (N_14512,N_14256,N_14077);
or U14513 (N_14513,N_14426,N_14349);
nand U14514 (N_14514,N_14121,N_14308);
or U14515 (N_14515,N_14322,N_14423);
and U14516 (N_14516,N_14115,N_14303);
nand U14517 (N_14517,N_14240,N_14025);
nor U14518 (N_14518,N_14345,N_14110);
or U14519 (N_14519,N_14038,N_14342);
xor U14520 (N_14520,N_14041,N_14058);
or U14521 (N_14521,N_14376,N_14022);
nand U14522 (N_14522,N_14436,N_14033);
nor U14523 (N_14523,N_14287,N_14245);
xnor U14524 (N_14524,N_14216,N_14408);
nor U14525 (N_14525,N_14036,N_14159);
nand U14526 (N_14526,N_14183,N_14312);
xor U14527 (N_14527,N_14283,N_14289);
or U14528 (N_14528,N_14052,N_14315);
xor U14529 (N_14529,N_14250,N_14450);
or U14530 (N_14530,N_14374,N_14141);
and U14531 (N_14531,N_14329,N_14059);
nor U14532 (N_14532,N_14390,N_14174);
nand U14533 (N_14533,N_14205,N_14292);
xnor U14534 (N_14534,N_14006,N_14073);
or U14535 (N_14535,N_14440,N_14421);
nand U14536 (N_14536,N_14184,N_14405);
or U14537 (N_14537,N_14392,N_14473);
nor U14538 (N_14538,N_14338,N_14065);
xnor U14539 (N_14539,N_14112,N_14359);
nand U14540 (N_14540,N_14053,N_14026);
and U14541 (N_14541,N_14075,N_14406);
and U14542 (N_14542,N_14215,N_14282);
nand U14543 (N_14543,N_14043,N_14049);
and U14544 (N_14544,N_14306,N_14062);
and U14545 (N_14545,N_14236,N_14424);
nand U14546 (N_14546,N_14437,N_14400);
or U14547 (N_14547,N_14251,N_14176);
nor U14548 (N_14548,N_14499,N_14275);
and U14549 (N_14549,N_14087,N_14464);
or U14550 (N_14550,N_14381,N_14407);
xnor U14551 (N_14551,N_14410,N_14323);
nor U14552 (N_14552,N_14317,N_14368);
nand U14553 (N_14553,N_14355,N_14101);
and U14554 (N_14554,N_14186,N_14116);
or U14555 (N_14555,N_14493,N_14199);
nor U14556 (N_14556,N_14401,N_14365);
nand U14557 (N_14557,N_14497,N_14311);
and U14558 (N_14558,N_14163,N_14181);
and U14559 (N_14559,N_14234,N_14459);
xnor U14560 (N_14560,N_14442,N_14462);
nor U14561 (N_14561,N_14238,N_14475);
nand U14562 (N_14562,N_14185,N_14285);
nand U14563 (N_14563,N_14331,N_14425);
nor U14564 (N_14564,N_14182,N_14291);
nand U14565 (N_14565,N_14372,N_14169);
or U14566 (N_14566,N_14258,N_14064);
and U14567 (N_14567,N_14347,N_14108);
or U14568 (N_14568,N_14427,N_14320);
nand U14569 (N_14569,N_14384,N_14123);
xor U14570 (N_14570,N_14265,N_14480);
nor U14571 (N_14571,N_14221,N_14498);
nand U14572 (N_14572,N_14445,N_14090);
xnor U14573 (N_14573,N_14330,N_14235);
xnor U14574 (N_14574,N_14286,N_14277);
xor U14575 (N_14575,N_14158,N_14161);
nor U14576 (N_14576,N_14146,N_14430);
nand U14577 (N_14577,N_14414,N_14003);
xnor U14578 (N_14578,N_14104,N_14492);
xnor U14579 (N_14579,N_14098,N_14363);
and U14580 (N_14580,N_14357,N_14337);
or U14581 (N_14581,N_14435,N_14370);
nor U14582 (N_14582,N_14488,N_14086);
nor U14583 (N_14583,N_14136,N_14203);
nand U14584 (N_14584,N_14242,N_14451);
xor U14585 (N_14585,N_14439,N_14079);
and U14586 (N_14586,N_14024,N_14230);
xnor U14587 (N_14587,N_14210,N_14126);
nor U14588 (N_14588,N_14180,N_14122);
or U14589 (N_14589,N_14485,N_14366);
xnor U14590 (N_14590,N_14102,N_14091);
and U14591 (N_14591,N_14231,N_14128);
or U14592 (N_14592,N_14481,N_14375);
nand U14593 (N_14593,N_14193,N_14188);
nor U14594 (N_14594,N_14070,N_14032);
nand U14595 (N_14595,N_14218,N_14016);
and U14596 (N_14596,N_14081,N_14300);
xor U14597 (N_14597,N_14164,N_14334);
xor U14598 (N_14598,N_14171,N_14200);
and U14599 (N_14599,N_14469,N_14018);
xor U14600 (N_14600,N_14268,N_14226);
or U14601 (N_14601,N_14348,N_14467);
nand U14602 (N_14602,N_14402,N_14155);
and U14603 (N_14603,N_14189,N_14061);
nand U14604 (N_14604,N_14044,N_14160);
and U14605 (N_14605,N_14449,N_14166);
or U14606 (N_14606,N_14132,N_14225);
xnor U14607 (N_14607,N_14325,N_14327);
nand U14608 (N_14608,N_14360,N_14274);
or U14609 (N_14609,N_14380,N_14153);
or U14610 (N_14610,N_14138,N_14432);
nand U14611 (N_14611,N_14220,N_14109);
or U14612 (N_14612,N_14391,N_14371);
and U14613 (N_14613,N_14448,N_14213);
and U14614 (N_14614,N_14000,N_14224);
and U14615 (N_14615,N_14496,N_14177);
nor U14616 (N_14616,N_14297,N_14394);
nand U14617 (N_14617,N_14309,N_14211);
and U14618 (N_14618,N_14027,N_14344);
nand U14619 (N_14619,N_14362,N_14120);
or U14620 (N_14620,N_14461,N_14143);
nand U14621 (N_14621,N_14444,N_14361);
and U14622 (N_14622,N_14054,N_14484);
xnor U14623 (N_14623,N_14422,N_14135);
nor U14624 (N_14624,N_14168,N_14051);
xor U14625 (N_14625,N_14139,N_14008);
xnor U14626 (N_14626,N_14244,N_14100);
xnor U14627 (N_14627,N_14209,N_14257);
xor U14628 (N_14628,N_14278,N_14118);
nand U14629 (N_14629,N_14253,N_14197);
or U14630 (N_14630,N_14261,N_14082);
nor U14631 (N_14631,N_14178,N_14191);
and U14632 (N_14632,N_14411,N_14145);
or U14633 (N_14633,N_14034,N_14310);
or U14634 (N_14634,N_14465,N_14294);
nor U14635 (N_14635,N_14269,N_14456);
nand U14636 (N_14636,N_14030,N_14105);
and U14637 (N_14637,N_14491,N_14068);
nor U14638 (N_14638,N_14170,N_14020);
or U14639 (N_14639,N_14195,N_14284);
and U14640 (N_14640,N_14096,N_14431);
and U14641 (N_14641,N_14117,N_14262);
nand U14642 (N_14642,N_14201,N_14005);
and U14643 (N_14643,N_14085,N_14013);
and U14644 (N_14644,N_14243,N_14364);
or U14645 (N_14645,N_14476,N_14252);
nand U14646 (N_14646,N_14395,N_14165);
and U14647 (N_14647,N_14055,N_14358);
xor U14648 (N_14648,N_14194,N_14388);
xnor U14649 (N_14649,N_14217,N_14202);
xnor U14650 (N_14650,N_14014,N_14125);
or U14651 (N_14651,N_14147,N_14222);
nor U14652 (N_14652,N_14047,N_14468);
xor U14653 (N_14653,N_14254,N_14088);
xnor U14654 (N_14654,N_14314,N_14057);
or U14655 (N_14655,N_14270,N_14264);
xnor U14656 (N_14656,N_14482,N_14346);
nand U14657 (N_14657,N_14490,N_14192);
nand U14658 (N_14658,N_14144,N_14420);
nor U14659 (N_14659,N_14271,N_14137);
xor U14660 (N_14660,N_14343,N_14288);
or U14661 (N_14661,N_14150,N_14389);
xor U14662 (N_14662,N_14304,N_14151);
xor U14663 (N_14663,N_14353,N_14012);
and U14664 (N_14664,N_14273,N_14399);
nand U14665 (N_14665,N_14037,N_14378);
nand U14666 (N_14666,N_14084,N_14318);
nand U14667 (N_14667,N_14204,N_14089);
nor U14668 (N_14668,N_14039,N_14233);
nor U14669 (N_14669,N_14048,N_14483);
and U14670 (N_14670,N_14131,N_14021);
and U14671 (N_14671,N_14272,N_14387);
and U14672 (N_14672,N_14023,N_14035);
or U14673 (N_14673,N_14083,N_14466);
or U14674 (N_14674,N_14248,N_14148);
nor U14675 (N_14675,N_14417,N_14263);
or U14676 (N_14676,N_14298,N_14114);
nor U14677 (N_14677,N_14214,N_14335);
or U14678 (N_14678,N_14232,N_14094);
nor U14679 (N_14679,N_14078,N_14259);
and U14680 (N_14680,N_14056,N_14479);
or U14681 (N_14681,N_14046,N_14129);
xnor U14682 (N_14682,N_14157,N_14393);
nor U14683 (N_14683,N_14433,N_14031);
and U14684 (N_14684,N_14339,N_14281);
or U14685 (N_14685,N_14419,N_14369);
and U14686 (N_14686,N_14472,N_14009);
and U14687 (N_14687,N_14247,N_14196);
nor U14688 (N_14688,N_14293,N_14463);
nor U14689 (N_14689,N_14296,N_14198);
nand U14690 (N_14690,N_14454,N_14187);
nor U14691 (N_14691,N_14332,N_14002);
nand U14692 (N_14692,N_14452,N_14301);
and U14693 (N_14693,N_14237,N_14396);
nand U14694 (N_14694,N_14060,N_14418);
or U14695 (N_14695,N_14477,N_14409);
or U14696 (N_14696,N_14453,N_14127);
nand U14697 (N_14697,N_14447,N_14228);
xor U14698 (N_14698,N_14340,N_14019);
nand U14699 (N_14699,N_14341,N_14076);
xnor U14700 (N_14700,N_14095,N_14212);
or U14701 (N_14701,N_14494,N_14471);
nor U14702 (N_14702,N_14313,N_14099);
nand U14703 (N_14703,N_14474,N_14154);
or U14704 (N_14704,N_14149,N_14072);
and U14705 (N_14705,N_14412,N_14103);
nor U14706 (N_14706,N_14067,N_14004);
and U14707 (N_14707,N_14373,N_14429);
nand U14708 (N_14708,N_14092,N_14190);
xnor U14709 (N_14709,N_14080,N_14460);
and U14710 (N_14710,N_14416,N_14350);
xor U14711 (N_14711,N_14133,N_14167);
and U14712 (N_14712,N_14403,N_14356);
nor U14713 (N_14713,N_14290,N_14260);
nor U14714 (N_14714,N_14207,N_14383);
xnor U14715 (N_14715,N_14011,N_14040);
nor U14716 (N_14716,N_14319,N_14229);
or U14717 (N_14717,N_14124,N_14354);
and U14718 (N_14718,N_14458,N_14074);
xor U14719 (N_14719,N_14324,N_14119);
nand U14720 (N_14720,N_14428,N_14093);
or U14721 (N_14721,N_14107,N_14175);
nor U14722 (N_14722,N_14336,N_14208);
nor U14723 (N_14723,N_14299,N_14489);
xnor U14724 (N_14724,N_14255,N_14066);
and U14725 (N_14725,N_14071,N_14280);
or U14726 (N_14726,N_14495,N_14326);
nor U14727 (N_14727,N_14305,N_14434);
nor U14728 (N_14728,N_14266,N_14302);
or U14729 (N_14729,N_14328,N_14316);
or U14730 (N_14730,N_14050,N_14333);
xor U14731 (N_14731,N_14045,N_14321);
nor U14732 (N_14732,N_14397,N_14069);
xnor U14733 (N_14733,N_14404,N_14111);
nand U14734 (N_14734,N_14246,N_14443);
nor U14735 (N_14735,N_14156,N_14295);
nand U14736 (N_14736,N_14377,N_14206);
nand U14737 (N_14737,N_14441,N_14142);
nor U14738 (N_14738,N_14415,N_14063);
and U14739 (N_14739,N_14172,N_14470);
nor U14740 (N_14740,N_14379,N_14385);
nor U14741 (N_14741,N_14015,N_14173);
xor U14742 (N_14742,N_14028,N_14438);
nor U14743 (N_14743,N_14140,N_14179);
or U14744 (N_14744,N_14241,N_14113);
nor U14745 (N_14745,N_14457,N_14134);
or U14746 (N_14746,N_14029,N_14486);
and U14747 (N_14747,N_14249,N_14017);
xnor U14748 (N_14748,N_14130,N_14307);
or U14749 (N_14749,N_14001,N_14382);
nor U14750 (N_14750,N_14371,N_14205);
nor U14751 (N_14751,N_14281,N_14303);
nor U14752 (N_14752,N_14094,N_14184);
xnor U14753 (N_14753,N_14463,N_14410);
or U14754 (N_14754,N_14221,N_14001);
or U14755 (N_14755,N_14266,N_14323);
xnor U14756 (N_14756,N_14069,N_14042);
nand U14757 (N_14757,N_14322,N_14468);
nor U14758 (N_14758,N_14186,N_14357);
nand U14759 (N_14759,N_14102,N_14235);
xnor U14760 (N_14760,N_14230,N_14081);
nor U14761 (N_14761,N_14134,N_14351);
and U14762 (N_14762,N_14227,N_14452);
nor U14763 (N_14763,N_14072,N_14083);
and U14764 (N_14764,N_14259,N_14043);
or U14765 (N_14765,N_14298,N_14382);
nor U14766 (N_14766,N_14347,N_14110);
or U14767 (N_14767,N_14321,N_14330);
nor U14768 (N_14768,N_14058,N_14232);
or U14769 (N_14769,N_14073,N_14146);
and U14770 (N_14770,N_14448,N_14462);
nor U14771 (N_14771,N_14079,N_14116);
and U14772 (N_14772,N_14282,N_14245);
nand U14773 (N_14773,N_14274,N_14153);
or U14774 (N_14774,N_14274,N_14231);
xnor U14775 (N_14775,N_14256,N_14095);
or U14776 (N_14776,N_14050,N_14470);
nand U14777 (N_14777,N_14151,N_14320);
xnor U14778 (N_14778,N_14274,N_14276);
or U14779 (N_14779,N_14390,N_14013);
nand U14780 (N_14780,N_14192,N_14333);
nor U14781 (N_14781,N_14390,N_14203);
nand U14782 (N_14782,N_14363,N_14143);
and U14783 (N_14783,N_14432,N_14372);
nand U14784 (N_14784,N_14126,N_14021);
or U14785 (N_14785,N_14248,N_14019);
nand U14786 (N_14786,N_14212,N_14101);
xor U14787 (N_14787,N_14044,N_14188);
and U14788 (N_14788,N_14252,N_14007);
nand U14789 (N_14789,N_14043,N_14409);
nand U14790 (N_14790,N_14056,N_14197);
xor U14791 (N_14791,N_14234,N_14400);
nand U14792 (N_14792,N_14039,N_14188);
xor U14793 (N_14793,N_14223,N_14212);
and U14794 (N_14794,N_14073,N_14132);
and U14795 (N_14795,N_14390,N_14339);
nand U14796 (N_14796,N_14057,N_14116);
nor U14797 (N_14797,N_14231,N_14366);
or U14798 (N_14798,N_14239,N_14031);
nor U14799 (N_14799,N_14170,N_14369);
or U14800 (N_14800,N_14006,N_14451);
nand U14801 (N_14801,N_14063,N_14480);
nand U14802 (N_14802,N_14225,N_14271);
nor U14803 (N_14803,N_14201,N_14461);
nand U14804 (N_14804,N_14201,N_14323);
or U14805 (N_14805,N_14241,N_14234);
nand U14806 (N_14806,N_14191,N_14172);
and U14807 (N_14807,N_14492,N_14273);
or U14808 (N_14808,N_14246,N_14277);
xor U14809 (N_14809,N_14371,N_14326);
or U14810 (N_14810,N_14013,N_14053);
or U14811 (N_14811,N_14498,N_14075);
nand U14812 (N_14812,N_14008,N_14359);
and U14813 (N_14813,N_14113,N_14314);
nor U14814 (N_14814,N_14030,N_14356);
nand U14815 (N_14815,N_14269,N_14230);
xnor U14816 (N_14816,N_14154,N_14236);
or U14817 (N_14817,N_14262,N_14409);
or U14818 (N_14818,N_14373,N_14300);
nor U14819 (N_14819,N_14381,N_14409);
nor U14820 (N_14820,N_14190,N_14238);
or U14821 (N_14821,N_14368,N_14384);
nand U14822 (N_14822,N_14199,N_14394);
and U14823 (N_14823,N_14348,N_14103);
xnor U14824 (N_14824,N_14374,N_14353);
xor U14825 (N_14825,N_14075,N_14490);
nand U14826 (N_14826,N_14407,N_14305);
nor U14827 (N_14827,N_14153,N_14394);
or U14828 (N_14828,N_14424,N_14290);
or U14829 (N_14829,N_14324,N_14441);
and U14830 (N_14830,N_14331,N_14197);
xor U14831 (N_14831,N_14362,N_14415);
nor U14832 (N_14832,N_14445,N_14421);
and U14833 (N_14833,N_14088,N_14167);
nand U14834 (N_14834,N_14303,N_14480);
xor U14835 (N_14835,N_14077,N_14205);
nor U14836 (N_14836,N_14299,N_14127);
nor U14837 (N_14837,N_14267,N_14404);
and U14838 (N_14838,N_14413,N_14137);
nor U14839 (N_14839,N_14046,N_14355);
or U14840 (N_14840,N_14219,N_14167);
or U14841 (N_14841,N_14498,N_14015);
xnor U14842 (N_14842,N_14018,N_14295);
nand U14843 (N_14843,N_14052,N_14441);
nor U14844 (N_14844,N_14019,N_14200);
and U14845 (N_14845,N_14400,N_14444);
xnor U14846 (N_14846,N_14263,N_14306);
and U14847 (N_14847,N_14313,N_14020);
nand U14848 (N_14848,N_14423,N_14165);
xnor U14849 (N_14849,N_14059,N_14084);
or U14850 (N_14850,N_14391,N_14489);
and U14851 (N_14851,N_14286,N_14368);
nor U14852 (N_14852,N_14377,N_14379);
or U14853 (N_14853,N_14190,N_14076);
nor U14854 (N_14854,N_14034,N_14427);
or U14855 (N_14855,N_14098,N_14200);
and U14856 (N_14856,N_14343,N_14222);
nor U14857 (N_14857,N_14075,N_14473);
nand U14858 (N_14858,N_14220,N_14332);
nand U14859 (N_14859,N_14068,N_14186);
nor U14860 (N_14860,N_14230,N_14316);
nor U14861 (N_14861,N_14031,N_14414);
nor U14862 (N_14862,N_14182,N_14321);
or U14863 (N_14863,N_14334,N_14131);
and U14864 (N_14864,N_14263,N_14255);
nand U14865 (N_14865,N_14263,N_14400);
or U14866 (N_14866,N_14187,N_14180);
nand U14867 (N_14867,N_14381,N_14295);
and U14868 (N_14868,N_14387,N_14217);
and U14869 (N_14869,N_14350,N_14051);
or U14870 (N_14870,N_14190,N_14334);
nor U14871 (N_14871,N_14045,N_14370);
and U14872 (N_14872,N_14262,N_14124);
or U14873 (N_14873,N_14256,N_14007);
xnor U14874 (N_14874,N_14435,N_14408);
and U14875 (N_14875,N_14130,N_14455);
xor U14876 (N_14876,N_14454,N_14427);
and U14877 (N_14877,N_14344,N_14346);
nand U14878 (N_14878,N_14152,N_14044);
xor U14879 (N_14879,N_14233,N_14291);
nand U14880 (N_14880,N_14078,N_14003);
xor U14881 (N_14881,N_14493,N_14342);
and U14882 (N_14882,N_14337,N_14153);
nand U14883 (N_14883,N_14362,N_14458);
and U14884 (N_14884,N_14443,N_14352);
nand U14885 (N_14885,N_14351,N_14099);
and U14886 (N_14886,N_14192,N_14393);
and U14887 (N_14887,N_14307,N_14386);
or U14888 (N_14888,N_14085,N_14098);
nor U14889 (N_14889,N_14371,N_14182);
nor U14890 (N_14890,N_14279,N_14093);
nand U14891 (N_14891,N_14199,N_14405);
or U14892 (N_14892,N_14086,N_14455);
or U14893 (N_14893,N_14176,N_14046);
or U14894 (N_14894,N_14115,N_14341);
nand U14895 (N_14895,N_14184,N_14306);
xor U14896 (N_14896,N_14007,N_14132);
and U14897 (N_14897,N_14336,N_14215);
nand U14898 (N_14898,N_14139,N_14054);
xnor U14899 (N_14899,N_14333,N_14290);
and U14900 (N_14900,N_14107,N_14282);
nand U14901 (N_14901,N_14178,N_14377);
nand U14902 (N_14902,N_14094,N_14433);
nand U14903 (N_14903,N_14340,N_14425);
nand U14904 (N_14904,N_14146,N_14110);
and U14905 (N_14905,N_14484,N_14373);
or U14906 (N_14906,N_14341,N_14349);
nand U14907 (N_14907,N_14293,N_14211);
or U14908 (N_14908,N_14119,N_14118);
or U14909 (N_14909,N_14071,N_14375);
or U14910 (N_14910,N_14448,N_14465);
or U14911 (N_14911,N_14124,N_14434);
nand U14912 (N_14912,N_14386,N_14086);
and U14913 (N_14913,N_14103,N_14440);
nor U14914 (N_14914,N_14321,N_14445);
nand U14915 (N_14915,N_14309,N_14494);
or U14916 (N_14916,N_14337,N_14328);
and U14917 (N_14917,N_14291,N_14049);
xor U14918 (N_14918,N_14469,N_14359);
nand U14919 (N_14919,N_14018,N_14412);
nand U14920 (N_14920,N_14164,N_14441);
nor U14921 (N_14921,N_14309,N_14117);
and U14922 (N_14922,N_14011,N_14426);
xor U14923 (N_14923,N_14107,N_14399);
nor U14924 (N_14924,N_14086,N_14096);
xor U14925 (N_14925,N_14379,N_14346);
xnor U14926 (N_14926,N_14316,N_14130);
and U14927 (N_14927,N_14268,N_14404);
xnor U14928 (N_14928,N_14439,N_14060);
or U14929 (N_14929,N_14260,N_14491);
or U14930 (N_14930,N_14308,N_14023);
nor U14931 (N_14931,N_14228,N_14411);
and U14932 (N_14932,N_14404,N_14340);
nor U14933 (N_14933,N_14483,N_14249);
nand U14934 (N_14934,N_14312,N_14235);
and U14935 (N_14935,N_14349,N_14324);
nand U14936 (N_14936,N_14381,N_14092);
or U14937 (N_14937,N_14361,N_14307);
nor U14938 (N_14938,N_14066,N_14347);
nand U14939 (N_14939,N_14088,N_14272);
xor U14940 (N_14940,N_14142,N_14235);
and U14941 (N_14941,N_14435,N_14299);
nor U14942 (N_14942,N_14365,N_14415);
nor U14943 (N_14943,N_14281,N_14227);
or U14944 (N_14944,N_14037,N_14466);
xor U14945 (N_14945,N_14122,N_14155);
nand U14946 (N_14946,N_14220,N_14170);
nand U14947 (N_14947,N_14359,N_14085);
and U14948 (N_14948,N_14212,N_14199);
nor U14949 (N_14949,N_14227,N_14166);
and U14950 (N_14950,N_14274,N_14230);
xor U14951 (N_14951,N_14072,N_14006);
xor U14952 (N_14952,N_14130,N_14045);
and U14953 (N_14953,N_14223,N_14460);
nand U14954 (N_14954,N_14314,N_14465);
nand U14955 (N_14955,N_14292,N_14044);
nand U14956 (N_14956,N_14247,N_14268);
and U14957 (N_14957,N_14315,N_14110);
nor U14958 (N_14958,N_14424,N_14353);
xor U14959 (N_14959,N_14257,N_14444);
and U14960 (N_14960,N_14169,N_14196);
nand U14961 (N_14961,N_14047,N_14280);
and U14962 (N_14962,N_14369,N_14473);
nor U14963 (N_14963,N_14478,N_14167);
xor U14964 (N_14964,N_14128,N_14224);
nor U14965 (N_14965,N_14488,N_14139);
nand U14966 (N_14966,N_14295,N_14299);
or U14967 (N_14967,N_14314,N_14160);
nor U14968 (N_14968,N_14260,N_14452);
and U14969 (N_14969,N_14275,N_14343);
nand U14970 (N_14970,N_14287,N_14332);
nand U14971 (N_14971,N_14035,N_14043);
xor U14972 (N_14972,N_14160,N_14396);
xor U14973 (N_14973,N_14305,N_14145);
nor U14974 (N_14974,N_14416,N_14133);
nor U14975 (N_14975,N_14459,N_14260);
or U14976 (N_14976,N_14460,N_14288);
nand U14977 (N_14977,N_14056,N_14372);
or U14978 (N_14978,N_14227,N_14111);
and U14979 (N_14979,N_14250,N_14417);
or U14980 (N_14980,N_14128,N_14006);
nand U14981 (N_14981,N_14328,N_14321);
nand U14982 (N_14982,N_14158,N_14153);
nand U14983 (N_14983,N_14200,N_14065);
nand U14984 (N_14984,N_14385,N_14299);
nand U14985 (N_14985,N_14206,N_14279);
nand U14986 (N_14986,N_14368,N_14038);
and U14987 (N_14987,N_14133,N_14006);
or U14988 (N_14988,N_14392,N_14378);
nand U14989 (N_14989,N_14136,N_14096);
xor U14990 (N_14990,N_14277,N_14442);
nor U14991 (N_14991,N_14442,N_14182);
and U14992 (N_14992,N_14499,N_14430);
or U14993 (N_14993,N_14498,N_14367);
nor U14994 (N_14994,N_14359,N_14366);
nand U14995 (N_14995,N_14210,N_14114);
nand U14996 (N_14996,N_14348,N_14025);
xor U14997 (N_14997,N_14381,N_14137);
xnor U14998 (N_14998,N_14137,N_14189);
nor U14999 (N_14999,N_14243,N_14415);
and U15000 (N_15000,N_14819,N_14817);
or U15001 (N_15001,N_14650,N_14839);
nor U15002 (N_15002,N_14659,N_14837);
xnor U15003 (N_15003,N_14713,N_14940);
and U15004 (N_15004,N_14739,N_14956);
nand U15005 (N_15005,N_14561,N_14647);
nand U15006 (N_15006,N_14676,N_14971);
xnor U15007 (N_15007,N_14637,N_14820);
or U15008 (N_15008,N_14856,N_14943);
and U15009 (N_15009,N_14830,N_14951);
or U15010 (N_15010,N_14807,N_14795);
or U15011 (N_15011,N_14576,N_14513);
xnor U15012 (N_15012,N_14707,N_14536);
or U15013 (N_15013,N_14598,N_14564);
nand U15014 (N_15014,N_14551,N_14841);
xnor U15015 (N_15015,N_14597,N_14699);
nand U15016 (N_15016,N_14808,N_14733);
or U15017 (N_15017,N_14648,N_14555);
nand U15018 (N_15018,N_14779,N_14579);
nor U15019 (N_15019,N_14588,N_14913);
nor U15020 (N_15020,N_14821,N_14757);
and U15021 (N_15021,N_14912,N_14553);
or U15022 (N_15022,N_14935,N_14881);
or U15023 (N_15023,N_14906,N_14697);
nor U15024 (N_15024,N_14734,N_14514);
xor U15025 (N_15025,N_14575,N_14934);
or U15026 (N_15026,N_14919,N_14716);
and U15027 (N_15027,N_14642,N_14688);
or U15028 (N_15028,N_14785,N_14723);
nor U15029 (N_15029,N_14886,N_14952);
or U15030 (N_15030,N_14986,N_14784);
and U15031 (N_15031,N_14834,N_14567);
nand U15032 (N_15032,N_14946,N_14915);
nor U15033 (N_15033,N_14735,N_14759);
xnor U15034 (N_15034,N_14968,N_14849);
and U15035 (N_15035,N_14869,N_14931);
and U15036 (N_15036,N_14972,N_14780);
nand U15037 (N_15037,N_14996,N_14570);
nand U15038 (N_15038,N_14541,N_14655);
and U15039 (N_15039,N_14621,N_14964);
nor U15040 (N_15040,N_14873,N_14674);
xor U15041 (N_15041,N_14715,N_14857);
nand U15042 (N_15042,N_14954,N_14748);
nand U15043 (N_15043,N_14680,N_14771);
and U15044 (N_15044,N_14772,N_14937);
or U15045 (N_15045,N_14522,N_14884);
nor U15046 (N_15046,N_14770,N_14617);
xor U15047 (N_15047,N_14920,N_14847);
nand U15048 (N_15048,N_14833,N_14526);
nor U15049 (N_15049,N_14994,N_14646);
nor U15050 (N_15050,N_14590,N_14731);
and U15051 (N_15051,N_14503,N_14634);
and U15052 (N_15052,N_14711,N_14729);
nor U15053 (N_15053,N_14801,N_14933);
and U15054 (N_15054,N_14622,N_14975);
xnor U15055 (N_15055,N_14753,N_14623);
nor U15056 (N_15056,N_14815,N_14721);
and U15057 (N_15057,N_14596,N_14507);
nand U15058 (N_15058,N_14727,N_14704);
nand U15059 (N_15059,N_14649,N_14864);
nand U15060 (N_15060,N_14569,N_14880);
and U15061 (N_15061,N_14632,N_14897);
nor U15062 (N_15062,N_14624,N_14700);
nand U15063 (N_15063,N_14749,N_14504);
nor U15064 (N_15064,N_14929,N_14728);
xnor U15065 (N_15065,N_14792,N_14629);
nor U15066 (N_15066,N_14928,N_14947);
or U15067 (N_15067,N_14515,N_14987);
nand U15068 (N_15068,N_14627,N_14828);
nor U15069 (N_15069,N_14584,N_14610);
xnor U15070 (N_15070,N_14794,N_14605);
or U15071 (N_15071,N_14898,N_14983);
or U15072 (N_15072,N_14914,N_14538);
or U15073 (N_15073,N_14595,N_14562);
nor U15074 (N_15074,N_14651,N_14774);
nor U15075 (N_15075,N_14766,N_14525);
and U15076 (N_15076,N_14822,N_14978);
and U15077 (N_15077,N_14568,N_14630);
xnor U15078 (N_15078,N_14758,N_14741);
nand U15079 (N_15079,N_14549,N_14944);
xor U15080 (N_15080,N_14916,N_14517);
or U15081 (N_15081,N_14652,N_14903);
nand U15082 (N_15082,N_14980,N_14950);
nand U15083 (N_15083,N_14922,N_14997);
nor U15084 (N_15084,N_14532,N_14752);
nor U15085 (N_15085,N_14602,N_14730);
and U15086 (N_15086,N_14874,N_14530);
nor U15087 (N_15087,N_14861,N_14683);
or U15088 (N_15088,N_14668,N_14671);
nor U15089 (N_15089,N_14523,N_14520);
nand U15090 (N_15090,N_14667,N_14724);
nand U15091 (N_15091,N_14781,N_14710);
nor U15092 (N_15092,N_14738,N_14835);
nand U15093 (N_15093,N_14974,N_14967);
xnor U15094 (N_15094,N_14926,N_14742);
xor U15095 (N_15095,N_14509,N_14677);
nand U15096 (N_15096,N_14945,N_14554);
nand U15097 (N_15097,N_14638,N_14628);
nand U15098 (N_15098,N_14641,N_14587);
nor U15099 (N_15099,N_14670,N_14959);
xor U15100 (N_15100,N_14559,N_14706);
and U15101 (N_15101,N_14802,N_14572);
or U15102 (N_15102,N_14705,N_14583);
nor U15103 (N_15103,N_14566,N_14644);
nand U15104 (N_15104,N_14692,N_14941);
nand U15105 (N_15105,N_14533,N_14556);
nor U15106 (N_15106,N_14798,N_14661);
and U15107 (N_15107,N_14720,N_14838);
or U15108 (N_15108,N_14672,N_14613);
xor U15109 (N_15109,N_14768,N_14845);
xnor U15110 (N_15110,N_14918,N_14546);
nor U15111 (N_15111,N_14603,N_14854);
nor U15112 (N_15112,N_14998,N_14501);
nand U15113 (N_15113,N_14901,N_14803);
nor U15114 (N_15114,N_14850,N_14657);
xor U15115 (N_15115,N_14879,N_14611);
and U15116 (N_15116,N_14889,N_14899);
xor U15117 (N_15117,N_14656,N_14762);
xor U15118 (N_15118,N_14930,N_14805);
or U15119 (N_15119,N_14535,N_14865);
nand U15120 (N_15120,N_14534,N_14842);
xnor U15121 (N_15121,N_14979,N_14718);
or U15122 (N_15122,N_14925,N_14927);
xnor U15123 (N_15123,N_14890,N_14577);
and U15124 (N_15124,N_14949,N_14722);
nand U15125 (N_15125,N_14851,N_14965);
xnor U15126 (N_15126,N_14574,N_14563);
and U15127 (N_15127,N_14558,N_14958);
or U15128 (N_15128,N_14957,N_14982);
nor U15129 (N_15129,N_14740,N_14776);
and U15130 (N_15130,N_14750,N_14924);
and U15131 (N_15131,N_14814,N_14764);
and U15132 (N_15132,N_14591,N_14846);
and U15133 (N_15133,N_14778,N_14787);
xor U15134 (N_15134,N_14663,N_14895);
or U15135 (N_15135,N_14519,N_14592);
xor U15136 (N_15136,N_14548,N_14678);
or U15137 (N_15137,N_14528,N_14755);
xor U15138 (N_15138,N_14995,N_14545);
xor U15139 (N_15139,N_14988,N_14827);
nor U15140 (N_15140,N_14858,N_14521);
or U15141 (N_15141,N_14760,N_14712);
or U15142 (N_15142,N_14581,N_14862);
nand U15143 (N_15143,N_14518,N_14806);
xnor U15144 (N_15144,N_14589,N_14686);
xor U15145 (N_15145,N_14506,N_14654);
xnor U15146 (N_15146,N_14769,N_14761);
nor U15147 (N_15147,N_14500,N_14608);
and U15148 (N_15148,N_14550,N_14796);
nand U15149 (N_15149,N_14527,N_14799);
xnor U15150 (N_15150,N_14786,N_14543);
nor U15151 (N_15151,N_14664,N_14948);
or U15152 (N_15152,N_14868,N_14844);
and U15153 (N_15153,N_14639,N_14653);
nor U15154 (N_15154,N_14557,N_14614);
and U15155 (N_15155,N_14618,N_14658);
and U15156 (N_15156,N_14875,N_14963);
nor U15157 (N_15157,N_14904,N_14871);
or U15158 (N_15158,N_14747,N_14900);
nor U15159 (N_15159,N_14966,N_14836);
nand U15160 (N_15160,N_14932,N_14696);
and U15161 (N_15161,N_14810,N_14872);
nand U15162 (N_15162,N_14985,N_14882);
and U15163 (N_15163,N_14910,N_14573);
nor U15164 (N_15164,N_14981,N_14607);
or U15165 (N_15165,N_14660,N_14789);
nor U15166 (N_15166,N_14703,N_14942);
and U15167 (N_15167,N_14508,N_14682);
xor U15168 (N_15168,N_14537,N_14812);
xnor U15169 (N_15169,N_14960,N_14679);
and U15170 (N_15170,N_14775,N_14560);
xnor U15171 (N_15171,N_14896,N_14600);
and U15172 (N_15172,N_14529,N_14708);
and U15173 (N_15173,N_14831,N_14593);
nand U15174 (N_15174,N_14826,N_14698);
nor U15175 (N_15175,N_14989,N_14685);
xnor U15176 (N_15176,N_14811,N_14797);
nor U15177 (N_15177,N_14876,N_14921);
and U15178 (N_15178,N_14645,N_14917);
nand U15179 (N_15179,N_14909,N_14544);
nand U15180 (N_15180,N_14961,N_14505);
xor U15181 (N_15181,N_14691,N_14743);
xnor U15182 (N_15182,N_14684,N_14791);
xor U15183 (N_15183,N_14782,N_14962);
nand U15184 (N_15184,N_14687,N_14636);
and U15185 (N_15185,N_14832,N_14976);
and U15186 (N_15186,N_14745,N_14620);
nand U15187 (N_15187,N_14823,N_14955);
or U15188 (N_15188,N_14580,N_14892);
xor U15189 (N_15189,N_14977,N_14907);
or U15190 (N_15190,N_14829,N_14969);
xor U15191 (N_15191,N_14582,N_14777);
or U15192 (N_15192,N_14726,N_14973);
or U15193 (N_15193,N_14984,N_14571);
xnor U15194 (N_15194,N_14908,N_14665);
xor U15195 (N_15195,N_14790,N_14751);
nand U15196 (N_15196,N_14824,N_14626);
xnor U15197 (N_15197,N_14631,N_14552);
and U15198 (N_15198,N_14640,N_14578);
and U15199 (N_15199,N_14788,N_14662);
nor U15200 (N_15200,N_14695,N_14719);
xor U15201 (N_15201,N_14635,N_14891);
or U15202 (N_15202,N_14714,N_14689);
nand U15203 (N_15203,N_14599,N_14502);
and U15204 (N_15204,N_14804,N_14601);
and U15205 (N_15205,N_14725,N_14606);
nor U15206 (N_15206,N_14911,N_14547);
nand U15207 (N_15207,N_14970,N_14609);
or U15208 (N_15208,N_14863,N_14717);
nor U15209 (N_15209,N_14887,N_14666);
or U15210 (N_15210,N_14754,N_14859);
nor U15211 (N_15211,N_14840,N_14643);
or U15212 (N_15212,N_14746,N_14512);
and U15213 (N_15213,N_14866,N_14673);
nor U15214 (N_15214,N_14737,N_14690);
or U15215 (N_15215,N_14936,N_14702);
or U15216 (N_15216,N_14999,N_14883);
nand U15217 (N_15217,N_14885,N_14539);
and U15218 (N_15218,N_14736,N_14675);
xnor U15219 (N_15219,N_14693,N_14992);
xnor U15220 (N_15220,N_14867,N_14585);
nor U15221 (N_15221,N_14767,N_14604);
xor U15222 (N_15222,N_14783,N_14991);
nor U15223 (N_15223,N_14870,N_14809);
nand U15224 (N_15224,N_14701,N_14793);
xnor U15225 (N_15225,N_14516,N_14616);
and U15226 (N_15226,N_14825,N_14939);
and U15227 (N_15227,N_14905,N_14902);
nand U15228 (N_15228,N_14732,N_14888);
nor U15229 (N_15229,N_14615,N_14853);
xor U15230 (N_15230,N_14531,N_14524);
nand U15231 (N_15231,N_14894,N_14800);
nand U15232 (N_15232,N_14669,N_14540);
nor U15233 (N_15233,N_14855,N_14511);
xor U15234 (N_15234,N_14993,N_14586);
and U15235 (N_15235,N_14542,N_14756);
or U15236 (N_15236,N_14877,N_14612);
or U15237 (N_15237,N_14625,N_14765);
nor U15238 (N_15238,N_14744,N_14878);
xor U15239 (N_15239,N_14565,N_14923);
and U15240 (N_15240,N_14990,N_14818);
xor U15241 (N_15241,N_14848,N_14816);
nand U15242 (N_15242,N_14510,N_14938);
or U15243 (N_15243,N_14953,N_14813);
or U15244 (N_15244,N_14893,N_14852);
xor U15245 (N_15245,N_14843,N_14694);
nand U15246 (N_15246,N_14860,N_14619);
nor U15247 (N_15247,N_14709,N_14773);
or U15248 (N_15248,N_14763,N_14681);
and U15249 (N_15249,N_14594,N_14633);
nand U15250 (N_15250,N_14919,N_14812);
nand U15251 (N_15251,N_14735,N_14663);
xor U15252 (N_15252,N_14802,N_14974);
or U15253 (N_15253,N_14745,N_14774);
and U15254 (N_15254,N_14691,N_14523);
nor U15255 (N_15255,N_14627,N_14941);
nand U15256 (N_15256,N_14655,N_14634);
xor U15257 (N_15257,N_14947,N_14643);
nor U15258 (N_15258,N_14793,N_14611);
xnor U15259 (N_15259,N_14588,N_14566);
nor U15260 (N_15260,N_14863,N_14670);
and U15261 (N_15261,N_14685,N_14548);
and U15262 (N_15262,N_14673,N_14692);
and U15263 (N_15263,N_14651,N_14950);
and U15264 (N_15264,N_14742,N_14512);
nand U15265 (N_15265,N_14543,N_14793);
and U15266 (N_15266,N_14754,N_14548);
or U15267 (N_15267,N_14894,N_14865);
nor U15268 (N_15268,N_14766,N_14767);
or U15269 (N_15269,N_14887,N_14703);
nor U15270 (N_15270,N_14937,N_14548);
xor U15271 (N_15271,N_14818,N_14560);
nand U15272 (N_15272,N_14715,N_14528);
nor U15273 (N_15273,N_14939,N_14787);
and U15274 (N_15274,N_14672,N_14920);
nand U15275 (N_15275,N_14845,N_14799);
nor U15276 (N_15276,N_14627,N_14995);
nor U15277 (N_15277,N_14641,N_14621);
nor U15278 (N_15278,N_14605,N_14513);
or U15279 (N_15279,N_14683,N_14618);
and U15280 (N_15280,N_14523,N_14604);
xnor U15281 (N_15281,N_14792,N_14787);
or U15282 (N_15282,N_14637,N_14869);
nand U15283 (N_15283,N_14835,N_14943);
xor U15284 (N_15284,N_14604,N_14913);
xor U15285 (N_15285,N_14902,N_14921);
xnor U15286 (N_15286,N_14989,N_14753);
nand U15287 (N_15287,N_14508,N_14543);
nor U15288 (N_15288,N_14806,N_14924);
nand U15289 (N_15289,N_14697,N_14754);
or U15290 (N_15290,N_14961,N_14525);
xor U15291 (N_15291,N_14904,N_14932);
xnor U15292 (N_15292,N_14511,N_14935);
or U15293 (N_15293,N_14637,N_14501);
and U15294 (N_15294,N_14575,N_14592);
and U15295 (N_15295,N_14951,N_14765);
nor U15296 (N_15296,N_14846,N_14782);
and U15297 (N_15297,N_14885,N_14860);
nand U15298 (N_15298,N_14789,N_14790);
or U15299 (N_15299,N_14521,N_14834);
xnor U15300 (N_15300,N_14916,N_14793);
nor U15301 (N_15301,N_14815,N_14679);
and U15302 (N_15302,N_14974,N_14980);
xnor U15303 (N_15303,N_14734,N_14923);
and U15304 (N_15304,N_14739,N_14537);
nand U15305 (N_15305,N_14889,N_14940);
nor U15306 (N_15306,N_14811,N_14529);
nor U15307 (N_15307,N_14609,N_14992);
and U15308 (N_15308,N_14557,N_14940);
nand U15309 (N_15309,N_14801,N_14929);
and U15310 (N_15310,N_14904,N_14740);
or U15311 (N_15311,N_14850,N_14516);
nand U15312 (N_15312,N_14571,N_14981);
nor U15313 (N_15313,N_14990,N_14599);
nor U15314 (N_15314,N_14751,N_14542);
and U15315 (N_15315,N_14673,N_14650);
nand U15316 (N_15316,N_14856,N_14724);
or U15317 (N_15317,N_14834,N_14517);
xnor U15318 (N_15318,N_14805,N_14799);
or U15319 (N_15319,N_14535,N_14621);
nand U15320 (N_15320,N_14756,N_14560);
nand U15321 (N_15321,N_14829,N_14559);
or U15322 (N_15322,N_14642,N_14833);
nand U15323 (N_15323,N_14761,N_14533);
xor U15324 (N_15324,N_14524,N_14530);
or U15325 (N_15325,N_14899,N_14701);
and U15326 (N_15326,N_14533,N_14882);
nor U15327 (N_15327,N_14581,N_14709);
xnor U15328 (N_15328,N_14591,N_14726);
nor U15329 (N_15329,N_14930,N_14989);
and U15330 (N_15330,N_14786,N_14778);
and U15331 (N_15331,N_14605,N_14664);
or U15332 (N_15332,N_14517,N_14595);
xnor U15333 (N_15333,N_14788,N_14950);
nand U15334 (N_15334,N_14550,N_14765);
nand U15335 (N_15335,N_14674,N_14937);
and U15336 (N_15336,N_14505,N_14658);
nor U15337 (N_15337,N_14985,N_14876);
and U15338 (N_15338,N_14832,N_14837);
or U15339 (N_15339,N_14743,N_14517);
xor U15340 (N_15340,N_14739,N_14538);
and U15341 (N_15341,N_14940,N_14737);
nand U15342 (N_15342,N_14884,N_14731);
nand U15343 (N_15343,N_14564,N_14845);
xor U15344 (N_15344,N_14606,N_14896);
or U15345 (N_15345,N_14579,N_14894);
or U15346 (N_15346,N_14707,N_14844);
or U15347 (N_15347,N_14894,N_14738);
nor U15348 (N_15348,N_14594,N_14788);
and U15349 (N_15349,N_14713,N_14811);
and U15350 (N_15350,N_14832,N_14944);
nand U15351 (N_15351,N_14647,N_14736);
xor U15352 (N_15352,N_14960,N_14604);
and U15353 (N_15353,N_14830,N_14538);
nor U15354 (N_15354,N_14986,N_14787);
nand U15355 (N_15355,N_14950,N_14779);
nor U15356 (N_15356,N_14704,N_14923);
nand U15357 (N_15357,N_14977,N_14647);
nand U15358 (N_15358,N_14956,N_14675);
xor U15359 (N_15359,N_14950,N_14813);
xnor U15360 (N_15360,N_14565,N_14888);
xnor U15361 (N_15361,N_14909,N_14795);
nor U15362 (N_15362,N_14664,N_14881);
nand U15363 (N_15363,N_14735,N_14678);
and U15364 (N_15364,N_14707,N_14566);
nand U15365 (N_15365,N_14668,N_14543);
nor U15366 (N_15366,N_14541,N_14849);
or U15367 (N_15367,N_14652,N_14785);
nand U15368 (N_15368,N_14749,N_14925);
nand U15369 (N_15369,N_14659,N_14839);
xnor U15370 (N_15370,N_14806,N_14792);
xnor U15371 (N_15371,N_14906,N_14552);
and U15372 (N_15372,N_14862,N_14726);
nor U15373 (N_15373,N_14985,N_14989);
and U15374 (N_15374,N_14631,N_14869);
or U15375 (N_15375,N_14572,N_14942);
or U15376 (N_15376,N_14765,N_14574);
nand U15377 (N_15377,N_14730,N_14956);
nor U15378 (N_15378,N_14676,N_14564);
nor U15379 (N_15379,N_14569,N_14565);
and U15380 (N_15380,N_14505,N_14521);
and U15381 (N_15381,N_14738,N_14503);
xor U15382 (N_15382,N_14868,N_14688);
nor U15383 (N_15383,N_14557,N_14511);
nand U15384 (N_15384,N_14993,N_14885);
nor U15385 (N_15385,N_14692,N_14851);
nor U15386 (N_15386,N_14813,N_14908);
or U15387 (N_15387,N_14864,N_14543);
nor U15388 (N_15388,N_14848,N_14650);
or U15389 (N_15389,N_14520,N_14777);
and U15390 (N_15390,N_14583,N_14843);
xnor U15391 (N_15391,N_14711,N_14762);
nand U15392 (N_15392,N_14585,N_14800);
or U15393 (N_15393,N_14972,N_14631);
or U15394 (N_15394,N_14656,N_14640);
nand U15395 (N_15395,N_14690,N_14796);
nor U15396 (N_15396,N_14707,N_14652);
nor U15397 (N_15397,N_14771,N_14627);
xor U15398 (N_15398,N_14713,N_14967);
or U15399 (N_15399,N_14647,N_14966);
or U15400 (N_15400,N_14941,N_14783);
and U15401 (N_15401,N_14715,N_14818);
nand U15402 (N_15402,N_14854,N_14908);
or U15403 (N_15403,N_14628,N_14676);
nor U15404 (N_15404,N_14698,N_14569);
nor U15405 (N_15405,N_14950,N_14530);
nor U15406 (N_15406,N_14822,N_14901);
and U15407 (N_15407,N_14541,N_14790);
xnor U15408 (N_15408,N_14552,N_14918);
nor U15409 (N_15409,N_14538,N_14782);
nor U15410 (N_15410,N_14701,N_14951);
nand U15411 (N_15411,N_14936,N_14520);
and U15412 (N_15412,N_14774,N_14870);
and U15413 (N_15413,N_14552,N_14927);
nor U15414 (N_15414,N_14951,N_14630);
and U15415 (N_15415,N_14827,N_14781);
xor U15416 (N_15416,N_14561,N_14671);
xor U15417 (N_15417,N_14580,N_14731);
or U15418 (N_15418,N_14659,N_14685);
nand U15419 (N_15419,N_14782,N_14753);
xor U15420 (N_15420,N_14707,N_14698);
nor U15421 (N_15421,N_14744,N_14963);
or U15422 (N_15422,N_14973,N_14985);
nand U15423 (N_15423,N_14957,N_14541);
xnor U15424 (N_15424,N_14735,N_14969);
or U15425 (N_15425,N_14710,N_14725);
or U15426 (N_15426,N_14933,N_14607);
or U15427 (N_15427,N_14876,N_14974);
xor U15428 (N_15428,N_14697,N_14803);
or U15429 (N_15429,N_14817,N_14717);
nand U15430 (N_15430,N_14916,N_14885);
nand U15431 (N_15431,N_14523,N_14618);
or U15432 (N_15432,N_14958,N_14781);
nand U15433 (N_15433,N_14535,N_14952);
and U15434 (N_15434,N_14835,N_14762);
nor U15435 (N_15435,N_14994,N_14551);
xor U15436 (N_15436,N_14734,N_14875);
or U15437 (N_15437,N_14977,N_14914);
xnor U15438 (N_15438,N_14613,N_14997);
nor U15439 (N_15439,N_14539,N_14827);
nand U15440 (N_15440,N_14877,N_14571);
nor U15441 (N_15441,N_14638,N_14652);
nand U15442 (N_15442,N_14742,N_14788);
nand U15443 (N_15443,N_14531,N_14682);
and U15444 (N_15444,N_14627,N_14940);
nand U15445 (N_15445,N_14633,N_14624);
or U15446 (N_15446,N_14879,N_14567);
and U15447 (N_15447,N_14644,N_14591);
and U15448 (N_15448,N_14557,N_14678);
or U15449 (N_15449,N_14952,N_14892);
nor U15450 (N_15450,N_14759,N_14855);
xor U15451 (N_15451,N_14853,N_14836);
xnor U15452 (N_15452,N_14752,N_14516);
nor U15453 (N_15453,N_14591,N_14952);
nor U15454 (N_15454,N_14942,N_14588);
nand U15455 (N_15455,N_14829,N_14945);
and U15456 (N_15456,N_14658,N_14672);
nand U15457 (N_15457,N_14912,N_14839);
and U15458 (N_15458,N_14946,N_14869);
nor U15459 (N_15459,N_14655,N_14894);
and U15460 (N_15460,N_14915,N_14733);
xor U15461 (N_15461,N_14748,N_14939);
or U15462 (N_15462,N_14856,N_14854);
and U15463 (N_15463,N_14611,N_14593);
and U15464 (N_15464,N_14620,N_14907);
nand U15465 (N_15465,N_14762,N_14596);
or U15466 (N_15466,N_14826,N_14706);
nand U15467 (N_15467,N_14807,N_14710);
nand U15468 (N_15468,N_14765,N_14871);
or U15469 (N_15469,N_14612,N_14869);
or U15470 (N_15470,N_14719,N_14707);
nand U15471 (N_15471,N_14911,N_14858);
xor U15472 (N_15472,N_14603,N_14979);
and U15473 (N_15473,N_14986,N_14611);
and U15474 (N_15474,N_14956,N_14957);
and U15475 (N_15475,N_14654,N_14644);
or U15476 (N_15476,N_14558,N_14831);
or U15477 (N_15477,N_14804,N_14754);
and U15478 (N_15478,N_14685,N_14738);
nor U15479 (N_15479,N_14938,N_14658);
nor U15480 (N_15480,N_14773,N_14760);
and U15481 (N_15481,N_14940,N_14572);
xnor U15482 (N_15482,N_14966,N_14607);
xnor U15483 (N_15483,N_14647,N_14964);
xor U15484 (N_15484,N_14562,N_14572);
nor U15485 (N_15485,N_14721,N_14679);
nor U15486 (N_15486,N_14877,N_14617);
and U15487 (N_15487,N_14847,N_14616);
xor U15488 (N_15488,N_14846,N_14752);
nor U15489 (N_15489,N_14942,N_14534);
nand U15490 (N_15490,N_14751,N_14597);
or U15491 (N_15491,N_14970,N_14735);
and U15492 (N_15492,N_14517,N_14945);
nor U15493 (N_15493,N_14826,N_14781);
nor U15494 (N_15494,N_14555,N_14777);
nor U15495 (N_15495,N_14608,N_14831);
nand U15496 (N_15496,N_14717,N_14503);
nand U15497 (N_15497,N_14891,N_14501);
or U15498 (N_15498,N_14654,N_14563);
and U15499 (N_15499,N_14858,N_14539);
nand U15500 (N_15500,N_15456,N_15361);
or U15501 (N_15501,N_15344,N_15014);
xor U15502 (N_15502,N_15418,N_15234);
and U15503 (N_15503,N_15003,N_15366);
xor U15504 (N_15504,N_15145,N_15296);
nand U15505 (N_15505,N_15368,N_15087);
and U15506 (N_15506,N_15293,N_15462);
or U15507 (N_15507,N_15070,N_15259);
nand U15508 (N_15508,N_15246,N_15480);
xnor U15509 (N_15509,N_15306,N_15044);
or U15510 (N_15510,N_15230,N_15185);
xor U15511 (N_15511,N_15433,N_15400);
nand U15512 (N_15512,N_15080,N_15357);
nand U15513 (N_15513,N_15432,N_15143);
nand U15514 (N_15514,N_15267,N_15369);
nand U15515 (N_15515,N_15364,N_15325);
and U15516 (N_15516,N_15064,N_15046);
and U15517 (N_15517,N_15022,N_15386);
nand U15518 (N_15518,N_15341,N_15180);
and U15519 (N_15519,N_15297,N_15471);
and U15520 (N_15520,N_15194,N_15453);
nor U15521 (N_15521,N_15193,N_15485);
xnor U15522 (N_15522,N_15329,N_15437);
xnor U15523 (N_15523,N_15127,N_15375);
or U15524 (N_15524,N_15388,N_15416);
and U15525 (N_15525,N_15481,N_15019);
nand U15526 (N_15526,N_15333,N_15255);
or U15527 (N_15527,N_15262,N_15034);
or U15528 (N_15528,N_15134,N_15382);
and U15529 (N_15529,N_15107,N_15041);
xor U15530 (N_15530,N_15397,N_15258);
nand U15531 (N_15531,N_15302,N_15410);
nor U15532 (N_15532,N_15187,N_15363);
and U15533 (N_15533,N_15222,N_15219);
nand U15534 (N_15534,N_15492,N_15280);
nor U15535 (N_15535,N_15252,N_15028);
and U15536 (N_15536,N_15441,N_15081);
and U15537 (N_15537,N_15128,N_15419);
nand U15538 (N_15538,N_15101,N_15459);
xnor U15539 (N_15539,N_15298,N_15343);
nor U15540 (N_15540,N_15015,N_15215);
nor U15541 (N_15541,N_15077,N_15159);
nor U15542 (N_15542,N_15443,N_15281);
or U15543 (N_15543,N_15115,N_15049);
nand U15544 (N_15544,N_15290,N_15042);
nor U15545 (N_15545,N_15496,N_15324);
xor U15546 (N_15546,N_15461,N_15109);
and U15547 (N_15547,N_15286,N_15263);
nor U15548 (N_15548,N_15444,N_15018);
and U15549 (N_15549,N_15378,N_15105);
nand U15550 (N_15550,N_15275,N_15299);
xor U15551 (N_15551,N_15289,N_15268);
or U15552 (N_15552,N_15106,N_15111);
xor U15553 (N_15553,N_15192,N_15057);
or U15554 (N_15554,N_15352,N_15204);
nor U15555 (N_15555,N_15477,N_15149);
and U15556 (N_15556,N_15318,N_15167);
nand U15557 (N_15557,N_15328,N_15142);
or U15558 (N_15558,N_15347,N_15276);
xor U15559 (N_15559,N_15054,N_15146);
nor U15560 (N_15560,N_15487,N_15332);
xnor U15561 (N_15561,N_15438,N_15284);
or U15562 (N_15562,N_15495,N_15300);
xnor U15563 (N_15563,N_15446,N_15068);
or U15564 (N_15564,N_15110,N_15227);
and U15565 (N_15565,N_15112,N_15448);
nor U15566 (N_15566,N_15322,N_15434);
xnor U15567 (N_15567,N_15147,N_15355);
nand U15568 (N_15568,N_15216,N_15002);
nand U15569 (N_15569,N_15083,N_15455);
and U15570 (N_15570,N_15164,N_15313);
xor U15571 (N_15571,N_15010,N_15336);
or U15572 (N_15572,N_15038,N_15218);
nor U15573 (N_15573,N_15220,N_15493);
nor U15574 (N_15574,N_15223,N_15316);
nand U15575 (N_15575,N_15210,N_15207);
nand U15576 (N_15576,N_15392,N_15211);
or U15577 (N_15577,N_15125,N_15024);
nor U15578 (N_15578,N_15285,N_15072);
xor U15579 (N_15579,N_15294,N_15183);
or U15580 (N_15580,N_15458,N_15061);
nand U15581 (N_15581,N_15413,N_15367);
nand U15582 (N_15582,N_15426,N_15374);
xor U15583 (N_15583,N_15191,N_15237);
or U15584 (N_15584,N_15165,N_15138);
nor U15585 (N_15585,N_15079,N_15148);
nand U15586 (N_15586,N_15354,N_15314);
or U15587 (N_15587,N_15043,N_15278);
xor U15588 (N_15588,N_15005,N_15157);
xnor U15589 (N_15589,N_15436,N_15182);
nand U15590 (N_15590,N_15498,N_15221);
nand U15591 (N_15591,N_15190,N_15139);
nor U15592 (N_15592,N_15169,N_15209);
nand U15593 (N_15593,N_15412,N_15279);
or U15594 (N_15594,N_15283,N_15345);
nor U15595 (N_15595,N_15175,N_15305);
or U15596 (N_15596,N_15136,N_15062);
nor U15597 (N_15597,N_15226,N_15086);
nand U15598 (N_15598,N_15452,N_15118);
or U15599 (N_15599,N_15051,N_15472);
nor U15600 (N_15600,N_15337,N_15162);
and U15601 (N_15601,N_15174,N_15383);
and U15602 (N_15602,N_15338,N_15260);
xor U15603 (N_15603,N_15120,N_15121);
or U15604 (N_15604,N_15409,N_15240);
and U15605 (N_15605,N_15342,N_15188);
nand U15606 (N_15606,N_15287,N_15399);
or U15607 (N_15607,N_15428,N_15168);
or U15608 (N_15608,N_15346,N_15025);
nand U15609 (N_15609,N_15256,N_15090);
nand U15610 (N_15610,N_15423,N_15060);
nor U15611 (N_15611,N_15173,N_15202);
nand U15612 (N_15612,N_15026,N_15292);
or U15613 (N_15613,N_15447,N_15253);
and U15614 (N_15614,N_15376,N_15103);
nand U15615 (N_15615,N_15084,N_15301);
nand U15616 (N_15616,N_15321,N_15454);
nor U15617 (N_15617,N_15295,N_15479);
xnor U15618 (N_15618,N_15108,N_15497);
or U15619 (N_15619,N_15449,N_15488);
nor U15620 (N_15620,N_15037,N_15425);
nand U15621 (N_15621,N_15312,N_15214);
or U15622 (N_15622,N_15095,N_15066);
nor U15623 (N_15623,N_15415,N_15360);
xnor U15624 (N_15624,N_15414,N_15144);
or U15625 (N_15625,N_15063,N_15248);
and U15626 (N_15626,N_15031,N_15265);
nor U15627 (N_15627,N_15251,N_15059);
nand U15628 (N_15628,N_15156,N_15116);
nor U15629 (N_15629,N_15451,N_15291);
nand U15630 (N_15630,N_15132,N_15135);
xor U15631 (N_15631,N_15007,N_15004);
or U15632 (N_15632,N_15391,N_15001);
nor U15633 (N_15633,N_15208,N_15273);
nand U15634 (N_15634,N_15151,N_15235);
nor U15635 (N_15635,N_15073,N_15331);
xor U15636 (N_15636,N_15310,N_15200);
xnor U15637 (N_15637,N_15104,N_15254);
or U15638 (N_15638,N_15179,N_15274);
and U15639 (N_15639,N_15431,N_15442);
nand U15640 (N_15640,N_15377,N_15071);
or U15641 (N_15641,N_15201,N_15243);
nand U15642 (N_15642,N_15404,N_15470);
and U15643 (N_15643,N_15197,N_15439);
nand U15644 (N_15644,N_15203,N_15236);
nand U15645 (N_15645,N_15430,N_15379);
nor U15646 (N_15646,N_15320,N_15393);
and U15647 (N_15647,N_15385,N_15365);
or U15648 (N_15648,N_15349,N_15123);
nor U15649 (N_15649,N_15372,N_15099);
and U15650 (N_15650,N_15161,N_15315);
or U15651 (N_15651,N_15303,N_15114);
and U15652 (N_15652,N_15069,N_15422);
or U15653 (N_15653,N_15098,N_15213);
or U15654 (N_15654,N_15140,N_15023);
xor U15655 (N_15655,N_15045,N_15170);
nand U15656 (N_15656,N_15427,N_15166);
nor U15657 (N_15657,N_15239,N_15027);
nand U15658 (N_15658,N_15089,N_15198);
nand U15659 (N_15659,N_15406,N_15473);
xor U15660 (N_15660,N_15006,N_15466);
or U15661 (N_15661,N_15020,N_15076);
xnor U15662 (N_15662,N_15241,N_15405);
or U15663 (N_15663,N_15421,N_15091);
and U15664 (N_15664,N_15356,N_15131);
nor U15665 (N_15665,N_15032,N_15052);
nand U15666 (N_15666,N_15067,N_15065);
or U15667 (N_15667,N_15238,N_15196);
xnor U15668 (N_15668,N_15094,N_15311);
xnor U15669 (N_15669,N_15154,N_15491);
or U15670 (N_15670,N_15074,N_15351);
xnor U15671 (N_15671,N_15308,N_15186);
and U15672 (N_15672,N_15249,N_15499);
and U15673 (N_15673,N_15171,N_15467);
and U15674 (N_15674,N_15224,N_15119);
and U15675 (N_15675,N_15195,N_15158);
xor U15676 (N_15676,N_15133,N_15460);
nor U15677 (N_15677,N_15396,N_15056);
xnor U15678 (N_15678,N_15484,N_15229);
nor U15679 (N_15679,N_15417,N_15464);
nand U15680 (N_15680,N_15160,N_15327);
or U15681 (N_15681,N_15058,N_15075);
or U15682 (N_15682,N_15177,N_15270);
or U15683 (N_15683,N_15011,N_15309);
nor U15684 (N_15684,N_15009,N_15129);
and U15685 (N_15685,N_15228,N_15247);
and U15686 (N_15686,N_15334,N_15326);
nand U15687 (N_15687,N_15130,N_15475);
and U15688 (N_15688,N_15212,N_15370);
or U15689 (N_15689,N_15100,N_15093);
nor U15690 (N_15690,N_15319,N_15282);
and U15691 (N_15691,N_15261,N_15150);
and U15692 (N_15692,N_15102,N_15029);
or U15693 (N_15693,N_15035,N_15463);
nand U15694 (N_15694,N_15040,N_15402);
nand U15695 (N_15695,N_15184,N_15486);
nand U15696 (N_15696,N_15153,N_15036);
or U15697 (N_15697,N_15047,N_15335);
nor U15698 (N_15698,N_15242,N_15232);
or U15699 (N_15699,N_15117,N_15494);
nor U15700 (N_15700,N_15181,N_15231);
nor U15701 (N_15701,N_15469,N_15272);
nand U15702 (N_15702,N_15137,N_15245);
xnor U15703 (N_15703,N_15264,N_15476);
nor U15704 (N_15704,N_15122,N_15092);
and U15705 (N_15705,N_15000,N_15163);
or U15706 (N_15706,N_15435,N_15257);
nor U15707 (N_15707,N_15362,N_15176);
xnor U15708 (N_15708,N_15317,N_15380);
and U15709 (N_15709,N_15055,N_15017);
or U15710 (N_15710,N_15373,N_15205);
and U15711 (N_15711,N_15350,N_15113);
nand U15712 (N_15712,N_15126,N_15053);
or U15713 (N_15713,N_15483,N_15353);
and U15714 (N_15714,N_15304,N_15096);
nor U15715 (N_15715,N_15288,N_15401);
xnor U15716 (N_15716,N_15398,N_15050);
nand U15717 (N_15717,N_15244,N_15457);
or U15718 (N_15718,N_15440,N_15384);
xor U15719 (N_15719,N_15124,N_15250);
nand U15720 (N_15720,N_15465,N_15078);
nand U15721 (N_15721,N_15403,N_15445);
and U15722 (N_15722,N_15474,N_15307);
and U15723 (N_15723,N_15482,N_15323);
nand U15724 (N_15724,N_15012,N_15088);
nor U15725 (N_15725,N_15371,N_15269);
xor U15726 (N_15726,N_15450,N_15199);
and U15727 (N_15727,N_15390,N_15420);
nand U15728 (N_15728,N_15266,N_15395);
and U15729 (N_15729,N_15478,N_15030);
xor U15730 (N_15730,N_15082,N_15155);
and U15731 (N_15731,N_15152,N_15021);
and U15732 (N_15732,N_15277,N_15429);
nand U15733 (N_15733,N_15389,N_15407);
nand U15734 (N_15734,N_15489,N_15206);
xnor U15735 (N_15735,N_15141,N_15048);
and U15736 (N_15736,N_15039,N_15358);
or U15737 (N_15737,N_15424,N_15348);
or U15738 (N_15738,N_15408,N_15330);
and U15739 (N_15739,N_15085,N_15490);
and U15740 (N_15740,N_15225,N_15411);
nand U15741 (N_15741,N_15097,N_15189);
and U15742 (N_15742,N_15172,N_15178);
nor U15743 (N_15743,N_15008,N_15217);
nand U15744 (N_15744,N_15468,N_15233);
or U15745 (N_15745,N_15016,N_15033);
nor U15746 (N_15746,N_15394,N_15359);
and U15747 (N_15747,N_15387,N_15381);
and U15748 (N_15748,N_15339,N_15013);
nand U15749 (N_15749,N_15340,N_15271);
xnor U15750 (N_15750,N_15246,N_15149);
and U15751 (N_15751,N_15202,N_15104);
xor U15752 (N_15752,N_15391,N_15335);
or U15753 (N_15753,N_15400,N_15255);
or U15754 (N_15754,N_15163,N_15018);
nand U15755 (N_15755,N_15152,N_15324);
nand U15756 (N_15756,N_15407,N_15426);
and U15757 (N_15757,N_15224,N_15200);
nor U15758 (N_15758,N_15385,N_15227);
or U15759 (N_15759,N_15486,N_15395);
nand U15760 (N_15760,N_15212,N_15296);
nand U15761 (N_15761,N_15291,N_15001);
xnor U15762 (N_15762,N_15224,N_15070);
nor U15763 (N_15763,N_15239,N_15322);
nor U15764 (N_15764,N_15349,N_15020);
or U15765 (N_15765,N_15247,N_15310);
or U15766 (N_15766,N_15167,N_15050);
xor U15767 (N_15767,N_15126,N_15055);
or U15768 (N_15768,N_15428,N_15003);
nand U15769 (N_15769,N_15200,N_15322);
or U15770 (N_15770,N_15441,N_15039);
or U15771 (N_15771,N_15374,N_15022);
nor U15772 (N_15772,N_15040,N_15317);
nand U15773 (N_15773,N_15445,N_15279);
xnor U15774 (N_15774,N_15153,N_15002);
nand U15775 (N_15775,N_15328,N_15162);
nand U15776 (N_15776,N_15125,N_15071);
nand U15777 (N_15777,N_15422,N_15273);
nor U15778 (N_15778,N_15474,N_15212);
nand U15779 (N_15779,N_15157,N_15082);
xnor U15780 (N_15780,N_15397,N_15449);
or U15781 (N_15781,N_15237,N_15054);
xnor U15782 (N_15782,N_15121,N_15354);
nand U15783 (N_15783,N_15131,N_15162);
nand U15784 (N_15784,N_15047,N_15404);
or U15785 (N_15785,N_15244,N_15152);
nand U15786 (N_15786,N_15089,N_15367);
nand U15787 (N_15787,N_15072,N_15174);
and U15788 (N_15788,N_15163,N_15264);
or U15789 (N_15789,N_15478,N_15109);
xor U15790 (N_15790,N_15440,N_15383);
or U15791 (N_15791,N_15083,N_15493);
xor U15792 (N_15792,N_15041,N_15151);
or U15793 (N_15793,N_15110,N_15223);
nand U15794 (N_15794,N_15001,N_15171);
nor U15795 (N_15795,N_15424,N_15037);
nand U15796 (N_15796,N_15381,N_15357);
and U15797 (N_15797,N_15341,N_15488);
nor U15798 (N_15798,N_15233,N_15018);
nor U15799 (N_15799,N_15488,N_15486);
nand U15800 (N_15800,N_15248,N_15420);
and U15801 (N_15801,N_15416,N_15264);
nor U15802 (N_15802,N_15474,N_15090);
xnor U15803 (N_15803,N_15160,N_15238);
and U15804 (N_15804,N_15142,N_15244);
xor U15805 (N_15805,N_15431,N_15039);
and U15806 (N_15806,N_15289,N_15106);
and U15807 (N_15807,N_15069,N_15023);
nor U15808 (N_15808,N_15261,N_15229);
and U15809 (N_15809,N_15320,N_15334);
xnor U15810 (N_15810,N_15140,N_15467);
or U15811 (N_15811,N_15429,N_15216);
nand U15812 (N_15812,N_15289,N_15213);
and U15813 (N_15813,N_15244,N_15432);
nor U15814 (N_15814,N_15253,N_15331);
xor U15815 (N_15815,N_15371,N_15202);
xnor U15816 (N_15816,N_15425,N_15299);
or U15817 (N_15817,N_15386,N_15214);
xor U15818 (N_15818,N_15109,N_15138);
xnor U15819 (N_15819,N_15187,N_15495);
or U15820 (N_15820,N_15429,N_15301);
xor U15821 (N_15821,N_15002,N_15000);
xnor U15822 (N_15822,N_15208,N_15230);
nand U15823 (N_15823,N_15454,N_15019);
nand U15824 (N_15824,N_15232,N_15370);
nand U15825 (N_15825,N_15472,N_15162);
or U15826 (N_15826,N_15429,N_15054);
nand U15827 (N_15827,N_15327,N_15298);
nor U15828 (N_15828,N_15084,N_15019);
nor U15829 (N_15829,N_15320,N_15499);
and U15830 (N_15830,N_15321,N_15166);
nor U15831 (N_15831,N_15405,N_15118);
and U15832 (N_15832,N_15419,N_15317);
or U15833 (N_15833,N_15233,N_15029);
nand U15834 (N_15834,N_15327,N_15249);
or U15835 (N_15835,N_15231,N_15206);
or U15836 (N_15836,N_15189,N_15334);
nand U15837 (N_15837,N_15484,N_15099);
nor U15838 (N_15838,N_15493,N_15023);
xor U15839 (N_15839,N_15465,N_15457);
and U15840 (N_15840,N_15118,N_15317);
and U15841 (N_15841,N_15423,N_15313);
nand U15842 (N_15842,N_15113,N_15313);
nand U15843 (N_15843,N_15138,N_15444);
or U15844 (N_15844,N_15124,N_15328);
xor U15845 (N_15845,N_15235,N_15469);
nor U15846 (N_15846,N_15065,N_15175);
xnor U15847 (N_15847,N_15199,N_15309);
and U15848 (N_15848,N_15080,N_15472);
nor U15849 (N_15849,N_15482,N_15443);
or U15850 (N_15850,N_15154,N_15483);
xor U15851 (N_15851,N_15441,N_15000);
or U15852 (N_15852,N_15086,N_15074);
or U15853 (N_15853,N_15176,N_15234);
xnor U15854 (N_15854,N_15295,N_15223);
and U15855 (N_15855,N_15468,N_15314);
nor U15856 (N_15856,N_15263,N_15016);
nor U15857 (N_15857,N_15198,N_15304);
xnor U15858 (N_15858,N_15045,N_15352);
or U15859 (N_15859,N_15195,N_15396);
nand U15860 (N_15860,N_15447,N_15069);
nand U15861 (N_15861,N_15434,N_15074);
nand U15862 (N_15862,N_15301,N_15119);
or U15863 (N_15863,N_15355,N_15360);
or U15864 (N_15864,N_15340,N_15416);
xor U15865 (N_15865,N_15499,N_15216);
nor U15866 (N_15866,N_15191,N_15407);
nand U15867 (N_15867,N_15463,N_15032);
nor U15868 (N_15868,N_15173,N_15472);
xor U15869 (N_15869,N_15428,N_15250);
and U15870 (N_15870,N_15478,N_15140);
nor U15871 (N_15871,N_15370,N_15135);
xnor U15872 (N_15872,N_15131,N_15019);
and U15873 (N_15873,N_15002,N_15387);
and U15874 (N_15874,N_15296,N_15422);
nand U15875 (N_15875,N_15250,N_15034);
and U15876 (N_15876,N_15228,N_15034);
xnor U15877 (N_15877,N_15282,N_15154);
nand U15878 (N_15878,N_15102,N_15382);
nor U15879 (N_15879,N_15191,N_15219);
and U15880 (N_15880,N_15043,N_15197);
xnor U15881 (N_15881,N_15482,N_15064);
and U15882 (N_15882,N_15170,N_15337);
nand U15883 (N_15883,N_15187,N_15209);
xor U15884 (N_15884,N_15295,N_15484);
or U15885 (N_15885,N_15495,N_15018);
nor U15886 (N_15886,N_15055,N_15297);
and U15887 (N_15887,N_15367,N_15047);
nand U15888 (N_15888,N_15492,N_15360);
xnor U15889 (N_15889,N_15241,N_15155);
nor U15890 (N_15890,N_15231,N_15377);
xor U15891 (N_15891,N_15200,N_15434);
nand U15892 (N_15892,N_15389,N_15002);
nor U15893 (N_15893,N_15280,N_15254);
or U15894 (N_15894,N_15296,N_15142);
nand U15895 (N_15895,N_15409,N_15157);
xnor U15896 (N_15896,N_15017,N_15419);
or U15897 (N_15897,N_15333,N_15448);
or U15898 (N_15898,N_15174,N_15365);
nor U15899 (N_15899,N_15243,N_15004);
or U15900 (N_15900,N_15398,N_15229);
nand U15901 (N_15901,N_15437,N_15448);
nand U15902 (N_15902,N_15356,N_15470);
and U15903 (N_15903,N_15195,N_15008);
or U15904 (N_15904,N_15072,N_15318);
and U15905 (N_15905,N_15091,N_15446);
or U15906 (N_15906,N_15118,N_15241);
and U15907 (N_15907,N_15235,N_15490);
xnor U15908 (N_15908,N_15474,N_15429);
or U15909 (N_15909,N_15057,N_15272);
and U15910 (N_15910,N_15130,N_15053);
or U15911 (N_15911,N_15291,N_15345);
nor U15912 (N_15912,N_15056,N_15092);
xor U15913 (N_15913,N_15051,N_15425);
nand U15914 (N_15914,N_15354,N_15358);
or U15915 (N_15915,N_15420,N_15172);
xor U15916 (N_15916,N_15051,N_15274);
nand U15917 (N_15917,N_15125,N_15243);
and U15918 (N_15918,N_15304,N_15483);
or U15919 (N_15919,N_15411,N_15286);
or U15920 (N_15920,N_15322,N_15234);
nand U15921 (N_15921,N_15389,N_15285);
nand U15922 (N_15922,N_15459,N_15468);
and U15923 (N_15923,N_15066,N_15424);
xnor U15924 (N_15924,N_15288,N_15234);
or U15925 (N_15925,N_15029,N_15017);
nand U15926 (N_15926,N_15063,N_15254);
nand U15927 (N_15927,N_15298,N_15326);
xnor U15928 (N_15928,N_15093,N_15034);
nand U15929 (N_15929,N_15358,N_15026);
and U15930 (N_15930,N_15259,N_15031);
nor U15931 (N_15931,N_15049,N_15365);
xor U15932 (N_15932,N_15023,N_15031);
or U15933 (N_15933,N_15291,N_15307);
xor U15934 (N_15934,N_15323,N_15404);
or U15935 (N_15935,N_15371,N_15334);
xor U15936 (N_15936,N_15185,N_15287);
and U15937 (N_15937,N_15314,N_15197);
or U15938 (N_15938,N_15479,N_15317);
or U15939 (N_15939,N_15445,N_15349);
nand U15940 (N_15940,N_15028,N_15146);
or U15941 (N_15941,N_15199,N_15364);
nand U15942 (N_15942,N_15471,N_15474);
nor U15943 (N_15943,N_15092,N_15320);
nand U15944 (N_15944,N_15290,N_15252);
nor U15945 (N_15945,N_15333,N_15471);
or U15946 (N_15946,N_15126,N_15170);
and U15947 (N_15947,N_15229,N_15295);
or U15948 (N_15948,N_15171,N_15477);
xor U15949 (N_15949,N_15134,N_15065);
nand U15950 (N_15950,N_15297,N_15281);
and U15951 (N_15951,N_15146,N_15474);
nand U15952 (N_15952,N_15048,N_15209);
nor U15953 (N_15953,N_15434,N_15124);
nand U15954 (N_15954,N_15222,N_15165);
xor U15955 (N_15955,N_15436,N_15221);
or U15956 (N_15956,N_15161,N_15449);
or U15957 (N_15957,N_15282,N_15333);
nand U15958 (N_15958,N_15031,N_15302);
or U15959 (N_15959,N_15351,N_15097);
or U15960 (N_15960,N_15328,N_15070);
nor U15961 (N_15961,N_15202,N_15065);
or U15962 (N_15962,N_15485,N_15013);
nor U15963 (N_15963,N_15485,N_15493);
nor U15964 (N_15964,N_15096,N_15439);
nor U15965 (N_15965,N_15385,N_15253);
nand U15966 (N_15966,N_15273,N_15414);
or U15967 (N_15967,N_15095,N_15361);
nor U15968 (N_15968,N_15228,N_15345);
nor U15969 (N_15969,N_15215,N_15284);
nor U15970 (N_15970,N_15404,N_15273);
nand U15971 (N_15971,N_15032,N_15152);
or U15972 (N_15972,N_15492,N_15252);
and U15973 (N_15973,N_15334,N_15191);
nor U15974 (N_15974,N_15262,N_15273);
or U15975 (N_15975,N_15168,N_15094);
xnor U15976 (N_15976,N_15016,N_15295);
nor U15977 (N_15977,N_15273,N_15008);
nand U15978 (N_15978,N_15355,N_15158);
xor U15979 (N_15979,N_15255,N_15477);
and U15980 (N_15980,N_15387,N_15255);
nor U15981 (N_15981,N_15231,N_15059);
nand U15982 (N_15982,N_15470,N_15082);
and U15983 (N_15983,N_15188,N_15100);
nand U15984 (N_15984,N_15305,N_15301);
nand U15985 (N_15985,N_15455,N_15267);
and U15986 (N_15986,N_15243,N_15337);
or U15987 (N_15987,N_15289,N_15129);
nor U15988 (N_15988,N_15010,N_15118);
xor U15989 (N_15989,N_15292,N_15308);
and U15990 (N_15990,N_15424,N_15360);
nand U15991 (N_15991,N_15050,N_15082);
and U15992 (N_15992,N_15359,N_15233);
xor U15993 (N_15993,N_15038,N_15266);
nor U15994 (N_15994,N_15249,N_15068);
or U15995 (N_15995,N_15204,N_15235);
or U15996 (N_15996,N_15377,N_15315);
or U15997 (N_15997,N_15419,N_15129);
xor U15998 (N_15998,N_15047,N_15063);
and U15999 (N_15999,N_15094,N_15161);
xor U16000 (N_16000,N_15966,N_15896);
and U16001 (N_16001,N_15993,N_15839);
xor U16002 (N_16002,N_15644,N_15987);
nor U16003 (N_16003,N_15822,N_15678);
nand U16004 (N_16004,N_15691,N_15542);
nand U16005 (N_16005,N_15507,N_15503);
or U16006 (N_16006,N_15878,N_15834);
nand U16007 (N_16007,N_15808,N_15932);
and U16008 (N_16008,N_15805,N_15587);
nor U16009 (N_16009,N_15957,N_15798);
xnor U16010 (N_16010,N_15622,N_15779);
or U16011 (N_16011,N_15649,N_15717);
or U16012 (N_16012,N_15860,N_15914);
or U16013 (N_16013,N_15601,N_15763);
and U16014 (N_16014,N_15929,N_15999);
and U16015 (N_16015,N_15652,N_15922);
or U16016 (N_16016,N_15845,N_15648);
xor U16017 (N_16017,N_15558,N_15597);
xor U16018 (N_16018,N_15603,N_15902);
nor U16019 (N_16019,N_15546,N_15982);
and U16020 (N_16020,N_15619,N_15864);
and U16021 (N_16021,N_15872,N_15515);
nand U16022 (N_16022,N_15826,N_15662);
nand U16023 (N_16023,N_15672,N_15547);
nand U16024 (N_16024,N_15856,N_15916);
or U16025 (N_16025,N_15959,N_15668);
xnor U16026 (N_16026,N_15623,N_15725);
xor U16027 (N_16027,N_15835,N_15752);
and U16028 (N_16028,N_15680,N_15727);
or U16029 (N_16029,N_15550,N_15733);
nor U16030 (N_16030,N_15536,N_15741);
xor U16031 (N_16031,N_15769,N_15640);
or U16032 (N_16032,N_15970,N_15998);
xor U16033 (N_16033,N_15683,N_15750);
nand U16034 (N_16034,N_15595,N_15947);
or U16035 (N_16035,N_15512,N_15833);
nor U16036 (N_16036,N_15992,N_15551);
or U16037 (N_16037,N_15608,N_15517);
nand U16038 (N_16038,N_15554,N_15905);
or U16039 (N_16039,N_15630,N_15876);
nand U16040 (N_16040,N_15949,N_15890);
or U16041 (N_16041,N_15961,N_15962);
nand U16042 (N_16042,N_15565,N_15730);
nor U16043 (N_16043,N_15837,N_15829);
nor U16044 (N_16044,N_15592,N_15624);
nand U16045 (N_16045,N_15761,N_15726);
and U16046 (N_16046,N_15765,N_15944);
nor U16047 (N_16047,N_15951,N_15943);
xnor U16048 (N_16048,N_15504,N_15548);
and U16049 (N_16049,N_15895,N_15768);
and U16050 (N_16050,N_15981,N_15851);
nor U16051 (N_16051,N_15607,N_15915);
xnor U16052 (N_16052,N_15852,N_15540);
nor U16053 (N_16053,N_15569,N_15994);
or U16054 (N_16054,N_15722,N_15718);
nand U16055 (N_16055,N_15816,N_15948);
nor U16056 (N_16056,N_15588,N_15828);
xor U16057 (N_16057,N_15917,N_15539);
or U16058 (N_16058,N_15582,N_15527);
nor U16059 (N_16059,N_15514,N_15973);
or U16060 (N_16060,N_15941,N_15656);
nand U16061 (N_16061,N_15921,N_15535);
or U16062 (N_16062,N_15964,N_15708);
nand U16063 (N_16063,N_15789,N_15575);
nand U16064 (N_16064,N_15931,N_15711);
xor U16065 (N_16065,N_15502,N_15907);
or U16066 (N_16066,N_15738,N_15759);
nand U16067 (N_16067,N_15781,N_15795);
nand U16068 (N_16068,N_15985,N_15628);
nand U16069 (N_16069,N_15681,N_15863);
nor U16070 (N_16070,N_15654,N_15563);
nor U16071 (N_16071,N_15918,N_15538);
nor U16072 (N_16072,N_15780,N_15745);
nor U16073 (N_16073,N_15661,N_15618);
xnor U16074 (N_16074,N_15614,N_15942);
and U16075 (N_16075,N_15885,N_15658);
and U16076 (N_16076,N_15511,N_15621);
or U16077 (N_16077,N_15785,N_15609);
and U16078 (N_16078,N_15653,N_15626);
nand U16079 (N_16079,N_15946,N_15616);
nand U16080 (N_16080,N_15685,N_15701);
or U16081 (N_16081,N_15743,N_15848);
nor U16082 (N_16082,N_15911,N_15841);
nand U16083 (N_16083,N_15854,N_15865);
nor U16084 (N_16084,N_15858,N_15663);
and U16085 (N_16085,N_15953,N_15713);
nand U16086 (N_16086,N_15632,N_15908);
and U16087 (N_16087,N_15500,N_15728);
nand U16088 (N_16088,N_15753,N_15742);
nor U16089 (N_16089,N_15818,N_15573);
or U16090 (N_16090,N_15593,N_15891);
xor U16091 (N_16091,N_15821,N_15716);
nand U16092 (N_16092,N_15843,N_15797);
or U16093 (N_16093,N_15576,N_15963);
nand U16094 (N_16094,N_15977,N_15846);
xor U16095 (N_16095,N_15838,N_15897);
nor U16096 (N_16096,N_15635,N_15506);
nand U16097 (N_16097,N_15710,N_15552);
or U16098 (N_16098,N_15901,N_15541);
nand U16099 (N_16099,N_15806,N_15887);
xor U16100 (N_16100,N_15651,N_15737);
xnor U16101 (N_16101,N_15572,N_15571);
nand U16102 (N_16102,N_15686,N_15699);
or U16103 (N_16103,N_15655,N_15937);
nand U16104 (N_16104,N_15873,N_15871);
nor U16105 (N_16105,N_15697,N_15862);
and U16106 (N_16106,N_15979,N_15849);
nor U16107 (N_16107,N_15602,N_15721);
nand U16108 (N_16108,N_15532,N_15620);
or U16109 (N_16109,N_15801,N_15700);
or U16110 (N_16110,N_15581,N_15513);
nand U16111 (N_16111,N_15978,N_15531);
and U16112 (N_16112,N_15804,N_15819);
or U16113 (N_16113,N_15952,N_15831);
and U16114 (N_16114,N_15731,N_15525);
and U16115 (N_16115,N_15612,N_15880);
nand U16116 (N_16116,N_15783,N_15799);
and U16117 (N_16117,N_15589,N_15800);
nor U16118 (N_16118,N_15936,N_15754);
or U16119 (N_16119,N_15583,N_15694);
and U16120 (N_16120,N_15639,N_15764);
nand U16121 (N_16121,N_15627,N_15928);
and U16122 (N_16122,N_15501,N_15671);
nand U16123 (N_16123,N_15776,N_15972);
xnor U16124 (N_16124,N_15996,N_15555);
xor U16125 (N_16125,N_15889,N_15631);
xor U16126 (N_16126,N_15762,N_15698);
and U16127 (N_16127,N_15598,N_15794);
nor U16128 (N_16128,N_15919,N_15886);
nor U16129 (N_16129,N_15903,N_15774);
or U16130 (N_16130,N_15590,N_15820);
nor U16131 (N_16131,N_15666,N_15969);
and U16132 (N_16132,N_15604,N_15874);
nor U16133 (N_16133,N_15770,N_15875);
nor U16134 (N_16134,N_15940,N_15657);
and U16135 (N_16135,N_15610,N_15773);
or U16136 (N_16136,N_15633,N_15732);
and U16137 (N_16137,N_15578,N_15545);
nand U16138 (N_16138,N_15677,N_15585);
or U16139 (N_16139,N_15850,N_15706);
nor U16140 (N_16140,N_15664,N_15958);
and U16141 (N_16141,N_15510,N_15667);
or U16142 (N_16142,N_15586,N_15508);
and U16143 (N_16143,N_15522,N_15720);
nand U16144 (N_16144,N_15778,N_15810);
and U16145 (N_16145,N_15559,N_15782);
nand U16146 (N_16146,N_15791,N_15647);
xor U16147 (N_16147,N_15636,N_15516);
nor U16148 (N_16148,N_15827,N_15988);
or U16149 (N_16149,N_15606,N_15520);
xor U16150 (N_16150,N_15910,N_15815);
xor U16151 (N_16151,N_15817,N_15809);
nor U16152 (N_16152,N_15509,N_15669);
nor U16153 (N_16153,N_15906,N_15719);
and U16154 (N_16154,N_15641,N_15986);
nor U16155 (N_16155,N_15983,N_15505);
or U16156 (N_16156,N_15675,N_15629);
xnor U16157 (N_16157,N_15847,N_15796);
or U16158 (N_16158,N_15660,N_15646);
or U16159 (N_16159,N_15557,N_15913);
or U16160 (N_16160,N_15784,N_15617);
nand U16161 (N_16161,N_15537,N_15574);
or U16162 (N_16162,N_15688,N_15830);
xor U16163 (N_16163,N_15549,N_15740);
xor U16164 (N_16164,N_15676,N_15637);
nor U16165 (N_16165,N_15645,N_15693);
and U16166 (N_16166,N_15855,N_15989);
xnor U16167 (N_16167,N_15923,N_15965);
and U16168 (N_16168,N_15634,N_15758);
xor U16169 (N_16169,N_15665,N_15591);
or U16170 (N_16170,N_15894,N_15904);
xor U16171 (N_16171,N_15544,N_15920);
xnor U16172 (N_16172,N_15939,N_15771);
and U16173 (N_16173,N_15570,N_15898);
or U16174 (N_16174,N_15812,N_15879);
xnor U16175 (N_16175,N_15735,N_15579);
nor U16176 (N_16176,N_15792,N_15926);
or U16177 (N_16177,N_15883,N_15682);
nand U16178 (N_16178,N_15975,N_15523);
nor U16179 (N_16179,N_15772,N_15567);
nor U16180 (N_16180,N_15811,N_15755);
xor U16181 (N_16181,N_15519,N_15705);
or U16182 (N_16182,N_15638,N_15802);
xnor U16183 (N_16183,N_15707,N_15956);
or U16184 (N_16184,N_15882,N_15980);
nand U16185 (N_16185,N_15611,N_15751);
xor U16186 (N_16186,N_15881,N_15560);
nand U16187 (N_16187,N_15533,N_15766);
and U16188 (N_16188,N_15723,N_15739);
and U16189 (N_16189,N_15518,N_15840);
and U16190 (N_16190,N_15909,N_15715);
nand U16191 (N_16191,N_15945,N_15642);
xor U16192 (N_16192,N_15788,N_15925);
nor U16193 (N_16193,N_15714,N_15692);
and U16194 (N_16194,N_15892,N_15775);
and U16195 (N_16195,N_15786,N_15674);
and U16196 (N_16196,N_15529,N_15613);
and U16197 (N_16197,N_15760,N_15704);
nor U16198 (N_16198,N_15553,N_15836);
nand U16199 (N_16199,N_15562,N_15596);
nor U16200 (N_16200,N_15859,N_15689);
xnor U16201 (N_16201,N_15971,N_15787);
xnor U16202 (N_16202,N_15884,N_15832);
or U16203 (N_16203,N_15927,N_15673);
nor U16204 (N_16204,N_15564,N_15561);
or U16205 (N_16205,N_15709,N_15568);
or U16206 (N_16206,N_15650,N_15934);
or U16207 (N_16207,N_15580,N_15955);
xor U16208 (N_16208,N_15659,N_15615);
nor U16209 (N_16209,N_15984,N_15991);
xnor U16210 (N_16210,N_15997,N_15748);
xor U16211 (N_16211,N_15777,N_15825);
xnor U16212 (N_16212,N_15888,N_15703);
nand U16213 (N_16213,N_15690,N_15756);
nand U16214 (N_16214,N_15950,N_15877);
xnor U16215 (N_16215,N_15670,N_15749);
or U16216 (N_16216,N_15790,N_15813);
nor U16217 (N_16217,N_15976,N_15767);
xnor U16218 (N_16218,N_15747,N_15857);
nor U16219 (N_16219,N_15967,N_15599);
nand U16220 (N_16220,N_15729,N_15930);
or U16221 (N_16221,N_15566,N_15974);
or U16222 (N_16222,N_15724,N_15534);
or U16223 (N_16223,N_15530,N_15679);
nand U16224 (N_16224,N_15995,N_15695);
xnor U16225 (N_16225,N_15844,N_15935);
xnor U16226 (N_16226,N_15600,N_15893);
or U16227 (N_16227,N_15900,N_15736);
xor U16228 (N_16228,N_15853,N_15861);
nand U16229 (N_16229,N_15757,N_15968);
nor U16230 (N_16230,N_15543,N_15990);
nor U16231 (N_16231,N_15869,N_15814);
xnor U16232 (N_16232,N_15556,N_15594);
xor U16233 (N_16233,N_15524,N_15521);
and U16234 (N_16234,N_15526,N_15528);
xnor U16235 (N_16235,N_15643,N_15954);
nor U16236 (N_16236,N_15866,N_15702);
or U16237 (N_16237,N_15734,N_15823);
nand U16238 (N_16238,N_15899,N_15868);
or U16239 (N_16239,N_15712,N_15867);
nor U16240 (N_16240,N_15824,N_15924);
nor U16241 (N_16241,N_15870,N_15625);
nor U16242 (N_16242,N_15744,N_15803);
or U16243 (N_16243,N_15746,N_15793);
or U16244 (N_16244,N_15577,N_15960);
nand U16245 (N_16245,N_15687,N_15696);
nor U16246 (N_16246,N_15938,N_15807);
and U16247 (N_16247,N_15605,N_15584);
or U16248 (N_16248,N_15912,N_15684);
and U16249 (N_16249,N_15842,N_15933);
nor U16250 (N_16250,N_15677,N_15790);
nand U16251 (N_16251,N_15519,N_15679);
nand U16252 (N_16252,N_15690,N_15651);
xor U16253 (N_16253,N_15849,N_15829);
or U16254 (N_16254,N_15719,N_15538);
xor U16255 (N_16255,N_15671,N_15761);
nor U16256 (N_16256,N_15926,N_15977);
nand U16257 (N_16257,N_15733,N_15999);
nand U16258 (N_16258,N_15730,N_15618);
or U16259 (N_16259,N_15929,N_15946);
nor U16260 (N_16260,N_15644,N_15688);
and U16261 (N_16261,N_15553,N_15882);
nor U16262 (N_16262,N_15758,N_15712);
xor U16263 (N_16263,N_15862,N_15950);
nor U16264 (N_16264,N_15724,N_15672);
and U16265 (N_16265,N_15509,N_15865);
or U16266 (N_16266,N_15747,N_15570);
nor U16267 (N_16267,N_15828,N_15684);
xor U16268 (N_16268,N_15773,N_15826);
or U16269 (N_16269,N_15966,N_15752);
xnor U16270 (N_16270,N_15569,N_15636);
and U16271 (N_16271,N_15609,N_15851);
nand U16272 (N_16272,N_15511,N_15802);
and U16273 (N_16273,N_15639,N_15840);
or U16274 (N_16274,N_15929,N_15905);
nand U16275 (N_16275,N_15511,N_15815);
xor U16276 (N_16276,N_15938,N_15850);
xor U16277 (N_16277,N_15522,N_15894);
xor U16278 (N_16278,N_15869,N_15641);
and U16279 (N_16279,N_15702,N_15679);
and U16280 (N_16280,N_15647,N_15557);
nor U16281 (N_16281,N_15755,N_15838);
nor U16282 (N_16282,N_15783,N_15986);
and U16283 (N_16283,N_15612,N_15819);
nand U16284 (N_16284,N_15565,N_15716);
nor U16285 (N_16285,N_15707,N_15891);
and U16286 (N_16286,N_15755,N_15870);
or U16287 (N_16287,N_15810,N_15794);
and U16288 (N_16288,N_15769,N_15995);
or U16289 (N_16289,N_15909,N_15660);
or U16290 (N_16290,N_15860,N_15836);
nor U16291 (N_16291,N_15508,N_15620);
nor U16292 (N_16292,N_15651,N_15998);
or U16293 (N_16293,N_15540,N_15934);
nor U16294 (N_16294,N_15571,N_15537);
xnor U16295 (N_16295,N_15866,N_15597);
and U16296 (N_16296,N_15920,N_15653);
nor U16297 (N_16297,N_15946,N_15711);
or U16298 (N_16298,N_15733,N_15520);
or U16299 (N_16299,N_15560,N_15548);
nor U16300 (N_16300,N_15708,N_15525);
nand U16301 (N_16301,N_15681,N_15896);
or U16302 (N_16302,N_15899,N_15623);
xnor U16303 (N_16303,N_15982,N_15758);
and U16304 (N_16304,N_15980,N_15951);
and U16305 (N_16305,N_15732,N_15940);
or U16306 (N_16306,N_15510,N_15695);
or U16307 (N_16307,N_15747,N_15513);
or U16308 (N_16308,N_15724,N_15775);
and U16309 (N_16309,N_15636,N_15760);
nand U16310 (N_16310,N_15530,N_15910);
nor U16311 (N_16311,N_15799,N_15807);
nand U16312 (N_16312,N_15567,N_15990);
nand U16313 (N_16313,N_15761,N_15631);
nor U16314 (N_16314,N_15851,N_15628);
xnor U16315 (N_16315,N_15976,N_15797);
nor U16316 (N_16316,N_15972,N_15757);
or U16317 (N_16317,N_15757,N_15839);
or U16318 (N_16318,N_15938,N_15653);
and U16319 (N_16319,N_15809,N_15955);
nor U16320 (N_16320,N_15639,N_15855);
nor U16321 (N_16321,N_15761,N_15734);
xnor U16322 (N_16322,N_15645,N_15910);
xnor U16323 (N_16323,N_15891,N_15773);
and U16324 (N_16324,N_15670,N_15943);
nor U16325 (N_16325,N_15696,N_15688);
and U16326 (N_16326,N_15531,N_15921);
nor U16327 (N_16327,N_15723,N_15668);
xnor U16328 (N_16328,N_15520,N_15668);
nand U16329 (N_16329,N_15956,N_15886);
nor U16330 (N_16330,N_15559,N_15760);
or U16331 (N_16331,N_15703,N_15853);
and U16332 (N_16332,N_15980,N_15953);
nand U16333 (N_16333,N_15672,N_15933);
and U16334 (N_16334,N_15597,N_15956);
nand U16335 (N_16335,N_15908,N_15827);
or U16336 (N_16336,N_15854,N_15810);
nand U16337 (N_16337,N_15754,N_15648);
xor U16338 (N_16338,N_15817,N_15551);
nor U16339 (N_16339,N_15564,N_15606);
and U16340 (N_16340,N_15518,N_15546);
nor U16341 (N_16341,N_15861,N_15832);
xor U16342 (N_16342,N_15569,N_15689);
nor U16343 (N_16343,N_15646,N_15948);
or U16344 (N_16344,N_15783,N_15980);
or U16345 (N_16345,N_15583,N_15999);
nor U16346 (N_16346,N_15811,N_15831);
nand U16347 (N_16347,N_15588,N_15535);
nor U16348 (N_16348,N_15906,N_15746);
xnor U16349 (N_16349,N_15815,N_15890);
and U16350 (N_16350,N_15638,N_15886);
xnor U16351 (N_16351,N_15752,N_15757);
or U16352 (N_16352,N_15990,N_15837);
or U16353 (N_16353,N_15718,N_15526);
or U16354 (N_16354,N_15928,N_15749);
xnor U16355 (N_16355,N_15567,N_15718);
xnor U16356 (N_16356,N_15762,N_15753);
nor U16357 (N_16357,N_15630,N_15774);
nor U16358 (N_16358,N_15880,N_15912);
and U16359 (N_16359,N_15849,N_15961);
and U16360 (N_16360,N_15641,N_15569);
nand U16361 (N_16361,N_15953,N_15507);
xnor U16362 (N_16362,N_15767,N_15761);
xor U16363 (N_16363,N_15532,N_15896);
xnor U16364 (N_16364,N_15866,N_15630);
nand U16365 (N_16365,N_15827,N_15951);
and U16366 (N_16366,N_15981,N_15859);
and U16367 (N_16367,N_15517,N_15797);
nand U16368 (N_16368,N_15501,N_15695);
or U16369 (N_16369,N_15690,N_15965);
xnor U16370 (N_16370,N_15659,N_15900);
nor U16371 (N_16371,N_15541,N_15757);
or U16372 (N_16372,N_15830,N_15600);
and U16373 (N_16373,N_15748,N_15681);
nand U16374 (N_16374,N_15680,N_15844);
nor U16375 (N_16375,N_15968,N_15530);
xor U16376 (N_16376,N_15919,N_15862);
or U16377 (N_16377,N_15939,N_15770);
and U16378 (N_16378,N_15761,N_15609);
or U16379 (N_16379,N_15851,N_15614);
or U16380 (N_16380,N_15921,N_15826);
xor U16381 (N_16381,N_15807,N_15864);
and U16382 (N_16382,N_15926,N_15598);
and U16383 (N_16383,N_15629,N_15598);
nand U16384 (N_16384,N_15724,N_15705);
xnor U16385 (N_16385,N_15729,N_15589);
and U16386 (N_16386,N_15528,N_15747);
and U16387 (N_16387,N_15849,N_15753);
nor U16388 (N_16388,N_15511,N_15721);
nor U16389 (N_16389,N_15899,N_15843);
xnor U16390 (N_16390,N_15714,N_15732);
xor U16391 (N_16391,N_15570,N_15890);
nand U16392 (N_16392,N_15594,N_15653);
or U16393 (N_16393,N_15707,N_15530);
or U16394 (N_16394,N_15750,N_15996);
and U16395 (N_16395,N_15852,N_15806);
or U16396 (N_16396,N_15527,N_15987);
or U16397 (N_16397,N_15758,N_15640);
nand U16398 (N_16398,N_15726,N_15708);
and U16399 (N_16399,N_15765,N_15615);
nand U16400 (N_16400,N_15686,N_15831);
and U16401 (N_16401,N_15900,N_15968);
nand U16402 (N_16402,N_15961,N_15972);
or U16403 (N_16403,N_15725,N_15935);
nor U16404 (N_16404,N_15655,N_15774);
and U16405 (N_16405,N_15707,N_15949);
nand U16406 (N_16406,N_15750,N_15924);
xor U16407 (N_16407,N_15668,N_15801);
nand U16408 (N_16408,N_15938,N_15806);
xor U16409 (N_16409,N_15854,N_15684);
nand U16410 (N_16410,N_15857,N_15852);
xnor U16411 (N_16411,N_15921,N_15528);
nor U16412 (N_16412,N_15628,N_15588);
xor U16413 (N_16413,N_15530,N_15589);
nand U16414 (N_16414,N_15941,N_15662);
nand U16415 (N_16415,N_15604,N_15501);
and U16416 (N_16416,N_15859,N_15677);
xnor U16417 (N_16417,N_15565,N_15580);
and U16418 (N_16418,N_15583,N_15884);
or U16419 (N_16419,N_15753,N_15632);
xnor U16420 (N_16420,N_15959,N_15717);
and U16421 (N_16421,N_15832,N_15767);
or U16422 (N_16422,N_15917,N_15965);
xor U16423 (N_16423,N_15528,N_15854);
nand U16424 (N_16424,N_15574,N_15730);
or U16425 (N_16425,N_15814,N_15888);
and U16426 (N_16426,N_15790,N_15664);
xnor U16427 (N_16427,N_15591,N_15701);
xnor U16428 (N_16428,N_15726,N_15512);
nor U16429 (N_16429,N_15682,N_15891);
xnor U16430 (N_16430,N_15870,N_15658);
nand U16431 (N_16431,N_15760,N_15861);
xnor U16432 (N_16432,N_15949,N_15694);
xnor U16433 (N_16433,N_15812,N_15821);
and U16434 (N_16434,N_15623,N_15668);
xnor U16435 (N_16435,N_15791,N_15969);
xnor U16436 (N_16436,N_15589,N_15780);
or U16437 (N_16437,N_15899,N_15746);
nand U16438 (N_16438,N_15855,N_15596);
nand U16439 (N_16439,N_15661,N_15943);
xnor U16440 (N_16440,N_15839,N_15511);
xnor U16441 (N_16441,N_15853,N_15798);
nor U16442 (N_16442,N_15503,N_15674);
nand U16443 (N_16443,N_15502,N_15655);
nand U16444 (N_16444,N_15981,N_15916);
xor U16445 (N_16445,N_15739,N_15814);
and U16446 (N_16446,N_15627,N_15825);
and U16447 (N_16447,N_15796,N_15610);
and U16448 (N_16448,N_15652,N_15785);
nor U16449 (N_16449,N_15867,N_15793);
nor U16450 (N_16450,N_15563,N_15517);
and U16451 (N_16451,N_15575,N_15777);
nor U16452 (N_16452,N_15679,N_15665);
xor U16453 (N_16453,N_15766,N_15655);
nand U16454 (N_16454,N_15884,N_15712);
xor U16455 (N_16455,N_15968,N_15771);
or U16456 (N_16456,N_15664,N_15658);
nor U16457 (N_16457,N_15674,N_15542);
nand U16458 (N_16458,N_15717,N_15806);
nor U16459 (N_16459,N_15962,N_15631);
or U16460 (N_16460,N_15909,N_15816);
nor U16461 (N_16461,N_15717,N_15626);
nor U16462 (N_16462,N_15767,N_15623);
and U16463 (N_16463,N_15962,N_15881);
nand U16464 (N_16464,N_15567,N_15674);
xor U16465 (N_16465,N_15512,N_15960);
xnor U16466 (N_16466,N_15506,N_15596);
and U16467 (N_16467,N_15903,N_15781);
xor U16468 (N_16468,N_15824,N_15990);
and U16469 (N_16469,N_15720,N_15930);
or U16470 (N_16470,N_15540,N_15727);
and U16471 (N_16471,N_15877,N_15868);
or U16472 (N_16472,N_15884,N_15932);
and U16473 (N_16473,N_15635,N_15799);
nor U16474 (N_16474,N_15929,N_15869);
and U16475 (N_16475,N_15829,N_15817);
or U16476 (N_16476,N_15682,N_15997);
nand U16477 (N_16477,N_15863,N_15569);
and U16478 (N_16478,N_15594,N_15652);
nand U16479 (N_16479,N_15543,N_15806);
nor U16480 (N_16480,N_15835,N_15959);
xor U16481 (N_16481,N_15981,N_15902);
and U16482 (N_16482,N_15693,N_15832);
nor U16483 (N_16483,N_15808,N_15964);
xor U16484 (N_16484,N_15694,N_15518);
nand U16485 (N_16485,N_15594,N_15898);
xnor U16486 (N_16486,N_15544,N_15797);
nand U16487 (N_16487,N_15540,N_15569);
xor U16488 (N_16488,N_15847,N_15908);
or U16489 (N_16489,N_15588,N_15882);
nand U16490 (N_16490,N_15794,N_15680);
xor U16491 (N_16491,N_15550,N_15830);
xor U16492 (N_16492,N_15579,N_15810);
nor U16493 (N_16493,N_15843,N_15806);
or U16494 (N_16494,N_15656,N_15910);
nor U16495 (N_16495,N_15682,N_15821);
or U16496 (N_16496,N_15553,N_15912);
or U16497 (N_16497,N_15835,N_15504);
nor U16498 (N_16498,N_15658,N_15743);
or U16499 (N_16499,N_15707,N_15559);
xor U16500 (N_16500,N_16168,N_16395);
nand U16501 (N_16501,N_16452,N_16137);
nand U16502 (N_16502,N_16025,N_16251);
or U16503 (N_16503,N_16293,N_16208);
or U16504 (N_16504,N_16071,N_16401);
or U16505 (N_16505,N_16441,N_16213);
or U16506 (N_16506,N_16299,N_16338);
nand U16507 (N_16507,N_16450,N_16291);
and U16508 (N_16508,N_16019,N_16434);
or U16509 (N_16509,N_16348,N_16244);
nand U16510 (N_16510,N_16379,N_16473);
and U16511 (N_16511,N_16167,N_16261);
xor U16512 (N_16512,N_16230,N_16009);
or U16513 (N_16513,N_16240,N_16377);
nor U16514 (N_16514,N_16467,N_16023);
or U16515 (N_16515,N_16257,N_16130);
or U16516 (N_16516,N_16346,N_16047);
and U16517 (N_16517,N_16253,N_16409);
and U16518 (N_16518,N_16435,N_16335);
xor U16519 (N_16519,N_16046,N_16172);
nand U16520 (N_16520,N_16022,N_16483);
nor U16521 (N_16521,N_16135,N_16081);
nand U16522 (N_16522,N_16196,N_16454);
and U16523 (N_16523,N_16497,N_16218);
nand U16524 (N_16524,N_16443,N_16316);
nand U16525 (N_16525,N_16292,N_16365);
or U16526 (N_16526,N_16481,N_16021);
xnor U16527 (N_16527,N_16352,N_16459);
nand U16528 (N_16528,N_16495,N_16354);
or U16529 (N_16529,N_16209,N_16212);
and U16530 (N_16530,N_16268,N_16279);
or U16531 (N_16531,N_16110,N_16060);
and U16532 (N_16532,N_16076,N_16033);
nor U16533 (N_16533,N_16256,N_16222);
nand U16534 (N_16534,N_16195,N_16038);
xor U16535 (N_16535,N_16158,N_16223);
nor U16536 (N_16536,N_16187,N_16465);
xor U16537 (N_16537,N_16057,N_16255);
or U16538 (N_16538,N_16082,N_16080);
nor U16539 (N_16539,N_16179,N_16098);
and U16540 (N_16540,N_16095,N_16093);
nand U16541 (N_16541,N_16417,N_16066);
or U16542 (N_16542,N_16312,N_16007);
and U16543 (N_16543,N_16152,N_16103);
nand U16544 (N_16544,N_16091,N_16486);
and U16545 (N_16545,N_16271,N_16433);
or U16546 (N_16546,N_16138,N_16242);
or U16547 (N_16547,N_16034,N_16406);
and U16548 (N_16548,N_16117,N_16421);
nor U16549 (N_16549,N_16400,N_16108);
or U16550 (N_16550,N_16120,N_16224);
and U16551 (N_16551,N_16324,N_16362);
or U16552 (N_16552,N_16074,N_16259);
xnor U16553 (N_16553,N_16493,N_16307);
and U16554 (N_16554,N_16102,N_16429);
xnor U16555 (N_16555,N_16188,N_16451);
nand U16556 (N_16556,N_16418,N_16125);
xor U16557 (N_16557,N_16478,N_16183);
or U16558 (N_16558,N_16144,N_16063);
xnor U16559 (N_16559,N_16380,N_16200);
xnor U16560 (N_16560,N_16479,N_16356);
or U16561 (N_16561,N_16036,N_16457);
or U16562 (N_16562,N_16109,N_16397);
or U16563 (N_16563,N_16373,N_16469);
xnor U16564 (N_16564,N_16001,N_16243);
and U16565 (N_16565,N_16190,N_16105);
or U16566 (N_16566,N_16330,N_16414);
or U16567 (N_16567,N_16068,N_16045);
nor U16568 (N_16568,N_16012,N_16410);
xor U16569 (N_16569,N_16077,N_16037);
nor U16570 (N_16570,N_16048,N_16425);
nor U16571 (N_16571,N_16442,N_16030);
nor U16572 (N_16572,N_16328,N_16482);
and U16573 (N_16573,N_16423,N_16067);
xnor U16574 (N_16574,N_16180,N_16297);
xor U16575 (N_16575,N_16357,N_16315);
and U16576 (N_16576,N_16027,N_16424);
or U16577 (N_16577,N_16258,N_16192);
nand U16578 (N_16578,N_16405,N_16359);
and U16579 (N_16579,N_16083,N_16003);
nor U16580 (N_16580,N_16378,N_16408);
and U16581 (N_16581,N_16387,N_16171);
xnor U16582 (N_16582,N_16126,N_16159);
and U16583 (N_16583,N_16282,N_16078);
nor U16584 (N_16584,N_16136,N_16094);
nand U16585 (N_16585,N_16402,N_16134);
xnor U16586 (N_16586,N_16131,N_16043);
nor U16587 (N_16587,N_16054,N_16000);
nand U16588 (N_16588,N_16403,N_16202);
and U16589 (N_16589,N_16341,N_16194);
nor U16590 (N_16590,N_16461,N_16132);
nand U16591 (N_16591,N_16466,N_16286);
nor U16592 (N_16592,N_16181,N_16308);
and U16593 (N_16593,N_16121,N_16235);
xor U16594 (N_16594,N_16221,N_16439);
and U16595 (N_16595,N_16254,N_16369);
nand U16596 (N_16596,N_16300,N_16332);
or U16597 (N_16597,N_16124,N_16284);
nor U16598 (N_16598,N_16232,N_16347);
nor U16599 (N_16599,N_16203,N_16013);
or U16600 (N_16600,N_16331,N_16295);
or U16601 (N_16601,N_16018,N_16384);
and U16602 (N_16602,N_16388,N_16140);
and U16603 (N_16603,N_16114,N_16236);
and U16604 (N_16604,N_16327,N_16164);
or U16605 (N_16605,N_16290,N_16306);
nand U16606 (N_16606,N_16026,N_16431);
nor U16607 (N_16607,N_16069,N_16129);
xnor U16608 (N_16608,N_16139,N_16337);
nand U16609 (N_16609,N_16028,N_16073);
nor U16610 (N_16610,N_16326,N_16062);
nand U16611 (N_16611,N_16407,N_16173);
and U16612 (N_16612,N_16247,N_16280);
and U16613 (N_16613,N_16170,N_16191);
nand U16614 (N_16614,N_16262,N_16220);
or U16615 (N_16615,N_16283,N_16264);
and U16616 (N_16616,N_16488,N_16107);
nand U16617 (N_16617,N_16151,N_16039);
and U16618 (N_16618,N_16006,N_16149);
nor U16619 (N_16619,N_16155,N_16336);
xor U16620 (N_16620,N_16372,N_16123);
or U16621 (N_16621,N_16368,N_16487);
xnor U16622 (N_16622,N_16396,N_16079);
and U16623 (N_16623,N_16344,N_16288);
and U16624 (N_16624,N_16016,N_16381);
and U16625 (N_16625,N_16175,N_16456);
xnor U16626 (N_16626,N_16474,N_16498);
nor U16627 (N_16627,N_16472,N_16376);
nand U16628 (N_16628,N_16334,N_16128);
nor U16629 (N_16629,N_16165,N_16041);
or U16630 (N_16630,N_16017,N_16374);
nor U16631 (N_16631,N_16070,N_16215);
xor U16632 (N_16632,N_16432,N_16391);
nor U16633 (N_16633,N_16427,N_16186);
nor U16634 (N_16634,N_16176,N_16490);
or U16635 (N_16635,N_16278,N_16345);
and U16636 (N_16636,N_16225,N_16275);
and U16637 (N_16637,N_16339,N_16411);
nand U16638 (N_16638,N_16298,N_16446);
xnor U16639 (N_16639,N_16398,N_16184);
nand U16640 (N_16640,N_16447,N_16445);
and U16641 (N_16641,N_16216,N_16207);
and U16642 (N_16642,N_16484,N_16426);
nand U16643 (N_16643,N_16040,N_16100);
xor U16644 (N_16644,N_16087,N_16383);
xnor U16645 (N_16645,N_16480,N_16106);
nand U16646 (N_16646,N_16499,N_16363);
nor U16647 (N_16647,N_16462,N_16088);
nand U16648 (N_16648,N_16044,N_16342);
or U16649 (N_16649,N_16303,N_16239);
and U16650 (N_16650,N_16096,N_16197);
nand U16651 (N_16651,N_16436,N_16350);
nor U16652 (N_16652,N_16064,N_16325);
and U16653 (N_16653,N_16389,N_16422);
nand U16654 (N_16654,N_16118,N_16148);
and U16655 (N_16655,N_16177,N_16267);
xor U16656 (N_16656,N_16169,N_16189);
and U16657 (N_16657,N_16428,N_16464);
xnor U16658 (N_16658,N_16349,N_16217);
or U16659 (N_16659,N_16246,N_16455);
and U16660 (N_16660,N_16101,N_16049);
nor U16661 (N_16661,N_16210,N_16056);
nor U16662 (N_16662,N_16296,N_16386);
xor U16663 (N_16663,N_16156,N_16153);
nor U16664 (N_16664,N_16182,N_16438);
nand U16665 (N_16665,N_16154,N_16496);
or U16666 (N_16666,N_16305,N_16143);
and U16667 (N_16667,N_16471,N_16227);
nor U16668 (N_16668,N_16231,N_16011);
xnor U16669 (N_16669,N_16437,N_16086);
xor U16670 (N_16670,N_16008,N_16112);
nor U16671 (N_16671,N_16449,N_16249);
xnor U16672 (N_16672,N_16470,N_16343);
nor U16673 (N_16673,N_16382,N_16185);
and U16674 (N_16674,N_16051,N_16444);
xnor U16675 (N_16675,N_16219,N_16020);
nor U16676 (N_16676,N_16150,N_16052);
nand U16677 (N_16677,N_16276,N_16201);
xor U16678 (N_16678,N_16329,N_16104);
xor U16679 (N_16679,N_16274,N_16206);
nand U16680 (N_16680,N_16085,N_16304);
nor U16681 (N_16681,N_16289,N_16214);
nor U16682 (N_16682,N_16002,N_16260);
nand U16683 (N_16683,N_16119,N_16116);
nand U16684 (N_16684,N_16265,N_16463);
nand U16685 (N_16685,N_16413,N_16375);
nand U16686 (N_16686,N_16092,N_16394);
nand U16687 (N_16687,N_16287,N_16309);
xor U16688 (N_16688,N_16485,N_16157);
nand U16689 (N_16689,N_16010,N_16238);
nand U16690 (N_16690,N_16113,N_16333);
nand U16691 (N_16691,N_16353,N_16266);
and U16692 (N_16692,N_16234,N_16166);
nand U16693 (N_16693,N_16491,N_16453);
nand U16694 (N_16694,N_16229,N_16178);
and U16695 (N_16695,N_16412,N_16489);
nand U16696 (N_16696,N_16111,N_16364);
or U16697 (N_16697,N_16174,N_16160);
and U16698 (N_16698,N_16277,N_16321);
and U16699 (N_16699,N_16233,N_16320);
nor U16700 (N_16700,N_16029,N_16351);
or U16701 (N_16701,N_16294,N_16055);
and U16702 (N_16702,N_16285,N_16468);
or U16703 (N_16703,N_16360,N_16237);
and U16704 (N_16704,N_16050,N_16361);
and U16705 (N_16705,N_16317,N_16115);
nor U16706 (N_16706,N_16099,N_16245);
xor U16707 (N_16707,N_16311,N_16031);
xor U16708 (N_16708,N_16024,N_16032);
or U16709 (N_16709,N_16142,N_16263);
nand U16710 (N_16710,N_16211,N_16477);
or U16711 (N_16711,N_16226,N_16015);
and U16712 (N_16712,N_16161,N_16272);
nand U16713 (N_16713,N_16370,N_16042);
and U16714 (N_16714,N_16269,N_16075);
nand U16715 (N_16715,N_16065,N_16313);
and U16716 (N_16716,N_16089,N_16193);
nor U16717 (N_16717,N_16476,N_16385);
nor U16718 (N_16718,N_16228,N_16358);
nand U16719 (N_16719,N_16241,N_16430);
nor U16720 (N_16720,N_16058,N_16273);
nor U16721 (N_16721,N_16133,N_16475);
xor U16722 (N_16722,N_16146,N_16367);
xnor U16723 (N_16723,N_16371,N_16390);
xnor U16724 (N_16724,N_16248,N_16310);
nand U16725 (N_16725,N_16340,N_16355);
xnor U16726 (N_16726,N_16141,N_16319);
xor U16727 (N_16727,N_16415,N_16005);
or U16728 (N_16728,N_16014,N_16392);
and U16729 (N_16729,N_16059,N_16053);
or U16730 (N_16730,N_16163,N_16072);
and U16731 (N_16731,N_16205,N_16145);
or U16732 (N_16732,N_16366,N_16147);
and U16733 (N_16733,N_16302,N_16090);
xnor U16734 (N_16734,N_16281,N_16420);
nand U16735 (N_16735,N_16314,N_16035);
nor U16736 (N_16736,N_16404,N_16270);
xor U16737 (N_16737,N_16448,N_16393);
or U16738 (N_16738,N_16004,N_16061);
or U16739 (N_16739,N_16127,N_16492);
or U16740 (N_16740,N_16204,N_16084);
xnor U16741 (N_16741,N_16250,N_16458);
nor U16742 (N_16742,N_16494,N_16399);
xor U16743 (N_16743,N_16440,N_16323);
nor U16744 (N_16744,N_16252,N_16322);
or U16745 (N_16745,N_16460,N_16162);
nand U16746 (N_16746,N_16318,N_16199);
xnor U16747 (N_16747,N_16198,N_16122);
xor U16748 (N_16748,N_16097,N_16419);
nor U16749 (N_16749,N_16416,N_16301);
xor U16750 (N_16750,N_16251,N_16289);
xnor U16751 (N_16751,N_16037,N_16031);
nor U16752 (N_16752,N_16285,N_16388);
nor U16753 (N_16753,N_16245,N_16279);
nand U16754 (N_16754,N_16181,N_16209);
or U16755 (N_16755,N_16061,N_16443);
nand U16756 (N_16756,N_16439,N_16064);
xor U16757 (N_16757,N_16224,N_16478);
nor U16758 (N_16758,N_16120,N_16282);
xor U16759 (N_16759,N_16179,N_16378);
nor U16760 (N_16760,N_16312,N_16493);
nor U16761 (N_16761,N_16076,N_16259);
and U16762 (N_16762,N_16224,N_16331);
xnor U16763 (N_16763,N_16119,N_16274);
nor U16764 (N_16764,N_16251,N_16104);
xnor U16765 (N_16765,N_16418,N_16002);
and U16766 (N_16766,N_16101,N_16349);
nand U16767 (N_16767,N_16325,N_16089);
xnor U16768 (N_16768,N_16460,N_16488);
or U16769 (N_16769,N_16490,N_16290);
nor U16770 (N_16770,N_16430,N_16072);
xnor U16771 (N_16771,N_16194,N_16113);
xor U16772 (N_16772,N_16035,N_16014);
nor U16773 (N_16773,N_16431,N_16336);
nand U16774 (N_16774,N_16001,N_16337);
nand U16775 (N_16775,N_16132,N_16394);
nor U16776 (N_16776,N_16238,N_16200);
nor U16777 (N_16777,N_16034,N_16443);
xnor U16778 (N_16778,N_16391,N_16008);
and U16779 (N_16779,N_16413,N_16000);
nand U16780 (N_16780,N_16231,N_16243);
or U16781 (N_16781,N_16364,N_16452);
or U16782 (N_16782,N_16192,N_16098);
or U16783 (N_16783,N_16267,N_16217);
nor U16784 (N_16784,N_16041,N_16184);
and U16785 (N_16785,N_16065,N_16025);
xor U16786 (N_16786,N_16389,N_16185);
or U16787 (N_16787,N_16331,N_16336);
and U16788 (N_16788,N_16246,N_16226);
and U16789 (N_16789,N_16136,N_16181);
or U16790 (N_16790,N_16122,N_16182);
nand U16791 (N_16791,N_16411,N_16112);
and U16792 (N_16792,N_16066,N_16421);
or U16793 (N_16793,N_16169,N_16121);
xor U16794 (N_16794,N_16497,N_16181);
xnor U16795 (N_16795,N_16125,N_16039);
nor U16796 (N_16796,N_16411,N_16270);
and U16797 (N_16797,N_16292,N_16170);
xor U16798 (N_16798,N_16284,N_16242);
xor U16799 (N_16799,N_16432,N_16430);
and U16800 (N_16800,N_16381,N_16256);
nor U16801 (N_16801,N_16085,N_16146);
xnor U16802 (N_16802,N_16083,N_16487);
or U16803 (N_16803,N_16172,N_16121);
and U16804 (N_16804,N_16483,N_16214);
and U16805 (N_16805,N_16049,N_16297);
nor U16806 (N_16806,N_16212,N_16281);
or U16807 (N_16807,N_16054,N_16300);
xor U16808 (N_16808,N_16151,N_16358);
xnor U16809 (N_16809,N_16290,N_16176);
nor U16810 (N_16810,N_16275,N_16333);
nand U16811 (N_16811,N_16048,N_16173);
xor U16812 (N_16812,N_16270,N_16167);
xnor U16813 (N_16813,N_16464,N_16370);
xnor U16814 (N_16814,N_16445,N_16004);
or U16815 (N_16815,N_16157,N_16414);
nand U16816 (N_16816,N_16228,N_16414);
nand U16817 (N_16817,N_16161,N_16396);
xnor U16818 (N_16818,N_16320,N_16370);
or U16819 (N_16819,N_16216,N_16024);
and U16820 (N_16820,N_16121,N_16463);
and U16821 (N_16821,N_16300,N_16436);
xor U16822 (N_16822,N_16402,N_16321);
nand U16823 (N_16823,N_16494,N_16473);
and U16824 (N_16824,N_16359,N_16089);
nand U16825 (N_16825,N_16340,N_16190);
nand U16826 (N_16826,N_16459,N_16490);
or U16827 (N_16827,N_16374,N_16262);
nor U16828 (N_16828,N_16032,N_16256);
xor U16829 (N_16829,N_16267,N_16402);
or U16830 (N_16830,N_16082,N_16102);
nor U16831 (N_16831,N_16194,N_16187);
nand U16832 (N_16832,N_16392,N_16275);
or U16833 (N_16833,N_16169,N_16177);
xnor U16834 (N_16834,N_16161,N_16425);
nor U16835 (N_16835,N_16095,N_16203);
nor U16836 (N_16836,N_16264,N_16322);
nor U16837 (N_16837,N_16386,N_16264);
nor U16838 (N_16838,N_16228,N_16336);
xor U16839 (N_16839,N_16001,N_16317);
and U16840 (N_16840,N_16410,N_16152);
nor U16841 (N_16841,N_16112,N_16302);
nor U16842 (N_16842,N_16194,N_16455);
xnor U16843 (N_16843,N_16062,N_16368);
or U16844 (N_16844,N_16117,N_16077);
nor U16845 (N_16845,N_16180,N_16483);
or U16846 (N_16846,N_16025,N_16407);
and U16847 (N_16847,N_16327,N_16196);
nand U16848 (N_16848,N_16118,N_16432);
nor U16849 (N_16849,N_16378,N_16458);
nand U16850 (N_16850,N_16100,N_16399);
nor U16851 (N_16851,N_16228,N_16153);
or U16852 (N_16852,N_16295,N_16126);
xor U16853 (N_16853,N_16344,N_16375);
nor U16854 (N_16854,N_16163,N_16336);
or U16855 (N_16855,N_16180,N_16173);
and U16856 (N_16856,N_16125,N_16379);
nand U16857 (N_16857,N_16408,N_16404);
xnor U16858 (N_16858,N_16171,N_16463);
xor U16859 (N_16859,N_16448,N_16130);
nand U16860 (N_16860,N_16303,N_16021);
nor U16861 (N_16861,N_16124,N_16432);
and U16862 (N_16862,N_16144,N_16338);
or U16863 (N_16863,N_16078,N_16238);
nor U16864 (N_16864,N_16113,N_16124);
xor U16865 (N_16865,N_16344,N_16086);
nand U16866 (N_16866,N_16210,N_16366);
xor U16867 (N_16867,N_16145,N_16218);
nor U16868 (N_16868,N_16017,N_16331);
xnor U16869 (N_16869,N_16082,N_16219);
xnor U16870 (N_16870,N_16349,N_16337);
nand U16871 (N_16871,N_16146,N_16035);
or U16872 (N_16872,N_16083,N_16022);
nor U16873 (N_16873,N_16492,N_16211);
or U16874 (N_16874,N_16230,N_16329);
nor U16875 (N_16875,N_16131,N_16417);
and U16876 (N_16876,N_16137,N_16044);
nor U16877 (N_16877,N_16131,N_16438);
nor U16878 (N_16878,N_16095,N_16447);
nor U16879 (N_16879,N_16063,N_16346);
or U16880 (N_16880,N_16450,N_16231);
and U16881 (N_16881,N_16385,N_16199);
nand U16882 (N_16882,N_16462,N_16459);
nand U16883 (N_16883,N_16425,N_16388);
nor U16884 (N_16884,N_16379,N_16004);
nand U16885 (N_16885,N_16023,N_16000);
or U16886 (N_16886,N_16103,N_16461);
and U16887 (N_16887,N_16336,N_16169);
nand U16888 (N_16888,N_16360,N_16495);
and U16889 (N_16889,N_16369,N_16258);
and U16890 (N_16890,N_16392,N_16220);
nor U16891 (N_16891,N_16489,N_16259);
and U16892 (N_16892,N_16430,N_16285);
or U16893 (N_16893,N_16053,N_16084);
xor U16894 (N_16894,N_16372,N_16091);
xnor U16895 (N_16895,N_16242,N_16190);
or U16896 (N_16896,N_16244,N_16165);
and U16897 (N_16897,N_16086,N_16293);
nor U16898 (N_16898,N_16213,N_16036);
nand U16899 (N_16899,N_16357,N_16448);
and U16900 (N_16900,N_16157,N_16043);
and U16901 (N_16901,N_16161,N_16214);
and U16902 (N_16902,N_16333,N_16366);
nor U16903 (N_16903,N_16324,N_16020);
xor U16904 (N_16904,N_16041,N_16371);
xnor U16905 (N_16905,N_16461,N_16054);
and U16906 (N_16906,N_16149,N_16211);
xnor U16907 (N_16907,N_16172,N_16257);
xor U16908 (N_16908,N_16137,N_16421);
and U16909 (N_16909,N_16065,N_16051);
nor U16910 (N_16910,N_16220,N_16287);
nor U16911 (N_16911,N_16454,N_16053);
nor U16912 (N_16912,N_16333,N_16312);
nand U16913 (N_16913,N_16411,N_16177);
and U16914 (N_16914,N_16145,N_16461);
nand U16915 (N_16915,N_16062,N_16222);
and U16916 (N_16916,N_16069,N_16330);
or U16917 (N_16917,N_16138,N_16260);
or U16918 (N_16918,N_16440,N_16449);
or U16919 (N_16919,N_16064,N_16360);
xnor U16920 (N_16920,N_16345,N_16257);
and U16921 (N_16921,N_16204,N_16019);
xor U16922 (N_16922,N_16196,N_16071);
or U16923 (N_16923,N_16490,N_16389);
and U16924 (N_16924,N_16255,N_16483);
or U16925 (N_16925,N_16445,N_16156);
nand U16926 (N_16926,N_16176,N_16173);
nor U16927 (N_16927,N_16062,N_16278);
xnor U16928 (N_16928,N_16295,N_16435);
nand U16929 (N_16929,N_16132,N_16072);
xnor U16930 (N_16930,N_16049,N_16070);
and U16931 (N_16931,N_16244,N_16059);
nand U16932 (N_16932,N_16109,N_16425);
and U16933 (N_16933,N_16138,N_16346);
xor U16934 (N_16934,N_16298,N_16478);
and U16935 (N_16935,N_16040,N_16381);
xnor U16936 (N_16936,N_16341,N_16004);
nor U16937 (N_16937,N_16429,N_16121);
nor U16938 (N_16938,N_16367,N_16329);
xor U16939 (N_16939,N_16431,N_16266);
or U16940 (N_16940,N_16360,N_16061);
or U16941 (N_16941,N_16242,N_16397);
and U16942 (N_16942,N_16487,N_16110);
nor U16943 (N_16943,N_16385,N_16095);
nor U16944 (N_16944,N_16331,N_16451);
nand U16945 (N_16945,N_16155,N_16361);
and U16946 (N_16946,N_16072,N_16499);
and U16947 (N_16947,N_16479,N_16190);
and U16948 (N_16948,N_16335,N_16206);
or U16949 (N_16949,N_16439,N_16253);
nor U16950 (N_16950,N_16005,N_16162);
xor U16951 (N_16951,N_16383,N_16329);
xnor U16952 (N_16952,N_16366,N_16012);
xnor U16953 (N_16953,N_16357,N_16178);
nor U16954 (N_16954,N_16030,N_16275);
and U16955 (N_16955,N_16279,N_16193);
or U16956 (N_16956,N_16449,N_16470);
nand U16957 (N_16957,N_16199,N_16183);
nor U16958 (N_16958,N_16288,N_16401);
xnor U16959 (N_16959,N_16018,N_16161);
nor U16960 (N_16960,N_16180,N_16283);
or U16961 (N_16961,N_16312,N_16352);
xor U16962 (N_16962,N_16240,N_16165);
or U16963 (N_16963,N_16075,N_16182);
xnor U16964 (N_16964,N_16223,N_16333);
nor U16965 (N_16965,N_16255,N_16116);
nor U16966 (N_16966,N_16036,N_16210);
nor U16967 (N_16967,N_16218,N_16344);
and U16968 (N_16968,N_16153,N_16353);
nor U16969 (N_16969,N_16039,N_16280);
nor U16970 (N_16970,N_16214,N_16484);
nand U16971 (N_16971,N_16045,N_16182);
or U16972 (N_16972,N_16058,N_16378);
nor U16973 (N_16973,N_16449,N_16455);
nor U16974 (N_16974,N_16478,N_16179);
and U16975 (N_16975,N_16045,N_16375);
and U16976 (N_16976,N_16354,N_16273);
nand U16977 (N_16977,N_16458,N_16231);
nand U16978 (N_16978,N_16066,N_16152);
and U16979 (N_16979,N_16046,N_16312);
and U16980 (N_16980,N_16289,N_16309);
xor U16981 (N_16981,N_16069,N_16023);
nand U16982 (N_16982,N_16330,N_16002);
or U16983 (N_16983,N_16470,N_16274);
nand U16984 (N_16984,N_16441,N_16265);
or U16985 (N_16985,N_16330,N_16497);
nand U16986 (N_16986,N_16030,N_16129);
or U16987 (N_16987,N_16400,N_16069);
xnor U16988 (N_16988,N_16134,N_16367);
nor U16989 (N_16989,N_16400,N_16489);
and U16990 (N_16990,N_16041,N_16076);
xnor U16991 (N_16991,N_16225,N_16353);
and U16992 (N_16992,N_16036,N_16440);
nor U16993 (N_16993,N_16045,N_16334);
nand U16994 (N_16994,N_16260,N_16445);
nand U16995 (N_16995,N_16040,N_16042);
nor U16996 (N_16996,N_16307,N_16170);
nand U16997 (N_16997,N_16073,N_16303);
nand U16998 (N_16998,N_16288,N_16284);
xor U16999 (N_16999,N_16127,N_16122);
and U17000 (N_17000,N_16748,N_16988);
nand U17001 (N_17001,N_16896,N_16804);
nor U17002 (N_17002,N_16705,N_16799);
nor U17003 (N_17003,N_16711,N_16826);
nor U17004 (N_17004,N_16907,N_16933);
xnor U17005 (N_17005,N_16681,N_16555);
nor U17006 (N_17006,N_16914,N_16978);
and U17007 (N_17007,N_16842,N_16740);
or U17008 (N_17008,N_16610,N_16834);
or U17009 (N_17009,N_16642,N_16609);
xor U17010 (N_17010,N_16549,N_16708);
or U17011 (N_17011,N_16924,N_16534);
nand U17012 (N_17012,N_16702,N_16682);
xor U17013 (N_17013,N_16593,N_16921);
and U17014 (N_17014,N_16837,N_16672);
xor U17015 (N_17015,N_16501,N_16965);
nand U17016 (N_17016,N_16531,N_16691);
or U17017 (N_17017,N_16538,N_16540);
xnor U17018 (N_17018,N_16923,N_16898);
nor U17019 (N_17019,N_16680,N_16871);
nand U17020 (N_17020,N_16920,N_16951);
or U17021 (N_17021,N_16636,N_16629);
xnor U17022 (N_17022,N_16582,N_16516);
or U17023 (N_17023,N_16692,N_16795);
or U17024 (N_17024,N_16851,N_16675);
and U17025 (N_17025,N_16602,N_16780);
nor U17026 (N_17026,N_16703,N_16628);
nor U17027 (N_17027,N_16752,N_16942);
xnor U17028 (N_17028,N_16743,N_16578);
nor U17029 (N_17029,N_16563,N_16747);
nand U17030 (N_17030,N_16759,N_16706);
nand U17031 (N_17031,N_16828,N_16577);
nor U17032 (N_17032,N_16754,N_16718);
or U17033 (N_17033,N_16627,N_16607);
nor U17034 (N_17034,N_16881,N_16587);
xnor U17035 (N_17035,N_16815,N_16912);
and U17036 (N_17036,N_16996,N_16971);
xor U17037 (N_17037,N_16961,N_16556);
nand U17038 (N_17038,N_16600,N_16806);
and U17039 (N_17039,N_16781,N_16664);
nor U17040 (N_17040,N_16758,N_16882);
xor U17041 (N_17041,N_16696,N_16742);
nor U17042 (N_17042,N_16635,N_16821);
and U17043 (N_17043,N_16559,N_16950);
or U17044 (N_17044,N_16713,N_16764);
or U17045 (N_17045,N_16503,N_16619);
nor U17046 (N_17046,N_16878,N_16760);
nand U17047 (N_17047,N_16707,N_16542);
nand U17048 (N_17048,N_16909,N_16983);
or U17049 (N_17049,N_16919,N_16990);
and U17050 (N_17050,N_16852,N_16993);
and U17051 (N_17051,N_16822,N_16512);
xnor U17052 (N_17052,N_16601,N_16893);
nor U17053 (N_17053,N_16551,N_16906);
and U17054 (N_17054,N_16856,N_16813);
nor U17055 (N_17055,N_16865,N_16997);
or U17056 (N_17056,N_16550,N_16622);
and U17057 (N_17057,N_16880,N_16830);
nand U17058 (N_17058,N_16645,N_16657);
xor U17059 (N_17059,N_16836,N_16753);
xor U17060 (N_17060,N_16571,N_16962);
nor U17061 (N_17061,N_16520,N_16947);
xor U17062 (N_17062,N_16676,N_16825);
nor U17063 (N_17063,N_16980,N_16528);
and U17064 (N_17064,N_16522,N_16803);
and U17065 (N_17065,N_16569,N_16631);
nor U17066 (N_17066,N_16514,N_16784);
nor U17067 (N_17067,N_16669,N_16936);
nor U17068 (N_17068,N_16573,N_16546);
nor U17069 (N_17069,N_16566,N_16615);
xnor U17070 (N_17070,N_16592,N_16938);
and U17071 (N_17071,N_16776,N_16637);
or U17072 (N_17072,N_16952,N_16969);
nand U17073 (N_17073,N_16889,N_16934);
nand U17074 (N_17074,N_16727,N_16908);
and U17075 (N_17075,N_16886,N_16500);
xnor U17076 (N_17076,N_16583,N_16720);
nand U17077 (N_17077,N_16598,N_16586);
xor U17078 (N_17078,N_16770,N_16979);
nand U17079 (N_17079,N_16626,N_16508);
nand U17080 (N_17080,N_16732,N_16939);
and U17081 (N_17081,N_16879,N_16771);
nand U17082 (N_17082,N_16543,N_16721);
and U17083 (N_17083,N_16839,N_16917);
and U17084 (N_17084,N_16639,N_16630);
and U17085 (N_17085,N_16509,N_16956);
xor U17086 (N_17086,N_16548,N_16562);
and U17087 (N_17087,N_16940,N_16810);
nor U17088 (N_17088,N_16957,N_16552);
xnor U17089 (N_17089,N_16994,N_16794);
nand U17090 (N_17090,N_16517,N_16717);
nand U17091 (N_17091,N_16521,N_16589);
and U17092 (N_17092,N_16633,N_16701);
and U17093 (N_17093,N_16590,N_16820);
xor U17094 (N_17094,N_16649,N_16805);
nor U17095 (N_17095,N_16975,N_16526);
and U17096 (N_17096,N_16674,N_16973);
or U17097 (N_17097,N_16850,N_16812);
xor U17098 (N_17098,N_16808,N_16722);
nand U17099 (N_17099,N_16605,N_16643);
and U17100 (N_17100,N_16561,N_16801);
nor U17101 (N_17101,N_16787,N_16591);
nand U17102 (N_17102,N_16741,N_16737);
or U17103 (N_17103,N_16665,N_16790);
or U17104 (N_17104,N_16868,N_16558);
nand U17105 (N_17105,N_16554,N_16927);
or U17106 (N_17106,N_16576,N_16838);
nor U17107 (N_17107,N_16855,N_16944);
xor U17108 (N_17108,N_16960,N_16567);
and U17109 (N_17109,N_16782,N_16966);
xor U17110 (N_17110,N_16824,N_16710);
and U17111 (N_17111,N_16854,N_16505);
and U17112 (N_17112,N_16697,N_16716);
or U17113 (N_17113,N_16553,N_16861);
nor U17114 (N_17114,N_16513,N_16831);
nor U17115 (N_17115,N_16928,N_16900);
nor U17116 (N_17116,N_16651,N_16890);
and U17117 (N_17117,N_16719,N_16653);
or U17118 (N_17118,N_16876,N_16809);
nor U17119 (N_17119,N_16902,N_16685);
xor U17120 (N_17120,N_16584,N_16945);
nor U17121 (N_17121,N_16866,N_16925);
and U17122 (N_17122,N_16547,N_16926);
nand U17123 (N_17123,N_16624,N_16800);
or U17124 (N_17124,N_16901,N_16905);
nor U17125 (N_17125,N_16617,N_16964);
xnor U17126 (N_17126,N_16730,N_16572);
xor U17127 (N_17127,N_16954,N_16768);
and U17128 (N_17128,N_16734,N_16857);
or U17129 (N_17129,N_16744,N_16725);
and U17130 (N_17130,N_16967,N_16527);
nand U17131 (N_17131,N_16606,N_16991);
or U17132 (N_17132,N_16666,N_16791);
or U17133 (N_17133,N_16916,N_16818);
and U17134 (N_17134,N_16510,N_16504);
nand U17135 (N_17135,N_16678,N_16723);
nand U17136 (N_17136,N_16767,N_16858);
nor U17137 (N_17137,N_16904,N_16564);
and U17138 (N_17138,N_16658,N_16798);
nand U17139 (N_17139,N_16603,N_16887);
nand U17140 (N_17140,N_16875,N_16999);
nor U17141 (N_17141,N_16621,N_16731);
or U17142 (N_17142,N_16982,N_16786);
or U17143 (N_17143,N_16544,N_16574);
xor U17144 (N_17144,N_16668,N_16968);
xnor U17145 (N_17145,N_16931,N_16937);
nand U17146 (N_17146,N_16918,N_16756);
nand U17147 (N_17147,N_16565,N_16844);
nand U17148 (N_17148,N_16816,N_16958);
or U17149 (N_17149,N_16539,N_16714);
and U17150 (N_17150,N_16557,N_16888);
or U17151 (N_17151,N_16864,N_16656);
nor U17152 (N_17152,N_16652,N_16618);
xnor U17153 (N_17153,N_16829,N_16763);
xnor U17154 (N_17154,N_16634,N_16532);
or U17155 (N_17155,N_16833,N_16699);
and U17156 (N_17156,N_16814,N_16762);
nor U17157 (N_17157,N_16775,N_16729);
or U17158 (N_17158,N_16683,N_16827);
or U17159 (N_17159,N_16687,N_16661);
nor U17160 (N_17160,N_16935,N_16894);
nand U17161 (N_17161,N_16910,N_16644);
xor U17162 (N_17162,N_16523,N_16646);
nand U17163 (N_17163,N_16774,N_16783);
nand U17164 (N_17164,N_16613,N_16872);
and U17165 (N_17165,N_16533,N_16673);
nand U17166 (N_17166,N_16860,N_16765);
and U17167 (N_17167,N_16671,N_16612);
or U17168 (N_17168,N_16853,N_16823);
nand U17169 (N_17169,N_16728,N_16611);
xor U17170 (N_17170,N_16797,N_16654);
or U17171 (N_17171,N_16884,N_16745);
nand U17172 (N_17172,N_16545,N_16941);
or U17173 (N_17173,N_16874,N_16616);
or U17174 (N_17174,N_16751,N_16739);
xnor U17175 (N_17175,N_16746,N_16625);
nor U17176 (N_17176,N_16955,N_16761);
xor U17177 (N_17177,N_16594,N_16749);
nor U17178 (N_17178,N_16655,N_16848);
and U17179 (N_17179,N_16529,N_16862);
or U17180 (N_17180,N_16614,N_16849);
and U17181 (N_17181,N_16677,N_16632);
and U17182 (N_17182,N_16981,N_16647);
and U17183 (N_17183,N_16502,N_16972);
nand U17184 (N_17184,N_16623,N_16793);
nor U17185 (N_17185,N_16873,N_16985);
xor U17186 (N_17186,N_16579,N_16897);
nand U17187 (N_17187,N_16946,N_16769);
and U17188 (N_17188,N_16779,N_16974);
or U17189 (N_17189,N_16995,N_16688);
or U17190 (N_17190,N_16929,N_16693);
or U17191 (N_17191,N_16596,N_16998);
or U17192 (N_17192,N_16686,N_16959);
xor U17193 (N_17193,N_16953,N_16840);
xor U17194 (N_17194,N_16733,N_16883);
and U17195 (N_17195,N_16949,N_16511);
nand U17196 (N_17196,N_16690,N_16575);
xnor U17197 (N_17197,N_16620,N_16835);
xor U17198 (N_17198,N_16895,N_16989);
nor U17199 (N_17199,N_16537,N_16515);
xnor U17200 (N_17200,N_16891,N_16641);
xor U17201 (N_17201,N_16506,N_16659);
nand U17202 (N_17202,N_16715,N_16662);
nor U17203 (N_17203,N_16541,N_16986);
nor U17204 (N_17204,N_16976,N_16585);
nand U17205 (N_17205,N_16788,N_16846);
or U17206 (N_17206,N_16913,N_16698);
nor U17207 (N_17207,N_16963,N_16597);
xnor U17208 (N_17208,N_16670,N_16599);
or U17209 (N_17209,N_16604,N_16738);
and U17210 (N_17210,N_16660,N_16712);
and U17211 (N_17211,N_16518,N_16694);
and U17212 (N_17212,N_16867,N_16581);
and U17213 (N_17213,N_16847,N_16977);
and U17214 (N_17214,N_16892,N_16588);
or U17215 (N_17215,N_16560,N_16802);
xor U17216 (N_17216,N_16750,N_16736);
nor U17217 (N_17217,N_16525,N_16755);
or U17218 (N_17218,N_16859,N_16885);
nand U17219 (N_17219,N_16899,N_16772);
nand U17220 (N_17220,N_16817,N_16789);
xnor U17221 (N_17221,N_16757,N_16843);
and U17222 (N_17222,N_16869,N_16984);
xor U17223 (N_17223,N_16679,N_16667);
nor U17224 (N_17224,N_16841,N_16519);
and U17225 (N_17225,N_16877,N_16663);
and U17226 (N_17226,N_16992,N_16700);
nand U17227 (N_17227,N_16948,N_16640);
or U17228 (N_17228,N_16684,N_16773);
and U17229 (N_17229,N_16570,N_16970);
and U17230 (N_17230,N_16922,N_16580);
xor U17231 (N_17231,N_16792,N_16689);
and U17232 (N_17232,N_16811,N_16807);
and U17233 (N_17233,N_16695,N_16735);
xnor U17234 (N_17234,N_16930,N_16819);
nand U17235 (N_17235,N_16704,N_16568);
or U17236 (N_17236,N_16536,N_16863);
and U17237 (N_17237,N_16766,N_16903);
xnor U17238 (N_17238,N_16911,N_16726);
nor U17239 (N_17239,N_16796,N_16778);
xnor U17240 (N_17240,N_16943,N_16524);
or U17241 (N_17241,N_16870,N_16638);
or U17242 (N_17242,N_16932,N_16507);
xnor U17243 (N_17243,N_16785,N_16650);
or U17244 (N_17244,N_16595,N_16608);
nand U17245 (N_17245,N_16777,N_16832);
nand U17246 (N_17246,N_16915,N_16709);
nor U17247 (N_17247,N_16530,N_16648);
nand U17248 (N_17248,N_16724,N_16535);
xnor U17249 (N_17249,N_16845,N_16987);
nor U17250 (N_17250,N_16510,N_16599);
xnor U17251 (N_17251,N_16763,N_16804);
nand U17252 (N_17252,N_16844,N_16891);
or U17253 (N_17253,N_16676,N_16757);
nand U17254 (N_17254,N_16513,N_16925);
or U17255 (N_17255,N_16720,N_16667);
or U17256 (N_17256,N_16878,N_16738);
nor U17257 (N_17257,N_16633,N_16788);
and U17258 (N_17258,N_16729,N_16950);
xnor U17259 (N_17259,N_16886,N_16597);
nor U17260 (N_17260,N_16935,N_16527);
and U17261 (N_17261,N_16830,N_16540);
or U17262 (N_17262,N_16844,N_16518);
or U17263 (N_17263,N_16603,N_16642);
and U17264 (N_17264,N_16541,N_16916);
and U17265 (N_17265,N_16655,N_16592);
and U17266 (N_17266,N_16956,N_16991);
nor U17267 (N_17267,N_16961,N_16771);
and U17268 (N_17268,N_16695,N_16977);
or U17269 (N_17269,N_16593,N_16963);
and U17270 (N_17270,N_16933,N_16671);
xor U17271 (N_17271,N_16984,N_16767);
nand U17272 (N_17272,N_16994,N_16863);
nand U17273 (N_17273,N_16894,N_16751);
and U17274 (N_17274,N_16628,N_16716);
or U17275 (N_17275,N_16812,N_16701);
and U17276 (N_17276,N_16882,N_16748);
nor U17277 (N_17277,N_16710,N_16623);
or U17278 (N_17278,N_16881,N_16991);
nor U17279 (N_17279,N_16573,N_16868);
nand U17280 (N_17280,N_16764,N_16579);
nand U17281 (N_17281,N_16567,N_16715);
nor U17282 (N_17282,N_16561,N_16779);
xor U17283 (N_17283,N_16501,N_16637);
and U17284 (N_17284,N_16661,N_16595);
xor U17285 (N_17285,N_16647,N_16950);
nand U17286 (N_17286,N_16981,N_16761);
or U17287 (N_17287,N_16910,N_16741);
xor U17288 (N_17288,N_16528,N_16824);
nor U17289 (N_17289,N_16674,N_16649);
nand U17290 (N_17290,N_16696,N_16870);
and U17291 (N_17291,N_16842,N_16871);
xor U17292 (N_17292,N_16987,N_16603);
or U17293 (N_17293,N_16933,N_16968);
and U17294 (N_17294,N_16782,N_16625);
nor U17295 (N_17295,N_16667,N_16748);
and U17296 (N_17296,N_16686,N_16677);
nand U17297 (N_17297,N_16605,N_16530);
xor U17298 (N_17298,N_16946,N_16898);
and U17299 (N_17299,N_16531,N_16519);
nor U17300 (N_17300,N_16857,N_16939);
nand U17301 (N_17301,N_16834,N_16757);
or U17302 (N_17302,N_16917,N_16604);
xnor U17303 (N_17303,N_16626,N_16953);
xnor U17304 (N_17304,N_16539,N_16835);
or U17305 (N_17305,N_16518,N_16930);
xor U17306 (N_17306,N_16883,N_16751);
or U17307 (N_17307,N_16963,N_16642);
xnor U17308 (N_17308,N_16697,N_16847);
and U17309 (N_17309,N_16827,N_16937);
and U17310 (N_17310,N_16933,N_16680);
and U17311 (N_17311,N_16611,N_16877);
nor U17312 (N_17312,N_16883,N_16660);
xor U17313 (N_17313,N_16846,N_16644);
nand U17314 (N_17314,N_16573,N_16881);
nand U17315 (N_17315,N_16571,N_16613);
and U17316 (N_17316,N_16863,N_16754);
or U17317 (N_17317,N_16765,N_16868);
nor U17318 (N_17318,N_16601,N_16538);
nor U17319 (N_17319,N_16758,N_16805);
and U17320 (N_17320,N_16967,N_16834);
nand U17321 (N_17321,N_16778,N_16545);
nand U17322 (N_17322,N_16680,N_16694);
nand U17323 (N_17323,N_16696,N_16501);
nand U17324 (N_17324,N_16899,N_16970);
or U17325 (N_17325,N_16691,N_16734);
or U17326 (N_17326,N_16540,N_16997);
xnor U17327 (N_17327,N_16678,N_16558);
xnor U17328 (N_17328,N_16645,N_16520);
xor U17329 (N_17329,N_16747,N_16965);
nand U17330 (N_17330,N_16506,N_16633);
nor U17331 (N_17331,N_16745,N_16594);
xor U17332 (N_17332,N_16770,N_16693);
and U17333 (N_17333,N_16833,N_16681);
and U17334 (N_17334,N_16564,N_16666);
or U17335 (N_17335,N_16585,N_16610);
nand U17336 (N_17336,N_16593,N_16742);
and U17337 (N_17337,N_16725,N_16771);
or U17338 (N_17338,N_16509,N_16738);
or U17339 (N_17339,N_16986,N_16628);
or U17340 (N_17340,N_16610,N_16543);
nand U17341 (N_17341,N_16636,N_16632);
xor U17342 (N_17342,N_16637,N_16943);
or U17343 (N_17343,N_16799,N_16775);
and U17344 (N_17344,N_16841,N_16676);
and U17345 (N_17345,N_16670,N_16623);
or U17346 (N_17346,N_16741,N_16619);
and U17347 (N_17347,N_16941,N_16785);
and U17348 (N_17348,N_16875,N_16765);
nor U17349 (N_17349,N_16719,N_16554);
nand U17350 (N_17350,N_16568,N_16867);
nand U17351 (N_17351,N_16657,N_16563);
nand U17352 (N_17352,N_16737,N_16701);
nor U17353 (N_17353,N_16563,N_16699);
nand U17354 (N_17354,N_16943,N_16594);
nand U17355 (N_17355,N_16894,N_16603);
xnor U17356 (N_17356,N_16854,N_16598);
or U17357 (N_17357,N_16681,N_16673);
nor U17358 (N_17358,N_16661,N_16683);
nand U17359 (N_17359,N_16682,N_16522);
xor U17360 (N_17360,N_16836,N_16826);
nor U17361 (N_17361,N_16834,N_16617);
xnor U17362 (N_17362,N_16949,N_16533);
nand U17363 (N_17363,N_16959,N_16820);
nor U17364 (N_17364,N_16666,N_16634);
or U17365 (N_17365,N_16561,N_16895);
nor U17366 (N_17366,N_16942,N_16982);
nor U17367 (N_17367,N_16698,N_16991);
nand U17368 (N_17368,N_16622,N_16735);
nand U17369 (N_17369,N_16719,N_16571);
and U17370 (N_17370,N_16590,N_16840);
and U17371 (N_17371,N_16745,N_16553);
nand U17372 (N_17372,N_16506,N_16776);
and U17373 (N_17373,N_16851,N_16850);
nand U17374 (N_17374,N_16871,N_16774);
nor U17375 (N_17375,N_16966,N_16638);
nor U17376 (N_17376,N_16711,N_16885);
or U17377 (N_17377,N_16588,N_16937);
or U17378 (N_17378,N_16548,N_16782);
and U17379 (N_17379,N_16836,N_16957);
nor U17380 (N_17380,N_16701,N_16919);
or U17381 (N_17381,N_16937,N_16701);
or U17382 (N_17382,N_16959,N_16615);
and U17383 (N_17383,N_16691,N_16698);
nor U17384 (N_17384,N_16974,N_16709);
and U17385 (N_17385,N_16724,N_16815);
nand U17386 (N_17386,N_16930,N_16587);
nand U17387 (N_17387,N_16581,N_16959);
and U17388 (N_17388,N_16844,N_16630);
nor U17389 (N_17389,N_16617,N_16898);
or U17390 (N_17390,N_16625,N_16764);
and U17391 (N_17391,N_16505,N_16693);
nand U17392 (N_17392,N_16695,N_16784);
or U17393 (N_17393,N_16971,N_16830);
nor U17394 (N_17394,N_16595,N_16956);
or U17395 (N_17395,N_16802,N_16572);
xnor U17396 (N_17396,N_16627,N_16628);
nand U17397 (N_17397,N_16758,N_16761);
or U17398 (N_17398,N_16885,N_16817);
nand U17399 (N_17399,N_16549,N_16634);
xnor U17400 (N_17400,N_16888,N_16998);
xnor U17401 (N_17401,N_16591,N_16555);
or U17402 (N_17402,N_16655,N_16562);
nor U17403 (N_17403,N_16799,N_16990);
nor U17404 (N_17404,N_16645,N_16741);
and U17405 (N_17405,N_16771,N_16694);
nand U17406 (N_17406,N_16803,N_16977);
nand U17407 (N_17407,N_16722,N_16872);
xnor U17408 (N_17408,N_16618,N_16627);
nor U17409 (N_17409,N_16779,N_16877);
nand U17410 (N_17410,N_16853,N_16777);
nor U17411 (N_17411,N_16853,N_16595);
xnor U17412 (N_17412,N_16732,N_16854);
nand U17413 (N_17413,N_16735,N_16613);
or U17414 (N_17414,N_16672,N_16824);
nor U17415 (N_17415,N_16603,N_16848);
xor U17416 (N_17416,N_16806,N_16930);
and U17417 (N_17417,N_16611,N_16655);
xnor U17418 (N_17418,N_16670,N_16893);
nor U17419 (N_17419,N_16555,N_16510);
nand U17420 (N_17420,N_16565,N_16610);
or U17421 (N_17421,N_16548,N_16997);
nand U17422 (N_17422,N_16685,N_16858);
or U17423 (N_17423,N_16724,N_16905);
nor U17424 (N_17424,N_16652,N_16918);
nand U17425 (N_17425,N_16803,N_16996);
or U17426 (N_17426,N_16927,N_16802);
xor U17427 (N_17427,N_16969,N_16922);
and U17428 (N_17428,N_16970,N_16790);
and U17429 (N_17429,N_16887,N_16944);
or U17430 (N_17430,N_16577,N_16818);
nand U17431 (N_17431,N_16663,N_16724);
nand U17432 (N_17432,N_16943,N_16810);
or U17433 (N_17433,N_16900,N_16818);
nor U17434 (N_17434,N_16642,N_16974);
nor U17435 (N_17435,N_16532,N_16937);
and U17436 (N_17436,N_16507,N_16606);
or U17437 (N_17437,N_16935,N_16640);
and U17438 (N_17438,N_16993,N_16761);
or U17439 (N_17439,N_16717,N_16918);
xnor U17440 (N_17440,N_16934,N_16592);
nor U17441 (N_17441,N_16947,N_16721);
nand U17442 (N_17442,N_16786,N_16827);
and U17443 (N_17443,N_16565,N_16523);
and U17444 (N_17444,N_16959,N_16771);
nand U17445 (N_17445,N_16571,N_16814);
nand U17446 (N_17446,N_16685,N_16609);
and U17447 (N_17447,N_16742,N_16627);
or U17448 (N_17448,N_16788,N_16908);
nand U17449 (N_17449,N_16502,N_16738);
nand U17450 (N_17450,N_16561,N_16954);
and U17451 (N_17451,N_16852,N_16986);
nand U17452 (N_17452,N_16599,N_16990);
nor U17453 (N_17453,N_16908,N_16558);
xor U17454 (N_17454,N_16502,N_16814);
or U17455 (N_17455,N_16894,N_16599);
and U17456 (N_17456,N_16951,N_16704);
nor U17457 (N_17457,N_16867,N_16855);
or U17458 (N_17458,N_16549,N_16702);
xnor U17459 (N_17459,N_16732,N_16615);
or U17460 (N_17460,N_16800,N_16575);
and U17461 (N_17461,N_16926,N_16731);
or U17462 (N_17462,N_16761,N_16987);
or U17463 (N_17463,N_16587,N_16580);
nand U17464 (N_17464,N_16866,N_16900);
xnor U17465 (N_17465,N_16839,N_16728);
xor U17466 (N_17466,N_16718,N_16828);
and U17467 (N_17467,N_16564,N_16801);
and U17468 (N_17468,N_16943,N_16852);
or U17469 (N_17469,N_16889,N_16690);
nor U17470 (N_17470,N_16582,N_16733);
or U17471 (N_17471,N_16535,N_16726);
nand U17472 (N_17472,N_16675,N_16540);
nor U17473 (N_17473,N_16557,N_16736);
nand U17474 (N_17474,N_16611,N_16910);
and U17475 (N_17475,N_16611,N_16746);
nand U17476 (N_17476,N_16663,N_16938);
xor U17477 (N_17477,N_16757,N_16635);
nand U17478 (N_17478,N_16775,N_16963);
and U17479 (N_17479,N_16673,N_16585);
nand U17480 (N_17480,N_16836,N_16560);
nor U17481 (N_17481,N_16624,N_16994);
nor U17482 (N_17482,N_16705,N_16780);
and U17483 (N_17483,N_16629,N_16795);
and U17484 (N_17484,N_16706,N_16572);
or U17485 (N_17485,N_16996,N_16815);
nand U17486 (N_17486,N_16505,N_16930);
or U17487 (N_17487,N_16573,N_16520);
nand U17488 (N_17488,N_16776,N_16675);
or U17489 (N_17489,N_16635,N_16693);
and U17490 (N_17490,N_16871,N_16552);
and U17491 (N_17491,N_16973,N_16672);
nor U17492 (N_17492,N_16929,N_16615);
or U17493 (N_17493,N_16521,N_16954);
and U17494 (N_17494,N_16952,N_16974);
xor U17495 (N_17495,N_16603,N_16711);
nand U17496 (N_17496,N_16919,N_16874);
nand U17497 (N_17497,N_16508,N_16907);
or U17498 (N_17498,N_16526,N_16680);
nor U17499 (N_17499,N_16910,N_16944);
nor U17500 (N_17500,N_17389,N_17419);
nor U17501 (N_17501,N_17217,N_17480);
and U17502 (N_17502,N_17344,N_17372);
nand U17503 (N_17503,N_17256,N_17357);
and U17504 (N_17504,N_17338,N_17122);
or U17505 (N_17505,N_17317,N_17220);
xor U17506 (N_17506,N_17386,N_17064);
and U17507 (N_17507,N_17424,N_17490);
and U17508 (N_17508,N_17112,N_17315);
and U17509 (N_17509,N_17226,N_17165);
nor U17510 (N_17510,N_17164,N_17396);
xnor U17511 (N_17511,N_17432,N_17313);
nand U17512 (N_17512,N_17002,N_17343);
or U17513 (N_17513,N_17113,N_17285);
or U17514 (N_17514,N_17463,N_17061);
nand U17515 (N_17515,N_17376,N_17416);
and U17516 (N_17516,N_17465,N_17262);
or U17517 (N_17517,N_17144,N_17489);
xnor U17518 (N_17518,N_17379,N_17231);
or U17519 (N_17519,N_17260,N_17156);
xnor U17520 (N_17520,N_17092,N_17019);
and U17521 (N_17521,N_17446,N_17183);
and U17522 (N_17522,N_17137,N_17460);
and U17523 (N_17523,N_17194,N_17373);
nand U17524 (N_17524,N_17232,N_17402);
xor U17525 (N_17525,N_17336,N_17190);
and U17526 (N_17526,N_17129,N_17299);
nor U17527 (N_17527,N_17420,N_17401);
and U17528 (N_17528,N_17210,N_17351);
xor U17529 (N_17529,N_17417,N_17304);
or U17530 (N_17530,N_17076,N_17230);
or U17531 (N_17531,N_17366,N_17300);
or U17532 (N_17532,N_17205,N_17244);
or U17533 (N_17533,N_17020,N_17038);
or U17534 (N_17534,N_17058,N_17130);
xnor U17535 (N_17535,N_17105,N_17314);
nand U17536 (N_17536,N_17140,N_17128);
xor U17537 (N_17537,N_17335,N_17282);
nand U17538 (N_17538,N_17108,N_17119);
and U17539 (N_17539,N_17384,N_17004);
xnor U17540 (N_17540,N_17451,N_17223);
and U17541 (N_17541,N_17136,N_17201);
nand U17542 (N_17542,N_17032,N_17365);
nor U17543 (N_17543,N_17184,N_17268);
or U17544 (N_17544,N_17007,N_17455);
nor U17545 (N_17545,N_17481,N_17425);
and U17546 (N_17546,N_17118,N_17153);
and U17547 (N_17547,N_17196,N_17193);
and U17548 (N_17548,N_17187,N_17227);
nand U17549 (N_17549,N_17388,N_17134);
nor U17550 (N_17550,N_17464,N_17155);
nand U17551 (N_17551,N_17272,N_17361);
nand U17552 (N_17552,N_17022,N_17025);
or U17553 (N_17553,N_17492,N_17041);
xor U17554 (N_17554,N_17470,N_17078);
and U17555 (N_17555,N_17243,N_17052);
xor U17556 (N_17556,N_17293,N_17473);
xnor U17557 (N_17557,N_17043,N_17498);
nand U17558 (N_17558,N_17375,N_17408);
or U17559 (N_17559,N_17218,N_17222);
nor U17560 (N_17560,N_17253,N_17409);
nor U17561 (N_17561,N_17281,N_17482);
nand U17562 (N_17562,N_17199,N_17477);
or U17563 (N_17563,N_17069,N_17269);
and U17564 (N_17564,N_17143,N_17146);
nor U17565 (N_17565,N_17127,N_17307);
nor U17566 (N_17566,N_17319,N_17279);
xor U17567 (N_17567,N_17060,N_17162);
nand U17568 (N_17568,N_17035,N_17147);
nand U17569 (N_17569,N_17342,N_17016);
nor U17570 (N_17570,N_17181,N_17085);
and U17571 (N_17571,N_17255,N_17192);
nor U17572 (N_17572,N_17132,N_17459);
and U17573 (N_17573,N_17185,N_17170);
or U17574 (N_17574,N_17142,N_17059);
xor U17575 (N_17575,N_17436,N_17221);
nor U17576 (N_17576,N_17213,N_17330);
and U17577 (N_17577,N_17415,N_17188);
xnor U17578 (N_17578,N_17021,N_17042);
nand U17579 (N_17579,N_17476,N_17349);
nor U17580 (N_17580,N_17249,N_17400);
xor U17581 (N_17581,N_17487,N_17467);
nand U17582 (N_17582,N_17242,N_17399);
or U17583 (N_17583,N_17421,N_17246);
or U17584 (N_17584,N_17318,N_17003);
and U17585 (N_17585,N_17278,N_17149);
xor U17586 (N_17586,N_17067,N_17308);
xor U17587 (N_17587,N_17006,N_17305);
xor U17588 (N_17588,N_17385,N_17054);
or U17589 (N_17589,N_17195,N_17339);
nand U17590 (N_17590,N_17238,N_17423);
xnor U17591 (N_17591,N_17018,N_17271);
xor U17592 (N_17592,N_17056,N_17049);
or U17593 (N_17593,N_17493,N_17478);
and U17594 (N_17594,N_17013,N_17131);
nand U17595 (N_17595,N_17448,N_17345);
nor U17596 (N_17596,N_17378,N_17090);
nand U17597 (N_17597,N_17074,N_17405);
or U17598 (N_17598,N_17011,N_17453);
or U17599 (N_17599,N_17206,N_17332);
nand U17600 (N_17600,N_17179,N_17086);
or U17601 (N_17601,N_17250,N_17191);
nand U17602 (N_17602,N_17053,N_17494);
nand U17603 (N_17603,N_17368,N_17075);
or U17604 (N_17604,N_17100,N_17241);
nand U17605 (N_17605,N_17261,N_17287);
and U17606 (N_17606,N_17440,N_17148);
nand U17607 (N_17607,N_17302,N_17447);
xor U17608 (N_17608,N_17333,N_17234);
or U17609 (N_17609,N_17087,N_17320);
xor U17610 (N_17610,N_17177,N_17387);
xor U17611 (N_17611,N_17171,N_17496);
or U17612 (N_17612,N_17203,N_17139);
nor U17613 (N_17613,N_17167,N_17257);
and U17614 (N_17614,N_17166,N_17207);
xor U17615 (N_17615,N_17267,N_17427);
xor U17616 (N_17616,N_17363,N_17353);
or U17617 (N_17617,N_17120,N_17469);
nand U17618 (N_17618,N_17175,N_17150);
xor U17619 (N_17619,N_17160,N_17377);
nand U17620 (N_17620,N_17245,N_17104);
and U17621 (N_17621,N_17010,N_17418);
nand U17622 (N_17622,N_17334,N_17431);
and U17623 (N_17623,N_17347,N_17173);
xor U17624 (N_17624,N_17495,N_17450);
nor U17625 (N_17625,N_17098,N_17371);
nor U17626 (N_17626,N_17110,N_17099);
or U17627 (N_17627,N_17286,N_17029);
nor U17628 (N_17628,N_17356,N_17340);
nor U17629 (N_17629,N_17324,N_17121);
or U17630 (N_17630,N_17024,N_17133);
nand U17631 (N_17631,N_17277,N_17039);
nand U17632 (N_17632,N_17101,N_17204);
nand U17633 (N_17633,N_17176,N_17198);
nand U17634 (N_17634,N_17102,N_17044);
xor U17635 (N_17635,N_17264,N_17224);
and U17636 (N_17636,N_17380,N_17283);
xnor U17637 (N_17637,N_17089,N_17433);
or U17638 (N_17638,N_17066,N_17251);
xor U17639 (N_17639,N_17051,N_17406);
or U17640 (N_17640,N_17135,N_17301);
or U17641 (N_17641,N_17145,N_17115);
xnor U17642 (N_17642,N_17040,N_17298);
xnor U17643 (N_17643,N_17214,N_17017);
xnor U17644 (N_17644,N_17458,N_17471);
and U17645 (N_17645,N_17093,N_17325);
or U17646 (N_17646,N_17082,N_17070);
xnor U17647 (N_17647,N_17352,N_17117);
nand U17648 (N_17648,N_17483,N_17275);
or U17649 (N_17649,N_17397,N_17321);
nand U17650 (N_17650,N_17186,N_17452);
or U17651 (N_17651,N_17284,N_17252);
or U17652 (N_17652,N_17172,N_17328);
or U17653 (N_17653,N_17354,N_17466);
nand U17654 (N_17654,N_17096,N_17084);
nand U17655 (N_17655,N_17414,N_17383);
nand U17656 (N_17656,N_17012,N_17296);
xor U17657 (N_17657,N_17265,N_17323);
nor U17658 (N_17658,N_17337,N_17233);
nand U17659 (N_17659,N_17410,N_17240);
or U17660 (N_17660,N_17393,N_17499);
and U17661 (N_17661,N_17216,N_17445);
nor U17662 (N_17662,N_17370,N_17292);
and U17663 (N_17663,N_17157,N_17033);
and U17664 (N_17664,N_17229,N_17331);
xnor U17665 (N_17665,N_17141,N_17063);
and U17666 (N_17666,N_17374,N_17030);
xnor U17667 (N_17667,N_17291,N_17106);
nor U17668 (N_17668,N_17200,N_17441);
xor U17669 (N_17669,N_17407,N_17014);
or U17670 (N_17670,N_17312,N_17273);
and U17671 (N_17671,N_17168,N_17348);
or U17672 (N_17672,N_17097,N_17479);
xnor U17673 (N_17673,N_17404,N_17116);
xor U17674 (N_17674,N_17202,N_17239);
nor U17675 (N_17675,N_17247,N_17047);
nor U17676 (N_17676,N_17077,N_17472);
xnor U17677 (N_17677,N_17485,N_17322);
nor U17678 (N_17678,N_17174,N_17484);
nand U17679 (N_17679,N_17208,N_17395);
and U17680 (N_17680,N_17444,N_17457);
xor U17681 (N_17681,N_17215,N_17235);
and U17682 (N_17682,N_17364,N_17057);
nor U17683 (N_17683,N_17182,N_17350);
and U17684 (N_17684,N_17071,N_17329);
nand U17685 (N_17685,N_17088,N_17091);
and U17686 (N_17686,N_17094,N_17326);
or U17687 (N_17687,N_17026,N_17412);
or U17688 (N_17688,N_17248,N_17189);
xnor U17689 (N_17689,N_17468,N_17311);
nor U17690 (N_17690,N_17028,N_17274);
nand U17691 (N_17691,N_17114,N_17398);
nand U17692 (N_17692,N_17341,N_17327);
or U17693 (N_17693,N_17358,N_17394);
or U17694 (N_17694,N_17295,N_17083);
or U17695 (N_17695,N_17095,N_17456);
and U17696 (N_17696,N_17294,N_17443);
or U17697 (N_17697,N_17454,N_17360);
nand U17698 (N_17698,N_17125,N_17355);
nand U17699 (N_17699,N_17236,N_17306);
nor U17700 (N_17700,N_17225,N_17000);
or U17701 (N_17701,N_17392,N_17434);
nand U17702 (N_17702,N_17288,N_17316);
and U17703 (N_17703,N_17266,N_17212);
and U17704 (N_17704,N_17126,N_17048);
xnor U17705 (N_17705,N_17023,N_17062);
or U17706 (N_17706,N_17346,N_17045);
xor U17707 (N_17707,N_17411,N_17034);
xor U17708 (N_17708,N_17237,N_17037);
or U17709 (N_17709,N_17209,N_17228);
nor U17710 (N_17710,N_17442,N_17031);
nand U17711 (N_17711,N_17362,N_17439);
and U17712 (N_17712,N_17163,N_17429);
or U17713 (N_17713,N_17065,N_17310);
or U17714 (N_17714,N_17280,N_17359);
nor U17715 (N_17715,N_17367,N_17254);
or U17716 (N_17716,N_17123,N_17462);
and U17717 (N_17717,N_17259,N_17152);
xor U17718 (N_17718,N_17297,N_17263);
and U17719 (N_17719,N_17497,N_17159);
nor U17720 (N_17720,N_17124,N_17008);
nor U17721 (N_17721,N_17461,N_17055);
and U17722 (N_17722,N_17276,N_17413);
and U17723 (N_17723,N_17435,N_17474);
xnor U17724 (N_17724,N_17391,N_17303);
nor U17725 (N_17725,N_17369,N_17027);
or U17726 (N_17726,N_17151,N_17449);
or U17727 (N_17727,N_17197,N_17403);
nor U17728 (N_17728,N_17158,N_17079);
xor U17729 (N_17729,N_17178,N_17050);
nand U17730 (N_17730,N_17390,N_17015);
nand U17731 (N_17731,N_17488,N_17426);
or U17732 (N_17732,N_17154,N_17211);
and U17733 (N_17733,N_17138,N_17107);
and U17734 (N_17734,N_17080,N_17073);
nand U17735 (N_17735,N_17309,N_17491);
nor U17736 (N_17736,N_17068,N_17290);
nand U17737 (N_17737,N_17081,N_17270);
and U17738 (N_17738,N_17103,N_17169);
nor U17739 (N_17739,N_17219,N_17437);
xnor U17740 (N_17740,N_17005,N_17180);
nor U17741 (N_17741,N_17161,N_17486);
or U17742 (N_17742,N_17001,N_17438);
or U17743 (N_17743,N_17428,N_17046);
nand U17744 (N_17744,N_17382,N_17258);
xor U17745 (N_17745,N_17381,N_17289);
or U17746 (N_17746,N_17036,N_17422);
and U17747 (N_17747,N_17430,N_17475);
xnor U17748 (N_17748,N_17009,N_17072);
nand U17749 (N_17749,N_17111,N_17109);
nor U17750 (N_17750,N_17490,N_17014);
or U17751 (N_17751,N_17208,N_17365);
or U17752 (N_17752,N_17311,N_17481);
or U17753 (N_17753,N_17034,N_17212);
xnor U17754 (N_17754,N_17484,N_17249);
or U17755 (N_17755,N_17097,N_17344);
nor U17756 (N_17756,N_17140,N_17087);
nor U17757 (N_17757,N_17241,N_17315);
and U17758 (N_17758,N_17127,N_17410);
or U17759 (N_17759,N_17199,N_17205);
nand U17760 (N_17760,N_17442,N_17287);
and U17761 (N_17761,N_17064,N_17233);
nor U17762 (N_17762,N_17203,N_17315);
or U17763 (N_17763,N_17378,N_17334);
nor U17764 (N_17764,N_17207,N_17004);
nand U17765 (N_17765,N_17281,N_17392);
nand U17766 (N_17766,N_17370,N_17350);
nand U17767 (N_17767,N_17414,N_17215);
nor U17768 (N_17768,N_17470,N_17392);
and U17769 (N_17769,N_17334,N_17085);
xnor U17770 (N_17770,N_17017,N_17143);
and U17771 (N_17771,N_17314,N_17217);
nand U17772 (N_17772,N_17013,N_17167);
nor U17773 (N_17773,N_17154,N_17434);
nor U17774 (N_17774,N_17052,N_17214);
and U17775 (N_17775,N_17457,N_17155);
or U17776 (N_17776,N_17063,N_17330);
or U17777 (N_17777,N_17178,N_17128);
nor U17778 (N_17778,N_17276,N_17458);
and U17779 (N_17779,N_17430,N_17354);
nor U17780 (N_17780,N_17171,N_17241);
or U17781 (N_17781,N_17431,N_17465);
and U17782 (N_17782,N_17341,N_17283);
and U17783 (N_17783,N_17226,N_17044);
nor U17784 (N_17784,N_17475,N_17498);
and U17785 (N_17785,N_17206,N_17132);
or U17786 (N_17786,N_17141,N_17458);
nor U17787 (N_17787,N_17134,N_17121);
or U17788 (N_17788,N_17368,N_17183);
nor U17789 (N_17789,N_17456,N_17497);
or U17790 (N_17790,N_17440,N_17456);
nand U17791 (N_17791,N_17186,N_17083);
nand U17792 (N_17792,N_17402,N_17488);
or U17793 (N_17793,N_17461,N_17108);
or U17794 (N_17794,N_17156,N_17428);
nand U17795 (N_17795,N_17409,N_17488);
nand U17796 (N_17796,N_17003,N_17293);
and U17797 (N_17797,N_17261,N_17436);
nand U17798 (N_17798,N_17092,N_17253);
or U17799 (N_17799,N_17188,N_17088);
or U17800 (N_17800,N_17401,N_17139);
xor U17801 (N_17801,N_17393,N_17015);
nor U17802 (N_17802,N_17236,N_17300);
or U17803 (N_17803,N_17279,N_17197);
and U17804 (N_17804,N_17344,N_17109);
and U17805 (N_17805,N_17282,N_17092);
xnor U17806 (N_17806,N_17097,N_17055);
xor U17807 (N_17807,N_17484,N_17152);
or U17808 (N_17808,N_17303,N_17015);
and U17809 (N_17809,N_17242,N_17439);
nor U17810 (N_17810,N_17339,N_17116);
or U17811 (N_17811,N_17459,N_17066);
xor U17812 (N_17812,N_17334,N_17205);
nor U17813 (N_17813,N_17470,N_17067);
or U17814 (N_17814,N_17270,N_17212);
or U17815 (N_17815,N_17103,N_17464);
nor U17816 (N_17816,N_17145,N_17003);
nand U17817 (N_17817,N_17473,N_17115);
nand U17818 (N_17818,N_17358,N_17192);
nand U17819 (N_17819,N_17200,N_17296);
xor U17820 (N_17820,N_17062,N_17193);
nand U17821 (N_17821,N_17240,N_17284);
or U17822 (N_17822,N_17189,N_17288);
or U17823 (N_17823,N_17277,N_17481);
nor U17824 (N_17824,N_17276,N_17208);
and U17825 (N_17825,N_17044,N_17496);
nor U17826 (N_17826,N_17463,N_17222);
and U17827 (N_17827,N_17468,N_17295);
nand U17828 (N_17828,N_17446,N_17262);
nor U17829 (N_17829,N_17296,N_17069);
xnor U17830 (N_17830,N_17298,N_17163);
and U17831 (N_17831,N_17441,N_17490);
nand U17832 (N_17832,N_17204,N_17482);
nand U17833 (N_17833,N_17068,N_17355);
nand U17834 (N_17834,N_17023,N_17332);
or U17835 (N_17835,N_17197,N_17051);
and U17836 (N_17836,N_17426,N_17111);
xnor U17837 (N_17837,N_17167,N_17333);
and U17838 (N_17838,N_17432,N_17182);
and U17839 (N_17839,N_17451,N_17051);
and U17840 (N_17840,N_17118,N_17152);
or U17841 (N_17841,N_17214,N_17173);
nand U17842 (N_17842,N_17008,N_17396);
xnor U17843 (N_17843,N_17045,N_17343);
and U17844 (N_17844,N_17168,N_17497);
nor U17845 (N_17845,N_17214,N_17198);
and U17846 (N_17846,N_17472,N_17265);
nand U17847 (N_17847,N_17152,N_17307);
and U17848 (N_17848,N_17426,N_17040);
nor U17849 (N_17849,N_17346,N_17221);
nand U17850 (N_17850,N_17024,N_17259);
nor U17851 (N_17851,N_17414,N_17379);
xor U17852 (N_17852,N_17125,N_17439);
xnor U17853 (N_17853,N_17059,N_17447);
xor U17854 (N_17854,N_17235,N_17086);
nand U17855 (N_17855,N_17080,N_17044);
or U17856 (N_17856,N_17263,N_17211);
nor U17857 (N_17857,N_17032,N_17149);
or U17858 (N_17858,N_17137,N_17062);
and U17859 (N_17859,N_17444,N_17143);
nor U17860 (N_17860,N_17002,N_17320);
and U17861 (N_17861,N_17151,N_17084);
nor U17862 (N_17862,N_17471,N_17475);
nand U17863 (N_17863,N_17105,N_17141);
xor U17864 (N_17864,N_17455,N_17042);
nand U17865 (N_17865,N_17012,N_17481);
and U17866 (N_17866,N_17066,N_17200);
or U17867 (N_17867,N_17137,N_17296);
or U17868 (N_17868,N_17120,N_17072);
nand U17869 (N_17869,N_17424,N_17133);
and U17870 (N_17870,N_17226,N_17170);
or U17871 (N_17871,N_17006,N_17490);
nand U17872 (N_17872,N_17135,N_17427);
and U17873 (N_17873,N_17013,N_17158);
nor U17874 (N_17874,N_17453,N_17247);
xnor U17875 (N_17875,N_17395,N_17022);
or U17876 (N_17876,N_17369,N_17206);
and U17877 (N_17877,N_17443,N_17447);
nor U17878 (N_17878,N_17481,N_17452);
nand U17879 (N_17879,N_17056,N_17247);
nor U17880 (N_17880,N_17302,N_17066);
and U17881 (N_17881,N_17389,N_17121);
nand U17882 (N_17882,N_17450,N_17102);
nor U17883 (N_17883,N_17385,N_17429);
or U17884 (N_17884,N_17474,N_17241);
nor U17885 (N_17885,N_17013,N_17344);
nand U17886 (N_17886,N_17300,N_17298);
or U17887 (N_17887,N_17326,N_17380);
or U17888 (N_17888,N_17407,N_17293);
xor U17889 (N_17889,N_17093,N_17308);
xor U17890 (N_17890,N_17354,N_17228);
nor U17891 (N_17891,N_17421,N_17168);
and U17892 (N_17892,N_17117,N_17025);
and U17893 (N_17893,N_17208,N_17053);
or U17894 (N_17894,N_17389,N_17186);
or U17895 (N_17895,N_17432,N_17463);
nand U17896 (N_17896,N_17456,N_17403);
and U17897 (N_17897,N_17136,N_17473);
or U17898 (N_17898,N_17187,N_17370);
and U17899 (N_17899,N_17113,N_17490);
nor U17900 (N_17900,N_17446,N_17479);
xor U17901 (N_17901,N_17037,N_17376);
or U17902 (N_17902,N_17312,N_17165);
xnor U17903 (N_17903,N_17172,N_17111);
nor U17904 (N_17904,N_17076,N_17480);
nor U17905 (N_17905,N_17267,N_17329);
or U17906 (N_17906,N_17020,N_17284);
nand U17907 (N_17907,N_17381,N_17290);
xnor U17908 (N_17908,N_17187,N_17047);
nor U17909 (N_17909,N_17469,N_17383);
or U17910 (N_17910,N_17145,N_17354);
and U17911 (N_17911,N_17062,N_17278);
xnor U17912 (N_17912,N_17264,N_17359);
and U17913 (N_17913,N_17138,N_17135);
nor U17914 (N_17914,N_17068,N_17323);
nand U17915 (N_17915,N_17220,N_17427);
nand U17916 (N_17916,N_17306,N_17302);
or U17917 (N_17917,N_17499,N_17221);
nor U17918 (N_17918,N_17023,N_17477);
xor U17919 (N_17919,N_17007,N_17469);
and U17920 (N_17920,N_17374,N_17365);
nor U17921 (N_17921,N_17135,N_17417);
xor U17922 (N_17922,N_17127,N_17178);
nor U17923 (N_17923,N_17070,N_17496);
nand U17924 (N_17924,N_17228,N_17345);
nor U17925 (N_17925,N_17296,N_17156);
xnor U17926 (N_17926,N_17349,N_17111);
and U17927 (N_17927,N_17186,N_17092);
xor U17928 (N_17928,N_17397,N_17220);
nor U17929 (N_17929,N_17194,N_17210);
and U17930 (N_17930,N_17470,N_17011);
nor U17931 (N_17931,N_17108,N_17160);
or U17932 (N_17932,N_17478,N_17370);
xor U17933 (N_17933,N_17405,N_17467);
nor U17934 (N_17934,N_17482,N_17085);
nor U17935 (N_17935,N_17385,N_17162);
nand U17936 (N_17936,N_17467,N_17179);
nor U17937 (N_17937,N_17042,N_17288);
nand U17938 (N_17938,N_17476,N_17009);
nand U17939 (N_17939,N_17365,N_17486);
and U17940 (N_17940,N_17006,N_17179);
and U17941 (N_17941,N_17080,N_17139);
or U17942 (N_17942,N_17254,N_17053);
or U17943 (N_17943,N_17247,N_17096);
nor U17944 (N_17944,N_17106,N_17479);
and U17945 (N_17945,N_17327,N_17136);
nor U17946 (N_17946,N_17372,N_17240);
nand U17947 (N_17947,N_17482,N_17011);
nand U17948 (N_17948,N_17334,N_17249);
and U17949 (N_17949,N_17024,N_17416);
xor U17950 (N_17950,N_17347,N_17307);
xnor U17951 (N_17951,N_17397,N_17365);
xor U17952 (N_17952,N_17358,N_17418);
or U17953 (N_17953,N_17134,N_17448);
nor U17954 (N_17954,N_17421,N_17076);
xor U17955 (N_17955,N_17194,N_17454);
and U17956 (N_17956,N_17349,N_17348);
xor U17957 (N_17957,N_17137,N_17111);
nor U17958 (N_17958,N_17157,N_17498);
and U17959 (N_17959,N_17342,N_17092);
nand U17960 (N_17960,N_17068,N_17368);
and U17961 (N_17961,N_17440,N_17028);
nor U17962 (N_17962,N_17015,N_17069);
or U17963 (N_17963,N_17267,N_17049);
and U17964 (N_17964,N_17290,N_17236);
nand U17965 (N_17965,N_17394,N_17211);
nor U17966 (N_17966,N_17463,N_17368);
nand U17967 (N_17967,N_17136,N_17373);
nand U17968 (N_17968,N_17419,N_17280);
xor U17969 (N_17969,N_17466,N_17175);
nor U17970 (N_17970,N_17021,N_17244);
and U17971 (N_17971,N_17469,N_17218);
or U17972 (N_17972,N_17279,N_17137);
nor U17973 (N_17973,N_17171,N_17317);
nand U17974 (N_17974,N_17016,N_17054);
or U17975 (N_17975,N_17093,N_17442);
xnor U17976 (N_17976,N_17260,N_17012);
xnor U17977 (N_17977,N_17404,N_17138);
nor U17978 (N_17978,N_17029,N_17287);
or U17979 (N_17979,N_17152,N_17046);
xnor U17980 (N_17980,N_17174,N_17276);
or U17981 (N_17981,N_17405,N_17129);
and U17982 (N_17982,N_17076,N_17409);
nor U17983 (N_17983,N_17457,N_17021);
and U17984 (N_17984,N_17022,N_17375);
nand U17985 (N_17985,N_17328,N_17010);
or U17986 (N_17986,N_17355,N_17167);
xnor U17987 (N_17987,N_17048,N_17257);
nor U17988 (N_17988,N_17181,N_17130);
and U17989 (N_17989,N_17409,N_17448);
or U17990 (N_17990,N_17178,N_17025);
and U17991 (N_17991,N_17410,N_17445);
or U17992 (N_17992,N_17292,N_17004);
or U17993 (N_17993,N_17364,N_17424);
nor U17994 (N_17994,N_17084,N_17121);
or U17995 (N_17995,N_17453,N_17030);
nor U17996 (N_17996,N_17208,N_17154);
nor U17997 (N_17997,N_17021,N_17143);
nand U17998 (N_17998,N_17200,N_17417);
and U17999 (N_17999,N_17044,N_17206);
or U18000 (N_18000,N_17724,N_17659);
xor U18001 (N_18001,N_17964,N_17882);
or U18002 (N_18002,N_17908,N_17609);
or U18003 (N_18003,N_17752,N_17878);
and U18004 (N_18004,N_17938,N_17906);
nor U18005 (N_18005,N_17656,N_17683);
nor U18006 (N_18006,N_17931,N_17976);
and U18007 (N_18007,N_17792,N_17751);
xor U18008 (N_18008,N_17860,N_17925);
xor U18009 (N_18009,N_17928,N_17841);
nor U18010 (N_18010,N_17970,N_17584);
xnor U18011 (N_18011,N_17746,N_17922);
nand U18012 (N_18012,N_17807,N_17885);
nand U18013 (N_18013,N_17610,N_17833);
nand U18014 (N_18014,N_17804,N_17978);
xnor U18015 (N_18015,N_17676,N_17822);
nand U18016 (N_18016,N_17814,N_17703);
xor U18017 (N_18017,N_17817,N_17681);
xnor U18018 (N_18018,N_17660,N_17783);
nand U18019 (N_18019,N_17962,N_17859);
nor U18020 (N_18020,N_17919,N_17762);
xor U18021 (N_18021,N_17825,N_17690);
xnor U18022 (N_18022,N_17876,N_17768);
and U18023 (N_18023,N_17716,N_17809);
and U18024 (N_18024,N_17877,N_17571);
xnor U18025 (N_18025,N_17636,N_17590);
nand U18026 (N_18026,N_17553,N_17616);
or U18027 (N_18027,N_17949,N_17510);
nand U18028 (N_18028,N_17969,N_17995);
or U18029 (N_18029,N_17558,N_17577);
and U18030 (N_18030,N_17950,N_17737);
nand U18031 (N_18031,N_17585,N_17945);
or U18032 (N_18032,N_17883,N_17805);
xor U18033 (N_18033,N_17845,N_17834);
and U18034 (N_18034,N_17791,N_17988);
nor U18035 (N_18035,N_17599,N_17898);
xor U18036 (N_18036,N_17530,N_17648);
and U18037 (N_18037,N_17588,N_17521);
nor U18038 (N_18038,N_17608,N_17559);
nand U18039 (N_18039,N_17879,N_17909);
or U18040 (N_18040,N_17920,N_17591);
nand U18041 (N_18041,N_17862,N_17789);
xnor U18042 (N_18042,N_17915,N_17910);
and U18043 (N_18043,N_17874,N_17687);
nand U18044 (N_18044,N_17547,N_17528);
or U18045 (N_18045,N_17890,N_17638);
or U18046 (N_18046,N_17646,N_17677);
and U18047 (N_18047,N_17798,N_17720);
xor U18048 (N_18048,N_17844,N_17843);
or U18049 (N_18049,N_17899,N_17569);
xor U18050 (N_18050,N_17996,N_17633);
xor U18051 (N_18051,N_17535,N_17719);
or U18052 (N_18052,N_17560,N_17722);
or U18053 (N_18053,N_17542,N_17598);
nand U18054 (N_18054,N_17575,N_17544);
xor U18055 (N_18055,N_17963,N_17937);
nand U18056 (N_18056,N_17820,N_17940);
nor U18057 (N_18057,N_17708,N_17960);
or U18058 (N_18058,N_17618,N_17733);
nand U18059 (N_18059,N_17939,N_17796);
nor U18060 (N_18060,N_17505,N_17582);
or U18061 (N_18061,N_17842,N_17948);
nand U18062 (N_18062,N_17873,N_17579);
or U18063 (N_18063,N_17731,N_17508);
or U18064 (N_18064,N_17568,N_17769);
xor U18065 (N_18065,N_17705,N_17797);
nor U18066 (N_18066,N_17852,N_17624);
nand U18067 (N_18067,N_17566,N_17975);
xnor U18068 (N_18068,N_17586,N_17861);
and U18069 (N_18069,N_17527,N_17642);
xor U18070 (N_18070,N_17515,N_17543);
and U18071 (N_18071,N_17835,N_17738);
and U18072 (N_18072,N_17854,N_17956);
xnor U18073 (N_18073,N_17765,N_17857);
nor U18074 (N_18074,N_17570,N_17786);
and U18075 (N_18075,N_17617,N_17800);
xor U18076 (N_18076,N_17525,N_17884);
and U18077 (N_18077,N_17847,N_17594);
or U18078 (N_18078,N_17605,N_17892);
nand U18079 (N_18079,N_17743,N_17750);
or U18080 (N_18080,N_17671,N_17604);
xnor U18081 (N_18081,N_17650,N_17704);
and U18082 (N_18082,N_17702,N_17574);
or U18083 (N_18083,N_17758,N_17697);
and U18084 (N_18084,N_17917,N_17987);
or U18085 (N_18085,N_17572,N_17790);
and U18086 (N_18086,N_17699,N_17897);
xnor U18087 (N_18087,N_17838,N_17710);
xnor U18088 (N_18088,N_17688,N_17649);
nor U18089 (N_18089,N_17596,N_17951);
or U18090 (N_18090,N_17548,N_17924);
or U18091 (N_18091,N_17851,N_17936);
nor U18092 (N_18092,N_17685,N_17562);
nor U18093 (N_18093,N_17721,N_17869);
nand U18094 (N_18094,N_17819,N_17853);
nor U18095 (N_18095,N_17932,N_17644);
xor U18096 (N_18096,N_17620,N_17652);
nor U18097 (N_18097,N_17918,N_17540);
nor U18098 (N_18098,N_17763,N_17546);
or U18099 (N_18099,N_17943,N_17739);
nor U18100 (N_18100,N_17868,N_17840);
nor U18101 (N_18101,N_17895,N_17564);
nand U18102 (N_18102,N_17523,N_17849);
nor U18103 (N_18103,N_17923,N_17679);
nand U18104 (N_18104,N_17985,N_17966);
nand U18105 (N_18105,N_17946,N_17997);
nand U18106 (N_18106,N_17771,N_17713);
nor U18107 (N_18107,N_17753,N_17576);
and U18108 (N_18108,N_17634,N_17669);
and U18109 (N_18109,N_17812,N_17696);
nor U18110 (N_18110,N_17593,N_17513);
xor U18111 (N_18111,N_17999,N_17782);
nor U18112 (N_18112,N_17781,N_17887);
xor U18113 (N_18113,N_17555,N_17955);
xnor U18114 (N_18114,N_17694,N_17886);
nor U18115 (N_18115,N_17779,N_17934);
and U18116 (N_18116,N_17767,N_17846);
and U18117 (N_18117,N_17651,N_17701);
nand U18118 (N_18118,N_17630,N_17600);
nand U18119 (N_18119,N_17803,N_17958);
nand U18120 (N_18120,N_17865,N_17640);
nand U18121 (N_18121,N_17902,N_17994);
nand U18122 (N_18122,N_17654,N_17941);
xnor U18123 (N_18123,N_17592,N_17580);
nor U18124 (N_18124,N_17889,N_17788);
xor U18125 (N_18125,N_17647,N_17631);
nor U18126 (N_18126,N_17602,N_17509);
xnor U18127 (N_18127,N_17992,N_17935);
xnor U18128 (N_18128,N_17666,N_17744);
and U18129 (N_18129,N_17664,N_17520);
and U18130 (N_18130,N_17824,N_17735);
nor U18131 (N_18131,N_17643,N_17611);
nand U18132 (N_18132,N_17871,N_17517);
xor U18133 (N_18133,N_17614,N_17848);
or U18134 (N_18134,N_17668,N_17748);
and U18135 (N_18135,N_17736,N_17828);
nor U18136 (N_18136,N_17619,N_17639);
and U18137 (N_18137,N_17982,N_17684);
nor U18138 (N_18138,N_17531,N_17545);
and U18139 (N_18139,N_17532,N_17691);
and U18140 (N_18140,N_17793,N_17866);
xnor U18141 (N_18141,N_17657,N_17637);
nand U18142 (N_18142,N_17711,N_17506);
xnor U18143 (N_18143,N_17799,N_17658);
nand U18144 (N_18144,N_17565,N_17749);
or U18145 (N_18145,N_17815,N_17726);
nor U18146 (N_18146,N_17759,N_17777);
or U18147 (N_18147,N_17893,N_17888);
xor U18148 (N_18148,N_17770,N_17794);
and U18149 (N_18149,N_17785,N_17551);
nand U18150 (N_18150,N_17529,N_17626);
xnor U18151 (N_18151,N_17811,N_17519);
nor U18152 (N_18152,N_17900,N_17755);
xor U18153 (N_18153,N_17732,N_17977);
nor U18154 (N_18154,N_17766,N_17926);
and U18155 (N_18155,N_17581,N_17730);
nand U18156 (N_18156,N_17891,N_17573);
and U18157 (N_18157,N_17795,N_17747);
or U18158 (N_18158,N_17990,N_17627);
nand U18159 (N_18159,N_17503,N_17801);
or U18160 (N_18160,N_17665,N_17533);
or U18161 (N_18161,N_17896,N_17511);
nand U18162 (N_18162,N_17603,N_17907);
nor U18163 (N_18163,N_17717,N_17622);
and U18164 (N_18164,N_17589,N_17556);
nor U18165 (N_18165,N_17635,N_17816);
xor U18166 (N_18166,N_17692,N_17641);
nand U18167 (N_18167,N_17615,N_17826);
or U18168 (N_18168,N_17818,N_17526);
and U18169 (N_18169,N_17813,N_17968);
or U18170 (N_18170,N_17552,N_17973);
nor U18171 (N_18171,N_17839,N_17921);
and U18172 (N_18172,N_17507,N_17780);
nand U18173 (N_18173,N_17903,N_17727);
xor U18174 (N_18174,N_17645,N_17864);
nand U18175 (N_18175,N_17612,N_17663);
nand U18176 (N_18176,N_17808,N_17723);
and U18177 (N_18177,N_17673,N_17881);
and U18178 (N_18178,N_17561,N_17662);
nand U18179 (N_18179,N_17742,N_17971);
and U18180 (N_18180,N_17991,N_17578);
nor U18181 (N_18181,N_17979,N_17672);
and U18182 (N_18182,N_17695,N_17778);
and U18183 (N_18183,N_17607,N_17855);
nand U18184 (N_18184,N_17764,N_17563);
xnor U18185 (N_18185,N_17952,N_17974);
and U18186 (N_18186,N_17534,N_17707);
nor U18187 (N_18187,N_17856,N_17823);
and U18188 (N_18188,N_17632,N_17725);
or U18189 (N_18189,N_17986,N_17601);
or U18190 (N_18190,N_17830,N_17550);
xor U18191 (N_18191,N_17912,N_17718);
nor U18192 (N_18192,N_17787,N_17712);
nor U18193 (N_18193,N_17698,N_17549);
xor U18194 (N_18194,N_17831,N_17942);
or U18195 (N_18195,N_17829,N_17518);
nand U18196 (N_18196,N_17858,N_17863);
nor U18197 (N_18197,N_17867,N_17901);
xnor U18198 (N_18198,N_17880,N_17983);
xnor U18199 (N_18199,N_17947,N_17514);
or U18200 (N_18200,N_17961,N_17827);
and U18201 (N_18201,N_17972,N_17537);
and U18202 (N_18202,N_17678,N_17980);
nand U18203 (N_18203,N_17595,N_17539);
xnor U18204 (N_18204,N_17745,N_17916);
and U18205 (N_18205,N_17541,N_17729);
xor U18206 (N_18206,N_17557,N_17714);
nor U18207 (N_18207,N_17965,N_17989);
and U18208 (N_18208,N_17554,N_17913);
nand U18209 (N_18209,N_17567,N_17728);
and U18210 (N_18210,N_17944,N_17773);
and U18211 (N_18211,N_17653,N_17760);
and U18212 (N_18212,N_17930,N_17894);
nor U18213 (N_18213,N_17606,N_17625);
nor U18214 (N_18214,N_17741,N_17583);
nor U18215 (N_18215,N_17904,N_17967);
nand U18216 (N_18216,N_17706,N_17802);
nand U18217 (N_18217,N_17772,N_17674);
and U18218 (N_18218,N_17621,N_17905);
or U18219 (N_18219,N_17500,N_17837);
nor U18220 (N_18220,N_17957,N_17998);
and U18221 (N_18221,N_17832,N_17501);
nand U18222 (N_18222,N_17689,N_17512);
nand U18223 (N_18223,N_17538,N_17524);
and U18224 (N_18224,N_17734,N_17613);
and U18225 (N_18225,N_17784,N_17911);
or U18226 (N_18226,N_17686,N_17502);
and U18227 (N_18227,N_17850,N_17821);
and U18228 (N_18228,N_17680,N_17927);
xor U18229 (N_18229,N_17516,N_17715);
nand U18230 (N_18230,N_17682,N_17628);
or U18231 (N_18231,N_17953,N_17693);
xor U18232 (N_18232,N_17954,N_17774);
and U18233 (N_18233,N_17522,N_17655);
xnor U18234 (N_18234,N_17984,N_17675);
and U18235 (N_18235,N_17629,N_17929);
xnor U18236 (N_18236,N_17667,N_17740);
xnor U18237 (N_18237,N_17775,N_17981);
and U18238 (N_18238,N_17709,N_17872);
or U18239 (N_18239,N_17587,N_17661);
nand U18240 (N_18240,N_17623,N_17914);
and U18241 (N_18241,N_17670,N_17536);
or U18242 (N_18242,N_17875,N_17959);
or U18243 (N_18243,N_17933,N_17754);
or U18244 (N_18244,N_17700,N_17993);
nor U18245 (N_18245,N_17757,N_17806);
nand U18246 (N_18246,N_17504,N_17761);
nand U18247 (N_18247,N_17756,N_17776);
and U18248 (N_18248,N_17597,N_17836);
xor U18249 (N_18249,N_17870,N_17810);
nor U18250 (N_18250,N_17977,N_17729);
nand U18251 (N_18251,N_17941,N_17892);
nand U18252 (N_18252,N_17754,N_17909);
nand U18253 (N_18253,N_17506,N_17982);
and U18254 (N_18254,N_17773,N_17982);
or U18255 (N_18255,N_17559,N_17712);
or U18256 (N_18256,N_17613,N_17870);
xnor U18257 (N_18257,N_17974,N_17599);
nand U18258 (N_18258,N_17632,N_17664);
nor U18259 (N_18259,N_17565,N_17668);
nor U18260 (N_18260,N_17888,N_17546);
xor U18261 (N_18261,N_17955,N_17805);
nand U18262 (N_18262,N_17561,N_17813);
or U18263 (N_18263,N_17535,N_17999);
or U18264 (N_18264,N_17968,N_17849);
and U18265 (N_18265,N_17788,N_17792);
and U18266 (N_18266,N_17956,N_17701);
nor U18267 (N_18267,N_17638,N_17576);
nand U18268 (N_18268,N_17566,N_17525);
nand U18269 (N_18269,N_17956,N_17943);
nor U18270 (N_18270,N_17846,N_17647);
xnor U18271 (N_18271,N_17615,N_17607);
and U18272 (N_18272,N_17617,N_17664);
xor U18273 (N_18273,N_17729,N_17587);
nand U18274 (N_18274,N_17737,N_17701);
nand U18275 (N_18275,N_17972,N_17878);
nor U18276 (N_18276,N_17584,N_17731);
nor U18277 (N_18277,N_17899,N_17918);
xnor U18278 (N_18278,N_17928,N_17748);
nor U18279 (N_18279,N_17855,N_17682);
or U18280 (N_18280,N_17997,N_17523);
and U18281 (N_18281,N_17905,N_17969);
or U18282 (N_18282,N_17661,N_17851);
xnor U18283 (N_18283,N_17703,N_17525);
and U18284 (N_18284,N_17792,N_17991);
nor U18285 (N_18285,N_17931,N_17948);
nor U18286 (N_18286,N_17821,N_17869);
or U18287 (N_18287,N_17955,N_17903);
or U18288 (N_18288,N_17922,N_17526);
nor U18289 (N_18289,N_17511,N_17845);
xnor U18290 (N_18290,N_17917,N_17876);
and U18291 (N_18291,N_17845,N_17595);
xor U18292 (N_18292,N_17596,N_17691);
nand U18293 (N_18293,N_17776,N_17767);
and U18294 (N_18294,N_17666,N_17779);
and U18295 (N_18295,N_17988,N_17608);
xnor U18296 (N_18296,N_17547,N_17550);
nand U18297 (N_18297,N_17612,N_17782);
nor U18298 (N_18298,N_17746,N_17957);
and U18299 (N_18299,N_17926,N_17957);
or U18300 (N_18300,N_17987,N_17925);
or U18301 (N_18301,N_17644,N_17984);
nand U18302 (N_18302,N_17600,N_17578);
nand U18303 (N_18303,N_17566,N_17983);
nand U18304 (N_18304,N_17556,N_17795);
xor U18305 (N_18305,N_17725,N_17901);
or U18306 (N_18306,N_17682,N_17690);
nor U18307 (N_18307,N_17631,N_17816);
xnor U18308 (N_18308,N_17655,N_17878);
nand U18309 (N_18309,N_17675,N_17539);
xnor U18310 (N_18310,N_17841,N_17670);
xor U18311 (N_18311,N_17858,N_17992);
nor U18312 (N_18312,N_17509,N_17848);
nand U18313 (N_18313,N_17553,N_17761);
nor U18314 (N_18314,N_17932,N_17659);
or U18315 (N_18315,N_17786,N_17753);
or U18316 (N_18316,N_17711,N_17832);
xnor U18317 (N_18317,N_17781,N_17804);
nor U18318 (N_18318,N_17812,N_17976);
nand U18319 (N_18319,N_17744,N_17891);
and U18320 (N_18320,N_17691,N_17743);
xor U18321 (N_18321,N_17778,N_17866);
and U18322 (N_18322,N_17552,N_17700);
nor U18323 (N_18323,N_17700,N_17626);
and U18324 (N_18324,N_17503,N_17611);
or U18325 (N_18325,N_17861,N_17859);
nand U18326 (N_18326,N_17546,N_17685);
nand U18327 (N_18327,N_17995,N_17773);
or U18328 (N_18328,N_17985,N_17607);
xnor U18329 (N_18329,N_17782,N_17540);
and U18330 (N_18330,N_17596,N_17772);
and U18331 (N_18331,N_17776,N_17517);
and U18332 (N_18332,N_17549,N_17623);
and U18333 (N_18333,N_17914,N_17760);
xor U18334 (N_18334,N_17896,N_17627);
or U18335 (N_18335,N_17791,N_17777);
xor U18336 (N_18336,N_17868,N_17764);
or U18337 (N_18337,N_17676,N_17745);
nand U18338 (N_18338,N_17552,N_17745);
and U18339 (N_18339,N_17564,N_17843);
and U18340 (N_18340,N_17542,N_17685);
nand U18341 (N_18341,N_17516,N_17751);
nand U18342 (N_18342,N_17943,N_17918);
nor U18343 (N_18343,N_17933,N_17889);
nor U18344 (N_18344,N_17871,N_17658);
xnor U18345 (N_18345,N_17553,N_17810);
and U18346 (N_18346,N_17554,N_17955);
nand U18347 (N_18347,N_17778,N_17762);
nor U18348 (N_18348,N_17719,N_17609);
xnor U18349 (N_18349,N_17754,N_17904);
nand U18350 (N_18350,N_17852,N_17612);
nand U18351 (N_18351,N_17896,N_17562);
or U18352 (N_18352,N_17543,N_17838);
or U18353 (N_18353,N_17968,N_17775);
nor U18354 (N_18354,N_17839,N_17655);
xor U18355 (N_18355,N_17626,N_17575);
nor U18356 (N_18356,N_17649,N_17568);
nand U18357 (N_18357,N_17510,N_17708);
or U18358 (N_18358,N_17842,N_17753);
and U18359 (N_18359,N_17874,N_17780);
or U18360 (N_18360,N_17887,N_17974);
and U18361 (N_18361,N_17714,N_17795);
and U18362 (N_18362,N_17552,N_17860);
nand U18363 (N_18363,N_17548,N_17919);
xor U18364 (N_18364,N_17857,N_17936);
nand U18365 (N_18365,N_17993,N_17948);
and U18366 (N_18366,N_17623,N_17963);
xor U18367 (N_18367,N_17612,N_17677);
or U18368 (N_18368,N_17712,N_17662);
xnor U18369 (N_18369,N_17732,N_17588);
nand U18370 (N_18370,N_17742,N_17522);
and U18371 (N_18371,N_17781,N_17634);
nand U18372 (N_18372,N_17568,N_17728);
or U18373 (N_18373,N_17757,N_17876);
xor U18374 (N_18374,N_17888,N_17996);
nand U18375 (N_18375,N_17908,N_17783);
or U18376 (N_18376,N_17706,N_17994);
or U18377 (N_18377,N_17500,N_17737);
nor U18378 (N_18378,N_17916,N_17897);
or U18379 (N_18379,N_17910,N_17962);
and U18380 (N_18380,N_17944,N_17585);
or U18381 (N_18381,N_17608,N_17952);
and U18382 (N_18382,N_17834,N_17509);
and U18383 (N_18383,N_17817,N_17529);
or U18384 (N_18384,N_17533,N_17643);
xor U18385 (N_18385,N_17502,N_17908);
or U18386 (N_18386,N_17918,N_17647);
and U18387 (N_18387,N_17526,N_17645);
nor U18388 (N_18388,N_17968,N_17671);
nor U18389 (N_18389,N_17860,N_17538);
or U18390 (N_18390,N_17848,N_17659);
nand U18391 (N_18391,N_17511,N_17539);
nand U18392 (N_18392,N_17830,N_17785);
xor U18393 (N_18393,N_17896,N_17859);
or U18394 (N_18394,N_17571,N_17761);
and U18395 (N_18395,N_17949,N_17693);
nor U18396 (N_18396,N_17847,N_17560);
xor U18397 (N_18397,N_17629,N_17694);
nor U18398 (N_18398,N_17725,N_17876);
nand U18399 (N_18399,N_17903,N_17718);
nor U18400 (N_18400,N_17671,N_17663);
or U18401 (N_18401,N_17790,N_17734);
and U18402 (N_18402,N_17780,N_17738);
nand U18403 (N_18403,N_17664,N_17727);
nand U18404 (N_18404,N_17670,N_17784);
xnor U18405 (N_18405,N_17803,N_17913);
and U18406 (N_18406,N_17935,N_17552);
and U18407 (N_18407,N_17753,N_17593);
or U18408 (N_18408,N_17983,N_17799);
nand U18409 (N_18409,N_17999,N_17517);
nand U18410 (N_18410,N_17934,N_17900);
nor U18411 (N_18411,N_17584,N_17610);
nand U18412 (N_18412,N_17961,N_17889);
or U18413 (N_18413,N_17609,N_17863);
nand U18414 (N_18414,N_17571,N_17654);
nand U18415 (N_18415,N_17555,N_17541);
or U18416 (N_18416,N_17611,N_17674);
nor U18417 (N_18417,N_17697,N_17667);
xor U18418 (N_18418,N_17589,N_17712);
or U18419 (N_18419,N_17803,N_17521);
nor U18420 (N_18420,N_17574,N_17641);
or U18421 (N_18421,N_17988,N_17625);
xor U18422 (N_18422,N_17809,N_17712);
nand U18423 (N_18423,N_17845,N_17893);
and U18424 (N_18424,N_17919,N_17531);
and U18425 (N_18425,N_17536,N_17968);
and U18426 (N_18426,N_17753,N_17890);
nand U18427 (N_18427,N_17649,N_17588);
nor U18428 (N_18428,N_17602,N_17700);
or U18429 (N_18429,N_17956,N_17914);
nand U18430 (N_18430,N_17569,N_17788);
and U18431 (N_18431,N_17956,N_17591);
and U18432 (N_18432,N_17868,N_17829);
or U18433 (N_18433,N_17915,N_17622);
xor U18434 (N_18434,N_17721,N_17632);
and U18435 (N_18435,N_17925,N_17972);
nor U18436 (N_18436,N_17529,N_17777);
and U18437 (N_18437,N_17868,N_17614);
nor U18438 (N_18438,N_17661,N_17889);
or U18439 (N_18439,N_17769,N_17754);
or U18440 (N_18440,N_17687,N_17860);
or U18441 (N_18441,N_17934,N_17656);
and U18442 (N_18442,N_17848,N_17604);
nor U18443 (N_18443,N_17974,N_17804);
nor U18444 (N_18444,N_17894,N_17622);
and U18445 (N_18445,N_17912,N_17689);
nor U18446 (N_18446,N_17627,N_17941);
xnor U18447 (N_18447,N_17786,N_17544);
nor U18448 (N_18448,N_17584,N_17662);
xor U18449 (N_18449,N_17871,N_17796);
or U18450 (N_18450,N_17525,N_17972);
and U18451 (N_18451,N_17583,N_17710);
xnor U18452 (N_18452,N_17892,N_17594);
nor U18453 (N_18453,N_17687,N_17847);
and U18454 (N_18454,N_17892,N_17580);
nor U18455 (N_18455,N_17676,N_17728);
and U18456 (N_18456,N_17673,N_17683);
and U18457 (N_18457,N_17950,N_17560);
nand U18458 (N_18458,N_17959,N_17892);
or U18459 (N_18459,N_17548,N_17646);
nand U18460 (N_18460,N_17833,N_17690);
or U18461 (N_18461,N_17626,N_17917);
xnor U18462 (N_18462,N_17715,N_17823);
or U18463 (N_18463,N_17803,N_17696);
nor U18464 (N_18464,N_17517,N_17990);
or U18465 (N_18465,N_17823,N_17661);
xor U18466 (N_18466,N_17733,N_17755);
and U18467 (N_18467,N_17526,N_17816);
nor U18468 (N_18468,N_17593,N_17938);
nor U18469 (N_18469,N_17859,N_17881);
nor U18470 (N_18470,N_17654,N_17920);
nand U18471 (N_18471,N_17591,N_17735);
nand U18472 (N_18472,N_17683,N_17609);
and U18473 (N_18473,N_17881,N_17761);
nor U18474 (N_18474,N_17756,N_17768);
and U18475 (N_18475,N_17812,N_17684);
or U18476 (N_18476,N_17539,N_17800);
xor U18477 (N_18477,N_17997,N_17604);
nor U18478 (N_18478,N_17936,N_17777);
or U18479 (N_18479,N_17992,N_17523);
nor U18480 (N_18480,N_17870,N_17680);
nor U18481 (N_18481,N_17605,N_17685);
and U18482 (N_18482,N_17695,N_17511);
and U18483 (N_18483,N_17515,N_17894);
nor U18484 (N_18484,N_17972,N_17962);
nand U18485 (N_18485,N_17652,N_17934);
nand U18486 (N_18486,N_17670,N_17960);
nand U18487 (N_18487,N_17913,N_17963);
xnor U18488 (N_18488,N_17674,N_17950);
or U18489 (N_18489,N_17817,N_17976);
nor U18490 (N_18490,N_17541,N_17655);
xor U18491 (N_18491,N_17828,N_17906);
and U18492 (N_18492,N_17625,N_17677);
nand U18493 (N_18493,N_17768,N_17532);
nor U18494 (N_18494,N_17684,N_17887);
and U18495 (N_18495,N_17731,N_17585);
nand U18496 (N_18496,N_17985,N_17531);
or U18497 (N_18497,N_17993,N_17706);
nor U18498 (N_18498,N_17676,N_17872);
and U18499 (N_18499,N_17735,N_17672);
or U18500 (N_18500,N_18079,N_18210);
nand U18501 (N_18501,N_18015,N_18440);
and U18502 (N_18502,N_18433,N_18185);
and U18503 (N_18503,N_18325,N_18051);
and U18504 (N_18504,N_18023,N_18019);
nor U18505 (N_18505,N_18038,N_18100);
or U18506 (N_18506,N_18491,N_18466);
or U18507 (N_18507,N_18447,N_18139);
nand U18508 (N_18508,N_18104,N_18160);
xor U18509 (N_18509,N_18076,N_18326);
nand U18510 (N_18510,N_18312,N_18146);
xnor U18511 (N_18511,N_18245,N_18263);
nor U18512 (N_18512,N_18112,N_18062);
nor U18513 (N_18513,N_18181,N_18443);
or U18514 (N_18514,N_18078,N_18054);
or U18515 (N_18515,N_18373,N_18480);
xor U18516 (N_18516,N_18095,N_18320);
or U18517 (N_18517,N_18022,N_18234);
xnor U18518 (N_18518,N_18262,N_18059);
nand U18519 (N_18519,N_18353,N_18232);
nand U18520 (N_18520,N_18183,N_18392);
xnor U18521 (N_18521,N_18220,N_18068);
and U18522 (N_18522,N_18401,N_18130);
xnor U18523 (N_18523,N_18282,N_18410);
xnor U18524 (N_18524,N_18006,N_18170);
and U18525 (N_18525,N_18377,N_18499);
or U18526 (N_18526,N_18350,N_18197);
xor U18527 (N_18527,N_18111,N_18148);
nor U18528 (N_18528,N_18364,N_18211);
nor U18529 (N_18529,N_18405,N_18028);
nand U18530 (N_18530,N_18150,N_18376);
or U18531 (N_18531,N_18286,N_18475);
nor U18532 (N_18532,N_18441,N_18287);
or U18533 (N_18533,N_18135,N_18463);
and U18534 (N_18534,N_18495,N_18238);
xnor U18535 (N_18535,N_18385,N_18123);
xor U18536 (N_18536,N_18159,N_18305);
and U18537 (N_18537,N_18196,N_18394);
nand U18538 (N_18538,N_18226,N_18106);
nor U18539 (N_18539,N_18348,N_18246);
or U18540 (N_18540,N_18310,N_18498);
xnor U18541 (N_18541,N_18343,N_18260);
nand U18542 (N_18542,N_18021,N_18296);
or U18543 (N_18543,N_18081,N_18249);
and U18544 (N_18544,N_18467,N_18424);
nand U18545 (N_18545,N_18285,N_18192);
or U18546 (N_18546,N_18259,N_18008);
nand U18547 (N_18547,N_18327,N_18203);
nand U18548 (N_18548,N_18026,N_18336);
nand U18549 (N_18549,N_18479,N_18046);
xor U18550 (N_18550,N_18142,N_18445);
nand U18551 (N_18551,N_18016,N_18360);
nand U18552 (N_18552,N_18031,N_18409);
and U18553 (N_18553,N_18332,N_18161);
or U18554 (N_18554,N_18254,N_18381);
or U18555 (N_18555,N_18184,N_18129);
or U18556 (N_18556,N_18153,N_18319);
and U18557 (N_18557,N_18302,N_18264);
nand U18558 (N_18558,N_18341,N_18363);
nand U18559 (N_18559,N_18241,N_18431);
xor U18560 (N_18560,N_18244,N_18036);
or U18561 (N_18561,N_18370,N_18041);
and U18562 (N_18562,N_18010,N_18261);
nor U18563 (N_18563,N_18290,N_18435);
nand U18564 (N_18564,N_18060,N_18012);
xnor U18565 (N_18565,N_18256,N_18057);
nand U18566 (N_18566,N_18411,N_18291);
xnor U18567 (N_18567,N_18149,N_18223);
or U18568 (N_18568,N_18248,N_18432);
nand U18569 (N_18569,N_18193,N_18400);
and U18570 (N_18570,N_18216,N_18255);
nand U18571 (N_18571,N_18283,N_18235);
xnor U18572 (N_18572,N_18453,N_18288);
and U18573 (N_18573,N_18090,N_18425);
nand U18574 (N_18574,N_18301,N_18404);
nand U18575 (N_18575,N_18276,N_18001);
nand U18576 (N_18576,N_18454,N_18087);
and U18577 (N_18577,N_18213,N_18346);
nor U18578 (N_18578,N_18240,N_18331);
nand U18579 (N_18579,N_18227,N_18329);
or U18580 (N_18580,N_18209,N_18049);
nand U18581 (N_18581,N_18141,N_18271);
or U18582 (N_18582,N_18176,N_18446);
nor U18583 (N_18583,N_18045,N_18250);
xor U18584 (N_18584,N_18243,N_18113);
or U18585 (N_18585,N_18422,N_18402);
nand U18586 (N_18586,N_18020,N_18187);
nor U18587 (N_18587,N_18473,N_18163);
xor U18588 (N_18588,N_18252,N_18205);
or U18589 (N_18589,N_18154,N_18103);
xnor U18590 (N_18590,N_18295,N_18011);
xor U18591 (N_18591,N_18217,N_18098);
xnor U18592 (N_18592,N_18390,N_18372);
and U18593 (N_18593,N_18125,N_18335);
or U18594 (N_18594,N_18471,N_18351);
and U18595 (N_18595,N_18304,N_18084);
nand U18596 (N_18596,N_18279,N_18116);
xnor U18597 (N_18597,N_18448,N_18053);
nor U18598 (N_18598,N_18439,N_18274);
and U18599 (N_18599,N_18228,N_18434);
and U18600 (N_18600,N_18455,N_18119);
xor U18601 (N_18601,N_18427,N_18464);
nand U18602 (N_18602,N_18229,N_18337);
nor U18603 (N_18603,N_18412,N_18052);
xnor U18604 (N_18604,N_18042,N_18316);
nor U18605 (N_18605,N_18131,N_18476);
nand U18606 (N_18606,N_18114,N_18027);
and U18607 (N_18607,N_18069,N_18124);
and U18608 (N_18608,N_18469,N_18225);
nand U18609 (N_18609,N_18147,N_18371);
and U18610 (N_18610,N_18395,N_18330);
or U18611 (N_18611,N_18494,N_18004);
nor U18612 (N_18612,N_18460,N_18474);
and U18613 (N_18613,N_18207,N_18089);
xnor U18614 (N_18614,N_18088,N_18175);
or U18615 (N_18615,N_18354,N_18050);
nand U18616 (N_18616,N_18338,N_18369);
or U18617 (N_18617,N_18292,N_18481);
xnor U18618 (N_18618,N_18270,N_18414);
and U18619 (N_18619,N_18085,N_18470);
and U18620 (N_18620,N_18315,N_18034);
xor U18621 (N_18621,N_18152,N_18167);
and U18622 (N_18622,N_18324,N_18449);
nand U18623 (N_18623,N_18105,N_18172);
or U18624 (N_18624,N_18362,N_18342);
or U18625 (N_18625,N_18014,N_18426);
nor U18626 (N_18626,N_18387,N_18191);
and U18627 (N_18627,N_18061,N_18365);
and U18628 (N_18628,N_18482,N_18265);
xnor U18629 (N_18629,N_18055,N_18236);
nor U18630 (N_18630,N_18430,N_18415);
nand U18631 (N_18631,N_18178,N_18025);
and U18632 (N_18632,N_18033,N_18194);
xor U18633 (N_18633,N_18321,N_18239);
nand U18634 (N_18634,N_18073,N_18115);
nand U18635 (N_18635,N_18155,N_18005);
nand U18636 (N_18636,N_18157,N_18413);
nand U18637 (N_18637,N_18328,N_18251);
xor U18638 (N_18638,N_18117,N_18110);
and U18639 (N_18639,N_18206,N_18037);
or U18640 (N_18640,N_18138,N_18029);
nand U18641 (N_18641,N_18201,N_18436);
xor U18642 (N_18642,N_18386,N_18009);
nand U18643 (N_18643,N_18397,N_18122);
and U18644 (N_18644,N_18035,N_18355);
xor U18645 (N_18645,N_18478,N_18429);
nand U18646 (N_18646,N_18275,N_18349);
nor U18647 (N_18647,N_18407,N_18000);
and U18648 (N_18648,N_18420,N_18379);
xnor U18649 (N_18649,N_18311,N_18177);
or U18650 (N_18650,N_18309,N_18039);
nand U18651 (N_18651,N_18438,N_18303);
nand U18652 (N_18652,N_18233,N_18323);
xnor U18653 (N_18653,N_18136,N_18202);
xnor U18654 (N_18654,N_18166,N_18314);
nand U18655 (N_18655,N_18273,N_18056);
nand U18656 (N_18656,N_18080,N_18374);
or U18657 (N_18657,N_18477,N_18195);
or U18658 (N_18658,N_18182,N_18483);
nor U18659 (N_18659,N_18472,N_18361);
or U18660 (N_18660,N_18272,N_18024);
nor U18661 (N_18661,N_18018,N_18452);
or U18662 (N_18662,N_18002,N_18490);
xor U18663 (N_18663,N_18082,N_18218);
nor U18664 (N_18664,N_18065,N_18189);
nor U18665 (N_18665,N_18007,N_18384);
xnor U18666 (N_18666,N_18318,N_18214);
xor U18667 (N_18667,N_18179,N_18118);
nand U18668 (N_18668,N_18486,N_18137);
and U18669 (N_18669,N_18269,N_18058);
and U18670 (N_18670,N_18066,N_18186);
xor U18671 (N_18671,N_18212,N_18442);
nand U18672 (N_18672,N_18382,N_18418);
xor U18673 (N_18673,N_18074,N_18493);
xor U18674 (N_18674,N_18278,N_18044);
or U18675 (N_18675,N_18307,N_18092);
nand U18676 (N_18676,N_18134,N_18064);
xnor U18677 (N_18677,N_18268,N_18333);
nand U18678 (N_18678,N_18322,N_18257);
or U18679 (N_18679,N_18253,N_18091);
xnor U18680 (N_18680,N_18222,N_18383);
nand U18681 (N_18681,N_18357,N_18067);
nor U18682 (N_18682,N_18168,N_18188);
xor U18683 (N_18683,N_18101,N_18126);
nor U18684 (N_18684,N_18231,N_18461);
and U18685 (N_18685,N_18120,N_18221);
or U18686 (N_18686,N_18204,N_18389);
nand U18687 (N_18687,N_18465,N_18171);
and U18688 (N_18688,N_18102,N_18145);
or U18689 (N_18689,N_18156,N_18094);
or U18690 (N_18690,N_18151,N_18047);
and U18691 (N_18691,N_18497,N_18419);
nand U18692 (N_18692,N_18180,N_18345);
xnor U18693 (N_18693,N_18109,N_18313);
and U18694 (N_18694,N_18366,N_18174);
nand U18695 (N_18695,N_18492,N_18070);
xor U18696 (N_18696,N_18284,N_18219);
xnor U18697 (N_18697,N_18396,N_18132);
nand U18698 (N_18698,N_18317,N_18421);
xor U18699 (N_18699,N_18200,N_18107);
nand U18700 (N_18700,N_18165,N_18398);
nor U18701 (N_18701,N_18017,N_18063);
or U18702 (N_18702,N_18451,N_18444);
or U18703 (N_18703,N_18198,N_18406);
nand U18704 (N_18704,N_18237,N_18300);
xnor U18705 (N_18705,N_18459,N_18352);
nor U18706 (N_18706,N_18380,N_18347);
xor U18707 (N_18707,N_18208,N_18485);
and U18708 (N_18708,N_18340,N_18266);
xnor U18709 (N_18709,N_18128,N_18496);
nor U18710 (N_18710,N_18391,N_18032);
nor U18711 (N_18711,N_18356,N_18294);
xnor U18712 (N_18712,N_18224,N_18158);
nand U18713 (N_18713,N_18281,N_18077);
and U18714 (N_18714,N_18367,N_18199);
and U18715 (N_18715,N_18484,N_18375);
nand U18716 (N_18716,N_18428,N_18456);
xor U18717 (N_18717,N_18099,N_18140);
or U18718 (N_18718,N_18030,N_18267);
or U18719 (N_18719,N_18277,N_18190);
or U18720 (N_18720,N_18230,N_18417);
nor U18721 (N_18721,N_18289,N_18040);
nor U18722 (N_18722,N_18308,N_18487);
or U18723 (N_18723,N_18450,N_18173);
and U18724 (N_18724,N_18457,N_18378);
xnor U18725 (N_18725,N_18403,N_18489);
or U18726 (N_18726,N_18162,N_18097);
nand U18727 (N_18727,N_18393,N_18071);
nor U18728 (N_18728,N_18408,N_18003);
xnor U18729 (N_18729,N_18164,N_18437);
nand U18730 (N_18730,N_18306,N_18242);
xor U18731 (N_18731,N_18344,N_18359);
nor U18732 (N_18732,N_18108,N_18093);
nor U18733 (N_18733,N_18468,N_18121);
nand U18734 (N_18734,N_18127,N_18416);
nor U18735 (N_18735,N_18462,N_18043);
or U18736 (N_18736,N_18358,N_18423);
nand U18737 (N_18737,N_18299,N_18247);
nor U18738 (N_18738,N_18013,N_18083);
or U18739 (N_18739,N_18280,N_18133);
or U18740 (N_18740,N_18293,N_18096);
and U18741 (N_18741,N_18339,N_18086);
and U18742 (N_18742,N_18334,N_18072);
nor U18743 (N_18743,N_18388,N_18075);
and U18744 (N_18744,N_18048,N_18458);
and U18745 (N_18745,N_18399,N_18169);
or U18746 (N_18746,N_18298,N_18143);
xor U18747 (N_18747,N_18488,N_18215);
and U18748 (N_18748,N_18297,N_18258);
xnor U18749 (N_18749,N_18368,N_18144);
or U18750 (N_18750,N_18060,N_18342);
nor U18751 (N_18751,N_18476,N_18109);
or U18752 (N_18752,N_18331,N_18007);
and U18753 (N_18753,N_18473,N_18314);
xnor U18754 (N_18754,N_18073,N_18468);
nand U18755 (N_18755,N_18355,N_18250);
or U18756 (N_18756,N_18378,N_18086);
xor U18757 (N_18757,N_18135,N_18069);
nand U18758 (N_18758,N_18067,N_18075);
xnor U18759 (N_18759,N_18467,N_18346);
nor U18760 (N_18760,N_18180,N_18357);
nand U18761 (N_18761,N_18349,N_18003);
and U18762 (N_18762,N_18379,N_18248);
or U18763 (N_18763,N_18091,N_18028);
nand U18764 (N_18764,N_18031,N_18074);
nor U18765 (N_18765,N_18403,N_18185);
xor U18766 (N_18766,N_18003,N_18485);
xor U18767 (N_18767,N_18314,N_18311);
nand U18768 (N_18768,N_18042,N_18025);
xnor U18769 (N_18769,N_18398,N_18139);
or U18770 (N_18770,N_18331,N_18096);
and U18771 (N_18771,N_18495,N_18222);
xor U18772 (N_18772,N_18291,N_18473);
nor U18773 (N_18773,N_18428,N_18379);
nand U18774 (N_18774,N_18462,N_18350);
xnor U18775 (N_18775,N_18137,N_18414);
xnor U18776 (N_18776,N_18279,N_18475);
or U18777 (N_18777,N_18206,N_18232);
xnor U18778 (N_18778,N_18452,N_18012);
xor U18779 (N_18779,N_18153,N_18170);
xnor U18780 (N_18780,N_18365,N_18439);
and U18781 (N_18781,N_18414,N_18440);
and U18782 (N_18782,N_18212,N_18423);
and U18783 (N_18783,N_18164,N_18111);
or U18784 (N_18784,N_18051,N_18421);
nor U18785 (N_18785,N_18497,N_18319);
xnor U18786 (N_18786,N_18031,N_18452);
xnor U18787 (N_18787,N_18325,N_18341);
nor U18788 (N_18788,N_18467,N_18450);
nand U18789 (N_18789,N_18497,N_18206);
xor U18790 (N_18790,N_18325,N_18402);
nor U18791 (N_18791,N_18453,N_18218);
or U18792 (N_18792,N_18155,N_18113);
nand U18793 (N_18793,N_18393,N_18193);
and U18794 (N_18794,N_18475,N_18166);
nand U18795 (N_18795,N_18392,N_18483);
nor U18796 (N_18796,N_18064,N_18381);
and U18797 (N_18797,N_18204,N_18399);
nand U18798 (N_18798,N_18413,N_18244);
nor U18799 (N_18799,N_18095,N_18237);
xnor U18800 (N_18800,N_18346,N_18124);
nand U18801 (N_18801,N_18273,N_18126);
nand U18802 (N_18802,N_18469,N_18490);
and U18803 (N_18803,N_18212,N_18064);
nor U18804 (N_18804,N_18192,N_18486);
or U18805 (N_18805,N_18498,N_18120);
nand U18806 (N_18806,N_18133,N_18377);
nor U18807 (N_18807,N_18411,N_18395);
or U18808 (N_18808,N_18465,N_18015);
nand U18809 (N_18809,N_18356,N_18447);
nor U18810 (N_18810,N_18450,N_18462);
nor U18811 (N_18811,N_18086,N_18274);
nor U18812 (N_18812,N_18012,N_18371);
or U18813 (N_18813,N_18188,N_18007);
xnor U18814 (N_18814,N_18153,N_18239);
nor U18815 (N_18815,N_18136,N_18266);
nand U18816 (N_18816,N_18227,N_18243);
xnor U18817 (N_18817,N_18451,N_18141);
or U18818 (N_18818,N_18257,N_18157);
or U18819 (N_18819,N_18049,N_18344);
nand U18820 (N_18820,N_18371,N_18468);
xor U18821 (N_18821,N_18401,N_18048);
nor U18822 (N_18822,N_18476,N_18016);
xor U18823 (N_18823,N_18019,N_18307);
nand U18824 (N_18824,N_18378,N_18438);
or U18825 (N_18825,N_18198,N_18074);
and U18826 (N_18826,N_18220,N_18266);
nand U18827 (N_18827,N_18312,N_18276);
xnor U18828 (N_18828,N_18493,N_18274);
nor U18829 (N_18829,N_18094,N_18086);
nand U18830 (N_18830,N_18487,N_18160);
nor U18831 (N_18831,N_18465,N_18467);
and U18832 (N_18832,N_18381,N_18111);
nor U18833 (N_18833,N_18080,N_18088);
xor U18834 (N_18834,N_18236,N_18140);
nand U18835 (N_18835,N_18183,N_18224);
and U18836 (N_18836,N_18189,N_18318);
xnor U18837 (N_18837,N_18475,N_18438);
or U18838 (N_18838,N_18387,N_18309);
and U18839 (N_18839,N_18120,N_18087);
and U18840 (N_18840,N_18334,N_18103);
or U18841 (N_18841,N_18091,N_18295);
or U18842 (N_18842,N_18394,N_18428);
xor U18843 (N_18843,N_18187,N_18308);
xor U18844 (N_18844,N_18253,N_18401);
nor U18845 (N_18845,N_18177,N_18478);
and U18846 (N_18846,N_18391,N_18249);
nand U18847 (N_18847,N_18458,N_18220);
and U18848 (N_18848,N_18061,N_18333);
nand U18849 (N_18849,N_18045,N_18248);
or U18850 (N_18850,N_18025,N_18362);
nor U18851 (N_18851,N_18396,N_18275);
nor U18852 (N_18852,N_18299,N_18329);
nand U18853 (N_18853,N_18471,N_18423);
and U18854 (N_18854,N_18409,N_18394);
and U18855 (N_18855,N_18147,N_18498);
nor U18856 (N_18856,N_18371,N_18137);
nor U18857 (N_18857,N_18379,N_18199);
xor U18858 (N_18858,N_18236,N_18380);
xnor U18859 (N_18859,N_18225,N_18227);
and U18860 (N_18860,N_18344,N_18384);
and U18861 (N_18861,N_18429,N_18449);
nor U18862 (N_18862,N_18234,N_18472);
or U18863 (N_18863,N_18395,N_18109);
nor U18864 (N_18864,N_18405,N_18456);
nor U18865 (N_18865,N_18286,N_18394);
and U18866 (N_18866,N_18316,N_18352);
and U18867 (N_18867,N_18204,N_18037);
nor U18868 (N_18868,N_18159,N_18384);
nand U18869 (N_18869,N_18105,N_18323);
xnor U18870 (N_18870,N_18328,N_18463);
or U18871 (N_18871,N_18013,N_18298);
nand U18872 (N_18872,N_18382,N_18410);
and U18873 (N_18873,N_18013,N_18250);
and U18874 (N_18874,N_18213,N_18326);
xnor U18875 (N_18875,N_18138,N_18484);
nor U18876 (N_18876,N_18170,N_18493);
and U18877 (N_18877,N_18066,N_18411);
xor U18878 (N_18878,N_18029,N_18320);
nand U18879 (N_18879,N_18342,N_18100);
nor U18880 (N_18880,N_18492,N_18463);
and U18881 (N_18881,N_18130,N_18024);
or U18882 (N_18882,N_18151,N_18269);
nor U18883 (N_18883,N_18145,N_18309);
or U18884 (N_18884,N_18351,N_18441);
nand U18885 (N_18885,N_18012,N_18466);
xnor U18886 (N_18886,N_18279,N_18282);
xor U18887 (N_18887,N_18140,N_18182);
xor U18888 (N_18888,N_18265,N_18199);
nand U18889 (N_18889,N_18360,N_18332);
xor U18890 (N_18890,N_18066,N_18275);
xnor U18891 (N_18891,N_18228,N_18481);
and U18892 (N_18892,N_18151,N_18274);
xnor U18893 (N_18893,N_18354,N_18360);
nand U18894 (N_18894,N_18260,N_18252);
nor U18895 (N_18895,N_18251,N_18421);
nand U18896 (N_18896,N_18428,N_18279);
or U18897 (N_18897,N_18253,N_18370);
xnor U18898 (N_18898,N_18144,N_18427);
nand U18899 (N_18899,N_18447,N_18456);
and U18900 (N_18900,N_18412,N_18271);
or U18901 (N_18901,N_18352,N_18119);
nor U18902 (N_18902,N_18452,N_18387);
xor U18903 (N_18903,N_18316,N_18234);
nor U18904 (N_18904,N_18381,N_18083);
xor U18905 (N_18905,N_18034,N_18172);
xor U18906 (N_18906,N_18387,N_18013);
nor U18907 (N_18907,N_18260,N_18338);
xnor U18908 (N_18908,N_18281,N_18487);
and U18909 (N_18909,N_18139,N_18389);
nand U18910 (N_18910,N_18307,N_18299);
nor U18911 (N_18911,N_18077,N_18499);
xor U18912 (N_18912,N_18424,N_18414);
xor U18913 (N_18913,N_18124,N_18157);
nor U18914 (N_18914,N_18286,N_18323);
or U18915 (N_18915,N_18248,N_18326);
nand U18916 (N_18916,N_18264,N_18233);
and U18917 (N_18917,N_18294,N_18107);
nor U18918 (N_18918,N_18166,N_18356);
and U18919 (N_18919,N_18391,N_18453);
and U18920 (N_18920,N_18445,N_18107);
nand U18921 (N_18921,N_18336,N_18283);
and U18922 (N_18922,N_18164,N_18434);
or U18923 (N_18923,N_18225,N_18054);
and U18924 (N_18924,N_18458,N_18114);
xor U18925 (N_18925,N_18176,N_18157);
nand U18926 (N_18926,N_18038,N_18144);
nand U18927 (N_18927,N_18419,N_18052);
or U18928 (N_18928,N_18092,N_18031);
nor U18929 (N_18929,N_18279,N_18093);
nor U18930 (N_18930,N_18011,N_18282);
nand U18931 (N_18931,N_18033,N_18133);
xnor U18932 (N_18932,N_18165,N_18372);
nand U18933 (N_18933,N_18480,N_18032);
or U18934 (N_18934,N_18069,N_18034);
xnor U18935 (N_18935,N_18022,N_18209);
and U18936 (N_18936,N_18428,N_18023);
or U18937 (N_18937,N_18175,N_18481);
or U18938 (N_18938,N_18075,N_18063);
or U18939 (N_18939,N_18068,N_18160);
nor U18940 (N_18940,N_18112,N_18175);
xnor U18941 (N_18941,N_18174,N_18296);
or U18942 (N_18942,N_18235,N_18072);
or U18943 (N_18943,N_18376,N_18045);
nand U18944 (N_18944,N_18388,N_18462);
xor U18945 (N_18945,N_18283,N_18054);
xor U18946 (N_18946,N_18458,N_18172);
or U18947 (N_18947,N_18179,N_18116);
xnor U18948 (N_18948,N_18296,N_18184);
nand U18949 (N_18949,N_18313,N_18183);
and U18950 (N_18950,N_18012,N_18131);
or U18951 (N_18951,N_18354,N_18187);
and U18952 (N_18952,N_18003,N_18370);
and U18953 (N_18953,N_18063,N_18304);
or U18954 (N_18954,N_18189,N_18431);
nor U18955 (N_18955,N_18388,N_18231);
nor U18956 (N_18956,N_18267,N_18119);
and U18957 (N_18957,N_18080,N_18455);
xor U18958 (N_18958,N_18374,N_18303);
nand U18959 (N_18959,N_18136,N_18495);
and U18960 (N_18960,N_18196,N_18315);
and U18961 (N_18961,N_18448,N_18461);
nor U18962 (N_18962,N_18090,N_18082);
and U18963 (N_18963,N_18117,N_18226);
xnor U18964 (N_18964,N_18492,N_18169);
nand U18965 (N_18965,N_18169,N_18441);
xnor U18966 (N_18966,N_18177,N_18426);
and U18967 (N_18967,N_18147,N_18331);
and U18968 (N_18968,N_18187,N_18056);
nand U18969 (N_18969,N_18107,N_18387);
xnor U18970 (N_18970,N_18371,N_18181);
and U18971 (N_18971,N_18003,N_18452);
or U18972 (N_18972,N_18229,N_18321);
and U18973 (N_18973,N_18319,N_18339);
or U18974 (N_18974,N_18308,N_18396);
nand U18975 (N_18975,N_18324,N_18471);
xor U18976 (N_18976,N_18124,N_18117);
and U18977 (N_18977,N_18161,N_18360);
nor U18978 (N_18978,N_18268,N_18229);
and U18979 (N_18979,N_18351,N_18379);
or U18980 (N_18980,N_18042,N_18088);
nor U18981 (N_18981,N_18148,N_18272);
or U18982 (N_18982,N_18112,N_18157);
or U18983 (N_18983,N_18136,N_18184);
and U18984 (N_18984,N_18148,N_18456);
or U18985 (N_18985,N_18338,N_18335);
nor U18986 (N_18986,N_18346,N_18432);
nor U18987 (N_18987,N_18049,N_18259);
and U18988 (N_18988,N_18431,N_18307);
nand U18989 (N_18989,N_18472,N_18387);
xnor U18990 (N_18990,N_18332,N_18152);
nor U18991 (N_18991,N_18479,N_18361);
and U18992 (N_18992,N_18496,N_18413);
nor U18993 (N_18993,N_18003,N_18320);
and U18994 (N_18994,N_18495,N_18418);
nor U18995 (N_18995,N_18077,N_18371);
or U18996 (N_18996,N_18330,N_18405);
nand U18997 (N_18997,N_18136,N_18181);
or U18998 (N_18998,N_18497,N_18205);
and U18999 (N_18999,N_18256,N_18469);
or U19000 (N_19000,N_18545,N_18641);
and U19001 (N_19001,N_18882,N_18554);
or U19002 (N_19002,N_18751,N_18549);
or U19003 (N_19003,N_18804,N_18834);
nand U19004 (N_19004,N_18857,N_18637);
or U19005 (N_19005,N_18952,N_18722);
and U19006 (N_19006,N_18672,N_18847);
xnor U19007 (N_19007,N_18979,N_18916);
nand U19008 (N_19008,N_18967,N_18803);
or U19009 (N_19009,N_18592,N_18521);
and U19010 (N_19010,N_18556,N_18874);
and U19011 (N_19011,N_18801,N_18575);
xor U19012 (N_19012,N_18809,N_18845);
xnor U19013 (N_19013,N_18824,N_18853);
or U19014 (N_19014,N_18741,N_18811);
or U19015 (N_19015,N_18535,N_18547);
or U19016 (N_19016,N_18669,N_18677);
and U19017 (N_19017,N_18897,N_18560);
or U19018 (N_19018,N_18955,N_18534);
or U19019 (N_19019,N_18623,N_18928);
nand U19020 (N_19020,N_18910,N_18912);
or U19021 (N_19021,N_18602,N_18686);
or U19022 (N_19022,N_18702,N_18848);
nand U19023 (N_19023,N_18694,N_18799);
nor U19024 (N_19024,N_18774,N_18517);
and U19025 (N_19025,N_18827,N_18524);
nor U19026 (N_19026,N_18611,N_18917);
or U19027 (N_19027,N_18745,N_18700);
and U19028 (N_19028,N_18533,N_18971);
xnor U19029 (N_19029,N_18783,N_18949);
nand U19030 (N_19030,N_18585,N_18918);
nor U19031 (N_19031,N_18643,N_18706);
xor U19032 (N_19032,N_18940,N_18660);
nor U19033 (N_19033,N_18957,N_18605);
or U19034 (N_19034,N_18557,N_18818);
xnor U19035 (N_19035,N_18586,N_18690);
nand U19036 (N_19036,N_18960,N_18851);
nand U19037 (N_19037,N_18567,N_18542);
and U19038 (N_19038,N_18929,N_18968);
nand U19039 (N_19039,N_18540,N_18919);
nor U19040 (N_19040,N_18973,N_18618);
nand U19041 (N_19041,N_18516,N_18899);
nor U19042 (N_19042,N_18599,N_18890);
xnor U19043 (N_19043,N_18757,N_18877);
and U19044 (N_19044,N_18836,N_18966);
nand U19045 (N_19045,N_18555,N_18691);
xor U19046 (N_19046,N_18584,N_18954);
and U19047 (N_19047,N_18770,N_18806);
nand U19048 (N_19048,N_18697,N_18775);
and U19049 (N_19049,N_18832,N_18797);
and U19050 (N_19050,N_18792,N_18679);
or U19051 (N_19051,N_18839,N_18662);
or U19052 (N_19052,N_18588,N_18872);
xnor U19053 (N_19053,N_18999,N_18552);
xnor U19054 (N_19054,N_18748,N_18959);
and U19055 (N_19055,N_18652,N_18932);
nand U19056 (N_19056,N_18656,N_18707);
xor U19057 (N_19057,N_18768,N_18849);
nor U19058 (N_19058,N_18944,N_18505);
or U19059 (N_19059,N_18536,N_18670);
nor U19060 (N_19060,N_18794,N_18996);
or U19061 (N_19061,N_18657,N_18561);
nor U19062 (N_19062,N_18525,N_18749);
or U19063 (N_19063,N_18914,N_18642);
nand U19064 (N_19064,N_18649,N_18788);
nor U19065 (N_19065,N_18989,N_18862);
nand U19066 (N_19066,N_18764,N_18684);
nand U19067 (N_19067,N_18746,N_18713);
nand U19068 (N_19068,N_18907,N_18509);
or U19069 (N_19069,N_18798,N_18664);
nor U19070 (N_19070,N_18568,N_18587);
or U19071 (N_19071,N_18993,N_18721);
and U19072 (N_19072,N_18913,N_18671);
and U19073 (N_19073,N_18895,N_18511);
and U19074 (N_19074,N_18667,N_18873);
and U19075 (N_19075,N_18889,N_18915);
and U19076 (N_19076,N_18850,N_18841);
or U19077 (N_19077,N_18503,N_18962);
nor U19078 (N_19078,N_18699,N_18590);
and U19079 (N_19079,N_18507,N_18926);
or U19080 (N_19080,N_18769,N_18682);
nor U19081 (N_19081,N_18953,N_18943);
xor U19082 (N_19082,N_18941,N_18674);
xor U19083 (N_19083,N_18761,N_18520);
nand U19084 (N_19084,N_18508,N_18796);
nand U19085 (N_19085,N_18992,N_18638);
or U19086 (N_19086,N_18815,N_18737);
xnor U19087 (N_19087,N_18566,N_18822);
and U19088 (N_19088,N_18879,N_18687);
nand U19089 (N_19089,N_18726,N_18763);
xnor U19090 (N_19090,N_18821,N_18778);
nand U19091 (N_19091,N_18978,N_18734);
xnor U19092 (N_19092,N_18595,N_18529);
xnor U19093 (N_19093,N_18972,N_18601);
nor U19094 (N_19094,N_18622,N_18728);
and U19095 (N_19095,N_18758,N_18784);
or U19096 (N_19096,N_18871,N_18695);
and U19097 (N_19097,N_18830,N_18647);
nor U19098 (N_19098,N_18842,N_18983);
nand U19099 (N_19099,N_18922,N_18578);
and U19100 (N_19100,N_18884,N_18984);
nand U19101 (N_19101,N_18522,N_18998);
nor U19102 (N_19102,N_18580,N_18501);
nor U19103 (N_19103,N_18886,N_18956);
nor U19104 (N_19104,N_18541,N_18630);
xnor U19105 (N_19105,N_18740,N_18854);
nand U19106 (N_19106,N_18885,N_18607);
and U19107 (N_19107,N_18573,N_18701);
or U19108 (N_19108,N_18987,N_18744);
nand U19109 (N_19109,N_18620,N_18712);
and U19110 (N_19110,N_18594,N_18985);
nor U19111 (N_19111,N_18869,N_18866);
xnor U19112 (N_19112,N_18709,N_18698);
nand U19113 (N_19113,N_18574,N_18583);
nor U19114 (N_19114,N_18760,N_18692);
nor U19115 (N_19115,N_18608,N_18891);
nor U19116 (N_19116,N_18844,N_18546);
or U19117 (N_19117,N_18961,N_18831);
or U19118 (N_19118,N_18894,N_18612);
nand U19119 (N_19119,N_18703,N_18793);
xor U19120 (N_19120,N_18924,N_18504);
and U19121 (N_19121,N_18970,N_18500);
and U19122 (N_19122,N_18859,N_18683);
and U19123 (N_19123,N_18523,N_18528);
nor U19124 (N_19124,N_18730,N_18655);
or U19125 (N_19125,N_18909,N_18743);
nor U19126 (N_19126,N_18990,N_18921);
and U19127 (N_19127,N_18765,N_18810);
nor U19128 (N_19128,N_18645,N_18777);
or U19129 (N_19129,N_18597,N_18781);
and U19130 (N_19130,N_18863,N_18668);
nor U19131 (N_19131,N_18988,N_18538);
and U19132 (N_19132,N_18846,N_18865);
xor U19133 (N_19133,N_18976,N_18807);
nor U19134 (N_19134,N_18565,N_18875);
and U19135 (N_19135,N_18878,N_18596);
xnor U19136 (N_19136,N_18950,N_18965);
nand U19137 (N_19137,N_18780,N_18515);
or U19138 (N_19138,N_18795,N_18958);
nand U19139 (N_19139,N_18994,N_18659);
xnor U19140 (N_19140,N_18736,N_18881);
or U19141 (N_19141,N_18654,N_18598);
xor U19142 (N_19142,N_18582,N_18579);
or U19143 (N_19143,N_18685,N_18661);
xor U19144 (N_19144,N_18820,N_18860);
xor U19145 (N_19145,N_18997,N_18593);
nand U19146 (N_19146,N_18902,N_18710);
xor U19147 (N_19147,N_18876,N_18982);
xor U19148 (N_19148,N_18742,N_18510);
or U19149 (N_19149,N_18964,N_18689);
or U19150 (N_19150,N_18813,N_18812);
xnor U19151 (N_19151,N_18880,N_18790);
and U19152 (N_19152,N_18723,N_18614);
xnor U19153 (N_19153,N_18938,N_18711);
xnor U19154 (N_19154,N_18581,N_18738);
nor U19155 (N_19155,N_18939,N_18782);
and U19156 (N_19156,N_18816,N_18603);
or U19157 (N_19157,N_18805,N_18644);
nor U19158 (N_19158,N_18753,N_18635);
and U19159 (N_19159,N_18925,N_18675);
nor U19160 (N_19160,N_18750,N_18840);
nand U19161 (N_19161,N_18786,N_18708);
nand U19162 (N_19162,N_18615,N_18986);
or U19163 (N_19163,N_18591,N_18864);
and U19164 (N_19164,N_18908,N_18977);
xnor U19165 (N_19165,N_18688,N_18530);
nor U19166 (N_19166,N_18969,N_18693);
nand U19167 (N_19167,N_18785,N_18651);
nand U19168 (N_19168,N_18532,N_18564);
xor U19169 (N_19169,N_18559,N_18773);
nand U19170 (N_19170,N_18893,N_18930);
nand U19171 (N_19171,N_18920,N_18828);
nor U19172 (N_19172,N_18762,N_18636);
and U19173 (N_19173,N_18858,N_18755);
and U19174 (N_19174,N_18727,N_18717);
nor U19175 (N_19175,N_18563,N_18613);
or U19176 (N_19176,N_18519,N_18543);
nand U19177 (N_19177,N_18817,N_18735);
or U19178 (N_19178,N_18826,N_18927);
xor U19179 (N_19179,N_18527,N_18896);
and U19180 (N_19180,N_18539,N_18576);
nand U19181 (N_19181,N_18906,N_18678);
or U19182 (N_19182,N_18759,N_18766);
xor U19183 (N_19183,N_18518,N_18629);
or U19184 (N_19184,N_18653,N_18756);
or U19185 (N_19185,N_18855,N_18548);
nor U19186 (N_19186,N_18888,N_18704);
and U19187 (N_19187,N_18901,N_18837);
nor U19188 (N_19188,N_18771,N_18600);
nand U19189 (N_19189,N_18696,N_18808);
nor U19190 (N_19190,N_18627,N_18719);
nand U19191 (N_19191,N_18892,N_18835);
and U19192 (N_19192,N_18610,N_18626);
nor U19193 (N_19193,N_18569,N_18772);
and U19194 (N_19194,N_18625,N_18904);
and U19195 (N_19195,N_18633,N_18658);
nand U19196 (N_19196,N_18621,N_18946);
nor U19197 (N_19197,N_18666,N_18550);
nor U19198 (N_19198,N_18604,N_18665);
nand U19199 (N_19199,N_18663,N_18752);
and U19200 (N_19200,N_18933,N_18923);
or U19201 (N_19201,N_18572,N_18852);
nand U19202 (N_19202,N_18963,N_18787);
xnor U19203 (N_19203,N_18619,N_18729);
and U19204 (N_19204,N_18947,N_18991);
or U19205 (N_19205,N_18948,N_18632);
and U19206 (N_19206,N_18676,N_18825);
nor U19207 (N_19207,N_18754,N_18937);
nand U19208 (N_19208,N_18789,N_18898);
and U19209 (N_19209,N_18980,N_18715);
and U19210 (N_19210,N_18570,N_18732);
nor U19211 (N_19211,N_18616,N_18861);
and U19212 (N_19212,N_18609,N_18823);
nand U19213 (N_19213,N_18526,N_18867);
xor U19214 (N_19214,N_18705,N_18791);
xnor U19215 (N_19215,N_18716,N_18995);
or U19216 (N_19216,N_18931,N_18634);
nor U19217 (N_19217,N_18838,N_18739);
nor U19218 (N_19218,N_18900,N_18631);
and U19219 (N_19219,N_18942,N_18681);
nor U19220 (N_19220,N_18856,N_18577);
nand U19221 (N_19221,N_18936,N_18639);
nor U19222 (N_19222,N_18617,N_18544);
nor U19223 (N_19223,N_18512,N_18829);
nor U19224 (N_19224,N_18537,N_18868);
nand U19225 (N_19225,N_18551,N_18628);
and U19226 (N_19226,N_18747,N_18945);
nand U19227 (N_19227,N_18718,N_18887);
xor U19228 (N_19228,N_18833,N_18975);
and U19229 (N_19229,N_18513,N_18640);
nand U19230 (N_19230,N_18571,N_18903);
or U19231 (N_19231,N_18802,N_18648);
nor U19232 (N_19232,N_18800,N_18814);
and U19233 (N_19233,N_18733,N_18562);
xor U19234 (N_19234,N_18589,N_18673);
nor U19235 (N_19235,N_18724,N_18720);
or U19236 (N_19236,N_18714,N_18506);
nand U19237 (N_19237,N_18981,N_18776);
nand U19238 (N_19238,N_18606,N_18502);
nand U19239 (N_19239,N_18883,N_18870);
nand U19240 (N_19240,N_18819,N_18935);
xnor U19241 (N_19241,N_18731,N_18553);
and U19242 (N_19242,N_18725,N_18624);
and U19243 (N_19243,N_18531,N_18650);
xor U19244 (N_19244,N_18974,N_18680);
nand U19245 (N_19245,N_18767,N_18934);
nor U19246 (N_19246,N_18779,N_18646);
or U19247 (N_19247,N_18911,N_18905);
nor U19248 (N_19248,N_18514,N_18843);
and U19249 (N_19249,N_18951,N_18558);
nor U19250 (N_19250,N_18782,N_18843);
nand U19251 (N_19251,N_18511,N_18719);
and U19252 (N_19252,N_18595,N_18645);
xor U19253 (N_19253,N_18587,N_18807);
and U19254 (N_19254,N_18733,N_18531);
xnor U19255 (N_19255,N_18918,N_18541);
nor U19256 (N_19256,N_18918,N_18980);
nand U19257 (N_19257,N_18829,N_18699);
or U19258 (N_19258,N_18722,N_18736);
and U19259 (N_19259,N_18520,N_18638);
nand U19260 (N_19260,N_18887,N_18921);
or U19261 (N_19261,N_18596,N_18986);
and U19262 (N_19262,N_18755,N_18974);
and U19263 (N_19263,N_18562,N_18511);
nor U19264 (N_19264,N_18913,N_18937);
nand U19265 (N_19265,N_18661,N_18996);
and U19266 (N_19266,N_18554,N_18556);
nor U19267 (N_19267,N_18849,N_18592);
nand U19268 (N_19268,N_18983,N_18958);
xnor U19269 (N_19269,N_18993,N_18621);
or U19270 (N_19270,N_18550,N_18898);
or U19271 (N_19271,N_18886,N_18825);
xor U19272 (N_19272,N_18694,N_18538);
xnor U19273 (N_19273,N_18883,N_18801);
nor U19274 (N_19274,N_18966,N_18853);
nor U19275 (N_19275,N_18508,N_18728);
xnor U19276 (N_19276,N_18999,N_18942);
nand U19277 (N_19277,N_18846,N_18987);
nand U19278 (N_19278,N_18593,N_18543);
nor U19279 (N_19279,N_18888,N_18891);
and U19280 (N_19280,N_18877,N_18684);
nand U19281 (N_19281,N_18553,N_18844);
xnor U19282 (N_19282,N_18880,N_18626);
nor U19283 (N_19283,N_18731,N_18535);
or U19284 (N_19284,N_18708,N_18654);
nand U19285 (N_19285,N_18836,N_18845);
nor U19286 (N_19286,N_18603,N_18778);
nand U19287 (N_19287,N_18940,N_18834);
xor U19288 (N_19288,N_18990,N_18774);
or U19289 (N_19289,N_18944,N_18700);
xnor U19290 (N_19290,N_18643,N_18894);
and U19291 (N_19291,N_18534,N_18708);
nor U19292 (N_19292,N_18548,N_18881);
and U19293 (N_19293,N_18776,N_18931);
nand U19294 (N_19294,N_18524,N_18753);
nand U19295 (N_19295,N_18797,N_18669);
nand U19296 (N_19296,N_18779,N_18911);
nand U19297 (N_19297,N_18985,N_18575);
nor U19298 (N_19298,N_18756,N_18800);
nand U19299 (N_19299,N_18899,N_18765);
xor U19300 (N_19300,N_18766,N_18693);
nor U19301 (N_19301,N_18613,N_18521);
or U19302 (N_19302,N_18683,N_18943);
or U19303 (N_19303,N_18588,N_18812);
xor U19304 (N_19304,N_18517,N_18550);
and U19305 (N_19305,N_18899,N_18563);
or U19306 (N_19306,N_18988,N_18841);
nand U19307 (N_19307,N_18561,N_18685);
nand U19308 (N_19308,N_18881,N_18884);
nor U19309 (N_19309,N_18611,N_18934);
nand U19310 (N_19310,N_18961,N_18882);
nand U19311 (N_19311,N_18548,N_18989);
nand U19312 (N_19312,N_18854,N_18663);
or U19313 (N_19313,N_18532,N_18735);
and U19314 (N_19314,N_18788,N_18528);
and U19315 (N_19315,N_18983,N_18538);
nand U19316 (N_19316,N_18569,N_18662);
nor U19317 (N_19317,N_18932,N_18663);
nor U19318 (N_19318,N_18839,N_18545);
and U19319 (N_19319,N_18881,N_18739);
xor U19320 (N_19320,N_18748,N_18501);
xnor U19321 (N_19321,N_18993,N_18985);
or U19322 (N_19322,N_18787,N_18659);
or U19323 (N_19323,N_18876,N_18804);
nor U19324 (N_19324,N_18955,N_18926);
and U19325 (N_19325,N_18974,N_18558);
nand U19326 (N_19326,N_18575,N_18562);
nand U19327 (N_19327,N_18546,N_18735);
or U19328 (N_19328,N_18956,N_18776);
nor U19329 (N_19329,N_18878,N_18724);
nor U19330 (N_19330,N_18737,N_18709);
and U19331 (N_19331,N_18630,N_18699);
or U19332 (N_19332,N_18600,N_18881);
and U19333 (N_19333,N_18979,N_18694);
and U19334 (N_19334,N_18842,N_18703);
and U19335 (N_19335,N_18840,N_18549);
xor U19336 (N_19336,N_18844,N_18849);
xor U19337 (N_19337,N_18504,N_18575);
or U19338 (N_19338,N_18608,N_18744);
xor U19339 (N_19339,N_18839,N_18524);
xor U19340 (N_19340,N_18906,N_18820);
and U19341 (N_19341,N_18954,N_18769);
nor U19342 (N_19342,N_18646,N_18612);
nand U19343 (N_19343,N_18976,N_18665);
and U19344 (N_19344,N_18560,N_18788);
nor U19345 (N_19345,N_18536,N_18574);
and U19346 (N_19346,N_18977,N_18784);
xnor U19347 (N_19347,N_18508,N_18871);
xor U19348 (N_19348,N_18966,N_18969);
xor U19349 (N_19349,N_18551,N_18797);
nand U19350 (N_19350,N_18876,N_18932);
nor U19351 (N_19351,N_18896,N_18833);
or U19352 (N_19352,N_18851,N_18732);
xor U19353 (N_19353,N_18885,N_18786);
xnor U19354 (N_19354,N_18603,N_18782);
nand U19355 (N_19355,N_18532,N_18699);
xnor U19356 (N_19356,N_18803,N_18601);
xnor U19357 (N_19357,N_18987,N_18623);
xor U19358 (N_19358,N_18679,N_18799);
nor U19359 (N_19359,N_18533,N_18603);
nand U19360 (N_19360,N_18879,N_18848);
nor U19361 (N_19361,N_18682,N_18683);
nor U19362 (N_19362,N_18578,N_18630);
and U19363 (N_19363,N_18820,N_18951);
nor U19364 (N_19364,N_18644,N_18630);
or U19365 (N_19365,N_18524,N_18793);
or U19366 (N_19366,N_18580,N_18812);
xnor U19367 (N_19367,N_18805,N_18963);
nor U19368 (N_19368,N_18757,N_18604);
xnor U19369 (N_19369,N_18531,N_18598);
nor U19370 (N_19370,N_18539,N_18980);
nor U19371 (N_19371,N_18803,N_18928);
nor U19372 (N_19372,N_18869,N_18824);
xor U19373 (N_19373,N_18547,N_18803);
and U19374 (N_19374,N_18727,N_18750);
or U19375 (N_19375,N_18856,N_18848);
and U19376 (N_19376,N_18699,N_18828);
xor U19377 (N_19377,N_18957,N_18604);
and U19378 (N_19378,N_18774,N_18761);
nor U19379 (N_19379,N_18981,N_18738);
xor U19380 (N_19380,N_18524,N_18697);
and U19381 (N_19381,N_18650,N_18523);
nand U19382 (N_19382,N_18580,N_18852);
or U19383 (N_19383,N_18839,N_18624);
xnor U19384 (N_19384,N_18664,N_18596);
xnor U19385 (N_19385,N_18631,N_18592);
and U19386 (N_19386,N_18522,N_18639);
nand U19387 (N_19387,N_18955,N_18623);
nand U19388 (N_19388,N_18500,N_18791);
or U19389 (N_19389,N_18909,N_18739);
xor U19390 (N_19390,N_18562,N_18551);
xor U19391 (N_19391,N_18775,N_18723);
nand U19392 (N_19392,N_18584,N_18640);
xnor U19393 (N_19393,N_18914,N_18548);
or U19394 (N_19394,N_18686,N_18703);
nand U19395 (N_19395,N_18547,N_18733);
nor U19396 (N_19396,N_18784,N_18645);
and U19397 (N_19397,N_18587,N_18939);
or U19398 (N_19398,N_18649,N_18733);
nand U19399 (N_19399,N_18835,N_18732);
nand U19400 (N_19400,N_18914,N_18669);
nand U19401 (N_19401,N_18821,N_18898);
or U19402 (N_19402,N_18864,N_18957);
and U19403 (N_19403,N_18601,N_18840);
or U19404 (N_19404,N_18602,N_18825);
nand U19405 (N_19405,N_18604,N_18924);
nor U19406 (N_19406,N_18819,N_18712);
nand U19407 (N_19407,N_18754,N_18583);
nand U19408 (N_19408,N_18778,N_18676);
xnor U19409 (N_19409,N_18982,N_18996);
xor U19410 (N_19410,N_18796,N_18550);
xor U19411 (N_19411,N_18717,N_18526);
or U19412 (N_19412,N_18531,N_18564);
and U19413 (N_19413,N_18741,N_18736);
nor U19414 (N_19414,N_18828,N_18566);
xnor U19415 (N_19415,N_18984,N_18946);
xnor U19416 (N_19416,N_18839,N_18615);
or U19417 (N_19417,N_18956,N_18546);
xor U19418 (N_19418,N_18896,N_18717);
and U19419 (N_19419,N_18872,N_18947);
xor U19420 (N_19420,N_18688,N_18531);
or U19421 (N_19421,N_18555,N_18871);
nand U19422 (N_19422,N_18736,N_18646);
nand U19423 (N_19423,N_18633,N_18920);
or U19424 (N_19424,N_18873,N_18696);
nand U19425 (N_19425,N_18615,N_18869);
xor U19426 (N_19426,N_18824,N_18874);
xor U19427 (N_19427,N_18819,N_18585);
and U19428 (N_19428,N_18777,N_18686);
and U19429 (N_19429,N_18504,N_18741);
nor U19430 (N_19430,N_18826,N_18514);
nor U19431 (N_19431,N_18737,N_18740);
xor U19432 (N_19432,N_18923,N_18830);
nor U19433 (N_19433,N_18533,N_18752);
and U19434 (N_19434,N_18847,N_18667);
nand U19435 (N_19435,N_18961,N_18967);
nand U19436 (N_19436,N_18554,N_18838);
nor U19437 (N_19437,N_18694,N_18928);
nand U19438 (N_19438,N_18717,N_18505);
xor U19439 (N_19439,N_18919,N_18649);
nor U19440 (N_19440,N_18604,N_18647);
nor U19441 (N_19441,N_18598,N_18926);
xnor U19442 (N_19442,N_18647,N_18817);
and U19443 (N_19443,N_18921,N_18658);
and U19444 (N_19444,N_18581,N_18930);
xnor U19445 (N_19445,N_18688,N_18776);
xnor U19446 (N_19446,N_18694,N_18511);
nor U19447 (N_19447,N_18744,N_18566);
or U19448 (N_19448,N_18637,N_18815);
xor U19449 (N_19449,N_18724,N_18980);
nand U19450 (N_19450,N_18579,N_18922);
or U19451 (N_19451,N_18983,N_18708);
and U19452 (N_19452,N_18841,N_18600);
or U19453 (N_19453,N_18725,N_18770);
nor U19454 (N_19454,N_18984,N_18673);
xnor U19455 (N_19455,N_18957,N_18584);
or U19456 (N_19456,N_18555,N_18617);
or U19457 (N_19457,N_18610,N_18655);
xnor U19458 (N_19458,N_18723,N_18774);
xnor U19459 (N_19459,N_18919,N_18911);
and U19460 (N_19460,N_18769,N_18551);
or U19461 (N_19461,N_18724,N_18565);
and U19462 (N_19462,N_18712,N_18840);
nor U19463 (N_19463,N_18712,N_18785);
nor U19464 (N_19464,N_18938,N_18887);
nand U19465 (N_19465,N_18503,N_18922);
nand U19466 (N_19466,N_18903,N_18909);
or U19467 (N_19467,N_18676,N_18708);
nor U19468 (N_19468,N_18853,N_18836);
xnor U19469 (N_19469,N_18523,N_18853);
nand U19470 (N_19470,N_18989,N_18917);
nor U19471 (N_19471,N_18870,N_18578);
nand U19472 (N_19472,N_18763,N_18505);
xnor U19473 (N_19473,N_18791,N_18922);
nand U19474 (N_19474,N_18550,N_18805);
xnor U19475 (N_19475,N_18590,N_18802);
nor U19476 (N_19476,N_18728,N_18715);
nand U19477 (N_19477,N_18534,N_18876);
nor U19478 (N_19478,N_18656,N_18556);
nand U19479 (N_19479,N_18595,N_18906);
xor U19480 (N_19480,N_18738,N_18790);
and U19481 (N_19481,N_18796,N_18578);
and U19482 (N_19482,N_18886,N_18954);
xnor U19483 (N_19483,N_18955,N_18767);
xor U19484 (N_19484,N_18627,N_18510);
nor U19485 (N_19485,N_18900,N_18568);
nand U19486 (N_19486,N_18876,N_18694);
and U19487 (N_19487,N_18883,N_18697);
xor U19488 (N_19488,N_18730,N_18684);
nand U19489 (N_19489,N_18733,N_18688);
nand U19490 (N_19490,N_18769,N_18612);
and U19491 (N_19491,N_18783,N_18581);
and U19492 (N_19492,N_18748,N_18584);
nand U19493 (N_19493,N_18539,N_18558);
nand U19494 (N_19494,N_18580,N_18845);
nand U19495 (N_19495,N_18578,N_18845);
nand U19496 (N_19496,N_18661,N_18553);
and U19497 (N_19497,N_18812,N_18691);
nor U19498 (N_19498,N_18856,N_18831);
xor U19499 (N_19499,N_18791,N_18646);
or U19500 (N_19500,N_19071,N_19349);
nor U19501 (N_19501,N_19313,N_19241);
or U19502 (N_19502,N_19486,N_19019);
and U19503 (N_19503,N_19386,N_19412);
and U19504 (N_19504,N_19244,N_19148);
nor U19505 (N_19505,N_19156,N_19339);
nor U19506 (N_19506,N_19322,N_19024);
or U19507 (N_19507,N_19065,N_19480);
and U19508 (N_19508,N_19410,N_19005);
xor U19509 (N_19509,N_19438,N_19272);
nor U19510 (N_19510,N_19429,N_19120);
nand U19511 (N_19511,N_19017,N_19149);
and U19512 (N_19512,N_19343,N_19111);
and U19513 (N_19513,N_19014,N_19176);
nor U19514 (N_19514,N_19205,N_19228);
xnor U19515 (N_19515,N_19471,N_19278);
and U19516 (N_19516,N_19021,N_19018);
nand U19517 (N_19517,N_19179,N_19215);
or U19518 (N_19518,N_19309,N_19100);
nor U19519 (N_19519,N_19105,N_19253);
or U19520 (N_19520,N_19183,N_19122);
nand U19521 (N_19521,N_19242,N_19012);
and U19522 (N_19522,N_19470,N_19328);
nand U19523 (N_19523,N_19033,N_19494);
nand U19524 (N_19524,N_19209,N_19321);
xor U19525 (N_19525,N_19364,N_19069);
xnor U19526 (N_19526,N_19393,N_19155);
nand U19527 (N_19527,N_19492,N_19308);
xnor U19528 (N_19528,N_19340,N_19239);
or U19529 (N_19529,N_19185,N_19295);
or U19530 (N_19530,N_19161,N_19384);
xnor U19531 (N_19531,N_19327,N_19367);
xnor U19532 (N_19532,N_19263,N_19459);
or U19533 (N_19533,N_19041,N_19271);
xor U19534 (N_19534,N_19398,N_19196);
xnor U19535 (N_19535,N_19468,N_19143);
nor U19536 (N_19536,N_19441,N_19455);
xnor U19537 (N_19537,N_19422,N_19286);
nor U19538 (N_19538,N_19277,N_19079);
and U19539 (N_19539,N_19366,N_19414);
or U19540 (N_19540,N_19056,N_19224);
xor U19541 (N_19541,N_19285,N_19227);
and U19542 (N_19542,N_19266,N_19391);
and U19543 (N_19543,N_19003,N_19302);
or U19544 (N_19544,N_19347,N_19469);
and U19545 (N_19545,N_19324,N_19119);
nand U19546 (N_19546,N_19448,N_19297);
nor U19547 (N_19547,N_19249,N_19274);
nor U19548 (N_19548,N_19118,N_19163);
or U19549 (N_19549,N_19446,N_19430);
nor U19550 (N_19550,N_19232,N_19081);
nand U19551 (N_19551,N_19117,N_19047);
or U19552 (N_19552,N_19315,N_19086);
nand U19553 (N_19553,N_19166,N_19445);
nor U19554 (N_19554,N_19058,N_19043);
nand U19555 (N_19555,N_19326,N_19057);
and U19556 (N_19556,N_19496,N_19000);
nand U19557 (N_19557,N_19475,N_19458);
nand U19558 (N_19558,N_19075,N_19354);
nor U19559 (N_19559,N_19035,N_19174);
xor U19560 (N_19560,N_19167,N_19137);
and U19561 (N_19561,N_19273,N_19235);
xor U19562 (N_19562,N_19423,N_19045);
and U19563 (N_19563,N_19067,N_19481);
nor U19564 (N_19564,N_19433,N_19332);
and U19565 (N_19565,N_19020,N_19076);
nand U19566 (N_19566,N_19390,N_19477);
xor U19567 (N_19567,N_19136,N_19029);
nor U19568 (N_19568,N_19304,N_19134);
nand U19569 (N_19569,N_19281,N_19098);
or U19570 (N_19570,N_19084,N_19046);
nor U19571 (N_19571,N_19157,N_19094);
or U19572 (N_19572,N_19038,N_19173);
nor U19573 (N_19573,N_19193,N_19026);
nand U19574 (N_19574,N_19030,N_19202);
nor U19575 (N_19575,N_19211,N_19415);
and U19576 (N_19576,N_19113,N_19397);
nor U19577 (N_19577,N_19307,N_19303);
or U19578 (N_19578,N_19437,N_19133);
or U19579 (N_19579,N_19497,N_19432);
nand U19580 (N_19580,N_19221,N_19087);
xor U19581 (N_19581,N_19452,N_19363);
or U19582 (N_19582,N_19400,N_19218);
nor U19583 (N_19583,N_19061,N_19187);
and U19584 (N_19584,N_19022,N_19395);
or U19585 (N_19585,N_19417,N_19311);
nand U19586 (N_19586,N_19060,N_19370);
nand U19587 (N_19587,N_19270,N_19381);
xnor U19588 (N_19588,N_19039,N_19219);
nor U19589 (N_19589,N_19288,N_19158);
nor U19590 (N_19590,N_19256,N_19368);
nand U19591 (N_19591,N_19210,N_19344);
or U19592 (N_19592,N_19376,N_19457);
and U19593 (N_19593,N_19225,N_19460);
nor U19594 (N_19594,N_19265,N_19341);
nor U19595 (N_19595,N_19170,N_19216);
xnor U19596 (N_19596,N_19154,N_19204);
xnor U19597 (N_19597,N_19255,N_19192);
xnor U19598 (N_19598,N_19290,N_19195);
nand U19599 (N_19599,N_19233,N_19015);
and U19600 (N_19600,N_19335,N_19392);
nor U19601 (N_19601,N_19032,N_19482);
or U19602 (N_19602,N_19372,N_19345);
xnor U19603 (N_19603,N_19403,N_19093);
and U19604 (N_19604,N_19431,N_19177);
and U19605 (N_19605,N_19007,N_19331);
and U19606 (N_19606,N_19254,N_19101);
and U19607 (N_19607,N_19449,N_19418);
nand U19608 (N_19608,N_19305,N_19329);
nand U19609 (N_19609,N_19048,N_19357);
or U19610 (N_19610,N_19108,N_19325);
and U19611 (N_19611,N_19268,N_19292);
and U19612 (N_19612,N_19055,N_19405);
and U19613 (N_19613,N_19251,N_19109);
nand U19614 (N_19614,N_19217,N_19451);
and U19615 (N_19615,N_19011,N_19054);
nor U19616 (N_19616,N_19352,N_19427);
xnor U19617 (N_19617,N_19258,N_19301);
or U19618 (N_19618,N_19495,N_19413);
nor U19619 (N_19619,N_19247,N_19106);
and U19620 (N_19620,N_19197,N_19236);
nand U19621 (N_19621,N_19178,N_19318);
xor U19622 (N_19622,N_19073,N_19359);
or U19623 (N_19623,N_19276,N_19159);
and U19624 (N_19624,N_19490,N_19262);
nor U19625 (N_19625,N_19131,N_19443);
and U19626 (N_19626,N_19394,N_19099);
xor U19627 (N_19627,N_19208,N_19411);
nand U19628 (N_19628,N_19483,N_19013);
or U19629 (N_19629,N_19385,N_19153);
nand U19630 (N_19630,N_19124,N_19097);
or U19631 (N_19631,N_19456,N_19378);
and U19632 (N_19632,N_19184,N_19186);
nor U19633 (N_19633,N_19072,N_19404);
and U19634 (N_19634,N_19004,N_19330);
and U19635 (N_19635,N_19213,N_19360);
nor U19636 (N_19636,N_19252,N_19289);
nand U19637 (N_19637,N_19487,N_19191);
and U19638 (N_19638,N_19280,N_19316);
and U19639 (N_19639,N_19127,N_19466);
xnor U19640 (N_19640,N_19478,N_19181);
nor U19641 (N_19641,N_19066,N_19006);
xor U19642 (N_19642,N_19267,N_19356);
or U19643 (N_19643,N_19031,N_19162);
nor U19644 (N_19644,N_19010,N_19375);
or U19645 (N_19645,N_19420,N_19214);
xnor U19646 (N_19646,N_19092,N_19474);
nand U19647 (N_19647,N_19287,N_19358);
or U19648 (N_19648,N_19189,N_19082);
nand U19649 (N_19649,N_19201,N_19409);
xor U19650 (N_19650,N_19231,N_19182);
or U19651 (N_19651,N_19426,N_19044);
xnor U19652 (N_19652,N_19485,N_19180);
or U19653 (N_19653,N_19028,N_19001);
xnor U19654 (N_19654,N_19257,N_19128);
nand U19655 (N_19655,N_19283,N_19190);
nor U19656 (N_19656,N_19051,N_19172);
or U19657 (N_19657,N_19425,N_19245);
or U19658 (N_19658,N_19034,N_19361);
and U19659 (N_19659,N_19453,N_19164);
nor U19660 (N_19660,N_19115,N_19104);
or U19661 (N_19661,N_19300,N_19317);
and U19662 (N_19662,N_19207,N_19473);
nand U19663 (N_19663,N_19291,N_19036);
xnor U19664 (N_19664,N_19234,N_19140);
nand U19665 (N_19665,N_19123,N_19248);
xor U19666 (N_19666,N_19279,N_19169);
nor U19667 (N_19667,N_19016,N_19171);
nand U19668 (N_19668,N_19447,N_19450);
nand U19669 (N_19669,N_19319,N_19440);
xnor U19670 (N_19670,N_19399,N_19095);
xor U19671 (N_19671,N_19064,N_19229);
or U19672 (N_19672,N_19063,N_19369);
xor U19673 (N_19673,N_19348,N_19489);
or U19674 (N_19674,N_19261,N_19306);
or U19675 (N_19675,N_19362,N_19238);
nand U19676 (N_19676,N_19121,N_19138);
xor U19677 (N_19677,N_19243,N_19275);
nor U19678 (N_19678,N_19371,N_19091);
nand U19679 (N_19679,N_19088,N_19042);
and U19680 (N_19680,N_19436,N_19342);
and U19681 (N_19681,N_19387,N_19152);
or U19682 (N_19682,N_19365,N_19346);
and U19683 (N_19683,N_19090,N_19223);
nand U19684 (N_19684,N_19078,N_19002);
nand U19685 (N_19685,N_19023,N_19025);
nand U19686 (N_19686,N_19135,N_19498);
nor U19687 (N_19687,N_19168,N_19132);
or U19688 (N_19688,N_19114,N_19424);
nor U19689 (N_19689,N_19040,N_19070);
and U19690 (N_19690,N_19008,N_19416);
nand U19691 (N_19691,N_19464,N_19350);
xor U19692 (N_19692,N_19454,N_19050);
xnor U19693 (N_19693,N_19080,N_19293);
xnor U19694 (N_19694,N_19334,N_19160);
and U19695 (N_19695,N_19260,N_19126);
xnor U19696 (N_19696,N_19408,N_19479);
or U19697 (N_19697,N_19298,N_19200);
and U19698 (N_19698,N_19491,N_19089);
and U19699 (N_19699,N_19151,N_19439);
and U19700 (N_19700,N_19062,N_19096);
and U19701 (N_19701,N_19467,N_19336);
nor U19702 (N_19702,N_19077,N_19246);
or U19703 (N_19703,N_19373,N_19310);
or U19704 (N_19704,N_19240,N_19389);
nor U19705 (N_19705,N_19442,N_19220);
nand U19706 (N_19706,N_19383,N_19259);
or U19707 (N_19707,N_19147,N_19052);
nor U19708 (N_19708,N_19027,N_19068);
and U19709 (N_19709,N_19338,N_19264);
nand U19710 (N_19710,N_19407,N_19421);
and U19711 (N_19711,N_19396,N_19484);
xor U19712 (N_19712,N_19203,N_19388);
xor U19713 (N_19713,N_19434,N_19296);
nor U19714 (N_19714,N_19382,N_19125);
or U19715 (N_19715,N_19226,N_19444);
and U19716 (N_19716,N_19112,N_19009);
xor U19717 (N_19717,N_19165,N_19435);
or U19718 (N_19718,N_19107,N_19102);
xor U19719 (N_19719,N_19103,N_19461);
nand U19720 (N_19720,N_19406,N_19472);
nand U19721 (N_19721,N_19146,N_19206);
nand U19722 (N_19722,N_19351,N_19476);
nand U19723 (N_19723,N_19199,N_19337);
xor U19724 (N_19724,N_19222,N_19499);
xor U19725 (N_19725,N_19463,N_19355);
nand U19726 (N_19726,N_19150,N_19379);
or U19727 (N_19727,N_19059,N_19074);
or U19728 (N_19728,N_19145,N_19462);
and U19729 (N_19729,N_19049,N_19333);
xnor U19730 (N_19730,N_19083,N_19250);
or U19731 (N_19731,N_19142,N_19037);
and U19732 (N_19732,N_19294,N_19188);
xor U19733 (N_19733,N_19320,N_19194);
nand U19734 (N_19734,N_19116,N_19465);
nand U19735 (N_19735,N_19237,N_19299);
xor U19736 (N_19736,N_19284,N_19269);
and U19737 (N_19737,N_19428,N_19401);
nand U19738 (N_19738,N_19130,N_19144);
nand U19739 (N_19739,N_19493,N_19419);
nand U19740 (N_19740,N_19380,N_19110);
or U19741 (N_19741,N_19053,N_19230);
or U19742 (N_19742,N_19402,N_19175);
or U19743 (N_19743,N_19488,N_19085);
or U19744 (N_19744,N_19312,N_19323);
xor U19745 (N_19745,N_19198,N_19314);
or U19746 (N_19746,N_19282,N_19374);
xor U19747 (N_19747,N_19129,N_19141);
nor U19748 (N_19748,N_19353,N_19377);
or U19749 (N_19749,N_19139,N_19212);
and U19750 (N_19750,N_19362,N_19218);
xor U19751 (N_19751,N_19356,N_19086);
xor U19752 (N_19752,N_19453,N_19037);
xor U19753 (N_19753,N_19390,N_19039);
nand U19754 (N_19754,N_19425,N_19262);
nor U19755 (N_19755,N_19459,N_19457);
and U19756 (N_19756,N_19337,N_19280);
or U19757 (N_19757,N_19426,N_19223);
or U19758 (N_19758,N_19478,N_19145);
xnor U19759 (N_19759,N_19418,N_19395);
nor U19760 (N_19760,N_19152,N_19136);
or U19761 (N_19761,N_19302,N_19276);
and U19762 (N_19762,N_19145,N_19287);
and U19763 (N_19763,N_19230,N_19112);
xnor U19764 (N_19764,N_19151,N_19043);
xnor U19765 (N_19765,N_19094,N_19421);
nor U19766 (N_19766,N_19491,N_19224);
xor U19767 (N_19767,N_19375,N_19141);
nand U19768 (N_19768,N_19120,N_19437);
nand U19769 (N_19769,N_19170,N_19389);
xor U19770 (N_19770,N_19191,N_19360);
or U19771 (N_19771,N_19046,N_19182);
and U19772 (N_19772,N_19306,N_19001);
and U19773 (N_19773,N_19401,N_19132);
nor U19774 (N_19774,N_19330,N_19318);
or U19775 (N_19775,N_19122,N_19311);
xor U19776 (N_19776,N_19001,N_19250);
or U19777 (N_19777,N_19074,N_19465);
nor U19778 (N_19778,N_19075,N_19439);
and U19779 (N_19779,N_19330,N_19380);
nor U19780 (N_19780,N_19400,N_19390);
nand U19781 (N_19781,N_19356,N_19384);
nor U19782 (N_19782,N_19456,N_19038);
and U19783 (N_19783,N_19466,N_19279);
nor U19784 (N_19784,N_19016,N_19428);
or U19785 (N_19785,N_19497,N_19452);
nor U19786 (N_19786,N_19199,N_19398);
nand U19787 (N_19787,N_19001,N_19082);
nor U19788 (N_19788,N_19043,N_19383);
and U19789 (N_19789,N_19399,N_19334);
nand U19790 (N_19790,N_19301,N_19222);
xor U19791 (N_19791,N_19207,N_19316);
nand U19792 (N_19792,N_19146,N_19160);
xnor U19793 (N_19793,N_19082,N_19025);
nand U19794 (N_19794,N_19049,N_19033);
or U19795 (N_19795,N_19487,N_19204);
and U19796 (N_19796,N_19354,N_19129);
nand U19797 (N_19797,N_19265,N_19145);
xor U19798 (N_19798,N_19173,N_19497);
xor U19799 (N_19799,N_19069,N_19354);
or U19800 (N_19800,N_19378,N_19331);
and U19801 (N_19801,N_19123,N_19273);
and U19802 (N_19802,N_19211,N_19379);
and U19803 (N_19803,N_19195,N_19081);
or U19804 (N_19804,N_19484,N_19394);
or U19805 (N_19805,N_19009,N_19453);
nor U19806 (N_19806,N_19242,N_19193);
or U19807 (N_19807,N_19088,N_19420);
or U19808 (N_19808,N_19107,N_19452);
nor U19809 (N_19809,N_19324,N_19202);
nor U19810 (N_19810,N_19191,N_19150);
or U19811 (N_19811,N_19130,N_19377);
and U19812 (N_19812,N_19485,N_19041);
and U19813 (N_19813,N_19331,N_19120);
nand U19814 (N_19814,N_19323,N_19344);
and U19815 (N_19815,N_19223,N_19325);
nand U19816 (N_19816,N_19466,N_19458);
nand U19817 (N_19817,N_19220,N_19461);
or U19818 (N_19818,N_19005,N_19068);
nor U19819 (N_19819,N_19369,N_19444);
nor U19820 (N_19820,N_19411,N_19455);
or U19821 (N_19821,N_19309,N_19190);
or U19822 (N_19822,N_19329,N_19417);
nand U19823 (N_19823,N_19024,N_19172);
and U19824 (N_19824,N_19218,N_19198);
or U19825 (N_19825,N_19327,N_19170);
nor U19826 (N_19826,N_19228,N_19473);
and U19827 (N_19827,N_19041,N_19424);
nor U19828 (N_19828,N_19202,N_19295);
nor U19829 (N_19829,N_19021,N_19345);
nand U19830 (N_19830,N_19152,N_19412);
and U19831 (N_19831,N_19448,N_19121);
nor U19832 (N_19832,N_19336,N_19407);
nor U19833 (N_19833,N_19050,N_19150);
or U19834 (N_19834,N_19114,N_19153);
nand U19835 (N_19835,N_19180,N_19297);
nand U19836 (N_19836,N_19336,N_19395);
nand U19837 (N_19837,N_19091,N_19471);
nand U19838 (N_19838,N_19186,N_19399);
or U19839 (N_19839,N_19442,N_19024);
and U19840 (N_19840,N_19398,N_19348);
nand U19841 (N_19841,N_19077,N_19254);
nor U19842 (N_19842,N_19201,N_19337);
nand U19843 (N_19843,N_19239,N_19285);
or U19844 (N_19844,N_19117,N_19411);
or U19845 (N_19845,N_19454,N_19016);
or U19846 (N_19846,N_19074,N_19144);
nand U19847 (N_19847,N_19114,N_19041);
or U19848 (N_19848,N_19223,N_19070);
or U19849 (N_19849,N_19263,N_19201);
nand U19850 (N_19850,N_19032,N_19497);
and U19851 (N_19851,N_19441,N_19340);
and U19852 (N_19852,N_19196,N_19014);
xnor U19853 (N_19853,N_19410,N_19095);
nand U19854 (N_19854,N_19360,N_19479);
nand U19855 (N_19855,N_19077,N_19134);
and U19856 (N_19856,N_19435,N_19173);
xor U19857 (N_19857,N_19270,N_19454);
xor U19858 (N_19858,N_19375,N_19464);
nor U19859 (N_19859,N_19029,N_19363);
or U19860 (N_19860,N_19471,N_19461);
xnor U19861 (N_19861,N_19376,N_19137);
or U19862 (N_19862,N_19154,N_19156);
or U19863 (N_19863,N_19198,N_19222);
nor U19864 (N_19864,N_19351,N_19233);
or U19865 (N_19865,N_19348,N_19340);
xor U19866 (N_19866,N_19294,N_19405);
nand U19867 (N_19867,N_19387,N_19023);
nand U19868 (N_19868,N_19440,N_19149);
xnor U19869 (N_19869,N_19051,N_19294);
and U19870 (N_19870,N_19066,N_19049);
or U19871 (N_19871,N_19382,N_19321);
or U19872 (N_19872,N_19339,N_19029);
xor U19873 (N_19873,N_19341,N_19364);
nor U19874 (N_19874,N_19091,N_19427);
nand U19875 (N_19875,N_19465,N_19453);
or U19876 (N_19876,N_19322,N_19006);
and U19877 (N_19877,N_19345,N_19351);
and U19878 (N_19878,N_19077,N_19030);
nand U19879 (N_19879,N_19349,N_19053);
and U19880 (N_19880,N_19197,N_19014);
nand U19881 (N_19881,N_19458,N_19075);
nand U19882 (N_19882,N_19486,N_19359);
nor U19883 (N_19883,N_19407,N_19192);
nor U19884 (N_19884,N_19086,N_19364);
and U19885 (N_19885,N_19203,N_19035);
nor U19886 (N_19886,N_19331,N_19215);
xor U19887 (N_19887,N_19290,N_19467);
nand U19888 (N_19888,N_19374,N_19436);
nor U19889 (N_19889,N_19010,N_19492);
nor U19890 (N_19890,N_19002,N_19167);
or U19891 (N_19891,N_19359,N_19047);
nor U19892 (N_19892,N_19012,N_19068);
nor U19893 (N_19893,N_19209,N_19076);
or U19894 (N_19894,N_19174,N_19462);
nor U19895 (N_19895,N_19221,N_19334);
nor U19896 (N_19896,N_19263,N_19216);
nor U19897 (N_19897,N_19056,N_19453);
xnor U19898 (N_19898,N_19264,N_19409);
xor U19899 (N_19899,N_19240,N_19338);
nand U19900 (N_19900,N_19439,N_19122);
xor U19901 (N_19901,N_19391,N_19209);
and U19902 (N_19902,N_19469,N_19306);
nand U19903 (N_19903,N_19267,N_19020);
nor U19904 (N_19904,N_19218,N_19002);
xor U19905 (N_19905,N_19231,N_19003);
or U19906 (N_19906,N_19235,N_19421);
and U19907 (N_19907,N_19387,N_19097);
or U19908 (N_19908,N_19465,N_19236);
and U19909 (N_19909,N_19044,N_19070);
and U19910 (N_19910,N_19365,N_19117);
nor U19911 (N_19911,N_19081,N_19447);
nand U19912 (N_19912,N_19279,N_19312);
and U19913 (N_19913,N_19218,N_19221);
xor U19914 (N_19914,N_19270,N_19334);
nor U19915 (N_19915,N_19209,N_19241);
and U19916 (N_19916,N_19098,N_19490);
xnor U19917 (N_19917,N_19194,N_19135);
or U19918 (N_19918,N_19490,N_19100);
nor U19919 (N_19919,N_19328,N_19247);
nor U19920 (N_19920,N_19410,N_19088);
and U19921 (N_19921,N_19318,N_19165);
nand U19922 (N_19922,N_19426,N_19254);
nor U19923 (N_19923,N_19233,N_19101);
or U19924 (N_19924,N_19265,N_19210);
nor U19925 (N_19925,N_19340,N_19251);
or U19926 (N_19926,N_19382,N_19472);
and U19927 (N_19927,N_19262,N_19267);
and U19928 (N_19928,N_19127,N_19076);
nor U19929 (N_19929,N_19039,N_19024);
xor U19930 (N_19930,N_19187,N_19159);
nand U19931 (N_19931,N_19371,N_19172);
nor U19932 (N_19932,N_19254,N_19232);
nor U19933 (N_19933,N_19210,N_19331);
nor U19934 (N_19934,N_19186,N_19419);
xnor U19935 (N_19935,N_19315,N_19472);
xnor U19936 (N_19936,N_19292,N_19497);
nand U19937 (N_19937,N_19397,N_19027);
nand U19938 (N_19938,N_19095,N_19012);
xor U19939 (N_19939,N_19018,N_19068);
nand U19940 (N_19940,N_19335,N_19399);
nand U19941 (N_19941,N_19464,N_19252);
xnor U19942 (N_19942,N_19092,N_19405);
nor U19943 (N_19943,N_19001,N_19168);
or U19944 (N_19944,N_19391,N_19300);
nand U19945 (N_19945,N_19168,N_19087);
nor U19946 (N_19946,N_19481,N_19065);
xnor U19947 (N_19947,N_19000,N_19110);
or U19948 (N_19948,N_19443,N_19143);
nor U19949 (N_19949,N_19165,N_19249);
nor U19950 (N_19950,N_19170,N_19137);
nand U19951 (N_19951,N_19075,N_19165);
nand U19952 (N_19952,N_19264,N_19020);
xor U19953 (N_19953,N_19361,N_19285);
xnor U19954 (N_19954,N_19156,N_19288);
nand U19955 (N_19955,N_19130,N_19163);
and U19956 (N_19956,N_19346,N_19361);
nand U19957 (N_19957,N_19393,N_19394);
nor U19958 (N_19958,N_19458,N_19423);
or U19959 (N_19959,N_19003,N_19078);
nor U19960 (N_19960,N_19254,N_19334);
xnor U19961 (N_19961,N_19032,N_19001);
or U19962 (N_19962,N_19326,N_19125);
xnor U19963 (N_19963,N_19167,N_19101);
and U19964 (N_19964,N_19000,N_19019);
xor U19965 (N_19965,N_19378,N_19469);
nand U19966 (N_19966,N_19266,N_19044);
or U19967 (N_19967,N_19172,N_19268);
or U19968 (N_19968,N_19453,N_19153);
nand U19969 (N_19969,N_19149,N_19279);
or U19970 (N_19970,N_19315,N_19105);
nor U19971 (N_19971,N_19284,N_19308);
nor U19972 (N_19972,N_19000,N_19351);
and U19973 (N_19973,N_19382,N_19437);
or U19974 (N_19974,N_19052,N_19089);
and U19975 (N_19975,N_19451,N_19387);
and U19976 (N_19976,N_19236,N_19090);
nand U19977 (N_19977,N_19227,N_19070);
xnor U19978 (N_19978,N_19167,N_19459);
nor U19979 (N_19979,N_19128,N_19146);
or U19980 (N_19980,N_19129,N_19426);
nor U19981 (N_19981,N_19315,N_19061);
nand U19982 (N_19982,N_19377,N_19151);
nor U19983 (N_19983,N_19488,N_19219);
nand U19984 (N_19984,N_19293,N_19349);
xor U19985 (N_19985,N_19308,N_19194);
nor U19986 (N_19986,N_19381,N_19144);
or U19987 (N_19987,N_19493,N_19452);
xnor U19988 (N_19988,N_19305,N_19206);
or U19989 (N_19989,N_19033,N_19045);
nand U19990 (N_19990,N_19253,N_19244);
and U19991 (N_19991,N_19328,N_19187);
or U19992 (N_19992,N_19001,N_19242);
or U19993 (N_19993,N_19182,N_19270);
nand U19994 (N_19994,N_19160,N_19117);
nor U19995 (N_19995,N_19225,N_19298);
or U19996 (N_19996,N_19180,N_19019);
nor U19997 (N_19997,N_19122,N_19129);
xor U19998 (N_19998,N_19306,N_19368);
nand U19999 (N_19999,N_19243,N_19421);
and U20000 (N_20000,N_19702,N_19721);
xnor U20001 (N_20001,N_19895,N_19736);
xnor U20002 (N_20002,N_19756,N_19598);
or U20003 (N_20003,N_19880,N_19913);
and U20004 (N_20004,N_19659,N_19796);
and U20005 (N_20005,N_19817,N_19653);
nor U20006 (N_20006,N_19690,N_19692);
and U20007 (N_20007,N_19576,N_19751);
nand U20008 (N_20008,N_19854,N_19818);
or U20009 (N_20009,N_19739,N_19514);
nor U20010 (N_20010,N_19633,N_19925);
and U20011 (N_20011,N_19816,N_19612);
nand U20012 (N_20012,N_19972,N_19681);
xor U20013 (N_20013,N_19984,N_19634);
and U20014 (N_20014,N_19503,N_19920);
and U20015 (N_20015,N_19559,N_19899);
or U20016 (N_20016,N_19539,N_19884);
or U20017 (N_20017,N_19752,N_19922);
or U20018 (N_20018,N_19955,N_19534);
xnor U20019 (N_20019,N_19630,N_19793);
nor U20020 (N_20020,N_19511,N_19757);
nand U20021 (N_20021,N_19778,N_19998);
or U20022 (N_20022,N_19629,N_19871);
xnor U20023 (N_20023,N_19932,N_19807);
and U20024 (N_20024,N_19996,N_19927);
nor U20025 (N_20025,N_19551,N_19640);
xnor U20026 (N_20026,N_19679,N_19620);
nand U20027 (N_20027,N_19815,N_19987);
xnor U20028 (N_20028,N_19574,N_19839);
and U20029 (N_20029,N_19621,N_19566);
and U20030 (N_20030,N_19542,N_19593);
or U20031 (N_20031,N_19768,N_19879);
nand U20032 (N_20032,N_19844,N_19905);
and U20033 (N_20033,N_19671,N_19767);
xor U20034 (N_20034,N_19892,N_19935);
nand U20035 (N_20035,N_19678,N_19637);
xnor U20036 (N_20036,N_19709,N_19942);
nor U20037 (N_20037,N_19952,N_19538);
xnor U20038 (N_20038,N_19744,N_19826);
xor U20039 (N_20039,N_19502,N_19575);
and U20040 (N_20040,N_19785,N_19657);
xnor U20041 (N_20041,N_19959,N_19587);
or U20042 (N_20042,N_19663,N_19532);
xor U20043 (N_20043,N_19779,N_19515);
nand U20044 (N_20044,N_19750,N_19792);
or U20045 (N_20045,N_19956,N_19774);
and U20046 (N_20046,N_19624,N_19572);
or U20047 (N_20047,N_19855,N_19706);
and U20048 (N_20048,N_19536,N_19990);
or U20049 (N_20049,N_19762,N_19594);
nand U20050 (N_20050,N_19582,N_19641);
xor U20051 (N_20051,N_19877,N_19921);
xor U20052 (N_20052,N_19609,N_19613);
nand U20053 (N_20053,N_19970,N_19896);
nand U20054 (N_20054,N_19909,N_19509);
and U20055 (N_20055,N_19766,N_19974);
and U20056 (N_20056,N_19527,N_19700);
nor U20057 (N_20057,N_19635,N_19686);
nor U20058 (N_20058,N_19810,N_19971);
nor U20059 (N_20059,N_19601,N_19628);
or U20060 (N_20060,N_19928,N_19869);
nand U20061 (N_20061,N_19872,N_19772);
and U20062 (N_20062,N_19724,N_19526);
and U20063 (N_20063,N_19851,N_19957);
nor U20064 (N_20064,N_19699,N_19507);
and U20065 (N_20065,N_19875,N_19760);
nor U20066 (N_20066,N_19558,N_19902);
xnor U20067 (N_20067,N_19623,N_19759);
or U20068 (N_20068,N_19619,N_19963);
nand U20069 (N_20069,N_19831,N_19941);
xnor U20070 (N_20070,N_19771,N_19936);
nand U20071 (N_20071,N_19652,N_19874);
xor U20072 (N_20072,N_19666,N_19830);
or U20073 (N_20073,N_19966,N_19517);
and U20074 (N_20074,N_19832,N_19660);
xor U20075 (N_20075,N_19632,N_19622);
nand U20076 (N_20076,N_19554,N_19876);
or U20077 (N_20077,N_19533,N_19821);
nor U20078 (N_20078,N_19579,N_19562);
nor U20079 (N_20079,N_19610,N_19898);
and U20080 (N_20080,N_19900,N_19791);
or U20081 (N_20081,N_19937,N_19662);
and U20082 (N_20082,N_19513,N_19933);
or U20083 (N_20083,N_19908,N_19833);
nor U20084 (N_20084,N_19697,N_19606);
nand U20085 (N_20085,N_19848,N_19518);
nand U20086 (N_20086,N_19856,N_19547);
and U20087 (N_20087,N_19599,N_19529);
nor U20088 (N_20088,N_19713,N_19853);
nand U20089 (N_20089,N_19967,N_19580);
and U20090 (N_20090,N_19703,N_19577);
nand U20091 (N_20091,N_19741,N_19746);
nor U20092 (N_20092,N_19638,N_19642);
nand U20093 (N_20093,N_19979,N_19894);
nand U20094 (N_20094,N_19790,N_19729);
and U20095 (N_20095,N_19858,N_19523);
or U20096 (N_20096,N_19591,N_19693);
or U20097 (N_20097,N_19893,N_19834);
xnor U20098 (N_20098,N_19584,N_19753);
nor U20099 (N_20099,N_19865,N_19688);
or U20100 (N_20100,N_19958,N_19983);
nand U20101 (N_20101,N_19737,N_19782);
and U20102 (N_20102,N_19573,N_19649);
nand U20103 (N_20103,N_19676,N_19835);
nor U20104 (N_20104,N_19545,N_19911);
and U20105 (N_20105,N_19596,N_19665);
nor U20106 (N_20106,N_19667,N_19720);
nor U20107 (N_20107,N_19516,N_19749);
nand U20108 (N_20108,N_19861,N_19951);
or U20109 (N_20109,N_19561,N_19560);
nand U20110 (N_20110,N_19565,N_19904);
xor U20111 (N_20111,N_19776,N_19930);
xnor U20112 (N_20112,N_19819,N_19543);
and U20113 (N_20113,N_19828,N_19647);
or U20114 (N_20114,N_19530,N_19969);
nor U20115 (N_20115,N_19891,N_19531);
xor U20116 (N_20116,N_19626,N_19578);
or U20117 (N_20117,N_19712,N_19730);
xor U20118 (N_20118,N_19801,N_19827);
nor U20119 (N_20119,N_19732,N_19748);
nor U20120 (N_20120,N_19814,N_19811);
or U20121 (N_20121,N_19675,N_19980);
or U20122 (N_20122,N_19975,N_19824);
nor U20123 (N_20123,N_19668,N_19780);
and U20124 (N_20124,N_19740,N_19687);
nor U20125 (N_20125,N_19803,N_19939);
nand U20126 (N_20126,N_19842,N_19581);
and U20127 (N_20127,N_19852,N_19643);
and U20128 (N_20128,N_19886,N_19696);
nand U20129 (N_20129,N_19655,N_19885);
xnor U20130 (N_20130,N_19617,N_19670);
nand U20131 (N_20131,N_19618,N_19938);
xor U20132 (N_20132,N_19995,N_19929);
and U20133 (N_20133,N_19999,N_19944);
nor U20134 (N_20134,N_19777,N_19781);
nand U20135 (N_20135,N_19717,N_19845);
or U20136 (N_20136,N_19590,N_19563);
and U20137 (N_20137,N_19520,N_19915);
nor U20138 (N_20138,N_19906,N_19631);
and U20139 (N_20139,N_19765,N_19548);
xnor U20140 (N_20140,N_19775,N_19718);
or U20141 (N_20141,N_19931,N_19537);
nand U20142 (N_20142,N_19889,N_19734);
xor U20143 (N_20143,N_19934,N_19866);
or U20144 (N_20144,N_19600,N_19683);
or U20145 (N_20145,N_19917,N_19604);
and U20146 (N_20146,N_19625,N_19754);
xnor U20147 (N_20147,N_19881,N_19727);
xor U20148 (N_20148,N_19962,N_19658);
nor U20149 (N_20149,N_19669,N_19564);
or U20150 (N_20150,N_19654,N_19639);
nand U20151 (N_20151,N_19950,N_19605);
xnor U20152 (N_20152,N_19924,N_19977);
nand U20153 (N_20153,N_19544,N_19627);
nor U20154 (N_20154,N_19812,N_19568);
and U20155 (N_20155,N_19820,N_19707);
and U20156 (N_20156,N_19747,N_19571);
nand U20157 (N_20157,N_19602,N_19673);
nor U20158 (N_20158,N_19809,N_19948);
xnor U20159 (N_20159,N_19714,N_19755);
nand U20160 (N_20160,N_19829,N_19661);
xnor U20161 (N_20161,N_19524,N_19731);
xor U20162 (N_20162,N_19910,N_19946);
nand U20163 (N_20163,N_19758,N_19773);
nand U20164 (N_20164,N_19680,N_19549);
nor U20165 (N_20165,N_19501,N_19505);
and U20166 (N_20166,N_19541,N_19822);
and U20167 (N_20167,N_19887,N_19918);
nand U20168 (N_20168,N_19556,N_19608);
xor U20169 (N_20169,N_19864,N_19570);
and U20170 (N_20170,N_19953,N_19764);
nor U20171 (N_20171,N_19795,N_19555);
nand U20172 (N_20172,N_19806,N_19888);
nand U20173 (N_20173,N_19636,N_19985);
xor U20174 (N_20174,N_19528,N_19973);
nand U20175 (N_20175,N_19651,N_19836);
nand U20176 (N_20176,N_19552,N_19850);
and U20177 (N_20177,N_19859,N_19823);
nor U20178 (N_20178,N_19677,N_19982);
and U20179 (N_20179,N_19698,N_19786);
nand U20180 (N_20180,N_19719,N_19849);
nor U20181 (N_20181,N_19770,N_19840);
or U20182 (N_20182,N_19802,N_19949);
and U20183 (N_20183,N_19607,N_19589);
nor U20184 (N_20184,N_19797,N_19728);
and U20185 (N_20185,N_19716,N_19926);
xor U20186 (N_20186,N_19592,N_19726);
nand U20187 (N_20187,N_19843,N_19711);
nor U20188 (N_20188,N_19689,N_19986);
and U20189 (N_20189,N_19997,N_19682);
or U20190 (N_20190,N_19912,N_19993);
xnor U20191 (N_20191,N_19868,N_19723);
xor U20192 (N_20192,N_19976,N_19540);
or U20193 (N_20193,N_19569,N_19787);
or U20194 (N_20194,N_19825,N_19883);
nand U20195 (N_20195,N_19783,N_19611);
nand U20196 (N_20196,N_19991,N_19837);
and U20197 (N_20197,N_19919,N_19616);
or U20198 (N_20198,N_19943,N_19512);
xor U20199 (N_20199,N_19738,N_19890);
and U20200 (N_20200,N_19788,N_19506);
or U20201 (N_20201,N_19954,N_19722);
and U20202 (N_20202,N_19901,N_19691);
xor U20203 (N_20203,N_19800,N_19743);
xor U20204 (N_20204,N_19557,N_19860);
nor U20205 (N_20205,N_19650,N_19794);
and U20206 (N_20206,N_19964,N_19978);
nor U20207 (N_20207,N_19525,N_19947);
nand U20208 (N_20208,N_19550,N_19704);
or U20209 (N_20209,N_19992,N_19870);
xor U20210 (N_20210,N_19546,N_19789);
nor U20211 (N_20211,N_19907,N_19586);
or U20212 (N_20212,N_19508,N_19672);
and U20213 (N_20213,N_19664,N_19857);
xor U20214 (N_20214,N_19603,N_19588);
or U20215 (N_20215,N_19994,N_19567);
nor U20216 (N_20216,N_19940,N_19945);
xnor U20217 (N_20217,N_19521,N_19808);
xnor U20218 (N_20218,N_19873,N_19583);
nand U20219 (N_20219,N_19656,N_19735);
xor U20220 (N_20220,N_19960,N_19715);
nand U20221 (N_20221,N_19614,N_19763);
or U20222 (N_20222,N_19916,N_19867);
nand U20223 (N_20223,N_19968,N_19914);
or U20224 (N_20224,N_19500,N_19644);
xor U20225 (N_20225,N_19701,N_19923);
and U20226 (N_20226,N_19847,N_19799);
or U20227 (N_20227,N_19897,N_19863);
or U20228 (N_20228,N_19798,N_19585);
nor U20229 (N_20229,N_19684,N_19841);
xor U20230 (N_20230,N_19745,N_19882);
and U20231 (N_20231,N_19903,N_19961);
nand U20232 (N_20232,N_19708,N_19805);
or U20233 (N_20233,N_19615,N_19674);
nand U20234 (N_20234,N_19761,N_19522);
nand U20235 (N_20235,N_19725,N_19742);
nor U20236 (N_20236,N_19784,N_19769);
xor U20237 (N_20237,N_19504,N_19535);
nand U20238 (N_20238,N_19510,N_19710);
and U20239 (N_20239,N_19846,N_19878);
and U20240 (N_20240,N_19553,N_19595);
xor U20241 (N_20241,N_19685,N_19813);
nand U20242 (N_20242,N_19981,N_19597);
and U20243 (N_20243,N_19965,N_19646);
nand U20244 (N_20244,N_19705,N_19838);
xnor U20245 (N_20245,N_19694,N_19988);
xor U20246 (N_20246,N_19648,N_19989);
nor U20247 (N_20247,N_19519,N_19695);
xnor U20248 (N_20248,N_19733,N_19862);
or U20249 (N_20249,N_19645,N_19804);
nand U20250 (N_20250,N_19942,N_19737);
nand U20251 (N_20251,N_19726,N_19865);
xnor U20252 (N_20252,N_19641,N_19521);
or U20253 (N_20253,N_19701,N_19907);
nor U20254 (N_20254,N_19882,N_19812);
nor U20255 (N_20255,N_19725,N_19629);
and U20256 (N_20256,N_19529,N_19564);
and U20257 (N_20257,N_19729,N_19837);
nor U20258 (N_20258,N_19663,N_19744);
and U20259 (N_20259,N_19982,N_19742);
and U20260 (N_20260,N_19915,N_19617);
nand U20261 (N_20261,N_19782,N_19699);
or U20262 (N_20262,N_19813,N_19731);
or U20263 (N_20263,N_19950,N_19861);
nand U20264 (N_20264,N_19956,N_19819);
xor U20265 (N_20265,N_19520,N_19726);
or U20266 (N_20266,N_19736,N_19708);
and U20267 (N_20267,N_19959,N_19840);
or U20268 (N_20268,N_19681,N_19912);
xor U20269 (N_20269,N_19693,N_19943);
nand U20270 (N_20270,N_19814,N_19776);
and U20271 (N_20271,N_19645,N_19868);
nand U20272 (N_20272,N_19918,N_19920);
or U20273 (N_20273,N_19552,N_19761);
or U20274 (N_20274,N_19997,N_19602);
xor U20275 (N_20275,N_19783,N_19598);
and U20276 (N_20276,N_19787,N_19688);
nand U20277 (N_20277,N_19573,N_19570);
and U20278 (N_20278,N_19870,N_19640);
and U20279 (N_20279,N_19894,N_19772);
and U20280 (N_20280,N_19930,N_19538);
xor U20281 (N_20281,N_19552,N_19730);
xor U20282 (N_20282,N_19601,N_19572);
and U20283 (N_20283,N_19627,N_19607);
nor U20284 (N_20284,N_19866,N_19987);
and U20285 (N_20285,N_19897,N_19548);
nand U20286 (N_20286,N_19995,N_19554);
xnor U20287 (N_20287,N_19739,N_19823);
xnor U20288 (N_20288,N_19706,N_19834);
nor U20289 (N_20289,N_19621,N_19655);
or U20290 (N_20290,N_19867,N_19850);
nand U20291 (N_20291,N_19625,N_19761);
nor U20292 (N_20292,N_19916,N_19523);
nor U20293 (N_20293,N_19725,N_19716);
nand U20294 (N_20294,N_19653,N_19535);
and U20295 (N_20295,N_19921,N_19611);
nor U20296 (N_20296,N_19849,N_19620);
nor U20297 (N_20297,N_19978,N_19693);
or U20298 (N_20298,N_19850,N_19879);
nand U20299 (N_20299,N_19784,N_19946);
xor U20300 (N_20300,N_19551,N_19973);
or U20301 (N_20301,N_19516,N_19792);
and U20302 (N_20302,N_19503,N_19598);
xnor U20303 (N_20303,N_19679,N_19598);
nand U20304 (N_20304,N_19857,N_19689);
nand U20305 (N_20305,N_19523,N_19997);
nand U20306 (N_20306,N_19948,N_19699);
and U20307 (N_20307,N_19831,N_19625);
nand U20308 (N_20308,N_19646,N_19595);
nand U20309 (N_20309,N_19545,N_19973);
nor U20310 (N_20310,N_19657,N_19712);
nand U20311 (N_20311,N_19571,N_19504);
nand U20312 (N_20312,N_19802,N_19912);
or U20313 (N_20313,N_19770,N_19742);
xnor U20314 (N_20314,N_19559,N_19585);
nand U20315 (N_20315,N_19795,N_19916);
nor U20316 (N_20316,N_19779,N_19728);
or U20317 (N_20317,N_19894,N_19741);
nor U20318 (N_20318,N_19862,N_19926);
xor U20319 (N_20319,N_19925,N_19962);
nor U20320 (N_20320,N_19854,N_19816);
and U20321 (N_20321,N_19956,N_19556);
and U20322 (N_20322,N_19570,N_19607);
nand U20323 (N_20323,N_19927,N_19854);
nand U20324 (N_20324,N_19952,N_19988);
xor U20325 (N_20325,N_19678,N_19977);
nand U20326 (N_20326,N_19585,N_19502);
or U20327 (N_20327,N_19669,N_19567);
nor U20328 (N_20328,N_19701,N_19556);
or U20329 (N_20329,N_19652,N_19772);
nor U20330 (N_20330,N_19867,N_19628);
nand U20331 (N_20331,N_19984,N_19963);
nand U20332 (N_20332,N_19865,N_19798);
and U20333 (N_20333,N_19916,N_19521);
or U20334 (N_20334,N_19983,N_19729);
nand U20335 (N_20335,N_19728,N_19884);
nor U20336 (N_20336,N_19743,N_19870);
or U20337 (N_20337,N_19914,N_19643);
nand U20338 (N_20338,N_19877,N_19852);
or U20339 (N_20339,N_19891,N_19529);
xor U20340 (N_20340,N_19504,N_19994);
nor U20341 (N_20341,N_19526,N_19663);
nand U20342 (N_20342,N_19504,N_19808);
and U20343 (N_20343,N_19508,N_19836);
nor U20344 (N_20344,N_19869,N_19531);
or U20345 (N_20345,N_19993,N_19511);
xnor U20346 (N_20346,N_19916,N_19522);
nor U20347 (N_20347,N_19560,N_19517);
xnor U20348 (N_20348,N_19667,N_19790);
or U20349 (N_20349,N_19595,N_19541);
and U20350 (N_20350,N_19906,N_19871);
nand U20351 (N_20351,N_19642,N_19778);
nand U20352 (N_20352,N_19844,N_19575);
xnor U20353 (N_20353,N_19596,N_19908);
xnor U20354 (N_20354,N_19937,N_19768);
xor U20355 (N_20355,N_19819,N_19713);
nor U20356 (N_20356,N_19567,N_19535);
and U20357 (N_20357,N_19929,N_19829);
nor U20358 (N_20358,N_19939,N_19662);
xor U20359 (N_20359,N_19806,N_19930);
and U20360 (N_20360,N_19801,N_19597);
nand U20361 (N_20361,N_19507,N_19771);
nor U20362 (N_20362,N_19871,N_19594);
or U20363 (N_20363,N_19550,N_19777);
xor U20364 (N_20364,N_19556,N_19663);
xor U20365 (N_20365,N_19773,N_19973);
nor U20366 (N_20366,N_19734,N_19725);
nor U20367 (N_20367,N_19502,N_19890);
nor U20368 (N_20368,N_19747,N_19699);
nand U20369 (N_20369,N_19863,N_19562);
xnor U20370 (N_20370,N_19992,N_19744);
nand U20371 (N_20371,N_19844,N_19799);
or U20372 (N_20372,N_19644,N_19803);
nand U20373 (N_20373,N_19831,N_19834);
nor U20374 (N_20374,N_19653,N_19663);
and U20375 (N_20375,N_19626,N_19541);
xnor U20376 (N_20376,N_19507,N_19894);
or U20377 (N_20377,N_19927,N_19749);
nor U20378 (N_20378,N_19777,N_19710);
and U20379 (N_20379,N_19744,N_19844);
nor U20380 (N_20380,N_19739,N_19737);
nor U20381 (N_20381,N_19573,N_19538);
nor U20382 (N_20382,N_19698,N_19759);
or U20383 (N_20383,N_19911,N_19775);
nor U20384 (N_20384,N_19856,N_19526);
or U20385 (N_20385,N_19591,N_19677);
xnor U20386 (N_20386,N_19922,N_19765);
nand U20387 (N_20387,N_19880,N_19918);
nor U20388 (N_20388,N_19557,N_19630);
xor U20389 (N_20389,N_19885,N_19634);
nor U20390 (N_20390,N_19704,N_19609);
nor U20391 (N_20391,N_19553,N_19522);
nor U20392 (N_20392,N_19660,N_19632);
nand U20393 (N_20393,N_19677,N_19981);
xnor U20394 (N_20394,N_19891,N_19690);
nand U20395 (N_20395,N_19968,N_19637);
and U20396 (N_20396,N_19732,N_19981);
xnor U20397 (N_20397,N_19740,N_19895);
or U20398 (N_20398,N_19960,N_19570);
xnor U20399 (N_20399,N_19947,N_19780);
or U20400 (N_20400,N_19540,N_19615);
nor U20401 (N_20401,N_19655,N_19577);
or U20402 (N_20402,N_19635,N_19574);
nor U20403 (N_20403,N_19677,N_19609);
and U20404 (N_20404,N_19914,N_19991);
nand U20405 (N_20405,N_19511,N_19562);
nor U20406 (N_20406,N_19863,N_19624);
or U20407 (N_20407,N_19616,N_19941);
nor U20408 (N_20408,N_19834,N_19805);
and U20409 (N_20409,N_19753,N_19850);
nand U20410 (N_20410,N_19975,N_19767);
and U20411 (N_20411,N_19916,N_19737);
xnor U20412 (N_20412,N_19942,N_19801);
xnor U20413 (N_20413,N_19950,N_19891);
or U20414 (N_20414,N_19788,N_19531);
or U20415 (N_20415,N_19657,N_19975);
and U20416 (N_20416,N_19683,N_19644);
and U20417 (N_20417,N_19980,N_19619);
or U20418 (N_20418,N_19970,N_19633);
nand U20419 (N_20419,N_19947,N_19649);
nor U20420 (N_20420,N_19909,N_19529);
and U20421 (N_20421,N_19726,N_19607);
or U20422 (N_20422,N_19605,N_19793);
xnor U20423 (N_20423,N_19773,N_19547);
nor U20424 (N_20424,N_19949,N_19983);
xnor U20425 (N_20425,N_19989,N_19517);
xnor U20426 (N_20426,N_19524,N_19555);
nand U20427 (N_20427,N_19756,N_19579);
nor U20428 (N_20428,N_19720,N_19776);
xnor U20429 (N_20429,N_19535,N_19735);
nor U20430 (N_20430,N_19793,N_19636);
or U20431 (N_20431,N_19695,N_19669);
xnor U20432 (N_20432,N_19629,N_19556);
nor U20433 (N_20433,N_19959,N_19821);
or U20434 (N_20434,N_19817,N_19965);
xnor U20435 (N_20435,N_19634,N_19947);
or U20436 (N_20436,N_19514,N_19506);
xnor U20437 (N_20437,N_19586,N_19859);
or U20438 (N_20438,N_19744,N_19753);
nand U20439 (N_20439,N_19993,N_19818);
or U20440 (N_20440,N_19680,N_19779);
nor U20441 (N_20441,N_19820,N_19701);
or U20442 (N_20442,N_19941,N_19759);
xor U20443 (N_20443,N_19878,N_19944);
nor U20444 (N_20444,N_19793,N_19503);
and U20445 (N_20445,N_19553,N_19816);
xor U20446 (N_20446,N_19657,N_19701);
or U20447 (N_20447,N_19785,N_19794);
xnor U20448 (N_20448,N_19731,N_19612);
nor U20449 (N_20449,N_19747,N_19982);
or U20450 (N_20450,N_19598,N_19623);
nor U20451 (N_20451,N_19715,N_19597);
nand U20452 (N_20452,N_19611,N_19922);
nor U20453 (N_20453,N_19929,N_19848);
nor U20454 (N_20454,N_19905,N_19517);
nor U20455 (N_20455,N_19950,N_19759);
nand U20456 (N_20456,N_19727,N_19927);
and U20457 (N_20457,N_19872,N_19688);
xor U20458 (N_20458,N_19613,N_19924);
or U20459 (N_20459,N_19975,N_19833);
or U20460 (N_20460,N_19922,N_19965);
xor U20461 (N_20461,N_19834,N_19684);
or U20462 (N_20462,N_19884,N_19864);
or U20463 (N_20463,N_19525,N_19653);
nor U20464 (N_20464,N_19680,N_19696);
nand U20465 (N_20465,N_19650,N_19635);
nor U20466 (N_20466,N_19957,N_19859);
xnor U20467 (N_20467,N_19974,N_19680);
or U20468 (N_20468,N_19565,N_19562);
nor U20469 (N_20469,N_19574,N_19744);
or U20470 (N_20470,N_19913,N_19988);
xnor U20471 (N_20471,N_19621,N_19933);
nor U20472 (N_20472,N_19986,N_19520);
nor U20473 (N_20473,N_19877,N_19534);
xnor U20474 (N_20474,N_19849,N_19781);
and U20475 (N_20475,N_19591,N_19614);
nand U20476 (N_20476,N_19670,N_19965);
xor U20477 (N_20477,N_19961,N_19724);
or U20478 (N_20478,N_19954,N_19581);
nor U20479 (N_20479,N_19717,N_19519);
and U20480 (N_20480,N_19974,N_19936);
nand U20481 (N_20481,N_19743,N_19803);
nand U20482 (N_20482,N_19513,N_19570);
and U20483 (N_20483,N_19900,N_19518);
or U20484 (N_20484,N_19645,N_19587);
or U20485 (N_20485,N_19994,N_19717);
nand U20486 (N_20486,N_19909,N_19676);
or U20487 (N_20487,N_19701,N_19683);
and U20488 (N_20488,N_19688,N_19759);
nand U20489 (N_20489,N_19519,N_19942);
nand U20490 (N_20490,N_19913,N_19763);
nand U20491 (N_20491,N_19735,N_19930);
xnor U20492 (N_20492,N_19639,N_19850);
nand U20493 (N_20493,N_19631,N_19963);
xnor U20494 (N_20494,N_19746,N_19618);
nand U20495 (N_20495,N_19512,N_19662);
or U20496 (N_20496,N_19572,N_19791);
nor U20497 (N_20497,N_19783,N_19633);
nand U20498 (N_20498,N_19857,N_19969);
nand U20499 (N_20499,N_19607,N_19639);
nand U20500 (N_20500,N_20384,N_20490);
nand U20501 (N_20501,N_20162,N_20426);
nand U20502 (N_20502,N_20050,N_20471);
xor U20503 (N_20503,N_20337,N_20168);
xor U20504 (N_20504,N_20335,N_20341);
xor U20505 (N_20505,N_20183,N_20416);
or U20506 (N_20506,N_20496,N_20425);
or U20507 (N_20507,N_20404,N_20339);
nor U20508 (N_20508,N_20305,N_20418);
nor U20509 (N_20509,N_20330,N_20027);
or U20510 (N_20510,N_20199,N_20097);
nor U20511 (N_20511,N_20234,N_20143);
nand U20512 (N_20512,N_20185,N_20212);
xor U20513 (N_20513,N_20283,N_20282);
or U20514 (N_20514,N_20014,N_20118);
or U20515 (N_20515,N_20427,N_20391);
and U20516 (N_20516,N_20035,N_20235);
or U20517 (N_20517,N_20280,N_20279);
or U20518 (N_20518,N_20026,N_20174);
nand U20519 (N_20519,N_20262,N_20211);
nor U20520 (N_20520,N_20184,N_20138);
and U20521 (N_20521,N_20017,N_20463);
nand U20522 (N_20522,N_20196,N_20030);
nand U20523 (N_20523,N_20344,N_20444);
and U20524 (N_20524,N_20461,N_20170);
xor U20525 (N_20525,N_20137,N_20166);
xor U20526 (N_20526,N_20289,N_20311);
xor U20527 (N_20527,N_20260,N_20160);
or U20528 (N_20528,N_20086,N_20098);
or U20529 (N_20529,N_20225,N_20263);
or U20530 (N_20530,N_20251,N_20328);
nand U20531 (N_20531,N_20356,N_20077);
or U20532 (N_20532,N_20308,N_20476);
and U20533 (N_20533,N_20430,N_20245);
nor U20534 (N_20534,N_20049,N_20271);
nor U20535 (N_20535,N_20150,N_20329);
nor U20536 (N_20536,N_20304,N_20039);
nor U20537 (N_20537,N_20291,N_20421);
nor U20538 (N_20538,N_20317,N_20115);
nand U20539 (N_20539,N_20024,N_20277);
nand U20540 (N_20540,N_20132,N_20075);
xor U20541 (N_20541,N_20470,N_20462);
nand U20542 (N_20542,N_20290,N_20485);
and U20543 (N_20543,N_20479,N_20101);
xor U20544 (N_20544,N_20422,N_20415);
nor U20545 (N_20545,N_20372,N_20197);
or U20546 (N_20546,N_20355,N_20210);
nand U20547 (N_20547,N_20071,N_20434);
xor U20548 (N_20548,N_20414,N_20207);
nand U20549 (N_20549,N_20056,N_20497);
and U20550 (N_20550,N_20413,N_20440);
nor U20551 (N_20551,N_20145,N_20193);
or U20552 (N_20552,N_20453,N_20043);
xnor U20553 (N_20553,N_20059,N_20257);
xor U20554 (N_20554,N_20127,N_20238);
nand U20555 (N_20555,N_20406,N_20319);
or U20556 (N_20556,N_20085,N_20468);
or U20557 (N_20557,N_20227,N_20200);
nor U20558 (N_20558,N_20078,N_20365);
nor U20559 (N_20559,N_20094,N_20044);
xnor U20560 (N_20560,N_20457,N_20155);
xnor U20561 (N_20561,N_20134,N_20186);
nor U20562 (N_20562,N_20424,N_20009);
nor U20563 (N_20563,N_20111,N_20057);
nand U20564 (N_20564,N_20405,N_20410);
or U20565 (N_20565,N_20036,N_20491);
nand U20566 (N_20566,N_20403,N_20368);
or U20567 (N_20567,N_20040,N_20108);
or U20568 (N_20568,N_20073,N_20128);
nor U20569 (N_20569,N_20306,N_20272);
nor U20570 (N_20570,N_20171,N_20109);
nand U20571 (N_20571,N_20439,N_20366);
and U20572 (N_20572,N_20361,N_20130);
xor U20573 (N_20573,N_20327,N_20244);
xnor U20574 (N_20574,N_20480,N_20489);
and U20575 (N_20575,N_20275,N_20045);
nand U20576 (N_20576,N_20343,N_20449);
xnor U20577 (N_20577,N_20437,N_20089);
and U20578 (N_20578,N_20158,N_20229);
and U20579 (N_20579,N_20123,N_20438);
nand U20580 (N_20580,N_20222,N_20103);
and U20581 (N_20581,N_20205,N_20250);
and U20582 (N_20582,N_20374,N_20081);
nand U20583 (N_20583,N_20446,N_20218);
nand U20584 (N_20584,N_20013,N_20357);
xor U20585 (N_20585,N_20003,N_20495);
nand U20586 (N_20586,N_20322,N_20249);
and U20587 (N_20587,N_20258,N_20006);
xnor U20588 (N_20588,N_20239,N_20389);
xnor U20589 (N_20589,N_20347,N_20002);
nor U20590 (N_20590,N_20012,N_20072);
nor U20591 (N_20591,N_20467,N_20033);
nor U20592 (N_20592,N_20063,N_20455);
or U20593 (N_20593,N_20448,N_20004);
or U20594 (N_20594,N_20248,N_20346);
nand U20595 (N_20595,N_20396,N_20302);
nor U20596 (N_20596,N_20371,N_20386);
nor U20597 (N_20597,N_20058,N_20061);
nor U20598 (N_20598,N_20079,N_20408);
and U20599 (N_20599,N_20474,N_20393);
nand U20600 (N_20600,N_20092,N_20281);
or U20601 (N_20601,N_20129,N_20095);
xnor U20602 (N_20602,N_20140,N_20454);
xnor U20603 (N_20603,N_20146,N_20215);
xnor U20604 (N_20604,N_20298,N_20019);
and U20605 (N_20605,N_20029,N_20164);
and U20606 (N_20606,N_20149,N_20090);
or U20607 (N_20607,N_20333,N_20312);
nor U20608 (N_20608,N_20436,N_20219);
nand U20609 (N_20609,N_20373,N_20267);
nor U20610 (N_20610,N_20053,N_20294);
nand U20611 (N_20611,N_20392,N_20156);
or U20612 (N_20612,N_20390,N_20121);
nand U20613 (N_20613,N_20214,N_20435);
or U20614 (N_20614,N_20323,N_20142);
and U20615 (N_20615,N_20202,N_20032);
nor U20616 (N_20616,N_20379,N_20301);
or U20617 (N_20617,N_20240,N_20124);
xnor U20618 (N_20618,N_20313,N_20482);
nand U20619 (N_20619,N_20131,N_20034);
and U20620 (N_20620,N_20175,N_20412);
or U20621 (N_20621,N_20220,N_20233);
or U20622 (N_20622,N_20102,N_20120);
nand U20623 (N_20623,N_20255,N_20028);
nor U20624 (N_20624,N_20377,N_20052);
and U20625 (N_20625,N_20342,N_20070);
and U20626 (N_20626,N_20402,N_20252);
xnor U20627 (N_20627,N_20083,N_20181);
xnor U20628 (N_20628,N_20278,N_20483);
xnor U20629 (N_20629,N_20189,N_20498);
nand U20630 (N_20630,N_20064,N_20069);
nand U20631 (N_20631,N_20400,N_20008);
xnor U20632 (N_20632,N_20314,N_20213);
or U20633 (N_20633,N_20242,N_20318);
nand U20634 (N_20634,N_20241,N_20025);
or U20635 (N_20635,N_20286,N_20338);
xnor U20636 (N_20636,N_20484,N_20100);
nand U20637 (N_20637,N_20472,N_20493);
nor U20638 (N_20638,N_20190,N_20136);
xnor U20639 (N_20639,N_20292,N_20096);
and U20640 (N_20640,N_20080,N_20091);
or U20641 (N_20641,N_20221,N_20180);
nor U20642 (N_20642,N_20261,N_20253);
nor U20643 (N_20643,N_20288,N_20477);
xnor U20644 (N_20644,N_20209,N_20047);
nor U20645 (N_20645,N_20217,N_20297);
or U20646 (N_20646,N_20487,N_20375);
nand U20647 (N_20647,N_20432,N_20176);
nor U20648 (N_20648,N_20481,N_20456);
or U20649 (N_20649,N_20246,N_20179);
or U20650 (N_20650,N_20107,N_20352);
and U20651 (N_20651,N_20119,N_20451);
nand U20652 (N_20652,N_20104,N_20144);
and U20653 (N_20653,N_20216,N_20247);
nor U20654 (N_20654,N_20037,N_20354);
xnor U20655 (N_20655,N_20324,N_20074);
nand U20656 (N_20656,N_20206,N_20204);
nand U20657 (N_20657,N_20362,N_20165);
and U20658 (N_20658,N_20203,N_20345);
xnor U20659 (N_20659,N_20237,N_20316);
nor U20660 (N_20660,N_20178,N_20106);
xnor U20661 (N_20661,N_20122,N_20125);
nand U20662 (N_20662,N_20062,N_20296);
and U20663 (N_20663,N_20000,N_20023);
xor U20664 (N_20664,N_20182,N_20154);
and U20665 (N_20665,N_20381,N_20151);
and U20666 (N_20666,N_20147,N_20167);
xor U20667 (N_20667,N_20208,N_20010);
xor U20668 (N_20668,N_20363,N_20172);
and U20669 (N_20669,N_20082,N_20236);
nand U20670 (N_20670,N_20159,N_20460);
and U20671 (N_20671,N_20370,N_20041);
or U20672 (N_20672,N_20114,N_20116);
xor U20673 (N_20673,N_20177,N_20011);
or U20674 (N_20674,N_20423,N_20016);
or U20675 (N_20675,N_20015,N_20494);
and U20676 (N_20676,N_20135,N_20420);
nor U20677 (N_20677,N_20042,N_20048);
nor U20678 (N_20678,N_20465,N_20473);
or U20679 (N_20679,N_20407,N_20265);
or U20680 (N_20680,N_20228,N_20350);
xnor U20681 (N_20681,N_20163,N_20287);
xnor U20682 (N_20682,N_20411,N_20469);
nand U20683 (N_20683,N_20088,N_20431);
xor U20684 (N_20684,N_20452,N_20068);
nor U20685 (N_20685,N_20447,N_20285);
or U20686 (N_20686,N_20117,N_20266);
and U20687 (N_20687,N_20325,N_20232);
and U20688 (N_20688,N_20488,N_20099);
or U20689 (N_20689,N_20274,N_20051);
or U20690 (N_20690,N_20020,N_20360);
nand U20691 (N_20691,N_20284,N_20169);
and U20692 (N_20692,N_20334,N_20367);
and U20693 (N_20693,N_20105,N_20055);
nor U20694 (N_20694,N_20340,N_20351);
or U20695 (N_20695,N_20409,N_20398);
nor U20696 (N_20696,N_20417,N_20307);
xnor U20697 (N_20697,N_20359,N_20475);
xor U20698 (N_20698,N_20348,N_20331);
nand U20699 (N_20699,N_20349,N_20152);
xnor U20700 (N_20700,N_20445,N_20065);
nor U20701 (N_20701,N_20067,N_20038);
nor U20702 (N_20702,N_20022,N_20388);
nor U20703 (N_20703,N_20126,N_20459);
xor U20704 (N_20704,N_20192,N_20315);
and U20705 (N_20705,N_20464,N_20397);
xor U20706 (N_20706,N_20259,N_20066);
or U20707 (N_20707,N_20358,N_20401);
xnor U20708 (N_20708,N_20383,N_20376);
or U20709 (N_20709,N_20054,N_20458);
and U20710 (N_20710,N_20187,N_20076);
nand U20711 (N_20711,N_20093,N_20326);
nand U20712 (N_20712,N_20450,N_20466);
or U20713 (N_20713,N_20223,N_20254);
xnor U20714 (N_20714,N_20226,N_20139);
and U20715 (N_20715,N_20492,N_20478);
nand U20716 (N_20716,N_20441,N_20320);
xnor U20717 (N_20717,N_20382,N_20194);
nand U20718 (N_20718,N_20191,N_20007);
nand U20719 (N_20719,N_20195,N_20110);
nand U20720 (N_20720,N_20005,N_20295);
or U20721 (N_20721,N_20224,N_20428);
and U20722 (N_20722,N_20161,N_20332);
or U20723 (N_20723,N_20031,N_20364);
nor U20724 (N_20724,N_20443,N_20273);
nor U20725 (N_20725,N_20188,N_20369);
xnor U20726 (N_20726,N_20087,N_20157);
xnor U20727 (N_20727,N_20113,N_20153);
nor U20728 (N_20728,N_20300,N_20310);
and U20729 (N_20729,N_20353,N_20433);
xnor U20730 (N_20730,N_20084,N_20378);
nor U20731 (N_20731,N_20380,N_20018);
or U20732 (N_20732,N_20231,N_20395);
nor U20733 (N_20733,N_20399,N_20173);
and U20734 (N_20734,N_20309,N_20429);
and U20735 (N_20735,N_20419,N_20269);
xnor U20736 (N_20736,N_20387,N_20499);
xnor U20737 (N_20737,N_20268,N_20385);
nand U20738 (N_20738,N_20112,N_20276);
or U20739 (N_20739,N_20442,N_20133);
and U20740 (N_20740,N_20060,N_20394);
or U20741 (N_20741,N_20001,N_20230);
nand U20742 (N_20742,N_20198,N_20148);
nand U20743 (N_20743,N_20046,N_20270);
and U20744 (N_20744,N_20299,N_20201);
nand U20745 (N_20745,N_20256,N_20303);
and U20746 (N_20746,N_20021,N_20243);
xnor U20747 (N_20747,N_20264,N_20336);
or U20748 (N_20748,N_20141,N_20293);
xor U20749 (N_20749,N_20321,N_20486);
and U20750 (N_20750,N_20397,N_20119);
nand U20751 (N_20751,N_20398,N_20049);
nand U20752 (N_20752,N_20225,N_20135);
and U20753 (N_20753,N_20346,N_20225);
nand U20754 (N_20754,N_20144,N_20472);
nor U20755 (N_20755,N_20136,N_20022);
and U20756 (N_20756,N_20205,N_20251);
or U20757 (N_20757,N_20497,N_20350);
nor U20758 (N_20758,N_20245,N_20429);
nand U20759 (N_20759,N_20280,N_20375);
xnor U20760 (N_20760,N_20162,N_20218);
or U20761 (N_20761,N_20354,N_20384);
xor U20762 (N_20762,N_20401,N_20314);
nor U20763 (N_20763,N_20076,N_20266);
nand U20764 (N_20764,N_20357,N_20491);
nor U20765 (N_20765,N_20488,N_20225);
xnor U20766 (N_20766,N_20044,N_20098);
or U20767 (N_20767,N_20270,N_20050);
or U20768 (N_20768,N_20181,N_20256);
xnor U20769 (N_20769,N_20293,N_20349);
or U20770 (N_20770,N_20020,N_20461);
nor U20771 (N_20771,N_20440,N_20110);
nand U20772 (N_20772,N_20132,N_20055);
and U20773 (N_20773,N_20366,N_20297);
xnor U20774 (N_20774,N_20044,N_20323);
and U20775 (N_20775,N_20243,N_20463);
nand U20776 (N_20776,N_20271,N_20402);
and U20777 (N_20777,N_20000,N_20399);
and U20778 (N_20778,N_20270,N_20025);
or U20779 (N_20779,N_20175,N_20373);
or U20780 (N_20780,N_20109,N_20352);
xor U20781 (N_20781,N_20073,N_20223);
xor U20782 (N_20782,N_20153,N_20047);
xor U20783 (N_20783,N_20477,N_20322);
and U20784 (N_20784,N_20398,N_20217);
and U20785 (N_20785,N_20230,N_20247);
or U20786 (N_20786,N_20307,N_20005);
and U20787 (N_20787,N_20302,N_20426);
nand U20788 (N_20788,N_20419,N_20404);
xor U20789 (N_20789,N_20189,N_20066);
or U20790 (N_20790,N_20162,N_20241);
or U20791 (N_20791,N_20085,N_20209);
nor U20792 (N_20792,N_20201,N_20343);
and U20793 (N_20793,N_20279,N_20314);
nand U20794 (N_20794,N_20140,N_20132);
or U20795 (N_20795,N_20407,N_20126);
xor U20796 (N_20796,N_20368,N_20178);
nand U20797 (N_20797,N_20288,N_20108);
and U20798 (N_20798,N_20019,N_20284);
and U20799 (N_20799,N_20265,N_20221);
xor U20800 (N_20800,N_20169,N_20213);
or U20801 (N_20801,N_20160,N_20133);
and U20802 (N_20802,N_20384,N_20152);
xnor U20803 (N_20803,N_20319,N_20114);
xnor U20804 (N_20804,N_20450,N_20110);
nor U20805 (N_20805,N_20041,N_20198);
nand U20806 (N_20806,N_20187,N_20400);
xor U20807 (N_20807,N_20276,N_20153);
and U20808 (N_20808,N_20389,N_20007);
and U20809 (N_20809,N_20114,N_20381);
and U20810 (N_20810,N_20341,N_20203);
nor U20811 (N_20811,N_20494,N_20378);
nand U20812 (N_20812,N_20186,N_20031);
and U20813 (N_20813,N_20255,N_20306);
xor U20814 (N_20814,N_20282,N_20005);
and U20815 (N_20815,N_20043,N_20143);
nand U20816 (N_20816,N_20075,N_20307);
and U20817 (N_20817,N_20472,N_20102);
xnor U20818 (N_20818,N_20260,N_20318);
nor U20819 (N_20819,N_20156,N_20440);
xor U20820 (N_20820,N_20106,N_20071);
or U20821 (N_20821,N_20130,N_20395);
nor U20822 (N_20822,N_20429,N_20336);
nand U20823 (N_20823,N_20196,N_20342);
or U20824 (N_20824,N_20341,N_20466);
xor U20825 (N_20825,N_20157,N_20373);
nor U20826 (N_20826,N_20070,N_20217);
nand U20827 (N_20827,N_20166,N_20331);
xnor U20828 (N_20828,N_20456,N_20362);
nor U20829 (N_20829,N_20178,N_20268);
and U20830 (N_20830,N_20096,N_20348);
or U20831 (N_20831,N_20336,N_20403);
and U20832 (N_20832,N_20496,N_20172);
xnor U20833 (N_20833,N_20494,N_20409);
xnor U20834 (N_20834,N_20102,N_20327);
and U20835 (N_20835,N_20098,N_20033);
nand U20836 (N_20836,N_20345,N_20354);
and U20837 (N_20837,N_20002,N_20000);
or U20838 (N_20838,N_20013,N_20422);
and U20839 (N_20839,N_20256,N_20000);
xor U20840 (N_20840,N_20225,N_20102);
or U20841 (N_20841,N_20313,N_20132);
nor U20842 (N_20842,N_20283,N_20227);
or U20843 (N_20843,N_20134,N_20331);
xnor U20844 (N_20844,N_20456,N_20014);
xor U20845 (N_20845,N_20211,N_20487);
or U20846 (N_20846,N_20393,N_20278);
or U20847 (N_20847,N_20073,N_20116);
and U20848 (N_20848,N_20425,N_20348);
nor U20849 (N_20849,N_20307,N_20189);
nand U20850 (N_20850,N_20474,N_20239);
nor U20851 (N_20851,N_20021,N_20147);
or U20852 (N_20852,N_20293,N_20089);
or U20853 (N_20853,N_20203,N_20013);
nand U20854 (N_20854,N_20017,N_20057);
xor U20855 (N_20855,N_20247,N_20368);
or U20856 (N_20856,N_20011,N_20202);
nand U20857 (N_20857,N_20268,N_20211);
nor U20858 (N_20858,N_20465,N_20042);
nand U20859 (N_20859,N_20202,N_20431);
nor U20860 (N_20860,N_20173,N_20401);
and U20861 (N_20861,N_20266,N_20428);
and U20862 (N_20862,N_20172,N_20006);
xnor U20863 (N_20863,N_20382,N_20192);
and U20864 (N_20864,N_20116,N_20193);
or U20865 (N_20865,N_20422,N_20042);
nor U20866 (N_20866,N_20048,N_20415);
nor U20867 (N_20867,N_20437,N_20384);
nand U20868 (N_20868,N_20234,N_20067);
and U20869 (N_20869,N_20419,N_20322);
xor U20870 (N_20870,N_20060,N_20129);
or U20871 (N_20871,N_20217,N_20091);
or U20872 (N_20872,N_20188,N_20147);
nand U20873 (N_20873,N_20371,N_20405);
xor U20874 (N_20874,N_20069,N_20326);
nand U20875 (N_20875,N_20394,N_20427);
nand U20876 (N_20876,N_20294,N_20395);
or U20877 (N_20877,N_20251,N_20394);
xor U20878 (N_20878,N_20247,N_20488);
or U20879 (N_20879,N_20241,N_20371);
and U20880 (N_20880,N_20079,N_20316);
and U20881 (N_20881,N_20440,N_20313);
xnor U20882 (N_20882,N_20105,N_20040);
or U20883 (N_20883,N_20099,N_20176);
nand U20884 (N_20884,N_20495,N_20155);
nand U20885 (N_20885,N_20119,N_20357);
nor U20886 (N_20886,N_20056,N_20365);
xnor U20887 (N_20887,N_20363,N_20238);
nor U20888 (N_20888,N_20181,N_20012);
nor U20889 (N_20889,N_20026,N_20437);
or U20890 (N_20890,N_20224,N_20122);
or U20891 (N_20891,N_20467,N_20021);
or U20892 (N_20892,N_20292,N_20293);
nor U20893 (N_20893,N_20132,N_20149);
nand U20894 (N_20894,N_20083,N_20332);
xor U20895 (N_20895,N_20291,N_20013);
or U20896 (N_20896,N_20190,N_20079);
nand U20897 (N_20897,N_20215,N_20095);
nor U20898 (N_20898,N_20195,N_20383);
or U20899 (N_20899,N_20426,N_20180);
and U20900 (N_20900,N_20004,N_20322);
xnor U20901 (N_20901,N_20111,N_20376);
nor U20902 (N_20902,N_20318,N_20445);
nor U20903 (N_20903,N_20406,N_20182);
nor U20904 (N_20904,N_20263,N_20182);
xor U20905 (N_20905,N_20204,N_20114);
or U20906 (N_20906,N_20099,N_20344);
nor U20907 (N_20907,N_20496,N_20247);
nand U20908 (N_20908,N_20061,N_20480);
nor U20909 (N_20909,N_20488,N_20312);
nand U20910 (N_20910,N_20095,N_20007);
or U20911 (N_20911,N_20179,N_20204);
xnor U20912 (N_20912,N_20226,N_20220);
or U20913 (N_20913,N_20063,N_20183);
xor U20914 (N_20914,N_20085,N_20462);
nand U20915 (N_20915,N_20064,N_20284);
and U20916 (N_20916,N_20439,N_20029);
nand U20917 (N_20917,N_20419,N_20434);
nor U20918 (N_20918,N_20031,N_20075);
nand U20919 (N_20919,N_20257,N_20427);
xor U20920 (N_20920,N_20093,N_20428);
nand U20921 (N_20921,N_20284,N_20232);
or U20922 (N_20922,N_20308,N_20378);
nand U20923 (N_20923,N_20340,N_20179);
nand U20924 (N_20924,N_20134,N_20108);
nor U20925 (N_20925,N_20150,N_20087);
and U20926 (N_20926,N_20130,N_20127);
nand U20927 (N_20927,N_20249,N_20426);
nand U20928 (N_20928,N_20084,N_20384);
xor U20929 (N_20929,N_20168,N_20278);
nor U20930 (N_20930,N_20305,N_20031);
nor U20931 (N_20931,N_20048,N_20254);
or U20932 (N_20932,N_20305,N_20436);
and U20933 (N_20933,N_20441,N_20063);
or U20934 (N_20934,N_20197,N_20260);
xor U20935 (N_20935,N_20495,N_20270);
nor U20936 (N_20936,N_20097,N_20496);
or U20937 (N_20937,N_20462,N_20324);
and U20938 (N_20938,N_20171,N_20005);
nor U20939 (N_20939,N_20445,N_20248);
nand U20940 (N_20940,N_20444,N_20303);
xnor U20941 (N_20941,N_20384,N_20429);
and U20942 (N_20942,N_20464,N_20169);
nand U20943 (N_20943,N_20147,N_20389);
or U20944 (N_20944,N_20305,N_20460);
nand U20945 (N_20945,N_20038,N_20404);
or U20946 (N_20946,N_20029,N_20392);
nor U20947 (N_20947,N_20174,N_20479);
xnor U20948 (N_20948,N_20128,N_20458);
nand U20949 (N_20949,N_20037,N_20452);
nor U20950 (N_20950,N_20275,N_20149);
xor U20951 (N_20951,N_20141,N_20285);
xnor U20952 (N_20952,N_20206,N_20205);
nor U20953 (N_20953,N_20370,N_20155);
nand U20954 (N_20954,N_20238,N_20489);
nor U20955 (N_20955,N_20347,N_20083);
and U20956 (N_20956,N_20347,N_20205);
nand U20957 (N_20957,N_20346,N_20411);
nand U20958 (N_20958,N_20430,N_20271);
xnor U20959 (N_20959,N_20353,N_20425);
nand U20960 (N_20960,N_20442,N_20253);
nand U20961 (N_20961,N_20385,N_20051);
and U20962 (N_20962,N_20382,N_20369);
nor U20963 (N_20963,N_20092,N_20253);
nor U20964 (N_20964,N_20436,N_20094);
nand U20965 (N_20965,N_20470,N_20295);
nand U20966 (N_20966,N_20381,N_20411);
xnor U20967 (N_20967,N_20214,N_20099);
and U20968 (N_20968,N_20347,N_20055);
nand U20969 (N_20969,N_20311,N_20472);
or U20970 (N_20970,N_20071,N_20039);
xor U20971 (N_20971,N_20072,N_20200);
xor U20972 (N_20972,N_20211,N_20026);
nand U20973 (N_20973,N_20429,N_20399);
and U20974 (N_20974,N_20212,N_20026);
nand U20975 (N_20975,N_20021,N_20181);
or U20976 (N_20976,N_20011,N_20496);
nand U20977 (N_20977,N_20238,N_20180);
nor U20978 (N_20978,N_20411,N_20440);
or U20979 (N_20979,N_20217,N_20239);
or U20980 (N_20980,N_20177,N_20468);
and U20981 (N_20981,N_20301,N_20199);
xor U20982 (N_20982,N_20228,N_20229);
nor U20983 (N_20983,N_20074,N_20457);
nor U20984 (N_20984,N_20140,N_20259);
xnor U20985 (N_20985,N_20469,N_20492);
or U20986 (N_20986,N_20145,N_20167);
nand U20987 (N_20987,N_20124,N_20398);
xor U20988 (N_20988,N_20343,N_20126);
xnor U20989 (N_20989,N_20424,N_20133);
or U20990 (N_20990,N_20069,N_20223);
nor U20991 (N_20991,N_20303,N_20451);
nand U20992 (N_20992,N_20265,N_20018);
or U20993 (N_20993,N_20362,N_20227);
and U20994 (N_20994,N_20169,N_20417);
nand U20995 (N_20995,N_20453,N_20109);
xor U20996 (N_20996,N_20430,N_20164);
or U20997 (N_20997,N_20418,N_20480);
xnor U20998 (N_20998,N_20166,N_20343);
xnor U20999 (N_20999,N_20478,N_20320);
and U21000 (N_21000,N_20956,N_20504);
or U21001 (N_21001,N_20680,N_20662);
and U21002 (N_21002,N_20694,N_20926);
or U21003 (N_21003,N_20549,N_20715);
nand U21004 (N_21004,N_20743,N_20897);
and U21005 (N_21005,N_20991,N_20859);
nor U21006 (N_21006,N_20821,N_20790);
xnor U21007 (N_21007,N_20669,N_20966);
and U21008 (N_21008,N_20634,N_20577);
nor U21009 (N_21009,N_20880,N_20614);
xor U21010 (N_21010,N_20685,N_20686);
nand U21011 (N_21011,N_20878,N_20898);
nand U21012 (N_21012,N_20633,N_20871);
and U21013 (N_21013,N_20709,N_20954);
or U21014 (N_21014,N_20908,N_20617);
or U21015 (N_21015,N_20658,N_20856);
and U21016 (N_21016,N_20759,N_20811);
or U21017 (N_21017,N_20713,N_20995);
or U21018 (N_21018,N_20833,N_20585);
and U21019 (N_21019,N_20844,N_20822);
nor U21020 (N_21020,N_20712,N_20719);
nor U21021 (N_21021,N_20944,N_20987);
nor U21022 (N_21022,N_20788,N_20802);
nor U21023 (N_21023,N_20730,N_20544);
or U21024 (N_21024,N_20762,N_20969);
nand U21025 (N_21025,N_20884,N_20541);
xor U21026 (N_21026,N_20665,N_20657);
nand U21027 (N_21027,N_20936,N_20958);
and U21028 (N_21028,N_20704,N_20804);
nand U21029 (N_21029,N_20621,N_20824);
nor U21030 (N_21030,N_20800,N_20953);
or U21031 (N_21031,N_20984,N_20961);
xor U21032 (N_21032,N_20866,N_20870);
nand U21033 (N_21033,N_20748,N_20645);
xor U21034 (N_21034,N_20643,N_20976);
or U21035 (N_21035,N_20553,N_20687);
xnor U21036 (N_21036,N_20533,N_20696);
xnor U21037 (N_21037,N_20588,N_20510);
xor U21038 (N_21038,N_20755,N_20530);
xnor U21039 (N_21039,N_20605,N_20938);
and U21040 (N_21040,N_20942,N_20823);
or U21041 (N_21041,N_20787,N_20767);
nor U21042 (N_21042,N_20916,N_20536);
or U21043 (N_21043,N_20814,N_20725);
or U21044 (N_21044,N_20933,N_20946);
and U21045 (N_21045,N_20807,N_20718);
and U21046 (N_21046,N_20932,N_20746);
and U21047 (N_21047,N_20988,N_20540);
nor U21048 (N_21048,N_20875,N_20637);
nand U21049 (N_21049,N_20603,N_20532);
xnor U21050 (N_21050,N_20611,N_20789);
and U21051 (N_21051,N_20728,N_20990);
and U21052 (N_21052,N_20769,N_20535);
xnor U21053 (N_21053,N_20766,N_20590);
nor U21054 (N_21054,N_20661,N_20992);
or U21055 (N_21055,N_20865,N_20838);
or U21056 (N_21056,N_20919,N_20613);
nand U21057 (N_21057,N_20862,N_20622);
nor U21058 (N_21058,N_20959,N_20597);
and U21059 (N_21059,N_20562,N_20798);
nand U21060 (N_21060,N_20945,N_20893);
nand U21061 (N_21061,N_20700,N_20595);
or U21062 (N_21062,N_20731,N_20981);
and U21063 (N_21063,N_20957,N_20881);
nand U21064 (N_21064,N_20503,N_20749);
or U21065 (N_21065,N_20628,N_20840);
or U21066 (N_21066,N_20950,N_20761);
nand U21067 (N_21067,N_20869,N_20774);
or U21068 (N_21068,N_20911,N_20776);
nor U21069 (N_21069,N_20778,N_20809);
nor U21070 (N_21070,N_20708,N_20918);
nor U21071 (N_21071,N_20683,N_20625);
nand U21072 (N_21072,N_20747,N_20501);
or U21073 (N_21073,N_20707,N_20519);
and U21074 (N_21074,N_20734,N_20513);
and U21075 (N_21075,N_20509,N_20592);
and U21076 (N_21076,N_20879,N_20529);
and U21077 (N_21077,N_20717,N_20786);
nand U21078 (N_21078,N_20819,N_20828);
nand U21079 (N_21079,N_20738,N_20854);
and U21080 (N_21080,N_20752,N_20905);
and U21081 (N_21081,N_20797,N_20967);
nand U21082 (N_21082,N_20754,N_20601);
and U21083 (N_21083,N_20805,N_20695);
and U21084 (N_21084,N_20985,N_20925);
nor U21085 (N_21085,N_20834,N_20745);
and U21086 (N_21086,N_20640,N_20975);
xnor U21087 (N_21087,N_20901,N_20500);
xnor U21088 (N_21088,N_20564,N_20937);
or U21089 (N_21089,N_20596,N_20554);
nor U21090 (N_21090,N_20829,N_20567);
and U21091 (N_21091,N_20599,N_20702);
or U21092 (N_21092,N_20785,N_20631);
or U21093 (N_21093,N_20593,N_20882);
nor U21094 (N_21094,N_20518,N_20545);
xnor U21095 (N_21095,N_20538,N_20960);
xnor U21096 (N_21096,N_20527,N_20861);
and U21097 (N_21097,N_20735,N_20896);
nor U21098 (N_21098,N_20656,N_20701);
nor U21099 (N_21099,N_20664,N_20779);
and U21100 (N_21100,N_20551,N_20955);
or U21101 (N_21101,N_20591,N_20550);
nand U21102 (N_21102,N_20575,N_20890);
and U21103 (N_21103,N_20569,N_20638);
nand U21104 (N_21104,N_20710,N_20803);
or U21105 (N_21105,N_20857,N_20703);
and U21106 (N_21106,N_20626,N_20934);
nand U21107 (N_21107,N_20511,N_20679);
nor U21108 (N_21108,N_20952,N_20733);
xnor U21109 (N_21109,N_20915,N_20777);
nand U21110 (N_21110,N_20516,N_20600);
nor U21111 (N_21111,N_20583,N_20741);
nand U21112 (N_21112,N_20773,N_20691);
nand U21113 (N_21113,N_20639,N_20855);
or U21114 (N_21114,N_20780,N_20760);
nand U21115 (N_21115,N_20993,N_20671);
or U21116 (N_21116,N_20682,N_20965);
and U21117 (N_21117,N_20624,N_20684);
and U21118 (N_21118,N_20506,N_20531);
nor U21119 (N_21119,N_20978,N_20817);
or U21120 (N_21120,N_20557,N_20806);
or U21121 (N_21121,N_20610,N_20581);
nor U21122 (N_21122,N_20598,N_20744);
nor U21123 (N_21123,N_20632,N_20943);
nand U21124 (N_21124,N_20563,N_20565);
nand U21125 (N_21125,N_20690,N_20722);
nand U21126 (N_21126,N_20589,N_20612);
and U21127 (N_21127,N_20989,N_20697);
xor U21128 (N_21128,N_20528,N_20693);
or U21129 (N_21129,N_20904,N_20826);
nor U21130 (N_21130,N_20566,N_20737);
and U21131 (N_21131,N_20572,N_20517);
nand U21132 (N_21132,N_20616,N_20968);
and U21133 (N_21133,N_20827,N_20860);
and U21134 (N_21134,N_20782,N_20921);
nand U21135 (N_21135,N_20852,N_20556);
xnor U21136 (N_21136,N_20729,N_20698);
nand U21137 (N_21137,N_20641,N_20524);
nand U21138 (N_21138,N_20765,N_20781);
xnor U21139 (N_21139,N_20820,N_20999);
and U21140 (N_21140,N_20512,N_20602);
or U21141 (N_21141,N_20587,N_20889);
xnor U21142 (N_21142,N_20832,N_20699);
and U21143 (N_21143,N_20654,N_20842);
xnor U21144 (N_21144,N_20724,N_20580);
and U21145 (N_21145,N_20913,N_20655);
or U21146 (N_21146,N_20615,N_20892);
and U21147 (N_21147,N_20848,N_20888);
nand U21148 (N_21148,N_20986,N_20674);
xor U21149 (N_21149,N_20977,N_20650);
or U21150 (N_21150,N_20931,N_20753);
xor U21151 (N_21151,N_20502,N_20652);
nor U21152 (N_21152,N_20594,N_20659);
xnor U21153 (N_21153,N_20973,N_20885);
and U21154 (N_21154,N_20830,N_20899);
xor U21155 (N_21155,N_20940,N_20505);
and U21156 (N_21156,N_20770,N_20740);
or U21157 (N_21157,N_20521,N_20979);
or U21158 (N_21158,N_20635,N_20983);
and U21159 (N_21159,N_20795,N_20850);
xor U21160 (N_21160,N_20548,N_20673);
nand U21161 (N_21161,N_20739,N_20623);
nor U21162 (N_21162,N_20876,N_20895);
and U21163 (N_21163,N_20792,N_20972);
xnor U21164 (N_21164,N_20742,N_20839);
xnor U21165 (N_21165,N_20974,N_20847);
nor U21166 (N_21166,N_20537,N_20676);
or U21167 (N_21167,N_20929,N_20873);
or U21168 (N_21168,N_20646,N_20508);
nor U21169 (N_21169,N_20574,N_20542);
nand U21170 (N_21170,N_20525,N_20845);
and U21171 (N_21171,N_20666,N_20607);
nor U21172 (N_21172,N_20948,N_20675);
nand U21173 (N_21173,N_20670,N_20606);
or U21174 (N_21174,N_20689,N_20757);
and U21175 (N_21175,N_20705,N_20835);
xor U21176 (N_21176,N_20947,N_20843);
xnor U21177 (N_21177,N_20677,N_20663);
nand U21178 (N_21178,N_20912,N_20570);
nor U21179 (N_21179,N_20799,N_20970);
xnor U21180 (N_21180,N_20681,N_20971);
nor U21181 (N_21181,N_20906,N_20836);
or U21182 (N_21182,N_20688,N_20526);
nand U21183 (N_21183,N_20692,N_20841);
xor U21184 (N_21184,N_20618,N_20507);
nor U21185 (N_21185,N_20863,N_20732);
nand U21186 (N_21186,N_20672,N_20808);
and U21187 (N_21187,N_20578,N_20815);
nor U21188 (N_21188,N_20520,N_20714);
nand U21189 (N_21189,N_20812,N_20608);
nand U21190 (N_21190,N_20964,N_20678);
or U21191 (N_21191,N_20796,N_20642);
or U21192 (N_21192,N_20558,N_20849);
xor U21193 (N_21193,N_20851,N_20930);
xor U21194 (N_21194,N_20867,N_20846);
nor U21195 (N_21195,N_20784,N_20910);
xor U21196 (N_21196,N_20764,N_20872);
xor U21197 (N_21197,N_20546,N_20887);
xnor U21198 (N_21198,N_20627,N_20772);
and U21199 (N_21199,N_20886,N_20914);
nand U21200 (N_21200,N_20922,N_20810);
or U21201 (N_21201,N_20941,N_20980);
nand U21202 (N_21202,N_20514,N_20920);
xnor U21203 (N_21203,N_20584,N_20620);
and U21204 (N_21204,N_20568,N_20825);
nand U21205 (N_21205,N_20903,N_20837);
nor U21206 (N_21206,N_20579,N_20868);
nor U21207 (N_21207,N_20571,N_20939);
xor U21208 (N_21208,N_20818,N_20582);
and U21209 (N_21209,N_20949,N_20660);
nor U21210 (N_21210,N_20924,N_20668);
nor U21211 (N_21211,N_20900,N_20726);
xnor U21212 (N_21212,N_20982,N_20647);
and U21213 (N_21213,N_20649,N_20736);
and U21214 (N_21214,N_20874,N_20927);
or U21215 (N_21215,N_20547,N_20864);
and U21216 (N_21216,N_20816,N_20877);
nor U21217 (N_21217,N_20515,N_20763);
and U21218 (N_21218,N_20667,N_20907);
xnor U21219 (N_21219,N_20751,N_20791);
nand U21220 (N_21220,N_20951,N_20923);
nand U21221 (N_21221,N_20750,N_20891);
and U21222 (N_21222,N_20651,N_20534);
and U21223 (N_21223,N_20648,N_20894);
nand U21224 (N_21224,N_20522,N_20928);
xor U21225 (N_21225,N_20555,N_20771);
or U21226 (N_21226,N_20576,N_20560);
and U21227 (N_21227,N_20813,N_20552);
and U21228 (N_21228,N_20559,N_20604);
nand U21229 (N_21229,N_20801,N_20523);
or U21230 (N_21230,N_20909,N_20543);
nand U21231 (N_21231,N_20727,N_20935);
and U21232 (N_21232,N_20883,N_20706);
nor U21233 (N_21233,N_20902,N_20586);
xor U21234 (N_21234,N_20768,N_20994);
or U21235 (N_21235,N_20783,N_20539);
nand U21236 (N_21236,N_20573,N_20629);
nor U21237 (N_21237,N_20917,N_20775);
or U21238 (N_21238,N_20716,N_20997);
xor U21239 (N_21239,N_20853,N_20998);
nor U21240 (N_21240,N_20609,N_20644);
nor U21241 (N_21241,N_20723,N_20996);
nand U21242 (N_21242,N_20858,N_20963);
xnor U21243 (N_21243,N_20721,N_20831);
nor U21244 (N_21244,N_20711,N_20794);
xnor U21245 (N_21245,N_20720,N_20962);
xor U21246 (N_21246,N_20793,N_20619);
nor U21247 (N_21247,N_20653,N_20630);
nand U21248 (N_21248,N_20758,N_20756);
or U21249 (N_21249,N_20636,N_20561);
or U21250 (N_21250,N_20522,N_20715);
nor U21251 (N_21251,N_20996,N_20622);
and U21252 (N_21252,N_20753,N_20792);
nand U21253 (N_21253,N_20504,N_20785);
nor U21254 (N_21254,N_20846,N_20616);
and U21255 (N_21255,N_20987,N_20744);
and U21256 (N_21256,N_20608,N_20766);
nand U21257 (N_21257,N_20887,N_20751);
or U21258 (N_21258,N_20760,N_20804);
xnor U21259 (N_21259,N_20649,N_20681);
nor U21260 (N_21260,N_20794,N_20831);
and U21261 (N_21261,N_20517,N_20522);
and U21262 (N_21262,N_20841,N_20584);
and U21263 (N_21263,N_20777,N_20771);
or U21264 (N_21264,N_20619,N_20902);
or U21265 (N_21265,N_20522,N_20796);
and U21266 (N_21266,N_20709,N_20759);
or U21267 (N_21267,N_20825,N_20579);
and U21268 (N_21268,N_20517,N_20636);
nor U21269 (N_21269,N_20570,N_20567);
or U21270 (N_21270,N_20636,N_20514);
xor U21271 (N_21271,N_20879,N_20695);
nor U21272 (N_21272,N_20677,N_20623);
nor U21273 (N_21273,N_20790,N_20530);
nor U21274 (N_21274,N_20735,N_20978);
nor U21275 (N_21275,N_20969,N_20821);
and U21276 (N_21276,N_20842,N_20611);
nand U21277 (N_21277,N_20798,N_20814);
xnor U21278 (N_21278,N_20853,N_20833);
nand U21279 (N_21279,N_20566,N_20653);
nand U21280 (N_21280,N_20576,N_20561);
nand U21281 (N_21281,N_20878,N_20602);
nand U21282 (N_21282,N_20684,N_20563);
xor U21283 (N_21283,N_20979,N_20593);
nor U21284 (N_21284,N_20839,N_20611);
xnor U21285 (N_21285,N_20790,N_20642);
nor U21286 (N_21286,N_20864,N_20865);
and U21287 (N_21287,N_20693,N_20633);
nand U21288 (N_21288,N_20863,N_20935);
nor U21289 (N_21289,N_20896,N_20804);
or U21290 (N_21290,N_20800,N_20661);
nor U21291 (N_21291,N_20691,N_20661);
nor U21292 (N_21292,N_20634,N_20674);
or U21293 (N_21293,N_20581,N_20604);
and U21294 (N_21294,N_20986,N_20805);
and U21295 (N_21295,N_20520,N_20747);
nor U21296 (N_21296,N_20851,N_20807);
nand U21297 (N_21297,N_20510,N_20764);
or U21298 (N_21298,N_20702,N_20846);
nand U21299 (N_21299,N_20742,N_20830);
or U21300 (N_21300,N_20544,N_20875);
nor U21301 (N_21301,N_20627,N_20795);
xor U21302 (N_21302,N_20887,N_20860);
nor U21303 (N_21303,N_20615,N_20906);
xor U21304 (N_21304,N_20757,N_20978);
nor U21305 (N_21305,N_20848,N_20626);
nand U21306 (N_21306,N_20807,N_20876);
nand U21307 (N_21307,N_20853,N_20842);
and U21308 (N_21308,N_20633,N_20838);
or U21309 (N_21309,N_20824,N_20858);
nand U21310 (N_21310,N_20798,N_20653);
and U21311 (N_21311,N_20815,N_20929);
or U21312 (N_21312,N_20635,N_20553);
nand U21313 (N_21313,N_20696,N_20881);
nor U21314 (N_21314,N_20602,N_20520);
nor U21315 (N_21315,N_20757,N_20967);
nor U21316 (N_21316,N_20885,N_20548);
nor U21317 (N_21317,N_20883,N_20620);
nor U21318 (N_21318,N_20737,N_20807);
or U21319 (N_21319,N_20913,N_20626);
nor U21320 (N_21320,N_20520,N_20766);
or U21321 (N_21321,N_20588,N_20770);
nor U21322 (N_21322,N_20776,N_20934);
nand U21323 (N_21323,N_20624,N_20530);
or U21324 (N_21324,N_20650,N_20916);
nand U21325 (N_21325,N_20698,N_20992);
xnor U21326 (N_21326,N_20694,N_20901);
nand U21327 (N_21327,N_20986,N_20821);
or U21328 (N_21328,N_20872,N_20913);
nor U21329 (N_21329,N_20738,N_20578);
nor U21330 (N_21330,N_20828,N_20734);
nor U21331 (N_21331,N_20793,N_20653);
and U21332 (N_21332,N_20660,N_20677);
and U21333 (N_21333,N_20550,N_20984);
nand U21334 (N_21334,N_20983,N_20750);
xor U21335 (N_21335,N_20540,N_20701);
nor U21336 (N_21336,N_20830,N_20883);
nand U21337 (N_21337,N_20801,N_20885);
nand U21338 (N_21338,N_20902,N_20735);
and U21339 (N_21339,N_20739,N_20793);
nor U21340 (N_21340,N_20877,N_20793);
nand U21341 (N_21341,N_20889,N_20842);
and U21342 (N_21342,N_20512,N_20707);
or U21343 (N_21343,N_20503,N_20744);
nor U21344 (N_21344,N_20687,N_20811);
nor U21345 (N_21345,N_20930,N_20546);
nand U21346 (N_21346,N_20629,N_20576);
xnor U21347 (N_21347,N_20985,N_20785);
nand U21348 (N_21348,N_20688,N_20947);
nor U21349 (N_21349,N_20666,N_20547);
or U21350 (N_21350,N_20762,N_20721);
and U21351 (N_21351,N_20779,N_20631);
nand U21352 (N_21352,N_20664,N_20704);
xor U21353 (N_21353,N_20771,N_20919);
nor U21354 (N_21354,N_20748,N_20540);
or U21355 (N_21355,N_20885,N_20977);
xnor U21356 (N_21356,N_20584,N_20703);
nor U21357 (N_21357,N_20668,N_20634);
nand U21358 (N_21358,N_20523,N_20808);
or U21359 (N_21359,N_20995,N_20967);
nand U21360 (N_21360,N_20727,N_20814);
nor U21361 (N_21361,N_20607,N_20606);
xor U21362 (N_21362,N_20701,N_20775);
nand U21363 (N_21363,N_20681,N_20868);
nand U21364 (N_21364,N_20986,N_20917);
nor U21365 (N_21365,N_20916,N_20586);
xor U21366 (N_21366,N_20572,N_20686);
nand U21367 (N_21367,N_20826,N_20531);
and U21368 (N_21368,N_20556,N_20953);
nand U21369 (N_21369,N_20786,N_20992);
xnor U21370 (N_21370,N_20651,N_20578);
or U21371 (N_21371,N_20698,N_20566);
xnor U21372 (N_21372,N_20793,N_20892);
xor U21373 (N_21373,N_20734,N_20559);
nor U21374 (N_21374,N_20544,N_20819);
nor U21375 (N_21375,N_20865,N_20981);
nor U21376 (N_21376,N_20761,N_20708);
nand U21377 (N_21377,N_20577,N_20873);
and U21378 (N_21378,N_20967,N_20606);
xnor U21379 (N_21379,N_20956,N_20540);
nor U21380 (N_21380,N_20790,N_20649);
nor U21381 (N_21381,N_20760,N_20899);
nand U21382 (N_21382,N_20617,N_20887);
nand U21383 (N_21383,N_20672,N_20528);
and U21384 (N_21384,N_20723,N_20565);
and U21385 (N_21385,N_20647,N_20995);
or U21386 (N_21386,N_20975,N_20657);
and U21387 (N_21387,N_20686,N_20564);
xor U21388 (N_21388,N_20642,N_20645);
xnor U21389 (N_21389,N_20893,N_20878);
xor U21390 (N_21390,N_20598,N_20784);
or U21391 (N_21391,N_20839,N_20595);
nand U21392 (N_21392,N_20921,N_20598);
and U21393 (N_21393,N_20547,N_20567);
nand U21394 (N_21394,N_20737,N_20688);
xor U21395 (N_21395,N_20731,N_20984);
nand U21396 (N_21396,N_20923,N_20586);
xor U21397 (N_21397,N_20768,N_20991);
or U21398 (N_21398,N_20900,N_20610);
nand U21399 (N_21399,N_20587,N_20695);
nand U21400 (N_21400,N_20894,N_20617);
xor U21401 (N_21401,N_20764,N_20793);
or U21402 (N_21402,N_20576,N_20714);
xnor U21403 (N_21403,N_20863,N_20605);
or U21404 (N_21404,N_20817,N_20556);
nor U21405 (N_21405,N_20915,N_20869);
and U21406 (N_21406,N_20615,N_20741);
xor U21407 (N_21407,N_20751,N_20584);
or U21408 (N_21408,N_20641,N_20698);
nand U21409 (N_21409,N_20943,N_20901);
nand U21410 (N_21410,N_20983,N_20825);
xnor U21411 (N_21411,N_20981,N_20685);
and U21412 (N_21412,N_20881,N_20673);
xnor U21413 (N_21413,N_20776,N_20953);
xnor U21414 (N_21414,N_20588,N_20918);
or U21415 (N_21415,N_20822,N_20691);
nand U21416 (N_21416,N_20754,N_20846);
xnor U21417 (N_21417,N_20644,N_20517);
xnor U21418 (N_21418,N_20692,N_20677);
nand U21419 (N_21419,N_20503,N_20641);
or U21420 (N_21420,N_20880,N_20521);
nor U21421 (N_21421,N_20549,N_20626);
or U21422 (N_21422,N_20603,N_20974);
nand U21423 (N_21423,N_20884,N_20518);
and U21424 (N_21424,N_20824,N_20748);
or U21425 (N_21425,N_20583,N_20662);
xnor U21426 (N_21426,N_20736,N_20575);
or U21427 (N_21427,N_20669,N_20985);
xnor U21428 (N_21428,N_20886,N_20665);
nor U21429 (N_21429,N_20636,N_20585);
nor U21430 (N_21430,N_20568,N_20910);
nand U21431 (N_21431,N_20723,N_20518);
nor U21432 (N_21432,N_20662,N_20923);
or U21433 (N_21433,N_20751,N_20803);
and U21434 (N_21434,N_20897,N_20809);
nor U21435 (N_21435,N_20781,N_20817);
or U21436 (N_21436,N_20796,N_20777);
or U21437 (N_21437,N_20523,N_20504);
or U21438 (N_21438,N_20909,N_20678);
or U21439 (N_21439,N_20816,N_20843);
and U21440 (N_21440,N_20695,N_20874);
or U21441 (N_21441,N_20843,N_20526);
or U21442 (N_21442,N_20764,N_20867);
nand U21443 (N_21443,N_20833,N_20934);
or U21444 (N_21444,N_20531,N_20761);
or U21445 (N_21445,N_20816,N_20824);
nand U21446 (N_21446,N_20830,N_20909);
or U21447 (N_21447,N_20566,N_20747);
nand U21448 (N_21448,N_20822,N_20640);
and U21449 (N_21449,N_20832,N_20996);
xor U21450 (N_21450,N_20799,N_20836);
nand U21451 (N_21451,N_20560,N_20563);
nand U21452 (N_21452,N_20673,N_20525);
and U21453 (N_21453,N_20719,N_20574);
xnor U21454 (N_21454,N_20951,N_20522);
and U21455 (N_21455,N_20655,N_20870);
or U21456 (N_21456,N_20613,N_20978);
nor U21457 (N_21457,N_20965,N_20638);
and U21458 (N_21458,N_20501,N_20507);
nand U21459 (N_21459,N_20875,N_20955);
nor U21460 (N_21460,N_20659,N_20682);
xor U21461 (N_21461,N_20911,N_20865);
or U21462 (N_21462,N_20560,N_20829);
nor U21463 (N_21463,N_20778,N_20568);
or U21464 (N_21464,N_20997,N_20982);
nor U21465 (N_21465,N_20532,N_20591);
xnor U21466 (N_21466,N_20764,N_20691);
nor U21467 (N_21467,N_20738,N_20938);
nor U21468 (N_21468,N_20756,N_20770);
xnor U21469 (N_21469,N_20821,N_20693);
or U21470 (N_21470,N_20988,N_20601);
xor U21471 (N_21471,N_20754,N_20713);
nor U21472 (N_21472,N_20664,N_20638);
nor U21473 (N_21473,N_20878,N_20792);
nor U21474 (N_21474,N_20888,N_20736);
nand U21475 (N_21475,N_20706,N_20768);
nand U21476 (N_21476,N_20799,N_20869);
and U21477 (N_21477,N_20957,N_20975);
or U21478 (N_21478,N_20546,N_20786);
nor U21479 (N_21479,N_20539,N_20747);
nor U21480 (N_21480,N_20776,N_20793);
nand U21481 (N_21481,N_20703,N_20506);
nand U21482 (N_21482,N_20809,N_20941);
or U21483 (N_21483,N_20712,N_20667);
xnor U21484 (N_21484,N_20800,N_20850);
or U21485 (N_21485,N_20515,N_20927);
xnor U21486 (N_21486,N_20937,N_20849);
nand U21487 (N_21487,N_20709,N_20746);
nand U21488 (N_21488,N_20831,N_20533);
xor U21489 (N_21489,N_20605,N_20736);
nand U21490 (N_21490,N_20639,N_20770);
and U21491 (N_21491,N_20937,N_20782);
and U21492 (N_21492,N_20958,N_20943);
xor U21493 (N_21493,N_20775,N_20515);
nand U21494 (N_21494,N_20835,N_20655);
nand U21495 (N_21495,N_20801,N_20925);
and U21496 (N_21496,N_20900,N_20860);
and U21497 (N_21497,N_20943,N_20674);
nor U21498 (N_21498,N_20779,N_20936);
nand U21499 (N_21499,N_20985,N_20637);
nor U21500 (N_21500,N_21371,N_21385);
nand U21501 (N_21501,N_21422,N_21022);
nand U21502 (N_21502,N_21414,N_21261);
and U21503 (N_21503,N_21127,N_21170);
xor U21504 (N_21504,N_21187,N_21193);
xor U21505 (N_21505,N_21000,N_21496);
and U21506 (N_21506,N_21205,N_21429);
or U21507 (N_21507,N_21292,N_21060);
and U21508 (N_21508,N_21472,N_21388);
xor U21509 (N_21509,N_21445,N_21207);
xnor U21510 (N_21510,N_21177,N_21419);
and U21511 (N_21511,N_21186,N_21120);
nor U21512 (N_21512,N_21399,N_21342);
and U21513 (N_21513,N_21267,N_21034);
or U21514 (N_21514,N_21158,N_21375);
xnor U21515 (N_21515,N_21173,N_21420);
nand U21516 (N_21516,N_21457,N_21286);
and U21517 (N_21517,N_21411,N_21454);
and U21518 (N_21518,N_21223,N_21161);
or U21519 (N_21519,N_21406,N_21288);
nand U21520 (N_21520,N_21356,N_21019);
nor U21521 (N_21521,N_21440,N_21243);
and U21522 (N_21522,N_21026,N_21255);
xor U21523 (N_21523,N_21183,N_21273);
nor U21524 (N_21524,N_21112,N_21113);
nand U21525 (N_21525,N_21485,N_21357);
nor U21526 (N_21526,N_21217,N_21297);
and U21527 (N_21527,N_21259,N_21095);
nand U21528 (N_21528,N_21413,N_21084);
nand U21529 (N_21529,N_21171,N_21244);
and U21530 (N_21530,N_21129,N_21133);
nand U21531 (N_21531,N_21262,N_21444);
nor U21532 (N_21532,N_21470,N_21097);
nor U21533 (N_21533,N_21073,N_21070);
nor U21534 (N_21534,N_21009,N_21322);
or U21535 (N_21535,N_21248,N_21380);
nand U21536 (N_21536,N_21085,N_21269);
nor U21537 (N_21537,N_21241,N_21032);
nand U21538 (N_21538,N_21037,N_21374);
and U21539 (N_21539,N_21305,N_21423);
xnor U21540 (N_21540,N_21099,N_21151);
and U21541 (N_21541,N_21434,N_21090);
and U21542 (N_21542,N_21483,N_21266);
nand U21543 (N_21543,N_21361,N_21105);
nor U21544 (N_21544,N_21108,N_21296);
nor U21545 (N_21545,N_21174,N_21114);
and U21546 (N_21546,N_21426,N_21004);
xnor U21547 (N_21547,N_21005,N_21447);
and U21548 (N_21548,N_21030,N_21017);
nor U21549 (N_21549,N_21013,N_21199);
and U21550 (N_21550,N_21143,N_21192);
or U21551 (N_21551,N_21263,N_21020);
or U21552 (N_21552,N_21140,N_21359);
nor U21553 (N_21553,N_21314,N_21442);
nor U21554 (N_21554,N_21221,N_21206);
xnor U21555 (N_21555,N_21274,N_21281);
xor U21556 (N_21556,N_21278,N_21401);
or U21557 (N_21557,N_21150,N_21325);
and U21558 (N_21558,N_21135,N_21093);
xor U21559 (N_21559,N_21308,N_21283);
xnor U21560 (N_21560,N_21246,N_21456);
nor U21561 (N_21561,N_21260,N_21110);
and U21562 (N_21562,N_21366,N_21229);
nand U21563 (N_21563,N_21491,N_21404);
nor U21564 (N_21564,N_21169,N_21332);
nand U21565 (N_21565,N_21088,N_21236);
and U21566 (N_21566,N_21346,N_21331);
xnor U21567 (N_21567,N_21036,N_21389);
nand U21568 (N_21568,N_21294,N_21204);
and U21569 (N_21569,N_21301,N_21490);
nor U21570 (N_21570,N_21035,N_21293);
xor U21571 (N_21571,N_21191,N_21068);
nand U21572 (N_21572,N_21144,N_21363);
nand U21573 (N_21573,N_21042,N_21317);
or U21574 (N_21574,N_21486,N_21280);
xor U21575 (N_21575,N_21272,N_21249);
nand U21576 (N_21576,N_21157,N_21118);
nand U21577 (N_21577,N_21290,N_21250);
or U21578 (N_21578,N_21117,N_21195);
nand U21579 (N_21579,N_21153,N_21450);
and U21580 (N_21580,N_21251,N_21387);
or U21581 (N_21581,N_21458,N_21462);
xor U21582 (N_21582,N_21446,N_21024);
and U21583 (N_21583,N_21130,N_21386);
nand U21584 (N_21584,N_21393,N_21175);
nand U21585 (N_21585,N_21015,N_21460);
or U21586 (N_21586,N_21010,N_21298);
and U21587 (N_21587,N_21333,N_21126);
and U21588 (N_21588,N_21424,N_21040);
and U21589 (N_21589,N_21482,N_21327);
xnor U21590 (N_21590,N_21358,N_21023);
or U21591 (N_21591,N_21289,N_21355);
or U21592 (N_21592,N_21448,N_21370);
xnor U21593 (N_21593,N_21237,N_21421);
and U21594 (N_21594,N_21218,N_21319);
nor U21595 (N_21595,N_21159,N_21451);
nand U21596 (N_21596,N_21392,N_21210);
xnor U21597 (N_21597,N_21466,N_21307);
nor U21598 (N_21598,N_21369,N_21344);
or U21599 (N_21599,N_21107,N_21235);
or U21600 (N_21600,N_21148,N_21196);
and U21601 (N_21601,N_21328,N_21043);
nor U21602 (N_21602,N_21203,N_21412);
nor U21603 (N_21603,N_21306,N_21165);
nand U21604 (N_21604,N_21116,N_21007);
xnor U21605 (N_21605,N_21123,N_21271);
nand U21606 (N_21606,N_21390,N_21141);
or U21607 (N_21607,N_21285,N_21189);
nor U21608 (N_21608,N_21179,N_21057);
nor U21609 (N_21609,N_21227,N_21498);
or U21610 (N_21610,N_21417,N_21018);
xnor U21611 (N_21611,N_21052,N_21152);
xnor U21612 (N_21612,N_21372,N_21348);
nand U21613 (N_21613,N_21418,N_21475);
xor U21614 (N_21614,N_21452,N_21086);
nand U21615 (N_21615,N_21339,N_21435);
nor U21616 (N_21616,N_21198,N_21051);
nor U21617 (N_21617,N_21131,N_21106);
nor U21618 (N_21618,N_21038,N_21295);
and U21619 (N_21619,N_21211,N_21087);
xor U21620 (N_21620,N_21337,N_21321);
xor U21621 (N_21621,N_21316,N_21416);
xnor U21622 (N_21622,N_21471,N_21438);
and U21623 (N_21623,N_21465,N_21076);
and U21624 (N_21624,N_21025,N_21313);
or U21625 (N_21625,N_21050,N_21493);
nand U21626 (N_21626,N_21326,N_21138);
nand U21627 (N_21627,N_21487,N_21125);
or U21628 (N_21628,N_21323,N_21265);
nor U21629 (N_21629,N_21154,N_21252);
xnor U21630 (N_21630,N_21464,N_21242);
and U21631 (N_21631,N_21232,N_21098);
or U21632 (N_21632,N_21433,N_21247);
and U21633 (N_21633,N_21058,N_21200);
nor U21634 (N_21634,N_21184,N_21484);
nand U21635 (N_21635,N_21489,N_21257);
and U21636 (N_21636,N_21347,N_21164);
and U21637 (N_21637,N_21228,N_21334);
or U21638 (N_21638,N_21176,N_21432);
and U21639 (N_21639,N_21335,N_21402);
or U21640 (N_21640,N_21391,N_21224);
nand U21641 (N_21641,N_21343,N_21100);
and U21642 (N_21642,N_21282,N_21081);
nand U21643 (N_21643,N_21029,N_21047);
nand U21644 (N_21644,N_21353,N_21378);
nor U21645 (N_21645,N_21222,N_21104);
or U21646 (N_21646,N_21202,N_21006);
nand U21647 (N_21647,N_21279,N_21453);
nor U21648 (N_21648,N_21270,N_21082);
and U21649 (N_21649,N_21056,N_21364);
nand U21650 (N_21650,N_21400,N_21080);
or U21651 (N_21651,N_21463,N_21049);
nand U21652 (N_21652,N_21373,N_21039);
nor U21653 (N_21653,N_21459,N_21311);
or U21654 (N_21654,N_21268,N_21415);
and U21655 (N_21655,N_21077,N_21044);
and U21656 (N_21656,N_21329,N_21155);
and U21657 (N_21657,N_21059,N_21405);
xnor U21658 (N_21658,N_21194,N_21443);
or U21659 (N_21659,N_21276,N_21383);
and U21660 (N_21660,N_21209,N_21368);
nor U21661 (N_21661,N_21254,N_21499);
and U21662 (N_21662,N_21461,N_21075);
or U21663 (N_21663,N_21381,N_21336);
xnor U21664 (N_21664,N_21479,N_21065);
nor U21665 (N_21665,N_21469,N_21309);
nor U21666 (N_21666,N_21384,N_21299);
xnor U21667 (N_21667,N_21287,N_21441);
and U21668 (N_21668,N_21312,N_21437);
and U21669 (N_21669,N_21233,N_21310);
and U21670 (N_21670,N_21041,N_21045);
nand U21671 (N_21671,N_21178,N_21338);
and U21672 (N_21672,N_21122,N_21008);
xnor U21673 (N_21673,N_21340,N_21215);
nand U21674 (N_21674,N_21407,N_21102);
or U21675 (N_21675,N_21495,N_21397);
and U21676 (N_21676,N_21324,N_21089);
xor U21677 (N_21677,N_21230,N_21197);
nand U21678 (N_21678,N_21330,N_21396);
nand U21679 (N_21679,N_21468,N_21239);
or U21680 (N_21680,N_21185,N_21003);
and U21681 (N_21681,N_21258,N_21220);
or U21682 (N_21682,N_21376,N_21067);
nand U21683 (N_21683,N_21403,N_21436);
xor U21684 (N_21684,N_21149,N_21395);
or U21685 (N_21685,N_21053,N_21014);
xor U21686 (N_21686,N_21360,N_21379);
or U21687 (N_21687,N_21101,N_21142);
or U21688 (N_21688,N_21264,N_21069);
nor U21689 (N_21689,N_21480,N_21428);
xnor U21690 (N_21690,N_21021,N_21449);
nor U21691 (N_21691,N_21066,N_21011);
and U21692 (N_21692,N_21354,N_21048);
nand U21693 (N_21693,N_21409,N_21061);
or U21694 (N_21694,N_21190,N_21352);
and U21695 (N_21695,N_21304,N_21094);
or U21696 (N_21696,N_21002,N_21033);
and U21697 (N_21697,N_21079,N_21072);
or U21698 (N_21698,N_21168,N_21341);
or U21699 (N_21699,N_21430,N_21427);
nor U21700 (N_21700,N_21062,N_21046);
nor U21701 (N_21701,N_21109,N_21147);
and U21702 (N_21702,N_21439,N_21367);
and U21703 (N_21703,N_21055,N_21492);
or U21704 (N_21704,N_21139,N_21284);
nor U21705 (N_21705,N_21172,N_21181);
or U21706 (N_21706,N_21477,N_21163);
and U21707 (N_21707,N_21398,N_21166);
nand U21708 (N_21708,N_21216,N_21382);
and U21709 (N_21709,N_21115,N_21256);
nand U21710 (N_21710,N_21027,N_21137);
or U21711 (N_21711,N_21128,N_21145);
nand U21712 (N_21712,N_21134,N_21208);
xor U21713 (N_21713,N_21488,N_21124);
and U21714 (N_21714,N_21291,N_21160);
or U21715 (N_21715,N_21362,N_21225);
nor U21716 (N_21716,N_21071,N_21119);
xnor U21717 (N_21717,N_21253,N_21240);
or U21718 (N_21718,N_21394,N_21092);
xnor U21719 (N_21719,N_21467,N_21078);
and U21720 (N_21720,N_21377,N_21365);
or U21721 (N_21721,N_21234,N_21146);
nand U21722 (N_21722,N_21303,N_21016);
or U21723 (N_21723,N_21156,N_21074);
nor U21724 (N_21724,N_21182,N_21238);
or U21725 (N_21725,N_21180,N_21214);
nor U21726 (N_21726,N_21497,N_21064);
or U21727 (N_21727,N_21231,N_21121);
nand U21728 (N_21728,N_21226,N_21001);
or U21729 (N_21729,N_21212,N_21474);
nand U21730 (N_21730,N_21476,N_21315);
nand U21731 (N_21731,N_21012,N_21083);
xor U21732 (N_21732,N_21103,N_21201);
or U21733 (N_21733,N_21219,N_21028);
xor U21734 (N_21734,N_21431,N_21345);
and U21735 (N_21735,N_21478,N_21245);
xor U21736 (N_21736,N_21320,N_21318);
and U21737 (N_21737,N_21350,N_21091);
xor U21738 (N_21738,N_21494,N_21136);
and U21739 (N_21739,N_21213,N_21277);
and U21740 (N_21740,N_21408,N_21351);
or U21741 (N_21741,N_21054,N_21167);
and U21742 (N_21742,N_21455,N_21425);
xor U21743 (N_21743,N_21481,N_21132);
nand U21744 (N_21744,N_21162,N_21410);
and U21745 (N_21745,N_21473,N_21300);
xor U21746 (N_21746,N_21349,N_21188);
nor U21747 (N_21747,N_21302,N_21096);
or U21748 (N_21748,N_21111,N_21063);
nand U21749 (N_21749,N_21031,N_21275);
nor U21750 (N_21750,N_21273,N_21349);
xnor U21751 (N_21751,N_21176,N_21067);
xnor U21752 (N_21752,N_21381,N_21144);
nand U21753 (N_21753,N_21481,N_21316);
xor U21754 (N_21754,N_21155,N_21473);
or U21755 (N_21755,N_21434,N_21234);
or U21756 (N_21756,N_21479,N_21478);
xor U21757 (N_21757,N_21119,N_21127);
nor U21758 (N_21758,N_21138,N_21144);
or U21759 (N_21759,N_21495,N_21177);
and U21760 (N_21760,N_21281,N_21324);
and U21761 (N_21761,N_21000,N_21495);
and U21762 (N_21762,N_21421,N_21263);
nand U21763 (N_21763,N_21404,N_21363);
and U21764 (N_21764,N_21391,N_21242);
nand U21765 (N_21765,N_21038,N_21196);
nor U21766 (N_21766,N_21465,N_21228);
or U21767 (N_21767,N_21181,N_21012);
and U21768 (N_21768,N_21114,N_21035);
xnor U21769 (N_21769,N_21232,N_21161);
xor U21770 (N_21770,N_21461,N_21118);
nand U21771 (N_21771,N_21194,N_21245);
and U21772 (N_21772,N_21470,N_21174);
xor U21773 (N_21773,N_21403,N_21272);
and U21774 (N_21774,N_21387,N_21369);
and U21775 (N_21775,N_21199,N_21258);
nand U21776 (N_21776,N_21299,N_21006);
xor U21777 (N_21777,N_21336,N_21143);
xor U21778 (N_21778,N_21276,N_21317);
nor U21779 (N_21779,N_21490,N_21031);
xor U21780 (N_21780,N_21312,N_21145);
and U21781 (N_21781,N_21405,N_21452);
nand U21782 (N_21782,N_21497,N_21211);
and U21783 (N_21783,N_21494,N_21083);
xnor U21784 (N_21784,N_21173,N_21016);
nand U21785 (N_21785,N_21328,N_21004);
or U21786 (N_21786,N_21109,N_21395);
or U21787 (N_21787,N_21228,N_21338);
xnor U21788 (N_21788,N_21378,N_21020);
nor U21789 (N_21789,N_21390,N_21217);
or U21790 (N_21790,N_21489,N_21120);
or U21791 (N_21791,N_21266,N_21042);
nor U21792 (N_21792,N_21380,N_21162);
or U21793 (N_21793,N_21209,N_21347);
xor U21794 (N_21794,N_21191,N_21344);
nor U21795 (N_21795,N_21116,N_21295);
nand U21796 (N_21796,N_21240,N_21156);
nand U21797 (N_21797,N_21363,N_21154);
xor U21798 (N_21798,N_21328,N_21230);
or U21799 (N_21799,N_21127,N_21035);
and U21800 (N_21800,N_21494,N_21058);
and U21801 (N_21801,N_21342,N_21008);
nand U21802 (N_21802,N_21441,N_21195);
nor U21803 (N_21803,N_21084,N_21453);
and U21804 (N_21804,N_21087,N_21075);
xnor U21805 (N_21805,N_21133,N_21319);
and U21806 (N_21806,N_21452,N_21138);
and U21807 (N_21807,N_21102,N_21307);
and U21808 (N_21808,N_21245,N_21451);
nor U21809 (N_21809,N_21381,N_21345);
nor U21810 (N_21810,N_21122,N_21223);
and U21811 (N_21811,N_21315,N_21010);
nor U21812 (N_21812,N_21340,N_21192);
nand U21813 (N_21813,N_21277,N_21256);
xnor U21814 (N_21814,N_21455,N_21458);
and U21815 (N_21815,N_21424,N_21116);
xor U21816 (N_21816,N_21349,N_21112);
nand U21817 (N_21817,N_21354,N_21197);
nand U21818 (N_21818,N_21383,N_21465);
and U21819 (N_21819,N_21139,N_21410);
nand U21820 (N_21820,N_21163,N_21468);
nor U21821 (N_21821,N_21133,N_21483);
xor U21822 (N_21822,N_21335,N_21147);
and U21823 (N_21823,N_21274,N_21126);
or U21824 (N_21824,N_21434,N_21174);
and U21825 (N_21825,N_21306,N_21396);
xor U21826 (N_21826,N_21423,N_21428);
or U21827 (N_21827,N_21175,N_21053);
nand U21828 (N_21828,N_21355,N_21215);
nand U21829 (N_21829,N_21082,N_21355);
or U21830 (N_21830,N_21307,N_21291);
nor U21831 (N_21831,N_21149,N_21283);
nor U21832 (N_21832,N_21217,N_21089);
or U21833 (N_21833,N_21122,N_21004);
or U21834 (N_21834,N_21088,N_21095);
nor U21835 (N_21835,N_21264,N_21048);
and U21836 (N_21836,N_21323,N_21345);
nor U21837 (N_21837,N_21473,N_21232);
nor U21838 (N_21838,N_21297,N_21396);
nor U21839 (N_21839,N_21172,N_21195);
or U21840 (N_21840,N_21158,N_21439);
or U21841 (N_21841,N_21182,N_21065);
nand U21842 (N_21842,N_21303,N_21424);
or U21843 (N_21843,N_21473,N_21471);
nand U21844 (N_21844,N_21050,N_21304);
xor U21845 (N_21845,N_21163,N_21316);
or U21846 (N_21846,N_21428,N_21055);
nand U21847 (N_21847,N_21023,N_21255);
nor U21848 (N_21848,N_21166,N_21190);
or U21849 (N_21849,N_21200,N_21395);
or U21850 (N_21850,N_21273,N_21326);
or U21851 (N_21851,N_21142,N_21280);
or U21852 (N_21852,N_21150,N_21393);
and U21853 (N_21853,N_21034,N_21217);
and U21854 (N_21854,N_21150,N_21379);
nor U21855 (N_21855,N_21085,N_21147);
or U21856 (N_21856,N_21301,N_21259);
and U21857 (N_21857,N_21114,N_21455);
xnor U21858 (N_21858,N_21418,N_21430);
or U21859 (N_21859,N_21336,N_21356);
xnor U21860 (N_21860,N_21182,N_21225);
nand U21861 (N_21861,N_21444,N_21126);
nand U21862 (N_21862,N_21330,N_21107);
nor U21863 (N_21863,N_21131,N_21349);
nand U21864 (N_21864,N_21360,N_21399);
nor U21865 (N_21865,N_21248,N_21249);
nor U21866 (N_21866,N_21148,N_21296);
nand U21867 (N_21867,N_21203,N_21268);
xor U21868 (N_21868,N_21464,N_21041);
nor U21869 (N_21869,N_21336,N_21032);
xnor U21870 (N_21870,N_21423,N_21352);
nor U21871 (N_21871,N_21149,N_21270);
nor U21872 (N_21872,N_21139,N_21187);
nand U21873 (N_21873,N_21277,N_21403);
and U21874 (N_21874,N_21429,N_21202);
nand U21875 (N_21875,N_21354,N_21043);
xor U21876 (N_21876,N_21081,N_21280);
and U21877 (N_21877,N_21430,N_21013);
or U21878 (N_21878,N_21117,N_21247);
and U21879 (N_21879,N_21095,N_21372);
xnor U21880 (N_21880,N_21236,N_21023);
xnor U21881 (N_21881,N_21078,N_21110);
nor U21882 (N_21882,N_21425,N_21364);
nor U21883 (N_21883,N_21009,N_21020);
nor U21884 (N_21884,N_21042,N_21491);
xor U21885 (N_21885,N_21123,N_21178);
nor U21886 (N_21886,N_21159,N_21070);
nor U21887 (N_21887,N_21136,N_21188);
or U21888 (N_21888,N_21441,N_21265);
nand U21889 (N_21889,N_21098,N_21178);
and U21890 (N_21890,N_21336,N_21017);
and U21891 (N_21891,N_21322,N_21256);
and U21892 (N_21892,N_21021,N_21447);
nand U21893 (N_21893,N_21373,N_21293);
or U21894 (N_21894,N_21454,N_21017);
xnor U21895 (N_21895,N_21339,N_21325);
or U21896 (N_21896,N_21301,N_21351);
and U21897 (N_21897,N_21000,N_21240);
and U21898 (N_21898,N_21007,N_21194);
and U21899 (N_21899,N_21047,N_21248);
xnor U21900 (N_21900,N_21315,N_21160);
and U21901 (N_21901,N_21060,N_21474);
or U21902 (N_21902,N_21422,N_21083);
or U21903 (N_21903,N_21075,N_21212);
nand U21904 (N_21904,N_21205,N_21356);
nand U21905 (N_21905,N_21254,N_21453);
or U21906 (N_21906,N_21225,N_21019);
and U21907 (N_21907,N_21061,N_21045);
and U21908 (N_21908,N_21191,N_21379);
nand U21909 (N_21909,N_21027,N_21133);
xor U21910 (N_21910,N_21074,N_21344);
and U21911 (N_21911,N_21220,N_21361);
and U21912 (N_21912,N_21472,N_21020);
and U21913 (N_21913,N_21184,N_21013);
or U21914 (N_21914,N_21132,N_21311);
nand U21915 (N_21915,N_21054,N_21264);
xor U21916 (N_21916,N_21057,N_21497);
nor U21917 (N_21917,N_21012,N_21431);
nor U21918 (N_21918,N_21194,N_21423);
xnor U21919 (N_21919,N_21323,N_21393);
nor U21920 (N_21920,N_21359,N_21038);
nor U21921 (N_21921,N_21060,N_21104);
nor U21922 (N_21922,N_21149,N_21207);
or U21923 (N_21923,N_21109,N_21131);
nand U21924 (N_21924,N_21363,N_21014);
and U21925 (N_21925,N_21114,N_21269);
nand U21926 (N_21926,N_21497,N_21069);
or U21927 (N_21927,N_21222,N_21354);
nor U21928 (N_21928,N_21096,N_21499);
or U21929 (N_21929,N_21092,N_21380);
and U21930 (N_21930,N_21480,N_21348);
or U21931 (N_21931,N_21323,N_21254);
nand U21932 (N_21932,N_21303,N_21450);
or U21933 (N_21933,N_21222,N_21264);
nand U21934 (N_21934,N_21479,N_21162);
xnor U21935 (N_21935,N_21227,N_21130);
nor U21936 (N_21936,N_21197,N_21065);
xnor U21937 (N_21937,N_21192,N_21141);
xor U21938 (N_21938,N_21141,N_21253);
xnor U21939 (N_21939,N_21210,N_21493);
nand U21940 (N_21940,N_21028,N_21482);
nand U21941 (N_21941,N_21154,N_21068);
or U21942 (N_21942,N_21388,N_21477);
xnor U21943 (N_21943,N_21113,N_21202);
xor U21944 (N_21944,N_21123,N_21154);
nor U21945 (N_21945,N_21355,N_21280);
nor U21946 (N_21946,N_21131,N_21450);
nor U21947 (N_21947,N_21062,N_21316);
xnor U21948 (N_21948,N_21238,N_21191);
xnor U21949 (N_21949,N_21048,N_21380);
and U21950 (N_21950,N_21374,N_21290);
nand U21951 (N_21951,N_21179,N_21134);
xor U21952 (N_21952,N_21403,N_21286);
and U21953 (N_21953,N_21057,N_21447);
xor U21954 (N_21954,N_21376,N_21410);
or U21955 (N_21955,N_21301,N_21229);
nor U21956 (N_21956,N_21285,N_21192);
or U21957 (N_21957,N_21212,N_21229);
or U21958 (N_21958,N_21340,N_21082);
xnor U21959 (N_21959,N_21185,N_21066);
xnor U21960 (N_21960,N_21316,N_21494);
nand U21961 (N_21961,N_21349,N_21343);
or U21962 (N_21962,N_21456,N_21413);
or U21963 (N_21963,N_21043,N_21059);
nor U21964 (N_21964,N_21334,N_21337);
nor U21965 (N_21965,N_21153,N_21234);
nand U21966 (N_21966,N_21024,N_21470);
nand U21967 (N_21967,N_21123,N_21284);
or U21968 (N_21968,N_21005,N_21425);
nand U21969 (N_21969,N_21028,N_21374);
xnor U21970 (N_21970,N_21099,N_21265);
nand U21971 (N_21971,N_21306,N_21214);
nor U21972 (N_21972,N_21440,N_21025);
or U21973 (N_21973,N_21327,N_21096);
xor U21974 (N_21974,N_21054,N_21410);
xnor U21975 (N_21975,N_21033,N_21428);
nor U21976 (N_21976,N_21247,N_21226);
nand U21977 (N_21977,N_21119,N_21146);
nand U21978 (N_21978,N_21302,N_21274);
nand U21979 (N_21979,N_21044,N_21147);
nor U21980 (N_21980,N_21339,N_21385);
nor U21981 (N_21981,N_21254,N_21199);
nand U21982 (N_21982,N_21003,N_21415);
nand U21983 (N_21983,N_21173,N_21066);
and U21984 (N_21984,N_21489,N_21161);
and U21985 (N_21985,N_21250,N_21177);
or U21986 (N_21986,N_21381,N_21224);
nand U21987 (N_21987,N_21457,N_21039);
nand U21988 (N_21988,N_21128,N_21151);
nand U21989 (N_21989,N_21368,N_21194);
nor U21990 (N_21990,N_21280,N_21430);
xnor U21991 (N_21991,N_21151,N_21176);
and U21992 (N_21992,N_21150,N_21491);
xnor U21993 (N_21993,N_21031,N_21394);
or U21994 (N_21994,N_21138,N_21180);
nor U21995 (N_21995,N_21025,N_21028);
xnor U21996 (N_21996,N_21100,N_21264);
nand U21997 (N_21997,N_21404,N_21300);
xnor U21998 (N_21998,N_21111,N_21191);
nand U21999 (N_21999,N_21168,N_21083);
xnor U22000 (N_22000,N_21779,N_21850);
and U22001 (N_22001,N_21794,N_21560);
and U22002 (N_22002,N_21562,N_21934);
or U22003 (N_22003,N_21645,N_21936);
and U22004 (N_22004,N_21993,N_21734);
nand U22005 (N_22005,N_21582,N_21827);
nand U22006 (N_22006,N_21762,N_21655);
and U22007 (N_22007,N_21553,N_21887);
or U22008 (N_22008,N_21835,N_21757);
xor U22009 (N_22009,N_21596,N_21960);
nor U22010 (N_22010,N_21601,N_21569);
and U22011 (N_22011,N_21909,N_21962);
and U22012 (N_22012,N_21573,N_21531);
and U22013 (N_22013,N_21978,N_21901);
or U22014 (N_22014,N_21672,N_21768);
nand U22015 (N_22015,N_21629,N_21654);
or U22016 (N_22016,N_21867,N_21931);
or U22017 (N_22017,N_21711,N_21519);
nor U22018 (N_22018,N_21876,N_21520);
and U22019 (N_22019,N_21988,N_21849);
nor U22020 (N_22020,N_21802,N_21597);
and U22021 (N_22021,N_21783,N_21566);
xor U22022 (N_22022,N_21511,N_21740);
or U22023 (N_22023,N_21682,N_21798);
nor U22024 (N_22024,N_21590,N_21907);
nor U22025 (N_22025,N_21980,N_21823);
and U22026 (N_22026,N_21615,N_21815);
xor U22027 (N_22027,N_21795,N_21700);
nand U22028 (N_22028,N_21610,N_21633);
and U22029 (N_22029,N_21838,N_21879);
or U22030 (N_22030,N_21656,N_21526);
and U22031 (N_22031,N_21780,N_21922);
nand U22032 (N_22032,N_21990,N_21657);
or U22033 (N_22033,N_21944,N_21549);
and U22034 (N_22034,N_21584,N_21819);
or U22035 (N_22035,N_21517,N_21735);
nor U22036 (N_22036,N_21646,N_21681);
and U22037 (N_22037,N_21644,N_21697);
nor U22038 (N_22038,N_21586,N_21699);
xnor U22039 (N_22039,N_21811,N_21774);
or U22040 (N_22040,N_21958,N_21955);
or U22041 (N_22041,N_21604,N_21754);
nor U22042 (N_22042,N_21982,N_21667);
xnor U22043 (N_22043,N_21996,N_21773);
and U22044 (N_22044,N_21576,N_21911);
or U22045 (N_22045,N_21719,N_21684);
nor U22046 (N_22046,N_21857,N_21525);
or U22047 (N_22047,N_21824,N_21809);
and U22048 (N_22048,N_21914,N_21659);
nor U22049 (N_22049,N_21686,N_21833);
or U22050 (N_22050,N_21895,N_21640);
nor U22051 (N_22051,N_21737,N_21885);
xor U22052 (N_22052,N_21705,N_21888);
nand U22053 (N_22053,N_21613,N_21623);
xor U22054 (N_22054,N_21583,N_21509);
and U22055 (N_22055,N_21539,N_21588);
nor U22056 (N_22056,N_21552,N_21891);
and U22057 (N_22057,N_21889,N_21653);
or U22058 (N_22058,N_21540,N_21598);
nand U22059 (N_22059,N_21919,N_21508);
and U22060 (N_22060,N_21935,N_21607);
or U22061 (N_22061,N_21899,N_21712);
xnor U22062 (N_22062,N_21845,N_21600);
or U22063 (N_22063,N_21842,N_21761);
and U22064 (N_22064,N_21991,N_21858);
nand U22065 (N_22065,N_21926,N_21832);
nand U22066 (N_22066,N_21679,N_21816);
or U22067 (N_22067,N_21637,N_21687);
or U22068 (N_22068,N_21942,N_21805);
nor U22069 (N_22069,N_21894,N_21591);
or U22070 (N_22070,N_21649,N_21866);
or U22071 (N_22071,N_21770,N_21671);
xor U22072 (N_22072,N_21886,N_21956);
nor U22073 (N_22073,N_21605,N_21967);
nand U22074 (N_22074,N_21963,N_21568);
nor U22075 (N_22075,N_21674,N_21543);
xor U22076 (N_22076,N_21846,N_21871);
nor U22077 (N_22077,N_21718,N_21972);
xor U22078 (N_22078,N_21592,N_21670);
nand U22079 (N_22079,N_21860,N_21567);
xor U22080 (N_22080,N_21621,N_21826);
nor U22081 (N_22081,N_21878,N_21751);
or U22082 (N_22082,N_21548,N_21853);
xnor U22083 (N_22083,N_21542,N_21665);
nand U22084 (N_22084,N_21896,N_21714);
xor U22085 (N_22085,N_21707,N_21863);
xnor U22086 (N_22086,N_21717,N_21787);
nor U22087 (N_22087,N_21785,N_21913);
nor U22088 (N_22088,N_21854,N_21694);
and U22089 (N_22089,N_21973,N_21500);
and U22090 (N_22090,N_21589,N_21766);
nand U22091 (N_22091,N_21535,N_21627);
nor U22092 (N_22092,N_21759,N_21528);
nand U22093 (N_22093,N_21504,N_21620);
and U22094 (N_22094,N_21917,N_21673);
and U22095 (N_22095,N_21954,N_21651);
or U22096 (N_22096,N_21938,N_21829);
nand U22097 (N_22097,N_21695,N_21728);
nand U22098 (N_22098,N_21581,N_21533);
nand U22099 (N_22099,N_21945,N_21564);
nand U22100 (N_22100,N_21666,N_21578);
nor U22101 (N_22101,N_21663,N_21703);
and U22102 (N_22102,N_21870,N_21776);
nor U22103 (N_22103,N_21769,N_21534);
or U22104 (N_22104,N_21808,N_21698);
nor U22105 (N_22105,N_21696,N_21987);
or U22106 (N_22106,N_21953,N_21940);
or U22107 (N_22107,N_21947,N_21507);
xnor U22108 (N_22108,N_21822,N_21561);
xnor U22109 (N_22109,N_21538,N_21618);
xor U22110 (N_22110,N_21632,N_21593);
or U22111 (N_22111,N_21585,N_21726);
and U22112 (N_22112,N_21710,N_21505);
nor U22113 (N_22113,N_21855,N_21658);
nor U22114 (N_22114,N_21792,N_21516);
nor U22115 (N_22115,N_21580,N_21760);
and U22116 (N_22116,N_21976,N_21579);
xnor U22117 (N_22117,N_21675,N_21959);
or U22118 (N_22118,N_21908,N_21738);
xor U22119 (N_22119,N_21558,N_21898);
and U22120 (N_22120,N_21796,N_21523);
xnor U22121 (N_22121,N_21716,N_21994);
xor U22122 (N_22122,N_21702,N_21793);
xnor U22123 (N_22123,N_21557,N_21704);
nand U22124 (N_22124,N_21890,N_21676);
xor U22125 (N_22125,N_21729,N_21758);
nand U22126 (N_22126,N_21950,N_21872);
or U22127 (N_22127,N_21814,N_21744);
or U22128 (N_22128,N_21844,N_21883);
xor U22129 (N_22129,N_21680,N_21606);
nand U22130 (N_22130,N_21943,N_21731);
nor U22131 (N_22131,N_21513,N_21652);
and U22132 (N_22132,N_21999,N_21884);
xor U22133 (N_22133,N_21951,N_21530);
and U22134 (N_22134,N_21817,N_21550);
nand U22135 (N_22135,N_21767,N_21949);
xnor U22136 (N_22136,N_21723,N_21957);
nand U22137 (N_22137,N_21724,N_21622);
nand U22138 (N_22138,N_21921,N_21932);
or U22139 (N_22139,N_21975,N_21873);
or U22140 (N_22140,N_21877,N_21952);
nor U22141 (N_22141,N_21522,N_21730);
xor U22142 (N_22142,N_21616,N_21800);
and U22143 (N_22143,N_21638,N_21986);
or U22144 (N_22144,N_21619,N_21970);
or U22145 (N_22145,N_21529,N_21727);
nor U22146 (N_22146,N_21903,N_21897);
and U22147 (N_22147,N_21918,N_21551);
nand U22148 (N_22148,N_21771,N_21625);
or U22149 (N_22149,N_21643,N_21752);
or U22150 (N_22150,N_21865,N_21961);
nor U22151 (N_22151,N_21688,N_21753);
or U22152 (N_22152,N_21764,N_21946);
and U22153 (N_22153,N_21574,N_21524);
or U22154 (N_22154,N_21924,N_21807);
or U22155 (N_22155,N_21628,N_21927);
nor U22156 (N_22156,N_21997,N_21839);
nand U22157 (N_22157,N_21851,N_21782);
or U22158 (N_22158,N_21741,N_21746);
nand U22159 (N_22159,N_21636,N_21781);
nor U22160 (N_22160,N_21852,N_21748);
nor U22161 (N_22161,N_21820,N_21880);
or U22162 (N_22162,N_21992,N_21547);
nor U22163 (N_22163,N_21841,N_21599);
nand U22164 (N_22164,N_21556,N_21571);
and U22165 (N_22165,N_21527,N_21609);
and U22166 (N_22166,N_21778,N_21691);
nor U22167 (N_22167,N_21541,N_21791);
xor U22168 (N_22168,N_21948,N_21570);
xor U22169 (N_22169,N_21544,N_21756);
or U22170 (N_22170,N_21818,N_21641);
nand U22171 (N_22171,N_21660,N_21998);
and U22172 (N_22172,N_21692,N_21555);
nor U22173 (N_22173,N_21969,N_21874);
nor U22174 (N_22174,N_21828,N_21869);
nor U22175 (N_22175,N_21929,N_21859);
and U22176 (N_22176,N_21985,N_21608);
or U22177 (N_22177,N_21515,N_21642);
nor U22178 (N_22178,N_21763,N_21806);
xnor U22179 (N_22179,N_21939,N_21906);
xor U22180 (N_22180,N_21634,N_21668);
nor U22181 (N_22181,N_21709,N_21789);
nand U22182 (N_22182,N_21893,N_21788);
xor U22183 (N_22183,N_21765,N_21813);
or U22184 (N_22184,N_21812,N_21977);
xnor U22185 (N_22185,N_21915,N_21941);
nand U22186 (N_22186,N_21706,N_21749);
and U22187 (N_22187,N_21678,N_21892);
and U22188 (N_22188,N_21834,N_21648);
and U22189 (N_22189,N_21964,N_21989);
nand U22190 (N_22190,N_21902,N_21830);
or U22191 (N_22191,N_21775,N_21565);
nand U22192 (N_22192,N_21587,N_21669);
and U22193 (N_22193,N_21647,N_21510);
and U22194 (N_22194,N_21790,N_21847);
nand U22195 (N_22195,N_21799,N_21572);
and U22196 (N_22196,N_21518,N_21512);
xor U22197 (N_22197,N_21821,N_21875);
xnor U22198 (N_22198,N_21501,N_21933);
and U22199 (N_22199,N_21603,N_21861);
nand U22200 (N_22200,N_21747,N_21554);
or U22201 (N_22201,N_21742,N_21693);
xnor U22202 (N_22202,N_21736,N_21503);
xnor U22203 (N_22203,N_21639,N_21635);
nand U22204 (N_22204,N_21966,N_21797);
and U22205 (N_22205,N_21974,N_21925);
nand U22206 (N_22206,N_21843,N_21905);
and U22207 (N_22207,N_21559,N_21968);
or U22208 (N_22208,N_21532,N_21928);
xor U22209 (N_22209,N_21720,N_21804);
and U22210 (N_22210,N_21837,N_21664);
xnor U22211 (N_22211,N_21784,N_21563);
xor U22212 (N_22212,N_21537,N_21739);
and U22213 (N_22213,N_21624,N_21912);
xor U22214 (N_22214,N_21722,N_21971);
or U22215 (N_22215,N_21732,N_21743);
nand U22216 (N_22216,N_21848,N_21545);
xnor U22217 (N_22217,N_21677,N_21650);
nor U22218 (N_22218,N_21777,N_21868);
nand U22219 (N_22219,N_21965,N_21725);
and U22220 (N_22220,N_21981,N_21602);
nor U22221 (N_22221,N_21626,N_21904);
or U22222 (N_22222,N_21614,N_21979);
and U22223 (N_22223,N_21882,N_21864);
nor U22224 (N_22224,N_21715,N_21577);
xor U22225 (N_22225,N_21983,N_21595);
nor U22226 (N_22226,N_21910,N_21689);
nor U22227 (N_22227,N_21611,N_21801);
and U22228 (N_22228,N_21750,N_21685);
and U22229 (N_22229,N_21772,N_21521);
nand U22230 (N_22230,N_21745,N_21514);
nand U22231 (N_22231,N_21733,N_21825);
nand U22232 (N_22232,N_21683,N_21930);
xnor U22233 (N_22233,N_21594,N_21708);
nand U22234 (N_22234,N_21612,N_21803);
xor U22235 (N_22235,N_21546,N_21617);
nor U22236 (N_22236,N_21502,N_21661);
nand U22237 (N_22237,N_21630,N_21721);
or U22238 (N_22238,N_21506,N_21701);
nand U22239 (N_22239,N_21920,N_21984);
or U22240 (N_22240,N_21575,N_21836);
xnor U22241 (N_22241,N_21786,N_21831);
or U22242 (N_22242,N_21713,N_21662);
xor U22243 (N_22243,N_21856,N_21755);
nand U22244 (N_22244,N_21690,N_21937);
xor U22245 (N_22245,N_21631,N_21900);
or U22246 (N_22246,N_21810,N_21923);
xor U22247 (N_22247,N_21840,N_21536);
xor U22248 (N_22248,N_21881,N_21916);
xnor U22249 (N_22249,N_21995,N_21862);
and U22250 (N_22250,N_21746,N_21865);
nand U22251 (N_22251,N_21876,N_21921);
and U22252 (N_22252,N_21737,N_21644);
or U22253 (N_22253,N_21695,N_21945);
xnor U22254 (N_22254,N_21558,N_21748);
nand U22255 (N_22255,N_21630,N_21843);
and U22256 (N_22256,N_21935,N_21960);
and U22257 (N_22257,N_21507,N_21891);
xnor U22258 (N_22258,N_21979,N_21673);
or U22259 (N_22259,N_21668,N_21575);
or U22260 (N_22260,N_21755,N_21863);
and U22261 (N_22261,N_21750,N_21613);
nor U22262 (N_22262,N_21727,N_21707);
xor U22263 (N_22263,N_21695,N_21525);
nand U22264 (N_22264,N_21856,N_21912);
and U22265 (N_22265,N_21902,N_21775);
and U22266 (N_22266,N_21707,N_21895);
nor U22267 (N_22267,N_21783,N_21527);
and U22268 (N_22268,N_21508,N_21748);
xnor U22269 (N_22269,N_21601,N_21919);
nand U22270 (N_22270,N_21742,N_21779);
or U22271 (N_22271,N_21958,N_21601);
nand U22272 (N_22272,N_21877,N_21862);
and U22273 (N_22273,N_21744,N_21623);
and U22274 (N_22274,N_21732,N_21985);
and U22275 (N_22275,N_21939,N_21878);
xnor U22276 (N_22276,N_21935,N_21665);
xnor U22277 (N_22277,N_21698,N_21934);
and U22278 (N_22278,N_21731,N_21634);
nor U22279 (N_22279,N_21830,N_21900);
xnor U22280 (N_22280,N_21689,N_21815);
or U22281 (N_22281,N_21510,N_21724);
nor U22282 (N_22282,N_21629,N_21768);
nor U22283 (N_22283,N_21581,N_21596);
nand U22284 (N_22284,N_21511,N_21736);
or U22285 (N_22285,N_21886,N_21715);
nor U22286 (N_22286,N_21921,N_21897);
nor U22287 (N_22287,N_21696,N_21911);
nor U22288 (N_22288,N_21891,N_21549);
nor U22289 (N_22289,N_21974,N_21857);
or U22290 (N_22290,N_21564,N_21520);
or U22291 (N_22291,N_21682,N_21756);
xor U22292 (N_22292,N_21767,N_21918);
and U22293 (N_22293,N_21771,N_21783);
and U22294 (N_22294,N_21595,N_21759);
nor U22295 (N_22295,N_21526,N_21551);
or U22296 (N_22296,N_21886,N_21663);
nor U22297 (N_22297,N_21674,N_21911);
nor U22298 (N_22298,N_21988,N_21614);
nor U22299 (N_22299,N_21891,N_21673);
or U22300 (N_22300,N_21904,N_21701);
xor U22301 (N_22301,N_21596,N_21529);
and U22302 (N_22302,N_21635,N_21802);
or U22303 (N_22303,N_21895,N_21586);
or U22304 (N_22304,N_21611,N_21662);
and U22305 (N_22305,N_21796,N_21728);
nor U22306 (N_22306,N_21984,N_21811);
or U22307 (N_22307,N_21703,N_21505);
and U22308 (N_22308,N_21891,N_21614);
nand U22309 (N_22309,N_21807,N_21990);
nand U22310 (N_22310,N_21903,N_21878);
nand U22311 (N_22311,N_21721,N_21762);
nor U22312 (N_22312,N_21716,N_21773);
xnor U22313 (N_22313,N_21506,N_21975);
nor U22314 (N_22314,N_21879,N_21582);
or U22315 (N_22315,N_21850,N_21567);
nor U22316 (N_22316,N_21915,N_21744);
nand U22317 (N_22317,N_21954,N_21582);
xnor U22318 (N_22318,N_21639,N_21637);
or U22319 (N_22319,N_21599,N_21692);
or U22320 (N_22320,N_21514,N_21824);
xnor U22321 (N_22321,N_21707,N_21705);
or U22322 (N_22322,N_21592,N_21501);
and U22323 (N_22323,N_21761,N_21774);
or U22324 (N_22324,N_21959,N_21977);
and U22325 (N_22325,N_21932,N_21938);
or U22326 (N_22326,N_21807,N_21766);
xor U22327 (N_22327,N_21917,N_21568);
and U22328 (N_22328,N_21810,N_21595);
xor U22329 (N_22329,N_21902,N_21699);
and U22330 (N_22330,N_21794,N_21596);
or U22331 (N_22331,N_21522,N_21891);
xor U22332 (N_22332,N_21893,N_21541);
nand U22333 (N_22333,N_21869,N_21891);
nand U22334 (N_22334,N_21688,N_21903);
and U22335 (N_22335,N_21869,N_21520);
xor U22336 (N_22336,N_21719,N_21923);
xor U22337 (N_22337,N_21798,N_21640);
xor U22338 (N_22338,N_21750,N_21607);
or U22339 (N_22339,N_21992,N_21527);
and U22340 (N_22340,N_21687,N_21930);
or U22341 (N_22341,N_21517,N_21761);
or U22342 (N_22342,N_21595,N_21924);
and U22343 (N_22343,N_21624,N_21709);
nand U22344 (N_22344,N_21848,N_21772);
or U22345 (N_22345,N_21988,N_21722);
nand U22346 (N_22346,N_21974,N_21991);
xnor U22347 (N_22347,N_21538,N_21890);
or U22348 (N_22348,N_21946,N_21710);
nand U22349 (N_22349,N_21677,N_21819);
xnor U22350 (N_22350,N_21902,N_21704);
and U22351 (N_22351,N_21615,N_21899);
nand U22352 (N_22352,N_21932,N_21766);
nor U22353 (N_22353,N_21507,N_21890);
or U22354 (N_22354,N_21599,N_21903);
or U22355 (N_22355,N_21985,N_21945);
nand U22356 (N_22356,N_21623,N_21552);
xnor U22357 (N_22357,N_21705,N_21828);
nand U22358 (N_22358,N_21859,N_21545);
or U22359 (N_22359,N_21552,N_21658);
nor U22360 (N_22360,N_21825,N_21513);
nand U22361 (N_22361,N_21633,N_21546);
or U22362 (N_22362,N_21707,N_21560);
or U22363 (N_22363,N_21614,N_21641);
nand U22364 (N_22364,N_21635,N_21718);
or U22365 (N_22365,N_21999,N_21804);
xnor U22366 (N_22366,N_21688,N_21572);
nor U22367 (N_22367,N_21594,N_21638);
nand U22368 (N_22368,N_21889,N_21722);
nand U22369 (N_22369,N_21594,N_21685);
xor U22370 (N_22370,N_21532,N_21761);
or U22371 (N_22371,N_21710,N_21745);
nor U22372 (N_22372,N_21663,N_21889);
xnor U22373 (N_22373,N_21563,N_21832);
nand U22374 (N_22374,N_21786,N_21986);
nor U22375 (N_22375,N_21790,N_21705);
or U22376 (N_22376,N_21543,N_21526);
nand U22377 (N_22377,N_21862,N_21660);
and U22378 (N_22378,N_21730,N_21619);
xnor U22379 (N_22379,N_21577,N_21557);
nor U22380 (N_22380,N_21583,N_21690);
or U22381 (N_22381,N_21937,N_21963);
and U22382 (N_22382,N_21809,N_21525);
and U22383 (N_22383,N_21707,N_21782);
nand U22384 (N_22384,N_21731,N_21589);
xnor U22385 (N_22385,N_21768,N_21517);
nand U22386 (N_22386,N_21748,N_21523);
nor U22387 (N_22387,N_21565,N_21752);
nand U22388 (N_22388,N_21885,N_21566);
and U22389 (N_22389,N_21586,N_21991);
xor U22390 (N_22390,N_21622,N_21926);
and U22391 (N_22391,N_21565,N_21911);
or U22392 (N_22392,N_21842,N_21714);
xor U22393 (N_22393,N_21615,N_21674);
and U22394 (N_22394,N_21798,N_21613);
nor U22395 (N_22395,N_21504,N_21841);
and U22396 (N_22396,N_21593,N_21777);
nor U22397 (N_22397,N_21631,N_21618);
or U22398 (N_22398,N_21669,N_21589);
and U22399 (N_22399,N_21701,N_21985);
xor U22400 (N_22400,N_21685,N_21860);
and U22401 (N_22401,N_21774,N_21746);
or U22402 (N_22402,N_21702,N_21519);
or U22403 (N_22403,N_21586,N_21510);
nor U22404 (N_22404,N_21888,N_21582);
nand U22405 (N_22405,N_21813,N_21827);
xnor U22406 (N_22406,N_21993,N_21778);
nor U22407 (N_22407,N_21851,N_21588);
and U22408 (N_22408,N_21707,N_21706);
nand U22409 (N_22409,N_21500,N_21855);
xnor U22410 (N_22410,N_21864,N_21701);
and U22411 (N_22411,N_21649,N_21742);
nand U22412 (N_22412,N_21561,N_21877);
and U22413 (N_22413,N_21826,N_21746);
nor U22414 (N_22414,N_21627,N_21709);
nor U22415 (N_22415,N_21944,N_21745);
nor U22416 (N_22416,N_21593,N_21891);
nor U22417 (N_22417,N_21787,N_21735);
xor U22418 (N_22418,N_21754,N_21943);
xor U22419 (N_22419,N_21529,N_21679);
nor U22420 (N_22420,N_21891,N_21706);
nor U22421 (N_22421,N_21676,N_21884);
nand U22422 (N_22422,N_21599,N_21962);
or U22423 (N_22423,N_21567,N_21578);
xnor U22424 (N_22424,N_21512,N_21888);
nand U22425 (N_22425,N_21609,N_21709);
nor U22426 (N_22426,N_21751,N_21957);
and U22427 (N_22427,N_21995,N_21772);
xor U22428 (N_22428,N_21795,N_21578);
nand U22429 (N_22429,N_21680,N_21715);
xor U22430 (N_22430,N_21745,N_21963);
nor U22431 (N_22431,N_21750,N_21906);
and U22432 (N_22432,N_21860,N_21527);
nand U22433 (N_22433,N_21743,N_21673);
nand U22434 (N_22434,N_21831,N_21793);
or U22435 (N_22435,N_21797,N_21597);
xnor U22436 (N_22436,N_21774,N_21781);
nor U22437 (N_22437,N_21925,N_21532);
or U22438 (N_22438,N_21747,N_21692);
xor U22439 (N_22439,N_21735,N_21906);
or U22440 (N_22440,N_21590,N_21514);
xnor U22441 (N_22441,N_21620,N_21758);
or U22442 (N_22442,N_21772,N_21752);
nand U22443 (N_22443,N_21930,N_21751);
and U22444 (N_22444,N_21709,N_21711);
nand U22445 (N_22445,N_21845,N_21880);
nor U22446 (N_22446,N_21832,N_21950);
and U22447 (N_22447,N_21974,N_21506);
xor U22448 (N_22448,N_21707,N_21684);
and U22449 (N_22449,N_21868,N_21855);
nand U22450 (N_22450,N_21750,N_21520);
or U22451 (N_22451,N_21932,N_21664);
xor U22452 (N_22452,N_21885,N_21733);
and U22453 (N_22453,N_21658,N_21865);
xnor U22454 (N_22454,N_21516,N_21653);
or U22455 (N_22455,N_21918,N_21785);
nor U22456 (N_22456,N_21602,N_21687);
or U22457 (N_22457,N_21517,N_21914);
nor U22458 (N_22458,N_21663,N_21902);
nand U22459 (N_22459,N_21991,N_21812);
nor U22460 (N_22460,N_21604,N_21730);
nor U22461 (N_22461,N_21768,N_21668);
xor U22462 (N_22462,N_21565,N_21655);
nor U22463 (N_22463,N_21839,N_21965);
xor U22464 (N_22464,N_21801,N_21923);
xor U22465 (N_22465,N_21641,N_21595);
xor U22466 (N_22466,N_21958,N_21634);
and U22467 (N_22467,N_21944,N_21813);
or U22468 (N_22468,N_21906,N_21757);
and U22469 (N_22469,N_21856,N_21926);
and U22470 (N_22470,N_21820,N_21919);
or U22471 (N_22471,N_21522,N_21828);
nand U22472 (N_22472,N_21808,N_21708);
nand U22473 (N_22473,N_21680,N_21764);
nand U22474 (N_22474,N_21550,N_21910);
and U22475 (N_22475,N_21590,N_21964);
nor U22476 (N_22476,N_21748,N_21866);
nand U22477 (N_22477,N_21624,N_21839);
nand U22478 (N_22478,N_21972,N_21629);
and U22479 (N_22479,N_21784,N_21811);
or U22480 (N_22480,N_21519,N_21844);
and U22481 (N_22481,N_21834,N_21606);
nand U22482 (N_22482,N_21628,N_21566);
nor U22483 (N_22483,N_21846,N_21621);
xor U22484 (N_22484,N_21844,N_21773);
nor U22485 (N_22485,N_21905,N_21934);
or U22486 (N_22486,N_21550,N_21644);
or U22487 (N_22487,N_21604,N_21763);
or U22488 (N_22488,N_21883,N_21876);
nand U22489 (N_22489,N_21578,N_21690);
or U22490 (N_22490,N_21785,N_21763);
nor U22491 (N_22491,N_21523,N_21846);
and U22492 (N_22492,N_21924,N_21987);
nand U22493 (N_22493,N_21568,N_21875);
nand U22494 (N_22494,N_21650,N_21985);
nor U22495 (N_22495,N_21769,N_21845);
xor U22496 (N_22496,N_21918,N_21507);
xor U22497 (N_22497,N_21530,N_21680);
nor U22498 (N_22498,N_21695,N_21670);
and U22499 (N_22499,N_21816,N_21608);
xor U22500 (N_22500,N_22421,N_22283);
and U22501 (N_22501,N_22413,N_22048);
nor U22502 (N_22502,N_22065,N_22443);
nand U22503 (N_22503,N_22030,N_22312);
nor U22504 (N_22504,N_22266,N_22394);
or U22505 (N_22505,N_22370,N_22407);
and U22506 (N_22506,N_22287,N_22158);
xnor U22507 (N_22507,N_22078,N_22044);
or U22508 (N_22508,N_22039,N_22476);
or U22509 (N_22509,N_22187,N_22079);
nand U22510 (N_22510,N_22398,N_22483);
or U22511 (N_22511,N_22325,N_22465);
xor U22512 (N_22512,N_22401,N_22128);
xor U22513 (N_22513,N_22264,N_22347);
and U22514 (N_22514,N_22029,N_22014);
and U22515 (N_22515,N_22049,N_22258);
nand U22516 (N_22516,N_22327,N_22136);
xnor U22517 (N_22517,N_22404,N_22367);
nand U22518 (N_22518,N_22383,N_22113);
and U22519 (N_22519,N_22038,N_22164);
or U22520 (N_22520,N_22084,N_22461);
or U22521 (N_22521,N_22174,N_22279);
or U22522 (N_22522,N_22234,N_22212);
nor U22523 (N_22523,N_22220,N_22442);
nand U22524 (N_22524,N_22425,N_22462);
and U22525 (N_22525,N_22345,N_22179);
or U22526 (N_22526,N_22356,N_22057);
xnor U22527 (N_22527,N_22467,N_22321);
xnor U22528 (N_22528,N_22286,N_22047);
or U22529 (N_22529,N_22458,N_22419);
and U22530 (N_22530,N_22184,N_22352);
or U22531 (N_22531,N_22351,N_22455);
nor U22532 (N_22532,N_22041,N_22357);
and U22533 (N_22533,N_22378,N_22021);
nor U22534 (N_22534,N_22059,N_22478);
or U22535 (N_22535,N_22097,N_22219);
xnor U22536 (N_22536,N_22228,N_22430);
or U22537 (N_22537,N_22449,N_22160);
or U22538 (N_22538,N_22484,N_22278);
nand U22539 (N_22539,N_22252,N_22306);
xor U22540 (N_22540,N_22472,N_22412);
nor U22541 (N_22541,N_22226,N_22077);
and U22542 (N_22542,N_22121,N_22124);
and U22543 (N_22543,N_22263,N_22218);
xnor U22544 (N_22544,N_22155,N_22410);
nor U22545 (N_22545,N_22199,N_22202);
or U22546 (N_22546,N_22067,N_22102);
nor U22547 (N_22547,N_22395,N_22365);
nand U22548 (N_22548,N_22125,N_22399);
nor U22549 (N_22549,N_22303,N_22471);
nor U22550 (N_22550,N_22388,N_22492);
nor U22551 (N_22551,N_22106,N_22093);
nor U22552 (N_22552,N_22230,N_22298);
and U22553 (N_22553,N_22181,N_22004);
or U22554 (N_22554,N_22046,N_22499);
nand U22555 (N_22555,N_22151,N_22115);
xor U22556 (N_22556,N_22104,N_22261);
xor U22557 (N_22557,N_22265,N_22469);
nor U22558 (N_22558,N_22320,N_22337);
or U22559 (N_22559,N_22364,N_22127);
or U22560 (N_22560,N_22451,N_22169);
nor U22561 (N_22561,N_22267,N_22387);
and U22562 (N_22562,N_22052,N_22223);
xnor U22563 (N_22563,N_22371,N_22050);
or U22564 (N_22564,N_22335,N_22385);
xnor U22565 (N_22565,N_22207,N_22361);
xnor U22566 (N_22566,N_22015,N_22118);
or U22567 (N_22567,N_22132,N_22200);
nand U22568 (N_22568,N_22488,N_22318);
nand U22569 (N_22569,N_22209,N_22232);
nand U22570 (N_22570,N_22354,N_22302);
and U22571 (N_22571,N_22444,N_22491);
or U22572 (N_22572,N_22073,N_22297);
nor U22573 (N_22573,N_22313,N_22391);
or U22574 (N_22574,N_22288,N_22058);
xnor U22575 (N_22575,N_22055,N_22149);
and U22576 (N_22576,N_22099,N_22482);
and U22577 (N_22577,N_22333,N_22344);
and U22578 (N_22578,N_22146,N_22315);
or U22579 (N_22579,N_22225,N_22418);
nor U22580 (N_22580,N_22109,N_22437);
nor U22581 (N_22581,N_22386,N_22075);
nand U22582 (N_22582,N_22245,N_22054);
xor U22583 (N_22583,N_22138,N_22163);
nand U22584 (N_22584,N_22363,N_22249);
xnor U22585 (N_22585,N_22002,N_22170);
nand U22586 (N_22586,N_22439,N_22331);
and U22587 (N_22587,N_22289,N_22020);
nand U22588 (N_22588,N_22142,N_22148);
xnor U22589 (N_22589,N_22456,N_22119);
xor U22590 (N_22590,N_22237,N_22446);
or U22591 (N_22591,N_22082,N_22305);
nand U22592 (N_22592,N_22229,N_22098);
or U22593 (N_22593,N_22427,N_22440);
or U22594 (N_22594,N_22380,N_22141);
xor U22595 (N_22595,N_22025,N_22396);
xnor U22596 (N_22596,N_22424,N_22248);
xor U22597 (N_22597,N_22271,N_22003);
nand U22598 (N_22598,N_22420,N_22019);
nand U22599 (N_22599,N_22296,N_22210);
nand U22600 (N_22600,N_22096,N_22080);
nor U22601 (N_22601,N_22022,N_22381);
xor U22602 (N_22602,N_22459,N_22417);
or U22603 (N_22603,N_22276,N_22183);
and U22604 (N_22604,N_22134,N_22092);
nand U22605 (N_22605,N_22193,N_22322);
nand U22606 (N_22606,N_22463,N_22208);
nor U22607 (N_22607,N_22088,N_22165);
nor U22608 (N_22608,N_22423,N_22368);
nand U22609 (N_22609,N_22076,N_22133);
nand U22610 (N_22610,N_22480,N_22262);
or U22611 (N_22611,N_22185,N_22481);
xor U22612 (N_22612,N_22013,N_22280);
or U22613 (N_22613,N_22091,N_22120);
nand U22614 (N_22614,N_22176,N_22285);
and U22615 (N_22615,N_22274,N_22194);
and U22616 (N_22616,N_22154,N_22445);
nor U22617 (N_22617,N_22301,N_22083);
nor U22618 (N_22618,N_22196,N_22317);
or U22619 (N_22619,N_22291,N_22172);
nor U22620 (N_22620,N_22246,N_22143);
nand U22621 (N_22621,N_22316,N_22206);
and U22622 (N_22622,N_22475,N_22485);
nor U22623 (N_22623,N_22253,N_22379);
nor U22624 (N_22624,N_22400,N_22338);
nor U22625 (N_22625,N_22374,N_22069);
nor U22626 (N_22626,N_22032,N_22498);
nand U22627 (N_22627,N_22175,N_22191);
nor U22628 (N_22628,N_22332,N_22457);
and U22629 (N_22629,N_22273,N_22023);
xor U22630 (N_22630,N_22006,N_22348);
or U22631 (N_22631,N_22366,N_22094);
nor U22632 (N_22632,N_22236,N_22086);
or U22633 (N_22633,N_22359,N_22182);
and U22634 (N_22634,N_22114,N_22043);
xnor U22635 (N_22635,N_22215,N_22438);
nand U22636 (N_22636,N_22240,N_22453);
nor U22637 (N_22637,N_22349,N_22275);
or U22638 (N_22638,N_22045,N_22452);
nand U22639 (N_22639,N_22064,N_22177);
xor U22640 (N_22640,N_22024,N_22293);
nor U22641 (N_22641,N_22190,N_22428);
or U22642 (N_22642,N_22493,N_22309);
nor U22643 (N_22643,N_22152,N_22000);
or U22644 (N_22644,N_22239,N_22355);
xor U22645 (N_22645,N_22435,N_22168);
nor U22646 (N_22646,N_22139,N_22340);
or U22647 (N_22647,N_22203,N_22072);
and U22648 (N_22648,N_22007,N_22161);
nand U22649 (N_22649,N_22429,N_22377);
nor U22650 (N_22650,N_22450,N_22005);
nor U22651 (N_22651,N_22147,N_22292);
nor U22652 (N_22652,N_22162,N_22254);
or U22653 (N_22653,N_22350,N_22300);
nand U22654 (N_22654,N_22495,N_22010);
xnor U22655 (N_22655,N_22235,N_22085);
nor U22656 (N_22656,N_22360,N_22295);
nand U22657 (N_22657,N_22108,N_22211);
nor U22658 (N_22658,N_22042,N_22342);
or U22659 (N_22659,N_22466,N_22105);
xor U22660 (N_22660,N_22403,N_22018);
nor U22661 (N_22661,N_22037,N_22195);
nor U22662 (N_22662,N_22402,N_22129);
nand U22663 (N_22663,N_22110,N_22216);
xnor U22664 (N_22664,N_22307,N_22408);
nor U22665 (N_22665,N_22397,N_22343);
nand U22666 (N_22666,N_22272,N_22330);
or U22667 (N_22667,N_22426,N_22101);
or U22668 (N_22668,N_22242,N_22479);
xnor U22669 (N_22669,N_22198,N_22173);
or U22670 (N_22670,N_22062,N_22081);
xnor U22671 (N_22671,N_22087,N_22167);
nand U22672 (N_22672,N_22411,N_22433);
xor U22673 (N_22673,N_22319,N_22066);
or U22674 (N_22674,N_22233,N_22497);
xor U22675 (N_22675,N_22329,N_22409);
or U22676 (N_22676,N_22178,N_22186);
nand U22677 (N_22677,N_22448,N_22474);
xor U22678 (N_22678,N_22157,N_22063);
nor U22679 (N_22679,N_22489,N_22144);
nor U22680 (N_22680,N_22323,N_22464);
nand U22681 (N_22681,N_22270,N_22434);
nand U22682 (N_22682,N_22454,N_22028);
and U22683 (N_22683,N_22334,N_22166);
nor U22684 (N_22684,N_22494,N_22221);
or U22685 (N_22685,N_22477,N_22375);
nand U22686 (N_22686,N_22192,N_22011);
and U22687 (N_22687,N_22369,N_22204);
xor U22688 (N_22688,N_22487,N_22432);
xnor U22689 (N_22689,N_22311,N_22040);
nor U22690 (N_22690,N_22036,N_22259);
and U22691 (N_22691,N_22009,N_22051);
xor U22692 (N_22692,N_22189,N_22470);
nor U22693 (N_22693,N_22241,N_22224);
or U22694 (N_22694,N_22071,N_22310);
nor U22695 (N_22695,N_22180,N_22460);
nor U22696 (N_22696,N_22447,N_22281);
or U22697 (N_22697,N_22415,N_22171);
xor U22698 (N_22698,N_22339,N_22089);
xnor U22699 (N_22699,N_22257,N_22214);
and U22700 (N_22700,N_22060,N_22314);
nand U22701 (N_22701,N_22358,N_22056);
xnor U22702 (N_22702,N_22269,N_22490);
and U22703 (N_22703,N_22250,N_22341);
nor U22704 (N_22704,N_22244,N_22131);
xnor U22705 (N_22705,N_22392,N_22103);
or U22706 (N_22706,N_22197,N_22393);
nor U22707 (N_22707,N_22243,N_22035);
and U22708 (N_22708,N_22008,N_22026);
nand U22709 (N_22709,N_22145,N_22255);
nor U22710 (N_22710,N_22227,N_22112);
and U22711 (N_22711,N_22390,N_22282);
and U22712 (N_22712,N_22140,N_22150);
xnor U22713 (N_22713,N_22441,N_22159);
nand U22714 (N_22714,N_22033,N_22473);
or U22715 (N_22715,N_22017,N_22130);
nand U22716 (N_22716,N_22336,N_22123);
or U22717 (N_22717,N_22111,N_22436);
nand U22718 (N_22718,N_22251,N_22308);
or U22719 (N_22719,N_22422,N_22362);
and U22720 (N_22720,N_22256,N_22486);
nor U22721 (N_22721,N_22290,N_22095);
nor U22722 (N_22722,N_22372,N_22012);
xnor U22723 (N_22723,N_22201,N_22496);
nor U22724 (N_22724,N_22034,N_22068);
and U22725 (N_22725,N_22299,N_22268);
xnor U22726 (N_22726,N_22090,N_22382);
or U22727 (N_22727,N_22326,N_22188);
and U22728 (N_22728,N_22294,N_22431);
nand U22729 (N_22729,N_22153,N_22070);
and U22730 (N_22730,N_22156,N_22414);
or U22731 (N_22731,N_22328,N_22061);
nor U22732 (N_22732,N_22031,N_22416);
or U22733 (N_22733,N_22406,N_22384);
nand U22734 (N_22734,N_22074,N_22137);
or U22735 (N_22735,N_22389,N_22053);
xnor U22736 (N_22736,N_22231,N_22222);
xor U22737 (N_22737,N_22260,N_22117);
xor U22738 (N_22738,N_22107,N_22213);
and U22739 (N_22739,N_22135,N_22284);
or U22740 (N_22740,N_22373,N_22122);
nand U22741 (N_22741,N_22217,N_22016);
nor U22742 (N_22742,N_22126,N_22277);
or U22743 (N_22743,N_22405,N_22324);
nor U22744 (N_22744,N_22001,N_22346);
and U22745 (N_22745,N_22100,N_22304);
nor U22746 (N_22746,N_22238,N_22247);
nand U22747 (N_22747,N_22353,N_22376);
nand U22748 (N_22748,N_22468,N_22027);
nand U22749 (N_22749,N_22205,N_22116);
or U22750 (N_22750,N_22350,N_22380);
xnor U22751 (N_22751,N_22121,N_22475);
xor U22752 (N_22752,N_22230,N_22426);
and U22753 (N_22753,N_22264,N_22390);
and U22754 (N_22754,N_22292,N_22458);
and U22755 (N_22755,N_22101,N_22120);
nand U22756 (N_22756,N_22010,N_22002);
nor U22757 (N_22757,N_22364,N_22295);
xnor U22758 (N_22758,N_22068,N_22373);
nand U22759 (N_22759,N_22156,N_22179);
nand U22760 (N_22760,N_22061,N_22038);
nor U22761 (N_22761,N_22088,N_22429);
xnor U22762 (N_22762,N_22497,N_22357);
nor U22763 (N_22763,N_22051,N_22469);
nor U22764 (N_22764,N_22082,N_22173);
nor U22765 (N_22765,N_22347,N_22260);
and U22766 (N_22766,N_22409,N_22191);
nor U22767 (N_22767,N_22478,N_22454);
nor U22768 (N_22768,N_22186,N_22068);
xor U22769 (N_22769,N_22029,N_22283);
and U22770 (N_22770,N_22498,N_22179);
or U22771 (N_22771,N_22477,N_22394);
or U22772 (N_22772,N_22061,N_22249);
xnor U22773 (N_22773,N_22352,N_22286);
nand U22774 (N_22774,N_22149,N_22200);
xnor U22775 (N_22775,N_22325,N_22045);
xor U22776 (N_22776,N_22148,N_22092);
or U22777 (N_22777,N_22489,N_22499);
nand U22778 (N_22778,N_22220,N_22091);
or U22779 (N_22779,N_22185,N_22162);
nand U22780 (N_22780,N_22245,N_22016);
xor U22781 (N_22781,N_22343,N_22069);
nor U22782 (N_22782,N_22322,N_22299);
nand U22783 (N_22783,N_22297,N_22159);
nor U22784 (N_22784,N_22429,N_22396);
xor U22785 (N_22785,N_22422,N_22026);
and U22786 (N_22786,N_22481,N_22304);
nand U22787 (N_22787,N_22155,N_22113);
or U22788 (N_22788,N_22208,N_22256);
xnor U22789 (N_22789,N_22204,N_22363);
nand U22790 (N_22790,N_22378,N_22101);
nor U22791 (N_22791,N_22449,N_22317);
and U22792 (N_22792,N_22222,N_22446);
xor U22793 (N_22793,N_22000,N_22376);
and U22794 (N_22794,N_22375,N_22354);
nand U22795 (N_22795,N_22424,N_22474);
xor U22796 (N_22796,N_22496,N_22418);
or U22797 (N_22797,N_22413,N_22194);
nor U22798 (N_22798,N_22393,N_22065);
or U22799 (N_22799,N_22192,N_22366);
nor U22800 (N_22800,N_22458,N_22453);
nand U22801 (N_22801,N_22056,N_22355);
nand U22802 (N_22802,N_22137,N_22133);
nor U22803 (N_22803,N_22092,N_22388);
and U22804 (N_22804,N_22229,N_22217);
nor U22805 (N_22805,N_22027,N_22035);
xor U22806 (N_22806,N_22110,N_22189);
and U22807 (N_22807,N_22047,N_22353);
nor U22808 (N_22808,N_22338,N_22444);
or U22809 (N_22809,N_22017,N_22254);
nand U22810 (N_22810,N_22359,N_22349);
nor U22811 (N_22811,N_22056,N_22396);
nor U22812 (N_22812,N_22224,N_22439);
xnor U22813 (N_22813,N_22391,N_22074);
and U22814 (N_22814,N_22455,N_22336);
and U22815 (N_22815,N_22274,N_22450);
nand U22816 (N_22816,N_22254,N_22048);
nor U22817 (N_22817,N_22159,N_22493);
xor U22818 (N_22818,N_22054,N_22374);
nand U22819 (N_22819,N_22265,N_22303);
and U22820 (N_22820,N_22276,N_22176);
or U22821 (N_22821,N_22398,N_22031);
xnor U22822 (N_22822,N_22304,N_22229);
and U22823 (N_22823,N_22180,N_22181);
nor U22824 (N_22824,N_22295,N_22344);
nor U22825 (N_22825,N_22190,N_22427);
and U22826 (N_22826,N_22263,N_22470);
xor U22827 (N_22827,N_22222,N_22358);
nor U22828 (N_22828,N_22368,N_22031);
nor U22829 (N_22829,N_22105,N_22249);
or U22830 (N_22830,N_22412,N_22422);
xnor U22831 (N_22831,N_22218,N_22195);
or U22832 (N_22832,N_22284,N_22181);
or U22833 (N_22833,N_22209,N_22255);
and U22834 (N_22834,N_22050,N_22196);
nand U22835 (N_22835,N_22216,N_22036);
nor U22836 (N_22836,N_22147,N_22041);
and U22837 (N_22837,N_22281,N_22023);
and U22838 (N_22838,N_22369,N_22366);
or U22839 (N_22839,N_22342,N_22225);
or U22840 (N_22840,N_22267,N_22021);
or U22841 (N_22841,N_22062,N_22044);
and U22842 (N_22842,N_22340,N_22467);
nor U22843 (N_22843,N_22199,N_22324);
or U22844 (N_22844,N_22399,N_22205);
nor U22845 (N_22845,N_22062,N_22257);
and U22846 (N_22846,N_22071,N_22050);
xnor U22847 (N_22847,N_22464,N_22236);
xor U22848 (N_22848,N_22397,N_22234);
nor U22849 (N_22849,N_22401,N_22258);
nand U22850 (N_22850,N_22495,N_22120);
nand U22851 (N_22851,N_22284,N_22064);
xnor U22852 (N_22852,N_22285,N_22452);
xnor U22853 (N_22853,N_22279,N_22113);
nor U22854 (N_22854,N_22300,N_22459);
or U22855 (N_22855,N_22035,N_22113);
nor U22856 (N_22856,N_22411,N_22152);
or U22857 (N_22857,N_22358,N_22046);
and U22858 (N_22858,N_22071,N_22260);
or U22859 (N_22859,N_22040,N_22220);
or U22860 (N_22860,N_22312,N_22042);
or U22861 (N_22861,N_22140,N_22072);
nand U22862 (N_22862,N_22272,N_22411);
xor U22863 (N_22863,N_22005,N_22402);
or U22864 (N_22864,N_22089,N_22479);
xor U22865 (N_22865,N_22080,N_22431);
nand U22866 (N_22866,N_22448,N_22195);
nand U22867 (N_22867,N_22188,N_22335);
or U22868 (N_22868,N_22142,N_22360);
nand U22869 (N_22869,N_22138,N_22342);
and U22870 (N_22870,N_22028,N_22439);
and U22871 (N_22871,N_22041,N_22196);
and U22872 (N_22872,N_22493,N_22387);
and U22873 (N_22873,N_22299,N_22053);
and U22874 (N_22874,N_22001,N_22294);
or U22875 (N_22875,N_22184,N_22454);
xnor U22876 (N_22876,N_22455,N_22248);
or U22877 (N_22877,N_22146,N_22015);
xor U22878 (N_22878,N_22356,N_22101);
xnor U22879 (N_22879,N_22417,N_22151);
nand U22880 (N_22880,N_22125,N_22243);
or U22881 (N_22881,N_22212,N_22102);
nand U22882 (N_22882,N_22376,N_22159);
xnor U22883 (N_22883,N_22136,N_22179);
xor U22884 (N_22884,N_22053,N_22218);
xnor U22885 (N_22885,N_22029,N_22438);
nor U22886 (N_22886,N_22153,N_22315);
nand U22887 (N_22887,N_22058,N_22208);
and U22888 (N_22888,N_22256,N_22250);
nor U22889 (N_22889,N_22457,N_22066);
xor U22890 (N_22890,N_22365,N_22225);
xor U22891 (N_22891,N_22057,N_22445);
nand U22892 (N_22892,N_22434,N_22032);
nand U22893 (N_22893,N_22138,N_22403);
nor U22894 (N_22894,N_22390,N_22468);
nand U22895 (N_22895,N_22183,N_22142);
nand U22896 (N_22896,N_22342,N_22398);
xor U22897 (N_22897,N_22375,N_22265);
nand U22898 (N_22898,N_22474,N_22056);
or U22899 (N_22899,N_22032,N_22277);
nand U22900 (N_22900,N_22372,N_22157);
or U22901 (N_22901,N_22186,N_22033);
or U22902 (N_22902,N_22288,N_22258);
nor U22903 (N_22903,N_22074,N_22065);
nor U22904 (N_22904,N_22236,N_22204);
and U22905 (N_22905,N_22465,N_22492);
xnor U22906 (N_22906,N_22207,N_22376);
nor U22907 (N_22907,N_22419,N_22469);
xnor U22908 (N_22908,N_22037,N_22058);
xnor U22909 (N_22909,N_22032,N_22058);
nor U22910 (N_22910,N_22448,N_22158);
and U22911 (N_22911,N_22072,N_22256);
or U22912 (N_22912,N_22385,N_22346);
and U22913 (N_22913,N_22065,N_22246);
and U22914 (N_22914,N_22087,N_22226);
or U22915 (N_22915,N_22150,N_22147);
nor U22916 (N_22916,N_22084,N_22137);
xnor U22917 (N_22917,N_22173,N_22277);
xor U22918 (N_22918,N_22348,N_22413);
xor U22919 (N_22919,N_22409,N_22127);
nor U22920 (N_22920,N_22461,N_22028);
xnor U22921 (N_22921,N_22160,N_22355);
and U22922 (N_22922,N_22101,N_22480);
and U22923 (N_22923,N_22178,N_22012);
and U22924 (N_22924,N_22258,N_22406);
nor U22925 (N_22925,N_22219,N_22423);
xnor U22926 (N_22926,N_22000,N_22213);
or U22927 (N_22927,N_22085,N_22194);
and U22928 (N_22928,N_22334,N_22336);
nand U22929 (N_22929,N_22229,N_22306);
nor U22930 (N_22930,N_22047,N_22114);
nand U22931 (N_22931,N_22183,N_22272);
nand U22932 (N_22932,N_22095,N_22051);
nor U22933 (N_22933,N_22039,N_22056);
nand U22934 (N_22934,N_22078,N_22124);
nand U22935 (N_22935,N_22140,N_22053);
or U22936 (N_22936,N_22076,N_22362);
xor U22937 (N_22937,N_22106,N_22071);
nor U22938 (N_22938,N_22483,N_22405);
nor U22939 (N_22939,N_22218,N_22424);
and U22940 (N_22940,N_22098,N_22039);
nand U22941 (N_22941,N_22113,N_22009);
and U22942 (N_22942,N_22029,N_22171);
nor U22943 (N_22943,N_22451,N_22125);
xnor U22944 (N_22944,N_22415,N_22462);
xor U22945 (N_22945,N_22396,N_22066);
xnor U22946 (N_22946,N_22497,N_22077);
xnor U22947 (N_22947,N_22200,N_22305);
nor U22948 (N_22948,N_22140,N_22001);
nor U22949 (N_22949,N_22327,N_22247);
xnor U22950 (N_22950,N_22201,N_22068);
xnor U22951 (N_22951,N_22031,N_22462);
xor U22952 (N_22952,N_22132,N_22193);
xnor U22953 (N_22953,N_22118,N_22489);
nand U22954 (N_22954,N_22233,N_22346);
nor U22955 (N_22955,N_22412,N_22005);
and U22956 (N_22956,N_22241,N_22220);
nor U22957 (N_22957,N_22456,N_22368);
nand U22958 (N_22958,N_22471,N_22386);
or U22959 (N_22959,N_22235,N_22019);
nand U22960 (N_22960,N_22343,N_22337);
or U22961 (N_22961,N_22130,N_22016);
nor U22962 (N_22962,N_22199,N_22092);
nand U22963 (N_22963,N_22140,N_22409);
and U22964 (N_22964,N_22370,N_22414);
nor U22965 (N_22965,N_22213,N_22313);
xor U22966 (N_22966,N_22406,N_22223);
xor U22967 (N_22967,N_22299,N_22104);
xnor U22968 (N_22968,N_22419,N_22128);
nor U22969 (N_22969,N_22426,N_22146);
nor U22970 (N_22970,N_22258,N_22256);
and U22971 (N_22971,N_22294,N_22315);
nor U22972 (N_22972,N_22158,N_22311);
and U22973 (N_22973,N_22395,N_22147);
and U22974 (N_22974,N_22385,N_22093);
nor U22975 (N_22975,N_22255,N_22312);
nor U22976 (N_22976,N_22346,N_22228);
nor U22977 (N_22977,N_22359,N_22317);
nand U22978 (N_22978,N_22255,N_22293);
nor U22979 (N_22979,N_22393,N_22439);
nand U22980 (N_22980,N_22427,N_22415);
nand U22981 (N_22981,N_22067,N_22440);
or U22982 (N_22982,N_22369,N_22032);
xor U22983 (N_22983,N_22203,N_22204);
xor U22984 (N_22984,N_22103,N_22284);
and U22985 (N_22985,N_22215,N_22497);
nand U22986 (N_22986,N_22043,N_22427);
nor U22987 (N_22987,N_22368,N_22088);
and U22988 (N_22988,N_22470,N_22382);
or U22989 (N_22989,N_22159,N_22417);
and U22990 (N_22990,N_22010,N_22294);
nor U22991 (N_22991,N_22135,N_22035);
and U22992 (N_22992,N_22176,N_22261);
or U22993 (N_22993,N_22313,N_22008);
and U22994 (N_22994,N_22319,N_22317);
or U22995 (N_22995,N_22412,N_22159);
nand U22996 (N_22996,N_22495,N_22001);
nand U22997 (N_22997,N_22396,N_22185);
nor U22998 (N_22998,N_22152,N_22165);
nor U22999 (N_22999,N_22146,N_22384);
xnor U23000 (N_23000,N_22835,N_22741);
xor U23001 (N_23001,N_22828,N_22543);
and U23002 (N_23002,N_22604,N_22790);
nand U23003 (N_23003,N_22903,N_22786);
nor U23004 (N_23004,N_22698,N_22662);
or U23005 (N_23005,N_22976,N_22535);
nor U23006 (N_23006,N_22996,N_22570);
xor U23007 (N_23007,N_22717,N_22630);
xnor U23008 (N_23008,N_22655,N_22985);
and U23009 (N_23009,N_22772,N_22555);
xnor U23010 (N_23010,N_22988,N_22765);
or U23011 (N_23011,N_22727,N_22631);
and U23012 (N_23012,N_22573,N_22796);
or U23013 (N_23013,N_22978,N_22914);
nor U23014 (N_23014,N_22856,N_22928);
nor U23015 (N_23015,N_22874,N_22798);
and U23016 (N_23016,N_22971,N_22587);
nand U23017 (N_23017,N_22615,N_22878);
xnor U23018 (N_23018,N_22730,N_22819);
xor U23019 (N_23019,N_22745,N_22838);
or U23020 (N_23020,N_22840,N_22957);
xnor U23021 (N_23021,N_22868,N_22692);
nand U23022 (N_23022,N_22725,N_22912);
and U23023 (N_23023,N_22743,N_22847);
nand U23024 (N_23024,N_22667,N_22677);
or U23025 (N_23025,N_22933,N_22645);
nor U23026 (N_23026,N_22536,N_22787);
xnor U23027 (N_23027,N_22523,N_22955);
or U23028 (N_23028,N_22782,N_22949);
or U23029 (N_23029,N_22580,N_22751);
or U23030 (N_23030,N_22824,N_22591);
and U23031 (N_23031,N_22624,N_22520);
xnor U23032 (N_23032,N_22884,N_22674);
and U23033 (N_23033,N_22590,N_22811);
and U23034 (N_23034,N_22930,N_22939);
nand U23035 (N_23035,N_22609,N_22929);
and U23036 (N_23036,N_22636,N_22813);
and U23037 (N_23037,N_22877,N_22697);
nor U23038 (N_23038,N_22529,N_22888);
and U23039 (N_23039,N_22920,N_22778);
nand U23040 (N_23040,N_22719,N_22739);
xnor U23041 (N_23041,N_22632,N_22718);
and U23042 (N_23042,N_22937,N_22788);
nand U23043 (N_23043,N_22647,N_22983);
nor U23044 (N_23044,N_22818,N_22825);
or U23045 (N_23045,N_22800,N_22746);
and U23046 (N_23046,N_22538,N_22972);
or U23047 (N_23047,N_22525,N_22548);
nor U23048 (N_23048,N_22889,N_22980);
nor U23049 (N_23049,N_22807,N_22742);
xnor U23050 (N_23050,N_22732,N_22962);
or U23051 (N_23051,N_22561,N_22654);
or U23052 (N_23052,N_22705,N_22945);
nor U23053 (N_23053,N_22669,N_22668);
nor U23054 (N_23054,N_22764,N_22648);
and U23055 (N_23055,N_22622,N_22897);
nor U23056 (N_23056,N_22894,N_22670);
nand U23057 (N_23057,N_22552,N_22612);
or U23058 (N_23058,N_22777,N_22517);
nor U23059 (N_23059,N_22756,N_22507);
nor U23060 (N_23060,N_22595,N_22923);
and U23061 (N_23061,N_22758,N_22922);
and U23062 (N_23062,N_22994,N_22673);
nor U23063 (N_23063,N_22829,N_22752);
and U23064 (N_23064,N_22537,N_22814);
and U23065 (N_23065,N_22857,N_22848);
nand U23066 (N_23066,N_22559,N_22816);
xor U23067 (N_23067,N_22560,N_22986);
nand U23068 (N_23068,N_22872,N_22505);
and U23069 (N_23069,N_22841,N_22823);
nor U23070 (N_23070,N_22905,N_22975);
or U23071 (N_23071,N_22837,N_22880);
nand U23072 (N_23072,N_22613,N_22927);
xnor U23073 (N_23073,N_22860,N_22821);
or U23074 (N_23074,N_22633,N_22576);
nor U23075 (N_23075,N_22794,N_22852);
nand U23076 (N_23076,N_22618,N_22513);
and U23077 (N_23077,N_22990,N_22554);
and U23078 (N_23078,N_22919,N_22569);
and U23079 (N_23079,N_22736,N_22755);
nor U23080 (N_23080,N_22979,N_22726);
nand U23081 (N_23081,N_22558,N_22557);
nor U23082 (N_23082,N_22577,N_22998);
nand U23083 (N_23083,N_22760,N_22926);
nand U23084 (N_23084,N_22831,N_22873);
xnor U23085 (N_23085,N_22849,N_22999);
nand U23086 (N_23086,N_22676,N_22773);
and U23087 (N_23087,N_22581,N_22691);
nor U23088 (N_23088,N_22634,N_22651);
xor U23089 (N_23089,N_22614,N_22579);
nor U23090 (N_23090,N_22958,N_22592);
and U23091 (N_23091,N_22617,N_22562);
nor U23092 (N_23092,N_22938,N_22968);
xor U23093 (N_23093,N_22509,N_22583);
nor U23094 (N_23094,N_22605,N_22516);
nor U23095 (N_23095,N_22508,N_22723);
xnor U23096 (N_23096,N_22593,N_22503);
nor U23097 (N_23097,N_22995,N_22693);
or U23098 (N_23098,N_22977,N_22871);
nor U23099 (N_23099,N_22540,N_22992);
xnor U23100 (N_23100,N_22853,N_22709);
nor U23101 (N_23101,N_22900,N_22941);
nand U23102 (N_23102,N_22965,N_22792);
xnor U23103 (N_23103,N_22943,N_22515);
xor U23104 (N_23104,N_22738,N_22907);
xnor U23105 (N_23105,N_22839,N_22733);
or U23106 (N_23106,N_22685,N_22909);
and U23107 (N_23107,N_22704,N_22808);
nor U23108 (N_23108,N_22785,N_22597);
nor U23109 (N_23109,N_22951,N_22659);
or U23110 (N_23110,N_22594,N_22585);
xnor U23111 (N_23111,N_22640,N_22721);
nand U23112 (N_23112,N_22602,N_22834);
nor U23113 (N_23113,N_22571,N_22961);
and U23114 (N_23114,N_22924,N_22506);
xnor U23115 (N_23115,N_22642,N_22551);
nor U23116 (N_23116,N_22896,N_22722);
xor U23117 (N_23117,N_22521,N_22895);
and U23118 (N_23118,N_22740,N_22661);
xor U23119 (N_23119,N_22522,N_22601);
nand U23120 (N_23120,N_22997,N_22628);
or U23121 (N_23121,N_22854,N_22600);
nor U23122 (N_23122,N_22750,N_22963);
nor U23123 (N_23123,N_22544,N_22759);
or U23124 (N_23124,N_22916,N_22703);
nand U23125 (N_23125,N_22588,N_22675);
nand U23126 (N_23126,N_22899,N_22969);
nor U23127 (N_23127,N_22641,N_22932);
and U23128 (N_23128,N_22846,N_22556);
or U23129 (N_23129,N_22524,N_22812);
xor U23130 (N_23130,N_22716,N_22547);
nand U23131 (N_23131,N_22578,N_22616);
and U23132 (N_23132,N_22973,N_22830);
nand U23133 (N_23133,N_22610,N_22694);
or U23134 (N_23134,N_22644,N_22657);
or U23135 (N_23135,N_22574,N_22954);
xnor U23136 (N_23136,N_22665,N_22776);
xor U23137 (N_23137,N_22864,N_22925);
and U23138 (N_23138,N_22737,N_22510);
nand U23139 (N_23139,N_22518,N_22886);
xnor U23140 (N_23140,N_22946,N_22827);
or U23141 (N_23141,N_22714,N_22934);
or U23142 (N_23142,N_22833,N_22680);
nand U23143 (N_23143,N_22708,N_22883);
and U23144 (N_23144,N_22845,N_22959);
and U23145 (N_23145,N_22890,N_22806);
nand U23146 (N_23146,N_22982,N_22715);
nor U23147 (N_23147,N_22836,N_22964);
nor U23148 (N_23148,N_22635,N_22809);
or U23149 (N_23149,N_22991,N_22687);
nor U23150 (N_23150,N_22950,N_22851);
or U23151 (N_23151,N_22512,N_22541);
or U23152 (N_23152,N_22566,N_22862);
nor U23153 (N_23153,N_22568,N_22710);
nand U23154 (N_23154,N_22817,N_22876);
or U23155 (N_23155,N_22918,N_22936);
and U23156 (N_23156,N_22966,N_22519);
or U23157 (N_23157,N_22917,N_22867);
and U23158 (N_23158,N_22660,N_22658);
xor U23159 (N_23159,N_22713,N_22861);
or U23160 (N_23160,N_22863,N_22542);
or U23161 (N_23161,N_22643,N_22689);
nor U23162 (N_23162,N_22620,N_22621);
nor U23163 (N_23163,N_22935,N_22753);
xor U23164 (N_23164,N_22953,N_22974);
or U23165 (N_23165,N_22993,N_22511);
or U23166 (N_23166,N_22649,N_22902);
and U23167 (N_23167,N_22885,N_22904);
and U23168 (N_23168,N_22619,N_22567);
nor U23169 (N_23169,N_22754,N_22940);
nand U23170 (N_23170,N_22948,N_22584);
nor U23171 (N_23171,N_22695,N_22607);
and U23172 (N_23172,N_22688,N_22815);
nand U23173 (N_23173,N_22627,N_22598);
nand U23174 (N_23174,N_22820,N_22720);
or U23175 (N_23175,N_22711,N_22781);
or U23176 (N_23176,N_22784,N_22767);
xor U23177 (N_23177,N_22672,N_22801);
nor U23178 (N_23178,N_22623,N_22504);
nor U23179 (N_23179,N_22989,N_22563);
nor U23180 (N_23180,N_22500,N_22822);
xor U23181 (N_23181,N_22639,N_22682);
and U23182 (N_23182,N_22881,N_22882);
nand U23183 (N_23183,N_22684,N_22629);
nand U23184 (N_23184,N_22768,N_22763);
xor U23185 (N_23185,N_22599,N_22652);
xor U23186 (N_23186,N_22810,N_22761);
nor U23187 (N_23187,N_22748,N_22783);
xor U23188 (N_23188,N_22915,N_22690);
nor U23189 (N_23189,N_22791,N_22795);
and U23190 (N_23190,N_22656,N_22549);
nor U23191 (N_23191,N_22892,N_22606);
xnor U23192 (N_23192,N_22683,N_22901);
or U23193 (N_23193,N_22843,N_22960);
and U23194 (N_23194,N_22671,N_22911);
or U23195 (N_23195,N_22545,N_22766);
xnor U23196 (N_23196,N_22553,N_22603);
xor U23197 (N_23197,N_22678,N_22646);
xnor U23198 (N_23198,N_22701,N_22865);
or U23199 (N_23199,N_22700,N_22626);
xor U23200 (N_23200,N_22531,N_22707);
or U23201 (N_23201,N_22729,N_22744);
and U23202 (N_23202,N_22696,N_22799);
or U23203 (N_23203,N_22844,N_22893);
xnor U23204 (N_23204,N_22870,N_22611);
nand U23205 (N_23205,N_22769,N_22803);
and U23206 (N_23206,N_22910,N_22650);
xor U23207 (N_23207,N_22637,N_22526);
and U23208 (N_23208,N_22780,N_22842);
nor U23209 (N_23209,N_22805,N_22789);
nand U23210 (N_23210,N_22734,N_22731);
nor U23211 (N_23211,N_22898,N_22770);
or U23212 (N_23212,N_22797,N_22582);
and U23213 (N_23213,N_22762,N_22921);
and U23214 (N_23214,N_22906,N_22502);
or U23215 (N_23215,N_22596,N_22728);
and U23216 (N_23216,N_22984,N_22944);
and U23217 (N_23217,N_22565,N_22747);
or U23218 (N_23218,N_22706,N_22956);
nand U23219 (N_23219,N_22532,N_22850);
or U23220 (N_23220,N_22702,N_22501);
or U23221 (N_23221,N_22663,N_22681);
or U23222 (N_23222,N_22858,N_22987);
or U23223 (N_23223,N_22913,N_22981);
xnor U23224 (N_23224,N_22564,N_22931);
nor U23225 (N_23225,N_22528,N_22572);
xor U23226 (N_23226,N_22908,N_22589);
or U23227 (N_23227,N_22859,N_22712);
and U23228 (N_23228,N_22638,N_22832);
and U23229 (N_23229,N_22793,N_22546);
and U23230 (N_23230,N_22653,N_22550);
nor U23231 (N_23231,N_22774,N_22664);
or U23232 (N_23232,N_22887,N_22539);
nand U23233 (N_23233,N_22869,N_22608);
and U23234 (N_23234,N_22826,N_22527);
or U23235 (N_23235,N_22804,N_22699);
and U23236 (N_23236,N_22534,N_22952);
and U23237 (N_23237,N_22879,N_22875);
xnor U23238 (N_23238,N_22586,N_22891);
nand U23239 (N_23239,N_22575,N_22735);
and U23240 (N_23240,N_22866,N_22967);
nand U23241 (N_23241,N_22942,N_22749);
and U23242 (N_23242,N_22625,N_22970);
xor U23243 (N_23243,N_22802,N_22779);
nand U23244 (N_23244,N_22724,N_22771);
nand U23245 (N_23245,N_22947,N_22686);
nand U23246 (N_23246,N_22533,N_22679);
nand U23247 (N_23247,N_22855,N_22666);
xnor U23248 (N_23248,N_22530,N_22757);
xor U23249 (N_23249,N_22514,N_22775);
or U23250 (N_23250,N_22708,N_22825);
nand U23251 (N_23251,N_22502,N_22608);
nor U23252 (N_23252,N_22972,N_22753);
xor U23253 (N_23253,N_22624,N_22838);
nor U23254 (N_23254,N_22894,N_22802);
nor U23255 (N_23255,N_22571,N_22682);
xor U23256 (N_23256,N_22997,N_22817);
and U23257 (N_23257,N_22704,N_22659);
or U23258 (N_23258,N_22889,N_22739);
xnor U23259 (N_23259,N_22522,N_22680);
nor U23260 (N_23260,N_22927,N_22775);
or U23261 (N_23261,N_22994,N_22765);
xor U23262 (N_23262,N_22552,N_22933);
and U23263 (N_23263,N_22712,N_22803);
nor U23264 (N_23264,N_22682,N_22887);
or U23265 (N_23265,N_22905,N_22855);
nand U23266 (N_23266,N_22895,N_22778);
and U23267 (N_23267,N_22745,N_22501);
nor U23268 (N_23268,N_22638,N_22647);
nand U23269 (N_23269,N_22682,N_22623);
and U23270 (N_23270,N_22791,N_22605);
nand U23271 (N_23271,N_22646,N_22628);
and U23272 (N_23272,N_22556,N_22586);
nand U23273 (N_23273,N_22596,N_22821);
nand U23274 (N_23274,N_22678,N_22983);
nor U23275 (N_23275,N_22737,N_22548);
nor U23276 (N_23276,N_22849,N_22557);
nand U23277 (N_23277,N_22729,N_22514);
or U23278 (N_23278,N_22740,N_22814);
nor U23279 (N_23279,N_22528,N_22995);
nor U23280 (N_23280,N_22621,N_22776);
and U23281 (N_23281,N_22557,N_22627);
nor U23282 (N_23282,N_22995,N_22982);
nand U23283 (N_23283,N_22645,N_22555);
nand U23284 (N_23284,N_22921,N_22960);
xnor U23285 (N_23285,N_22568,N_22664);
and U23286 (N_23286,N_22701,N_22659);
or U23287 (N_23287,N_22955,N_22537);
nor U23288 (N_23288,N_22925,N_22824);
and U23289 (N_23289,N_22929,N_22850);
nand U23290 (N_23290,N_22878,N_22764);
nand U23291 (N_23291,N_22900,N_22619);
and U23292 (N_23292,N_22770,N_22761);
nand U23293 (N_23293,N_22546,N_22626);
nand U23294 (N_23294,N_22841,N_22595);
nor U23295 (N_23295,N_22843,N_22995);
nand U23296 (N_23296,N_22761,N_22842);
nor U23297 (N_23297,N_22941,N_22746);
or U23298 (N_23298,N_22702,N_22685);
nor U23299 (N_23299,N_22966,N_22647);
nand U23300 (N_23300,N_22894,N_22891);
and U23301 (N_23301,N_22640,N_22658);
xor U23302 (N_23302,N_22815,N_22603);
or U23303 (N_23303,N_22990,N_22968);
nand U23304 (N_23304,N_22982,N_22587);
nand U23305 (N_23305,N_22562,N_22734);
or U23306 (N_23306,N_22502,N_22799);
nor U23307 (N_23307,N_22952,N_22900);
or U23308 (N_23308,N_22702,N_22551);
xor U23309 (N_23309,N_22647,N_22893);
xnor U23310 (N_23310,N_22638,N_22912);
nand U23311 (N_23311,N_22977,N_22561);
nand U23312 (N_23312,N_22718,N_22943);
and U23313 (N_23313,N_22994,N_22990);
or U23314 (N_23314,N_22964,N_22912);
nand U23315 (N_23315,N_22970,N_22923);
and U23316 (N_23316,N_22544,N_22695);
xnor U23317 (N_23317,N_22503,N_22531);
or U23318 (N_23318,N_22653,N_22954);
nand U23319 (N_23319,N_22796,N_22583);
xnor U23320 (N_23320,N_22762,N_22686);
nand U23321 (N_23321,N_22591,N_22978);
or U23322 (N_23322,N_22863,N_22671);
nand U23323 (N_23323,N_22927,N_22668);
and U23324 (N_23324,N_22613,N_22799);
and U23325 (N_23325,N_22783,N_22553);
nand U23326 (N_23326,N_22756,N_22642);
xor U23327 (N_23327,N_22672,N_22910);
or U23328 (N_23328,N_22572,N_22906);
or U23329 (N_23329,N_22749,N_22860);
xor U23330 (N_23330,N_22623,N_22547);
nor U23331 (N_23331,N_22867,N_22971);
or U23332 (N_23332,N_22651,N_22718);
nand U23333 (N_23333,N_22736,N_22893);
nor U23334 (N_23334,N_22629,N_22549);
or U23335 (N_23335,N_22560,N_22760);
nor U23336 (N_23336,N_22623,N_22794);
nor U23337 (N_23337,N_22716,N_22753);
xor U23338 (N_23338,N_22947,N_22820);
xnor U23339 (N_23339,N_22688,N_22690);
and U23340 (N_23340,N_22516,N_22511);
nand U23341 (N_23341,N_22662,N_22771);
or U23342 (N_23342,N_22800,N_22778);
xor U23343 (N_23343,N_22649,N_22919);
nor U23344 (N_23344,N_22998,N_22930);
and U23345 (N_23345,N_22686,N_22813);
or U23346 (N_23346,N_22727,N_22779);
and U23347 (N_23347,N_22885,N_22882);
nor U23348 (N_23348,N_22977,N_22849);
and U23349 (N_23349,N_22516,N_22960);
nor U23350 (N_23350,N_22943,N_22982);
xnor U23351 (N_23351,N_22921,N_22918);
nor U23352 (N_23352,N_22528,N_22797);
and U23353 (N_23353,N_22549,N_22609);
or U23354 (N_23354,N_22846,N_22931);
nand U23355 (N_23355,N_22764,N_22739);
or U23356 (N_23356,N_22658,N_22709);
xnor U23357 (N_23357,N_22540,N_22743);
or U23358 (N_23358,N_22800,N_22741);
nor U23359 (N_23359,N_22942,N_22560);
nor U23360 (N_23360,N_22852,N_22640);
and U23361 (N_23361,N_22867,N_22855);
or U23362 (N_23362,N_22697,N_22682);
xnor U23363 (N_23363,N_22577,N_22985);
xnor U23364 (N_23364,N_22777,N_22917);
nand U23365 (N_23365,N_22824,N_22594);
or U23366 (N_23366,N_22747,N_22916);
nor U23367 (N_23367,N_22615,N_22632);
xor U23368 (N_23368,N_22679,N_22887);
or U23369 (N_23369,N_22960,N_22930);
or U23370 (N_23370,N_22851,N_22791);
nor U23371 (N_23371,N_22697,N_22629);
nand U23372 (N_23372,N_22976,N_22692);
and U23373 (N_23373,N_22896,N_22633);
xor U23374 (N_23374,N_22719,N_22888);
nor U23375 (N_23375,N_22502,N_22503);
and U23376 (N_23376,N_22620,N_22908);
nor U23377 (N_23377,N_22528,N_22958);
xnor U23378 (N_23378,N_22989,N_22715);
nand U23379 (N_23379,N_22583,N_22527);
nor U23380 (N_23380,N_22573,N_22583);
nor U23381 (N_23381,N_22687,N_22664);
xor U23382 (N_23382,N_22614,N_22538);
and U23383 (N_23383,N_22592,N_22940);
xnor U23384 (N_23384,N_22701,N_22756);
or U23385 (N_23385,N_22599,N_22788);
and U23386 (N_23386,N_22540,N_22837);
xor U23387 (N_23387,N_22818,N_22528);
nand U23388 (N_23388,N_22909,N_22555);
nor U23389 (N_23389,N_22561,N_22990);
and U23390 (N_23390,N_22948,N_22889);
or U23391 (N_23391,N_22585,N_22557);
nand U23392 (N_23392,N_22949,N_22997);
xor U23393 (N_23393,N_22646,N_22677);
or U23394 (N_23394,N_22913,N_22744);
xnor U23395 (N_23395,N_22826,N_22761);
xor U23396 (N_23396,N_22681,N_22934);
nor U23397 (N_23397,N_22629,N_22871);
and U23398 (N_23398,N_22531,N_22963);
and U23399 (N_23399,N_22917,N_22888);
xnor U23400 (N_23400,N_22780,N_22967);
or U23401 (N_23401,N_22653,N_22744);
nor U23402 (N_23402,N_22643,N_22842);
and U23403 (N_23403,N_22574,N_22678);
nor U23404 (N_23404,N_22995,N_22599);
nor U23405 (N_23405,N_22667,N_22988);
nor U23406 (N_23406,N_22618,N_22745);
nor U23407 (N_23407,N_22618,N_22935);
xor U23408 (N_23408,N_22617,N_22944);
xnor U23409 (N_23409,N_22512,N_22852);
nor U23410 (N_23410,N_22547,N_22925);
nor U23411 (N_23411,N_22802,N_22569);
or U23412 (N_23412,N_22802,N_22781);
xor U23413 (N_23413,N_22603,N_22698);
and U23414 (N_23414,N_22627,N_22680);
or U23415 (N_23415,N_22754,N_22613);
xor U23416 (N_23416,N_22552,N_22632);
or U23417 (N_23417,N_22550,N_22780);
nand U23418 (N_23418,N_22827,N_22683);
or U23419 (N_23419,N_22747,N_22740);
xnor U23420 (N_23420,N_22566,N_22883);
xnor U23421 (N_23421,N_22658,N_22882);
nand U23422 (N_23422,N_22909,N_22689);
and U23423 (N_23423,N_22517,N_22794);
nor U23424 (N_23424,N_22964,N_22501);
nor U23425 (N_23425,N_22869,N_22713);
or U23426 (N_23426,N_22688,N_22547);
xor U23427 (N_23427,N_22862,N_22637);
nand U23428 (N_23428,N_22957,N_22913);
or U23429 (N_23429,N_22968,N_22742);
xor U23430 (N_23430,N_22684,N_22696);
xnor U23431 (N_23431,N_22619,N_22754);
and U23432 (N_23432,N_22568,N_22875);
nand U23433 (N_23433,N_22629,N_22646);
nand U23434 (N_23434,N_22664,N_22599);
or U23435 (N_23435,N_22514,N_22791);
or U23436 (N_23436,N_22943,N_22539);
or U23437 (N_23437,N_22544,N_22929);
or U23438 (N_23438,N_22638,N_22518);
xnor U23439 (N_23439,N_22517,N_22915);
or U23440 (N_23440,N_22887,N_22844);
xnor U23441 (N_23441,N_22907,N_22939);
nand U23442 (N_23442,N_22835,N_22844);
or U23443 (N_23443,N_22636,N_22587);
nor U23444 (N_23444,N_22712,N_22851);
xor U23445 (N_23445,N_22873,N_22813);
xor U23446 (N_23446,N_22500,N_22810);
or U23447 (N_23447,N_22769,N_22798);
and U23448 (N_23448,N_22720,N_22980);
nand U23449 (N_23449,N_22663,N_22833);
nand U23450 (N_23450,N_22596,N_22875);
nand U23451 (N_23451,N_22996,N_22882);
nand U23452 (N_23452,N_22738,N_22785);
nand U23453 (N_23453,N_22708,N_22507);
or U23454 (N_23454,N_22972,N_22958);
nand U23455 (N_23455,N_22822,N_22741);
nand U23456 (N_23456,N_22543,N_22722);
and U23457 (N_23457,N_22530,N_22817);
or U23458 (N_23458,N_22640,N_22832);
xor U23459 (N_23459,N_22835,N_22786);
or U23460 (N_23460,N_22907,N_22917);
nor U23461 (N_23461,N_22845,N_22992);
xnor U23462 (N_23462,N_22881,N_22610);
or U23463 (N_23463,N_22975,N_22631);
nor U23464 (N_23464,N_22511,N_22895);
or U23465 (N_23465,N_22876,N_22836);
xor U23466 (N_23466,N_22622,N_22754);
nand U23467 (N_23467,N_22509,N_22628);
nor U23468 (N_23468,N_22566,N_22877);
xnor U23469 (N_23469,N_22916,N_22616);
xor U23470 (N_23470,N_22871,N_22776);
or U23471 (N_23471,N_22968,N_22988);
nor U23472 (N_23472,N_22890,N_22632);
nor U23473 (N_23473,N_22589,N_22591);
xor U23474 (N_23474,N_22715,N_22542);
or U23475 (N_23475,N_22754,N_22881);
nand U23476 (N_23476,N_22952,N_22932);
and U23477 (N_23477,N_22633,N_22532);
or U23478 (N_23478,N_22792,N_22777);
and U23479 (N_23479,N_22681,N_22686);
nor U23480 (N_23480,N_22768,N_22636);
or U23481 (N_23481,N_22597,N_22787);
nor U23482 (N_23482,N_22516,N_22924);
or U23483 (N_23483,N_22925,N_22520);
xnor U23484 (N_23484,N_22997,N_22670);
nor U23485 (N_23485,N_22789,N_22853);
xnor U23486 (N_23486,N_22998,N_22955);
nor U23487 (N_23487,N_22844,N_22649);
or U23488 (N_23488,N_22929,N_22529);
nor U23489 (N_23489,N_22580,N_22721);
nor U23490 (N_23490,N_22759,N_22552);
or U23491 (N_23491,N_22702,N_22789);
nand U23492 (N_23492,N_22940,N_22572);
nand U23493 (N_23493,N_22757,N_22911);
nand U23494 (N_23494,N_22962,N_22811);
and U23495 (N_23495,N_22689,N_22991);
nor U23496 (N_23496,N_22728,N_22959);
or U23497 (N_23497,N_22767,N_22558);
or U23498 (N_23498,N_22992,N_22909);
xor U23499 (N_23499,N_22991,N_22839);
nor U23500 (N_23500,N_23233,N_23121);
nor U23501 (N_23501,N_23170,N_23462);
nand U23502 (N_23502,N_23117,N_23421);
xnor U23503 (N_23503,N_23212,N_23153);
and U23504 (N_23504,N_23068,N_23495);
nor U23505 (N_23505,N_23210,N_23156);
and U23506 (N_23506,N_23418,N_23100);
and U23507 (N_23507,N_23040,N_23102);
and U23508 (N_23508,N_23087,N_23248);
nor U23509 (N_23509,N_23486,N_23055);
or U23510 (N_23510,N_23157,N_23174);
and U23511 (N_23511,N_23145,N_23026);
nand U23512 (N_23512,N_23084,N_23176);
nor U23513 (N_23513,N_23337,N_23038);
nor U23514 (N_23514,N_23478,N_23479);
nor U23515 (N_23515,N_23195,N_23315);
xnor U23516 (N_23516,N_23410,N_23065);
or U23517 (N_23517,N_23060,N_23280);
and U23518 (N_23518,N_23198,N_23439);
nor U23519 (N_23519,N_23096,N_23132);
nor U23520 (N_23520,N_23464,N_23034);
or U23521 (N_23521,N_23115,N_23049);
and U23522 (N_23522,N_23203,N_23357);
nor U23523 (N_23523,N_23420,N_23274);
or U23524 (N_23524,N_23028,N_23309);
or U23525 (N_23525,N_23159,N_23336);
xnor U23526 (N_23526,N_23445,N_23128);
nand U23527 (N_23527,N_23425,N_23191);
nor U23528 (N_23528,N_23139,N_23490);
or U23529 (N_23529,N_23154,N_23222);
nand U23530 (N_23530,N_23260,N_23291);
nand U23531 (N_23531,N_23067,N_23384);
and U23532 (N_23532,N_23392,N_23207);
nand U23533 (N_23533,N_23214,N_23349);
nand U23534 (N_23534,N_23369,N_23449);
nor U23535 (N_23535,N_23048,N_23390);
and U23536 (N_23536,N_23202,N_23404);
xnor U23537 (N_23537,N_23296,N_23124);
and U23538 (N_23538,N_23230,N_23411);
and U23539 (N_23539,N_23002,N_23211);
xnor U23540 (N_23540,N_23224,N_23467);
xor U23541 (N_23541,N_23360,N_23249);
nand U23542 (N_23542,N_23213,N_23167);
and U23543 (N_23543,N_23466,N_23489);
nor U23544 (N_23544,N_23456,N_23234);
nor U23545 (N_23545,N_23030,N_23304);
nor U23546 (N_23546,N_23039,N_23220);
nor U23547 (N_23547,N_23064,N_23162);
and U23548 (N_23548,N_23373,N_23245);
nor U23549 (N_23549,N_23081,N_23386);
or U23550 (N_23550,N_23221,N_23272);
nor U23551 (N_23551,N_23253,N_23423);
nor U23552 (N_23552,N_23085,N_23056);
xnor U23553 (N_23553,N_23165,N_23334);
nand U23554 (N_23554,N_23442,N_23459);
and U23555 (N_23555,N_23018,N_23118);
nor U23556 (N_23556,N_23152,N_23484);
or U23557 (N_23557,N_23453,N_23474);
or U23558 (N_23558,N_23239,N_23074);
xor U23559 (N_23559,N_23090,N_23393);
nor U23560 (N_23560,N_23427,N_23236);
xor U23561 (N_23561,N_23316,N_23023);
nand U23562 (N_23562,N_23440,N_23146);
xor U23563 (N_23563,N_23052,N_23497);
xnor U23564 (N_23564,N_23250,N_23340);
nand U23565 (N_23565,N_23168,N_23308);
nor U23566 (N_23566,N_23077,N_23394);
nor U23567 (N_23567,N_23235,N_23218);
or U23568 (N_23568,N_23299,N_23380);
nand U23569 (N_23569,N_23240,N_23092);
xnor U23570 (N_23570,N_23172,N_23348);
and U23571 (N_23571,N_23252,N_23494);
or U23572 (N_23572,N_23322,N_23182);
and U23573 (N_23573,N_23256,N_23244);
or U23574 (N_23574,N_23416,N_23109);
or U23575 (N_23575,N_23119,N_23492);
nor U23576 (N_23576,N_23382,N_23398);
xor U23577 (N_23577,N_23199,N_23258);
or U23578 (N_23578,N_23059,N_23350);
and U23579 (N_23579,N_23365,N_23454);
nor U23580 (N_23580,N_23103,N_23330);
nor U23581 (N_23581,N_23385,N_23073);
nand U23582 (N_23582,N_23407,N_23364);
nor U23583 (N_23583,N_23205,N_23080);
xor U23584 (N_23584,N_23187,N_23408);
nand U23585 (N_23585,N_23051,N_23447);
nand U23586 (N_23586,N_23430,N_23241);
nand U23587 (N_23587,N_23223,N_23284);
nor U23588 (N_23588,N_23282,N_23275);
nand U23589 (N_23589,N_23376,N_23201);
xnor U23590 (N_23590,N_23114,N_23397);
xor U23591 (N_23591,N_23032,N_23247);
xor U23592 (N_23592,N_23166,N_23290);
and U23593 (N_23593,N_23317,N_23004);
nand U23594 (N_23594,N_23149,N_23110);
xnor U23595 (N_23595,N_23475,N_23196);
or U23596 (N_23596,N_23089,N_23000);
or U23597 (N_23597,N_23129,N_23131);
or U23598 (N_23598,N_23457,N_23158);
xor U23599 (N_23599,N_23434,N_23400);
nor U23600 (N_23600,N_23151,N_23116);
or U23601 (N_23601,N_23413,N_23135);
and U23602 (N_23602,N_23070,N_23126);
nand U23603 (N_23603,N_23352,N_23257);
or U23604 (N_23604,N_23363,N_23231);
and U23605 (N_23605,N_23086,N_23343);
nand U23606 (N_23606,N_23452,N_23232);
or U23607 (N_23607,N_23262,N_23345);
nand U23608 (N_23608,N_23485,N_23079);
nand U23609 (N_23609,N_23431,N_23061);
and U23610 (N_23610,N_23259,N_23477);
and U23611 (N_23611,N_23078,N_23396);
xor U23612 (N_23612,N_23189,N_23058);
and U23613 (N_23613,N_23123,N_23424);
xor U23614 (N_23614,N_23142,N_23361);
xor U23615 (N_23615,N_23335,N_23325);
and U23616 (N_23616,N_23193,N_23375);
nand U23617 (N_23617,N_23009,N_23403);
xnor U23618 (N_23618,N_23406,N_23496);
nand U23619 (N_23619,N_23082,N_23044);
or U23620 (N_23620,N_23267,N_23066);
xnor U23621 (N_23621,N_23185,N_23379);
and U23622 (N_23622,N_23412,N_23285);
or U23623 (N_23623,N_23219,N_23371);
nand U23624 (N_23624,N_23083,N_23037);
xnor U23625 (N_23625,N_23057,N_23164);
nand U23626 (N_23626,N_23209,N_23399);
or U23627 (N_23627,N_23271,N_23300);
xor U23628 (N_23628,N_23053,N_23428);
or U23629 (N_23629,N_23306,N_23419);
nor U23630 (N_23630,N_23141,N_23091);
nor U23631 (N_23631,N_23472,N_23307);
and U23632 (N_23632,N_23264,N_23169);
nand U23633 (N_23633,N_23127,N_23329);
xor U23634 (N_23634,N_23362,N_23292);
nor U23635 (N_23635,N_23108,N_23188);
nor U23636 (N_23636,N_23217,N_23438);
or U23637 (N_23637,N_23075,N_23181);
nand U23638 (N_23638,N_23254,N_23225);
nand U23639 (N_23639,N_23206,N_23179);
and U23640 (N_23640,N_23338,N_23025);
and U23641 (N_23641,N_23273,N_23354);
nor U23642 (N_23642,N_23372,N_23093);
nor U23643 (N_23643,N_23033,N_23024);
xnor U23644 (N_23644,N_23279,N_23183);
xnor U23645 (N_23645,N_23005,N_23339);
nor U23646 (N_23646,N_23368,N_23483);
and U23647 (N_23647,N_23021,N_23328);
xnor U23648 (N_23648,N_23173,N_23289);
and U23649 (N_23649,N_23043,N_23331);
xor U23650 (N_23650,N_23358,N_23332);
nor U23651 (N_23651,N_23045,N_23041);
nand U23652 (N_23652,N_23022,N_23441);
or U23653 (N_23653,N_23318,N_23270);
or U23654 (N_23654,N_23113,N_23229);
or U23655 (N_23655,N_23194,N_23042);
nor U23656 (N_23656,N_23488,N_23122);
or U23657 (N_23657,N_23178,N_23106);
nand U23658 (N_23658,N_23161,N_23251);
or U23659 (N_23659,N_23098,N_23072);
or U23660 (N_23660,N_23293,N_23377);
xor U23661 (N_23661,N_23101,N_23163);
nand U23662 (N_23662,N_23095,N_23294);
nor U23663 (N_23663,N_23303,N_23498);
or U23664 (N_23664,N_23155,N_23414);
nor U23665 (N_23665,N_23437,N_23326);
nand U23666 (N_23666,N_23266,N_23402);
nor U23667 (N_23667,N_23197,N_23016);
nor U23668 (N_23668,N_23076,N_23277);
xor U23669 (N_23669,N_23237,N_23177);
xor U23670 (N_23670,N_23001,N_23006);
xor U23671 (N_23671,N_23134,N_23031);
xnor U23672 (N_23672,N_23295,N_23133);
nor U23673 (N_23673,N_23226,N_23227);
nand U23674 (N_23674,N_23346,N_23099);
or U23675 (N_23675,N_23367,N_23320);
nand U23676 (N_23676,N_23125,N_23344);
nand U23677 (N_23677,N_23341,N_23389);
and U23678 (N_23678,N_23036,N_23228);
and U23679 (N_23679,N_23480,N_23192);
and U23680 (N_23680,N_23017,N_23011);
nor U23681 (N_23681,N_23286,N_23138);
xnor U23682 (N_23682,N_23415,N_23324);
and U23683 (N_23683,N_23027,N_23265);
nand U23684 (N_23684,N_23062,N_23473);
nand U23685 (N_23685,N_23463,N_23120);
xor U23686 (N_23686,N_23409,N_23448);
nor U23687 (N_23687,N_23148,N_23417);
xnor U23688 (N_23688,N_23136,N_23255);
nand U23689 (N_23689,N_23276,N_23238);
and U23690 (N_23690,N_23029,N_23327);
nand U23691 (N_23691,N_23310,N_23374);
xor U23692 (N_23692,N_23493,N_23395);
or U23693 (N_23693,N_23471,N_23347);
or U23694 (N_23694,N_23481,N_23246);
nand U23695 (N_23695,N_23112,N_23469);
or U23696 (N_23696,N_23283,N_23460);
or U23697 (N_23697,N_23387,N_23104);
or U23698 (N_23698,N_23186,N_23150);
nand U23699 (N_23699,N_23137,N_23499);
nor U23700 (N_23700,N_23391,N_23401);
nand U23701 (N_23701,N_23140,N_23047);
nand U23702 (N_23702,N_23071,N_23147);
xnor U23703 (N_23703,N_23487,N_23455);
nand U23704 (N_23704,N_23429,N_23444);
nand U23705 (N_23705,N_23461,N_23007);
and U23706 (N_23706,N_23144,N_23008);
xnor U23707 (N_23707,N_23355,N_23215);
or U23708 (N_23708,N_23301,N_23171);
nor U23709 (N_23709,N_23190,N_23436);
or U23710 (N_23710,N_23383,N_23312);
nor U23711 (N_23711,N_23184,N_23451);
xnor U23712 (N_23712,N_23458,N_23366);
nor U23713 (N_23713,N_23450,N_23269);
nand U23714 (N_23714,N_23242,N_23014);
and U23715 (N_23715,N_23208,N_23470);
or U23716 (N_23716,N_23263,N_23356);
and U23717 (N_23717,N_23297,N_23314);
xor U23718 (N_23718,N_23054,N_23160);
or U23719 (N_23719,N_23063,N_23204);
or U23720 (N_23720,N_23313,N_23465);
or U23721 (N_23721,N_23287,N_23035);
nor U23722 (N_23722,N_23015,N_23143);
and U23723 (N_23723,N_23351,N_23046);
and U23724 (N_23724,N_23130,N_23012);
and U23725 (N_23725,N_23426,N_23180);
nand U23726 (N_23726,N_23288,N_23050);
nand U23727 (N_23727,N_23278,N_23261);
xor U23728 (N_23728,N_23491,N_23305);
nor U23729 (N_23729,N_23020,N_23370);
xnor U23730 (N_23730,N_23476,N_23433);
and U23731 (N_23731,N_23281,N_23422);
and U23732 (N_23732,N_23200,N_23107);
nor U23733 (N_23733,N_23432,N_23388);
xor U23734 (N_23734,N_23302,N_23435);
and U23735 (N_23735,N_23405,N_23468);
xnor U23736 (N_23736,N_23446,N_23443);
and U23737 (N_23737,N_23069,N_23097);
xor U23738 (N_23738,N_23482,N_23321);
and U23739 (N_23739,N_23342,N_23019);
and U23740 (N_23740,N_23359,N_23243);
xnor U23741 (N_23741,N_23013,N_23088);
nand U23742 (N_23742,N_23311,N_23378);
nand U23743 (N_23743,N_23111,N_23319);
xnor U23744 (N_23744,N_23381,N_23216);
and U23745 (N_23745,N_23105,N_23175);
xor U23746 (N_23746,N_23003,N_23268);
or U23747 (N_23747,N_23298,N_23010);
nand U23748 (N_23748,N_23353,N_23094);
xnor U23749 (N_23749,N_23333,N_23323);
nand U23750 (N_23750,N_23332,N_23279);
or U23751 (N_23751,N_23354,N_23498);
or U23752 (N_23752,N_23099,N_23483);
or U23753 (N_23753,N_23122,N_23425);
and U23754 (N_23754,N_23194,N_23211);
nand U23755 (N_23755,N_23342,N_23163);
xnor U23756 (N_23756,N_23108,N_23033);
nor U23757 (N_23757,N_23213,N_23269);
nor U23758 (N_23758,N_23193,N_23497);
nand U23759 (N_23759,N_23240,N_23175);
and U23760 (N_23760,N_23406,N_23106);
xnor U23761 (N_23761,N_23308,N_23236);
nand U23762 (N_23762,N_23078,N_23446);
or U23763 (N_23763,N_23304,N_23057);
nor U23764 (N_23764,N_23291,N_23405);
or U23765 (N_23765,N_23012,N_23109);
xor U23766 (N_23766,N_23156,N_23257);
and U23767 (N_23767,N_23483,N_23460);
or U23768 (N_23768,N_23226,N_23355);
nor U23769 (N_23769,N_23298,N_23277);
nor U23770 (N_23770,N_23210,N_23144);
xnor U23771 (N_23771,N_23118,N_23355);
nand U23772 (N_23772,N_23250,N_23348);
or U23773 (N_23773,N_23128,N_23049);
or U23774 (N_23774,N_23032,N_23310);
or U23775 (N_23775,N_23224,N_23451);
nor U23776 (N_23776,N_23423,N_23031);
or U23777 (N_23777,N_23010,N_23467);
or U23778 (N_23778,N_23314,N_23444);
and U23779 (N_23779,N_23058,N_23308);
nand U23780 (N_23780,N_23187,N_23322);
xnor U23781 (N_23781,N_23383,N_23355);
xor U23782 (N_23782,N_23364,N_23326);
nor U23783 (N_23783,N_23317,N_23101);
xor U23784 (N_23784,N_23242,N_23400);
nor U23785 (N_23785,N_23067,N_23445);
nor U23786 (N_23786,N_23312,N_23359);
xor U23787 (N_23787,N_23306,N_23089);
nor U23788 (N_23788,N_23139,N_23091);
nor U23789 (N_23789,N_23271,N_23127);
nand U23790 (N_23790,N_23196,N_23076);
and U23791 (N_23791,N_23375,N_23376);
or U23792 (N_23792,N_23315,N_23427);
and U23793 (N_23793,N_23349,N_23343);
or U23794 (N_23794,N_23454,N_23328);
and U23795 (N_23795,N_23159,N_23422);
xor U23796 (N_23796,N_23339,N_23407);
nor U23797 (N_23797,N_23263,N_23300);
nand U23798 (N_23798,N_23275,N_23413);
or U23799 (N_23799,N_23377,N_23301);
or U23800 (N_23800,N_23075,N_23440);
or U23801 (N_23801,N_23342,N_23234);
nand U23802 (N_23802,N_23366,N_23168);
nor U23803 (N_23803,N_23227,N_23497);
or U23804 (N_23804,N_23283,N_23341);
xor U23805 (N_23805,N_23026,N_23182);
nand U23806 (N_23806,N_23295,N_23233);
and U23807 (N_23807,N_23112,N_23419);
xnor U23808 (N_23808,N_23106,N_23088);
xnor U23809 (N_23809,N_23490,N_23414);
nand U23810 (N_23810,N_23197,N_23065);
or U23811 (N_23811,N_23357,N_23303);
xor U23812 (N_23812,N_23048,N_23158);
and U23813 (N_23813,N_23269,N_23178);
nor U23814 (N_23814,N_23224,N_23106);
xnor U23815 (N_23815,N_23028,N_23270);
xor U23816 (N_23816,N_23362,N_23326);
nor U23817 (N_23817,N_23463,N_23237);
nand U23818 (N_23818,N_23440,N_23044);
and U23819 (N_23819,N_23461,N_23142);
xor U23820 (N_23820,N_23482,N_23276);
xor U23821 (N_23821,N_23284,N_23208);
nand U23822 (N_23822,N_23063,N_23403);
nand U23823 (N_23823,N_23435,N_23262);
nand U23824 (N_23824,N_23398,N_23268);
nor U23825 (N_23825,N_23030,N_23338);
and U23826 (N_23826,N_23252,N_23354);
or U23827 (N_23827,N_23201,N_23314);
nor U23828 (N_23828,N_23202,N_23401);
or U23829 (N_23829,N_23252,N_23232);
and U23830 (N_23830,N_23195,N_23199);
and U23831 (N_23831,N_23436,N_23415);
xnor U23832 (N_23832,N_23243,N_23066);
nor U23833 (N_23833,N_23453,N_23023);
nand U23834 (N_23834,N_23136,N_23181);
nand U23835 (N_23835,N_23137,N_23446);
and U23836 (N_23836,N_23433,N_23456);
or U23837 (N_23837,N_23304,N_23121);
nor U23838 (N_23838,N_23449,N_23249);
xor U23839 (N_23839,N_23208,N_23370);
xor U23840 (N_23840,N_23083,N_23366);
and U23841 (N_23841,N_23074,N_23231);
nor U23842 (N_23842,N_23269,N_23165);
xnor U23843 (N_23843,N_23282,N_23307);
xnor U23844 (N_23844,N_23420,N_23100);
nor U23845 (N_23845,N_23363,N_23086);
nand U23846 (N_23846,N_23032,N_23437);
nor U23847 (N_23847,N_23189,N_23104);
nand U23848 (N_23848,N_23072,N_23196);
xnor U23849 (N_23849,N_23083,N_23129);
or U23850 (N_23850,N_23419,N_23197);
xnor U23851 (N_23851,N_23256,N_23000);
nor U23852 (N_23852,N_23391,N_23390);
or U23853 (N_23853,N_23107,N_23210);
xnor U23854 (N_23854,N_23411,N_23253);
or U23855 (N_23855,N_23350,N_23300);
nor U23856 (N_23856,N_23099,N_23227);
nand U23857 (N_23857,N_23225,N_23147);
or U23858 (N_23858,N_23001,N_23242);
or U23859 (N_23859,N_23493,N_23087);
nand U23860 (N_23860,N_23322,N_23358);
xor U23861 (N_23861,N_23210,N_23495);
xor U23862 (N_23862,N_23069,N_23338);
nand U23863 (N_23863,N_23059,N_23468);
or U23864 (N_23864,N_23335,N_23187);
nand U23865 (N_23865,N_23450,N_23003);
xor U23866 (N_23866,N_23342,N_23143);
nand U23867 (N_23867,N_23497,N_23120);
nor U23868 (N_23868,N_23331,N_23068);
or U23869 (N_23869,N_23103,N_23485);
nor U23870 (N_23870,N_23424,N_23044);
or U23871 (N_23871,N_23141,N_23095);
xnor U23872 (N_23872,N_23344,N_23145);
nand U23873 (N_23873,N_23048,N_23278);
xor U23874 (N_23874,N_23067,N_23438);
or U23875 (N_23875,N_23063,N_23385);
and U23876 (N_23876,N_23406,N_23389);
or U23877 (N_23877,N_23378,N_23331);
and U23878 (N_23878,N_23326,N_23360);
nand U23879 (N_23879,N_23376,N_23045);
and U23880 (N_23880,N_23002,N_23080);
and U23881 (N_23881,N_23408,N_23209);
nor U23882 (N_23882,N_23403,N_23012);
or U23883 (N_23883,N_23046,N_23394);
and U23884 (N_23884,N_23440,N_23357);
nand U23885 (N_23885,N_23168,N_23202);
nor U23886 (N_23886,N_23367,N_23250);
nor U23887 (N_23887,N_23060,N_23085);
nand U23888 (N_23888,N_23097,N_23117);
xor U23889 (N_23889,N_23215,N_23067);
nor U23890 (N_23890,N_23220,N_23284);
or U23891 (N_23891,N_23081,N_23404);
and U23892 (N_23892,N_23001,N_23201);
or U23893 (N_23893,N_23049,N_23216);
and U23894 (N_23894,N_23020,N_23064);
and U23895 (N_23895,N_23346,N_23356);
or U23896 (N_23896,N_23385,N_23206);
or U23897 (N_23897,N_23345,N_23496);
xor U23898 (N_23898,N_23062,N_23245);
or U23899 (N_23899,N_23042,N_23327);
nor U23900 (N_23900,N_23494,N_23467);
xnor U23901 (N_23901,N_23150,N_23363);
xor U23902 (N_23902,N_23407,N_23133);
or U23903 (N_23903,N_23245,N_23351);
and U23904 (N_23904,N_23433,N_23247);
xor U23905 (N_23905,N_23041,N_23149);
xnor U23906 (N_23906,N_23470,N_23155);
and U23907 (N_23907,N_23042,N_23110);
and U23908 (N_23908,N_23162,N_23288);
xor U23909 (N_23909,N_23289,N_23316);
xnor U23910 (N_23910,N_23156,N_23335);
xor U23911 (N_23911,N_23185,N_23157);
nor U23912 (N_23912,N_23035,N_23239);
nor U23913 (N_23913,N_23290,N_23307);
nand U23914 (N_23914,N_23496,N_23450);
and U23915 (N_23915,N_23430,N_23498);
or U23916 (N_23916,N_23304,N_23411);
or U23917 (N_23917,N_23433,N_23029);
nand U23918 (N_23918,N_23159,N_23455);
xnor U23919 (N_23919,N_23100,N_23389);
xnor U23920 (N_23920,N_23018,N_23014);
or U23921 (N_23921,N_23261,N_23390);
or U23922 (N_23922,N_23462,N_23360);
or U23923 (N_23923,N_23017,N_23161);
or U23924 (N_23924,N_23250,N_23128);
or U23925 (N_23925,N_23451,N_23234);
and U23926 (N_23926,N_23439,N_23411);
xor U23927 (N_23927,N_23364,N_23454);
and U23928 (N_23928,N_23141,N_23105);
or U23929 (N_23929,N_23033,N_23232);
or U23930 (N_23930,N_23356,N_23216);
nor U23931 (N_23931,N_23310,N_23059);
nor U23932 (N_23932,N_23242,N_23025);
xnor U23933 (N_23933,N_23328,N_23182);
nor U23934 (N_23934,N_23438,N_23346);
and U23935 (N_23935,N_23235,N_23175);
xor U23936 (N_23936,N_23118,N_23074);
nor U23937 (N_23937,N_23042,N_23389);
or U23938 (N_23938,N_23321,N_23499);
nor U23939 (N_23939,N_23346,N_23304);
nor U23940 (N_23940,N_23297,N_23119);
or U23941 (N_23941,N_23387,N_23177);
or U23942 (N_23942,N_23467,N_23404);
or U23943 (N_23943,N_23021,N_23434);
or U23944 (N_23944,N_23381,N_23408);
or U23945 (N_23945,N_23404,N_23093);
xor U23946 (N_23946,N_23000,N_23301);
and U23947 (N_23947,N_23015,N_23073);
nand U23948 (N_23948,N_23497,N_23421);
nor U23949 (N_23949,N_23456,N_23483);
or U23950 (N_23950,N_23313,N_23482);
and U23951 (N_23951,N_23452,N_23387);
or U23952 (N_23952,N_23283,N_23251);
nor U23953 (N_23953,N_23477,N_23076);
nor U23954 (N_23954,N_23038,N_23087);
xor U23955 (N_23955,N_23024,N_23482);
xor U23956 (N_23956,N_23138,N_23130);
or U23957 (N_23957,N_23343,N_23434);
nor U23958 (N_23958,N_23328,N_23114);
or U23959 (N_23959,N_23491,N_23308);
nand U23960 (N_23960,N_23229,N_23211);
nor U23961 (N_23961,N_23217,N_23483);
nand U23962 (N_23962,N_23252,N_23152);
xor U23963 (N_23963,N_23036,N_23288);
and U23964 (N_23964,N_23376,N_23252);
nand U23965 (N_23965,N_23310,N_23270);
nor U23966 (N_23966,N_23450,N_23253);
xnor U23967 (N_23967,N_23432,N_23123);
and U23968 (N_23968,N_23196,N_23439);
and U23969 (N_23969,N_23293,N_23397);
xor U23970 (N_23970,N_23065,N_23250);
and U23971 (N_23971,N_23344,N_23290);
xnor U23972 (N_23972,N_23287,N_23029);
nand U23973 (N_23973,N_23036,N_23468);
xnor U23974 (N_23974,N_23374,N_23233);
nand U23975 (N_23975,N_23077,N_23311);
and U23976 (N_23976,N_23424,N_23031);
nor U23977 (N_23977,N_23137,N_23012);
nand U23978 (N_23978,N_23352,N_23292);
xnor U23979 (N_23979,N_23428,N_23276);
nor U23980 (N_23980,N_23468,N_23320);
and U23981 (N_23981,N_23273,N_23289);
xnor U23982 (N_23982,N_23047,N_23006);
and U23983 (N_23983,N_23234,N_23024);
nor U23984 (N_23984,N_23348,N_23018);
and U23985 (N_23985,N_23098,N_23410);
or U23986 (N_23986,N_23237,N_23419);
and U23987 (N_23987,N_23446,N_23432);
or U23988 (N_23988,N_23179,N_23135);
and U23989 (N_23989,N_23152,N_23116);
or U23990 (N_23990,N_23069,N_23253);
nor U23991 (N_23991,N_23308,N_23335);
or U23992 (N_23992,N_23067,N_23226);
xnor U23993 (N_23993,N_23111,N_23376);
xnor U23994 (N_23994,N_23457,N_23288);
nand U23995 (N_23995,N_23310,N_23056);
nor U23996 (N_23996,N_23369,N_23297);
and U23997 (N_23997,N_23009,N_23284);
and U23998 (N_23998,N_23437,N_23103);
and U23999 (N_23999,N_23293,N_23095);
xor U24000 (N_24000,N_23772,N_23681);
xor U24001 (N_24001,N_23859,N_23792);
and U24002 (N_24002,N_23846,N_23694);
and U24003 (N_24003,N_23755,N_23515);
or U24004 (N_24004,N_23973,N_23750);
and U24005 (N_24005,N_23672,N_23726);
or U24006 (N_24006,N_23967,N_23976);
nand U24007 (N_24007,N_23702,N_23985);
xnor U24008 (N_24008,N_23524,N_23791);
nor U24009 (N_24009,N_23674,N_23910);
and U24010 (N_24010,N_23598,N_23829);
xnor U24011 (N_24011,N_23686,N_23748);
xor U24012 (N_24012,N_23966,N_23535);
or U24013 (N_24013,N_23532,N_23586);
nand U24014 (N_24014,N_23899,N_23502);
and U24015 (N_24015,N_23897,N_23774);
xor U24016 (N_24016,N_23991,N_23602);
or U24017 (N_24017,N_23522,N_23877);
and U24018 (N_24018,N_23962,N_23545);
nand U24019 (N_24019,N_23907,N_23731);
xnor U24020 (N_24020,N_23560,N_23990);
nor U24021 (N_24021,N_23787,N_23730);
nor U24022 (N_24022,N_23604,N_23823);
and U24023 (N_24023,N_23749,N_23824);
and U24024 (N_24024,N_23510,N_23504);
and U24025 (N_24025,N_23762,N_23743);
xor U24026 (N_24026,N_23878,N_23646);
xor U24027 (N_24027,N_23876,N_23756);
nor U24028 (N_24028,N_23941,N_23732);
nand U24029 (N_24029,N_23719,N_23570);
nor U24030 (N_24030,N_23572,N_23815);
nor U24031 (N_24031,N_23668,N_23553);
or U24032 (N_24032,N_23869,N_23884);
or U24033 (N_24033,N_23549,N_23698);
xnor U24034 (N_24034,N_23905,N_23630);
and U24035 (N_24035,N_23875,N_23605);
nor U24036 (N_24036,N_23800,N_23600);
or U24037 (N_24037,N_23595,N_23541);
nor U24038 (N_24038,N_23701,N_23561);
nor U24039 (N_24039,N_23710,N_23663);
nor U24040 (N_24040,N_23953,N_23937);
xnor U24041 (N_24041,N_23757,N_23925);
nor U24042 (N_24042,N_23518,N_23709);
and U24043 (N_24043,N_23921,N_23758);
or U24044 (N_24044,N_23667,N_23608);
xnor U24045 (N_24045,N_23814,N_23989);
nand U24046 (N_24046,N_23920,N_23769);
and U24047 (N_24047,N_23851,N_23759);
nor U24048 (N_24048,N_23995,N_23754);
xnor U24049 (N_24049,N_23554,N_23746);
nor U24050 (N_24050,N_23854,N_23507);
and U24051 (N_24051,N_23635,N_23705);
or U24052 (N_24052,N_23901,N_23728);
nand U24053 (N_24053,N_23652,N_23874);
or U24054 (N_24054,N_23948,N_23569);
or U24055 (N_24055,N_23813,N_23785);
xor U24056 (N_24056,N_23676,N_23588);
xnor U24057 (N_24057,N_23795,N_23853);
and U24058 (N_24058,N_23651,N_23960);
nand U24059 (N_24059,N_23850,N_23512);
or U24060 (N_24060,N_23655,N_23678);
and U24061 (N_24061,N_23537,N_23793);
or U24062 (N_24062,N_23831,N_23776);
nor U24063 (N_24063,N_23856,N_23890);
nand U24064 (N_24064,N_23665,N_23514);
and U24065 (N_24065,N_23519,N_23885);
xnor U24066 (N_24066,N_23645,N_23855);
or U24067 (N_24067,N_23913,N_23817);
or U24068 (N_24068,N_23611,N_23596);
nor U24069 (N_24069,N_23888,N_23993);
and U24070 (N_24070,N_23734,N_23530);
nand U24071 (N_24071,N_23697,N_23898);
and U24072 (N_24072,N_23741,N_23503);
nor U24073 (N_24073,N_23879,N_23805);
or U24074 (N_24074,N_23808,N_23559);
xor U24075 (N_24075,N_23650,N_23609);
xnor U24076 (N_24076,N_23896,N_23615);
xor U24077 (N_24077,N_23523,N_23725);
nand U24078 (N_24078,N_23685,N_23603);
nor U24079 (N_24079,N_23675,N_23871);
nor U24080 (N_24080,N_23834,N_23919);
nor U24081 (N_24081,N_23822,N_23575);
xnor U24082 (N_24082,N_23547,N_23689);
and U24083 (N_24083,N_23752,N_23724);
and U24084 (N_24084,N_23648,N_23939);
nor U24085 (N_24085,N_23556,N_23627);
nand U24086 (N_24086,N_23927,N_23544);
nand U24087 (N_24087,N_23527,N_23526);
nand U24088 (N_24088,N_23924,N_23696);
or U24089 (N_24089,N_23505,N_23566);
nor U24090 (N_24090,N_23971,N_23688);
nand U24091 (N_24091,N_23912,N_23857);
nand U24092 (N_24092,N_23640,N_23649);
nor U24093 (N_24093,N_23770,N_23657);
nand U24094 (N_24094,N_23908,N_23677);
or U24095 (N_24095,N_23789,N_23836);
xor U24096 (N_24096,N_23811,N_23914);
and U24097 (N_24097,N_23521,N_23695);
xor U24098 (N_24098,N_23830,N_23771);
nand U24099 (N_24099,N_23832,N_23543);
and U24100 (N_24100,N_23825,N_23906);
xnor U24101 (N_24101,N_23969,N_23622);
nand U24102 (N_24102,N_23552,N_23629);
nor U24103 (N_24103,N_23916,N_23911);
nand U24104 (N_24104,N_23614,N_23781);
nor U24105 (N_24105,N_23712,N_23928);
nand U24106 (N_24106,N_23606,N_23849);
and U24107 (N_24107,N_23716,N_23509);
nand U24108 (N_24108,N_23639,N_23722);
xor U24109 (N_24109,N_23740,N_23634);
and U24110 (N_24110,N_23958,N_23607);
nand U24111 (N_24111,N_23867,N_23893);
nand U24112 (N_24112,N_23964,N_23567);
or U24113 (N_24113,N_23729,N_23986);
nand U24114 (N_24114,N_23520,N_23571);
and U24115 (N_24115,N_23858,N_23508);
nand U24116 (N_24116,N_23506,N_23786);
and U24117 (N_24117,N_23816,N_23778);
nand U24118 (N_24118,N_23718,N_23643);
or U24119 (N_24119,N_23558,N_23880);
nor U24120 (N_24120,N_23513,N_23972);
nand U24121 (N_24121,N_23847,N_23660);
xor U24122 (N_24122,N_23943,N_23982);
and U24123 (N_24123,N_23947,N_23766);
nand U24124 (N_24124,N_23700,N_23577);
xnor U24125 (N_24125,N_23801,N_23818);
or U24126 (N_24126,N_23938,N_23592);
nand U24127 (N_24127,N_23994,N_23782);
nor U24128 (N_24128,N_23804,N_23803);
and U24129 (N_24129,N_23654,N_23659);
or U24130 (N_24130,N_23579,N_23866);
or U24131 (N_24131,N_23717,N_23926);
and U24132 (N_24132,N_23624,N_23810);
and U24133 (N_24133,N_23662,N_23690);
and U24134 (N_24134,N_23658,N_23670);
nor U24135 (N_24135,N_23861,N_23979);
or U24136 (N_24136,N_23955,N_23961);
or U24137 (N_24137,N_23839,N_23929);
nand U24138 (N_24138,N_23739,N_23863);
or U24139 (N_24139,N_23599,N_23934);
or U24140 (N_24140,N_23583,N_23721);
or U24141 (N_24141,N_23631,N_23628);
or U24142 (N_24142,N_23687,N_23872);
or U24143 (N_24143,N_23841,N_23796);
nand U24144 (N_24144,N_23852,N_23983);
nand U24145 (N_24145,N_23568,N_23642);
xor U24146 (N_24146,N_23843,N_23711);
nor U24147 (N_24147,N_23768,N_23669);
xnor U24148 (N_24148,N_23998,N_23761);
nand U24149 (N_24149,N_23915,N_23744);
and U24150 (N_24150,N_23773,N_23827);
and U24151 (N_24151,N_23632,N_23970);
nand U24152 (N_24152,N_23533,N_23984);
and U24153 (N_24153,N_23809,N_23661);
and U24154 (N_24154,N_23623,N_23620);
xnor U24155 (N_24155,N_23974,N_23963);
nor U24156 (N_24156,N_23565,N_23935);
xor U24157 (N_24157,N_23587,N_23715);
nor U24158 (N_24158,N_23723,N_23840);
or U24159 (N_24159,N_23922,N_23584);
nand U24160 (N_24160,N_23633,N_23992);
xnor U24161 (N_24161,N_23653,N_23531);
nand U24162 (N_24162,N_23977,N_23736);
nand U24163 (N_24163,N_23904,N_23555);
nand U24164 (N_24164,N_23594,N_23673);
nor U24165 (N_24165,N_23644,N_23968);
nor U24166 (N_24166,N_23838,N_23763);
nand U24167 (N_24167,N_23807,N_23954);
nand U24168 (N_24168,N_23574,N_23613);
nor U24169 (N_24169,N_23589,N_23638);
and U24170 (N_24170,N_23767,N_23868);
nand U24171 (N_24171,N_23957,N_23610);
xor U24172 (N_24172,N_23656,N_23597);
xor U24173 (N_24173,N_23889,N_23933);
xnor U24174 (N_24174,N_23738,N_23917);
nor U24175 (N_24175,N_23704,N_23618);
nand U24176 (N_24176,N_23747,N_23797);
nor U24177 (N_24177,N_23517,N_23946);
and U24178 (N_24178,N_23636,N_23548);
and U24179 (N_24179,N_23842,N_23525);
and U24180 (N_24180,N_23802,N_23798);
nand U24181 (N_24181,N_23788,N_23720);
or U24182 (N_24182,N_23625,N_23996);
xnor U24183 (N_24183,N_23637,N_23784);
nor U24184 (N_24184,N_23956,N_23591);
xnor U24185 (N_24185,N_23923,N_23894);
nand U24186 (N_24186,N_23981,N_23987);
nand U24187 (N_24187,N_23909,N_23865);
nand U24188 (N_24188,N_23682,N_23593);
and U24189 (N_24189,N_23882,N_23619);
xor U24190 (N_24190,N_23581,N_23978);
or U24191 (N_24191,N_23783,N_23563);
xnor U24192 (N_24192,N_23745,N_23980);
and U24193 (N_24193,N_23936,N_23918);
xor U24194 (N_24194,N_23886,N_23988);
and U24195 (N_24195,N_23848,N_23580);
or U24196 (N_24196,N_23806,N_23501);
xnor U24197 (N_24197,N_23903,N_23799);
nand U24198 (N_24198,N_23870,N_23887);
and U24199 (N_24199,N_23952,N_23551);
xor U24200 (N_24200,N_23965,N_23837);
and U24201 (N_24201,N_23737,N_23542);
or U24202 (N_24202,N_23683,N_23895);
or U24203 (N_24203,N_23536,N_23641);
nand U24204 (N_24204,N_23699,N_23621);
or U24205 (N_24205,N_23949,N_23902);
nor U24206 (N_24206,N_23828,N_23573);
or U24207 (N_24207,N_23873,N_23820);
nor U24208 (N_24208,N_23706,N_23835);
xnor U24209 (N_24209,N_23692,N_23647);
xor U24210 (N_24210,N_23760,N_23585);
nand U24211 (N_24211,N_23578,N_23564);
and U24212 (N_24212,N_23626,N_23777);
nand U24213 (N_24213,N_23950,N_23945);
or U24214 (N_24214,N_23844,N_23534);
nor U24215 (N_24215,N_23664,N_23826);
nor U24216 (N_24216,N_23751,N_23765);
nor U24217 (N_24217,N_23550,N_23680);
nor U24218 (N_24218,N_23612,N_23516);
or U24219 (N_24219,N_23576,N_23819);
nor U24220 (N_24220,N_23693,N_23691);
nand U24221 (N_24221,N_23864,N_23959);
nor U24222 (N_24222,N_23708,N_23511);
nor U24223 (N_24223,N_23900,N_23779);
nor U24224 (N_24224,N_23742,N_23821);
or U24225 (N_24225,N_23940,N_23713);
nor U24226 (N_24226,N_23733,N_23529);
xnor U24227 (N_24227,N_23833,N_23735);
nand U24228 (N_24228,N_23727,N_23951);
xnor U24229 (N_24229,N_23679,N_23942);
or U24230 (N_24230,N_23891,N_23975);
nor U24231 (N_24231,N_23997,N_23539);
xnor U24232 (N_24232,N_23794,N_23703);
or U24233 (N_24233,N_23500,N_23790);
and U24234 (N_24234,N_23764,N_23707);
nand U24235 (N_24235,N_23562,N_23546);
and U24236 (N_24236,N_23617,N_23528);
nor U24237 (N_24237,N_23862,N_23753);
xor U24238 (N_24238,N_23601,N_23931);
nand U24239 (N_24239,N_23557,N_23860);
nor U24240 (N_24240,N_23930,N_23881);
nand U24241 (N_24241,N_23775,N_23944);
and U24242 (N_24242,N_23684,N_23932);
and U24243 (N_24243,N_23671,N_23883);
nand U24244 (N_24244,N_23616,N_23590);
or U24245 (N_24245,N_23538,N_23845);
nor U24246 (N_24246,N_23540,N_23812);
xnor U24247 (N_24247,N_23892,N_23714);
nand U24248 (N_24248,N_23999,N_23780);
nor U24249 (N_24249,N_23666,N_23582);
and U24250 (N_24250,N_23611,N_23939);
nor U24251 (N_24251,N_23823,N_23858);
nand U24252 (N_24252,N_23810,N_23866);
and U24253 (N_24253,N_23574,N_23717);
nand U24254 (N_24254,N_23545,N_23634);
xnor U24255 (N_24255,N_23678,N_23813);
nor U24256 (N_24256,N_23811,N_23526);
and U24257 (N_24257,N_23780,N_23734);
or U24258 (N_24258,N_23981,N_23563);
and U24259 (N_24259,N_23607,N_23964);
nand U24260 (N_24260,N_23856,N_23777);
nor U24261 (N_24261,N_23864,N_23609);
and U24262 (N_24262,N_23506,N_23744);
nor U24263 (N_24263,N_23679,N_23601);
xnor U24264 (N_24264,N_23819,N_23755);
and U24265 (N_24265,N_23683,N_23905);
and U24266 (N_24266,N_23794,N_23615);
or U24267 (N_24267,N_23637,N_23594);
xnor U24268 (N_24268,N_23974,N_23502);
xnor U24269 (N_24269,N_23516,N_23557);
and U24270 (N_24270,N_23803,N_23801);
xor U24271 (N_24271,N_23651,N_23537);
and U24272 (N_24272,N_23792,N_23777);
nor U24273 (N_24273,N_23879,N_23760);
nor U24274 (N_24274,N_23502,N_23733);
or U24275 (N_24275,N_23823,N_23953);
or U24276 (N_24276,N_23500,N_23822);
nand U24277 (N_24277,N_23649,N_23542);
xnor U24278 (N_24278,N_23807,N_23774);
xor U24279 (N_24279,N_23943,N_23880);
nand U24280 (N_24280,N_23945,N_23943);
nand U24281 (N_24281,N_23510,N_23815);
and U24282 (N_24282,N_23817,N_23744);
nor U24283 (N_24283,N_23860,N_23768);
xnor U24284 (N_24284,N_23596,N_23675);
xor U24285 (N_24285,N_23986,N_23671);
and U24286 (N_24286,N_23626,N_23821);
nand U24287 (N_24287,N_23970,N_23519);
nor U24288 (N_24288,N_23774,N_23828);
nand U24289 (N_24289,N_23942,N_23801);
nand U24290 (N_24290,N_23771,N_23719);
xnor U24291 (N_24291,N_23981,N_23658);
nor U24292 (N_24292,N_23522,N_23723);
nor U24293 (N_24293,N_23957,N_23947);
nand U24294 (N_24294,N_23674,N_23620);
nor U24295 (N_24295,N_23672,N_23887);
or U24296 (N_24296,N_23793,N_23635);
nor U24297 (N_24297,N_23714,N_23941);
nor U24298 (N_24298,N_23652,N_23830);
or U24299 (N_24299,N_23749,N_23680);
xor U24300 (N_24300,N_23604,N_23981);
and U24301 (N_24301,N_23757,N_23744);
xnor U24302 (N_24302,N_23773,N_23829);
and U24303 (N_24303,N_23657,N_23656);
or U24304 (N_24304,N_23811,N_23762);
nand U24305 (N_24305,N_23842,N_23536);
nor U24306 (N_24306,N_23821,N_23514);
and U24307 (N_24307,N_23681,N_23783);
nand U24308 (N_24308,N_23580,N_23758);
nor U24309 (N_24309,N_23830,N_23996);
nor U24310 (N_24310,N_23764,N_23713);
and U24311 (N_24311,N_23961,N_23690);
and U24312 (N_24312,N_23605,N_23831);
and U24313 (N_24313,N_23656,N_23969);
nor U24314 (N_24314,N_23902,N_23609);
nor U24315 (N_24315,N_23856,N_23747);
and U24316 (N_24316,N_23516,N_23809);
nand U24317 (N_24317,N_23573,N_23811);
nor U24318 (N_24318,N_23913,N_23733);
and U24319 (N_24319,N_23752,N_23896);
and U24320 (N_24320,N_23998,N_23875);
nand U24321 (N_24321,N_23924,N_23606);
xnor U24322 (N_24322,N_23755,N_23597);
or U24323 (N_24323,N_23988,N_23742);
nand U24324 (N_24324,N_23847,N_23819);
and U24325 (N_24325,N_23751,N_23513);
xor U24326 (N_24326,N_23579,N_23772);
or U24327 (N_24327,N_23552,N_23793);
nor U24328 (N_24328,N_23874,N_23742);
nand U24329 (N_24329,N_23741,N_23744);
and U24330 (N_24330,N_23520,N_23732);
or U24331 (N_24331,N_23703,N_23829);
or U24332 (N_24332,N_23890,N_23548);
nor U24333 (N_24333,N_23503,N_23850);
and U24334 (N_24334,N_23681,N_23886);
and U24335 (N_24335,N_23687,N_23585);
xnor U24336 (N_24336,N_23727,N_23927);
xnor U24337 (N_24337,N_23671,N_23923);
and U24338 (N_24338,N_23961,N_23654);
or U24339 (N_24339,N_23519,N_23549);
or U24340 (N_24340,N_23844,N_23716);
xor U24341 (N_24341,N_23724,N_23746);
xnor U24342 (N_24342,N_23676,N_23827);
or U24343 (N_24343,N_23721,N_23639);
and U24344 (N_24344,N_23997,N_23694);
or U24345 (N_24345,N_23601,N_23851);
and U24346 (N_24346,N_23742,N_23762);
nor U24347 (N_24347,N_23546,N_23778);
or U24348 (N_24348,N_23550,N_23617);
or U24349 (N_24349,N_23846,N_23702);
and U24350 (N_24350,N_23603,N_23601);
and U24351 (N_24351,N_23965,N_23870);
or U24352 (N_24352,N_23824,N_23915);
xnor U24353 (N_24353,N_23649,N_23917);
xor U24354 (N_24354,N_23941,N_23913);
xnor U24355 (N_24355,N_23616,N_23562);
xor U24356 (N_24356,N_23989,N_23901);
and U24357 (N_24357,N_23873,N_23882);
nor U24358 (N_24358,N_23503,N_23727);
xor U24359 (N_24359,N_23827,N_23972);
and U24360 (N_24360,N_23566,N_23508);
xnor U24361 (N_24361,N_23531,N_23911);
nand U24362 (N_24362,N_23578,N_23996);
xor U24363 (N_24363,N_23518,N_23641);
nand U24364 (N_24364,N_23994,N_23918);
and U24365 (N_24365,N_23716,N_23694);
and U24366 (N_24366,N_23503,N_23546);
or U24367 (N_24367,N_23903,N_23500);
nor U24368 (N_24368,N_23976,N_23725);
nor U24369 (N_24369,N_23723,N_23987);
nor U24370 (N_24370,N_23795,N_23938);
nand U24371 (N_24371,N_23741,N_23546);
and U24372 (N_24372,N_23885,N_23599);
nor U24373 (N_24373,N_23713,N_23891);
and U24374 (N_24374,N_23889,N_23714);
and U24375 (N_24375,N_23642,N_23929);
xnor U24376 (N_24376,N_23786,N_23817);
nand U24377 (N_24377,N_23770,N_23541);
or U24378 (N_24378,N_23663,N_23755);
nor U24379 (N_24379,N_23833,N_23613);
and U24380 (N_24380,N_23700,N_23548);
or U24381 (N_24381,N_23791,N_23501);
and U24382 (N_24382,N_23869,N_23728);
and U24383 (N_24383,N_23946,N_23531);
nor U24384 (N_24384,N_23912,N_23720);
nand U24385 (N_24385,N_23724,N_23661);
xnor U24386 (N_24386,N_23533,N_23850);
and U24387 (N_24387,N_23929,N_23589);
nand U24388 (N_24388,N_23712,N_23596);
and U24389 (N_24389,N_23630,N_23785);
nor U24390 (N_24390,N_23942,N_23888);
nor U24391 (N_24391,N_23512,N_23922);
nand U24392 (N_24392,N_23578,N_23523);
or U24393 (N_24393,N_23828,N_23834);
and U24394 (N_24394,N_23758,N_23964);
or U24395 (N_24395,N_23616,N_23531);
nand U24396 (N_24396,N_23723,N_23976);
nor U24397 (N_24397,N_23897,N_23829);
and U24398 (N_24398,N_23918,N_23536);
xnor U24399 (N_24399,N_23580,N_23555);
and U24400 (N_24400,N_23746,N_23728);
or U24401 (N_24401,N_23865,N_23820);
and U24402 (N_24402,N_23579,N_23756);
nor U24403 (N_24403,N_23863,N_23824);
nor U24404 (N_24404,N_23567,N_23884);
and U24405 (N_24405,N_23580,N_23906);
xor U24406 (N_24406,N_23756,N_23640);
nor U24407 (N_24407,N_23977,N_23912);
and U24408 (N_24408,N_23808,N_23618);
nand U24409 (N_24409,N_23989,N_23945);
or U24410 (N_24410,N_23819,N_23942);
and U24411 (N_24411,N_23756,N_23859);
and U24412 (N_24412,N_23803,N_23596);
or U24413 (N_24413,N_23548,N_23710);
or U24414 (N_24414,N_23573,N_23684);
nand U24415 (N_24415,N_23746,N_23645);
and U24416 (N_24416,N_23854,N_23604);
or U24417 (N_24417,N_23785,N_23535);
or U24418 (N_24418,N_23512,N_23972);
nand U24419 (N_24419,N_23831,N_23952);
and U24420 (N_24420,N_23682,N_23931);
or U24421 (N_24421,N_23692,N_23673);
or U24422 (N_24422,N_23682,N_23743);
or U24423 (N_24423,N_23670,N_23654);
nand U24424 (N_24424,N_23882,N_23953);
nand U24425 (N_24425,N_23602,N_23775);
or U24426 (N_24426,N_23742,N_23637);
or U24427 (N_24427,N_23987,N_23738);
and U24428 (N_24428,N_23804,N_23833);
and U24429 (N_24429,N_23536,N_23712);
or U24430 (N_24430,N_23533,N_23681);
and U24431 (N_24431,N_23688,N_23604);
and U24432 (N_24432,N_23570,N_23635);
or U24433 (N_24433,N_23704,N_23824);
xor U24434 (N_24434,N_23558,N_23631);
or U24435 (N_24435,N_23589,N_23652);
or U24436 (N_24436,N_23503,N_23626);
nand U24437 (N_24437,N_23511,N_23538);
or U24438 (N_24438,N_23521,N_23975);
nand U24439 (N_24439,N_23833,N_23746);
or U24440 (N_24440,N_23657,N_23912);
nand U24441 (N_24441,N_23601,N_23855);
xnor U24442 (N_24442,N_23881,N_23527);
nor U24443 (N_24443,N_23777,N_23524);
xnor U24444 (N_24444,N_23812,N_23998);
xnor U24445 (N_24445,N_23946,N_23750);
and U24446 (N_24446,N_23961,N_23779);
nor U24447 (N_24447,N_23795,N_23605);
xnor U24448 (N_24448,N_23903,N_23917);
xnor U24449 (N_24449,N_23952,N_23824);
xor U24450 (N_24450,N_23803,N_23796);
nor U24451 (N_24451,N_23562,N_23808);
xnor U24452 (N_24452,N_23670,N_23831);
and U24453 (N_24453,N_23712,N_23873);
and U24454 (N_24454,N_23669,N_23705);
nor U24455 (N_24455,N_23901,N_23918);
xnor U24456 (N_24456,N_23545,N_23949);
or U24457 (N_24457,N_23889,N_23672);
or U24458 (N_24458,N_23675,N_23828);
xnor U24459 (N_24459,N_23672,N_23921);
xnor U24460 (N_24460,N_23764,N_23507);
nand U24461 (N_24461,N_23882,N_23643);
or U24462 (N_24462,N_23719,N_23500);
nor U24463 (N_24463,N_23741,N_23560);
or U24464 (N_24464,N_23912,N_23813);
and U24465 (N_24465,N_23903,N_23603);
nor U24466 (N_24466,N_23811,N_23742);
nor U24467 (N_24467,N_23503,N_23704);
xor U24468 (N_24468,N_23707,N_23691);
nand U24469 (N_24469,N_23640,N_23696);
xor U24470 (N_24470,N_23684,N_23720);
nand U24471 (N_24471,N_23859,N_23601);
nand U24472 (N_24472,N_23558,N_23972);
nor U24473 (N_24473,N_23604,N_23964);
or U24474 (N_24474,N_23681,N_23626);
and U24475 (N_24475,N_23911,N_23746);
or U24476 (N_24476,N_23568,N_23769);
xnor U24477 (N_24477,N_23820,N_23960);
xnor U24478 (N_24478,N_23971,N_23505);
nand U24479 (N_24479,N_23558,N_23747);
xor U24480 (N_24480,N_23650,N_23646);
xnor U24481 (N_24481,N_23695,N_23651);
nor U24482 (N_24482,N_23743,N_23669);
xnor U24483 (N_24483,N_23526,N_23788);
or U24484 (N_24484,N_23527,N_23636);
nand U24485 (N_24485,N_23589,N_23920);
xnor U24486 (N_24486,N_23566,N_23979);
xnor U24487 (N_24487,N_23583,N_23846);
and U24488 (N_24488,N_23895,N_23736);
or U24489 (N_24489,N_23832,N_23979);
nand U24490 (N_24490,N_23737,N_23937);
or U24491 (N_24491,N_23763,N_23758);
xor U24492 (N_24492,N_23993,N_23689);
nor U24493 (N_24493,N_23802,N_23770);
and U24494 (N_24494,N_23609,N_23556);
xor U24495 (N_24495,N_23974,N_23504);
xor U24496 (N_24496,N_23906,N_23636);
xor U24497 (N_24497,N_23867,N_23876);
nand U24498 (N_24498,N_23784,N_23895);
xnor U24499 (N_24499,N_23834,N_23872);
nand U24500 (N_24500,N_24044,N_24459);
or U24501 (N_24501,N_24370,N_24445);
nor U24502 (N_24502,N_24292,N_24121);
xnor U24503 (N_24503,N_24275,N_24230);
nand U24504 (N_24504,N_24216,N_24439);
nand U24505 (N_24505,N_24012,N_24355);
and U24506 (N_24506,N_24351,N_24429);
or U24507 (N_24507,N_24239,N_24327);
nor U24508 (N_24508,N_24184,N_24455);
and U24509 (N_24509,N_24022,N_24109);
xnor U24510 (N_24510,N_24110,N_24463);
nand U24511 (N_24511,N_24343,N_24192);
or U24512 (N_24512,N_24176,N_24423);
xor U24513 (N_24513,N_24381,N_24209);
nor U24514 (N_24514,N_24251,N_24193);
nor U24515 (N_24515,N_24257,N_24099);
nor U24516 (N_24516,N_24433,N_24362);
or U24517 (N_24517,N_24268,N_24454);
nand U24518 (N_24518,N_24220,N_24419);
nor U24519 (N_24519,N_24051,N_24364);
and U24520 (N_24520,N_24217,N_24005);
or U24521 (N_24521,N_24400,N_24206);
xor U24522 (N_24522,N_24138,N_24287);
and U24523 (N_24523,N_24213,N_24108);
nand U24524 (N_24524,N_24170,N_24160);
or U24525 (N_24525,N_24368,N_24376);
nand U24526 (N_24526,N_24396,N_24322);
or U24527 (N_24527,N_24117,N_24414);
nand U24528 (N_24528,N_24353,N_24191);
nor U24529 (N_24529,N_24481,N_24175);
xnor U24530 (N_24530,N_24179,N_24134);
nand U24531 (N_24531,N_24395,N_24360);
xor U24532 (N_24532,N_24237,N_24332);
nor U24533 (N_24533,N_24348,N_24072);
xor U24534 (N_24534,N_24369,N_24350);
nand U24535 (N_24535,N_24168,N_24276);
nand U24536 (N_24536,N_24073,N_24470);
xnor U24537 (N_24537,N_24201,N_24382);
nand U24538 (N_24538,N_24076,N_24035);
nand U24539 (N_24539,N_24060,N_24159);
xor U24540 (N_24540,N_24386,N_24366);
or U24541 (N_24541,N_24185,N_24393);
nand U24542 (N_24542,N_24173,N_24180);
or U24543 (N_24543,N_24267,N_24405);
or U24544 (N_24544,N_24390,N_24290);
and U24545 (N_24545,N_24352,N_24320);
and U24546 (N_24546,N_24065,N_24443);
or U24547 (N_24547,N_24023,N_24247);
nor U24548 (N_24548,N_24085,N_24158);
nand U24549 (N_24549,N_24358,N_24460);
or U24550 (N_24550,N_24272,N_24204);
nand U24551 (N_24551,N_24324,N_24027);
nor U24552 (N_24552,N_24190,N_24256);
or U24553 (N_24553,N_24141,N_24208);
or U24554 (N_24554,N_24335,N_24222);
xor U24555 (N_24555,N_24248,N_24436);
xor U24556 (N_24556,N_24152,N_24171);
xnor U24557 (N_24557,N_24224,N_24140);
and U24558 (N_24558,N_24323,N_24384);
nor U24559 (N_24559,N_24069,N_24079);
and U24560 (N_24560,N_24434,N_24377);
or U24561 (N_24561,N_24032,N_24422);
nor U24562 (N_24562,N_24330,N_24318);
xnor U24563 (N_24563,N_24447,N_24467);
and U24564 (N_24564,N_24286,N_24294);
or U24565 (N_24565,N_24489,N_24404);
xnor U24566 (N_24566,N_24280,N_24244);
or U24567 (N_24567,N_24302,N_24042);
or U24568 (N_24568,N_24094,N_24164);
nor U24569 (N_24569,N_24097,N_24389);
nand U24570 (N_24570,N_24372,N_24078);
nand U24571 (N_24571,N_24071,N_24483);
xnor U24572 (N_24572,N_24137,N_24356);
or U24573 (N_24573,N_24167,N_24084);
nor U24574 (N_24574,N_24210,N_24407);
nor U24575 (N_24575,N_24034,N_24341);
and U24576 (N_24576,N_24049,N_24309);
xnor U24577 (N_24577,N_24361,N_24482);
nand U24578 (N_24578,N_24006,N_24089);
and U24579 (N_24579,N_24342,N_24145);
and U24580 (N_24580,N_24187,N_24437);
nand U24581 (N_24581,N_24004,N_24345);
xor U24582 (N_24582,N_24014,N_24074);
or U24583 (N_24583,N_24139,N_24298);
or U24584 (N_24584,N_24003,N_24253);
nand U24585 (N_24585,N_24178,N_24315);
nor U24586 (N_24586,N_24354,N_24040);
and U24587 (N_24587,N_24231,N_24314);
nor U24588 (N_24588,N_24056,N_24043);
nand U24589 (N_24589,N_24046,N_24091);
xor U24590 (N_24590,N_24313,N_24162);
nand U24591 (N_24591,N_24144,N_24235);
nor U24592 (N_24592,N_24474,N_24277);
xnor U24593 (N_24593,N_24106,N_24111);
xor U24594 (N_24594,N_24061,N_24449);
and U24595 (N_24595,N_24258,N_24096);
or U24596 (N_24596,N_24157,N_24103);
nor U24597 (N_24597,N_24234,N_24402);
and U24598 (N_24598,N_24118,N_24095);
and U24599 (N_24599,N_24226,N_24126);
xnor U24600 (N_24600,N_24128,N_24207);
and U24601 (N_24601,N_24189,N_24462);
and U24602 (N_24602,N_24435,N_24050);
xnor U24603 (N_24603,N_24497,N_24048);
nand U24604 (N_24604,N_24245,N_24221);
nand U24605 (N_24605,N_24306,N_24303);
nand U24606 (N_24606,N_24321,N_24365);
and U24607 (N_24607,N_24194,N_24392);
and U24608 (N_24608,N_24344,N_24143);
and U24609 (N_24609,N_24054,N_24359);
xor U24610 (N_24610,N_24196,N_24147);
nor U24611 (N_24611,N_24397,N_24293);
nand U24612 (N_24612,N_24347,N_24053);
and U24613 (N_24613,N_24485,N_24146);
nor U24614 (N_24614,N_24200,N_24086);
nand U24615 (N_24615,N_24476,N_24255);
nand U24616 (N_24616,N_24018,N_24241);
xnor U24617 (N_24617,N_24197,N_24148);
and U24618 (N_24618,N_24181,N_24457);
nor U24619 (N_24619,N_24047,N_24249);
nand U24620 (N_24620,N_24316,N_24112);
and U24621 (N_24621,N_24409,N_24172);
nor U24622 (N_24622,N_24163,N_24448);
nor U24623 (N_24623,N_24310,N_24100);
nand U24624 (N_24624,N_24289,N_24438);
nor U24625 (N_24625,N_24024,N_24278);
and U24626 (N_24626,N_24471,N_24312);
xor U24627 (N_24627,N_24317,N_24420);
nand U24628 (N_24628,N_24016,N_24093);
xnor U24629 (N_24629,N_24406,N_24031);
nand U24630 (N_24630,N_24285,N_24122);
and U24631 (N_24631,N_24464,N_24233);
nand U24632 (N_24632,N_24385,N_24057);
nor U24633 (N_24633,N_24379,N_24301);
xnor U24634 (N_24634,N_24304,N_24166);
nor U24635 (N_24635,N_24215,N_24300);
and U24636 (N_24636,N_24183,N_24487);
nor U24637 (N_24637,N_24064,N_24263);
and U24638 (N_24638,N_24388,N_24426);
or U24639 (N_24639,N_24349,N_24119);
nand U24640 (N_24640,N_24068,N_24161);
nor U24641 (N_24641,N_24446,N_24142);
nor U24642 (N_24642,N_24266,N_24199);
nand U24643 (N_24643,N_24001,N_24416);
xor U24644 (N_24644,N_24363,N_24188);
xor U24645 (N_24645,N_24123,N_24228);
nand U24646 (N_24646,N_24325,N_24214);
nand U24647 (N_24647,N_24394,N_24334);
and U24648 (N_24648,N_24410,N_24299);
nand U24649 (N_24649,N_24088,N_24262);
and U24650 (N_24650,N_24480,N_24424);
or U24651 (N_24651,N_24430,N_24092);
xor U24652 (N_24652,N_24133,N_24261);
and U24653 (N_24653,N_24038,N_24432);
or U24654 (N_24654,N_24329,N_24367);
xnor U24655 (N_24655,N_24479,N_24259);
and U24656 (N_24656,N_24378,N_24328);
and U24657 (N_24657,N_24254,N_24127);
and U24658 (N_24658,N_24337,N_24130);
and U24659 (N_24659,N_24223,N_24295);
nand U24660 (N_24660,N_24296,N_24002);
or U24661 (N_24661,N_24154,N_24490);
xor U24662 (N_24662,N_24177,N_24427);
or U24663 (N_24663,N_24113,N_24238);
and U24664 (N_24664,N_24486,N_24101);
nand U24665 (N_24665,N_24075,N_24475);
and U24666 (N_24666,N_24131,N_24013);
or U24667 (N_24667,N_24284,N_24346);
nand U24668 (N_24668,N_24339,N_24391);
nor U24669 (N_24669,N_24403,N_24058);
nand U24670 (N_24670,N_24205,N_24399);
xor U24671 (N_24671,N_24070,N_24030);
or U24672 (N_24672,N_24492,N_24229);
nand U24673 (N_24673,N_24020,N_24059);
xor U24674 (N_24674,N_24007,N_24311);
and U24675 (N_24675,N_24288,N_24431);
xnor U24676 (N_24676,N_24107,N_24270);
and U24677 (N_24677,N_24246,N_24124);
and U24678 (N_24678,N_24308,N_24104);
or U24679 (N_24679,N_24375,N_24102);
nand U24680 (N_24680,N_24491,N_24029);
nor U24681 (N_24681,N_24331,N_24062);
nor U24682 (N_24682,N_24472,N_24273);
nor U24683 (N_24683,N_24036,N_24469);
nand U24684 (N_24684,N_24252,N_24212);
nor U24685 (N_24685,N_24081,N_24495);
nand U24686 (N_24686,N_24225,N_24488);
nor U24687 (N_24687,N_24498,N_24105);
nand U24688 (N_24688,N_24125,N_24153);
or U24689 (N_24689,N_24452,N_24473);
nand U24690 (N_24690,N_24037,N_24045);
nand U24691 (N_24691,N_24242,N_24319);
or U24692 (N_24692,N_24440,N_24282);
and U24693 (N_24693,N_24357,N_24465);
nor U24694 (N_24694,N_24082,N_24418);
and U24695 (N_24695,N_24067,N_24456);
nor U24696 (N_24696,N_24371,N_24401);
and U24697 (N_24697,N_24063,N_24307);
and U24698 (N_24698,N_24496,N_24055);
xnor U24699 (N_24699,N_24417,N_24198);
nor U24700 (N_24700,N_24466,N_24265);
or U24701 (N_24701,N_24033,N_24236);
xnor U24702 (N_24702,N_24129,N_24116);
and U24703 (N_24703,N_24039,N_24305);
or U24704 (N_24704,N_24203,N_24021);
or U24705 (N_24705,N_24136,N_24494);
nand U24706 (N_24706,N_24428,N_24009);
and U24707 (N_24707,N_24413,N_24383);
xor U24708 (N_24708,N_24019,N_24380);
or U24709 (N_24709,N_24291,N_24408);
nand U24710 (N_24710,N_24015,N_24468);
and U24711 (N_24711,N_24477,N_24442);
or U24712 (N_24712,N_24326,N_24011);
nand U24713 (N_24713,N_24010,N_24269);
nor U24714 (N_24714,N_24333,N_24398);
and U24715 (N_24715,N_24336,N_24340);
xor U24716 (N_24716,N_24120,N_24098);
or U24717 (N_24717,N_24374,N_24115);
nor U24718 (N_24718,N_24026,N_24151);
or U24719 (N_24719,N_24260,N_24425);
nor U24720 (N_24720,N_24025,N_24274);
nand U24721 (N_24721,N_24017,N_24411);
and U24722 (N_24722,N_24493,N_24297);
or U24723 (N_24723,N_24090,N_24000);
xor U24724 (N_24724,N_24271,N_24202);
nor U24725 (N_24725,N_24165,N_24232);
xor U24726 (N_24726,N_24132,N_24499);
xor U24727 (N_24727,N_24387,N_24373);
and U24728 (N_24728,N_24484,N_24087);
or U24729 (N_24729,N_24250,N_24135);
xor U24730 (N_24730,N_24338,N_24169);
and U24731 (N_24731,N_24243,N_24114);
nand U24732 (N_24732,N_24450,N_24008);
and U24733 (N_24733,N_24195,N_24066);
nor U24734 (N_24734,N_24451,N_24458);
nor U24735 (N_24735,N_24052,N_24461);
or U24736 (N_24736,N_24149,N_24279);
nand U24737 (N_24737,N_24441,N_24211);
nor U24738 (N_24738,N_24264,N_24444);
nand U24739 (N_24739,N_24421,N_24240);
nor U24740 (N_24740,N_24186,N_24283);
nand U24741 (N_24741,N_24156,N_24028);
nand U24742 (N_24742,N_24227,N_24041);
xor U24743 (N_24743,N_24219,N_24453);
or U24744 (N_24744,N_24080,N_24174);
or U24745 (N_24745,N_24182,N_24155);
or U24746 (N_24746,N_24478,N_24218);
and U24747 (N_24747,N_24077,N_24412);
xnor U24748 (N_24748,N_24150,N_24281);
xor U24749 (N_24749,N_24083,N_24415);
and U24750 (N_24750,N_24467,N_24458);
xor U24751 (N_24751,N_24422,N_24154);
nand U24752 (N_24752,N_24333,N_24117);
and U24753 (N_24753,N_24444,N_24077);
nor U24754 (N_24754,N_24332,N_24301);
xnor U24755 (N_24755,N_24266,N_24280);
and U24756 (N_24756,N_24486,N_24022);
and U24757 (N_24757,N_24235,N_24391);
nand U24758 (N_24758,N_24222,N_24381);
nor U24759 (N_24759,N_24285,N_24397);
and U24760 (N_24760,N_24184,N_24334);
nand U24761 (N_24761,N_24164,N_24203);
nand U24762 (N_24762,N_24188,N_24136);
nand U24763 (N_24763,N_24130,N_24164);
xor U24764 (N_24764,N_24187,N_24479);
xor U24765 (N_24765,N_24458,N_24212);
nand U24766 (N_24766,N_24296,N_24484);
or U24767 (N_24767,N_24044,N_24113);
nand U24768 (N_24768,N_24123,N_24379);
and U24769 (N_24769,N_24178,N_24330);
nor U24770 (N_24770,N_24432,N_24095);
xnor U24771 (N_24771,N_24401,N_24196);
xor U24772 (N_24772,N_24420,N_24446);
nor U24773 (N_24773,N_24085,N_24340);
xnor U24774 (N_24774,N_24453,N_24345);
nor U24775 (N_24775,N_24381,N_24238);
xnor U24776 (N_24776,N_24437,N_24412);
xor U24777 (N_24777,N_24045,N_24309);
nand U24778 (N_24778,N_24254,N_24246);
xnor U24779 (N_24779,N_24292,N_24319);
and U24780 (N_24780,N_24057,N_24201);
nand U24781 (N_24781,N_24281,N_24298);
nor U24782 (N_24782,N_24207,N_24027);
and U24783 (N_24783,N_24308,N_24120);
and U24784 (N_24784,N_24457,N_24417);
or U24785 (N_24785,N_24189,N_24024);
or U24786 (N_24786,N_24475,N_24027);
or U24787 (N_24787,N_24348,N_24107);
nand U24788 (N_24788,N_24362,N_24039);
nor U24789 (N_24789,N_24220,N_24217);
and U24790 (N_24790,N_24107,N_24173);
xnor U24791 (N_24791,N_24135,N_24001);
xor U24792 (N_24792,N_24309,N_24484);
nor U24793 (N_24793,N_24199,N_24289);
nand U24794 (N_24794,N_24215,N_24035);
nand U24795 (N_24795,N_24264,N_24107);
nand U24796 (N_24796,N_24136,N_24403);
or U24797 (N_24797,N_24352,N_24159);
nor U24798 (N_24798,N_24294,N_24312);
or U24799 (N_24799,N_24173,N_24441);
xor U24800 (N_24800,N_24418,N_24205);
and U24801 (N_24801,N_24203,N_24044);
nor U24802 (N_24802,N_24432,N_24482);
and U24803 (N_24803,N_24110,N_24023);
and U24804 (N_24804,N_24429,N_24041);
xnor U24805 (N_24805,N_24071,N_24043);
xnor U24806 (N_24806,N_24230,N_24003);
and U24807 (N_24807,N_24267,N_24416);
xnor U24808 (N_24808,N_24448,N_24309);
and U24809 (N_24809,N_24348,N_24428);
and U24810 (N_24810,N_24083,N_24361);
nor U24811 (N_24811,N_24468,N_24052);
xor U24812 (N_24812,N_24494,N_24109);
and U24813 (N_24813,N_24404,N_24017);
or U24814 (N_24814,N_24107,N_24098);
nor U24815 (N_24815,N_24150,N_24027);
or U24816 (N_24816,N_24375,N_24420);
or U24817 (N_24817,N_24080,N_24327);
nor U24818 (N_24818,N_24127,N_24100);
and U24819 (N_24819,N_24042,N_24182);
xor U24820 (N_24820,N_24168,N_24413);
nand U24821 (N_24821,N_24248,N_24475);
nor U24822 (N_24822,N_24469,N_24145);
and U24823 (N_24823,N_24267,N_24356);
and U24824 (N_24824,N_24175,N_24248);
or U24825 (N_24825,N_24375,N_24142);
nand U24826 (N_24826,N_24178,N_24496);
xor U24827 (N_24827,N_24042,N_24169);
and U24828 (N_24828,N_24463,N_24029);
xnor U24829 (N_24829,N_24103,N_24149);
xor U24830 (N_24830,N_24391,N_24177);
and U24831 (N_24831,N_24300,N_24331);
nor U24832 (N_24832,N_24072,N_24344);
nor U24833 (N_24833,N_24221,N_24357);
xor U24834 (N_24834,N_24357,N_24127);
nor U24835 (N_24835,N_24169,N_24126);
or U24836 (N_24836,N_24010,N_24393);
nand U24837 (N_24837,N_24045,N_24133);
nor U24838 (N_24838,N_24494,N_24015);
nor U24839 (N_24839,N_24161,N_24426);
or U24840 (N_24840,N_24015,N_24389);
nand U24841 (N_24841,N_24370,N_24120);
and U24842 (N_24842,N_24410,N_24106);
nand U24843 (N_24843,N_24144,N_24217);
xor U24844 (N_24844,N_24121,N_24207);
nor U24845 (N_24845,N_24104,N_24074);
or U24846 (N_24846,N_24392,N_24453);
nor U24847 (N_24847,N_24332,N_24484);
and U24848 (N_24848,N_24469,N_24492);
nand U24849 (N_24849,N_24143,N_24360);
and U24850 (N_24850,N_24021,N_24499);
xor U24851 (N_24851,N_24339,N_24121);
or U24852 (N_24852,N_24000,N_24439);
xnor U24853 (N_24853,N_24077,N_24061);
xor U24854 (N_24854,N_24127,N_24225);
or U24855 (N_24855,N_24196,N_24358);
nor U24856 (N_24856,N_24252,N_24048);
and U24857 (N_24857,N_24160,N_24493);
nand U24858 (N_24858,N_24122,N_24154);
or U24859 (N_24859,N_24238,N_24248);
and U24860 (N_24860,N_24374,N_24386);
or U24861 (N_24861,N_24195,N_24285);
nand U24862 (N_24862,N_24067,N_24083);
and U24863 (N_24863,N_24413,N_24222);
nand U24864 (N_24864,N_24283,N_24431);
nor U24865 (N_24865,N_24455,N_24303);
nor U24866 (N_24866,N_24021,N_24413);
xnor U24867 (N_24867,N_24487,N_24198);
nor U24868 (N_24868,N_24138,N_24484);
nand U24869 (N_24869,N_24411,N_24254);
xor U24870 (N_24870,N_24232,N_24144);
xor U24871 (N_24871,N_24010,N_24494);
and U24872 (N_24872,N_24196,N_24270);
or U24873 (N_24873,N_24482,N_24161);
or U24874 (N_24874,N_24437,N_24001);
or U24875 (N_24875,N_24039,N_24365);
nand U24876 (N_24876,N_24417,N_24094);
nand U24877 (N_24877,N_24399,N_24274);
and U24878 (N_24878,N_24257,N_24411);
nor U24879 (N_24879,N_24177,N_24162);
and U24880 (N_24880,N_24474,N_24425);
and U24881 (N_24881,N_24417,N_24360);
nor U24882 (N_24882,N_24437,N_24395);
and U24883 (N_24883,N_24014,N_24307);
nor U24884 (N_24884,N_24184,N_24438);
xor U24885 (N_24885,N_24360,N_24462);
or U24886 (N_24886,N_24113,N_24339);
nor U24887 (N_24887,N_24030,N_24389);
or U24888 (N_24888,N_24212,N_24067);
or U24889 (N_24889,N_24109,N_24331);
nor U24890 (N_24890,N_24016,N_24124);
or U24891 (N_24891,N_24308,N_24003);
xnor U24892 (N_24892,N_24289,N_24377);
nor U24893 (N_24893,N_24400,N_24402);
or U24894 (N_24894,N_24354,N_24232);
nand U24895 (N_24895,N_24084,N_24378);
and U24896 (N_24896,N_24399,N_24271);
nand U24897 (N_24897,N_24144,N_24264);
nor U24898 (N_24898,N_24424,N_24320);
nor U24899 (N_24899,N_24395,N_24024);
or U24900 (N_24900,N_24340,N_24181);
or U24901 (N_24901,N_24317,N_24028);
nor U24902 (N_24902,N_24008,N_24223);
or U24903 (N_24903,N_24391,N_24223);
nor U24904 (N_24904,N_24166,N_24049);
nor U24905 (N_24905,N_24005,N_24193);
and U24906 (N_24906,N_24000,N_24166);
xnor U24907 (N_24907,N_24214,N_24033);
and U24908 (N_24908,N_24204,N_24488);
or U24909 (N_24909,N_24380,N_24090);
or U24910 (N_24910,N_24111,N_24115);
nand U24911 (N_24911,N_24025,N_24370);
and U24912 (N_24912,N_24035,N_24287);
and U24913 (N_24913,N_24075,N_24402);
nor U24914 (N_24914,N_24293,N_24303);
xor U24915 (N_24915,N_24014,N_24478);
and U24916 (N_24916,N_24186,N_24219);
and U24917 (N_24917,N_24395,N_24031);
or U24918 (N_24918,N_24061,N_24429);
or U24919 (N_24919,N_24068,N_24391);
nor U24920 (N_24920,N_24141,N_24425);
xnor U24921 (N_24921,N_24153,N_24096);
xor U24922 (N_24922,N_24143,N_24054);
xor U24923 (N_24923,N_24208,N_24432);
nor U24924 (N_24924,N_24383,N_24135);
or U24925 (N_24925,N_24489,N_24119);
nor U24926 (N_24926,N_24471,N_24291);
xor U24927 (N_24927,N_24422,N_24181);
or U24928 (N_24928,N_24134,N_24211);
nor U24929 (N_24929,N_24488,N_24041);
or U24930 (N_24930,N_24138,N_24034);
xor U24931 (N_24931,N_24023,N_24037);
nor U24932 (N_24932,N_24315,N_24448);
xor U24933 (N_24933,N_24067,N_24284);
nor U24934 (N_24934,N_24097,N_24049);
or U24935 (N_24935,N_24308,N_24354);
and U24936 (N_24936,N_24318,N_24391);
and U24937 (N_24937,N_24359,N_24304);
nor U24938 (N_24938,N_24054,N_24432);
nor U24939 (N_24939,N_24379,N_24276);
nor U24940 (N_24940,N_24417,N_24341);
nor U24941 (N_24941,N_24121,N_24478);
nor U24942 (N_24942,N_24194,N_24404);
nand U24943 (N_24943,N_24367,N_24472);
and U24944 (N_24944,N_24243,N_24129);
and U24945 (N_24945,N_24077,N_24346);
and U24946 (N_24946,N_24229,N_24064);
and U24947 (N_24947,N_24483,N_24143);
nor U24948 (N_24948,N_24290,N_24166);
or U24949 (N_24949,N_24414,N_24261);
or U24950 (N_24950,N_24252,N_24495);
nor U24951 (N_24951,N_24017,N_24324);
and U24952 (N_24952,N_24084,N_24400);
or U24953 (N_24953,N_24053,N_24429);
xnor U24954 (N_24954,N_24481,N_24061);
xor U24955 (N_24955,N_24271,N_24361);
and U24956 (N_24956,N_24162,N_24462);
nand U24957 (N_24957,N_24061,N_24355);
or U24958 (N_24958,N_24381,N_24094);
nand U24959 (N_24959,N_24439,N_24355);
and U24960 (N_24960,N_24124,N_24495);
or U24961 (N_24961,N_24045,N_24044);
and U24962 (N_24962,N_24260,N_24012);
or U24963 (N_24963,N_24257,N_24175);
and U24964 (N_24964,N_24118,N_24224);
nand U24965 (N_24965,N_24214,N_24054);
nor U24966 (N_24966,N_24210,N_24017);
nand U24967 (N_24967,N_24375,N_24214);
xnor U24968 (N_24968,N_24247,N_24350);
nand U24969 (N_24969,N_24330,N_24327);
xnor U24970 (N_24970,N_24141,N_24130);
or U24971 (N_24971,N_24054,N_24125);
and U24972 (N_24972,N_24264,N_24461);
xor U24973 (N_24973,N_24494,N_24454);
nor U24974 (N_24974,N_24232,N_24195);
and U24975 (N_24975,N_24465,N_24241);
nor U24976 (N_24976,N_24325,N_24382);
and U24977 (N_24977,N_24258,N_24458);
xor U24978 (N_24978,N_24089,N_24366);
nor U24979 (N_24979,N_24233,N_24486);
nor U24980 (N_24980,N_24278,N_24322);
nor U24981 (N_24981,N_24111,N_24469);
nor U24982 (N_24982,N_24250,N_24130);
or U24983 (N_24983,N_24332,N_24153);
or U24984 (N_24984,N_24208,N_24225);
nor U24985 (N_24985,N_24276,N_24458);
and U24986 (N_24986,N_24328,N_24389);
and U24987 (N_24987,N_24075,N_24240);
xor U24988 (N_24988,N_24468,N_24443);
nand U24989 (N_24989,N_24380,N_24386);
and U24990 (N_24990,N_24491,N_24246);
nand U24991 (N_24991,N_24365,N_24341);
or U24992 (N_24992,N_24463,N_24292);
nor U24993 (N_24993,N_24353,N_24355);
and U24994 (N_24994,N_24146,N_24103);
nand U24995 (N_24995,N_24386,N_24468);
xnor U24996 (N_24996,N_24351,N_24041);
and U24997 (N_24997,N_24261,N_24016);
nand U24998 (N_24998,N_24453,N_24498);
xor U24999 (N_24999,N_24064,N_24212);
xnor UO_0 (O_0,N_24838,N_24821);
and UO_1 (O_1,N_24706,N_24971);
or UO_2 (O_2,N_24962,N_24806);
nor UO_3 (O_3,N_24635,N_24647);
and UO_4 (O_4,N_24568,N_24809);
and UO_5 (O_5,N_24612,N_24674);
and UO_6 (O_6,N_24856,N_24965);
nand UO_7 (O_7,N_24650,N_24883);
or UO_8 (O_8,N_24508,N_24756);
and UO_9 (O_9,N_24571,N_24894);
and UO_10 (O_10,N_24545,N_24517);
xnor UO_11 (O_11,N_24890,N_24524);
nor UO_12 (O_12,N_24614,N_24819);
xnor UO_13 (O_13,N_24727,N_24698);
and UO_14 (O_14,N_24736,N_24699);
xor UO_15 (O_15,N_24666,N_24749);
xor UO_16 (O_16,N_24818,N_24869);
nor UO_17 (O_17,N_24795,N_24866);
and UO_18 (O_18,N_24774,N_24880);
xnor UO_19 (O_19,N_24903,N_24624);
and UO_20 (O_20,N_24623,N_24832);
or UO_21 (O_21,N_24796,N_24874);
or UO_22 (O_22,N_24574,N_24501);
or UO_23 (O_23,N_24948,N_24695);
nor UO_24 (O_24,N_24569,N_24761);
xor UO_25 (O_25,N_24802,N_24520);
nor UO_26 (O_26,N_24692,N_24788);
or UO_27 (O_27,N_24608,N_24533);
nand UO_28 (O_28,N_24630,N_24743);
nand UO_29 (O_29,N_24675,N_24567);
nand UO_30 (O_30,N_24741,N_24987);
nand UO_31 (O_31,N_24912,N_24882);
nor UO_32 (O_32,N_24844,N_24931);
xor UO_33 (O_33,N_24689,N_24671);
xor UO_34 (O_34,N_24585,N_24813);
nand UO_35 (O_35,N_24824,N_24629);
nand UO_36 (O_36,N_24747,N_24872);
nand UO_37 (O_37,N_24785,N_24851);
nor UO_38 (O_38,N_24507,N_24729);
nor UO_39 (O_39,N_24922,N_24678);
or UO_40 (O_40,N_24937,N_24659);
xor UO_41 (O_41,N_24786,N_24591);
nand UO_42 (O_42,N_24921,N_24999);
and UO_43 (O_43,N_24713,N_24564);
or UO_44 (O_44,N_24976,N_24864);
nor UO_45 (O_45,N_24655,N_24817);
nor UO_46 (O_46,N_24970,N_24925);
or UO_47 (O_47,N_24897,N_24710);
and UO_48 (O_48,N_24980,N_24611);
and UO_49 (O_49,N_24943,N_24810);
and UO_50 (O_50,N_24535,N_24904);
nand UO_51 (O_51,N_24836,N_24783);
xor UO_52 (O_52,N_24557,N_24654);
nand UO_53 (O_53,N_24870,N_24637);
or UO_54 (O_54,N_24909,N_24621);
nand UO_55 (O_55,N_24530,N_24670);
and UO_56 (O_56,N_24771,N_24644);
nor UO_57 (O_57,N_24900,N_24748);
and UO_58 (O_58,N_24638,N_24827);
xnor UO_59 (O_59,N_24561,N_24934);
nand UO_60 (O_60,N_24893,N_24791);
nand UO_61 (O_61,N_24515,N_24724);
nor UO_62 (O_62,N_24661,N_24878);
nand UO_63 (O_63,N_24757,N_24526);
and UO_64 (O_64,N_24553,N_24738);
xnor UO_65 (O_65,N_24728,N_24512);
nor UO_66 (O_66,N_24660,N_24719);
or UO_67 (O_67,N_24594,N_24596);
and UO_68 (O_68,N_24688,N_24877);
nor UO_69 (O_69,N_24677,N_24812);
nor UO_70 (O_70,N_24717,N_24841);
nand UO_71 (O_71,N_24926,N_24718);
and UO_72 (O_72,N_24589,N_24981);
and UO_73 (O_73,N_24775,N_24627);
or UO_74 (O_74,N_24658,N_24899);
nand UO_75 (O_75,N_24684,N_24781);
or UO_76 (O_76,N_24763,N_24834);
xnor UO_77 (O_77,N_24576,N_24952);
nor UO_78 (O_78,N_24853,N_24509);
and UO_79 (O_79,N_24665,N_24816);
nor UO_80 (O_80,N_24750,N_24735);
nand UO_81 (O_81,N_24707,N_24805);
or UO_82 (O_82,N_24759,N_24914);
and UO_83 (O_83,N_24908,N_24973);
and UO_84 (O_84,N_24778,N_24544);
nand UO_85 (O_85,N_24703,N_24930);
nand UO_86 (O_86,N_24811,N_24680);
or UO_87 (O_87,N_24823,N_24598);
nor UO_88 (O_88,N_24601,N_24705);
and UO_89 (O_89,N_24850,N_24798);
or UO_90 (O_90,N_24579,N_24932);
nor UO_91 (O_91,N_24541,N_24807);
nor UO_92 (O_92,N_24839,N_24907);
or UO_93 (O_93,N_24984,N_24988);
and UO_94 (O_94,N_24975,N_24694);
or UO_95 (O_95,N_24620,N_24780);
or UO_96 (O_96,N_24822,N_24875);
or UO_97 (O_97,N_24708,N_24916);
and UO_98 (O_98,N_24825,N_24518);
or UO_99 (O_99,N_24646,N_24935);
nand UO_100 (O_100,N_24527,N_24887);
nor UO_101 (O_101,N_24986,N_24969);
xor UO_102 (O_102,N_24884,N_24555);
or UO_103 (O_103,N_24672,N_24599);
xor UO_104 (O_104,N_24504,N_24842);
or UO_105 (O_105,N_24927,N_24577);
and UO_106 (O_106,N_24615,N_24733);
nor UO_107 (O_107,N_24691,N_24686);
nand UO_108 (O_108,N_24919,N_24715);
or UO_109 (O_109,N_24978,N_24732);
nand UO_110 (O_110,N_24559,N_24529);
or UO_111 (O_111,N_24920,N_24974);
nor UO_112 (O_112,N_24828,N_24998);
and UO_113 (O_113,N_24833,N_24632);
and UO_114 (O_114,N_24901,N_24863);
nor UO_115 (O_115,N_24871,N_24889);
and UO_116 (O_116,N_24516,N_24714);
xnor UO_117 (O_117,N_24702,N_24803);
nand UO_118 (O_118,N_24928,N_24860);
or UO_119 (O_119,N_24967,N_24959);
and UO_120 (O_120,N_24613,N_24896);
or UO_121 (O_121,N_24633,N_24622);
and UO_122 (O_122,N_24610,N_24532);
and UO_123 (O_123,N_24575,N_24996);
or UO_124 (O_124,N_24603,N_24657);
and UO_125 (O_125,N_24709,N_24949);
or UO_126 (O_126,N_24794,N_24734);
nand UO_127 (O_127,N_24991,N_24543);
nor UO_128 (O_128,N_24641,N_24906);
or UO_129 (O_129,N_24751,N_24500);
or UO_130 (O_130,N_24945,N_24835);
and UO_131 (O_131,N_24606,N_24799);
nor UO_132 (O_132,N_24639,N_24837);
and UO_133 (O_133,N_24848,N_24563);
and UO_134 (O_134,N_24859,N_24740);
and UO_135 (O_135,N_24958,N_24886);
and UO_136 (O_136,N_24548,N_24525);
and UO_137 (O_137,N_24755,N_24720);
and UO_138 (O_138,N_24942,N_24595);
nand UO_139 (O_139,N_24626,N_24648);
and UO_140 (O_140,N_24804,N_24829);
nand UO_141 (O_141,N_24768,N_24854);
nand UO_142 (O_142,N_24843,N_24765);
or UO_143 (O_143,N_24770,N_24873);
nand UO_144 (O_144,N_24929,N_24772);
and UO_145 (O_145,N_24766,N_24523);
or UO_146 (O_146,N_24676,N_24982);
nand UO_147 (O_147,N_24951,N_24570);
nand UO_148 (O_148,N_24550,N_24704);
or UO_149 (O_149,N_24528,N_24862);
xor UO_150 (O_150,N_24885,N_24552);
and UO_151 (O_151,N_24513,N_24597);
or UO_152 (O_152,N_24690,N_24793);
and UO_153 (O_153,N_24956,N_24989);
xor UO_154 (O_154,N_24721,N_24669);
nand UO_155 (O_155,N_24994,N_24758);
and UO_156 (O_156,N_24769,N_24584);
or UO_157 (O_157,N_24754,N_24619);
and UO_158 (O_158,N_24915,N_24737);
nand UO_159 (O_159,N_24673,N_24918);
nand UO_160 (O_160,N_24681,N_24801);
or UO_161 (O_161,N_24587,N_24968);
xor UO_162 (O_162,N_24815,N_24602);
xnor UO_163 (O_163,N_24726,N_24779);
nor UO_164 (O_164,N_24685,N_24618);
or UO_165 (O_165,N_24782,N_24723);
or UO_166 (O_166,N_24540,N_24852);
or UO_167 (O_167,N_24511,N_24583);
xnor UO_168 (O_168,N_24826,N_24663);
or UO_169 (O_169,N_24784,N_24536);
or UO_170 (O_170,N_24867,N_24955);
nor UO_171 (O_171,N_24933,N_24963);
and UO_172 (O_172,N_24985,N_24865);
or UO_173 (O_173,N_24742,N_24725);
or UO_174 (O_174,N_24600,N_24653);
nand UO_175 (O_175,N_24566,N_24607);
and UO_176 (O_176,N_24898,N_24554);
nand UO_177 (O_177,N_24712,N_24891);
and UO_178 (O_178,N_24957,N_24503);
or UO_179 (O_179,N_24652,N_24972);
nand UO_180 (O_180,N_24664,N_24911);
or UO_181 (O_181,N_24776,N_24643);
and UO_182 (O_182,N_24917,N_24616);
xnor UO_183 (O_183,N_24551,N_24902);
and UO_184 (O_184,N_24745,N_24879);
nor UO_185 (O_185,N_24605,N_24683);
nand UO_186 (O_186,N_24938,N_24580);
nand UO_187 (O_187,N_24868,N_24667);
nand UO_188 (O_188,N_24831,N_24961);
and UO_189 (O_189,N_24954,N_24990);
xnor UO_190 (O_190,N_24840,N_24792);
nor UO_191 (O_191,N_24966,N_24876);
nand UO_192 (O_192,N_24855,N_24939);
or UO_193 (O_193,N_24744,N_24790);
nor UO_194 (O_194,N_24546,N_24913);
xnor UO_195 (O_195,N_24510,N_24716);
and UO_196 (O_196,N_24617,N_24642);
nand UO_197 (O_197,N_24547,N_24950);
nor UO_198 (O_198,N_24977,N_24604);
xor UO_199 (O_199,N_24997,N_24502);
nand UO_200 (O_200,N_24861,N_24960);
or UO_201 (O_201,N_24910,N_24941);
and UO_202 (O_202,N_24592,N_24506);
nor UO_203 (O_203,N_24519,N_24701);
xor UO_204 (O_204,N_24746,N_24777);
xor UO_205 (O_205,N_24522,N_24808);
and UO_206 (O_206,N_24892,N_24542);
and UO_207 (O_207,N_24722,N_24995);
nand UO_208 (O_208,N_24662,N_24797);
or UO_209 (O_209,N_24696,N_24590);
nor UO_210 (O_210,N_24953,N_24905);
or UO_211 (O_211,N_24625,N_24773);
xnor UO_212 (O_212,N_24923,N_24531);
xor UO_213 (O_213,N_24752,N_24847);
or UO_214 (O_214,N_24505,N_24845);
or UO_215 (O_215,N_24636,N_24586);
and UO_216 (O_216,N_24562,N_24537);
nand UO_217 (O_217,N_24881,N_24538);
xnor UO_218 (O_218,N_24521,N_24634);
and UO_219 (O_219,N_24731,N_24760);
nand UO_220 (O_220,N_24693,N_24983);
or UO_221 (O_221,N_24944,N_24687);
nor UO_222 (O_222,N_24609,N_24578);
xnor UO_223 (O_223,N_24762,N_24549);
xor UO_224 (O_224,N_24651,N_24560);
xnor UO_225 (O_225,N_24558,N_24649);
or UO_226 (O_226,N_24820,N_24753);
or UO_227 (O_227,N_24940,N_24857);
nor UO_228 (O_228,N_24858,N_24711);
nand UO_229 (O_229,N_24789,N_24573);
and UO_230 (O_230,N_24767,N_24739);
nand UO_231 (O_231,N_24668,N_24645);
or UO_232 (O_232,N_24697,N_24764);
or UO_233 (O_233,N_24539,N_24936);
or UO_234 (O_234,N_24700,N_24993);
nand UO_235 (O_235,N_24572,N_24979);
or UO_236 (O_236,N_24964,N_24534);
nor UO_237 (O_237,N_24679,N_24628);
or UO_238 (O_238,N_24846,N_24800);
nand UO_239 (O_239,N_24830,N_24514);
nand UO_240 (O_240,N_24814,N_24588);
and UO_241 (O_241,N_24593,N_24631);
nand UO_242 (O_242,N_24924,N_24581);
xor UO_243 (O_243,N_24849,N_24895);
xor UO_244 (O_244,N_24992,N_24888);
or UO_245 (O_245,N_24556,N_24947);
and UO_246 (O_246,N_24730,N_24656);
and UO_247 (O_247,N_24582,N_24946);
and UO_248 (O_248,N_24787,N_24565);
xnor UO_249 (O_249,N_24682,N_24640);
and UO_250 (O_250,N_24517,N_24807);
nor UO_251 (O_251,N_24679,N_24939);
nor UO_252 (O_252,N_24805,N_24507);
xnor UO_253 (O_253,N_24843,N_24658);
and UO_254 (O_254,N_24969,N_24673);
or UO_255 (O_255,N_24780,N_24714);
or UO_256 (O_256,N_24839,N_24634);
nand UO_257 (O_257,N_24828,N_24883);
xor UO_258 (O_258,N_24695,N_24506);
or UO_259 (O_259,N_24774,N_24818);
or UO_260 (O_260,N_24718,N_24699);
xor UO_261 (O_261,N_24952,N_24507);
nor UO_262 (O_262,N_24878,N_24869);
nand UO_263 (O_263,N_24769,N_24726);
or UO_264 (O_264,N_24791,N_24573);
or UO_265 (O_265,N_24855,N_24886);
xor UO_266 (O_266,N_24715,N_24637);
xor UO_267 (O_267,N_24512,N_24595);
or UO_268 (O_268,N_24847,N_24917);
nand UO_269 (O_269,N_24587,N_24700);
xnor UO_270 (O_270,N_24838,N_24886);
nand UO_271 (O_271,N_24517,N_24522);
xor UO_272 (O_272,N_24616,N_24554);
xnor UO_273 (O_273,N_24854,N_24728);
xor UO_274 (O_274,N_24591,N_24653);
nand UO_275 (O_275,N_24642,N_24528);
or UO_276 (O_276,N_24547,N_24787);
nand UO_277 (O_277,N_24540,N_24660);
nor UO_278 (O_278,N_24865,N_24714);
nand UO_279 (O_279,N_24519,N_24667);
xnor UO_280 (O_280,N_24560,N_24500);
xnor UO_281 (O_281,N_24909,N_24701);
xor UO_282 (O_282,N_24823,N_24648);
nor UO_283 (O_283,N_24598,N_24945);
nor UO_284 (O_284,N_24791,N_24523);
nand UO_285 (O_285,N_24725,N_24529);
nand UO_286 (O_286,N_24508,N_24775);
xnor UO_287 (O_287,N_24871,N_24792);
or UO_288 (O_288,N_24528,N_24669);
nand UO_289 (O_289,N_24501,N_24900);
or UO_290 (O_290,N_24873,N_24745);
nand UO_291 (O_291,N_24752,N_24695);
nor UO_292 (O_292,N_24702,N_24523);
nor UO_293 (O_293,N_24966,N_24651);
or UO_294 (O_294,N_24609,N_24937);
and UO_295 (O_295,N_24635,N_24524);
nor UO_296 (O_296,N_24786,N_24773);
nor UO_297 (O_297,N_24824,N_24913);
or UO_298 (O_298,N_24983,N_24554);
nand UO_299 (O_299,N_24816,N_24609);
or UO_300 (O_300,N_24633,N_24587);
and UO_301 (O_301,N_24890,N_24545);
or UO_302 (O_302,N_24812,N_24700);
or UO_303 (O_303,N_24896,N_24941);
nand UO_304 (O_304,N_24998,N_24664);
and UO_305 (O_305,N_24503,N_24693);
xnor UO_306 (O_306,N_24636,N_24675);
and UO_307 (O_307,N_24514,N_24545);
nor UO_308 (O_308,N_24695,N_24562);
or UO_309 (O_309,N_24992,N_24909);
or UO_310 (O_310,N_24588,N_24779);
and UO_311 (O_311,N_24634,N_24609);
and UO_312 (O_312,N_24509,N_24685);
or UO_313 (O_313,N_24881,N_24708);
xor UO_314 (O_314,N_24846,N_24620);
and UO_315 (O_315,N_24995,N_24934);
or UO_316 (O_316,N_24846,N_24549);
xnor UO_317 (O_317,N_24751,N_24711);
and UO_318 (O_318,N_24703,N_24666);
nor UO_319 (O_319,N_24808,N_24807);
nor UO_320 (O_320,N_24544,N_24938);
xnor UO_321 (O_321,N_24875,N_24731);
or UO_322 (O_322,N_24936,N_24696);
or UO_323 (O_323,N_24754,N_24855);
nor UO_324 (O_324,N_24666,N_24626);
xor UO_325 (O_325,N_24697,N_24511);
and UO_326 (O_326,N_24985,N_24854);
and UO_327 (O_327,N_24829,N_24722);
nor UO_328 (O_328,N_24582,N_24870);
xor UO_329 (O_329,N_24669,N_24752);
nand UO_330 (O_330,N_24759,N_24995);
nand UO_331 (O_331,N_24702,N_24904);
and UO_332 (O_332,N_24995,N_24694);
nand UO_333 (O_333,N_24616,N_24719);
and UO_334 (O_334,N_24527,N_24622);
nor UO_335 (O_335,N_24698,N_24612);
or UO_336 (O_336,N_24930,N_24621);
nor UO_337 (O_337,N_24530,N_24801);
nor UO_338 (O_338,N_24535,N_24729);
nand UO_339 (O_339,N_24848,N_24758);
nand UO_340 (O_340,N_24800,N_24878);
xor UO_341 (O_341,N_24925,N_24508);
nor UO_342 (O_342,N_24947,N_24868);
nor UO_343 (O_343,N_24820,N_24963);
and UO_344 (O_344,N_24650,N_24544);
and UO_345 (O_345,N_24992,N_24522);
nand UO_346 (O_346,N_24614,N_24791);
and UO_347 (O_347,N_24856,N_24603);
or UO_348 (O_348,N_24889,N_24502);
and UO_349 (O_349,N_24800,N_24986);
nand UO_350 (O_350,N_24726,N_24535);
and UO_351 (O_351,N_24952,N_24942);
nand UO_352 (O_352,N_24612,N_24961);
nor UO_353 (O_353,N_24501,N_24783);
or UO_354 (O_354,N_24826,N_24682);
xnor UO_355 (O_355,N_24728,N_24664);
and UO_356 (O_356,N_24858,N_24972);
nand UO_357 (O_357,N_24746,N_24533);
or UO_358 (O_358,N_24744,N_24524);
or UO_359 (O_359,N_24527,N_24957);
nand UO_360 (O_360,N_24616,N_24926);
nor UO_361 (O_361,N_24818,N_24990);
and UO_362 (O_362,N_24607,N_24624);
xor UO_363 (O_363,N_24889,N_24862);
and UO_364 (O_364,N_24706,N_24939);
nand UO_365 (O_365,N_24785,N_24775);
xor UO_366 (O_366,N_24531,N_24659);
nand UO_367 (O_367,N_24832,N_24754);
xor UO_368 (O_368,N_24719,N_24658);
xnor UO_369 (O_369,N_24782,N_24501);
or UO_370 (O_370,N_24682,N_24877);
xor UO_371 (O_371,N_24659,N_24708);
nand UO_372 (O_372,N_24783,N_24716);
nor UO_373 (O_373,N_24963,N_24804);
nand UO_374 (O_374,N_24610,N_24767);
and UO_375 (O_375,N_24571,N_24551);
and UO_376 (O_376,N_24701,N_24566);
nor UO_377 (O_377,N_24676,N_24602);
and UO_378 (O_378,N_24584,N_24514);
nand UO_379 (O_379,N_24789,N_24506);
and UO_380 (O_380,N_24756,N_24525);
nor UO_381 (O_381,N_24909,N_24873);
or UO_382 (O_382,N_24866,N_24880);
or UO_383 (O_383,N_24952,N_24726);
and UO_384 (O_384,N_24596,N_24983);
and UO_385 (O_385,N_24525,N_24501);
or UO_386 (O_386,N_24816,N_24706);
or UO_387 (O_387,N_24806,N_24735);
or UO_388 (O_388,N_24582,N_24544);
nand UO_389 (O_389,N_24678,N_24703);
xnor UO_390 (O_390,N_24996,N_24978);
and UO_391 (O_391,N_24815,N_24832);
or UO_392 (O_392,N_24668,N_24944);
nor UO_393 (O_393,N_24841,N_24844);
nor UO_394 (O_394,N_24636,N_24602);
xnor UO_395 (O_395,N_24776,N_24733);
xor UO_396 (O_396,N_24877,N_24645);
or UO_397 (O_397,N_24758,N_24942);
and UO_398 (O_398,N_24500,N_24762);
or UO_399 (O_399,N_24612,N_24609);
and UO_400 (O_400,N_24600,N_24867);
xor UO_401 (O_401,N_24538,N_24765);
and UO_402 (O_402,N_24876,N_24812);
xor UO_403 (O_403,N_24603,N_24979);
xor UO_404 (O_404,N_24744,N_24976);
or UO_405 (O_405,N_24705,N_24762);
nand UO_406 (O_406,N_24525,N_24785);
nand UO_407 (O_407,N_24940,N_24898);
nand UO_408 (O_408,N_24924,N_24670);
or UO_409 (O_409,N_24624,N_24657);
or UO_410 (O_410,N_24982,N_24866);
xor UO_411 (O_411,N_24578,N_24660);
and UO_412 (O_412,N_24668,N_24833);
and UO_413 (O_413,N_24857,N_24616);
xnor UO_414 (O_414,N_24770,N_24739);
nand UO_415 (O_415,N_24733,N_24523);
and UO_416 (O_416,N_24968,N_24617);
nand UO_417 (O_417,N_24604,N_24708);
nand UO_418 (O_418,N_24966,N_24806);
xor UO_419 (O_419,N_24912,N_24588);
and UO_420 (O_420,N_24758,N_24944);
xor UO_421 (O_421,N_24500,N_24958);
and UO_422 (O_422,N_24616,N_24788);
nand UO_423 (O_423,N_24864,N_24779);
nand UO_424 (O_424,N_24776,N_24716);
or UO_425 (O_425,N_24756,N_24719);
xnor UO_426 (O_426,N_24927,N_24683);
nor UO_427 (O_427,N_24729,N_24964);
nor UO_428 (O_428,N_24539,N_24949);
nand UO_429 (O_429,N_24664,N_24995);
and UO_430 (O_430,N_24581,N_24785);
xor UO_431 (O_431,N_24601,N_24691);
xor UO_432 (O_432,N_24900,N_24801);
or UO_433 (O_433,N_24558,N_24802);
nand UO_434 (O_434,N_24848,N_24627);
or UO_435 (O_435,N_24830,N_24918);
nor UO_436 (O_436,N_24864,N_24875);
and UO_437 (O_437,N_24688,N_24712);
or UO_438 (O_438,N_24576,N_24570);
and UO_439 (O_439,N_24738,N_24653);
xor UO_440 (O_440,N_24767,N_24846);
nand UO_441 (O_441,N_24922,N_24684);
xor UO_442 (O_442,N_24615,N_24789);
and UO_443 (O_443,N_24702,N_24874);
xor UO_444 (O_444,N_24541,N_24878);
nand UO_445 (O_445,N_24581,N_24932);
nor UO_446 (O_446,N_24856,N_24804);
xor UO_447 (O_447,N_24774,N_24938);
nor UO_448 (O_448,N_24911,N_24854);
nor UO_449 (O_449,N_24990,N_24709);
and UO_450 (O_450,N_24959,N_24641);
nor UO_451 (O_451,N_24992,N_24816);
nand UO_452 (O_452,N_24847,N_24699);
xor UO_453 (O_453,N_24617,N_24786);
and UO_454 (O_454,N_24811,N_24622);
and UO_455 (O_455,N_24537,N_24704);
xnor UO_456 (O_456,N_24716,N_24587);
nor UO_457 (O_457,N_24519,N_24935);
and UO_458 (O_458,N_24978,N_24612);
nand UO_459 (O_459,N_24751,N_24929);
nand UO_460 (O_460,N_24830,N_24615);
or UO_461 (O_461,N_24860,N_24955);
nand UO_462 (O_462,N_24862,N_24738);
or UO_463 (O_463,N_24820,N_24586);
nand UO_464 (O_464,N_24856,N_24752);
nor UO_465 (O_465,N_24951,N_24723);
nand UO_466 (O_466,N_24623,N_24534);
xnor UO_467 (O_467,N_24516,N_24708);
nand UO_468 (O_468,N_24776,N_24925);
nand UO_469 (O_469,N_24589,N_24532);
or UO_470 (O_470,N_24677,N_24739);
or UO_471 (O_471,N_24728,N_24935);
and UO_472 (O_472,N_24686,N_24571);
and UO_473 (O_473,N_24959,N_24953);
nor UO_474 (O_474,N_24835,N_24748);
xnor UO_475 (O_475,N_24670,N_24867);
xor UO_476 (O_476,N_24879,N_24599);
nor UO_477 (O_477,N_24627,N_24810);
and UO_478 (O_478,N_24681,N_24726);
xor UO_479 (O_479,N_24876,N_24597);
nor UO_480 (O_480,N_24829,N_24852);
or UO_481 (O_481,N_24539,N_24959);
xor UO_482 (O_482,N_24519,N_24605);
nor UO_483 (O_483,N_24504,N_24801);
nor UO_484 (O_484,N_24647,N_24791);
or UO_485 (O_485,N_24959,N_24517);
nand UO_486 (O_486,N_24972,N_24892);
or UO_487 (O_487,N_24940,N_24829);
nand UO_488 (O_488,N_24849,N_24650);
nor UO_489 (O_489,N_24741,N_24997);
nand UO_490 (O_490,N_24875,N_24714);
and UO_491 (O_491,N_24592,N_24708);
or UO_492 (O_492,N_24796,N_24798);
xor UO_493 (O_493,N_24606,N_24788);
xnor UO_494 (O_494,N_24567,N_24833);
nor UO_495 (O_495,N_24726,N_24733);
or UO_496 (O_496,N_24604,N_24655);
nand UO_497 (O_497,N_24801,N_24673);
nor UO_498 (O_498,N_24765,N_24715);
nor UO_499 (O_499,N_24988,N_24934);
nand UO_500 (O_500,N_24503,N_24622);
nand UO_501 (O_501,N_24596,N_24554);
nand UO_502 (O_502,N_24787,N_24642);
nor UO_503 (O_503,N_24823,N_24595);
and UO_504 (O_504,N_24531,N_24905);
or UO_505 (O_505,N_24693,N_24650);
nand UO_506 (O_506,N_24594,N_24901);
xor UO_507 (O_507,N_24661,N_24504);
or UO_508 (O_508,N_24849,N_24743);
nand UO_509 (O_509,N_24623,N_24894);
nor UO_510 (O_510,N_24732,N_24541);
nand UO_511 (O_511,N_24846,N_24902);
nand UO_512 (O_512,N_24724,N_24657);
nand UO_513 (O_513,N_24573,N_24851);
nor UO_514 (O_514,N_24698,N_24561);
and UO_515 (O_515,N_24764,N_24873);
nor UO_516 (O_516,N_24618,N_24731);
nand UO_517 (O_517,N_24716,N_24755);
nand UO_518 (O_518,N_24856,N_24556);
xor UO_519 (O_519,N_24944,N_24922);
xor UO_520 (O_520,N_24678,N_24835);
nand UO_521 (O_521,N_24806,N_24775);
and UO_522 (O_522,N_24507,N_24940);
and UO_523 (O_523,N_24824,N_24517);
nor UO_524 (O_524,N_24555,N_24895);
nand UO_525 (O_525,N_24936,N_24597);
nor UO_526 (O_526,N_24557,N_24754);
nand UO_527 (O_527,N_24847,N_24745);
xor UO_528 (O_528,N_24905,N_24666);
nor UO_529 (O_529,N_24835,N_24656);
nand UO_530 (O_530,N_24736,N_24914);
nor UO_531 (O_531,N_24888,N_24832);
or UO_532 (O_532,N_24726,N_24855);
xnor UO_533 (O_533,N_24915,N_24932);
nor UO_534 (O_534,N_24872,N_24784);
nand UO_535 (O_535,N_24715,N_24514);
nor UO_536 (O_536,N_24703,N_24679);
xor UO_537 (O_537,N_24752,N_24861);
or UO_538 (O_538,N_24851,N_24965);
nor UO_539 (O_539,N_24996,N_24942);
nand UO_540 (O_540,N_24809,N_24912);
or UO_541 (O_541,N_24774,N_24604);
nand UO_542 (O_542,N_24894,N_24728);
xnor UO_543 (O_543,N_24637,N_24767);
or UO_544 (O_544,N_24887,N_24679);
and UO_545 (O_545,N_24758,N_24896);
or UO_546 (O_546,N_24702,N_24891);
nor UO_547 (O_547,N_24614,N_24572);
xor UO_548 (O_548,N_24648,N_24833);
nand UO_549 (O_549,N_24795,N_24586);
or UO_550 (O_550,N_24635,N_24548);
nor UO_551 (O_551,N_24885,N_24519);
xor UO_552 (O_552,N_24628,N_24785);
nor UO_553 (O_553,N_24500,N_24550);
or UO_554 (O_554,N_24646,N_24815);
nor UO_555 (O_555,N_24659,N_24632);
nor UO_556 (O_556,N_24610,N_24929);
nor UO_557 (O_557,N_24821,N_24515);
and UO_558 (O_558,N_24835,N_24618);
nor UO_559 (O_559,N_24678,N_24984);
or UO_560 (O_560,N_24984,N_24822);
nand UO_561 (O_561,N_24571,N_24848);
nand UO_562 (O_562,N_24586,N_24854);
and UO_563 (O_563,N_24502,N_24711);
xnor UO_564 (O_564,N_24559,N_24821);
nor UO_565 (O_565,N_24672,N_24847);
nand UO_566 (O_566,N_24892,N_24646);
nor UO_567 (O_567,N_24837,N_24569);
nor UO_568 (O_568,N_24612,N_24696);
xnor UO_569 (O_569,N_24868,N_24723);
xor UO_570 (O_570,N_24750,N_24647);
or UO_571 (O_571,N_24889,N_24603);
nor UO_572 (O_572,N_24517,N_24540);
or UO_573 (O_573,N_24689,N_24927);
xnor UO_574 (O_574,N_24611,N_24579);
or UO_575 (O_575,N_24684,N_24593);
nand UO_576 (O_576,N_24837,N_24744);
nor UO_577 (O_577,N_24718,N_24607);
nand UO_578 (O_578,N_24680,N_24568);
and UO_579 (O_579,N_24950,N_24801);
or UO_580 (O_580,N_24887,N_24805);
nor UO_581 (O_581,N_24852,N_24989);
xnor UO_582 (O_582,N_24821,N_24842);
and UO_583 (O_583,N_24739,N_24890);
nand UO_584 (O_584,N_24512,N_24770);
or UO_585 (O_585,N_24510,N_24847);
xnor UO_586 (O_586,N_24993,N_24904);
xnor UO_587 (O_587,N_24710,N_24953);
or UO_588 (O_588,N_24949,N_24606);
nand UO_589 (O_589,N_24811,N_24685);
nor UO_590 (O_590,N_24986,N_24948);
or UO_591 (O_591,N_24657,N_24555);
or UO_592 (O_592,N_24692,N_24578);
nor UO_593 (O_593,N_24919,N_24753);
nor UO_594 (O_594,N_24730,N_24729);
and UO_595 (O_595,N_24734,N_24975);
nor UO_596 (O_596,N_24596,N_24728);
and UO_597 (O_597,N_24647,N_24510);
xor UO_598 (O_598,N_24703,N_24921);
and UO_599 (O_599,N_24629,N_24837);
and UO_600 (O_600,N_24508,N_24872);
and UO_601 (O_601,N_24667,N_24840);
or UO_602 (O_602,N_24570,N_24954);
and UO_603 (O_603,N_24870,N_24556);
xnor UO_604 (O_604,N_24730,N_24890);
or UO_605 (O_605,N_24527,N_24580);
or UO_606 (O_606,N_24776,N_24954);
or UO_607 (O_607,N_24711,N_24745);
and UO_608 (O_608,N_24935,N_24831);
nand UO_609 (O_609,N_24935,N_24752);
or UO_610 (O_610,N_24925,N_24920);
nor UO_611 (O_611,N_24652,N_24668);
xnor UO_612 (O_612,N_24860,N_24505);
nand UO_613 (O_613,N_24908,N_24925);
xnor UO_614 (O_614,N_24508,N_24674);
xnor UO_615 (O_615,N_24695,N_24545);
nand UO_616 (O_616,N_24769,N_24893);
nor UO_617 (O_617,N_24692,N_24812);
nand UO_618 (O_618,N_24748,N_24875);
or UO_619 (O_619,N_24834,N_24611);
or UO_620 (O_620,N_24663,N_24918);
nand UO_621 (O_621,N_24509,N_24862);
or UO_622 (O_622,N_24514,N_24880);
nand UO_623 (O_623,N_24531,N_24581);
xor UO_624 (O_624,N_24975,N_24781);
nand UO_625 (O_625,N_24727,N_24760);
xor UO_626 (O_626,N_24887,N_24754);
xor UO_627 (O_627,N_24939,N_24540);
xnor UO_628 (O_628,N_24575,N_24879);
and UO_629 (O_629,N_24790,N_24754);
nand UO_630 (O_630,N_24611,N_24701);
nor UO_631 (O_631,N_24622,N_24845);
nor UO_632 (O_632,N_24644,N_24610);
and UO_633 (O_633,N_24755,N_24692);
nor UO_634 (O_634,N_24726,N_24962);
nor UO_635 (O_635,N_24789,N_24530);
and UO_636 (O_636,N_24865,N_24746);
or UO_637 (O_637,N_24572,N_24719);
xnor UO_638 (O_638,N_24576,N_24642);
and UO_639 (O_639,N_24863,N_24925);
or UO_640 (O_640,N_24679,N_24503);
nand UO_641 (O_641,N_24802,N_24637);
xnor UO_642 (O_642,N_24987,N_24910);
and UO_643 (O_643,N_24784,N_24822);
and UO_644 (O_644,N_24523,N_24967);
or UO_645 (O_645,N_24689,N_24645);
xnor UO_646 (O_646,N_24612,N_24932);
nor UO_647 (O_647,N_24607,N_24536);
nor UO_648 (O_648,N_24519,N_24704);
and UO_649 (O_649,N_24872,N_24598);
or UO_650 (O_650,N_24552,N_24798);
or UO_651 (O_651,N_24973,N_24904);
nand UO_652 (O_652,N_24741,N_24762);
and UO_653 (O_653,N_24526,N_24736);
or UO_654 (O_654,N_24788,N_24999);
nand UO_655 (O_655,N_24670,N_24953);
nor UO_656 (O_656,N_24541,N_24909);
or UO_657 (O_657,N_24951,N_24640);
nand UO_658 (O_658,N_24535,N_24788);
and UO_659 (O_659,N_24622,N_24848);
xnor UO_660 (O_660,N_24645,N_24814);
or UO_661 (O_661,N_24754,N_24515);
nor UO_662 (O_662,N_24748,N_24785);
or UO_663 (O_663,N_24989,N_24926);
nor UO_664 (O_664,N_24772,N_24710);
and UO_665 (O_665,N_24575,N_24641);
and UO_666 (O_666,N_24558,N_24766);
nor UO_667 (O_667,N_24900,N_24950);
xor UO_668 (O_668,N_24965,N_24669);
nand UO_669 (O_669,N_24836,N_24706);
xnor UO_670 (O_670,N_24569,N_24898);
and UO_671 (O_671,N_24612,N_24522);
nor UO_672 (O_672,N_24906,N_24950);
and UO_673 (O_673,N_24955,N_24774);
or UO_674 (O_674,N_24842,N_24585);
and UO_675 (O_675,N_24754,N_24615);
or UO_676 (O_676,N_24555,N_24517);
xnor UO_677 (O_677,N_24675,N_24888);
nor UO_678 (O_678,N_24889,N_24826);
nor UO_679 (O_679,N_24546,N_24543);
and UO_680 (O_680,N_24743,N_24673);
and UO_681 (O_681,N_24627,N_24696);
or UO_682 (O_682,N_24850,N_24906);
nor UO_683 (O_683,N_24769,N_24995);
nor UO_684 (O_684,N_24876,N_24932);
and UO_685 (O_685,N_24813,N_24906);
or UO_686 (O_686,N_24678,N_24873);
nor UO_687 (O_687,N_24513,N_24949);
or UO_688 (O_688,N_24698,N_24845);
and UO_689 (O_689,N_24905,N_24717);
and UO_690 (O_690,N_24883,N_24831);
or UO_691 (O_691,N_24723,N_24506);
nand UO_692 (O_692,N_24855,N_24526);
xnor UO_693 (O_693,N_24563,N_24520);
xnor UO_694 (O_694,N_24749,N_24855);
xnor UO_695 (O_695,N_24549,N_24635);
nand UO_696 (O_696,N_24768,N_24757);
or UO_697 (O_697,N_24660,N_24536);
and UO_698 (O_698,N_24942,N_24626);
nor UO_699 (O_699,N_24573,N_24765);
xor UO_700 (O_700,N_24809,N_24823);
nand UO_701 (O_701,N_24786,N_24729);
nor UO_702 (O_702,N_24527,N_24558);
xor UO_703 (O_703,N_24525,N_24993);
and UO_704 (O_704,N_24587,N_24563);
or UO_705 (O_705,N_24546,N_24695);
or UO_706 (O_706,N_24619,N_24747);
nor UO_707 (O_707,N_24539,N_24892);
xnor UO_708 (O_708,N_24694,N_24732);
nand UO_709 (O_709,N_24946,N_24627);
or UO_710 (O_710,N_24983,N_24986);
nor UO_711 (O_711,N_24504,N_24656);
and UO_712 (O_712,N_24523,N_24925);
and UO_713 (O_713,N_24971,N_24998);
nand UO_714 (O_714,N_24630,N_24807);
and UO_715 (O_715,N_24651,N_24829);
nor UO_716 (O_716,N_24792,N_24735);
nand UO_717 (O_717,N_24529,N_24953);
nor UO_718 (O_718,N_24932,N_24703);
and UO_719 (O_719,N_24875,N_24781);
xnor UO_720 (O_720,N_24924,N_24777);
and UO_721 (O_721,N_24964,N_24553);
or UO_722 (O_722,N_24686,N_24815);
or UO_723 (O_723,N_24557,N_24567);
xnor UO_724 (O_724,N_24758,N_24658);
and UO_725 (O_725,N_24535,N_24964);
nand UO_726 (O_726,N_24722,N_24841);
nand UO_727 (O_727,N_24837,N_24768);
and UO_728 (O_728,N_24559,N_24857);
nand UO_729 (O_729,N_24567,N_24617);
nand UO_730 (O_730,N_24646,N_24949);
xor UO_731 (O_731,N_24808,N_24536);
nor UO_732 (O_732,N_24922,N_24659);
xnor UO_733 (O_733,N_24788,N_24532);
or UO_734 (O_734,N_24951,N_24828);
nor UO_735 (O_735,N_24974,N_24741);
nand UO_736 (O_736,N_24657,N_24924);
and UO_737 (O_737,N_24599,N_24845);
nand UO_738 (O_738,N_24877,N_24820);
nand UO_739 (O_739,N_24731,N_24820);
nor UO_740 (O_740,N_24724,N_24637);
nor UO_741 (O_741,N_24676,N_24881);
and UO_742 (O_742,N_24679,N_24748);
and UO_743 (O_743,N_24518,N_24663);
xnor UO_744 (O_744,N_24703,N_24657);
nand UO_745 (O_745,N_24791,N_24561);
and UO_746 (O_746,N_24978,N_24678);
xor UO_747 (O_747,N_24537,N_24663);
and UO_748 (O_748,N_24613,N_24803);
nor UO_749 (O_749,N_24576,N_24560);
or UO_750 (O_750,N_24893,N_24808);
nor UO_751 (O_751,N_24515,N_24506);
xor UO_752 (O_752,N_24567,N_24934);
or UO_753 (O_753,N_24547,N_24540);
nor UO_754 (O_754,N_24730,N_24557);
or UO_755 (O_755,N_24540,N_24614);
xnor UO_756 (O_756,N_24976,N_24603);
nor UO_757 (O_757,N_24848,N_24945);
nor UO_758 (O_758,N_24500,N_24870);
nand UO_759 (O_759,N_24597,N_24966);
and UO_760 (O_760,N_24779,N_24711);
or UO_761 (O_761,N_24586,N_24748);
nand UO_762 (O_762,N_24791,N_24628);
nand UO_763 (O_763,N_24698,N_24575);
nor UO_764 (O_764,N_24808,N_24568);
or UO_765 (O_765,N_24530,N_24537);
and UO_766 (O_766,N_24825,N_24527);
or UO_767 (O_767,N_24506,N_24645);
nand UO_768 (O_768,N_24782,N_24930);
nor UO_769 (O_769,N_24606,N_24572);
and UO_770 (O_770,N_24592,N_24872);
or UO_771 (O_771,N_24892,N_24872);
nand UO_772 (O_772,N_24803,N_24812);
or UO_773 (O_773,N_24575,N_24876);
or UO_774 (O_774,N_24631,N_24551);
or UO_775 (O_775,N_24656,N_24716);
or UO_776 (O_776,N_24797,N_24559);
nand UO_777 (O_777,N_24705,N_24996);
nand UO_778 (O_778,N_24580,N_24855);
nand UO_779 (O_779,N_24929,N_24694);
xnor UO_780 (O_780,N_24672,N_24985);
and UO_781 (O_781,N_24920,N_24519);
xnor UO_782 (O_782,N_24969,N_24903);
and UO_783 (O_783,N_24828,N_24867);
nor UO_784 (O_784,N_24703,N_24872);
and UO_785 (O_785,N_24922,N_24637);
nor UO_786 (O_786,N_24935,N_24648);
xnor UO_787 (O_787,N_24976,N_24927);
and UO_788 (O_788,N_24547,N_24800);
xor UO_789 (O_789,N_24534,N_24785);
nor UO_790 (O_790,N_24730,N_24680);
xnor UO_791 (O_791,N_24672,N_24892);
nor UO_792 (O_792,N_24916,N_24539);
or UO_793 (O_793,N_24596,N_24681);
and UO_794 (O_794,N_24832,N_24958);
xnor UO_795 (O_795,N_24562,N_24603);
xnor UO_796 (O_796,N_24889,N_24994);
xor UO_797 (O_797,N_24858,N_24701);
or UO_798 (O_798,N_24765,N_24529);
nand UO_799 (O_799,N_24837,N_24957);
nand UO_800 (O_800,N_24708,N_24837);
nor UO_801 (O_801,N_24901,N_24880);
nor UO_802 (O_802,N_24611,N_24572);
and UO_803 (O_803,N_24811,N_24894);
or UO_804 (O_804,N_24979,N_24926);
nor UO_805 (O_805,N_24679,N_24865);
and UO_806 (O_806,N_24916,N_24805);
and UO_807 (O_807,N_24746,N_24907);
nand UO_808 (O_808,N_24523,N_24811);
or UO_809 (O_809,N_24536,N_24920);
xnor UO_810 (O_810,N_24544,N_24623);
nor UO_811 (O_811,N_24548,N_24633);
xor UO_812 (O_812,N_24646,N_24630);
xor UO_813 (O_813,N_24938,N_24915);
or UO_814 (O_814,N_24673,N_24966);
or UO_815 (O_815,N_24716,N_24629);
nand UO_816 (O_816,N_24850,N_24976);
nand UO_817 (O_817,N_24907,N_24906);
nand UO_818 (O_818,N_24728,N_24739);
or UO_819 (O_819,N_24574,N_24565);
xor UO_820 (O_820,N_24716,N_24704);
and UO_821 (O_821,N_24979,N_24884);
nand UO_822 (O_822,N_24741,N_24835);
or UO_823 (O_823,N_24577,N_24715);
or UO_824 (O_824,N_24719,N_24913);
nand UO_825 (O_825,N_24744,N_24690);
nor UO_826 (O_826,N_24724,N_24834);
nor UO_827 (O_827,N_24906,N_24840);
and UO_828 (O_828,N_24761,N_24918);
or UO_829 (O_829,N_24897,N_24553);
and UO_830 (O_830,N_24865,N_24859);
xnor UO_831 (O_831,N_24673,N_24636);
xnor UO_832 (O_832,N_24865,N_24526);
nand UO_833 (O_833,N_24893,N_24778);
xor UO_834 (O_834,N_24536,N_24597);
xnor UO_835 (O_835,N_24913,N_24933);
nor UO_836 (O_836,N_24719,N_24535);
and UO_837 (O_837,N_24884,N_24831);
nand UO_838 (O_838,N_24880,N_24615);
nor UO_839 (O_839,N_24852,N_24796);
and UO_840 (O_840,N_24843,N_24759);
or UO_841 (O_841,N_24795,N_24851);
nand UO_842 (O_842,N_24757,N_24520);
nand UO_843 (O_843,N_24743,N_24556);
xor UO_844 (O_844,N_24865,N_24641);
and UO_845 (O_845,N_24615,N_24979);
or UO_846 (O_846,N_24648,N_24507);
xnor UO_847 (O_847,N_24719,N_24721);
nand UO_848 (O_848,N_24632,N_24982);
nand UO_849 (O_849,N_24791,N_24751);
xnor UO_850 (O_850,N_24633,N_24918);
nor UO_851 (O_851,N_24872,N_24710);
xnor UO_852 (O_852,N_24712,N_24634);
or UO_853 (O_853,N_24731,N_24556);
nor UO_854 (O_854,N_24961,N_24705);
xor UO_855 (O_855,N_24846,N_24944);
xnor UO_856 (O_856,N_24992,N_24838);
or UO_857 (O_857,N_24744,N_24525);
and UO_858 (O_858,N_24543,N_24848);
and UO_859 (O_859,N_24691,N_24774);
nor UO_860 (O_860,N_24646,N_24739);
nor UO_861 (O_861,N_24632,N_24898);
nand UO_862 (O_862,N_24607,N_24744);
nand UO_863 (O_863,N_24686,N_24735);
xor UO_864 (O_864,N_24687,N_24522);
nand UO_865 (O_865,N_24986,N_24657);
nor UO_866 (O_866,N_24901,N_24721);
or UO_867 (O_867,N_24851,N_24866);
and UO_868 (O_868,N_24633,N_24691);
nor UO_869 (O_869,N_24519,N_24689);
or UO_870 (O_870,N_24617,N_24627);
and UO_871 (O_871,N_24518,N_24921);
or UO_872 (O_872,N_24745,N_24625);
nor UO_873 (O_873,N_24724,N_24964);
nor UO_874 (O_874,N_24635,N_24822);
or UO_875 (O_875,N_24965,N_24786);
xor UO_876 (O_876,N_24557,N_24550);
or UO_877 (O_877,N_24629,N_24798);
nand UO_878 (O_878,N_24778,N_24516);
and UO_879 (O_879,N_24740,N_24982);
or UO_880 (O_880,N_24623,N_24969);
or UO_881 (O_881,N_24928,N_24702);
nand UO_882 (O_882,N_24780,N_24697);
and UO_883 (O_883,N_24622,N_24500);
and UO_884 (O_884,N_24714,N_24595);
and UO_885 (O_885,N_24641,N_24716);
or UO_886 (O_886,N_24563,N_24857);
or UO_887 (O_887,N_24838,N_24981);
nand UO_888 (O_888,N_24588,N_24942);
or UO_889 (O_889,N_24559,N_24673);
nand UO_890 (O_890,N_24535,N_24908);
xnor UO_891 (O_891,N_24504,N_24567);
nand UO_892 (O_892,N_24992,N_24554);
and UO_893 (O_893,N_24935,N_24534);
nand UO_894 (O_894,N_24666,N_24545);
xnor UO_895 (O_895,N_24558,N_24569);
nor UO_896 (O_896,N_24910,N_24701);
nand UO_897 (O_897,N_24518,N_24697);
xnor UO_898 (O_898,N_24698,N_24863);
xor UO_899 (O_899,N_24606,N_24903);
nand UO_900 (O_900,N_24758,N_24647);
and UO_901 (O_901,N_24682,N_24624);
nor UO_902 (O_902,N_24922,N_24832);
nor UO_903 (O_903,N_24570,N_24955);
xnor UO_904 (O_904,N_24727,N_24552);
nor UO_905 (O_905,N_24959,N_24642);
nand UO_906 (O_906,N_24798,N_24737);
xor UO_907 (O_907,N_24874,N_24746);
xor UO_908 (O_908,N_24598,N_24558);
nor UO_909 (O_909,N_24718,N_24584);
xor UO_910 (O_910,N_24815,N_24714);
xor UO_911 (O_911,N_24835,N_24653);
nand UO_912 (O_912,N_24914,N_24761);
xor UO_913 (O_913,N_24997,N_24980);
nor UO_914 (O_914,N_24591,N_24651);
nand UO_915 (O_915,N_24521,N_24699);
xnor UO_916 (O_916,N_24985,N_24671);
nor UO_917 (O_917,N_24919,N_24509);
xor UO_918 (O_918,N_24991,N_24610);
and UO_919 (O_919,N_24508,N_24614);
nor UO_920 (O_920,N_24829,N_24996);
and UO_921 (O_921,N_24837,N_24646);
and UO_922 (O_922,N_24552,N_24566);
nand UO_923 (O_923,N_24866,N_24983);
xor UO_924 (O_924,N_24776,N_24931);
or UO_925 (O_925,N_24848,N_24878);
and UO_926 (O_926,N_24799,N_24719);
or UO_927 (O_927,N_24604,N_24761);
nand UO_928 (O_928,N_24834,N_24635);
and UO_929 (O_929,N_24784,N_24578);
or UO_930 (O_930,N_24912,N_24810);
xor UO_931 (O_931,N_24892,N_24947);
and UO_932 (O_932,N_24747,N_24882);
nor UO_933 (O_933,N_24518,N_24767);
or UO_934 (O_934,N_24638,N_24616);
nand UO_935 (O_935,N_24993,N_24959);
and UO_936 (O_936,N_24521,N_24696);
nand UO_937 (O_937,N_24991,N_24556);
and UO_938 (O_938,N_24943,N_24514);
or UO_939 (O_939,N_24672,N_24648);
or UO_940 (O_940,N_24841,N_24832);
nor UO_941 (O_941,N_24586,N_24617);
nand UO_942 (O_942,N_24713,N_24629);
xnor UO_943 (O_943,N_24952,N_24609);
xor UO_944 (O_944,N_24769,N_24993);
or UO_945 (O_945,N_24891,N_24850);
nand UO_946 (O_946,N_24644,N_24586);
or UO_947 (O_947,N_24841,N_24501);
xnor UO_948 (O_948,N_24984,N_24583);
and UO_949 (O_949,N_24854,N_24626);
or UO_950 (O_950,N_24873,N_24731);
nand UO_951 (O_951,N_24500,N_24841);
or UO_952 (O_952,N_24519,N_24786);
and UO_953 (O_953,N_24877,N_24846);
nand UO_954 (O_954,N_24781,N_24712);
and UO_955 (O_955,N_24585,N_24970);
nor UO_956 (O_956,N_24743,N_24933);
nor UO_957 (O_957,N_24806,N_24804);
and UO_958 (O_958,N_24679,N_24948);
nand UO_959 (O_959,N_24996,N_24694);
nand UO_960 (O_960,N_24789,N_24756);
xnor UO_961 (O_961,N_24596,N_24769);
nand UO_962 (O_962,N_24525,N_24896);
or UO_963 (O_963,N_24797,N_24861);
and UO_964 (O_964,N_24890,N_24878);
nor UO_965 (O_965,N_24779,N_24942);
and UO_966 (O_966,N_24568,N_24905);
and UO_967 (O_967,N_24894,N_24775);
nor UO_968 (O_968,N_24514,N_24908);
and UO_969 (O_969,N_24795,N_24824);
nor UO_970 (O_970,N_24697,N_24991);
nor UO_971 (O_971,N_24604,N_24728);
and UO_972 (O_972,N_24854,N_24666);
or UO_973 (O_973,N_24580,N_24990);
or UO_974 (O_974,N_24664,N_24948);
xnor UO_975 (O_975,N_24855,N_24782);
xor UO_976 (O_976,N_24936,N_24831);
or UO_977 (O_977,N_24555,N_24904);
and UO_978 (O_978,N_24928,N_24550);
or UO_979 (O_979,N_24645,N_24951);
or UO_980 (O_980,N_24580,N_24507);
xor UO_981 (O_981,N_24612,N_24558);
nand UO_982 (O_982,N_24931,N_24834);
or UO_983 (O_983,N_24515,N_24768);
or UO_984 (O_984,N_24770,N_24640);
or UO_985 (O_985,N_24629,N_24779);
or UO_986 (O_986,N_24983,N_24960);
or UO_987 (O_987,N_24911,N_24653);
nand UO_988 (O_988,N_24509,N_24547);
xnor UO_989 (O_989,N_24586,N_24988);
nor UO_990 (O_990,N_24629,N_24760);
and UO_991 (O_991,N_24675,N_24633);
and UO_992 (O_992,N_24913,N_24748);
or UO_993 (O_993,N_24646,N_24546);
nor UO_994 (O_994,N_24882,N_24746);
nand UO_995 (O_995,N_24934,N_24907);
or UO_996 (O_996,N_24710,N_24898);
and UO_997 (O_997,N_24796,N_24884);
xor UO_998 (O_998,N_24656,N_24771);
xnor UO_999 (O_999,N_24772,N_24899);
xor UO_1000 (O_1000,N_24655,N_24974);
xnor UO_1001 (O_1001,N_24555,N_24675);
nand UO_1002 (O_1002,N_24862,N_24711);
nor UO_1003 (O_1003,N_24846,N_24597);
xnor UO_1004 (O_1004,N_24867,N_24626);
or UO_1005 (O_1005,N_24568,N_24980);
and UO_1006 (O_1006,N_24704,N_24712);
or UO_1007 (O_1007,N_24963,N_24864);
xor UO_1008 (O_1008,N_24636,N_24671);
xnor UO_1009 (O_1009,N_24508,N_24860);
nor UO_1010 (O_1010,N_24753,N_24995);
and UO_1011 (O_1011,N_24790,N_24583);
or UO_1012 (O_1012,N_24976,N_24554);
and UO_1013 (O_1013,N_24899,N_24785);
nor UO_1014 (O_1014,N_24967,N_24638);
nor UO_1015 (O_1015,N_24714,N_24554);
nor UO_1016 (O_1016,N_24905,N_24635);
nand UO_1017 (O_1017,N_24789,N_24842);
nor UO_1018 (O_1018,N_24604,N_24605);
and UO_1019 (O_1019,N_24522,N_24739);
xnor UO_1020 (O_1020,N_24583,N_24535);
or UO_1021 (O_1021,N_24904,N_24896);
nor UO_1022 (O_1022,N_24681,N_24650);
and UO_1023 (O_1023,N_24617,N_24736);
nor UO_1024 (O_1024,N_24943,N_24956);
nand UO_1025 (O_1025,N_24651,N_24745);
and UO_1026 (O_1026,N_24908,N_24600);
nand UO_1027 (O_1027,N_24553,N_24861);
nor UO_1028 (O_1028,N_24955,N_24807);
nor UO_1029 (O_1029,N_24747,N_24901);
nand UO_1030 (O_1030,N_24505,N_24707);
nand UO_1031 (O_1031,N_24882,N_24769);
nor UO_1032 (O_1032,N_24951,N_24686);
and UO_1033 (O_1033,N_24928,N_24794);
nor UO_1034 (O_1034,N_24737,N_24920);
nor UO_1035 (O_1035,N_24790,N_24851);
and UO_1036 (O_1036,N_24784,N_24614);
and UO_1037 (O_1037,N_24590,N_24912);
xnor UO_1038 (O_1038,N_24930,N_24924);
or UO_1039 (O_1039,N_24549,N_24886);
or UO_1040 (O_1040,N_24753,N_24989);
and UO_1041 (O_1041,N_24518,N_24830);
xor UO_1042 (O_1042,N_24920,N_24704);
xnor UO_1043 (O_1043,N_24955,N_24887);
xor UO_1044 (O_1044,N_24586,N_24720);
xnor UO_1045 (O_1045,N_24612,N_24684);
nand UO_1046 (O_1046,N_24796,N_24503);
and UO_1047 (O_1047,N_24802,N_24689);
or UO_1048 (O_1048,N_24583,N_24670);
nor UO_1049 (O_1049,N_24556,N_24527);
nand UO_1050 (O_1050,N_24716,N_24624);
and UO_1051 (O_1051,N_24586,N_24853);
and UO_1052 (O_1052,N_24611,N_24658);
and UO_1053 (O_1053,N_24554,N_24796);
or UO_1054 (O_1054,N_24520,N_24514);
and UO_1055 (O_1055,N_24654,N_24987);
nand UO_1056 (O_1056,N_24664,N_24822);
and UO_1057 (O_1057,N_24538,N_24649);
and UO_1058 (O_1058,N_24876,N_24732);
nand UO_1059 (O_1059,N_24738,N_24949);
or UO_1060 (O_1060,N_24963,N_24724);
xor UO_1061 (O_1061,N_24664,N_24561);
and UO_1062 (O_1062,N_24905,N_24713);
nand UO_1063 (O_1063,N_24582,N_24676);
and UO_1064 (O_1064,N_24698,N_24559);
nand UO_1065 (O_1065,N_24792,N_24886);
nand UO_1066 (O_1066,N_24585,N_24683);
nand UO_1067 (O_1067,N_24981,N_24794);
xnor UO_1068 (O_1068,N_24885,N_24580);
xor UO_1069 (O_1069,N_24874,N_24621);
xnor UO_1070 (O_1070,N_24937,N_24886);
xnor UO_1071 (O_1071,N_24977,N_24539);
xor UO_1072 (O_1072,N_24911,N_24561);
nand UO_1073 (O_1073,N_24642,N_24639);
nor UO_1074 (O_1074,N_24667,N_24715);
or UO_1075 (O_1075,N_24566,N_24906);
nand UO_1076 (O_1076,N_24866,N_24959);
xnor UO_1077 (O_1077,N_24659,N_24782);
xor UO_1078 (O_1078,N_24641,N_24534);
or UO_1079 (O_1079,N_24575,N_24888);
nor UO_1080 (O_1080,N_24667,N_24846);
and UO_1081 (O_1081,N_24916,N_24781);
nand UO_1082 (O_1082,N_24967,N_24839);
nand UO_1083 (O_1083,N_24750,N_24508);
nor UO_1084 (O_1084,N_24867,N_24692);
nor UO_1085 (O_1085,N_24958,N_24568);
xor UO_1086 (O_1086,N_24892,N_24734);
or UO_1087 (O_1087,N_24984,N_24662);
nor UO_1088 (O_1088,N_24810,N_24685);
or UO_1089 (O_1089,N_24755,N_24833);
nand UO_1090 (O_1090,N_24547,N_24586);
or UO_1091 (O_1091,N_24753,N_24563);
xor UO_1092 (O_1092,N_24906,N_24809);
and UO_1093 (O_1093,N_24949,N_24733);
xnor UO_1094 (O_1094,N_24825,N_24745);
nor UO_1095 (O_1095,N_24905,N_24693);
and UO_1096 (O_1096,N_24725,N_24878);
and UO_1097 (O_1097,N_24557,N_24936);
xor UO_1098 (O_1098,N_24637,N_24744);
and UO_1099 (O_1099,N_24798,N_24568);
nor UO_1100 (O_1100,N_24635,N_24862);
xnor UO_1101 (O_1101,N_24992,N_24891);
nor UO_1102 (O_1102,N_24878,N_24561);
xnor UO_1103 (O_1103,N_24913,N_24622);
xnor UO_1104 (O_1104,N_24935,N_24614);
nor UO_1105 (O_1105,N_24648,N_24656);
nor UO_1106 (O_1106,N_24767,N_24531);
xor UO_1107 (O_1107,N_24757,N_24511);
or UO_1108 (O_1108,N_24740,N_24960);
xor UO_1109 (O_1109,N_24726,N_24979);
nor UO_1110 (O_1110,N_24645,N_24652);
or UO_1111 (O_1111,N_24994,N_24990);
and UO_1112 (O_1112,N_24928,N_24552);
xnor UO_1113 (O_1113,N_24608,N_24534);
nor UO_1114 (O_1114,N_24998,N_24624);
xor UO_1115 (O_1115,N_24754,N_24652);
nor UO_1116 (O_1116,N_24741,N_24643);
and UO_1117 (O_1117,N_24841,N_24532);
nor UO_1118 (O_1118,N_24875,N_24567);
xnor UO_1119 (O_1119,N_24931,N_24531);
nor UO_1120 (O_1120,N_24593,N_24624);
nand UO_1121 (O_1121,N_24965,N_24571);
and UO_1122 (O_1122,N_24769,N_24711);
nand UO_1123 (O_1123,N_24817,N_24757);
and UO_1124 (O_1124,N_24933,N_24824);
or UO_1125 (O_1125,N_24985,N_24858);
nor UO_1126 (O_1126,N_24908,N_24810);
or UO_1127 (O_1127,N_24534,N_24566);
or UO_1128 (O_1128,N_24580,N_24945);
or UO_1129 (O_1129,N_24683,N_24886);
nand UO_1130 (O_1130,N_24518,N_24606);
nand UO_1131 (O_1131,N_24594,N_24508);
and UO_1132 (O_1132,N_24525,N_24957);
xor UO_1133 (O_1133,N_24501,N_24810);
xor UO_1134 (O_1134,N_24841,N_24613);
nor UO_1135 (O_1135,N_24862,N_24693);
xnor UO_1136 (O_1136,N_24670,N_24795);
xor UO_1137 (O_1137,N_24725,N_24576);
xor UO_1138 (O_1138,N_24918,N_24587);
xor UO_1139 (O_1139,N_24787,N_24614);
nor UO_1140 (O_1140,N_24704,N_24625);
and UO_1141 (O_1141,N_24525,N_24528);
nand UO_1142 (O_1142,N_24635,N_24947);
nor UO_1143 (O_1143,N_24937,N_24858);
or UO_1144 (O_1144,N_24889,N_24657);
and UO_1145 (O_1145,N_24774,N_24503);
or UO_1146 (O_1146,N_24949,N_24744);
or UO_1147 (O_1147,N_24526,N_24771);
and UO_1148 (O_1148,N_24716,N_24577);
xnor UO_1149 (O_1149,N_24880,N_24641);
nor UO_1150 (O_1150,N_24544,N_24724);
nor UO_1151 (O_1151,N_24602,N_24920);
and UO_1152 (O_1152,N_24667,N_24764);
xnor UO_1153 (O_1153,N_24631,N_24799);
or UO_1154 (O_1154,N_24972,N_24738);
nand UO_1155 (O_1155,N_24779,N_24925);
xnor UO_1156 (O_1156,N_24871,N_24517);
xor UO_1157 (O_1157,N_24505,N_24809);
nor UO_1158 (O_1158,N_24890,N_24635);
nor UO_1159 (O_1159,N_24566,N_24554);
nor UO_1160 (O_1160,N_24765,N_24984);
or UO_1161 (O_1161,N_24987,N_24975);
nor UO_1162 (O_1162,N_24596,N_24975);
nand UO_1163 (O_1163,N_24563,N_24910);
nor UO_1164 (O_1164,N_24718,N_24655);
or UO_1165 (O_1165,N_24627,N_24975);
and UO_1166 (O_1166,N_24941,N_24580);
and UO_1167 (O_1167,N_24854,N_24630);
nor UO_1168 (O_1168,N_24703,N_24955);
xnor UO_1169 (O_1169,N_24786,N_24623);
and UO_1170 (O_1170,N_24651,N_24812);
and UO_1171 (O_1171,N_24677,N_24973);
nand UO_1172 (O_1172,N_24715,N_24863);
nor UO_1173 (O_1173,N_24654,N_24757);
xnor UO_1174 (O_1174,N_24960,N_24939);
and UO_1175 (O_1175,N_24628,N_24864);
or UO_1176 (O_1176,N_24936,N_24957);
xnor UO_1177 (O_1177,N_24939,N_24807);
nand UO_1178 (O_1178,N_24864,N_24920);
nand UO_1179 (O_1179,N_24837,N_24791);
nand UO_1180 (O_1180,N_24735,N_24789);
nor UO_1181 (O_1181,N_24556,N_24761);
and UO_1182 (O_1182,N_24768,N_24786);
nor UO_1183 (O_1183,N_24830,N_24814);
or UO_1184 (O_1184,N_24887,N_24706);
nor UO_1185 (O_1185,N_24935,N_24511);
and UO_1186 (O_1186,N_24750,N_24905);
nor UO_1187 (O_1187,N_24620,N_24878);
xor UO_1188 (O_1188,N_24547,N_24999);
or UO_1189 (O_1189,N_24591,N_24989);
xor UO_1190 (O_1190,N_24512,N_24939);
xor UO_1191 (O_1191,N_24852,N_24723);
nor UO_1192 (O_1192,N_24861,N_24990);
and UO_1193 (O_1193,N_24838,N_24578);
nor UO_1194 (O_1194,N_24969,N_24759);
xnor UO_1195 (O_1195,N_24851,N_24850);
nand UO_1196 (O_1196,N_24591,N_24825);
xnor UO_1197 (O_1197,N_24616,N_24685);
and UO_1198 (O_1198,N_24550,N_24766);
nand UO_1199 (O_1199,N_24503,N_24524);
or UO_1200 (O_1200,N_24710,N_24901);
and UO_1201 (O_1201,N_24594,N_24800);
and UO_1202 (O_1202,N_24641,N_24967);
xor UO_1203 (O_1203,N_24746,N_24901);
nand UO_1204 (O_1204,N_24680,N_24619);
and UO_1205 (O_1205,N_24546,N_24859);
nand UO_1206 (O_1206,N_24827,N_24584);
xnor UO_1207 (O_1207,N_24908,N_24739);
and UO_1208 (O_1208,N_24561,N_24699);
nand UO_1209 (O_1209,N_24518,N_24578);
or UO_1210 (O_1210,N_24793,N_24604);
or UO_1211 (O_1211,N_24663,N_24832);
and UO_1212 (O_1212,N_24595,N_24820);
or UO_1213 (O_1213,N_24850,N_24809);
xor UO_1214 (O_1214,N_24594,N_24942);
nand UO_1215 (O_1215,N_24658,N_24780);
and UO_1216 (O_1216,N_24586,N_24797);
nand UO_1217 (O_1217,N_24758,N_24759);
or UO_1218 (O_1218,N_24716,N_24705);
or UO_1219 (O_1219,N_24922,N_24919);
nand UO_1220 (O_1220,N_24749,N_24951);
xor UO_1221 (O_1221,N_24999,N_24792);
and UO_1222 (O_1222,N_24612,N_24943);
and UO_1223 (O_1223,N_24985,N_24665);
nor UO_1224 (O_1224,N_24854,N_24682);
nand UO_1225 (O_1225,N_24525,N_24982);
or UO_1226 (O_1226,N_24552,N_24922);
and UO_1227 (O_1227,N_24662,N_24736);
xnor UO_1228 (O_1228,N_24916,N_24696);
xnor UO_1229 (O_1229,N_24966,N_24712);
and UO_1230 (O_1230,N_24818,N_24765);
or UO_1231 (O_1231,N_24886,N_24503);
xor UO_1232 (O_1232,N_24694,N_24723);
xor UO_1233 (O_1233,N_24741,N_24840);
nand UO_1234 (O_1234,N_24526,N_24848);
nor UO_1235 (O_1235,N_24525,N_24947);
and UO_1236 (O_1236,N_24897,N_24751);
nand UO_1237 (O_1237,N_24778,N_24641);
xor UO_1238 (O_1238,N_24831,N_24596);
xnor UO_1239 (O_1239,N_24974,N_24725);
or UO_1240 (O_1240,N_24647,N_24535);
or UO_1241 (O_1241,N_24814,N_24924);
nand UO_1242 (O_1242,N_24875,N_24908);
nand UO_1243 (O_1243,N_24753,N_24648);
and UO_1244 (O_1244,N_24987,N_24673);
xor UO_1245 (O_1245,N_24563,N_24833);
nand UO_1246 (O_1246,N_24936,N_24694);
and UO_1247 (O_1247,N_24583,N_24887);
or UO_1248 (O_1248,N_24838,N_24853);
and UO_1249 (O_1249,N_24557,N_24679);
nand UO_1250 (O_1250,N_24971,N_24548);
or UO_1251 (O_1251,N_24708,N_24821);
nor UO_1252 (O_1252,N_24909,N_24884);
xor UO_1253 (O_1253,N_24567,N_24744);
xnor UO_1254 (O_1254,N_24886,N_24947);
and UO_1255 (O_1255,N_24869,N_24549);
and UO_1256 (O_1256,N_24935,N_24556);
xor UO_1257 (O_1257,N_24988,N_24619);
nand UO_1258 (O_1258,N_24954,N_24509);
nand UO_1259 (O_1259,N_24554,N_24794);
or UO_1260 (O_1260,N_24911,N_24795);
and UO_1261 (O_1261,N_24575,N_24522);
or UO_1262 (O_1262,N_24979,N_24526);
nor UO_1263 (O_1263,N_24582,N_24600);
or UO_1264 (O_1264,N_24855,N_24830);
nor UO_1265 (O_1265,N_24898,N_24741);
or UO_1266 (O_1266,N_24915,N_24922);
nand UO_1267 (O_1267,N_24790,N_24818);
and UO_1268 (O_1268,N_24951,N_24617);
nand UO_1269 (O_1269,N_24906,N_24626);
nand UO_1270 (O_1270,N_24727,N_24751);
and UO_1271 (O_1271,N_24993,N_24540);
and UO_1272 (O_1272,N_24554,N_24912);
nor UO_1273 (O_1273,N_24727,N_24838);
and UO_1274 (O_1274,N_24752,N_24531);
and UO_1275 (O_1275,N_24721,N_24892);
and UO_1276 (O_1276,N_24629,N_24516);
and UO_1277 (O_1277,N_24649,N_24563);
nor UO_1278 (O_1278,N_24745,N_24970);
nand UO_1279 (O_1279,N_24605,N_24580);
xor UO_1280 (O_1280,N_24951,N_24857);
xnor UO_1281 (O_1281,N_24902,N_24770);
and UO_1282 (O_1282,N_24831,N_24796);
or UO_1283 (O_1283,N_24893,N_24824);
nor UO_1284 (O_1284,N_24558,N_24972);
xor UO_1285 (O_1285,N_24916,N_24627);
or UO_1286 (O_1286,N_24847,N_24963);
xor UO_1287 (O_1287,N_24865,N_24864);
nand UO_1288 (O_1288,N_24617,N_24536);
xor UO_1289 (O_1289,N_24671,N_24725);
xor UO_1290 (O_1290,N_24925,N_24610);
and UO_1291 (O_1291,N_24508,N_24575);
nand UO_1292 (O_1292,N_24899,N_24815);
xor UO_1293 (O_1293,N_24681,N_24747);
xnor UO_1294 (O_1294,N_24676,N_24537);
xor UO_1295 (O_1295,N_24502,N_24960);
xor UO_1296 (O_1296,N_24549,N_24870);
nor UO_1297 (O_1297,N_24792,N_24634);
xnor UO_1298 (O_1298,N_24923,N_24910);
and UO_1299 (O_1299,N_24675,N_24626);
and UO_1300 (O_1300,N_24636,N_24727);
nor UO_1301 (O_1301,N_24950,N_24855);
xor UO_1302 (O_1302,N_24777,N_24751);
or UO_1303 (O_1303,N_24779,N_24813);
xor UO_1304 (O_1304,N_24763,N_24801);
nor UO_1305 (O_1305,N_24696,N_24947);
or UO_1306 (O_1306,N_24869,N_24888);
nor UO_1307 (O_1307,N_24850,N_24569);
or UO_1308 (O_1308,N_24824,N_24731);
and UO_1309 (O_1309,N_24579,N_24946);
and UO_1310 (O_1310,N_24548,N_24569);
and UO_1311 (O_1311,N_24912,N_24532);
nor UO_1312 (O_1312,N_24654,N_24967);
or UO_1313 (O_1313,N_24514,N_24690);
xnor UO_1314 (O_1314,N_24895,N_24993);
or UO_1315 (O_1315,N_24754,N_24808);
and UO_1316 (O_1316,N_24533,N_24928);
xor UO_1317 (O_1317,N_24658,N_24734);
nor UO_1318 (O_1318,N_24983,N_24602);
and UO_1319 (O_1319,N_24936,N_24993);
nor UO_1320 (O_1320,N_24954,N_24580);
and UO_1321 (O_1321,N_24754,N_24793);
xor UO_1322 (O_1322,N_24800,N_24788);
nand UO_1323 (O_1323,N_24707,N_24533);
nand UO_1324 (O_1324,N_24570,N_24601);
and UO_1325 (O_1325,N_24535,N_24705);
xor UO_1326 (O_1326,N_24645,N_24930);
and UO_1327 (O_1327,N_24748,N_24961);
nor UO_1328 (O_1328,N_24988,N_24990);
and UO_1329 (O_1329,N_24994,N_24825);
nand UO_1330 (O_1330,N_24570,N_24579);
nor UO_1331 (O_1331,N_24560,N_24669);
nand UO_1332 (O_1332,N_24943,N_24726);
nand UO_1333 (O_1333,N_24807,N_24719);
nand UO_1334 (O_1334,N_24694,N_24659);
nand UO_1335 (O_1335,N_24710,N_24608);
and UO_1336 (O_1336,N_24508,N_24821);
nor UO_1337 (O_1337,N_24583,N_24841);
xor UO_1338 (O_1338,N_24911,N_24516);
and UO_1339 (O_1339,N_24590,N_24515);
or UO_1340 (O_1340,N_24952,N_24845);
nand UO_1341 (O_1341,N_24533,N_24619);
and UO_1342 (O_1342,N_24935,N_24621);
nor UO_1343 (O_1343,N_24804,N_24570);
nor UO_1344 (O_1344,N_24904,N_24987);
nand UO_1345 (O_1345,N_24518,N_24512);
xnor UO_1346 (O_1346,N_24665,N_24765);
and UO_1347 (O_1347,N_24680,N_24625);
nand UO_1348 (O_1348,N_24874,N_24501);
or UO_1349 (O_1349,N_24793,N_24648);
nor UO_1350 (O_1350,N_24990,N_24579);
and UO_1351 (O_1351,N_24645,N_24553);
xor UO_1352 (O_1352,N_24550,N_24869);
nand UO_1353 (O_1353,N_24710,N_24724);
nand UO_1354 (O_1354,N_24608,N_24962);
nor UO_1355 (O_1355,N_24889,N_24685);
or UO_1356 (O_1356,N_24763,N_24614);
nor UO_1357 (O_1357,N_24667,N_24701);
nor UO_1358 (O_1358,N_24524,N_24735);
nand UO_1359 (O_1359,N_24578,N_24762);
nand UO_1360 (O_1360,N_24517,N_24622);
or UO_1361 (O_1361,N_24969,N_24642);
nor UO_1362 (O_1362,N_24648,N_24710);
and UO_1363 (O_1363,N_24579,N_24714);
or UO_1364 (O_1364,N_24817,N_24769);
xor UO_1365 (O_1365,N_24847,N_24555);
and UO_1366 (O_1366,N_24623,N_24981);
nor UO_1367 (O_1367,N_24614,N_24910);
and UO_1368 (O_1368,N_24600,N_24765);
nor UO_1369 (O_1369,N_24656,N_24590);
nor UO_1370 (O_1370,N_24591,N_24514);
and UO_1371 (O_1371,N_24924,N_24576);
xnor UO_1372 (O_1372,N_24863,N_24856);
and UO_1373 (O_1373,N_24881,N_24817);
or UO_1374 (O_1374,N_24696,N_24873);
or UO_1375 (O_1375,N_24801,N_24656);
nand UO_1376 (O_1376,N_24857,N_24535);
xor UO_1377 (O_1377,N_24645,N_24862);
xnor UO_1378 (O_1378,N_24782,N_24984);
xor UO_1379 (O_1379,N_24929,N_24551);
xor UO_1380 (O_1380,N_24866,N_24892);
nand UO_1381 (O_1381,N_24500,N_24809);
nand UO_1382 (O_1382,N_24676,N_24818);
nor UO_1383 (O_1383,N_24613,N_24581);
and UO_1384 (O_1384,N_24628,N_24625);
and UO_1385 (O_1385,N_24833,N_24522);
xor UO_1386 (O_1386,N_24844,N_24508);
and UO_1387 (O_1387,N_24551,N_24777);
nor UO_1388 (O_1388,N_24621,N_24513);
or UO_1389 (O_1389,N_24987,N_24888);
or UO_1390 (O_1390,N_24949,N_24848);
and UO_1391 (O_1391,N_24605,N_24927);
nand UO_1392 (O_1392,N_24983,N_24662);
or UO_1393 (O_1393,N_24986,N_24813);
nand UO_1394 (O_1394,N_24889,N_24630);
xnor UO_1395 (O_1395,N_24974,N_24510);
nor UO_1396 (O_1396,N_24564,N_24663);
nor UO_1397 (O_1397,N_24781,N_24636);
nor UO_1398 (O_1398,N_24560,N_24924);
xor UO_1399 (O_1399,N_24817,N_24637);
nor UO_1400 (O_1400,N_24778,N_24792);
xor UO_1401 (O_1401,N_24875,N_24526);
or UO_1402 (O_1402,N_24816,N_24657);
nand UO_1403 (O_1403,N_24776,N_24962);
nor UO_1404 (O_1404,N_24700,N_24711);
xor UO_1405 (O_1405,N_24630,N_24699);
nand UO_1406 (O_1406,N_24730,N_24645);
nand UO_1407 (O_1407,N_24762,N_24873);
xnor UO_1408 (O_1408,N_24796,N_24764);
or UO_1409 (O_1409,N_24539,N_24603);
nor UO_1410 (O_1410,N_24680,N_24660);
or UO_1411 (O_1411,N_24506,N_24964);
nand UO_1412 (O_1412,N_24521,N_24664);
nor UO_1413 (O_1413,N_24826,N_24944);
nand UO_1414 (O_1414,N_24796,N_24904);
nor UO_1415 (O_1415,N_24812,N_24503);
xnor UO_1416 (O_1416,N_24944,N_24729);
xor UO_1417 (O_1417,N_24795,N_24527);
xor UO_1418 (O_1418,N_24525,N_24745);
and UO_1419 (O_1419,N_24542,N_24821);
and UO_1420 (O_1420,N_24678,N_24637);
nand UO_1421 (O_1421,N_24899,N_24554);
or UO_1422 (O_1422,N_24615,N_24928);
nor UO_1423 (O_1423,N_24555,N_24839);
nor UO_1424 (O_1424,N_24561,N_24661);
xnor UO_1425 (O_1425,N_24910,N_24675);
nand UO_1426 (O_1426,N_24793,N_24520);
or UO_1427 (O_1427,N_24751,N_24835);
nor UO_1428 (O_1428,N_24629,N_24752);
and UO_1429 (O_1429,N_24515,N_24893);
nand UO_1430 (O_1430,N_24574,N_24825);
nor UO_1431 (O_1431,N_24629,N_24505);
nand UO_1432 (O_1432,N_24940,N_24773);
or UO_1433 (O_1433,N_24566,N_24720);
xnor UO_1434 (O_1434,N_24911,N_24676);
and UO_1435 (O_1435,N_24663,N_24669);
nor UO_1436 (O_1436,N_24956,N_24578);
or UO_1437 (O_1437,N_24854,N_24504);
nor UO_1438 (O_1438,N_24967,N_24679);
and UO_1439 (O_1439,N_24733,N_24913);
and UO_1440 (O_1440,N_24987,N_24750);
and UO_1441 (O_1441,N_24643,N_24628);
or UO_1442 (O_1442,N_24834,N_24576);
and UO_1443 (O_1443,N_24751,N_24515);
and UO_1444 (O_1444,N_24925,N_24987);
nor UO_1445 (O_1445,N_24693,N_24561);
and UO_1446 (O_1446,N_24662,N_24629);
or UO_1447 (O_1447,N_24922,N_24599);
xnor UO_1448 (O_1448,N_24770,N_24678);
and UO_1449 (O_1449,N_24556,N_24791);
nand UO_1450 (O_1450,N_24895,N_24680);
and UO_1451 (O_1451,N_24990,N_24824);
nand UO_1452 (O_1452,N_24607,N_24732);
and UO_1453 (O_1453,N_24996,N_24579);
or UO_1454 (O_1454,N_24872,N_24685);
and UO_1455 (O_1455,N_24695,N_24871);
or UO_1456 (O_1456,N_24538,N_24589);
and UO_1457 (O_1457,N_24512,N_24991);
nand UO_1458 (O_1458,N_24662,N_24691);
and UO_1459 (O_1459,N_24997,N_24906);
and UO_1460 (O_1460,N_24724,N_24930);
and UO_1461 (O_1461,N_24758,N_24574);
nor UO_1462 (O_1462,N_24884,N_24851);
nor UO_1463 (O_1463,N_24887,N_24597);
or UO_1464 (O_1464,N_24597,N_24554);
nand UO_1465 (O_1465,N_24632,N_24950);
and UO_1466 (O_1466,N_24991,N_24829);
nand UO_1467 (O_1467,N_24672,N_24500);
nor UO_1468 (O_1468,N_24663,N_24664);
and UO_1469 (O_1469,N_24924,N_24573);
nand UO_1470 (O_1470,N_24637,N_24845);
nand UO_1471 (O_1471,N_24826,N_24535);
xor UO_1472 (O_1472,N_24724,N_24977);
or UO_1473 (O_1473,N_24569,N_24701);
or UO_1474 (O_1474,N_24863,N_24928);
xor UO_1475 (O_1475,N_24752,N_24643);
nand UO_1476 (O_1476,N_24689,N_24974);
or UO_1477 (O_1477,N_24644,N_24949);
or UO_1478 (O_1478,N_24512,N_24705);
xnor UO_1479 (O_1479,N_24652,N_24819);
and UO_1480 (O_1480,N_24655,N_24667);
nor UO_1481 (O_1481,N_24843,N_24670);
and UO_1482 (O_1482,N_24980,N_24531);
or UO_1483 (O_1483,N_24690,N_24995);
and UO_1484 (O_1484,N_24620,N_24786);
xor UO_1485 (O_1485,N_24633,N_24667);
or UO_1486 (O_1486,N_24668,N_24547);
or UO_1487 (O_1487,N_24945,N_24807);
or UO_1488 (O_1488,N_24753,N_24641);
nand UO_1489 (O_1489,N_24719,N_24936);
or UO_1490 (O_1490,N_24626,N_24595);
and UO_1491 (O_1491,N_24763,N_24537);
and UO_1492 (O_1492,N_24621,N_24500);
nor UO_1493 (O_1493,N_24840,N_24531);
or UO_1494 (O_1494,N_24705,N_24850);
nand UO_1495 (O_1495,N_24860,N_24889);
and UO_1496 (O_1496,N_24770,N_24946);
nand UO_1497 (O_1497,N_24886,N_24801);
nor UO_1498 (O_1498,N_24553,N_24667);
xor UO_1499 (O_1499,N_24758,N_24576);
nand UO_1500 (O_1500,N_24577,N_24694);
nand UO_1501 (O_1501,N_24595,N_24892);
and UO_1502 (O_1502,N_24886,N_24849);
or UO_1503 (O_1503,N_24584,N_24818);
nor UO_1504 (O_1504,N_24917,N_24732);
nor UO_1505 (O_1505,N_24634,N_24662);
and UO_1506 (O_1506,N_24942,N_24754);
and UO_1507 (O_1507,N_24991,N_24806);
or UO_1508 (O_1508,N_24641,N_24767);
nand UO_1509 (O_1509,N_24961,N_24602);
or UO_1510 (O_1510,N_24875,N_24999);
or UO_1511 (O_1511,N_24936,N_24623);
xnor UO_1512 (O_1512,N_24817,N_24945);
nor UO_1513 (O_1513,N_24625,N_24983);
nand UO_1514 (O_1514,N_24786,N_24515);
nor UO_1515 (O_1515,N_24814,N_24973);
nor UO_1516 (O_1516,N_24885,N_24819);
nand UO_1517 (O_1517,N_24775,N_24938);
xnor UO_1518 (O_1518,N_24542,N_24732);
or UO_1519 (O_1519,N_24521,N_24755);
and UO_1520 (O_1520,N_24944,N_24726);
or UO_1521 (O_1521,N_24532,N_24838);
nand UO_1522 (O_1522,N_24514,N_24984);
nand UO_1523 (O_1523,N_24863,N_24957);
xor UO_1524 (O_1524,N_24631,N_24606);
or UO_1525 (O_1525,N_24967,N_24881);
nand UO_1526 (O_1526,N_24859,N_24816);
or UO_1527 (O_1527,N_24601,N_24775);
or UO_1528 (O_1528,N_24514,N_24601);
xnor UO_1529 (O_1529,N_24594,N_24815);
and UO_1530 (O_1530,N_24715,N_24525);
nor UO_1531 (O_1531,N_24858,N_24561);
and UO_1532 (O_1532,N_24783,N_24744);
nor UO_1533 (O_1533,N_24531,N_24832);
nand UO_1534 (O_1534,N_24738,N_24929);
xnor UO_1535 (O_1535,N_24645,N_24664);
or UO_1536 (O_1536,N_24565,N_24847);
nand UO_1537 (O_1537,N_24982,N_24962);
or UO_1538 (O_1538,N_24670,N_24807);
nand UO_1539 (O_1539,N_24703,N_24706);
or UO_1540 (O_1540,N_24925,N_24652);
or UO_1541 (O_1541,N_24950,N_24677);
nor UO_1542 (O_1542,N_24670,N_24683);
xor UO_1543 (O_1543,N_24817,N_24840);
xnor UO_1544 (O_1544,N_24526,N_24969);
nand UO_1545 (O_1545,N_24767,N_24770);
or UO_1546 (O_1546,N_24611,N_24566);
xnor UO_1547 (O_1547,N_24879,N_24755);
nand UO_1548 (O_1548,N_24705,N_24516);
nor UO_1549 (O_1549,N_24549,N_24853);
and UO_1550 (O_1550,N_24598,N_24982);
nor UO_1551 (O_1551,N_24556,N_24832);
nand UO_1552 (O_1552,N_24585,N_24870);
nor UO_1553 (O_1553,N_24743,N_24620);
nor UO_1554 (O_1554,N_24832,N_24636);
and UO_1555 (O_1555,N_24762,N_24604);
and UO_1556 (O_1556,N_24944,N_24774);
nand UO_1557 (O_1557,N_24859,N_24978);
or UO_1558 (O_1558,N_24644,N_24955);
nand UO_1559 (O_1559,N_24648,N_24655);
and UO_1560 (O_1560,N_24538,N_24844);
or UO_1561 (O_1561,N_24718,N_24601);
nor UO_1562 (O_1562,N_24515,N_24594);
xor UO_1563 (O_1563,N_24852,N_24702);
or UO_1564 (O_1564,N_24801,N_24704);
xor UO_1565 (O_1565,N_24755,N_24835);
nand UO_1566 (O_1566,N_24689,N_24798);
nand UO_1567 (O_1567,N_24948,N_24508);
xor UO_1568 (O_1568,N_24536,N_24532);
xnor UO_1569 (O_1569,N_24965,N_24599);
xnor UO_1570 (O_1570,N_24944,N_24827);
xnor UO_1571 (O_1571,N_24873,N_24708);
xor UO_1572 (O_1572,N_24784,N_24791);
or UO_1573 (O_1573,N_24796,N_24700);
nor UO_1574 (O_1574,N_24829,N_24616);
nor UO_1575 (O_1575,N_24659,N_24584);
nand UO_1576 (O_1576,N_24844,N_24854);
nand UO_1577 (O_1577,N_24797,N_24704);
nor UO_1578 (O_1578,N_24733,N_24868);
xnor UO_1579 (O_1579,N_24852,N_24856);
xor UO_1580 (O_1580,N_24681,N_24751);
and UO_1581 (O_1581,N_24916,N_24702);
xor UO_1582 (O_1582,N_24715,N_24778);
and UO_1583 (O_1583,N_24644,N_24914);
nor UO_1584 (O_1584,N_24838,N_24519);
xor UO_1585 (O_1585,N_24856,N_24995);
nor UO_1586 (O_1586,N_24933,N_24750);
nor UO_1587 (O_1587,N_24795,N_24636);
or UO_1588 (O_1588,N_24947,N_24855);
xnor UO_1589 (O_1589,N_24841,N_24764);
xor UO_1590 (O_1590,N_24971,N_24697);
nand UO_1591 (O_1591,N_24642,N_24857);
or UO_1592 (O_1592,N_24875,N_24809);
or UO_1593 (O_1593,N_24580,N_24767);
xor UO_1594 (O_1594,N_24875,N_24927);
or UO_1595 (O_1595,N_24629,N_24514);
nor UO_1596 (O_1596,N_24564,N_24560);
nor UO_1597 (O_1597,N_24711,N_24578);
nor UO_1598 (O_1598,N_24577,N_24735);
nand UO_1599 (O_1599,N_24759,N_24819);
or UO_1600 (O_1600,N_24932,N_24680);
nand UO_1601 (O_1601,N_24836,N_24580);
xnor UO_1602 (O_1602,N_24567,N_24598);
xnor UO_1603 (O_1603,N_24856,N_24685);
nor UO_1604 (O_1604,N_24843,N_24980);
nand UO_1605 (O_1605,N_24751,N_24838);
nor UO_1606 (O_1606,N_24773,N_24628);
nand UO_1607 (O_1607,N_24867,N_24533);
xnor UO_1608 (O_1608,N_24885,N_24562);
or UO_1609 (O_1609,N_24966,N_24804);
xor UO_1610 (O_1610,N_24945,N_24556);
nand UO_1611 (O_1611,N_24545,N_24569);
or UO_1612 (O_1612,N_24716,N_24870);
or UO_1613 (O_1613,N_24824,N_24525);
nor UO_1614 (O_1614,N_24959,N_24518);
nor UO_1615 (O_1615,N_24652,N_24641);
nor UO_1616 (O_1616,N_24700,N_24697);
and UO_1617 (O_1617,N_24799,N_24795);
and UO_1618 (O_1618,N_24946,N_24705);
and UO_1619 (O_1619,N_24865,N_24978);
xnor UO_1620 (O_1620,N_24931,N_24880);
or UO_1621 (O_1621,N_24747,N_24573);
xnor UO_1622 (O_1622,N_24634,N_24523);
or UO_1623 (O_1623,N_24873,N_24672);
nor UO_1624 (O_1624,N_24850,N_24610);
or UO_1625 (O_1625,N_24565,N_24849);
xor UO_1626 (O_1626,N_24971,N_24806);
nand UO_1627 (O_1627,N_24829,N_24972);
nor UO_1628 (O_1628,N_24748,N_24530);
nand UO_1629 (O_1629,N_24849,N_24629);
nor UO_1630 (O_1630,N_24717,N_24904);
nand UO_1631 (O_1631,N_24773,N_24850);
or UO_1632 (O_1632,N_24897,N_24918);
and UO_1633 (O_1633,N_24663,N_24747);
and UO_1634 (O_1634,N_24835,N_24912);
nand UO_1635 (O_1635,N_24624,N_24531);
or UO_1636 (O_1636,N_24584,N_24970);
or UO_1637 (O_1637,N_24522,N_24639);
nand UO_1638 (O_1638,N_24598,N_24978);
nand UO_1639 (O_1639,N_24892,N_24698);
xnor UO_1640 (O_1640,N_24823,N_24861);
nor UO_1641 (O_1641,N_24549,N_24545);
and UO_1642 (O_1642,N_24595,N_24633);
and UO_1643 (O_1643,N_24785,N_24711);
and UO_1644 (O_1644,N_24776,N_24953);
nor UO_1645 (O_1645,N_24927,N_24543);
nand UO_1646 (O_1646,N_24561,N_24621);
nor UO_1647 (O_1647,N_24952,N_24534);
or UO_1648 (O_1648,N_24586,N_24696);
nor UO_1649 (O_1649,N_24818,N_24557);
and UO_1650 (O_1650,N_24978,N_24602);
and UO_1651 (O_1651,N_24533,N_24765);
nor UO_1652 (O_1652,N_24764,N_24692);
xnor UO_1653 (O_1653,N_24814,N_24623);
nor UO_1654 (O_1654,N_24569,N_24907);
nand UO_1655 (O_1655,N_24961,N_24758);
nand UO_1656 (O_1656,N_24723,N_24990);
and UO_1657 (O_1657,N_24653,N_24614);
or UO_1658 (O_1658,N_24999,N_24694);
xnor UO_1659 (O_1659,N_24969,N_24505);
and UO_1660 (O_1660,N_24813,N_24553);
xnor UO_1661 (O_1661,N_24634,N_24883);
nand UO_1662 (O_1662,N_24983,N_24984);
or UO_1663 (O_1663,N_24784,N_24580);
or UO_1664 (O_1664,N_24600,N_24875);
nor UO_1665 (O_1665,N_24789,N_24919);
nand UO_1666 (O_1666,N_24560,N_24622);
xor UO_1667 (O_1667,N_24744,N_24852);
or UO_1668 (O_1668,N_24889,N_24571);
xnor UO_1669 (O_1669,N_24746,N_24555);
xor UO_1670 (O_1670,N_24726,N_24524);
xor UO_1671 (O_1671,N_24604,N_24985);
xor UO_1672 (O_1672,N_24693,N_24714);
nand UO_1673 (O_1673,N_24982,N_24758);
nor UO_1674 (O_1674,N_24873,N_24882);
nand UO_1675 (O_1675,N_24622,N_24544);
nand UO_1676 (O_1676,N_24913,N_24974);
or UO_1677 (O_1677,N_24754,N_24682);
nand UO_1678 (O_1678,N_24714,N_24752);
xnor UO_1679 (O_1679,N_24887,N_24742);
and UO_1680 (O_1680,N_24770,N_24930);
and UO_1681 (O_1681,N_24862,N_24754);
nand UO_1682 (O_1682,N_24819,N_24949);
xnor UO_1683 (O_1683,N_24553,N_24578);
nor UO_1684 (O_1684,N_24744,N_24760);
and UO_1685 (O_1685,N_24510,N_24648);
nand UO_1686 (O_1686,N_24691,N_24511);
or UO_1687 (O_1687,N_24706,N_24898);
nand UO_1688 (O_1688,N_24527,N_24638);
nand UO_1689 (O_1689,N_24600,N_24633);
nand UO_1690 (O_1690,N_24557,N_24642);
xnor UO_1691 (O_1691,N_24780,N_24539);
nand UO_1692 (O_1692,N_24500,N_24612);
or UO_1693 (O_1693,N_24524,N_24516);
and UO_1694 (O_1694,N_24567,N_24986);
xnor UO_1695 (O_1695,N_24763,N_24859);
or UO_1696 (O_1696,N_24846,N_24844);
or UO_1697 (O_1697,N_24550,N_24937);
or UO_1698 (O_1698,N_24974,N_24965);
or UO_1699 (O_1699,N_24606,N_24508);
nand UO_1700 (O_1700,N_24601,N_24841);
nor UO_1701 (O_1701,N_24846,N_24946);
and UO_1702 (O_1702,N_24904,N_24829);
nand UO_1703 (O_1703,N_24554,N_24633);
nand UO_1704 (O_1704,N_24576,N_24880);
nand UO_1705 (O_1705,N_24724,N_24763);
nand UO_1706 (O_1706,N_24684,N_24577);
nand UO_1707 (O_1707,N_24582,N_24734);
nand UO_1708 (O_1708,N_24724,N_24576);
nand UO_1709 (O_1709,N_24712,N_24812);
or UO_1710 (O_1710,N_24841,N_24678);
nand UO_1711 (O_1711,N_24901,N_24687);
nor UO_1712 (O_1712,N_24690,N_24856);
xor UO_1713 (O_1713,N_24685,N_24631);
nor UO_1714 (O_1714,N_24503,N_24514);
and UO_1715 (O_1715,N_24657,N_24643);
and UO_1716 (O_1716,N_24661,N_24609);
and UO_1717 (O_1717,N_24854,N_24608);
or UO_1718 (O_1718,N_24519,N_24918);
and UO_1719 (O_1719,N_24543,N_24617);
or UO_1720 (O_1720,N_24746,N_24817);
xnor UO_1721 (O_1721,N_24997,N_24744);
nor UO_1722 (O_1722,N_24929,N_24653);
or UO_1723 (O_1723,N_24625,N_24824);
and UO_1724 (O_1724,N_24802,N_24614);
xor UO_1725 (O_1725,N_24847,N_24815);
or UO_1726 (O_1726,N_24877,N_24993);
nand UO_1727 (O_1727,N_24932,N_24530);
or UO_1728 (O_1728,N_24865,N_24512);
nor UO_1729 (O_1729,N_24842,N_24508);
and UO_1730 (O_1730,N_24521,N_24608);
and UO_1731 (O_1731,N_24856,N_24639);
xnor UO_1732 (O_1732,N_24515,N_24592);
and UO_1733 (O_1733,N_24691,N_24682);
nand UO_1734 (O_1734,N_24626,N_24871);
and UO_1735 (O_1735,N_24789,N_24659);
and UO_1736 (O_1736,N_24966,N_24638);
and UO_1737 (O_1737,N_24756,N_24648);
or UO_1738 (O_1738,N_24575,N_24842);
nor UO_1739 (O_1739,N_24944,N_24544);
or UO_1740 (O_1740,N_24570,N_24832);
nand UO_1741 (O_1741,N_24686,N_24944);
and UO_1742 (O_1742,N_24706,N_24652);
nor UO_1743 (O_1743,N_24977,N_24536);
xnor UO_1744 (O_1744,N_24697,N_24924);
nor UO_1745 (O_1745,N_24619,N_24727);
and UO_1746 (O_1746,N_24570,N_24823);
or UO_1747 (O_1747,N_24722,N_24613);
xnor UO_1748 (O_1748,N_24584,N_24697);
nor UO_1749 (O_1749,N_24954,N_24773);
xor UO_1750 (O_1750,N_24802,N_24554);
or UO_1751 (O_1751,N_24507,N_24666);
nor UO_1752 (O_1752,N_24617,N_24840);
and UO_1753 (O_1753,N_24680,N_24740);
or UO_1754 (O_1754,N_24981,N_24810);
or UO_1755 (O_1755,N_24711,N_24504);
and UO_1756 (O_1756,N_24870,N_24996);
nand UO_1757 (O_1757,N_24895,N_24836);
nand UO_1758 (O_1758,N_24943,N_24587);
nor UO_1759 (O_1759,N_24767,N_24867);
and UO_1760 (O_1760,N_24508,N_24898);
and UO_1761 (O_1761,N_24750,N_24714);
xnor UO_1762 (O_1762,N_24888,N_24680);
nor UO_1763 (O_1763,N_24599,N_24561);
nand UO_1764 (O_1764,N_24553,N_24896);
xor UO_1765 (O_1765,N_24971,N_24763);
or UO_1766 (O_1766,N_24667,N_24525);
or UO_1767 (O_1767,N_24718,N_24975);
nand UO_1768 (O_1768,N_24583,N_24935);
or UO_1769 (O_1769,N_24740,N_24936);
and UO_1770 (O_1770,N_24744,N_24572);
or UO_1771 (O_1771,N_24507,N_24641);
nor UO_1772 (O_1772,N_24697,N_24513);
nor UO_1773 (O_1773,N_24931,N_24583);
or UO_1774 (O_1774,N_24695,N_24932);
nor UO_1775 (O_1775,N_24709,N_24804);
nand UO_1776 (O_1776,N_24774,N_24533);
or UO_1777 (O_1777,N_24959,N_24534);
nand UO_1778 (O_1778,N_24538,N_24919);
nor UO_1779 (O_1779,N_24848,N_24625);
xnor UO_1780 (O_1780,N_24835,N_24811);
or UO_1781 (O_1781,N_24506,N_24846);
xor UO_1782 (O_1782,N_24959,N_24520);
and UO_1783 (O_1783,N_24728,N_24769);
and UO_1784 (O_1784,N_24923,N_24930);
nand UO_1785 (O_1785,N_24545,N_24663);
xnor UO_1786 (O_1786,N_24639,N_24635);
and UO_1787 (O_1787,N_24977,N_24630);
xor UO_1788 (O_1788,N_24766,N_24921);
or UO_1789 (O_1789,N_24792,N_24986);
xor UO_1790 (O_1790,N_24817,N_24912);
xor UO_1791 (O_1791,N_24555,N_24900);
nor UO_1792 (O_1792,N_24854,N_24848);
or UO_1793 (O_1793,N_24909,N_24561);
nand UO_1794 (O_1794,N_24869,N_24614);
nand UO_1795 (O_1795,N_24976,N_24599);
xor UO_1796 (O_1796,N_24626,N_24890);
or UO_1797 (O_1797,N_24765,N_24954);
nand UO_1798 (O_1798,N_24534,N_24819);
nor UO_1799 (O_1799,N_24921,N_24590);
nor UO_1800 (O_1800,N_24653,N_24930);
or UO_1801 (O_1801,N_24611,N_24690);
xnor UO_1802 (O_1802,N_24673,N_24780);
nor UO_1803 (O_1803,N_24686,N_24748);
xor UO_1804 (O_1804,N_24901,N_24691);
and UO_1805 (O_1805,N_24629,N_24592);
xnor UO_1806 (O_1806,N_24975,N_24700);
xnor UO_1807 (O_1807,N_24591,N_24984);
and UO_1808 (O_1808,N_24585,N_24608);
nor UO_1809 (O_1809,N_24952,N_24747);
nor UO_1810 (O_1810,N_24776,N_24549);
or UO_1811 (O_1811,N_24877,N_24795);
and UO_1812 (O_1812,N_24891,N_24669);
nand UO_1813 (O_1813,N_24673,N_24593);
and UO_1814 (O_1814,N_24752,N_24660);
xnor UO_1815 (O_1815,N_24642,N_24628);
nand UO_1816 (O_1816,N_24689,N_24785);
nor UO_1817 (O_1817,N_24852,N_24649);
nor UO_1818 (O_1818,N_24903,N_24802);
and UO_1819 (O_1819,N_24590,N_24636);
or UO_1820 (O_1820,N_24591,N_24933);
nor UO_1821 (O_1821,N_24730,N_24710);
or UO_1822 (O_1822,N_24503,N_24890);
or UO_1823 (O_1823,N_24950,N_24806);
nor UO_1824 (O_1824,N_24520,N_24531);
and UO_1825 (O_1825,N_24599,N_24516);
or UO_1826 (O_1826,N_24913,N_24516);
nor UO_1827 (O_1827,N_24747,N_24843);
nand UO_1828 (O_1828,N_24969,N_24900);
and UO_1829 (O_1829,N_24750,N_24771);
and UO_1830 (O_1830,N_24553,N_24573);
xnor UO_1831 (O_1831,N_24656,N_24980);
and UO_1832 (O_1832,N_24639,N_24536);
nand UO_1833 (O_1833,N_24676,N_24662);
nor UO_1834 (O_1834,N_24666,N_24740);
nor UO_1835 (O_1835,N_24781,N_24830);
xnor UO_1836 (O_1836,N_24806,N_24829);
and UO_1837 (O_1837,N_24523,N_24571);
and UO_1838 (O_1838,N_24993,N_24507);
nor UO_1839 (O_1839,N_24814,N_24506);
xnor UO_1840 (O_1840,N_24843,N_24793);
and UO_1841 (O_1841,N_24538,N_24502);
or UO_1842 (O_1842,N_24867,N_24563);
and UO_1843 (O_1843,N_24592,N_24603);
or UO_1844 (O_1844,N_24545,N_24883);
nor UO_1845 (O_1845,N_24820,N_24746);
and UO_1846 (O_1846,N_24758,N_24572);
nor UO_1847 (O_1847,N_24961,N_24643);
nand UO_1848 (O_1848,N_24944,N_24892);
or UO_1849 (O_1849,N_24878,N_24540);
nor UO_1850 (O_1850,N_24742,N_24549);
and UO_1851 (O_1851,N_24733,N_24889);
or UO_1852 (O_1852,N_24502,N_24720);
nand UO_1853 (O_1853,N_24631,N_24908);
or UO_1854 (O_1854,N_24758,N_24804);
and UO_1855 (O_1855,N_24936,N_24652);
or UO_1856 (O_1856,N_24813,N_24848);
nand UO_1857 (O_1857,N_24523,N_24616);
nor UO_1858 (O_1858,N_24927,N_24563);
nand UO_1859 (O_1859,N_24832,N_24915);
and UO_1860 (O_1860,N_24732,N_24840);
and UO_1861 (O_1861,N_24781,N_24745);
and UO_1862 (O_1862,N_24756,N_24641);
nor UO_1863 (O_1863,N_24698,N_24560);
nand UO_1864 (O_1864,N_24738,N_24657);
nand UO_1865 (O_1865,N_24668,N_24809);
xnor UO_1866 (O_1866,N_24757,N_24566);
or UO_1867 (O_1867,N_24547,N_24649);
nor UO_1868 (O_1868,N_24981,N_24914);
xnor UO_1869 (O_1869,N_24544,N_24504);
or UO_1870 (O_1870,N_24609,N_24630);
xnor UO_1871 (O_1871,N_24907,N_24932);
xor UO_1872 (O_1872,N_24661,N_24683);
or UO_1873 (O_1873,N_24782,N_24779);
nor UO_1874 (O_1874,N_24943,N_24571);
nand UO_1875 (O_1875,N_24801,N_24623);
nand UO_1876 (O_1876,N_24965,N_24932);
xor UO_1877 (O_1877,N_24519,N_24817);
nand UO_1878 (O_1878,N_24745,N_24519);
and UO_1879 (O_1879,N_24624,N_24719);
nor UO_1880 (O_1880,N_24694,N_24878);
nand UO_1881 (O_1881,N_24737,N_24942);
nand UO_1882 (O_1882,N_24897,N_24680);
nand UO_1883 (O_1883,N_24607,N_24841);
xor UO_1884 (O_1884,N_24818,N_24932);
xnor UO_1885 (O_1885,N_24595,N_24562);
and UO_1886 (O_1886,N_24818,N_24887);
or UO_1887 (O_1887,N_24856,N_24595);
xnor UO_1888 (O_1888,N_24900,N_24629);
or UO_1889 (O_1889,N_24733,N_24769);
and UO_1890 (O_1890,N_24766,N_24761);
xor UO_1891 (O_1891,N_24902,N_24973);
and UO_1892 (O_1892,N_24555,N_24654);
nand UO_1893 (O_1893,N_24851,N_24989);
or UO_1894 (O_1894,N_24736,N_24727);
and UO_1895 (O_1895,N_24659,N_24512);
or UO_1896 (O_1896,N_24878,N_24923);
xor UO_1897 (O_1897,N_24816,N_24724);
nand UO_1898 (O_1898,N_24979,N_24831);
or UO_1899 (O_1899,N_24593,N_24709);
nand UO_1900 (O_1900,N_24663,N_24946);
nand UO_1901 (O_1901,N_24947,N_24597);
nor UO_1902 (O_1902,N_24752,N_24500);
xor UO_1903 (O_1903,N_24592,N_24510);
xor UO_1904 (O_1904,N_24899,N_24644);
xnor UO_1905 (O_1905,N_24902,N_24861);
nor UO_1906 (O_1906,N_24926,N_24601);
nor UO_1907 (O_1907,N_24659,N_24750);
nand UO_1908 (O_1908,N_24837,N_24788);
and UO_1909 (O_1909,N_24765,N_24646);
or UO_1910 (O_1910,N_24517,N_24703);
nor UO_1911 (O_1911,N_24697,N_24894);
nand UO_1912 (O_1912,N_24804,N_24590);
nor UO_1913 (O_1913,N_24885,N_24804);
xnor UO_1914 (O_1914,N_24742,N_24701);
nor UO_1915 (O_1915,N_24608,N_24570);
nand UO_1916 (O_1916,N_24960,N_24898);
xor UO_1917 (O_1917,N_24915,N_24827);
nor UO_1918 (O_1918,N_24810,N_24771);
or UO_1919 (O_1919,N_24670,N_24808);
nand UO_1920 (O_1920,N_24744,N_24509);
or UO_1921 (O_1921,N_24687,N_24984);
or UO_1922 (O_1922,N_24609,N_24954);
nor UO_1923 (O_1923,N_24677,N_24668);
nor UO_1924 (O_1924,N_24539,N_24733);
and UO_1925 (O_1925,N_24586,N_24693);
nor UO_1926 (O_1926,N_24578,N_24714);
nor UO_1927 (O_1927,N_24909,N_24650);
and UO_1928 (O_1928,N_24528,N_24985);
nand UO_1929 (O_1929,N_24672,N_24948);
and UO_1930 (O_1930,N_24752,N_24571);
nor UO_1931 (O_1931,N_24757,N_24948);
or UO_1932 (O_1932,N_24701,N_24639);
xor UO_1933 (O_1933,N_24626,N_24564);
nor UO_1934 (O_1934,N_24876,N_24994);
or UO_1935 (O_1935,N_24584,N_24743);
and UO_1936 (O_1936,N_24584,N_24802);
nor UO_1937 (O_1937,N_24938,N_24946);
nor UO_1938 (O_1938,N_24881,N_24615);
xnor UO_1939 (O_1939,N_24780,N_24846);
xor UO_1940 (O_1940,N_24795,N_24712);
xor UO_1941 (O_1941,N_24890,N_24535);
and UO_1942 (O_1942,N_24786,N_24628);
nor UO_1943 (O_1943,N_24529,N_24694);
nand UO_1944 (O_1944,N_24583,N_24854);
nor UO_1945 (O_1945,N_24737,N_24700);
or UO_1946 (O_1946,N_24726,N_24933);
and UO_1947 (O_1947,N_24660,N_24834);
or UO_1948 (O_1948,N_24574,N_24918);
or UO_1949 (O_1949,N_24976,N_24728);
xor UO_1950 (O_1950,N_24501,N_24629);
and UO_1951 (O_1951,N_24533,N_24849);
xnor UO_1952 (O_1952,N_24544,N_24593);
nor UO_1953 (O_1953,N_24644,N_24808);
nand UO_1954 (O_1954,N_24842,N_24996);
and UO_1955 (O_1955,N_24581,N_24794);
nand UO_1956 (O_1956,N_24668,N_24554);
and UO_1957 (O_1957,N_24600,N_24866);
xnor UO_1958 (O_1958,N_24896,N_24635);
nand UO_1959 (O_1959,N_24922,N_24921);
and UO_1960 (O_1960,N_24880,N_24593);
or UO_1961 (O_1961,N_24539,N_24924);
or UO_1962 (O_1962,N_24878,N_24843);
nand UO_1963 (O_1963,N_24502,N_24535);
nand UO_1964 (O_1964,N_24594,N_24863);
nor UO_1965 (O_1965,N_24800,N_24677);
nand UO_1966 (O_1966,N_24514,N_24866);
and UO_1967 (O_1967,N_24807,N_24776);
and UO_1968 (O_1968,N_24864,N_24789);
xor UO_1969 (O_1969,N_24528,N_24572);
nand UO_1970 (O_1970,N_24611,N_24654);
xor UO_1971 (O_1971,N_24781,N_24918);
and UO_1972 (O_1972,N_24692,N_24922);
nand UO_1973 (O_1973,N_24812,N_24618);
and UO_1974 (O_1974,N_24573,N_24699);
xnor UO_1975 (O_1975,N_24735,N_24952);
nor UO_1976 (O_1976,N_24516,N_24591);
and UO_1977 (O_1977,N_24833,N_24692);
xnor UO_1978 (O_1978,N_24593,N_24591);
xor UO_1979 (O_1979,N_24783,N_24738);
xnor UO_1980 (O_1980,N_24687,N_24632);
nor UO_1981 (O_1981,N_24620,N_24764);
xnor UO_1982 (O_1982,N_24623,N_24820);
nand UO_1983 (O_1983,N_24947,N_24902);
and UO_1984 (O_1984,N_24926,N_24901);
or UO_1985 (O_1985,N_24587,N_24565);
xnor UO_1986 (O_1986,N_24770,N_24999);
xor UO_1987 (O_1987,N_24826,N_24891);
xnor UO_1988 (O_1988,N_24516,N_24697);
nor UO_1989 (O_1989,N_24880,N_24907);
xnor UO_1990 (O_1990,N_24890,N_24691);
and UO_1991 (O_1991,N_24921,N_24739);
nor UO_1992 (O_1992,N_24578,N_24787);
nand UO_1993 (O_1993,N_24732,N_24503);
nand UO_1994 (O_1994,N_24653,N_24848);
nor UO_1995 (O_1995,N_24705,N_24979);
nand UO_1996 (O_1996,N_24501,N_24832);
nor UO_1997 (O_1997,N_24934,N_24608);
nand UO_1998 (O_1998,N_24980,N_24912);
nand UO_1999 (O_1999,N_24904,N_24737);
nor UO_2000 (O_2000,N_24834,N_24717);
or UO_2001 (O_2001,N_24781,N_24806);
nand UO_2002 (O_2002,N_24565,N_24839);
or UO_2003 (O_2003,N_24903,N_24676);
and UO_2004 (O_2004,N_24515,N_24987);
or UO_2005 (O_2005,N_24921,N_24715);
or UO_2006 (O_2006,N_24866,N_24604);
nor UO_2007 (O_2007,N_24884,N_24893);
nor UO_2008 (O_2008,N_24891,N_24544);
nand UO_2009 (O_2009,N_24542,N_24753);
xnor UO_2010 (O_2010,N_24826,N_24825);
nand UO_2011 (O_2011,N_24998,N_24774);
nand UO_2012 (O_2012,N_24624,N_24728);
nor UO_2013 (O_2013,N_24914,N_24576);
or UO_2014 (O_2014,N_24853,N_24721);
nor UO_2015 (O_2015,N_24574,N_24663);
or UO_2016 (O_2016,N_24572,N_24590);
nand UO_2017 (O_2017,N_24837,N_24664);
nor UO_2018 (O_2018,N_24666,N_24919);
or UO_2019 (O_2019,N_24825,N_24814);
or UO_2020 (O_2020,N_24944,N_24689);
xor UO_2021 (O_2021,N_24533,N_24925);
nor UO_2022 (O_2022,N_24920,N_24839);
nor UO_2023 (O_2023,N_24842,N_24925);
and UO_2024 (O_2024,N_24984,N_24537);
or UO_2025 (O_2025,N_24588,N_24807);
and UO_2026 (O_2026,N_24835,N_24707);
and UO_2027 (O_2027,N_24543,N_24524);
and UO_2028 (O_2028,N_24889,N_24855);
or UO_2029 (O_2029,N_24701,N_24975);
or UO_2030 (O_2030,N_24621,N_24680);
or UO_2031 (O_2031,N_24788,N_24773);
or UO_2032 (O_2032,N_24570,N_24653);
nand UO_2033 (O_2033,N_24765,N_24605);
nor UO_2034 (O_2034,N_24995,N_24835);
nand UO_2035 (O_2035,N_24746,N_24854);
or UO_2036 (O_2036,N_24721,N_24646);
and UO_2037 (O_2037,N_24766,N_24580);
nand UO_2038 (O_2038,N_24830,N_24929);
or UO_2039 (O_2039,N_24871,N_24555);
nor UO_2040 (O_2040,N_24982,N_24897);
or UO_2041 (O_2041,N_24585,N_24988);
nand UO_2042 (O_2042,N_24937,N_24910);
nor UO_2043 (O_2043,N_24609,N_24784);
nor UO_2044 (O_2044,N_24713,N_24878);
and UO_2045 (O_2045,N_24608,N_24851);
nand UO_2046 (O_2046,N_24779,N_24510);
nor UO_2047 (O_2047,N_24514,N_24778);
and UO_2048 (O_2048,N_24930,N_24761);
or UO_2049 (O_2049,N_24978,N_24810);
and UO_2050 (O_2050,N_24626,N_24620);
xor UO_2051 (O_2051,N_24724,N_24831);
nand UO_2052 (O_2052,N_24671,N_24547);
xor UO_2053 (O_2053,N_24697,N_24709);
nor UO_2054 (O_2054,N_24555,N_24899);
nand UO_2055 (O_2055,N_24617,N_24510);
and UO_2056 (O_2056,N_24840,N_24884);
and UO_2057 (O_2057,N_24631,N_24641);
xnor UO_2058 (O_2058,N_24942,N_24865);
nor UO_2059 (O_2059,N_24792,N_24757);
nor UO_2060 (O_2060,N_24727,N_24612);
and UO_2061 (O_2061,N_24934,N_24651);
nand UO_2062 (O_2062,N_24957,N_24760);
nor UO_2063 (O_2063,N_24505,N_24599);
nand UO_2064 (O_2064,N_24819,N_24539);
xnor UO_2065 (O_2065,N_24804,N_24554);
nor UO_2066 (O_2066,N_24730,N_24892);
xnor UO_2067 (O_2067,N_24743,N_24875);
nand UO_2068 (O_2068,N_24828,N_24640);
nand UO_2069 (O_2069,N_24534,N_24556);
or UO_2070 (O_2070,N_24926,N_24592);
and UO_2071 (O_2071,N_24795,N_24765);
xnor UO_2072 (O_2072,N_24782,N_24576);
and UO_2073 (O_2073,N_24955,N_24613);
xnor UO_2074 (O_2074,N_24625,N_24984);
xnor UO_2075 (O_2075,N_24807,N_24852);
nor UO_2076 (O_2076,N_24537,N_24590);
and UO_2077 (O_2077,N_24866,N_24645);
and UO_2078 (O_2078,N_24700,N_24612);
and UO_2079 (O_2079,N_24680,N_24947);
nand UO_2080 (O_2080,N_24970,N_24656);
or UO_2081 (O_2081,N_24771,N_24565);
nor UO_2082 (O_2082,N_24566,N_24932);
nor UO_2083 (O_2083,N_24965,N_24530);
and UO_2084 (O_2084,N_24739,N_24970);
xor UO_2085 (O_2085,N_24578,N_24766);
or UO_2086 (O_2086,N_24774,N_24536);
or UO_2087 (O_2087,N_24533,N_24715);
nand UO_2088 (O_2088,N_24846,N_24515);
nor UO_2089 (O_2089,N_24936,N_24754);
nor UO_2090 (O_2090,N_24575,N_24734);
nor UO_2091 (O_2091,N_24843,N_24740);
xor UO_2092 (O_2092,N_24778,N_24867);
nor UO_2093 (O_2093,N_24753,N_24528);
xnor UO_2094 (O_2094,N_24949,N_24525);
nand UO_2095 (O_2095,N_24558,N_24713);
nor UO_2096 (O_2096,N_24544,N_24921);
nor UO_2097 (O_2097,N_24949,N_24578);
nor UO_2098 (O_2098,N_24695,N_24885);
nand UO_2099 (O_2099,N_24852,N_24749);
nor UO_2100 (O_2100,N_24772,N_24896);
and UO_2101 (O_2101,N_24807,N_24986);
or UO_2102 (O_2102,N_24562,N_24999);
nand UO_2103 (O_2103,N_24687,N_24957);
nor UO_2104 (O_2104,N_24500,N_24649);
nand UO_2105 (O_2105,N_24769,N_24656);
nand UO_2106 (O_2106,N_24880,N_24929);
nor UO_2107 (O_2107,N_24829,N_24647);
or UO_2108 (O_2108,N_24618,N_24622);
nand UO_2109 (O_2109,N_24635,N_24547);
nand UO_2110 (O_2110,N_24903,N_24876);
nor UO_2111 (O_2111,N_24595,N_24566);
and UO_2112 (O_2112,N_24898,N_24685);
xor UO_2113 (O_2113,N_24785,N_24832);
nor UO_2114 (O_2114,N_24648,N_24500);
nor UO_2115 (O_2115,N_24553,N_24806);
nand UO_2116 (O_2116,N_24919,N_24580);
and UO_2117 (O_2117,N_24704,N_24975);
nand UO_2118 (O_2118,N_24760,N_24862);
and UO_2119 (O_2119,N_24826,N_24511);
xor UO_2120 (O_2120,N_24766,N_24838);
and UO_2121 (O_2121,N_24893,N_24961);
or UO_2122 (O_2122,N_24944,N_24862);
or UO_2123 (O_2123,N_24732,N_24587);
or UO_2124 (O_2124,N_24749,N_24546);
nand UO_2125 (O_2125,N_24920,N_24657);
nand UO_2126 (O_2126,N_24644,N_24803);
nand UO_2127 (O_2127,N_24753,N_24768);
nand UO_2128 (O_2128,N_24622,N_24871);
and UO_2129 (O_2129,N_24874,N_24935);
xnor UO_2130 (O_2130,N_24902,N_24726);
nor UO_2131 (O_2131,N_24695,N_24605);
nor UO_2132 (O_2132,N_24545,N_24729);
or UO_2133 (O_2133,N_24770,N_24774);
nor UO_2134 (O_2134,N_24958,N_24880);
nand UO_2135 (O_2135,N_24833,N_24961);
and UO_2136 (O_2136,N_24912,N_24612);
and UO_2137 (O_2137,N_24856,N_24817);
or UO_2138 (O_2138,N_24957,N_24653);
xor UO_2139 (O_2139,N_24638,N_24772);
xor UO_2140 (O_2140,N_24788,N_24921);
or UO_2141 (O_2141,N_24738,N_24836);
nand UO_2142 (O_2142,N_24573,N_24948);
or UO_2143 (O_2143,N_24510,N_24798);
xor UO_2144 (O_2144,N_24621,N_24871);
or UO_2145 (O_2145,N_24686,N_24590);
xor UO_2146 (O_2146,N_24858,N_24507);
or UO_2147 (O_2147,N_24700,N_24584);
or UO_2148 (O_2148,N_24713,N_24613);
xnor UO_2149 (O_2149,N_24597,N_24826);
xnor UO_2150 (O_2150,N_24628,N_24709);
and UO_2151 (O_2151,N_24836,N_24769);
nor UO_2152 (O_2152,N_24526,N_24791);
xor UO_2153 (O_2153,N_24785,N_24652);
and UO_2154 (O_2154,N_24980,N_24932);
or UO_2155 (O_2155,N_24648,N_24555);
xnor UO_2156 (O_2156,N_24615,N_24525);
nand UO_2157 (O_2157,N_24606,N_24855);
and UO_2158 (O_2158,N_24763,N_24575);
nor UO_2159 (O_2159,N_24626,N_24698);
or UO_2160 (O_2160,N_24723,N_24762);
or UO_2161 (O_2161,N_24511,N_24689);
or UO_2162 (O_2162,N_24920,N_24512);
xnor UO_2163 (O_2163,N_24742,N_24509);
xor UO_2164 (O_2164,N_24694,N_24834);
nand UO_2165 (O_2165,N_24594,N_24930);
and UO_2166 (O_2166,N_24594,N_24929);
and UO_2167 (O_2167,N_24776,N_24682);
or UO_2168 (O_2168,N_24520,N_24804);
nand UO_2169 (O_2169,N_24986,N_24898);
nor UO_2170 (O_2170,N_24777,N_24973);
or UO_2171 (O_2171,N_24588,N_24539);
and UO_2172 (O_2172,N_24838,N_24634);
and UO_2173 (O_2173,N_24902,N_24559);
xnor UO_2174 (O_2174,N_24787,N_24510);
and UO_2175 (O_2175,N_24682,N_24753);
and UO_2176 (O_2176,N_24663,N_24700);
nor UO_2177 (O_2177,N_24582,N_24796);
xor UO_2178 (O_2178,N_24605,N_24995);
and UO_2179 (O_2179,N_24587,N_24501);
nor UO_2180 (O_2180,N_24534,N_24695);
xor UO_2181 (O_2181,N_24802,N_24987);
and UO_2182 (O_2182,N_24836,N_24913);
and UO_2183 (O_2183,N_24992,N_24531);
nor UO_2184 (O_2184,N_24862,N_24967);
or UO_2185 (O_2185,N_24997,N_24797);
nand UO_2186 (O_2186,N_24921,N_24674);
xor UO_2187 (O_2187,N_24903,N_24797);
or UO_2188 (O_2188,N_24641,N_24881);
nand UO_2189 (O_2189,N_24534,N_24755);
xnor UO_2190 (O_2190,N_24986,N_24699);
nand UO_2191 (O_2191,N_24731,N_24520);
or UO_2192 (O_2192,N_24881,N_24714);
xnor UO_2193 (O_2193,N_24625,N_24612);
nor UO_2194 (O_2194,N_24826,N_24999);
nor UO_2195 (O_2195,N_24575,N_24926);
nor UO_2196 (O_2196,N_24584,N_24670);
and UO_2197 (O_2197,N_24932,N_24763);
and UO_2198 (O_2198,N_24560,N_24551);
xor UO_2199 (O_2199,N_24557,N_24545);
and UO_2200 (O_2200,N_24647,N_24553);
nand UO_2201 (O_2201,N_24827,N_24599);
and UO_2202 (O_2202,N_24520,N_24914);
and UO_2203 (O_2203,N_24523,N_24780);
nor UO_2204 (O_2204,N_24814,N_24664);
nand UO_2205 (O_2205,N_24854,N_24705);
nand UO_2206 (O_2206,N_24581,N_24980);
or UO_2207 (O_2207,N_24560,N_24690);
xnor UO_2208 (O_2208,N_24797,N_24744);
or UO_2209 (O_2209,N_24993,N_24814);
or UO_2210 (O_2210,N_24598,N_24857);
nor UO_2211 (O_2211,N_24662,N_24746);
nor UO_2212 (O_2212,N_24660,N_24753);
and UO_2213 (O_2213,N_24575,N_24704);
nand UO_2214 (O_2214,N_24912,N_24982);
nand UO_2215 (O_2215,N_24537,N_24501);
xor UO_2216 (O_2216,N_24975,N_24584);
and UO_2217 (O_2217,N_24891,N_24678);
nand UO_2218 (O_2218,N_24888,N_24911);
nor UO_2219 (O_2219,N_24782,N_24535);
and UO_2220 (O_2220,N_24959,N_24695);
nor UO_2221 (O_2221,N_24841,N_24847);
nor UO_2222 (O_2222,N_24723,N_24666);
nor UO_2223 (O_2223,N_24671,N_24804);
or UO_2224 (O_2224,N_24892,N_24685);
or UO_2225 (O_2225,N_24821,N_24640);
and UO_2226 (O_2226,N_24528,N_24740);
xnor UO_2227 (O_2227,N_24805,N_24585);
nand UO_2228 (O_2228,N_24664,N_24721);
xor UO_2229 (O_2229,N_24656,N_24681);
and UO_2230 (O_2230,N_24792,N_24709);
nand UO_2231 (O_2231,N_24684,N_24626);
nor UO_2232 (O_2232,N_24623,N_24851);
or UO_2233 (O_2233,N_24975,N_24739);
and UO_2234 (O_2234,N_24912,N_24777);
nor UO_2235 (O_2235,N_24680,N_24880);
or UO_2236 (O_2236,N_24707,N_24704);
nand UO_2237 (O_2237,N_24653,N_24824);
xor UO_2238 (O_2238,N_24821,N_24785);
nor UO_2239 (O_2239,N_24831,N_24692);
nand UO_2240 (O_2240,N_24740,N_24728);
and UO_2241 (O_2241,N_24944,N_24888);
xor UO_2242 (O_2242,N_24546,N_24808);
xor UO_2243 (O_2243,N_24578,N_24771);
nand UO_2244 (O_2244,N_24940,N_24944);
or UO_2245 (O_2245,N_24676,N_24887);
nand UO_2246 (O_2246,N_24745,N_24682);
nor UO_2247 (O_2247,N_24916,N_24833);
or UO_2248 (O_2248,N_24735,N_24518);
nor UO_2249 (O_2249,N_24596,N_24722);
or UO_2250 (O_2250,N_24635,N_24980);
nor UO_2251 (O_2251,N_24958,N_24874);
and UO_2252 (O_2252,N_24941,N_24763);
and UO_2253 (O_2253,N_24714,N_24746);
nor UO_2254 (O_2254,N_24591,N_24657);
or UO_2255 (O_2255,N_24745,N_24520);
or UO_2256 (O_2256,N_24995,N_24565);
nor UO_2257 (O_2257,N_24852,N_24848);
nand UO_2258 (O_2258,N_24908,N_24701);
nor UO_2259 (O_2259,N_24791,N_24636);
or UO_2260 (O_2260,N_24546,N_24716);
xnor UO_2261 (O_2261,N_24592,N_24753);
or UO_2262 (O_2262,N_24878,N_24949);
nand UO_2263 (O_2263,N_24599,N_24547);
xnor UO_2264 (O_2264,N_24838,N_24917);
nand UO_2265 (O_2265,N_24772,N_24948);
nor UO_2266 (O_2266,N_24690,N_24548);
and UO_2267 (O_2267,N_24882,N_24673);
or UO_2268 (O_2268,N_24888,N_24641);
and UO_2269 (O_2269,N_24561,N_24828);
nand UO_2270 (O_2270,N_24805,N_24927);
nor UO_2271 (O_2271,N_24874,N_24722);
nand UO_2272 (O_2272,N_24822,N_24508);
nand UO_2273 (O_2273,N_24894,N_24629);
and UO_2274 (O_2274,N_24932,N_24735);
nand UO_2275 (O_2275,N_24828,N_24999);
and UO_2276 (O_2276,N_24790,N_24544);
nor UO_2277 (O_2277,N_24640,N_24539);
nand UO_2278 (O_2278,N_24778,N_24734);
xor UO_2279 (O_2279,N_24785,N_24734);
nor UO_2280 (O_2280,N_24790,N_24935);
nand UO_2281 (O_2281,N_24656,N_24968);
or UO_2282 (O_2282,N_24906,N_24818);
xor UO_2283 (O_2283,N_24515,N_24939);
and UO_2284 (O_2284,N_24885,N_24849);
or UO_2285 (O_2285,N_24565,N_24745);
xor UO_2286 (O_2286,N_24830,N_24664);
nor UO_2287 (O_2287,N_24889,N_24878);
nor UO_2288 (O_2288,N_24976,N_24769);
and UO_2289 (O_2289,N_24999,N_24669);
nand UO_2290 (O_2290,N_24747,N_24943);
xor UO_2291 (O_2291,N_24601,N_24862);
nor UO_2292 (O_2292,N_24554,N_24982);
nand UO_2293 (O_2293,N_24758,N_24740);
or UO_2294 (O_2294,N_24904,N_24982);
and UO_2295 (O_2295,N_24692,N_24956);
or UO_2296 (O_2296,N_24607,N_24818);
xnor UO_2297 (O_2297,N_24968,N_24740);
and UO_2298 (O_2298,N_24910,N_24744);
xor UO_2299 (O_2299,N_24552,N_24544);
and UO_2300 (O_2300,N_24567,N_24777);
nand UO_2301 (O_2301,N_24686,N_24532);
and UO_2302 (O_2302,N_24871,N_24523);
xnor UO_2303 (O_2303,N_24722,N_24813);
xor UO_2304 (O_2304,N_24602,N_24877);
nor UO_2305 (O_2305,N_24916,N_24939);
nor UO_2306 (O_2306,N_24904,N_24734);
and UO_2307 (O_2307,N_24800,N_24956);
xor UO_2308 (O_2308,N_24691,N_24812);
or UO_2309 (O_2309,N_24841,N_24796);
and UO_2310 (O_2310,N_24691,N_24558);
nor UO_2311 (O_2311,N_24716,N_24823);
xnor UO_2312 (O_2312,N_24765,N_24526);
nor UO_2313 (O_2313,N_24559,N_24631);
nand UO_2314 (O_2314,N_24662,N_24709);
or UO_2315 (O_2315,N_24597,N_24735);
or UO_2316 (O_2316,N_24853,N_24570);
nor UO_2317 (O_2317,N_24711,N_24897);
xor UO_2318 (O_2318,N_24887,N_24834);
and UO_2319 (O_2319,N_24845,N_24932);
or UO_2320 (O_2320,N_24779,N_24761);
or UO_2321 (O_2321,N_24971,N_24999);
or UO_2322 (O_2322,N_24547,N_24920);
xor UO_2323 (O_2323,N_24735,N_24613);
or UO_2324 (O_2324,N_24851,N_24779);
nor UO_2325 (O_2325,N_24730,N_24628);
or UO_2326 (O_2326,N_24930,N_24502);
nor UO_2327 (O_2327,N_24607,N_24551);
nor UO_2328 (O_2328,N_24897,N_24677);
nor UO_2329 (O_2329,N_24556,N_24885);
nor UO_2330 (O_2330,N_24560,N_24601);
nor UO_2331 (O_2331,N_24919,N_24934);
nor UO_2332 (O_2332,N_24809,N_24907);
or UO_2333 (O_2333,N_24801,N_24691);
and UO_2334 (O_2334,N_24859,N_24947);
nor UO_2335 (O_2335,N_24608,N_24575);
nor UO_2336 (O_2336,N_24645,N_24890);
xor UO_2337 (O_2337,N_24506,N_24803);
nand UO_2338 (O_2338,N_24729,N_24915);
xnor UO_2339 (O_2339,N_24744,N_24631);
or UO_2340 (O_2340,N_24996,N_24807);
and UO_2341 (O_2341,N_24911,N_24910);
or UO_2342 (O_2342,N_24701,N_24878);
or UO_2343 (O_2343,N_24577,N_24599);
and UO_2344 (O_2344,N_24718,N_24549);
or UO_2345 (O_2345,N_24720,N_24570);
nor UO_2346 (O_2346,N_24920,N_24711);
and UO_2347 (O_2347,N_24944,N_24680);
and UO_2348 (O_2348,N_24525,N_24912);
or UO_2349 (O_2349,N_24512,N_24917);
and UO_2350 (O_2350,N_24663,N_24939);
nand UO_2351 (O_2351,N_24856,N_24994);
xnor UO_2352 (O_2352,N_24934,N_24939);
xor UO_2353 (O_2353,N_24575,N_24860);
nand UO_2354 (O_2354,N_24564,N_24792);
or UO_2355 (O_2355,N_24514,N_24977);
or UO_2356 (O_2356,N_24736,N_24908);
and UO_2357 (O_2357,N_24862,N_24547);
and UO_2358 (O_2358,N_24830,N_24708);
and UO_2359 (O_2359,N_24647,N_24512);
xor UO_2360 (O_2360,N_24630,N_24611);
and UO_2361 (O_2361,N_24699,N_24902);
nand UO_2362 (O_2362,N_24662,N_24696);
nor UO_2363 (O_2363,N_24692,N_24882);
or UO_2364 (O_2364,N_24865,N_24565);
and UO_2365 (O_2365,N_24776,N_24595);
xnor UO_2366 (O_2366,N_24706,N_24594);
and UO_2367 (O_2367,N_24503,N_24874);
xnor UO_2368 (O_2368,N_24545,N_24538);
and UO_2369 (O_2369,N_24725,N_24957);
nor UO_2370 (O_2370,N_24881,N_24933);
or UO_2371 (O_2371,N_24653,N_24619);
and UO_2372 (O_2372,N_24527,N_24593);
nand UO_2373 (O_2373,N_24532,N_24575);
xnor UO_2374 (O_2374,N_24628,N_24706);
xor UO_2375 (O_2375,N_24568,N_24541);
xor UO_2376 (O_2376,N_24924,N_24678);
nand UO_2377 (O_2377,N_24781,N_24772);
nand UO_2378 (O_2378,N_24548,N_24896);
or UO_2379 (O_2379,N_24596,N_24717);
and UO_2380 (O_2380,N_24866,N_24566);
nor UO_2381 (O_2381,N_24608,N_24819);
nor UO_2382 (O_2382,N_24669,N_24538);
or UO_2383 (O_2383,N_24828,N_24818);
nand UO_2384 (O_2384,N_24671,N_24990);
and UO_2385 (O_2385,N_24993,N_24794);
nand UO_2386 (O_2386,N_24654,N_24731);
nand UO_2387 (O_2387,N_24605,N_24693);
xnor UO_2388 (O_2388,N_24602,N_24588);
nand UO_2389 (O_2389,N_24502,N_24944);
nand UO_2390 (O_2390,N_24552,N_24895);
nand UO_2391 (O_2391,N_24942,N_24809);
nor UO_2392 (O_2392,N_24641,N_24829);
nand UO_2393 (O_2393,N_24875,N_24597);
or UO_2394 (O_2394,N_24603,N_24509);
nand UO_2395 (O_2395,N_24746,N_24651);
nor UO_2396 (O_2396,N_24611,N_24708);
and UO_2397 (O_2397,N_24847,N_24870);
and UO_2398 (O_2398,N_24673,N_24560);
xnor UO_2399 (O_2399,N_24784,N_24913);
and UO_2400 (O_2400,N_24772,N_24632);
xor UO_2401 (O_2401,N_24673,N_24989);
nand UO_2402 (O_2402,N_24529,N_24867);
xor UO_2403 (O_2403,N_24591,N_24693);
nor UO_2404 (O_2404,N_24572,N_24539);
nand UO_2405 (O_2405,N_24669,N_24766);
and UO_2406 (O_2406,N_24764,N_24646);
or UO_2407 (O_2407,N_24929,N_24689);
or UO_2408 (O_2408,N_24618,N_24970);
and UO_2409 (O_2409,N_24609,N_24867);
xnor UO_2410 (O_2410,N_24875,N_24720);
nor UO_2411 (O_2411,N_24549,N_24639);
xnor UO_2412 (O_2412,N_24756,N_24674);
or UO_2413 (O_2413,N_24884,N_24898);
xnor UO_2414 (O_2414,N_24683,N_24739);
xnor UO_2415 (O_2415,N_24550,N_24785);
or UO_2416 (O_2416,N_24975,N_24810);
or UO_2417 (O_2417,N_24774,N_24805);
nor UO_2418 (O_2418,N_24540,N_24594);
and UO_2419 (O_2419,N_24762,N_24850);
or UO_2420 (O_2420,N_24707,N_24555);
and UO_2421 (O_2421,N_24630,N_24963);
nand UO_2422 (O_2422,N_24946,N_24916);
nand UO_2423 (O_2423,N_24903,N_24943);
nand UO_2424 (O_2424,N_24809,N_24898);
or UO_2425 (O_2425,N_24789,N_24665);
nor UO_2426 (O_2426,N_24624,N_24613);
or UO_2427 (O_2427,N_24812,N_24818);
and UO_2428 (O_2428,N_24770,N_24606);
xnor UO_2429 (O_2429,N_24597,N_24508);
nand UO_2430 (O_2430,N_24870,N_24866);
xnor UO_2431 (O_2431,N_24702,N_24550);
xnor UO_2432 (O_2432,N_24980,N_24804);
nand UO_2433 (O_2433,N_24524,N_24648);
xor UO_2434 (O_2434,N_24799,N_24629);
xor UO_2435 (O_2435,N_24855,N_24838);
nand UO_2436 (O_2436,N_24597,N_24636);
nor UO_2437 (O_2437,N_24880,N_24805);
nand UO_2438 (O_2438,N_24716,N_24771);
xor UO_2439 (O_2439,N_24760,N_24780);
or UO_2440 (O_2440,N_24862,N_24551);
nand UO_2441 (O_2441,N_24642,N_24766);
nand UO_2442 (O_2442,N_24767,N_24624);
nor UO_2443 (O_2443,N_24514,N_24522);
or UO_2444 (O_2444,N_24783,N_24567);
xnor UO_2445 (O_2445,N_24962,N_24694);
and UO_2446 (O_2446,N_24904,N_24729);
and UO_2447 (O_2447,N_24654,N_24798);
nor UO_2448 (O_2448,N_24699,N_24691);
or UO_2449 (O_2449,N_24547,N_24840);
nand UO_2450 (O_2450,N_24911,N_24812);
or UO_2451 (O_2451,N_24773,N_24661);
xnor UO_2452 (O_2452,N_24795,N_24935);
nand UO_2453 (O_2453,N_24732,N_24523);
or UO_2454 (O_2454,N_24800,N_24533);
and UO_2455 (O_2455,N_24974,N_24921);
nor UO_2456 (O_2456,N_24535,N_24823);
nor UO_2457 (O_2457,N_24893,N_24964);
nor UO_2458 (O_2458,N_24692,N_24800);
and UO_2459 (O_2459,N_24888,N_24971);
xnor UO_2460 (O_2460,N_24650,N_24510);
or UO_2461 (O_2461,N_24651,N_24595);
or UO_2462 (O_2462,N_24872,N_24800);
nand UO_2463 (O_2463,N_24579,N_24800);
xnor UO_2464 (O_2464,N_24701,N_24518);
or UO_2465 (O_2465,N_24645,N_24549);
nand UO_2466 (O_2466,N_24680,N_24594);
nand UO_2467 (O_2467,N_24566,N_24792);
xnor UO_2468 (O_2468,N_24576,N_24982);
nand UO_2469 (O_2469,N_24917,N_24975);
and UO_2470 (O_2470,N_24551,N_24725);
nand UO_2471 (O_2471,N_24675,N_24994);
nand UO_2472 (O_2472,N_24650,N_24599);
nand UO_2473 (O_2473,N_24827,N_24580);
or UO_2474 (O_2474,N_24558,N_24700);
or UO_2475 (O_2475,N_24661,N_24927);
or UO_2476 (O_2476,N_24757,N_24954);
nor UO_2477 (O_2477,N_24964,N_24821);
or UO_2478 (O_2478,N_24803,N_24791);
nor UO_2479 (O_2479,N_24848,N_24518);
xor UO_2480 (O_2480,N_24692,N_24797);
xor UO_2481 (O_2481,N_24714,N_24648);
nand UO_2482 (O_2482,N_24503,N_24985);
nor UO_2483 (O_2483,N_24631,N_24574);
nor UO_2484 (O_2484,N_24582,N_24777);
and UO_2485 (O_2485,N_24603,N_24972);
xnor UO_2486 (O_2486,N_24794,N_24584);
nor UO_2487 (O_2487,N_24838,N_24518);
nand UO_2488 (O_2488,N_24763,N_24706);
xnor UO_2489 (O_2489,N_24750,N_24535);
xor UO_2490 (O_2490,N_24572,N_24934);
xnor UO_2491 (O_2491,N_24728,N_24831);
or UO_2492 (O_2492,N_24652,N_24934);
and UO_2493 (O_2493,N_24647,N_24976);
xor UO_2494 (O_2494,N_24624,N_24689);
nand UO_2495 (O_2495,N_24910,N_24573);
nand UO_2496 (O_2496,N_24572,N_24817);
xor UO_2497 (O_2497,N_24855,N_24792);
or UO_2498 (O_2498,N_24747,N_24713);
xor UO_2499 (O_2499,N_24779,N_24589);
and UO_2500 (O_2500,N_24528,N_24884);
nand UO_2501 (O_2501,N_24729,N_24695);
and UO_2502 (O_2502,N_24931,N_24792);
or UO_2503 (O_2503,N_24827,N_24523);
nor UO_2504 (O_2504,N_24520,N_24870);
and UO_2505 (O_2505,N_24742,N_24866);
nor UO_2506 (O_2506,N_24683,N_24859);
and UO_2507 (O_2507,N_24880,N_24926);
xnor UO_2508 (O_2508,N_24699,N_24703);
or UO_2509 (O_2509,N_24588,N_24663);
and UO_2510 (O_2510,N_24711,N_24529);
nor UO_2511 (O_2511,N_24972,N_24909);
and UO_2512 (O_2512,N_24962,N_24552);
nand UO_2513 (O_2513,N_24694,N_24518);
nand UO_2514 (O_2514,N_24911,N_24871);
xor UO_2515 (O_2515,N_24920,N_24852);
xor UO_2516 (O_2516,N_24867,N_24526);
and UO_2517 (O_2517,N_24514,N_24643);
nand UO_2518 (O_2518,N_24521,N_24920);
nand UO_2519 (O_2519,N_24578,N_24732);
nand UO_2520 (O_2520,N_24728,N_24920);
or UO_2521 (O_2521,N_24736,N_24795);
and UO_2522 (O_2522,N_24880,N_24968);
nor UO_2523 (O_2523,N_24502,N_24542);
or UO_2524 (O_2524,N_24680,N_24541);
and UO_2525 (O_2525,N_24919,N_24599);
xnor UO_2526 (O_2526,N_24974,N_24898);
or UO_2527 (O_2527,N_24811,N_24924);
or UO_2528 (O_2528,N_24589,N_24613);
nand UO_2529 (O_2529,N_24596,N_24999);
nor UO_2530 (O_2530,N_24840,N_24633);
nor UO_2531 (O_2531,N_24822,N_24725);
nand UO_2532 (O_2532,N_24593,N_24808);
nand UO_2533 (O_2533,N_24788,N_24502);
or UO_2534 (O_2534,N_24872,N_24505);
xnor UO_2535 (O_2535,N_24873,N_24783);
or UO_2536 (O_2536,N_24819,N_24789);
nor UO_2537 (O_2537,N_24991,N_24853);
and UO_2538 (O_2538,N_24839,N_24528);
nor UO_2539 (O_2539,N_24610,N_24867);
or UO_2540 (O_2540,N_24937,N_24982);
nor UO_2541 (O_2541,N_24611,N_24773);
xnor UO_2542 (O_2542,N_24980,N_24520);
nor UO_2543 (O_2543,N_24682,N_24990);
or UO_2544 (O_2544,N_24623,N_24887);
nor UO_2545 (O_2545,N_24813,N_24982);
xor UO_2546 (O_2546,N_24705,N_24853);
or UO_2547 (O_2547,N_24715,N_24817);
and UO_2548 (O_2548,N_24947,N_24631);
nand UO_2549 (O_2549,N_24757,N_24700);
or UO_2550 (O_2550,N_24529,N_24626);
or UO_2551 (O_2551,N_24744,N_24941);
nand UO_2552 (O_2552,N_24795,N_24873);
or UO_2553 (O_2553,N_24959,N_24699);
xor UO_2554 (O_2554,N_24886,N_24562);
nor UO_2555 (O_2555,N_24907,N_24987);
nand UO_2556 (O_2556,N_24680,N_24921);
xnor UO_2557 (O_2557,N_24950,N_24723);
and UO_2558 (O_2558,N_24736,N_24825);
xor UO_2559 (O_2559,N_24629,N_24518);
nor UO_2560 (O_2560,N_24587,N_24704);
or UO_2561 (O_2561,N_24752,N_24618);
nor UO_2562 (O_2562,N_24816,N_24850);
nand UO_2563 (O_2563,N_24762,N_24617);
xnor UO_2564 (O_2564,N_24862,N_24830);
xor UO_2565 (O_2565,N_24803,N_24909);
nand UO_2566 (O_2566,N_24717,N_24722);
nor UO_2567 (O_2567,N_24605,N_24711);
or UO_2568 (O_2568,N_24753,N_24505);
or UO_2569 (O_2569,N_24568,N_24823);
or UO_2570 (O_2570,N_24591,N_24599);
or UO_2571 (O_2571,N_24844,N_24607);
or UO_2572 (O_2572,N_24712,N_24943);
nor UO_2573 (O_2573,N_24832,N_24818);
xnor UO_2574 (O_2574,N_24512,N_24924);
nand UO_2575 (O_2575,N_24708,N_24766);
nor UO_2576 (O_2576,N_24663,N_24670);
nor UO_2577 (O_2577,N_24669,N_24544);
nand UO_2578 (O_2578,N_24567,N_24939);
nand UO_2579 (O_2579,N_24938,N_24809);
and UO_2580 (O_2580,N_24815,N_24921);
nor UO_2581 (O_2581,N_24757,N_24953);
xnor UO_2582 (O_2582,N_24521,N_24986);
xnor UO_2583 (O_2583,N_24720,N_24614);
xor UO_2584 (O_2584,N_24547,N_24627);
and UO_2585 (O_2585,N_24852,N_24893);
or UO_2586 (O_2586,N_24708,N_24811);
or UO_2587 (O_2587,N_24793,N_24964);
xor UO_2588 (O_2588,N_24876,N_24636);
nor UO_2589 (O_2589,N_24725,N_24502);
or UO_2590 (O_2590,N_24673,N_24817);
and UO_2591 (O_2591,N_24905,N_24565);
and UO_2592 (O_2592,N_24716,N_24847);
xnor UO_2593 (O_2593,N_24992,N_24764);
xnor UO_2594 (O_2594,N_24530,N_24627);
nor UO_2595 (O_2595,N_24881,N_24962);
or UO_2596 (O_2596,N_24513,N_24807);
or UO_2597 (O_2597,N_24516,N_24704);
xnor UO_2598 (O_2598,N_24808,N_24931);
nor UO_2599 (O_2599,N_24630,N_24597);
xor UO_2600 (O_2600,N_24789,N_24894);
nand UO_2601 (O_2601,N_24798,N_24607);
nand UO_2602 (O_2602,N_24914,N_24939);
or UO_2603 (O_2603,N_24536,N_24544);
and UO_2604 (O_2604,N_24625,N_24934);
and UO_2605 (O_2605,N_24735,N_24543);
nor UO_2606 (O_2606,N_24717,N_24909);
and UO_2607 (O_2607,N_24760,N_24798);
nor UO_2608 (O_2608,N_24682,N_24980);
xor UO_2609 (O_2609,N_24837,N_24688);
nand UO_2610 (O_2610,N_24939,N_24533);
nand UO_2611 (O_2611,N_24954,N_24564);
xor UO_2612 (O_2612,N_24699,N_24728);
xor UO_2613 (O_2613,N_24923,N_24633);
nor UO_2614 (O_2614,N_24779,N_24817);
nand UO_2615 (O_2615,N_24803,N_24890);
or UO_2616 (O_2616,N_24913,N_24509);
or UO_2617 (O_2617,N_24711,N_24663);
nor UO_2618 (O_2618,N_24912,N_24829);
or UO_2619 (O_2619,N_24752,N_24778);
xor UO_2620 (O_2620,N_24665,N_24900);
nand UO_2621 (O_2621,N_24828,N_24551);
or UO_2622 (O_2622,N_24684,N_24963);
or UO_2623 (O_2623,N_24540,N_24546);
and UO_2624 (O_2624,N_24953,N_24860);
or UO_2625 (O_2625,N_24552,N_24746);
or UO_2626 (O_2626,N_24742,N_24550);
or UO_2627 (O_2627,N_24731,N_24569);
nand UO_2628 (O_2628,N_24666,N_24918);
xor UO_2629 (O_2629,N_24967,N_24563);
nor UO_2630 (O_2630,N_24947,N_24739);
and UO_2631 (O_2631,N_24892,N_24868);
nor UO_2632 (O_2632,N_24937,N_24898);
xnor UO_2633 (O_2633,N_24866,N_24833);
nand UO_2634 (O_2634,N_24667,N_24528);
xor UO_2635 (O_2635,N_24933,N_24871);
nand UO_2636 (O_2636,N_24942,N_24583);
or UO_2637 (O_2637,N_24787,N_24851);
nand UO_2638 (O_2638,N_24622,N_24987);
nor UO_2639 (O_2639,N_24648,N_24540);
or UO_2640 (O_2640,N_24761,N_24916);
xnor UO_2641 (O_2641,N_24834,N_24780);
and UO_2642 (O_2642,N_24934,N_24765);
and UO_2643 (O_2643,N_24982,N_24551);
nor UO_2644 (O_2644,N_24837,N_24522);
nor UO_2645 (O_2645,N_24655,N_24676);
or UO_2646 (O_2646,N_24822,N_24660);
and UO_2647 (O_2647,N_24819,N_24926);
and UO_2648 (O_2648,N_24976,N_24807);
nor UO_2649 (O_2649,N_24578,N_24667);
and UO_2650 (O_2650,N_24707,N_24802);
and UO_2651 (O_2651,N_24526,N_24667);
nor UO_2652 (O_2652,N_24549,N_24765);
xnor UO_2653 (O_2653,N_24580,N_24879);
xor UO_2654 (O_2654,N_24502,N_24998);
nand UO_2655 (O_2655,N_24525,N_24791);
and UO_2656 (O_2656,N_24950,N_24962);
or UO_2657 (O_2657,N_24566,N_24748);
nor UO_2658 (O_2658,N_24760,N_24553);
and UO_2659 (O_2659,N_24527,N_24716);
and UO_2660 (O_2660,N_24611,N_24930);
and UO_2661 (O_2661,N_24549,N_24723);
nor UO_2662 (O_2662,N_24792,N_24756);
nor UO_2663 (O_2663,N_24774,N_24962);
and UO_2664 (O_2664,N_24631,N_24518);
or UO_2665 (O_2665,N_24741,N_24712);
or UO_2666 (O_2666,N_24543,N_24990);
nand UO_2667 (O_2667,N_24784,N_24740);
xor UO_2668 (O_2668,N_24844,N_24599);
nor UO_2669 (O_2669,N_24677,N_24550);
xor UO_2670 (O_2670,N_24938,N_24570);
nand UO_2671 (O_2671,N_24977,N_24839);
and UO_2672 (O_2672,N_24863,N_24888);
xnor UO_2673 (O_2673,N_24941,N_24860);
or UO_2674 (O_2674,N_24780,N_24638);
or UO_2675 (O_2675,N_24514,N_24767);
nor UO_2676 (O_2676,N_24659,N_24509);
or UO_2677 (O_2677,N_24812,N_24594);
and UO_2678 (O_2678,N_24873,N_24932);
xnor UO_2679 (O_2679,N_24797,N_24854);
nand UO_2680 (O_2680,N_24777,N_24983);
nand UO_2681 (O_2681,N_24848,N_24736);
xnor UO_2682 (O_2682,N_24732,N_24551);
nor UO_2683 (O_2683,N_24790,N_24802);
and UO_2684 (O_2684,N_24587,N_24915);
or UO_2685 (O_2685,N_24964,N_24565);
and UO_2686 (O_2686,N_24724,N_24627);
or UO_2687 (O_2687,N_24835,N_24862);
and UO_2688 (O_2688,N_24701,N_24746);
nand UO_2689 (O_2689,N_24854,N_24691);
or UO_2690 (O_2690,N_24783,N_24578);
xnor UO_2691 (O_2691,N_24567,N_24925);
nor UO_2692 (O_2692,N_24987,N_24839);
xnor UO_2693 (O_2693,N_24826,N_24836);
xnor UO_2694 (O_2694,N_24644,N_24845);
or UO_2695 (O_2695,N_24524,N_24515);
xor UO_2696 (O_2696,N_24716,N_24787);
nor UO_2697 (O_2697,N_24718,N_24938);
nor UO_2698 (O_2698,N_24874,N_24633);
or UO_2699 (O_2699,N_24500,N_24693);
xnor UO_2700 (O_2700,N_24649,N_24799);
nand UO_2701 (O_2701,N_24926,N_24680);
nor UO_2702 (O_2702,N_24866,N_24610);
and UO_2703 (O_2703,N_24847,N_24996);
or UO_2704 (O_2704,N_24737,N_24797);
nand UO_2705 (O_2705,N_24982,N_24920);
and UO_2706 (O_2706,N_24577,N_24871);
and UO_2707 (O_2707,N_24565,N_24811);
xnor UO_2708 (O_2708,N_24625,N_24525);
nand UO_2709 (O_2709,N_24612,N_24919);
or UO_2710 (O_2710,N_24637,N_24853);
xor UO_2711 (O_2711,N_24825,N_24705);
nand UO_2712 (O_2712,N_24764,N_24920);
or UO_2713 (O_2713,N_24845,N_24864);
and UO_2714 (O_2714,N_24704,N_24890);
xor UO_2715 (O_2715,N_24970,N_24520);
nand UO_2716 (O_2716,N_24876,N_24962);
or UO_2717 (O_2717,N_24554,N_24734);
or UO_2718 (O_2718,N_24758,N_24880);
or UO_2719 (O_2719,N_24799,N_24819);
xor UO_2720 (O_2720,N_24935,N_24914);
and UO_2721 (O_2721,N_24715,N_24870);
nor UO_2722 (O_2722,N_24636,N_24969);
nor UO_2723 (O_2723,N_24826,N_24925);
and UO_2724 (O_2724,N_24803,N_24757);
nand UO_2725 (O_2725,N_24943,N_24902);
and UO_2726 (O_2726,N_24566,N_24999);
nand UO_2727 (O_2727,N_24622,N_24713);
xor UO_2728 (O_2728,N_24933,N_24571);
nor UO_2729 (O_2729,N_24736,N_24538);
and UO_2730 (O_2730,N_24589,N_24835);
or UO_2731 (O_2731,N_24846,N_24624);
and UO_2732 (O_2732,N_24592,N_24943);
xor UO_2733 (O_2733,N_24621,N_24663);
nand UO_2734 (O_2734,N_24975,N_24729);
xor UO_2735 (O_2735,N_24526,N_24717);
or UO_2736 (O_2736,N_24560,N_24909);
or UO_2737 (O_2737,N_24650,N_24857);
and UO_2738 (O_2738,N_24753,N_24728);
and UO_2739 (O_2739,N_24532,N_24601);
nand UO_2740 (O_2740,N_24537,N_24653);
or UO_2741 (O_2741,N_24557,N_24799);
nor UO_2742 (O_2742,N_24530,N_24722);
and UO_2743 (O_2743,N_24801,N_24582);
xor UO_2744 (O_2744,N_24943,N_24839);
and UO_2745 (O_2745,N_24573,N_24905);
nor UO_2746 (O_2746,N_24727,N_24759);
xor UO_2747 (O_2747,N_24968,N_24961);
xor UO_2748 (O_2748,N_24847,N_24714);
and UO_2749 (O_2749,N_24735,N_24507);
and UO_2750 (O_2750,N_24930,N_24818);
nor UO_2751 (O_2751,N_24887,N_24781);
and UO_2752 (O_2752,N_24756,N_24805);
nand UO_2753 (O_2753,N_24565,N_24570);
nand UO_2754 (O_2754,N_24909,N_24559);
xor UO_2755 (O_2755,N_24870,N_24663);
or UO_2756 (O_2756,N_24518,N_24750);
and UO_2757 (O_2757,N_24779,N_24762);
xor UO_2758 (O_2758,N_24850,N_24613);
nand UO_2759 (O_2759,N_24867,N_24659);
nor UO_2760 (O_2760,N_24586,N_24918);
and UO_2761 (O_2761,N_24707,N_24899);
and UO_2762 (O_2762,N_24602,N_24508);
xor UO_2763 (O_2763,N_24606,N_24652);
and UO_2764 (O_2764,N_24757,N_24619);
xor UO_2765 (O_2765,N_24772,N_24890);
nor UO_2766 (O_2766,N_24735,N_24509);
xnor UO_2767 (O_2767,N_24822,N_24632);
nand UO_2768 (O_2768,N_24551,N_24743);
xnor UO_2769 (O_2769,N_24891,N_24628);
or UO_2770 (O_2770,N_24726,N_24850);
nor UO_2771 (O_2771,N_24675,N_24606);
xnor UO_2772 (O_2772,N_24862,N_24876);
nor UO_2773 (O_2773,N_24959,N_24757);
xnor UO_2774 (O_2774,N_24702,N_24788);
nor UO_2775 (O_2775,N_24551,N_24695);
nand UO_2776 (O_2776,N_24607,N_24620);
nand UO_2777 (O_2777,N_24784,N_24721);
and UO_2778 (O_2778,N_24546,N_24611);
xor UO_2779 (O_2779,N_24700,N_24886);
nor UO_2780 (O_2780,N_24536,N_24729);
or UO_2781 (O_2781,N_24832,N_24684);
nor UO_2782 (O_2782,N_24705,N_24911);
and UO_2783 (O_2783,N_24593,N_24871);
nor UO_2784 (O_2784,N_24763,N_24674);
xor UO_2785 (O_2785,N_24803,N_24511);
nand UO_2786 (O_2786,N_24881,N_24610);
or UO_2787 (O_2787,N_24665,N_24684);
and UO_2788 (O_2788,N_24872,N_24919);
and UO_2789 (O_2789,N_24567,N_24931);
or UO_2790 (O_2790,N_24976,N_24862);
or UO_2791 (O_2791,N_24540,N_24986);
nand UO_2792 (O_2792,N_24793,N_24512);
xor UO_2793 (O_2793,N_24909,N_24599);
xor UO_2794 (O_2794,N_24747,N_24889);
nor UO_2795 (O_2795,N_24597,N_24559);
and UO_2796 (O_2796,N_24701,N_24554);
or UO_2797 (O_2797,N_24734,N_24624);
nor UO_2798 (O_2798,N_24592,N_24757);
xor UO_2799 (O_2799,N_24582,N_24617);
and UO_2800 (O_2800,N_24776,N_24786);
or UO_2801 (O_2801,N_24776,N_24824);
or UO_2802 (O_2802,N_24702,N_24901);
nor UO_2803 (O_2803,N_24830,N_24684);
or UO_2804 (O_2804,N_24828,N_24648);
xnor UO_2805 (O_2805,N_24931,N_24995);
or UO_2806 (O_2806,N_24999,N_24804);
nand UO_2807 (O_2807,N_24905,N_24855);
nand UO_2808 (O_2808,N_24869,N_24586);
and UO_2809 (O_2809,N_24833,N_24997);
nor UO_2810 (O_2810,N_24566,N_24871);
xnor UO_2811 (O_2811,N_24936,N_24774);
or UO_2812 (O_2812,N_24678,N_24755);
and UO_2813 (O_2813,N_24614,N_24659);
and UO_2814 (O_2814,N_24519,N_24626);
and UO_2815 (O_2815,N_24647,N_24752);
or UO_2816 (O_2816,N_24929,N_24715);
xnor UO_2817 (O_2817,N_24994,N_24550);
and UO_2818 (O_2818,N_24641,N_24545);
and UO_2819 (O_2819,N_24927,N_24759);
nand UO_2820 (O_2820,N_24801,N_24641);
nand UO_2821 (O_2821,N_24844,N_24857);
nor UO_2822 (O_2822,N_24870,N_24824);
xnor UO_2823 (O_2823,N_24608,N_24866);
xor UO_2824 (O_2824,N_24768,N_24901);
or UO_2825 (O_2825,N_24870,N_24960);
xnor UO_2826 (O_2826,N_24690,N_24966);
and UO_2827 (O_2827,N_24775,N_24912);
xor UO_2828 (O_2828,N_24540,N_24785);
and UO_2829 (O_2829,N_24893,N_24966);
or UO_2830 (O_2830,N_24663,N_24602);
nand UO_2831 (O_2831,N_24645,N_24998);
or UO_2832 (O_2832,N_24738,N_24914);
xnor UO_2833 (O_2833,N_24836,N_24923);
nor UO_2834 (O_2834,N_24806,N_24995);
and UO_2835 (O_2835,N_24815,N_24577);
nand UO_2836 (O_2836,N_24830,N_24634);
nor UO_2837 (O_2837,N_24898,N_24866);
nand UO_2838 (O_2838,N_24827,N_24935);
nand UO_2839 (O_2839,N_24577,N_24537);
xnor UO_2840 (O_2840,N_24934,N_24928);
and UO_2841 (O_2841,N_24574,N_24717);
nand UO_2842 (O_2842,N_24529,N_24958);
or UO_2843 (O_2843,N_24952,N_24754);
xnor UO_2844 (O_2844,N_24777,N_24879);
nand UO_2845 (O_2845,N_24829,N_24627);
nor UO_2846 (O_2846,N_24814,N_24621);
nor UO_2847 (O_2847,N_24933,N_24652);
nand UO_2848 (O_2848,N_24817,N_24970);
or UO_2849 (O_2849,N_24580,N_24786);
nand UO_2850 (O_2850,N_24589,N_24872);
xnor UO_2851 (O_2851,N_24905,N_24744);
nor UO_2852 (O_2852,N_24767,N_24558);
or UO_2853 (O_2853,N_24887,N_24830);
nand UO_2854 (O_2854,N_24740,N_24552);
xnor UO_2855 (O_2855,N_24722,N_24728);
xnor UO_2856 (O_2856,N_24800,N_24791);
and UO_2857 (O_2857,N_24583,N_24650);
or UO_2858 (O_2858,N_24891,N_24535);
and UO_2859 (O_2859,N_24809,N_24970);
and UO_2860 (O_2860,N_24809,N_24956);
or UO_2861 (O_2861,N_24563,N_24889);
nand UO_2862 (O_2862,N_24809,N_24838);
nand UO_2863 (O_2863,N_24712,N_24596);
nor UO_2864 (O_2864,N_24835,N_24577);
xor UO_2865 (O_2865,N_24973,N_24578);
nor UO_2866 (O_2866,N_24526,N_24610);
xnor UO_2867 (O_2867,N_24615,N_24617);
xor UO_2868 (O_2868,N_24988,N_24987);
and UO_2869 (O_2869,N_24920,N_24841);
nand UO_2870 (O_2870,N_24728,N_24579);
nand UO_2871 (O_2871,N_24674,N_24920);
or UO_2872 (O_2872,N_24703,N_24819);
or UO_2873 (O_2873,N_24906,N_24841);
nand UO_2874 (O_2874,N_24720,N_24804);
nand UO_2875 (O_2875,N_24588,N_24563);
xnor UO_2876 (O_2876,N_24723,N_24758);
nor UO_2877 (O_2877,N_24640,N_24918);
or UO_2878 (O_2878,N_24919,N_24938);
or UO_2879 (O_2879,N_24943,N_24686);
and UO_2880 (O_2880,N_24870,N_24579);
xor UO_2881 (O_2881,N_24602,N_24680);
nor UO_2882 (O_2882,N_24792,N_24633);
nand UO_2883 (O_2883,N_24529,N_24940);
and UO_2884 (O_2884,N_24950,N_24694);
nor UO_2885 (O_2885,N_24951,N_24720);
and UO_2886 (O_2886,N_24898,N_24675);
nor UO_2887 (O_2887,N_24781,N_24890);
nor UO_2888 (O_2888,N_24575,N_24614);
xor UO_2889 (O_2889,N_24933,N_24944);
nand UO_2890 (O_2890,N_24917,N_24710);
or UO_2891 (O_2891,N_24741,N_24871);
nand UO_2892 (O_2892,N_24636,N_24849);
or UO_2893 (O_2893,N_24878,N_24788);
or UO_2894 (O_2894,N_24714,N_24593);
and UO_2895 (O_2895,N_24703,N_24727);
nand UO_2896 (O_2896,N_24579,N_24764);
or UO_2897 (O_2897,N_24776,N_24951);
nand UO_2898 (O_2898,N_24576,N_24973);
nand UO_2899 (O_2899,N_24756,N_24649);
or UO_2900 (O_2900,N_24620,N_24767);
nor UO_2901 (O_2901,N_24858,N_24705);
xnor UO_2902 (O_2902,N_24724,N_24683);
nor UO_2903 (O_2903,N_24647,N_24972);
or UO_2904 (O_2904,N_24955,N_24699);
or UO_2905 (O_2905,N_24554,N_24783);
nor UO_2906 (O_2906,N_24655,N_24597);
nor UO_2907 (O_2907,N_24843,N_24981);
xor UO_2908 (O_2908,N_24882,N_24914);
nand UO_2909 (O_2909,N_24920,N_24773);
xor UO_2910 (O_2910,N_24862,N_24667);
and UO_2911 (O_2911,N_24512,N_24667);
nor UO_2912 (O_2912,N_24623,N_24690);
nand UO_2913 (O_2913,N_24649,N_24630);
xnor UO_2914 (O_2914,N_24948,N_24565);
xor UO_2915 (O_2915,N_24954,N_24863);
nor UO_2916 (O_2916,N_24588,N_24676);
and UO_2917 (O_2917,N_24858,N_24765);
and UO_2918 (O_2918,N_24761,N_24995);
nor UO_2919 (O_2919,N_24754,N_24724);
and UO_2920 (O_2920,N_24733,N_24545);
and UO_2921 (O_2921,N_24828,N_24968);
nor UO_2922 (O_2922,N_24632,N_24569);
nor UO_2923 (O_2923,N_24859,N_24580);
nor UO_2924 (O_2924,N_24647,N_24908);
or UO_2925 (O_2925,N_24931,N_24872);
or UO_2926 (O_2926,N_24787,N_24918);
nor UO_2927 (O_2927,N_24590,N_24592);
xnor UO_2928 (O_2928,N_24785,N_24691);
nor UO_2929 (O_2929,N_24639,N_24936);
and UO_2930 (O_2930,N_24551,N_24875);
or UO_2931 (O_2931,N_24964,N_24568);
or UO_2932 (O_2932,N_24545,N_24594);
xor UO_2933 (O_2933,N_24852,N_24615);
xor UO_2934 (O_2934,N_24689,N_24784);
or UO_2935 (O_2935,N_24526,N_24531);
xnor UO_2936 (O_2936,N_24783,N_24735);
xor UO_2937 (O_2937,N_24964,N_24638);
nor UO_2938 (O_2938,N_24807,N_24963);
xor UO_2939 (O_2939,N_24661,N_24549);
and UO_2940 (O_2940,N_24678,N_24711);
or UO_2941 (O_2941,N_24667,N_24865);
xnor UO_2942 (O_2942,N_24526,N_24953);
or UO_2943 (O_2943,N_24707,N_24881);
xnor UO_2944 (O_2944,N_24725,N_24887);
and UO_2945 (O_2945,N_24851,N_24528);
nand UO_2946 (O_2946,N_24538,N_24855);
xnor UO_2947 (O_2947,N_24695,N_24694);
or UO_2948 (O_2948,N_24778,N_24946);
nand UO_2949 (O_2949,N_24762,N_24618);
and UO_2950 (O_2950,N_24942,N_24922);
nor UO_2951 (O_2951,N_24832,N_24773);
xor UO_2952 (O_2952,N_24858,N_24739);
nor UO_2953 (O_2953,N_24736,N_24987);
or UO_2954 (O_2954,N_24581,N_24771);
or UO_2955 (O_2955,N_24696,N_24780);
and UO_2956 (O_2956,N_24650,N_24769);
or UO_2957 (O_2957,N_24946,N_24827);
or UO_2958 (O_2958,N_24617,N_24575);
xnor UO_2959 (O_2959,N_24569,N_24891);
or UO_2960 (O_2960,N_24559,N_24900);
xor UO_2961 (O_2961,N_24812,N_24962);
and UO_2962 (O_2962,N_24673,N_24595);
or UO_2963 (O_2963,N_24532,N_24514);
nor UO_2964 (O_2964,N_24961,N_24977);
nor UO_2965 (O_2965,N_24533,N_24749);
and UO_2966 (O_2966,N_24543,N_24864);
and UO_2967 (O_2967,N_24831,N_24792);
nand UO_2968 (O_2968,N_24636,N_24826);
or UO_2969 (O_2969,N_24827,N_24973);
and UO_2970 (O_2970,N_24682,N_24710);
xnor UO_2971 (O_2971,N_24789,N_24832);
or UO_2972 (O_2972,N_24810,N_24526);
or UO_2973 (O_2973,N_24972,N_24808);
nand UO_2974 (O_2974,N_24515,N_24878);
nand UO_2975 (O_2975,N_24761,N_24820);
and UO_2976 (O_2976,N_24677,N_24741);
nand UO_2977 (O_2977,N_24867,N_24908);
nor UO_2978 (O_2978,N_24687,N_24665);
nor UO_2979 (O_2979,N_24506,N_24625);
and UO_2980 (O_2980,N_24930,N_24964);
nor UO_2981 (O_2981,N_24638,N_24572);
nor UO_2982 (O_2982,N_24813,N_24611);
or UO_2983 (O_2983,N_24821,N_24906);
nor UO_2984 (O_2984,N_24953,N_24719);
nand UO_2985 (O_2985,N_24803,N_24564);
nand UO_2986 (O_2986,N_24946,N_24933);
or UO_2987 (O_2987,N_24567,N_24928);
or UO_2988 (O_2988,N_24674,N_24706);
xor UO_2989 (O_2989,N_24501,N_24901);
or UO_2990 (O_2990,N_24697,N_24736);
xor UO_2991 (O_2991,N_24706,N_24694);
nand UO_2992 (O_2992,N_24972,N_24838);
or UO_2993 (O_2993,N_24762,N_24594);
xnor UO_2994 (O_2994,N_24701,N_24946);
xnor UO_2995 (O_2995,N_24607,N_24995);
and UO_2996 (O_2996,N_24620,N_24900);
nand UO_2997 (O_2997,N_24529,N_24579);
and UO_2998 (O_2998,N_24741,N_24558);
xnor UO_2999 (O_2999,N_24998,N_24603);
endmodule