module basic_2500_25000_3000_125_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_833,In_577);
and U1 (N_1,In_408,In_778);
or U2 (N_2,In_1616,In_649);
or U3 (N_3,In_544,In_1940);
nor U4 (N_4,In_154,In_1949);
nor U5 (N_5,In_1208,In_1202);
and U6 (N_6,In_1061,In_821);
or U7 (N_7,In_105,In_921);
or U8 (N_8,In_2212,In_362);
and U9 (N_9,In_1529,In_622);
nor U10 (N_10,In_1994,In_911);
nand U11 (N_11,In_2392,In_78);
or U12 (N_12,In_1337,In_2209);
nor U13 (N_13,In_487,In_2373);
and U14 (N_14,In_2383,In_576);
nor U15 (N_15,In_1967,In_218);
or U16 (N_16,In_1142,In_2476);
nor U17 (N_17,In_2360,In_45);
nor U18 (N_18,In_2498,In_1565);
and U19 (N_19,In_2322,In_1872);
nor U20 (N_20,In_1917,In_2204);
or U21 (N_21,In_1423,In_694);
and U22 (N_22,In_514,In_1245);
or U23 (N_23,In_231,In_667);
or U24 (N_24,In_1653,In_860);
nand U25 (N_25,In_438,In_1100);
nand U26 (N_26,In_799,In_555);
nand U27 (N_27,In_2479,In_181);
or U28 (N_28,In_1329,In_1869);
or U29 (N_29,In_1422,In_25);
and U30 (N_30,In_779,In_1841);
nand U31 (N_31,In_197,In_542);
and U32 (N_32,In_2012,In_2188);
nor U33 (N_33,In_2077,In_342);
nand U34 (N_34,In_1961,In_2251);
nor U35 (N_35,In_1448,In_52);
and U36 (N_36,In_2494,In_334);
or U37 (N_37,In_1235,In_171);
nand U38 (N_38,In_1608,In_2279);
nand U39 (N_39,In_1186,In_1993);
nand U40 (N_40,In_769,In_1705);
or U41 (N_41,In_2300,In_1192);
and U42 (N_42,In_612,In_807);
nor U43 (N_43,In_2109,In_1487);
nand U44 (N_44,In_1319,In_1982);
and U45 (N_45,In_282,In_2018);
nor U46 (N_46,In_2369,In_286);
nand U47 (N_47,In_1883,In_1720);
and U48 (N_48,In_793,In_1861);
nor U49 (N_49,In_364,In_2223);
nor U50 (N_50,In_2100,In_1758);
or U51 (N_51,In_463,In_2217);
or U52 (N_52,In_431,In_2073);
nand U53 (N_53,In_843,In_1643);
nand U54 (N_54,In_1385,In_2182);
nor U55 (N_55,In_1988,In_589);
or U56 (N_56,In_2296,In_272);
and U57 (N_57,In_764,In_1928);
and U58 (N_58,In_497,In_521);
nand U59 (N_59,In_24,In_1727);
nand U60 (N_60,In_955,In_855);
nand U61 (N_61,In_685,In_1991);
nor U62 (N_62,In_1469,In_1747);
and U63 (N_63,In_9,In_1766);
nand U64 (N_64,In_2291,In_1969);
nand U65 (N_65,In_977,In_1849);
nand U66 (N_66,In_363,In_459);
and U67 (N_67,In_88,In_652);
or U68 (N_68,In_2004,In_787);
or U69 (N_69,In_810,In_2189);
nand U70 (N_70,In_2164,In_1101);
or U71 (N_71,In_991,In_1382);
nand U72 (N_72,In_691,In_2042);
nand U73 (N_73,In_1343,In_2178);
and U74 (N_74,In_829,In_590);
nor U75 (N_75,In_1907,In_189);
nor U76 (N_76,In_639,In_403);
nand U77 (N_77,In_376,In_191);
and U78 (N_78,In_1615,In_1791);
and U79 (N_79,In_2332,In_321);
nand U80 (N_80,In_15,In_1012);
or U81 (N_81,In_2440,In_1312);
or U82 (N_82,In_222,In_2314);
nor U83 (N_83,In_2493,In_2441);
nor U84 (N_84,In_1203,In_2427);
nor U85 (N_85,In_1297,In_1730);
or U86 (N_86,In_1158,In_2413);
nor U87 (N_87,In_184,In_2348);
or U88 (N_88,In_1145,In_1147);
nand U89 (N_89,In_2031,In_1318);
nand U90 (N_90,In_1217,In_1259);
or U91 (N_91,In_1115,In_512);
nor U92 (N_92,In_611,In_1335);
or U93 (N_93,In_2231,In_2305);
nand U94 (N_94,In_1496,In_2262);
nand U95 (N_95,In_1709,In_842);
nand U96 (N_96,In_2264,In_1160);
and U97 (N_97,In_389,In_588);
or U98 (N_98,In_699,In_1294);
xnor U99 (N_99,In_1104,In_1067);
and U100 (N_100,In_1708,In_1728);
or U101 (N_101,In_2410,In_1621);
nand U102 (N_102,In_1472,In_1211);
or U103 (N_103,In_2245,In_526);
nand U104 (N_104,In_396,In_398);
nand U105 (N_105,In_1692,In_934);
nor U106 (N_106,In_304,In_1904);
nand U107 (N_107,In_1131,In_2066);
and U108 (N_108,In_1953,In_1734);
or U109 (N_109,In_425,In_624);
and U110 (N_110,In_1739,In_1984);
nand U111 (N_111,In_2345,In_1999);
nor U112 (N_112,In_199,In_1786);
and U113 (N_113,In_618,In_637);
nor U114 (N_114,In_739,In_2453);
nand U115 (N_115,In_194,In_655);
nand U116 (N_116,In_1336,In_872);
nor U117 (N_117,In_1305,In_580);
nor U118 (N_118,In_695,In_1238);
and U119 (N_119,In_2026,In_781);
nand U120 (N_120,In_1572,In_236);
or U121 (N_121,In_1626,In_2450);
or U122 (N_122,In_2195,In_1645);
and U123 (N_123,In_2108,In_1687);
nor U124 (N_124,In_1224,In_1398);
nand U125 (N_125,In_1702,In_40);
nor U126 (N_126,In_1772,In_1710);
or U127 (N_127,In_2495,In_758);
or U128 (N_128,In_887,In_2497);
nor U129 (N_129,In_2342,In_2478);
nor U130 (N_130,In_66,In_1241);
nand U131 (N_131,In_2320,In_1926);
or U132 (N_132,In_491,In_1737);
and U133 (N_133,In_920,In_1668);
nand U134 (N_134,In_7,In_460);
nor U135 (N_135,In_566,In_1461);
or U136 (N_136,In_1252,In_2078);
nand U137 (N_137,In_702,In_583);
nor U138 (N_138,In_2139,In_1954);
nor U139 (N_139,In_1411,In_1395);
or U140 (N_140,In_615,In_2242);
nor U141 (N_141,In_1020,In_1860);
and U142 (N_142,In_2101,In_2040);
or U143 (N_143,In_482,In_516);
nand U144 (N_144,In_992,In_2379);
nor U145 (N_145,In_503,In_76);
nand U146 (N_146,In_405,In_1644);
nand U147 (N_147,In_1001,In_2086);
nand U148 (N_148,In_1146,In_241);
nor U149 (N_149,In_136,In_1344);
or U150 (N_150,In_816,In_2458);
nand U151 (N_151,In_504,In_960);
nor U152 (N_152,In_414,In_1268);
nor U153 (N_153,In_1512,In_628);
and U154 (N_154,In_493,In_182);
nor U155 (N_155,In_323,In_1015);
nand U156 (N_156,In_1435,In_610);
and U157 (N_157,In_868,In_211);
nand U158 (N_158,In_2404,In_735);
or U159 (N_159,In_1361,In_257);
nor U160 (N_160,In_1414,In_1918);
nand U161 (N_161,In_578,In_1074);
and U162 (N_162,In_2187,In_1378);
nor U163 (N_163,In_2033,In_1449);
or U164 (N_164,In_956,In_1484);
and U165 (N_165,In_2420,In_2225);
and U166 (N_166,In_1379,In_951);
or U167 (N_167,In_159,In_1955);
nor U168 (N_168,In_2173,In_2341);
and U169 (N_169,In_1591,In_243);
nand U170 (N_170,In_1190,In_294);
and U171 (N_171,In_1602,In_748);
and U172 (N_172,In_1286,In_1228);
nand U173 (N_173,In_4,In_1108);
and U174 (N_174,In_1083,In_886);
and U175 (N_175,In_1106,In_2051);
xor U176 (N_176,In_745,In_1025);
nor U177 (N_177,In_2290,In_308);
xor U178 (N_178,In_114,In_902);
nor U179 (N_179,In_3,In_1938);
or U180 (N_180,In_1444,In_1059);
nor U181 (N_181,In_486,In_2009);
and U182 (N_182,In_1912,In_1442);
nor U183 (N_183,In_1897,In_708);
or U184 (N_184,In_1165,In_721);
nand U185 (N_185,In_1409,In_791);
nor U186 (N_186,In_1139,In_123);
nor U187 (N_187,In_770,In_891);
nand U188 (N_188,In_1289,In_82);
nor U189 (N_189,In_2435,In_269);
nand U190 (N_190,In_744,In_1497);
nand U191 (N_191,In_1221,In_982);
nor U192 (N_192,In_1604,In_1298);
nor U193 (N_193,In_680,In_2390);
or U194 (N_194,In_1769,In_1227);
nor U195 (N_195,In_2130,In_2003);
or U196 (N_196,In_1826,In_1486);
nand U197 (N_197,In_1743,In_2255);
nor U198 (N_198,In_1871,In_756);
nor U199 (N_199,In_1813,In_994);
nand U200 (N_200,In_742,In_1779);
nand U201 (N_201,In_264,In_1296);
or U202 (N_202,N_166,In_2105);
nor U203 (N_203,In_234,In_1367);
and U204 (N_204,In_1478,In_1845);
nand U205 (N_205,In_1506,In_621);
and U206 (N_206,In_1882,N_87);
or U207 (N_207,In_2277,In_1617);
nand U208 (N_208,In_2093,In_2213);
nor U209 (N_209,In_1915,In_2253);
and U210 (N_210,In_146,In_1452);
nand U211 (N_211,N_68,In_100);
and U212 (N_212,N_155,In_185);
nand U213 (N_213,N_160,In_677);
or U214 (N_214,In_18,In_550);
nor U215 (N_215,In_2241,In_444);
nor U216 (N_216,In_523,In_2252);
and U217 (N_217,In_1008,In_1886);
and U218 (N_218,N_126,In_1263);
nand U219 (N_219,N_28,In_1096);
or U220 (N_220,In_926,In_1076);
nand U221 (N_221,In_1253,In_881);
nand U222 (N_222,In_897,In_1426);
and U223 (N_223,In_1117,N_34);
and U224 (N_224,In_1153,In_495);
nor U225 (N_225,In_1906,In_68);
nor U226 (N_226,In_210,In_889);
and U227 (N_227,In_736,N_168);
or U228 (N_228,In_151,In_2168);
and U229 (N_229,In_1574,In_1630);
and U230 (N_230,In_229,In_1729);
and U231 (N_231,In_545,In_79);
and U232 (N_232,In_2125,In_2153);
nor U233 (N_233,In_638,In_77);
or U234 (N_234,In_1119,In_174);
and U235 (N_235,In_1243,In_524);
and U236 (N_236,In_2468,N_4);
and U237 (N_237,In_2271,In_988);
and U238 (N_238,In_1821,In_73);
nor U239 (N_239,In_1544,In_2384);
or U240 (N_240,In_2488,In_1471);
nor U241 (N_241,In_360,In_119);
and U242 (N_242,In_274,In_947);
nor U243 (N_243,N_51,In_1292);
or U244 (N_244,In_604,In_2315);
nor U245 (N_245,In_217,In_733);
nor U246 (N_246,In_2025,In_761);
nor U247 (N_247,In_270,In_98);
nand U248 (N_248,In_375,In_666);
nand U249 (N_249,In_1995,In_1855);
nor U250 (N_250,In_2483,In_1844);
or U251 (N_251,In_922,In_1971);
or U252 (N_252,In_2050,In_2247);
nand U253 (N_253,In_2462,In_135);
nand U254 (N_254,In_1479,In_630);
nand U255 (N_255,In_1102,In_2470);
or U256 (N_256,In_300,N_62);
nand U257 (N_257,In_147,In_2287);
or U258 (N_258,In_1019,In_1642);
nand U259 (N_259,In_2049,N_82);
or U260 (N_260,In_267,In_1375);
nor U261 (N_261,In_957,In_1612);
nand U262 (N_262,In_1780,In_1016);
or U263 (N_263,N_110,In_161);
or U264 (N_264,In_971,In_2380);
nor U265 (N_265,In_832,In_2371);
nand U266 (N_266,In_696,In_1870);
nand U267 (N_267,In_2196,In_58);
and U268 (N_268,N_21,In_1919);
nor U269 (N_269,In_1688,In_2344);
and U270 (N_270,In_1814,In_1762);
nand U271 (N_271,In_475,In_1637);
and U272 (N_272,In_1771,In_2285);
nand U273 (N_273,In_1859,In_1966);
or U274 (N_274,In_1194,In_2375);
nand U275 (N_275,In_1418,In_1427);
or U276 (N_276,In_1686,N_134);
nor U277 (N_277,In_1032,In_1068);
nand U278 (N_278,In_1164,In_23);
nand U279 (N_279,In_1664,In_1287);
nor U280 (N_280,In_1552,In_1460);
or U281 (N_281,N_111,In_2334);
nor U282 (N_282,N_147,In_723);
or U283 (N_283,In_775,In_731);
nand U284 (N_284,In_941,In_1364);
nor U285 (N_285,In_502,In_1090);
or U286 (N_286,In_232,In_844);
nor U287 (N_287,In_2218,In_1658);
or U288 (N_288,In_266,In_1371);
nor U289 (N_289,In_1468,In_2349);
nor U290 (N_290,In_1459,In_538);
nand U291 (N_291,In_1789,In_1451);
and U292 (N_292,In_1921,In_386);
nand U293 (N_293,In_1261,In_2183);
and U294 (N_294,N_199,In_1755);
nand U295 (N_295,In_1233,In_1521);
and U296 (N_296,In_297,In_2240);
nor U297 (N_297,In_490,In_824);
and U298 (N_298,In_1187,In_1856);
and U299 (N_299,In_1745,In_1528);
xor U300 (N_300,In_647,In_1910);
or U301 (N_301,In_2013,N_27);
or U302 (N_302,In_1500,In_543);
or U303 (N_303,In_187,In_158);
nor U304 (N_304,In_1669,In_1788);
and U305 (N_305,In_1050,In_511);
nor U306 (N_306,In_468,In_87);
and U307 (N_307,In_1156,In_1639);
nor U308 (N_308,In_1663,In_1925);
or U309 (N_309,In_1601,In_533);
nor U310 (N_310,In_600,N_167);
nor U311 (N_311,In_1566,In_380);
nand U312 (N_312,In_1097,In_1588);
nor U313 (N_313,N_156,In_1952);
or U314 (N_314,In_551,N_47);
nor U315 (N_315,In_395,In_1774);
or U316 (N_316,In_1080,In_2323);
or U317 (N_317,In_296,In_1873);
nor U318 (N_318,In_716,In_1699);
nor U319 (N_319,In_1597,In_130);
nand U320 (N_320,In_1892,In_1118);
and U321 (N_321,In_1392,In_2146);
nand U322 (N_322,In_1569,In_928);
and U323 (N_323,In_1944,In_290);
nor U324 (N_324,In_1081,N_101);
nor U325 (N_325,In_1888,In_1432);
or U326 (N_326,In_2472,In_2317);
or U327 (N_327,In_216,In_950);
or U328 (N_328,In_295,In_1126);
nor U329 (N_329,In_1679,N_63);
nor U330 (N_330,In_1741,In_1004);
nand U331 (N_331,In_1620,In_2457);
nor U332 (N_332,In_738,In_763);
and U333 (N_333,In_1443,N_11);
or U334 (N_334,In_1429,In_2079);
nand U335 (N_335,In_230,In_355);
nor U336 (N_336,N_59,In_2327);
nor U337 (N_337,In_1748,In_530);
nor U338 (N_338,In_1124,In_894);
and U339 (N_339,In_1537,In_1776);
and U340 (N_340,In_857,In_2363);
and U341 (N_341,N_198,In_806);
nor U342 (N_342,In_2274,In_640);
and U343 (N_343,In_1144,In_340);
nand U344 (N_344,In_773,In_1532);
and U345 (N_345,In_1510,In_1561);
nor U346 (N_346,In_2112,In_676);
and U347 (N_347,In_1136,In_2133);
or U348 (N_348,In_1111,N_159);
and U349 (N_349,In_1689,In_1030);
or U350 (N_350,In_2198,In_237);
nor U351 (N_351,In_1998,In_2214);
nor U352 (N_352,In_743,In_1802);
and U353 (N_353,In_1633,N_127);
or U354 (N_354,In_1848,In_1899);
nand U355 (N_355,In_620,N_100);
nor U356 (N_356,N_152,In_57);
nand U357 (N_357,N_123,In_552);
xnor U358 (N_358,In_1718,In_97);
or U359 (N_359,In_1191,In_1070);
nor U360 (N_360,In_394,In_741);
or U361 (N_361,In_1764,In_69);
nand U362 (N_362,In_287,In_265);
nand U363 (N_363,In_1666,In_1948);
nor U364 (N_364,In_2162,In_506);
or U365 (N_365,In_1738,In_795);
or U366 (N_366,In_548,In_1437);
nor U367 (N_367,In_2303,In_1488);
and U368 (N_368,In_301,In_121);
nor U369 (N_369,In_1933,In_567);
nor U370 (N_370,In_268,In_406);
nor U371 (N_371,In_2163,In_75);
nor U372 (N_372,In_2313,In_454);
nand U373 (N_373,In_1960,In_2286);
and U374 (N_374,N_132,N_31);
nor U375 (N_375,In_8,In_1744);
nor U376 (N_376,In_379,In_1505);
nor U377 (N_377,In_1338,In_21);
nor U378 (N_378,In_71,In_2176);
or U379 (N_379,In_796,In_707);
nand U380 (N_380,In_1750,N_108);
or U381 (N_381,In_1567,In_1244);
nor U382 (N_382,In_1697,In_255);
nand U383 (N_383,In_1977,In_423);
or U384 (N_384,In_867,In_2043);
nor U385 (N_385,In_420,In_2455);
nand U386 (N_386,In_927,N_70);
and U387 (N_387,In_1333,In_285);
and U388 (N_388,In_1322,In_1943);
and U389 (N_389,In_1924,In_1400);
and U390 (N_390,In_1308,In_1033);
or U391 (N_391,In_1481,In_800);
nor U392 (N_392,In_1576,In_348);
nor U393 (N_393,In_209,In_93);
nand U394 (N_394,In_678,N_124);
nor U395 (N_395,In_1373,N_189);
and U396 (N_396,In_441,In_333);
nand U397 (N_397,N_102,In_276);
or U398 (N_398,In_2090,In_986);
nor U399 (N_399,In_574,In_416);
nand U400 (N_400,In_5,In_1985);
and U401 (N_401,In_38,In_2350);
nor U402 (N_402,In_623,In_2280);
nor U403 (N_403,In_1498,In_325);
and U404 (N_404,In_834,In_2382);
nand U405 (N_405,In_1315,In_2408);
and U406 (N_406,N_107,In_385);
and U407 (N_407,In_1386,In_785);
nand U408 (N_408,In_2008,In_349);
nand U409 (N_409,In_1133,In_115);
or U410 (N_410,In_1733,In_1857);
and U411 (N_411,In_593,In_359);
or U412 (N_412,In_985,In_1210);
nor U413 (N_413,N_224,N_240);
or U414 (N_414,N_92,In_2421);
nand U415 (N_415,In_1480,In_2210);
and U416 (N_416,N_86,In_2473);
or U417 (N_417,In_2486,N_317);
nor U418 (N_418,In_1260,N_360);
or U419 (N_419,N_311,In_718);
xnor U420 (N_420,In_2160,In_312);
or U421 (N_421,N_364,In_1514);
nor U422 (N_422,In_2368,In_1874);
nand U423 (N_423,In_1321,In_1204);
or U424 (N_424,In_2268,In_1575);
nor U425 (N_425,N_251,N_273);
nand U426 (N_426,In_306,In_248);
and U427 (N_427,In_2122,N_210);
nor U428 (N_428,N_359,In_2481);
nor U429 (N_429,In_1800,In_317);
or U430 (N_430,In_898,In_2325);
nor U431 (N_431,In_2249,In_433);
nand U432 (N_432,In_2174,In_726);
nor U433 (N_433,In_2131,In_1018);
or U434 (N_434,In_1060,In_1526);
nand U435 (N_435,In_483,In_1179);
or U436 (N_436,In_1794,N_384);
and U437 (N_437,In_1503,In_2069);
or U438 (N_438,In_239,In_2299);
and U439 (N_439,N_24,In_609);
or U440 (N_440,In_126,In_1970);
nand U441 (N_441,In_2124,In_1958);
nor U442 (N_442,In_1288,N_347);
nor U443 (N_443,N_18,In_1513);
nor U444 (N_444,N_381,N_386);
nand U445 (N_445,N_348,In_173);
nand U446 (N_446,In_865,In_2035);
or U447 (N_447,In_2094,In_56);
nor U448 (N_448,N_60,In_125);
nand U449 (N_449,In_2396,N_308);
nor U450 (N_450,In_1041,N_2);
nand U451 (N_451,In_81,In_1258);
nand U452 (N_452,In_457,N_125);
or U453 (N_453,In_1058,In_1600);
nor U454 (N_454,In_1129,In_2418);
or U455 (N_455,In_582,In_427);
or U456 (N_456,In_365,In_2104);
or U457 (N_457,In_603,In_535);
nand U458 (N_458,N_307,In_1717);
or U459 (N_459,In_1089,In_1013);
nor U460 (N_460,In_1223,In_108);
and U461 (N_461,In_2443,In_1754);
nor U462 (N_462,In_1868,In_1197);
nand U463 (N_463,In_1225,In_2005);
nor U464 (N_464,In_1279,In_1670);
and U465 (N_465,In_1055,In_1785);
nand U466 (N_466,N_378,In_651);
or U467 (N_467,In_607,N_323);
nand U468 (N_468,In_1078,In_2063);
and U469 (N_469,In_1300,In_1130);
nand U470 (N_470,In_1834,In_1307);
nor U471 (N_471,N_93,N_339);
nand U472 (N_472,In_2192,In_2097);
and U473 (N_473,N_276,In_109);
and U474 (N_474,In_474,In_1775);
nor U475 (N_475,In_179,In_1370);
and U476 (N_476,In_1934,In_1638);
nor U477 (N_477,In_1808,In_307);
nand U478 (N_478,In_1579,In_752);
and U479 (N_479,N_131,In_1736);
or U480 (N_480,In_2321,In_1135);
and U481 (N_481,In_1704,In_2318);
and U482 (N_482,In_1820,In_626);
or U483 (N_483,In_1362,In_1508);
and U484 (N_484,In_1843,In_1181);
and U485 (N_485,In_143,In_1176);
and U486 (N_486,In_1393,In_874);
and U487 (N_487,In_2205,N_377);
and U488 (N_488,In_836,N_52);
nor U489 (N_489,In_1979,In_1439);
and U490 (N_490,In_1332,In_220);
or U491 (N_491,In_419,In_966);
and U492 (N_492,In_1879,N_398);
and U493 (N_493,In_26,In_1193);
nand U494 (N_494,N_8,N_71);
and U495 (N_495,In_1595,In_1964);
nor U496 (N_496,N_164,In_61);
or U497 (N_497,In_2439,In_1177);
nor U498 (N_498,N_80,In_1441);
or U499 (N_499,N_154,In_489);
and U500 (N_500,In_2419,In_462);
or U501 (N_501,In_1352,In_1340);
nand U502 (N_502,In_2061,In_1858);
or U503 (N_503,In_2311,In_44);
nor U504 (N_504,In_850,In_2310);
and U505 (N_505,In_1433,In_737);
or U506 (N_506,In_2248,In_1784);
nor U507 (N_507,In_2219,In_2415);
nand U508 (N_508,In_1757,In_631);
and U509 (N_509,N_367,In_839);
or U510 (N_510,In_2181,In_2145);
xnor U511 (N_511,In_2394,In_488);
nor U512 (N_512,In_908,In_1463);
or U513 (N_513,In_1072,N_88);
nor U514 (N_514,In_2308,N_226);
nor U515 (N_515,N_183,In_768);
nor U516 (N_516,N_121,In_1137);
or U517 (N_517,In_817,In_629);
xnor U518 (N_518,N_206,In_1796);
nor U519 (N_519,In_1920,In_2144);
nand U520 (N_520,In_1495,In_1309);
nor U521 (N_521,In_1835,In_110);
nand U522 (N_522,In_1341,In_1493);
nor U523 (N_523,N_202,In_1935);
nor U524 (N_524,In_2149,In_2460);
nand U525 (N_525,In_1006,In_2374);
nand U526 (N_526,In_167,In_1563);
nor U527 (N_527,In_1116,N_5);
and U528 (N_528,In_664,In_650);
nor U529 (N_529,N_256,N_331);
nand U530 (N_530,In_563,In_965);
xor U531 (N_531,In_2007,In_835);
and U532 (N_532,In_1103,In_828);
or U533 (N_533,In_2402,N_122);
nor U534 (N_534,In_2067,In_46);
and U535 (N_535,N_91,In_780);
and U536 (N_536,In_1079,In_1401);
or U537 (N_537,In_2467,In_1045);
nand U538 (N_538,In_201,In_734);
or U539 (N_539,In_2024,In_183);
or U540 (N_540,In_1562,N_355);
nand U541 (N_541,In_970,N_228);
or U542 (N_542,In_671,In_442);
or U543 (N_543,In_549,In_428);
nand U544 (N_544,In_240,N_242);
or U545 (N_545,In_341,In_1171);
nand U546 (N_546,In_1084,N_368);
nor U547 (N_547,In_352,In_354);
nor U548 (N_548,In_2237,N_136);
and U549 (N_549,In_1434,In_95);
nand U550 (N_550,In_1099,In_2234);
and U551 (N_551,N_312,In_84);
or U552 (N_552,In_90,N_294);
nor U553 (N_553,In_841,N_266);
nor U554 (N_554,In_2169,In_1007);
nor U555 (N_555,In_1863,In_112);
or U556 (N_556,N_177,In_2326);
nand U557 (N_557,N_109,In_314);
nor U558 (N_558,N_246,In_1180);
and U559 (N_559,N_248,N_345);
or U560 (N_560,In_2250,In_1029);
and U561 (N_561,In_409,In_2211);
nor U562 (N_562,In_2480,In_2155);
nor U563 (N_563,N_74,In_1278);
nor U564 (N_564,In_613,In_2273);
nor U565 (N_565,In_665,N_116);
nor U566 (N_566,In_750,N_218);
and U567 (N_567,In_569,In_924);
or U568 (N_568,In_275,In_27);
or U569 (N_569,In_1655,In_2400);
or U570 (N_570,In_917,In_193);
nand U571 (N_571,In_547,In_80);
or U572 (N_572,In_1242,In_1706);
or U573 (N_573,In_1207,In_2193);
or U574 (N_574,In_30,In_166);
nand U575 (N_575,In_1962,N_238);
nand U576 (N_576,N_252,N_334);
or U577 (N_577,In_2084,In_877);
and U578 (N_578,In_1759,In_2362);
nand U579 (N_579,In_1063,N_341);
nor U580 (N_580,In_399,In_455);
nand U581 (N_581,In_2276,In_1299);
and U582 (N_582,N_103,N_362);
or U583 (N_583,In_632,In_203);
nor U584 (N_584,In_1151,In_776);
and U585 (N_585,In_1696,In_157);
nand U586 (N_586,In_453,In_1010);
nor U587 (N_587,In_2170,In_432);
nor U588 (N_588,In_954,In_851);
or U589 (N_589,N_151,N_64);
nand U590 (N_590,In_1822,In_1327);
and U591 (N_591,In_1787,In_213);
nand U592 (N_592,In_1819,In_958);
nor U593 (N_593,In_2083,In_579);
nand U594 (N_594,In_430,In_2474);
and U595 (N_595,In_658,In_1929);
nor U596 (N_596,In_2257,In_765);
and U597 (N_597,In_1968,In_1182);
or U598 (N_598,In_1276,In_1685);
or U599 (N_599,In_1363,In_1254);
or U600 (N_600,In_1355,In_256);
nor U601 (N_601,In_2387,In_2222);
nand U602 (N_602,N_216,N_143);
nand U603 (N_603,In_1066,In_139);
or U604 (N_604,In_1684,In_401);
nor U605 (N_605,In_1266,In_2120);
xor U606 (N_606,N_414,N_576);
or U607 (N_607,In_1660,In_1402);
nor U608 (N_608,In_888,In_1389);
or U609 (N_609,N_482,In_895);
and U610 (N_610,In_591,N_436);
nand U611 (N_611,In_1980,In_480);
nand U612 (N_612,In_2466,In_2129);
nor U613 (N_613,N_408,In_1937);
or U614 (N_614,In_309,In_443);
nand U615 (N_615,In_1075,In_1284);
or U616 (N_616,In_1219,N_493);
and U617 (N_617,In_517,In_374);
or U618 (N_618,In_997,N_244);
and U619 (N_619,In_1148,In_1110);
nor U620 (N_620,N_292,N_561);
nand U621 (N_621,In_1265,In_305);
or U622 (N_622,In_2397,In_856);
nand U623 (N_623,N_346,N_506);
nor U624 (N_624,In_1046,N_40);
nand U625 (N_625,In_668,N_452);
or U626 (N_626,N_443,In_539);
nand U627 (N_627,In_1196,In_1951);
and U628 (N_628,In_2194,In_556);
or U629 (N_629,In_13,In_697);
nor U630 (N_630,In_2254,In_1582);
nand U631 (N_631,In_499,In_1793);
nand U632 (N_632,In_978,In_1399);
and U633 (N_633,In_673,In_2201);
and U634 (N_634,In_570,N_221);
nor U635 (N_635,N_395,N_545);
nand U636 (N_636,In_2337,In_2331);
and U637 (N_637,In_2278,In_2366);
and U638 (N_638,N_402,In_633);
nor U639 (N_639,N_535,N_579);
or U640 (N_640,In_2316,In_2484);
nor U641 (N_641,In_1248,N_598);
or U642 (N_642,In_1085,In_1695);
nor U643 (N_643,In_722,In_2378);
and U644 (N_644,N_117,In_2020);
and U645 (N_645,In_2465,In_1425);
nor U646 (N_646,In_1342,In_1770);
or U647 (N_647,In_2148,In_1665);
and U648 (N_648,In_37,In_250);
and U649 (N_649,In_675,In_204);
nand U650 (N_650,In_1310,In_1358);
or U651 (N_651,N_278,In_117);
or U652 (N_652,N_550,In_1167);
nor U653 (N_653,In_525,In_2275);
nand U654 (N_654,In_1350,In_2142);
nand U655 (N_655,In_1587,N_342);
or U656 (N_656,In_160,In_228);
nor U657 (N_657,N_37,In_1540);
nor U658 (N_658,In_54,N_192);
or U659 (N_659,N_591,In_1383);
nand U660 (N_660,In_1271,In_2220);
nand U661 (N_661,In_2202,In_152);
nand U662 (N_662,In_2405,In_2229);
and U663 (N_663,In_1522,In_2191);
nand U664 (N_664,In_440,In_1516);
nor U665 (N_665,In_1365,In_1541);
nor U666 (N_666,In_1125,In_2171);
nor U667 (N_667,In_2235,N_470);
or U668 (N_668,In_1239,In_1731);
or U669 (N_669,In_2499,In_2372);
nand U670 (N_670,In_1992,In_1605);
nand U671 (N_671,N_146,N_400);
or U672 (N_672,In_89,In_33);
nand U673 (N_673,In_1489,In_1809);
nand U674 (N_674,In_1905,In_162);
nand U675 (N_675,In_1234,N_245);
nand U676 (N_676,In_1878,N_567);
nor U677 (N_677,In_472,N_453);
and U678 (N_678,In_1316,In_2259);
nand U679 (N_679,N_95,In_448);
or U680 (N_680,In_2364,In_827);
nor U681 (N_681,In_804,In_2054);
or U682 (N_682,In_498,In_2283);
or U683 (N_683,N_434,In_1038);
and U684 (N_684,In_2057,In_1817);
and U685 (N_685,In_2449,N_504);
nor U686 (N_686,In_1157,In_661);
nand U687 (N_687,N_69,In_571);
and U688 (N_688,In_128,In_2463);
nand U689 (N_689,N_212,In_936);
and U690 (N_690,In_2064,In_1624);
or U691 (N_691,N_525,In_2388);
nand U692 (N_692,In_559,In_519);
nor U693 (N_693,In_2432,N_511);
and U694 (N_694,In_2353,In_1417);
nor U695 (N_695,N_176,In_1589);
nor U696 (N_696,In_1458,In_1749);
or U697 (N_697,In_809,N_289);
or U698 (N_698,N_532,N_337);
nand U699 (N_699,In_1438,In_1956);
or U700 (N_700,In_1530,In_273);
nand U701 (N_701,In_690,In_1087);
nand U702 (N_702,In_47,N_73);
nand U703 (N_703,In_2143,In_2416);
nand U704 (N_704,N_445,In_1519);
and U705 (N_705,N_137,In_35);
nand U706 (N_706,In_1564,In_2270);
or U707 (N_707,In_858,In_1499);
nand U708 (N_708,In_1816,In_1580);
or U709 (N_709,In_1014,In_2092);
nand U710 (N_710,N_358,In_1824);
and U711 (N_711,N_344,In_1445);
nand U712 (N_712,In_2329,In_208);
or U713 (N_713,In_1676,In_648);
and U714 (N_714,N_225,In_2166);
or U715 (N_715,In_2330,In_2336);
or U716 (N_716,In_1405,In_1065);
or U717 (N_717,N_321,In_1965);
nand U718 (N_718,In_1901,In_452);
nor U719 (N_719,N_544,In_2110);
nand U720 (N_720,In_34,In_602);
or U721 (N_721,In_407,In_49);
and U722 (N_722,In_1751,In_2106);
and U723 (N_723,N_29,In_2376);
and U724 (N_724,In_1916,N_23);
nor U725 (N_725,N_354,In_215);
nor U726 (N_726,In_727,In_863);
and U727 (N_727,In_481,In_890);
or U728 (N_728,In_605,N_481);
and U729 (N_729,In_1138,In_202);
or U730 (N_730,N_547,In_2281);
and U731 (N_731,In_1351,In_869);
or U732 (N_732,In_940,In_2016);
and U733 (N_733,N_376,In_1555);
nor U734 (N_734,In_2123,N_188);
and U735 (N_735,N_528,In_332);
nand U736 (N_736,In_1742,N_55);
or U737 (N_737,In_2047,In_2284);
nor U738 (N_738,In_1957,In_20);
nor U739 (N_739,In_382,N_410);
and U740 (N_740,N_196,N_518);
or U741 (N_741,N_26,N_81);
nor U742 (N_742,N_205,N_223);
and U743 (N_743,In_2041,N_84);
xor U744 (N_744,In_862,In_1680);
and U745 (N_745,N_399,In_2414);
or U746 (N_746,In_1545,In_302);
nand U747 (N_747,In_1501,In_447);
or U748 (N_748,In_2113,In_2088);
nand U749 (N_749,In_1161,N_370);
or U750 (N_750,In_1377,In_259);
or U751 (N_751,In_794,N_444);
or U752 (N_752,In_1485,In_2469);
or U753 (N_753,In_2244,In_1792);
nand U754 (N_754,In_2053,In_1037);
or U755 (N_755,In_777,In_774);
and U756 (N_756,In_2452,N_465);
nand U757 (N_757,In_2433,In_2208);
nor U758 (N_758,In_2152,N_520);
or U759 (N_759,In_1986,N_293);
nor U760 (N_760,In_1881,N_304);
and U761 (N_761,In_155,In_984);
nand U762 (N_762,In_1390,In_418);
nor U763 (N_763,In_271,In_751);
nor U764 (N_764,In_1270,In_1475);
or U765 (N_765,N_229,N_516);
or U766 (N_766,N_578,In_1651);
nand U767 (N_767,In_585,N_302);
nor U768 (N_768,N_427,In_879);
or U769 (N_769,In_326,In_935);
and U770 (N_770,In_62,In_1746);
or U771 (N_771,In_1216,N_329);
nand U772 (N_772,In_263,In_760);
or U773 (N_773,In_2406,In_1491);
or U774 (N_774,In_1255,In_1768);
and U775 (N_775,In_2172,N_382);
nand U776 (N_776,N_477,In_391);
or U777 (N_777,In_1213,In_1406);
or U778 (N_778,N_573,In_2103);
or U779 (N_779,In_1573,In_2409);
nand U780 (N_780,In_350,In_561);
nand U781 (N_781,In_2411,N_114);
nand U782 (N_782,N_409,N_241);
or U783 (N_783,N_597,N_66);
nand U784 (N_784,In_1105,In_2070);
and U785 (N_785,N_112,In_635);
or U786 (N_786,N_282,In_1978);
or U787 (N_787,In_1273,In_1936);
or U788 (N_788,In_1613,In_1455);
nand U789 (N_789,In_2436,N_17);
nor U790 (N_790,In_278,In_279);
or U791 (N_791,N_194,In_1549);
or U792 (N_792,In_2180,In_1875);
nor U793 (N_793,N_315,N_388);
or U794 (N_794,N_264,N_429);
or U795 (N_795,N_15,In_2346);
nor U796 (N_796,In_823,In_144);
or U797 (N_797,In_1672,In_905);
or U798 (N_798,N_239,In_2354);
nor U799 (N_799,In_564,N_247);
and U800 (N_800,In_2438,In_1570);
or U801 (N_801,In_2307,N_314);
nor U802 (N_802,N_694,N_723);
nand U803 (N_803,In_180,In_2448);
nor U804 (N_804,In_242,In_1502);
nand U805 (N_805,In_1250,N_169);
nand U806 (N_806,N_653,In_1893);
and U807 (N_807,In_730,In_1683);
nand U808 (N_808,In_1652,In_356);
or U809 (N_809,N_458,In_1467);
nand U810 (N_810,N_500,In_1973);
or U811 (N_811,In_127,In_2);
nor U812 (N_812,N_495,In_1884);
nor U813 (N_813,In_729,In_104);
nand U814 (N_814,In_705,N_72);
nor U815 (N_815,In_500,N_700);
or U816 (N_816,In_1724,N_42);
nor U817 (N_817,In_1440,In_688);
or U818 (N_818,In_435,N_335);
and U819 (N_819,In_1034,In_1162);
and U820 (N_820,N_227,N_413);
nand U821 (N_821,In_1301,In_2203);
or U822 (N_822,In_2072,In_501);
nand U823 (N_823,In_1811,N_75);
or U824 (N_824,In_1853,In_196);
nor U825 (N_825,N_36,In_2076);
nor U826 (N_826,In_700,In_1551);
and U827 (N_827,In_1150,In_2358);
nand U828 (N_828,In_1807,In_2186);
nor U829 (N_829,N_719,In_598);
nor U830 (N_830,N_585,N_449);
nand U831 (N_831,N_46,In_188);
nor U832 (N_832,In_2027,In_2111);
or U833 (N_833,In_1852,In_83);
or U834 (N_834,N_474,In_1114);
xnor U835 (N_835,In_914,In_1535);
and U836 (N_836,N_526,In_1583);
nor U837 (N_837,N_417,In_2292);
nand U838 (N_838,In_14,In_627);
nand U839 (N_839,In_2243,In_949);
nand U840 (N_840,N_601,In_948);
nor U841 (N_841,In_320,In_581);
xor U842 (N_842,In_1132,In_789);
or U843 (N_843,In_281,In_813);
nor U844 (N_844,N_451,N_697);
and U845 (N_845,N_745,In_446);
nor U846 (N_846,In_2134,In_1267);
nand U847 (N_847,In_1703,N_274);
and U848 (N_848,In_710,N_552);
and U849 (N_849,In_1782,N_648);
and U850 (N_850,In_2288,In_1262);
nor U851 (N_851,In_510,N_799);
nor U852 (N_852,N_157,N_351);
or U853 (N_853,In_2328,N_566);
nor U854 (N_854,N_654,N_610);
nor U855 (N_855,In_53,N_447);
nor U856 (N_856,N_717,N_390);
and U857 (N_857,N_698,In_1778);
or U858 (N_858,N_153,In_1618);
or U859 (N_859,In_2361,In_802);
nor U860 (N_860,N_666,In_134);
and U861 (N_861,In_1381,In_712);
or U862 (N_862,In_1996,N_372);
and U863 (N_863,In_1281,In_1781);
or U864 (N_864,In_412,N_633);
nor U865 (N_865,N_462,In_254);
or U866 (N_866,In_1831,In_1215);
nand U867 (N_867,In_2107,In_2434);
and U868 (N_868,In_1866,In_150);
or U869 (N_869,In_1172,N_180);
or U870 (N_870,In_820,In_1773);
nand U871 (N_871,In_687,In_870);
and U872 (N_872,N_213,N_673);
or U873 (N_873,In_660,N_480);
nand U874 (N_874,N_207,N_557);
nand U875 (N_875,In_1654,In_1293);
and U876 (N_876,In_2293,N_626);
nor U877 (N_877,In_757,N_336);
nand U878 (N_878,In_713,In_22);
or U879 (N_879,In_369,In_2232);
nand U880 (N_880,N_538,N_527);
nand U881 (N_881,In_693,In_1447);
nand U882 (N_882,In_515,In_1546);
nand U883 (N_883,In_805,In_2011);
nand U884 (N_884,In_303,In_709);
or U885 (N_885,In_1715,N_237);
nand U886 (N_886,N_599,N_539);
or U887 (N_887,In_207,In_1677);
or U888 (N_888,In_1723,N_796);
and U889 (N_889,In_1578,In_1908);
and U890 (N_890,In_1584,In_107);
and U891 (N_891,In_1698,N_0);
or U892 (N_892,N_668,In_1509);
and U893 (N_893,In_1656,In_2045);
nand U894 (N_894,In_2233,In_422);
xor U895 (N_895,N_419,In_509);
nor U896 (N_896,N_99,N_30);
nor U897 (N_897,In_1719,In_42);
or U898 (N_898,In_479,In_1726);
or U899 (N_899,In_1107,In_646);
nor U900 (N_900,N_787,N_230);
and U901 (N_901,N_328,In_1880);
nand U902 (N_902,In_324,N_772);
and U903 (N_903,In_1113,In_1963);
nand U904 (N_904,N_514,N_373);
nor U905 (N_905,N_508,N_200);
xor U906 (N_906,In_1975,In_2039);
nand U907 (N_907,In_2048,In_1825);
nand U908 (N_908,N_13,In_2002);
or U909 (N_909,In_1518,In_2475);
and U910 (N_910,In_1028,In_625);
or U911 (N_911,In_1889,In_1838);
nand U912 (N_912,In_1374,N_473);
nor U913 (N_913,N_716,N_318);
nor U914 (N_914,In_913,In_1035);
nand U915 (N_915,In_1031,In_2301);
and U916 (N_916,In_683,In_849);
or U917 (N_917,N_298,N_686);
nand U918 (N_918,In_864,N_701);
nand U919 (N_919,In_192,N_469);
or U920 (N_920,N_138,N_178);
nand U921 (N_921,In_906,N_624);
or U922 (N_922,In_2207,In_1446);
nand U923 (N_923,In_719,N_14);
nor U924 (N_924,N_760,In_65);
and U925 (N_925,In_32,In_2200);
nand U926 (N_926,N_352,In_492);
nor U927 (N_927,In_715,N_714);
nor U928 (N_928,In_2019,In_2444);
or U929 (N_929,N_448,In_124);
nand U930 (N_930,In_1044,In_2246);
and U931 (N_931,N_466,In_930);
or U932 (N_932,N_691,In_1415);
or U933 (N_933,In_1627,N_65);
nor U934 (N_934,In_2403,In_1152);
nor U935 (N_935,N_795,In_1464);
or U936 (N_936,N_676,N_365);
nand U937 (N_937,In_476,N_590);
nand U938 (N_938,N_709,In_1803);
or U939 (N_939,N_450,In_1990);
nand U940 (N_940,In_706,In_478);
or U941 (N_941,In_1212,N_534);
nand U942 (N_942,In_1885,In_387);
or U943 (N_943,In_1407,N_478);
nand U944 (N_944,N_727,In_2431);
and U945 (N_945,N_732,In_2261);
and U946 (N_946,In_1640,In_672);
nor U947 (N_947,N_530,In_2095);
nand U948 (N_948,In_728,In_258);
and U949 (N_949,In_912,In_2343);
or U950 (N_950,In_251,In_2091);
nor U951 (N_951,N_607,In_436);
or U952 (N_952,In_1345,In_102);
and U953 (N_953,In_1183,N_327);
nor U954 (N_954,N_637,In_1777);
nand U955 (N_955,N_253,N_670);
nor U956 (N_956,In_2014,In_893);
and U957 (N_957,In_122,In_2381);
nand U958 (N_958,In_469,N_9);
or U959 (N_959,In_2230,In_113);
nor U960 (N_960,In_532,In_1842);
or U961 (N_961,In_2424,In_919);
and U962 (N_962,In_214,N_476);
or U963 (N_963,In_1122,In_12);
or U964 (N_964,In_260,In_458);
or U965 (N_965,N_262,In_2485);
nand U966 (N_966,N_142,In_2391);
nand U967 (N_967,N_641,In_1353);
nand U968 (N_968,In_1877,N_739);
or U969 (N_969,In_449,In_654);
and U970 (N_970,In_1366,In_467);
and U971 (N_971,In_2459,In_2442);
or U972 (N_972,N_757,N_515);
nand U973 (N_973,N_285,N_297);
nor U974 (N_974,In_190,In_1581);
nand U975 (N_975,In_883,In_138);
or U976 (N_976,In_1430,N_163);
or U977 (N_977,N_678,N_394);
and U978 (N_978,N_371,In_558);
and U979 (N_979,N_788,N_777);
or U980 (N_980,In_831,In_1641);
nand U981 (N_981,In_546,N_770);
and U982 (N_982,N_517,In_1865);
or U983 (N_983,In_473,In_1178);
nor U984 (N_984,In_1120,N_735);
and U985 (N_985,In_417,In_2385);
or U986 (N_986,N_185,In_1457);
and U987 (N_987,N_265,N_589);
or U988 (N_988,In_410,In_1052);
and U989 (N_989,In_145,In_1818);
and U990 (N_990,In_2158,In_1610);
nor U991 (N_991,In_246,N_662);
and U992 (N_992,In_2121,In_565);
or U993 (N_993,In_1163,In_1357);
nand U994 (N_994,N_193,In_786);
xor U995 (N_995,In_262,In_1024);
nand U996 (N_996,In_1946,In_541);
nand U997 (N_997,In_2136,N_496);
or U998 (N_998,In_2038,In_289);
and U999 (N_999,In_837,In_1222);
or U1000 (N_1000,In_848,In_973);
and U1001 (N_1001,N_272,In_2141);
and U1002 (N_1002,N_971,N_741);
and U1003 (N_1003,In_996,In_225);
nor U1004 (N_1004,N_197,In_1098);
or U1005 (N_1005,In_1611,In_1836);
nor U1006 (N_1006,N_35,N_261);
or U1007 (N_1007,In_450,N_860);
and U1008 (N_1008,N_674,In_505);
or U1009 (N_1009,In_1372,N_862);
and U1010 (N_1010,N_280,N_537);
nor U1011 (N_1011,In_221,N_785);
and U1012 (N_1012,In_724,N_190);
nand U1013 (N_1013,In_319,In_2239);
and U1014 (N_1014,N_375,In_464);
xnor U1015 (N_1015,In_1127,N_858);
nand U1016 (N_1016,In_129,In_1662);
and U1017 (N_1017,N_222,In_244);
nand U1018 (N_1018,In_2137,In_826);
or U1019 (N_1019,In_1247,N_671);
and U1020 (N_1020,In_1902,N_89);
nor U1021 (N_1021,In_1397,In_2082);
nor U1022 (N_1022,In_528,In_2447);
nor U1023 (N_1023,In_2365,In_2074);
nand U1024 (N_1024,In_2289,In_1713);
and U1025 (N_1025,In_1314,N_140);
and U1026 (N_1026,In_1851,In_1175);
nand U1027 (N_1027,N_366,In_292);
and U1028 (N_1028,N_96,N_595);
and U1029 (N_1029,N_379,In_892);
nor U1030 (N_1030,N_505,N_503);
or U1031 (N_1031,N_295,N_584);
or U1032 (N_1032,N_659,N_809);
nor U1033 (N_1033,In_72,In_2351);
nand U1034 (N_1034,In_168,N_774);
or U1035 (N_1035,N_316,In_1246);
nand U1036 (N_1036,In_522,In_681);
nand U1037 (N_1037,N_353,In_797);
nor U1038 (N_1038,N_864,N_905);
nor U1039 (N_1039,In_1767,In_1056);
or U1040 (N_1040,N_681,N_913);
or U1041 (N_1041,In_725,In_1547);
and U1042 (N_1042,In_1542,In_1251);
or U1043 (N_1043,N_827,In_2269);
nor U1044 (N_1044,In_2052,N_7);
and U1045 (N_1045,N_819,N_300);
and U1046 (N_1046,In_669,In_1220);
nand U1047 (N_1047,In_368,In_1003);
nor U1048 (N_1048,N_554,N_20);
and U1049 (N_1049,In_939,N_521);
or U1050 (N_1050,N_914,In_291);
nand U1051 (N_1051,In_2258,N_179);
and U1052 (N_1052,In_1173,In_2036);
or U1053 (N_1053,N_997,N_890);
and U1054 (N_1054,In_392,In_1557);
and U1055 (N_1055,In_2080,In_1832);
and U1056 (N_1056,In_1629,In_1805);
or U1057 (N_1057,In_1042,In_1040);
nor U1058 (N_1058,N_78,N_941);
and U1059 (N_1059,N_428,N_612);
and U1060 (N_1060,In_1783,N_921);
and U1061 (N_1061,N_559,N_911);
or U1062 (N_1062,In_1369,N_992);
nor U1063 (N_1063,N_338,In_1507);
or U1064 (N_1064,In_2338,N_811);
nand U1065 (N_1065,In_198,N_571);
and U1066 (N_1066,N_254,N_423);
nor U1067 (N_1067,In_819,N_243);
xnor U1068 (N_1068,In_2065,In_99);
and U1069 (N_1069,In_133,N_446);
nand U1070 (N_1070,In_103,In_2022);
nor U1071 (N_1071,In_245,N_768);
nand U1072 (N_1072,In_2282,N_76);
and U1073 (N_1073,N_118,In_330);
and U1074 (N_1074,N_543,In_953);
nand U1075 (N_1075,N_978,In_2304);
or U1076 (N_1076,N_821,N_588);
or U1077 (N_1077,In_1077,In_1675);
or U1078 (N_1078,In_1285,N_215);
nor U1079 (N_1079,In_1911,N_460);
or U1080 (N_1080,In_1712,N_931);
nand U1081 (N_1081,N_652,N_541);
nor U1082 (N_1082,N_290,N_989);
nand U1083 (N_1083,N_724,N_467);
nor U1084 (N_1084,N_565,In_1295);
nand U1085 (N_1085,N_431,In_2099);
nand U1086 (N_1086,In_227,N_263);
nand U1087 (N_1087,In_361,In_1229);
nand U1088 (N_1088,In_1586,In_2272);
and U1089 (N_1089,In_1349,N_948);
nor U1090 (N_1090,N_269,In_353);
nand U1091 (N_1091,In_1134,N_791);
or U1092 (N_1092,N_270,In_645);
nand U1093 (N_1093,In_689,In_801);
nand U1094 (N_1094,In_1839,In_2482);
and U1095 (N_1095,N_743,N_617);
and U1096 (N_1096,In_1011,N_549);
nand U1097 (N_1097,N_214,N_814);
nor U1098 (N_1098,N_58,N_929);
nand U1099 (N_1099,In_2157,N_523);
nor U1100 (N_1100,N_930,In_1667);
nand U1101 (N_1101,N_792,N_171);
nand U1102 (N_1102,N_484,In_2477);
and U1103 (N_1103,In_50,N_77);
or U1104 (N_1104,N_425,In_812);
or U1105 (N_1105,In_2399,In_641);
and U1106 (N_1106,N_816,In_2236);
nor U1107 (N_1107,N_483,N_203);
or U1108 (N_1108,In_1473,N_640);
nand U1109 (N_1109,N_490,In_404);
and U1110 (N_1110,In_1959,N_440);
and U1111 (N_1111,In_617,In_682);
nand U1112 (N_1112,In_859,N_546);
nor U1113 (N_1113,In_1939,N_846);
or U1114 (N_1114,In_2185,In_608);
nand U1115 (N_1115,In_916,N_385);
or U1116 (N_1116,In_378,In_1989);
and U1117 (N_1117,N_249,N_357);
and U1118 (N_1118,N_897,In_165);
or U1119 (N_1119,In_1725,In_2216);
nand U1120 (N_1120,N_679,In_2417);
or U1121 (N_1121,In_2037,In_560);
or U1122 (N_1122,N_966,In_825);
nor U1123 (N_1123,In_31,N_977);
or U1124 (N_1124,In_156,N_710);
nor U1125 (N_1125,In_2190,In_749);
nor U1126 (N_1126,N_533,In_1659);
nor U1127 (N_1127,In_830,In_2046);
and U1128 (N_1128,N_441,N_79);
nand U1129 (N_1129,In_1681,In_747);
nand U1130 (N_1130,In_1420,In_178);
or U1131 (N_1131,N_857,N_522);
nor U1132 (N_1132,N_350,In_1466);
and U1133 (N_1133,N_904,In_2490);
nor U1134 (N_1134,In_513,N_259);
nand U1135 (N_1135,In_1051,N_845);
nor U1136 (N_1136,In_999,In_536);
and U1137 (N_1137,In_224,In_318);
or U1138 (N_1138,N_407,N_492);
and U1139 (N_1139,N_824,In_70);
nand U1140 (N_1140,In_2118,In_1380);
and U1141 (N_1141,In_937,N_753);
or U1142 (N_1142,In_2393,In_1829);
nor U1143 (N_1143,N_893,N_658);
xnor U1144 (N_1144,In_2059,N_487);
nand U1145 (N_1145,In_1806,N_435);
nor U1146 (N_1146,N_629,N_850);
and U1147 (N_1147,In_335,N_471);
and U1148 (N_1148,In_2356,In_1649);
nand U1149 (N_1149,In_39,In_871);
nor U1150 (N_1150,In_11,N_442);
and U1151 (N_1151,N_608,In_2306);
or U1152 (N_1152,N_863,In_1291);
nand U1153 (N_1153,N_832,In_1230);
and U1154 (N_1154,In_1431,N_749);
and U1155 (N_1155,N_947,N_938);
or U1156 (N_1156,N_455,N_489);
nor U1157 (N_1157,In_540,N_656);
nor U1158 (N_1158,In_1862,In_692);
nor U1159 (N_1159,In_790,In_337);
and U1160 (N_1160,N_936,In_397);
or U1161 (N_1161,N_778,In_2177);
and U1162 (N_1162,In_1876,In_1376);
or U1163 (N_1163,In_529,In_818);
nand U1164 (N_1164,In_1534,In_2102);
or U1165 (N_1165,In_1812,In_2297);
nor U1166 (N_1166,In_1256,N_106);
nand U1167 (N_1167,N_524,In_910);
nor U1168 (N_1168,In_1311,In_659);
nand U1169 (N_1169,In_1149,N_479);
nor U1170 (N_1170,In_931,N_220);
nor U1171 (N_1171,N_271,In_1048);
nand U1172 (N_1172,In_1909,In_439);
nand U1173 (N_1173,N_767,In_1592);
nand U1174 (N_1174,In_351,In_1790);
nand U1175 (N_1175,N_619,N_783);
and U1176 (N_1176,In_1632,N_10);
or U1177 (N_1177,In_1527,In_357);
nand U1178 (N_1178,In_553,In_67);
or U1179 (N_1179,N_880,In_1454);
or U1180 (N_1180,N_150,N_882);
nand U1181 (N_1181,In_424,In_1209);
or U1182 (N_1182,In_1554,In_2055);
and U1183 (N_1183,N_191,In_2446);
nand U1184 (N_1184,N_628,In_331);
or U1185 (N_1185,N_405,In_972);
or U1186 (N_1186,In_1607,N_990);
nand U1187 (N_1187,In_367,N_884);
or U1188 (N_1188,N_582,N_885);
nor U1189 (N_1189,N_403,N_49);
and U1190 (N_1190,In_1154,N_141);
nand U1191 (N_1191,N_631,In_223);
and U1192 (N_1192,N_708,N_291);
and U1193 (N_1193,N_830,N_606);
nor U1194 (N_1194,N_16,In_656);
or U1195 (N_1195,N_915,N_615);
or U1196 (N_1196,In_587,In_1021);
nand U1197 (N_1197,N_564,In_1648);
or U1198 (N_1198,N_306,In_59);
and U1199 (N_1199,In_2056,N_472);
xnor U1200 (N_1200,In_1005,In_2128);
or U1201 (N_1201,In_1086,N_67);
and U1202 (N_1202,N_332,N_1029);
or U1203 (N_1203,N_392,N_94);
nand U1204 (N_1204,N_683,N_1152);
nor U1205 (N_1205,In_853,N_1178);
or U1206 (N_1206,N_260,In_967);
and U1207 (N_1207,N_883,In_1093);
nor U1208 (N_1208,In_1403,In_784);
nand U1209 (N_1209,N_750,In_1553);
and U1210 (N_1210,In_1269,In_2312);
nor U1211 (N_1211,N_286,N_1036);
nand U1212 (N_1212,N_211,N_1065);
and U1213 (N_1213,N_841,N_438);
nor U1214 (N_1214,In_847,In_1049);
and U1215 (N_1215,In_2487,N_896);
nand U1216 (N_1216,In_814,N_208);
and U1217 (N_1217,N_964,N_1033);
and U1218 (N_1218,In_1282,In_1864);
or U1219 (N_1219,N_1025,N_926);
and U1220 (N_1220,N_889,N_794);
and U1221 (N_1221,In_1828,In_1571);
nand U1222 (N_1222,In_788,N_1128);
and U1223 (N_1223,In_1619,In_2161);
nor U1224 (N_1224,N_1096,N_693);
or U1225 (N_1225,In_1701,In_235);
or U1226 (N_1226,In_2294,In_366);
and U1227 (N_1227,N_1172,N_1177);
nand U1228 (N_1228,In_170,N_754);
nand U1229 (N_1229,N_1105,N_958);
nor U1230 (N_1230,In_1396,N_820);
and U1231 (N_1231,N_963,N_422);
nor U1232 (N_1232,In_186,N_313);
or U1233 (N_1233,N_1008,In_1707);
or U1234 (N_1234,In_1511,In_322);
nor U1235 (N_1235,In_1023,N_643);
nand U1236 (N_1236,In_703,N_720);
or U1237 (N_1237,In_2115,N_935);
nor U1238 (N_1238,N_1141,N_925);
or U1239 (N_1239,In_1932,In_1283);
or U1240 (N_1240,N_1089,N_497);
nand U1241 (N_1241,In_1492,N_634);
or U1242 (N_1242,In_175,N_1085);
or U1243 (N_1243,N_1088,In_1594);
xnor U1244 (N_1244,In_1436,N_861);
or U1245 (N_1245,N_1199,N_1050);
nor U1246 (N_1246,In_1558,N_333);
nand U1247 (N_1247,In_86,In_2032);
or U1248 (N_1248,N_764,In_2352);
nor U1249 (N_1249,N_962,N_622);
or U1250 (N_1250,N_995,In_717);
or U1251 (N_1251,In_2359,In_2199);
and U1252 (N_1252,N_1045,N_919);
and U1253 (N_1253,In_1476,N_50);
and U1254 (N_1254,In_2226,In_1474);
nand U1255 (N_1255,In_1690,In_643);
nor U1256 (N_1256,N_736,N_695);
and U1257 (N_1257,N_113,N_1149);
and U1258 (N_1258,In_132,In_1354);
nor U1259 (N_1259,N_878,In_1827);
and U1260 (N_1260,In_575,In_584);
and U1261 (N_1261,In_1328,N_976);
and U1262 (N_1262,In_339,In_686);
or U1263 (N_1263,In_2021,N_115);
and U1264 (N_1264,In_901,In_968);
nor U1265 (N_1265,In_932,In_852);
or U1266 (N_1266,In_1453,N_660);
and U1267 (N_1267,N_856,N_464);
or U1268 (N_1268,In_1200,N_742);
and U1269 (N_1269,N_721,N_551);
or U1270 (N_1270,N_982,In_929);
or U1271 (N_1271,In_1560,N_1067);
and U1272 (N_1272,N_991,N_85);
nor U1273 (N_1273,In_2295,In_2075);
and U1274 (N_1274,N_927,In_1206);
or U1275 (N_1275,N_804,N_604);
and U1276 (N_1276,N_1161,In_1650);
nor U1277 (N_1277,N_972,N_1038);
nor U1278 (N_1278,In_946,N_1119);
nand U1279 (N_1279,N_689,N_960);
nor U1280 (N_1280,N_303,In_1974);
nor U1281 (N_1281,N_301,In_470);
nor U1282 (N_1282,N_1188,In_137);
and U1283 (N_1283,In_2150,N_815);
and U1284 (N_1284,N_130,In_1556);
or U1285 (N_1285,In_477,N_747);
and U1286 (N_1286,N_430,In_990);
or U1287 (N_1287,In_1324,N_800);
nor U1288 (N_1288,N_90,In_2068);
and U1289 (N_1289,In_2445,In_1470);
or U1290 (N_1290,In_942,N_954);
nor U1291 (N_1291,N_1126,N_340);
nor U1292 (N_1292,N_718,In_28);
and U1293 (N_1293,In_2398,In_2114);
nor U1294 (N_1294,In_885,N_848);
nor U1295 (N_1295,N_956,N_912);
nand U1296 (N_1296,N_713,In_740);
and U1297 (N_1297,N_391,In_1073);
nand U1298 (N_1298,In_2140,N_1080);
or U1299 (N_1299,In_2215,In_338);
and U1300 (N_1300,N_319,N_1003);
nand U1301 (N_1301,In_1735,In_1823);
nor U1302 (N_1302,In_1797,N_840);
or U1303 (N_1303,In_2071,In_153);
and U1304 (N_1304,In_1833,N_1097);
and U1305 (N_1305,N_343,N_822);
nand U1306 (N_1306,N_174,N_1173);
or U1307 (N_1307,In_1306,N_437);
and U1308 (N_1308,In_815,In_336);
or U1309 (N_1309,N_1022,N_25);
nand U1310 (N_1310,In_311,In_1721);
nor U1311 (N_1311,N_53,In_2309);
nand U1312 (N_1312,In_2430,In_923);
or U1313 (N_1313,In_601,In_315);
or U1314 (N_1314,N_1118,In_838);
nand U1315 (N_1315,N_548,N_39);
nor U1316 (N_1316,In_2029,N_933);
nand U1317 (N_1317,In_1413,N_969);
nor U1318 (N_1318,N_910,In_2451);
or U1319 (N_1319,N_835,N_1021);
and U1320 (N_1320,N_491,In_2461);
and U1321 (N_1321,N_195,In_1082);
and U1322 (N_1322,N_1001,N_849);
nor U1323 (N_1323,N_1018,In_811);
and U1324 (N_1324,In_1890,N_513);
and U1325 (N_1325,In_1760,In_1525);
nand U1326 (N_1326,N_851,N_623);
nor U1327 (N_1327,N_219,In_85);
nand U1328 (N_1328,N_672,N_762);
or U1329 (N_1329,N_1084,In_998);
or U1330 (N_1330,In_2116,N_771);
nand U1331 (N_1331,In_595,In_597);
nand U1332 (N_1332,N_711,N_684);
and U1333 (N_1333,N_83,N_1047);
and U1334 (N_1334,N_1049,In_983);
and U1335 (N_1335,N_877,N_773);
and U1336 (N_1336,N_870,In_943);
nor U1337 (N_1337,N_793,N_187);
and U1338 (N_1338,In_531,In_1185);
and U1339 (N_1339,N_1012,N_876);
xor U1340 (N_1340,N_54,In_1593);
nor U1341 (N_1341,In_1410,In_219);
nand U1342 (N_1342,In_1039,N_955);
nor U1343 (N_1343,N_1010,N_1171);
nor U1344 (N_1344,In_766,In_2324);
nand U1345 (N_1345,N_605,In_51);
or U1346 (N_1346,N_255,In_48);
and U1347 (N_1347,N_602,In_2147);
nor U1348 (N_1348,In_2227,N_507);
and U1349 (N_1349,In_1981,N_498);
nand U1350 (N_1350,N_1190,N_837);
and U1351 (N_1351,N_609,In_507);
nand U1352 (N_1352,In_854,N_330);
and U1353 (N_1353,N_1051,In_1504);
nand U1354 (N_1354,N_984,N_1125);
nor U1355 (N_1355,N_690,N_581);
xnor U1356 (N_1356,N_572,N_32);
nor U1357 (N_1357,In_1515,N_1023);
nor U1358 (N_1358,N_940,N_3);
nand U1359 (N_1359,N_236,In_979);
or U1360 (N_1360,In_993,N_784);
nor U1361 (N_1361,In_293,N_139);
nand U1362 (N_1362,N_866,In_1914);
and U1363 (N_1363,N_855,In_280);
and U1364 (N_1364,N_1048,N_1019);
nor U1365 (N_1365,N_1066,In_372);
or U1366 (N_1366,In_1673,In_527);
and U1367 (N_1367,N_411,In_653);
nor U1368 (N_1368,In_822,N_983);
or U1369 (N_1369,N_61,In_662);
nor U1370 (N_1370,In_1517,In_670);
or U1371 (N_1371,N_133,In_704);
nor U1372 (N_1372,In_537,In_2096);
or U1373 (N_1373,N_275,In_346);
or U1374 (N_1374,In_2028,N_874);
nand U1375 (N_1375,In_568,N_744);
or U1376 (N_1376,N_600,In_1972);
nor U1377 (N_1377,In_1026,In_798);
nand U1378 (N_1378,In_2197,In_753);
and U1379 (N_1379,N_175,In_732);
nor U1380 (N_1380,In_1900,N_558);
or U1381 (N_1381,N_209,N_486);
nor U1382 (N_1382,N_951,In_164);
and U1383 (N_1383,N_722,N_1176);
nor U1384 (N_1384,N_728,In_461);
or U1385 (N_1385,N_798,N_844);
nor U1386 (N_1386,In_1388,N_393);
or U1387 (N_1387,In_1174,In_1303);
nor U1388 (N_1388,In_2089,In_904);
nand U1389 (N_1389,N_1044,N_993);
or U1390 (N_1390,N_937,In_2489);
and U1391 (N_1391,In_1671,N_568);
nand U1392 (N_1392,In_2034,N_1020);
nand U1393 (N_1393,N_1132,N_943);
and U1394 (N_1394,In_19,N_1034);
nand U1395 (N_1395,N_1043,N_779);
and U1396 (N_1396,In_1166,N_692);
nor U1397 (N_1397,N_325,N_1150);
nor U1398 (N_1398,In_880,In_1320);
or U1399 (N_1399,In_959,N_920);
nor U1400 (N_1400,In_1568,N_529);
and U1401 (N_1401,N_810,N_730);
nand U1402 (N_1402,N_574,N_1269);
nor U1403 (N_1403,In_2339,In_74);
nand U1404 (N_1404,In_899,In_1360);
nor U1405 (N_1405,In_1169,In_1198);
nand U1406 (N_1406,In_485,N_1129);
and U1407 (N_1407,N_1325,N_1081);
nand U1408 (N_1408,N_1277,N_201);
and U1409 (N_1409,N_387,In_1304);
nor U1410 (N_1410,In_1421,In_572);
nand U1411 (N_1411,N_1379,N_1207);
nand U1412 (N_1412,N_847,N_1356);
nand U1413 (N_1413,In_2023,N_1298);
nand U1414 (N_1414,In_1057,In_1143);
or U1415 (N_1415,N_1288,In_1694);
nand U1416 (N_1416,N_1253,In_94);
nor U1417 (N_1417,N_1328,N_1095);
nor U1418 (N_1418,In_261,In_1700);
nor U1419 (N_1419,N_1373,In_938);
or U1420 (N_1420,In_1062,In_384);
nand U1421 (N_1421,N_781,In_1347);
or U1422 (N_1422,In_16,In_140);
or U1423 (N_1423,N_592,N_1071);
and U1424 (N_1424,In_1419,N_45);
nor U1425 (N_1425,N_801,N_1341);
nor U1426 (N_1426,N_1109,In_1);
nand U1427 (N_1427,N_424,In_1274);
nand U1428 (N_1428,In_141,N_1323);
or U1429 (N_1429,In_106,N_33);
or U1430 (N_1430,In_1231,N_928);
nor U1431 (N_1431,N_279,N_868);
or U1432 (N_1432,N_1005,N_1344);
nand U1433 (N_1433,In_200,N_267);
nand U1434 (N_1434,N_1294,In_2298);
nand U1435 (N_1435,In_1538,N_1165);
nor U1436 (N_1436,N_776,In_1922);
nand U1437 (N_1437,In_1313,In_2015);
or U1438 (N_1438,N_618,In_2154);
or U1439 (N_1439,N_1395,N_1114);
and U1440 (N_1440,In_299,In_876);
nor U1441 (N_1441,In_1275,In_1128);
or U1442 (N_1442,N_1120,N_512);
nor U1443 (N_1443,N_186,N_233);
and U1444 (N_1444,In_981,N_433);
nand U1445 (N_1445,N_702,N_611);
or U1446 (N_1446,In_1837,In_2423);
or U1447 (N_1447,In_343,N_461);
nor U1448 (N_1448,N_872,N_831);
nor U1449 (N_1449,N_1307,N_1060);
or U1450 (N_1450,In_2256,In_1325);
nand U1451 (N_1451,N_1310,In_2426);
or U1452 (N_1452,In_101,In_1840);
and U1453 (N_1453,In_657,In_866);
nand U1454 (N_1454,In_2179,N_587);
and U1455 (N_1455,In_1095,In_176);
nand U1456 (N_1456,N_105,N_57);
or U1457 (N_1457,In_909,In_371);
nor U1458 (N_1458,In_1359,N_726);
and U1459 (N_1459,N_1371,N_287);
or U1460 (N_1460,N_1224,In_1188);
nand U1461 (N_1461,In_400,In_1903);
or U1462 (N_1462,In_252,N_1316);
nand U1463 (N_1463,N_1345,In_1536);
and U1464 (N_1464,N_1321,In_1631);
nand U1465 (N_1465,In_426,N_1350);
and U1466 (N_1466,In_1577,N_705);
nor U1467 (N_1467,N_1197,In_1272);
or U1468 (N_1468,N_1092,N_120);
or U1469 (N_1469,In_1140,N_594);
nand U1470 (N_1470,In_2425,N_1013);
nand U1471 (N_1471,In_1524,N_1210);
xnor U1472 (N_1472,In_195,N_737);
nor U1473 (N_1473,In_1931,N_994);
nand U1474 (N_1474,In_415,N_1247);
and U1475 (N_1475,In_6,In_1348);
nor U1476 (N_1476,In_163,In_347);
and U1477 (N_1477,N_1332,In_1623);
or U1478 (N_1478,N_1107,N_1216);
nand U1479 (N_1479,In_1218,N_1343);
or U1480 (N_1480,N_906,N_1157);
nor U1481 (N_1481,N_1367,In_2260);
and U1482 (N_1482,N_1239,In_2006);
and U1483 (N_1483,In_1894,In_1983);
or U1484 (N_1484,In_845,In_1609);
nor U1485 (N_1485,In_2437,N_135);
or U1486 (N_1486,N_324,N_765);
nand U1487 (N_1487,In_2001,N_128);
nand U1488 (N_1488,In_1091,N_1103);
nor U1489 (N_1489,In_1416,N_420);
nor U1490 (N_1490,In_1533,In_310);
nand U1491 (N_1491,In_1752,In_746);
nand U1492 (N_1492,In_148,In_149);
nor U1493 (N_1493,In_1237,N_12);
or U1494 (N_1494,In_2221,N_1189);
nand U1495 (N_1495,In_118,N_968);
nor U1496 (N_1496,N_903,In_792);
and U1497 (N_1497,In_1071,In_2370);
nor U1498 (N_1498,N_900,In_2357);
nand U1499 (N_1499,N_852,In_1384);
nand U1500 (N_1500,N_1218,N_1070);
nand U1501 (N_1501,In_2395,N_908);
xnor U1502 (N_1502,N_145,N_1226);
nand U1503 (N_1503,In_2347,In_1326);
or U1504 (N_1504,N_828,N_593);
and U1505 (N_1505,In_782,N_853);
nand U1506 (N_1506,N_1093,In_2224);
or U1507 (N_1507,N_1381,In_1520);
nand U1508 (N_1508,N_1100,N_975);
nand U1509 (N_1509,N_1258,N_1232);
and U1510 (N_1510,In_614,N_1311);
nor U1511 (N_1511,N_1063,N_677);
nor U1512 (N_1512,N_184,In_0);
nand U1513 (N_1513,N_1254,N_542);
and U1514 (N_1514,N_682,In_1450);
nand U1515 (N_1515,N_669,In_345);
nand U1516 (N_1516,N_1348,In_1691);
nand U1517 (N_1517,In_402,In_226);
and U1518 (N_1518,In_41,N_1208);
or U1519 (N_1519,N_1077,In_1141);
and U1520 (N_1520,N_1282,N_310);
nor U1521 (N_1521,In_987,In_969);
or U1522 (N_1522,In_1830,N_182);
nor U1523 (N_1523,N_1182,N_635);
and U1524 (N_1524,N_1156,N_829);
and U1525 (N_1525,N_1369,N_1153);
or U1526 (N_1526,N_945,N_510);
or U1527 (N_1527,In_964,In_1622);
or U1528 (N_1528,N_1243,N_1397);
or U1529 (N_1529,In_878,N_946);
and U1530 (N_1530,In_2060,N_1074);
and U1531 (N_1531,In_619,In_1674);
nor U1532 (N_1532,In_2030,N_494);
and U1533 (N_1533,In_586,N_1192);
xnor U1534 (N_1534,N_1259,N_258);
or U1535 (N_1535,N_1180,In_1523);
and U1536 (N_1536,N_1275,N_1073);
nand U1537 (N_1537,In_1264,N_959);
nor U1538 (N_1538,In_1317,In_2175);
nand U1539 (N_1539,In_772,N_43);
and U1540 (N_1540,In_177,N_1388);
or U1541 (N_1541,N_934,N_1279);
or U1542 (N_1542,N_899,N_257);
xnor U1543 (N_1543,N_887,N_1135);
nor U1544 (N_1544,N_1322,In_1846);
and U1545 (N_1545,In_1214,N_1370);
nand U1546 (N_1546,In_2429,N_894);
or U1547 (N_1547,N_454,N_1290);
or U1548 (N_1548,N_97,In_131);
and U1549 (N_1549,In_1184,N_1193);
and U1550 (N_1550,N_942,N_1244);
nor U1551 (N_1551,N_1015,N_562);
or U1552 (N_1552,N_6,N_1195);
and U1553 (N_1553,N_1235,N_1333);
nor U1554 (N_1554,In_2428,In_945);
nand U1555 (N_1555,N_1295,N_1204);
and U1556 (N_1556,N_1317,N_1398);
nor U1557 (N_1557,In_249,In_60);
nor U1558 (N_1558,N_1168,N_891);
nor U1559 (N_1559,N_1145,In_933);
or U1560 (N_1560,N_1355,N_651);
or U1561 (N_1561,N_1364,In_1898);
nand U1562 (N_1562,N_459,N_661);
and U1563 (N_1563,N_531,N_1312);
nand U1564 (N_1564,In_1277,N_1280);
and U1565 (N_1565,N_1375,N_833);
nand U1566 (N_1566,In_1896,N_952);
nor U1567 (N_1567,In_91,In_925);
nand U1568 (N_1568,N_647,N_1265);
and U1569 (N_1569,In_2081,N_636);
and U1570 (N_1570,N_755,N_1236);
and U1571 (N_1571,N_356,In_1199);
nor U1572 (N_1572,In_679,In_2135);
nand U1573 (N_1573,N_879,In_43);
nand U1574 (N_1574,N_485,N_706);
and U1575 (N_1575,N_104,In_1941);
or U1576 (N_1576,N_144,In_111);
nand U1577 (N_1577,In_840,N_1255);
nand U1578 (N_1578,In_1009,N_1035);
and U1579 (N_1579,In_283,In_995);
and U1580 (N_1580,N_575,N_780);
and U1581 (N_1581,In_2184,In_233);
nor U1582 (N_1582,In_1391,In_383);
nand U1583 (N_1583,In_1765,N_627);
or U1584 (N_1584,N_806,In_1109);
or U1585 (N_1585,N_1305,N_1342);
or U1586 (N_1586,N_1072,In_2127);
or U1587 (N_1587,N_1201,In_96);
and U1588 (N_1588,N_663,In_1539);
or U1589 (N_1589,N_1124,N_596);
nor U1590 (N_1590,In_1795,In_1798);
or U1591 (N_1591,N_234,In_1543);
nor U1592 (N_1592,N_1148,N_807);
nor U1593 (N_1593,In_2017,In_2098);
nand U1594 (N_1594,N_888,N_1301);
or U1595 (N_1595,In_1069,In_1657);
or U1596 (N_1596,N_501,In_2058);
xnor U1597 (N_1597,N_404,N_1336);
nand U1598 (N_1598,N_746,In_884);
or U1599 (N_1599,N_1315,In_238);
nand U1600 (N_1600,N_1514,N_1440);
and U1601 (N_1601,N_1558,N_1237);
nor U1602 (N_1602,In_437,In_1170);
or U1603 (N_1603,N_1469,N_1249);
nor U1604 (N_1604,N_1593,N_1598);
and U1605 (N_1605,N_129,N_457);
or U1606 (N_1606,In_767,In_1598);
xor U1607 (N_1607,In_1628,N_1458);
nand U1608 (N_1608,N_48,N_553);
nand U1609 (N_1609,In_1043,N_1211);
or U1610 (N_1610,N_1335,In_206);
nor U1611 (N_1611,N_873,N_1594);
nor U1612 (N_1612,N_644,N_638);
nor U1613 (N_1613,N_1098,N_775);
nor U1614 (N_1614,In_1047,N_1166);
or U1615 (N_1615,In_1585,N_412);
and U1616 (N_1616,N_1031,N_1041);
nand U1617 (N_1617,In_1195,N_1291);
and U1618 (N_1618,N_620,N_1209);
or U1619 (N_1619,In_1761,N_803);
and U1620 (N_1620,In_714,In_2265);
nor U1621 (N_1621,In_1027,N_1409);
nor U1622 (N_1622,N_556,N_397);
nand U1623 (N_1623,In_759,N_1581);
or U1624 (N_1624,N_1554,N_158);
or U1625 (N_1625,In_1054,N_1303);
nor U1626 (N_1626,N_383,N_1139);
or U1627 (N_1627,N_165,N_204);
and U1628 (N_1628,N_1205,In_1801);
and U1629 (N_1629,N_250,N_1389);
and U1630 (N_1630,In_1606,N_1430);
nand U1631 (N_1631,N_1075,N_1412);
or U1632 (N_1632,In_284,N_1360);
nor U1633 (N_1633,N_1361,In_1482);
and U1634 (N_1634,N_1574,N_1160);
nor U1635 (N_1635,N_731,N_970);
nor U1636 (N_1636,In_1053,N_119);
nor U1637 (N_1637,N_950,In_1356);
and U1638 (N_1638,In_1155,In_1531);
and U1639 (N_1639,N_1252,N_839);
nor U1640 (N_1640,In_2464,In_1404);
nand U1641 (N_1641,In_1854,N_1091);
nor U1642 (N_1642,N_1272,N_1387);
and U1643 (N_1643,N_1459,N_1543);
and U1644 (N_1644,In_1887,N_1308);
nor U1645 (N_1645,N_1014,N_98);
nor U1646 (N_1646,In_1121,N_1421);
or U1647 (N_1647,N_998,In_1590);
nand U1648 (N_1648,N_1569,N_688);
and U1649 (N_1649,N_1278,N_1200);
nand U1650 (N_1650,In_520,N_1492);
and U1651 (N_1651,N_1503,N_996);
nor U1652 (N_1652,N_1382,In_2340);
nor U1653 (N_1653,N_1556,In_644);
and U1654 (N_1654,In_1331,N_1589);
or U1655 (N_1655,In_2491,N_1434);
and U1656 (N_1656,N_1144,In_2238);
or U1657 (N_1657,In_2471,N_1147);
nand U1658 (N_1658,N_1560,In_298);
nand U1659 (N_1659,In_1330,N_881);
and U1660 (N_1660,In_63,N_1476);
nand U1661 (N_1661,In_616,N_1596);
nand U1662 (N_1662,N_463,In_808);
or U1663 (N_1663,In_1559,N_1219);
nor U1664 (N_1664,N_1573,N_577);
and U1665 (N_1665,In_2119,N_1539);
nor U1666 (N_1666,N_1505,N_1108);
nand U1667 (N_1667,N_1525,N_1580);
or U1668 (N_1668,In_1714,N_696);
and U1669 (N_1669,N_1546,N_1597);
or U1670 (N_1670,In_2085,In_2496);
nand U1671 (N_1671,In_1462,N_823);
and U1672 (N_1672,N_1122,N_162);
and U1673 (N_1673,N_1502,In_1923);
and U1674 (N_1674,In_2206,In_64);
and U1675 (N_1675,N_1473,N_1475);
and U1676 (N_1676,N_1214,N_704);
or U1677 (N_1677,N_1358,N_838);
and U1678 (N_1678,N_826,In_2333);
nand U1679 (N_1679,N_632,N_733);
and U1680 (N_1680,N_1498,N_1309);
nand U1681 (N_1681,N_613,In_1716);
nor U1682 (N_1682,N_1042,In_247);
or U1683 (N_1683,In_2389,N_1497);
nand U1684 (N_1684,N_1386,N_985);
nor U1685 (N_1685,N_1338,In_2151);
or U1686 (N_1686,N_1396,N_1270);
and U1687 (N_1687,N_909,N_1198);
nor U1688 (N_1688,In_783,N_1304);
nand U1689 (N_1689,N_1024,N_1327);
nand U1690 (N_1690,N_642,N_734);
nand U1691 (N_1691,N_1582,N_1284);
and U1692 (N_1692,N_1585,N_1376);
nand U1693 (N_1693,N_1414,N_540);
nand U1694 (N_1694,In_1891,N_867);
and U1695 (N_1695,N_1056,N_901);
nand U1696 (N_1696,N_813,N_687);
and U1697 (N_1697,N_570,In_771);
nand U1698 (N_1698,N_616,In_1732);
nand U1699 (N_1699,N_875,N_322);
and U1700 (N_1700,N_944,N_284);
nand U1701 (N_1701,In_606,N_917);
and U1702 (N_1702,N_231,N_1164);
nand U1703 (N_1703,In_962,N_1130);
nand U1704 (N_1704,In_421,N_1472);
nand U1705 (N_1705,N_961,N_1079);
or U1706 (N_1706,N_1453,In_2367);
or U1707 (N_1707,In_172,N_1553);
nor U1708 (N_1708,N_1545,N_1537);
nand U1709 (N_1709,N_825,In_413);
nor U1710 (N_1710,N_871,N_1086);
nor U1711 (N_1711,In_10,In_2412);
or U1712 (N_1712,N_667,N_1424);
nor U1713 (N_1713,N_1590,In_1682);
nor U1714 (N_1714,N_898,In_1847);
nand U1715 (N_1715,In_1678,N_1167);
nor U1716 (N_1716,N_369,N_1368);
and U1717 (N_1717,In_316,In_508);
or U1718 (N_1718,N_1299,N_895);
nor U1719 (N_1719,N_869,N_1465);
and U1720 (N_1720,N_1400,In_755);
nand U1721 (N_1721,N_1531,In_2319);
or U1722 (N_1722,N_1579,N_1474);
nand U1723 (N_1723,N_751,In_1257);
nand U1724 (N_1724,N_1540,N_1154);
or U1725 (N_1725,N_1046,N_1257);
nor U1726 (N_1726,In_1412,In_915);
nand U1727 (N_1727,In_429,N_1587);
nor U1728 (N_1728,N_1487,N_1155);
and U1729 (N_1729,N_1061,N_740);
nand U1730 (N_1730,N_1331,In_1799);
nor U1731 (N_1731,In_1625,N_1271);
nand U1732 (N_1732,N_756,N_922);
nand U1733 (N_1733,N_1549,In_2044);
nand U1734 (N_1734,N_1488,N_1240);
nand U1735 (N_1735,In_1168,N_1276);
nand U1736 (N_1736,In_212,N_475);
and U1737 (N_1737,N_758,In_2010);
nor U1738 (N_1738,N_1286,N_406);
nor U1739 (N_1739,In_1599,In_327);
nand U1740 (N_1740,N_1442,N_1470);
or U1741 (N_1741,In_1930,N_1245);
nand U1742 (N_1742,N_1099,In_2228);
and U1743 (N_1743,N_1002,N_1563);
or U1744 (N_1744,N_1551,N_277);
and U1745 (N_1745,N_1455,In_2407);
nor U1746 (N_1746,N_1445,In_907);
and U1747 (N_1747,N_1541,N_1584);
nand U1748 (N_1748,In_55,N_1471);
nor U1749 (N_1749,N_426,N_1489);
nand U1750 (N_1750,N_1527,N_1111);
xor U1751 (N_1751,In_557,N_1169);
nor U1752 (N_1752,N_1524,N_1565);
and U1753 (N_1753,N_1491,N_1196);
and U1754 (N_1754,N_802,N_707);
xor U1755 (N_1755,In_1596,N_1510);
nor U1756 (N_1756,In_1205,N_761);
or U1757 (N_1757,In_277,N_1365);
nand U1758 (N_1758,In_2454,N_1428);
and U1759 (N_1759,N_1007,N_712);
or U1760 (N_1760,In_961,In_846);
nor U1761 (N_1761,N_401,N_1532);
or U1762 (N_1762,N_1564,N_232);
nand U1763 (N_1763,N_1246,N_1289);
nor U1764 (N_1764,N_1112,N_421);
nor U1765 (N_1765,In_205,N_1319);
and U1766 (N_1766,In_496,N_1444);
nand U1767 (N_1767,N_1142,N_967);
or U1768 (N_1768,N_748,N_1354);
nand U1769 (N_1769,N_349,In_2355);
nor U1770 (N_1770,N_1116,N_1529);
and U1771 (N_1771,N_583,N_1501);
nand U1772 (N_1772,N_1561,In_2302);
and U1773 (N_1773,N_1425,N_170);
nor U1774 (N_1774,N_1004,N_1220);
nor U1775 (N_1775,N_621,N_782);
or U1776 (N_1776,In_1323,N_519);
nand U1777 (N_1777,In_1913,N_1203);
nor U1778 (N_1778,In_1722,N_1123);
nand U1779 (N_1779,N_1030,N_1181);
nand U1780 (N_1780,N_759,N_1595);
and U1781 (N_1781,N_639,N_468);
or U1782 (N_1782,N_1485,In_663);
nor U1783 (N_1783,N_1550,N_1185);
or U1784 (N_1784,In_1232,N_1206);
or U1785 (N_1785,N_1405,N_1377);
nand U1786 (N_1786,In_2267,N_625);
or U1787 (N_1787,N_949,N_1260);
nor U1788 (N_1788,In_373,N_1223);
nor U1789 (N_1789,In_451,N_1117);
nand U1790 (N_1790,N_1583,In_594);
and U1791 (N_1791,In_599,N_1330);
and U1792 (N_1792,In_288,N_1578);
nor U1793 (N_1793,N_859,In_329);
and U1794 (N_1794,N_1432,In_2159);
or U1795 (N_1795,N_305,In_1092);
nand U1796 (N_1796,In_1387,N_1230);
or U1797 (N_1797,N_675,N_1566);
or U1798 (N_1798,In_484,N_1411);
nand U1799 (N_1799,N_1057,In_1249);
nor U1800 (N_1800,N_1776,N_1535);
and U1801 (N_1801,N_432,N_1461);
and U1802 (N_1802,N_1062,In_370);
nor U1803 (N_1803,N_1624,N_374);
or U1804 (N_1804,N_1710,N_974);
nand U1805 (N_1805,N_1625,In_494);
xor U1806 (N_1806,N_1454,N_630);
and U1807 (N_1807,N_1570,N_1138);
or U1808 (N_1808,N_560,N_1179);
nand U1809 (N_1809,N_1384,N_1456);
nand U1810 (N_1810,N_1522,N_1619);
nand U1811 (N_1811,In_875,N_1659);
or U1812 (N_1812,In_975,N_1774);
or U1813 (N_1813,N_363,N_1426);
nor U1814 (N_1814,N_1747,N_1394);
nor U1815 (N_1815,In_873,N_886);
nand U1816 (N_1816,N_1266,N_1686);
and U1817 (N_1817,N_1763,In_1000);
or U1818 (N_1818,N_1242,In_989);
and U1819 (N_1819,N_1691,In_1088);
or U1820 (N_1820,In_518,N_1293);
nor U1821 (N_1821,N_1146,In_456);
or U1822 (N_1822,N_1642,N_1137);
or U1823 (N_1823,In_2062,N_923);
or U1824 (N_1824,In_2117,N_1302);
nor U1825 (N_1825,N_1359,N_1517);
or U1826 (N_1826,In_1456,In_596);
or U1827 (N_1827,N_766,N_1076);
or U1828 (N_1828,N_892,In_1634);
and U1829 (N_1829,N_1542,In_1483);
and U1830 (N_1830,N_1287,N_932);
or U1831 (N_1831,In_1236,N_1521);
or U1832 (N_1832,In_554,N_1727);
nor U1833 (N_1833,N_1324,N_1533);
nand U1834 (N_1834,N_1017,N_1158);
xnor U1835 (N_1835,N_1795,N_1643);
nor U1836 (N_1836,N_1334,N_1407);
nand U1837 (N_1837,N_161,N_1221);
and U1838 (N_1838,In_642,N_1136);
nor U1839 (N_1839,In_674,N_1133);
and U1840 (N_1840,N_1264,In_762);
nor U1841 (N_1841,N_1314,N_1761);
or U1842 (N_1842,In_1753,N_1788);
or U1843 (N_1843,N_1,N_1785);
and U1844 (N_1844,N_217,N_1651);
and U1845 (N_1845,N_1682,N_1054);
or U1846 (N_1846,N_1256,In_1302);
and U1847 (N_1847,N_1339,N_664);
and U1848 (N_1848,N_680,N_1706);
nand U1849 (N_1849,In_1804,N_1673);
nand U1850 (N_1850,N_1443,N_1660);
nor U1851 (N_1851,N_1053,N_1423);
and U1852 (N_1852,In_1123,In_974);
or U1853 (N_1853,N_296,N_1758);
nor U1854 (N_1854,N_1602,N_1599);
or U1855 (N_1855,N_715,N_488);
and U1856 (N_1856,N_1757,N_1562);
or U1857 (N_1857,N_1520,N_1571);
or U1858 (N_1858,N_1496,In_861);
and U1859 (N_1859,N_1495,N_769);
nor U1860 (N_1860,N_19,N_1450);
nor U1861 (N_1861,In_1201,N_1605);
nor U1862 (N_1862,N_1151,N_1016);
or U1863 (N_1863,N_1552,N_1684);
nor U1864 (N_1864,N_1499,N_1600);
nor U1865 (N_1865,N_965,N_1717);
xor U1866 (N_1866,In_2156,N_1357);
nor U1867 (N_1867,In_1763,N_1320);
nand U1868 (N_1868,N_1351,N_1478);
and U1869 (N_1869,N_1748,N_973);
or U1870 (N_1870,N_1131,N_1313);
and U1871 (N_1871,N_1745,N_657);
nor U1872 (N_1872,In_1490,N_1751);
or U1873 (N_1873,N_1764,N_1262);
nor U1874 (N_1874,N_1500,N_1712);
nor U1875 (N_1875,In_1947,In_1550);
and U1876 (N_1876,N_1739,N_1631);
nor U1877 (N_1877,N_1713,N_614);
or U1878 (N_1878,In_1094,N_1231);
or U1879 (N_1879,N_1422,N_502);
nand U1880 (N_1880,N_1796,N_1729);
and U1881 (N_1881,N_1457,N_1352);
and U1882 (N_1882,N_980,N_1534);
nand U1883 (N_1883,N_1055,N_1121);
nand U1884 (N_1884,In_434,N_1679);
nor U1885 (N_1885,N_1363,N_1756);
and U1886 (N_1886,In_534,N_645);
and U1887 (N_1887,N_1202,N_1481);
or U1888 (N_1888,N_1027,N_685);
nand U1889 (N_1889,N_1467,In_36);
nand U1890 (N_1890,N_1513,N_1744);
nor U1891 (N_1891,N_1466,N_1134);
or U1892 (N_1892,N_1752,N_1300);
nand U1893 (N_1893,N_1058,N_1792);
and U1894 (N_1894,N_1462,N_1702);
nand U1895 (N_1895,In_2335,N_1725);
nor U1896 (N_1896,In_471,N_1069);
and U1897 (N_1897,N_1484,N_1174);
or U1898 (N_1898,N_1380,N_1087);
and U1899 (N_1899,N_456,N_752);
and U1900 (N_1900,In_711,N_1678);
and U1901 (N_1901,N_1618,In_1339);
or U1902 (N_1902,N_1490,N_1616);
nand U1903 (N_1903,N_1438,N_1509);
nor U1904 (N_1904,N_1175,N_1538);
nand U1905 (N_1905,N_790,N_1685);
nand U1906 (N_1906,N_1567,N_1746);
and U1907 (N_1907,N_1617,N_1479);
or U1908 (N_1908,N_1775,N_1383);
nor U1909 (N_1909,In_636,N_729);
nand U1910 (N_1910,In_1465,N_1612);
nand U1911 (N_1911,N_1720,In_1226);
and U1912 (N_1912,N_1296,N_902);
nand U1913 (N_1913,In_466,N_1762);
nand U1914 (N_1914,N_1482,In_952);
nand U1915 (N_1915,N_1039,In_390);
and U1916 (N_1916,N_1568,N_1635);
nor U1917 (N_1917,N_1704,In_120);
and U1918 (N_1918,In_169,N_1692);
or U1919 (N_1919,N_1420,N_299);
nand U1920 (N_1920,N_1011,N_1222);
and U1921 (N_1921,In_963,N_1464);
nand U1922 (N_1922,N_1609,N_1408);
or U1923 (N_1923,N_1734,N_1715);
nor U1924 (N_1924,N_149,N_1634);
or U1925 (N_1925,N_361,N_1614);
nand U1926 (N_1926,N_1772,N_1447);
or U1927 (N_1927,N_1228,N_1771);
or U1928 (N_1928,N_1113,N_1576);
and U1929 (N_1929,In_2132,N_1786);
nand U1930 (N_1930,In_116,N_1468);
or U1931 (N_1931,N_1460,In_903);
or U1932 (N_1932,N_1480,N_738);
or U1933 (N_1933,N_646,In_1661);
and U1934 (N_1934,N_650,N_1652);
or U1935 (N_1935,In_465,N_1668);
nand U1936 (N_1936,N_1263,N_1391);
or U1937 (N_1937,N_1693,N_918);
nand U1938 (N_1938,N_1696,N_1234);
or U1939 (N_1939,N_1390,In_2401);
nor U1940 (N_1940,N_808,N_1749);
or U1941 (N_1941,N_1664,N_818);
and U1942 (N_1942,N_1705,N_1791);
xor U1943 (N_1943,N_1186,N_1733);
nand U1944 (N_1944,N_1028,N_1716);
and U1945 (N_1945,N_1451,In_2456);
nand U1946 (N_1946,N_1187,N_1274);
nor U1947 (N_1947,N_1787,N_586);
and U1948 (N_1948,N_1658,N_1688);
nor U1949 (N_1949,In_377,N_1402);
nand U1950 (N_1950,N_1507,In_1290);
or U1951 (N_1951,N_1059,N_1779);
and U1952 (N_1952,N_1268,N_1183);
and U1953 (N_1953,N_1511,N_1799);
or U1954 (N_1954,In_1646,N_1229);
nand U1955 (N_1955,N_1640,N_1689);
nand U1956 (N_1956,N_1780,N_1225);
and U1957 (N_1957,N_1697,N_1768);
nor U1958 (N_1958,In_1895,N_1374);
or U1959 (N_1959,In_1740,N_979);
or U1960 (N_1960,N_1738,N_1233);
nand U1961 (N_1961,N_1449,N_1700);
or U1962 (N_1962,In_944,N_1431);
and U1963 (N_1963,In_142,N_1329);
xnor U1964 (N_1964,N_981,N_1418);
or U1965 (N_1965,N_1415,N_1657);
nand U1966 (N_1966,N_1740,N_1639);
nand U1967 (N_1967,In_896,N_1645);
nand U1968 (N_1968,N_1680,In_1976);
or U1969 (N_1969,N_1504,N_1159);
and U1970 (N_1970,N_842,In_1159);
and U1971 (N_1971,In_1548,N_1767);
nand U1972 (N_1972,N_38,N_389);
or U1973 (N_1973,N_703,In_720);
nor U1974 (N_1974,N_1603,N_1090);
nor U1975 (N_1975,N_41,N_439);
and U1976 (N_1976,N_44,In_1815);
and U1977 (N_1977,In_1614,N_1703);
nor U1978 (N_1978,In_754,N_1721);
and U1979 (N_1979,N_1346,N_1604);
nor U1980 (N_1980,In_803,N_1675);
nand U1981 (N_1981,N_1106,N_1104);
and U1982 (N_1982,N_1687,N_817);
and U1983 (N_1983,N_1575,N_1493);
nor U1984 (N_1984,In_1927,N_1102);
or U1985 (N_1985,N_1385,N_1769);
and U1986 (N_1986,N_1674,In_1477);
and U1987 (N_1987,N_22,N_1064);
and U1988 (N_1988,N_1281,N_1040);
or U1989 (N_1989,N_1406,N_173);
nand U1990 (N_1990,N_1646,N_1068);
nor U1991 (N_1991,N_1736,N_1006);
and U1992 (N_1992,N_603,N_939);
nor U1993 (N_1993,N_1722,In_1112);
and U1994 (N_1994,N_1777,N_1663);
nor U1995 (N_1995,In_2165,N_1110);
or U1996 (N_1996,N_1217,N_1592);
nand U1997 (N_1997,In_900,N_1452);
and U1998 (N_1998,In_701,N_1163);
nor U1999 (N_1999,N_1753,N_1718);
or U2000 (N_2000,N_1923,N_1881);
nand U2001 (N_2001,N_1848,N_1913);
nor U2002 (N_2002,N_1760,In_592);
or U2003 (N_2003,N_1918,N_1413);
nand U2004 (N_2004,N_1586,N_1427);
nor U2005 (N_2005,N_1078,N_1804);
or U2006 (N_2006,N_1790,N_1676);
nor U2007 (N_2007,N_1963,N_1935);
nand U2008 (N_2008,In_328,N_1677);
or U2009 (N_2009,N_1856,N_569);
or U2010 (N_2010,In_1850,In_1346);
and U2011 (N_2011,N_1750,N_1661);
nor U2012 (N_2012,N_812,N_649);
nor U2013 (N_2013,N_988,N_1983);
or U2014 (N_2014,N_1809,N_1961);
nor U2015 (N_2015,In_381,N_1026);
nand U2016 (N_2016,N_235,In_1002);
or U2017 (N_2017,N_56,N_1820);
nand U2018 (N_2018,N_1666,N_1816);
nand U2019 (N_2019,N_1759,N_1337);
and U2020 (N_2020,N_1726,In_1334);
and U2021 (N_2021,N_1506,N_1261);
nor U2022 (N_2022,N_1857,N_1912);
nor U2023 (N_2023,In_1064,N_580);
or U2024 (N_2024,N_1735,In_2422);
or U2025 (N_2025,In_634,N_1934);
nand U2026 (N_2026,In_882,N_1942);
or U2027 (N_2027,N_1823,N_1832);
and U2028 (N_2028,N_1670,N_1948);
nand U2029 (N_2029,In_411,N_786);
and U2030 (N_2030,N_1694,N_1866);
nand U2031 (N_2031,N_1793,N_1101);
and U2032 (N_2032,N_1519,N_1698);
nand U2033 (N_2033,N_1800,N_1837);
nand U2034 (N_2034,N_1184,N_1858);
nand U2035 (N_2035,N_1914,N_1885);
nand U2036 (N_2036,N_1836,N_999);
or U2037 (N_2037,N_1623,In_1603);
and U2038 (N_2038,N_1633,N_1784);
nor U2039 (N_2039,N_1681,N_1655);
nor U2040 (N_2040,N_1250,N_1886);
nand U2041 (N_2041,N_1362,N_1731);
or U2042 (N_2042,N_1901,N_1824);
and U2043 (N_2043,N_1000,N_1714);
nand U2044 (N_2044,N_1446,In_17);
or U2045 (N_2045,N_1251,N_1854);
nor U2046 (N_2046,N_1656,N_1009);
and U2047 (N_2047,N_1815,N_843);
and U2048 (N_2048,N_1672,In_1424);
or U2049 (N_2049,N_1628,N_1765);
or U2050 (N_2050,N_1083,N_1755);
or U2051 (N_2051,N_1907,N_1778);
and U2052 (N_2052,N_1477,In_1647);
nand U2053 (N_2053,N_1872,N_1494);
and U2054 (N_2054,N_1821,In_573);
and U2055 (N_2055,N_1884,N_1835);
nor U2056 (N_2056,In_1017,N_1958);
nor U2057 (N_2057,N_1805,N_1052);
nor U2058 (N_2058,N_1649,N_1283);
or U2059 (N_2059,In_1022,N_499);
or U2060 (N_2060,N_1833,N_1548);
and U2061 (N_2061,N_1921,In_684);
or U2062 (N_2062,N_1648,N_1990);
and U2063 (N_2063,N_1879,N_1647);
or U2064 (N_2064,N_1911,N_1996);
nor U2065 (N_2065,N_1536,N_1944);
nor U2066 (N_2066,N_1895,N_1973);
nand U2067 (N_2067,In_562,N_1976);
and U2068 (N_2068,In_1394,N_1906);
xnor U2069 (N_2069,N_1813,N_1708);
and U2070 (N_2070,N_1993,N_1789);
nand U2071 (N_2071,N_1238,N_1518);
or U2072 (N_2072,N_1830,N_1898);
or U2073 (N_2073,N_1707,N_1900);
nor U2074 (N_2074,N_1318,N_288);
and U2075 (N_2075,N_1213,In_388);
or U2076 (N_2076,In_918,N_1241);
nor U2077 (N_2077,N_1436,N_1530);
nand U2078 (N_2078,N_1340,N_1897);
nor U2079 (N_2079,N_1927,N_1770);
and U2080 (N_2080,N_1860,N_1851);
or U2081 (N_2081,N_1591,N_1831);
or U2082 (N_2082,N_1626,N_1227);
nor U2083 (N_2083,N_1577,N_1399);
nor U2084 (N_2084,N_1994,N_1326);
and U2085 (N_2085,N_1435,N_1671);
nand U2086 (N_2086,In_2386,In_698);
or U2087 (N_2087,N_1847,N_1127);
nand U2088 (N_2088,N_1743,N_1957);
and U2089 (N_2089,N_1641,N_1938);
or U2090 (N_2090,N_1807,N_1806);
or U2091 (N_2091,N_181,N_1855);
and U2092 (N_2092,N_1867,N_1933);
and U2093 (N_2093,N_1512,N_1437);
nor U2094 (N_2094,In_1036,N_1797);
nor U2095 (N_2095,N_907,N_1995);
nand U2096 (N_2096,N_1699,In_1810);
nand U2097 (N_2097,N_1878,N_1638);
nor U2098 (N_2098,N_1644,N_1925);
nand U2099 (N_2099,N_1987,N_1992);
nor U2100 (N_2100,N_1695,N_1819);
nor U2101 (N_2101,In_1987,N_1728);
or U2102 (N_2102,N_1931,N_1985);
or U2103 (N_2103,N_1873,In_1867);
nand U2104 (N_2104,In_1756,In_1950);
nor U2105 (N_2105,In_358,N_1378);
nor U2106 (N_2106,In_2266,N_1930);
or U2107 (N_2107,N_1723,N_1846);
and U2108 (N_2108,N_1191,N_1811);
nor U2109 (N_2109,N_1941,N_1975);
nand U2110 (N_2110,N_1834,N_1862);
nor U2111 (N_2111,N_1915,N_1711);
or U2112 (N_2112,N_1888,N_1667);
nand U2113 (N_2113,N_1654,N_1621);
or U2114 (N_2114,N_1952,N_1801);
and U2115 (N_2115,N_1630,N_1909);
nand U2116 (N_2116,N_1353,N_1732);
and U2117 (N_2117,N_834,N_1964);
or U2118 (N_2118,N_1874,N_1523);
nor U2119 (N_2119,In_344,N_1606);
or U2120 (N_2120,N_1890,In_1368);
nor U2121 (N_2121,N_1297,N_1861);
or U2122 (N_2122,N_1248,N_1140);
or U2123 (N_2123,N_380,N_1920);
nor U2124 (N_2124,N_1620,N_1808);
or U2125 (N_2125,N_1939,N_1417);
or U2126 (N_2126,N_1588,N_1916);
or U2127 (N_2127,N_1889,N_1627);
nand U2128 (N_2128,N_1528,In_1189);
and U2129 (N_2129,N_415,N_1853);
nor U2130 (N_2130,N_1843,N_1719);
or U2131 (N_2131,In_445,N_1863);
nand U2132 (N_2132,N_1410,N_1970);
nor U2133 (N_2133,N_1908,N_1959);
or U2134 (N_2134,In_2126,N_1842);
and U2135 (N_2135,N_1947,N_1653);
and U2136 (N_2136,N_1267,N_1803);
nand U2137 (N_2137,N_1094,N_665);
and U2138 (N_2138,N_1852,N_1962);
nor U2139 (N_2139,N_1929,N_1636);
nor U2140 (N_2140,N_836,N_1783);
nand U2141 (N_2141,N_1960,N_1972);
or U2142 (N_2142,N_1829,N_1928);
or U2143 (N_2143,N_1215,N_536);
and U2144 (N_2144,In_1945,In_1997);
nor U2145 (N_2145,In_2263,N_1037);
nand U2146 (N_2146,In_1494,In_393);
nor U2147 (N_2147,N_1943,N_1984);
nor U2148 (N_2148,N_1559,N_1392);
nor U2149 (N_2149,N_1429,N_1419);
xnor U2150 (N_2150,N_986,N_1966);
and U2151 (N_2151,N_1611,N_1956);
nor U2152 (N_2152,N_1969,N_1544);
nand U2153 (N_2153,In_1942,In_2377);
nand U2154 (N_2154,N_1416,N_655);
and U2155 (N_2155,N_563,N_320);
nand U2156 (N_2156,N_1812,N_1839);
nor U2157 (N_2157,N_725,N_1572);
and U2158 (N_2158,N_1817,N_1876);
nor U2159 (N_2159,N_1986,In_2138);
or U2160 (N_2160,N_1991,N_1865);
nor U2161 (N_2161,N_1981,N_1601);
or U2162 (N_2162,N_1683,In_29);
or U2163 (N_2163,N_1486,N_1547);
or U2164 (N_2164,In_253,N_1439);
nand U2165 (N_2165,N_953,N_1622);
nand U2166 (N_2166,N_1115,N_1893);
and U2167 (N_2167,N_805,N_1869);
nand U2168 (N_2168,N_1974,N_1508);
or U2169 (N_2169,N_1950,N_1999);
nor U2170 (N_2170,N_1850,N_1742);
and U2171 (N_2171,N_699,N_1404);
xor U2172 (N_2172,N_1965,N_1650);
or U2173 (N_2173,N_1347,N_1882);
nand U2174 (N_2174,N_1741,N_1905);
nand U2175 (N_2175,N_1526,N_1838);
nand U2176 (N_2176,N_1690,N_797);
and U2177 (N_2177,N_1818,In_976);
nand U2178 (N_2178,N_1880,N_1978);
or U2179 (N_2179,N_1868,In_1428);
nor U2180 (N_2180,N_1170,N_1613);
nand U2181 (N_2181,N_1871,N_1903);
nand U2182 (N_2182,N_1212,N_1401);
nand U2183 (N_2183,N_924,N_1926);
nor U2184 (N_2184,N_1988,N_1946);
nand U2185 (N_2185,In_2492,N_309);
nand U2186 (N_2186,N_1285,N_281);
nor U2187 (N_2187,N_1798,In_92);
or U2188 (N_2188,N_1949,N_1782);
nand U2189 (N_2189,In_2167,In_1635);
nor U2190 (N_2190,N_1980,N_1730);
nor U2191 (N_2191,N_1977,N_1955);
and U2192 (N_2192,N_172,N_1924);
or U2193 (N_2193,N_1766,N_916);
or U2194 (N_2194,N_1937,N_268);
nand U2195 (N_2195,N_1828,N_1936);
or U2196 (N_2196,N_1463,N_1841);
and U2197 (N_2197,N_1162,N_1632);
and U2198 (N_2198,N_1615,N_1932);
nor U2199 (N_2199,N_1724,N_396);
and U2200 (N_2200,N_2139,N_2080);
and U2201 (N_2201,N_2022,N_1709);
nor U2202 (N_2202,N_2165,N_2060);
or U2203 (N_2203,N_2064,N_2023);
nor U2204 (N_2204,N_1968,N_2054);
xnor U2205 (N_2205,N_1665,N_2052);
nand U2206 (N_2206,N_2051,N_2142);
xnor U2207 (N_2207,N_2078,N_2172);
and U2208 (N_2208,N_2129,N_1366);
nor U2209 (N_2209,N_2162,N_1864);
nor U2210 (N_2210,N_1143,N_2081);
nor U2211 (N_2211,N_2163,N_2041);
or U2212 (N_2212,N_1997,N_2198);
and U2213 (N_2213,N_1902,N_2176);
or U2214 (N_2214,N_2017,N_1892);
and U2215 (N_2215,N_2106,N_1516);
nand U2216 (N_2216,N_2047,N_2079);
and U2217 (N_2217,N_2055,N_2149);
or U2218 (N_2218,N_555,N_2037);
nor U2219 (N_2219,N_2007,N_2192);
nor U2220 (N_2220,In_1408,N_2164);
and U2221 (N_2221,N_2018,N_1701);
and U2222 (N_2222,N_865,N_2095);
nor U2223 (N_2223,N_2133,N_2073);
or U2224 (N_2224,N_326,N_2189);
nand U2225 (N_2225,N_2045,N_1032);
nand U2226 (N_2226,N_1953,N_2148);
and U2227 (N_2227,N_2026,N_2025);
and U2228 (N_2228,N_2152,N_2140);
nand U2229 (N_2229,N_1607,N_2085);
nand U2230 (N_2230,N_2027,N_2090);
and U2231 (N_2231,In_980,N_2053);
and U2232 (N_2232,N_2115,N_2122);
nand U2233 (N_2233,N_1870,N_2035);
nor U2234 (N_2234,N_2084,N_2182);
nor U2235 (N_2235,N_2002,N_1669);
and U2236 (N_2236,In_1711,N_2087);
and U2237 (N_2237,N_1971,N_2157);
and U2238 (N_2238,N_1372,N_2156);
nand U2239 (N_2239,N_1951,N_2150);
nor U2240 (N_2240,N_2160,N_2098);
nand U2241 (N_2241,N_2191,N_1825);
nand U2242 (N_2242,N_2030,N_2061);
and U2243 (N_2243,N_2128,N_2135);
or U2244 (N_2244,N_2102,N_2067);
nor U2245 (N_2245,N_2144,N_2046);
nor U2246 (N_2246,N_2119,N_2174);
nand U2247 (N_2247,In_1280,N_2170);
nand U2248 (N_2248,N_2190,N_2092);
nor U2249 (N_2249,N_2010,N_283);
and U2250 (N_2250,N_2063,N_2159);
nand U2251 (N_2251,N_2101,N_1849);
nor U2252 (N_2252,N_2068,N_2145);
and U2253 (N_2253,N_2109,N_2187);
nand U2254 (N_2254,N_1555,N_1448);
nor U2255 (N_2255,N_2143,N_1917);
and U2256 (N_2256,N_418,N_2088);
nand U2257 (N_2257,N_2108,N_1826);
nand U2258 (N_2258,N_2123,N_1194);
and U2259 (N_2259,N_1989,N_1393);
or U2260 (N_2260,N_2118,N_1845);
nor U2261 (N_2261,N_1940,N_2169);
nand U2262 (N_2262,N_2093,N_2071);
nor U2263 (N_2263,N_2036,N_2146);
nand U2264 (N_2264,N_2040,N_2062);
nand U2265 (N_2265,N_2117,N_2179);
or U2266 (N_2266,N_2141,N_2197);
and U2267 (N_2267,N_1433,N_148);
and U2268 (N_2268,N_2155,N_2094);
nand U2269 (N_2269,N_1349,N_1998);
or U2270 (N_2270,N_2183,N_2012);
and U2271 (N_2271,N_1979,In_313);
nand U2272 (N_2272,N_2136,In_1693);
or U2273 (N_2273,N_2154,N_2011);
and U2274 (N_2274,N_789,N_2181);
nor U2275 (N_2275,N_2184,N_1292);
nor U2276 (N_2276,N_2056,N_2089);
nand U2277 (N_2277,N_2173,N_1794);
nand U2278 (N_2278,N_2131,N_1754);
nand U2279 (N_2279,N_1919,N_509);
nand U2280 (N_2280,N_1883,N_2130);
and U2281 (N_2281,N_2199,N_1441);
or U2282 (N_2282,N_2058,N_2075);
nand U2283 (N_2283,N_2104,N_416);
and U2284 (N_2284,N_2153,N_2147);
or U2285 (N_2285,N_2004,N_2057);
nor U2286 (N_2286,In_1240,N_1557);
nor U2287 (N_2287,N_2194,N_2166);
nor U2288 (N_2288,N_2070,N_2178);
or U2289 (N_2289,N_2097,N_1904);
and U2290 (N_2290,N_2031,N_2014);
nand U2291 (N_2291,N_2114,N_957);
nand U2292 (N_2292,N_2161,N_1967);
nor U2293 (N_2293,N_2121,N_1844);
or U2294 (N_2294,N_2005,N_1515);
nand U2295 (N_2295,N_2065,N_2124);
nor U2296 (N_2296,N_2193,N_1827);
nor U2297 (N_2297,N_2076,N_2167);
and U2298 (N_2298,N_2059,N_2105);
nor U2299 (N_2299,N_2015,N_1608);
or U2300 (N_2300,N_1737,N_2126);
or U2301 (N_2301,N_2049,N_2033);
and U2302 (N_2302,N_2008,N_2134);
or U2303 (N_2303,N_763,N_2069);
and U2304 (N_2304,N_2168,N_2074);
nand U2305 (N_2305,N_2066,N_2107);
and U2306 (N_2306,In_2000,N_1840);
or U2307 (N_2307,N_2028,N_2020);
and U2308 (N_2308,N_2116,N_2110);
nand U2309 (N_2309,N_1822,N_2111);
xor U2310 (N_2310,N_1922,N_2096);
and U2311 (N_2311,N_2175,N_2077);
or U2312 (N_2312,N_2132,N_2083);
nor U2313 (N_2313,N_2006,N_2188);
nor U2314 (N_2314,N_2137,N_2082);
or U2315 (N_2315,N_1875,N_2021);
or U2316 (N_2316,N_1877,N_2072);
and U2317 (N_2317,N_2050,N_1899);
nand U2318 (N_2318,N_2038,N_1859);
nor U2319 (N_2319,N_2125,N_1637);
and U2320 (N_2320,N_1887,In_2087);
and U2321 (N_2321,N_2024,N_2112);
nand U2322 (N_2322,N_2171,N_987);
or U2323 (N_2323,N_1945,N_1954);
and U2324 (N_2324,N_2091,N_1896);
and U2325 (N_2325,N_2099,N_2186);
nand U2326 (N_2326,N_1403,N_1483);
nor U2327 (N_2327,N_1910,N_1802);
nand U2328 (N_2328,N_2000,N_2113);
nand U2329 (N_2329,N_1781,N_2003);
and U2330 (N_2330,N_2043,N_2195);
nor U2331 (N_2331,N_1814,N_2120);
or U2332 (N_2332,N_1306,N_1894);
or U2333 (N_2333,N_2009,N_2086);
nor U2334 (N_2334,N_2177,N_2016);
and U2335 (N_2335,N_2185,N_2180);
and U2336 (N_2336,N_2158,N_2100);
nand U2337 (N_2337,N_2103,N_2001);
nor U2338 (N_2338,N_2196,N_2034);
and U2339 (N_2339,N_1082,N_2127);
nand U2340 (N_2340,N_1273,N_2013);
and U2341 (N_2341,N_1810,N_1773);
nor U2342 (N_2342,N_854,N_1982);
or U2343 (N_2343,N_2039,N_2044);
nand U2344 (N_2344,In_1636,N_2138);
or U2345 (N_2345,N_2048,N_1610);
nand U2346 (N_2346,N_2032,N_1662);
nor U2347 (N_2347,N_2019,N_2151);
nor U2348 (N_2348,N_1629,N_1891);
and U2349 (N_2349,N_2029,N_2042);
and U2350 (N_2350,N_2052,N_2045);
and U2351 (N_2351,N_2026,N_2192);
nand U2352 (N_2352,N_1516,In_1693);
or U2353 (N_2353,N_2189,N_2070);
nand U2354 (N_2354,N_2054,N_2116);
and U2355 (N_2355,N_2198,N_2111);
nand U2356 (N_2356,N_1896,N_1393);
nand U2357 (N_2357,N_2161,N_2099);
and U2358 (N_2358,N_2029,N_2184);
nand U2359 (N_2359,N_2199,N_2032);
nand U2360 (N_2360,N_2069,N_2134);
nand U2361 (N_2361,N_2132,N_2086);
nor U2362 (N_2362,N_2049,N_2149);
nand U2363 (N_2363,N_2113,N_1849);
nand U2364 (N_2364,In_313,N_1629);
nor U2365 (N_2365,N_2182,N_2035);
nand U2366 (N_2366,N_2147,N_2000);
nor U2367 (N_2367,N_2006,N_1403);
or U2368 (N_2368,N_2041,N_2068);
nor U2369 (N_2369,N_2078,N_2100);
or U2370 (N_2370,N_2014,N_1864);
nand U2371 (N_2371,N_2072,N_2094);
and U2372 (N_2372,N_2004,N_2154);
nand U2373 (N_2373,N_1555,N_2016);
nand U2374 (N_2374,N_2099,N_2158);
nor U2375 (N_2375,N_2027,N_2002);
or U2376 (N_2376,N_1979,N_2000);
and U2377 (N_2377,N_2074,N_2143);
and U2378 (N_2378,N_865,In_2087);
xnor U2379 (N_2379,N_2193,N_2019);
and U2380 (N_2380,N_148,N_1273);
and U2381 (N_2381,N_2157,N_2090);
or U2382 (N_2382,N_2099,N_2049);
or U2383 (N_2383,N_2188,N_1899);
or U2384 (N_2384,N_2138,N_2039);
nor U2385 (N_2385,N_1629,N_1896);
nor U2386 (N_2386,N_2084,N_2031);
nand U2387 (N_2387,N_1669,N_1637);
nor U2388 (N_2388,N_2167,N_2080);
or U2389 (N_2389,N_865,N_2199);
nor U2390 (N_2390,N_2042,N_2002);
nand U2391 (N_2391,N_2069,N_2079);
nand U2392 (N_2392,N_1802,N_2155);
nand U2393 (N_2393,N_2148,N_1945);
nand U2394 (N_2394,N_2070,N_1945);
and U2395 (N_2395,N_1403,N_2154);
and U2396 (N_2396,N_2093,N_2096);
or U2397 (N_2397,N_326,N_2142);
or U2398 (N_2398,N_2148,N_1840);
nor U2399 (N_2399,N_2005,N_2159);
or U2400 (N_2400,N_2326,N_2225);
nor U2401 (N_2401,N_2209,N_2360);
or U2402 (N_2402,N_2345,N_2297);
or U2403 (N_2403,N_2372,N_2342);
nor U2404 (N_2404,N_2281,N_2299);
and U2405 (N_2405,N_2271,N_2266);
and U2406 (N_2406,N_2368,N_2277);
nand U2407 (N_2407,N_2397,N_2331);
and U2408 (N_2408,N_2233,N_2239);
nor U2409 (N_2409,N_2229,N_2340);
and U2410 (N_2410,N_2384,N_2390);
nand U2411 (N_2411,N_2247,N_2371);
or U2412 (N_2412,N_2231,N_2308);
or U2413 (N_2413,N_2203,N_2291);
and U2414 (N_2414,N_2278,N_2248);
nor U2415 (N_2415,N_2254,N_2389);
nand U2416 (N_2416,N_2215,N_2353);
nand U2417 (N_2417,N_2363,N_2232);
nor U2418 (N_2418,N_2374,N_2208);
nor U2419 (N_2419,N_2301,N_2369);
or U2420 (N_2420,N_2314,N_2381);
nand U2421 (N_2421,N_2263,N_2241);
nand U2422 (N_2422,N_2223,N_2348);
nand U2423 (N_2423,N_2329,N_2334);
nand U2424 (N_2424,N_2216,N_2321);
nand U2425 (N_2425,N_2366,N_2265);
or U2426 (N_2426,N_2205,N_2243);
nor U2427 (N_2427,N_2391,N_2398);
nor U2428 (N_2428,N_2212,N_2325);
or U2429 (N_2429,N_2394,N_2396);
nor U2430 (N_2430,N_2349,N_2304);
nor U2431 (N_2431,N_2283,N_2260);
or U2432 (N_2432,N_2286,N_2282);
nand U2433 (N_2433,N_2399,N_2284);
nor U2434 (N_2434,N_2309,N_2395);
nor U2435 (N_2435,N_2289,N_2259);
or U2436 (N_2436,N_2327,N_2312);
nor U2437 (N_2437,N_2382,N_2279);
and U2438 (N_2438,N_2272,N_2201);
or U2439 (N_2439,N_2288,N_2373);
nor U2440 (N_2440,N_2214,N_2356);
nor U2441 (N_2441,N_2253,N_2204);
or U2442 (N_2442,N_2298,N_2306);
nor U2443 (N_2443,N_2235,N_2350);
nor U2444 (N_2444,N_2285,N_2220);
or U2445 (N_2445,N_2351,N_2352);
nor U2446 (N_2446,N_2287,N_2268);
and U2447 (N_2447,N_2386,N_2267);
and U2448 (N_2448,N_2237,N_2238);
or U2449 (N_2449,N_2339,N_2246);
or U2450 (N_2450,N_2269,N_2375);
or U2451 (N_2451,N_2388,N_2295);
and U2452 (N_2452,N_2347,N_2328);
nand U2453 (N_2453,N_2370,N_2311);
or U2454 (N_2454,N_2383,N_2317);
and U2455 (N_2455,N_2290,N_2310);
or U2456 (N_2456,N_2362,N_2315);
nand U2457 (N_2457,N_2392,N_2202);
nor U2458 (N_2458,N_2346,N_2207);
nand U2459 (N_2459,N_2227,N_2255);
nor U2460 (N_2460,N_2385,N_2274);
nand U2461 (N_2461,N_2320,N_2261);
nor U2462 (N_2462,N_2367,N_2234);
nand U2463 (N_2463,N_2357,N_2313);
or U2464 (N_2464,N_2275,N_2377);
xnor U2465 (N_2465,N_2249,N_2262);
or U2466 (N_2466,N_2376,N_2222);
nand U2467 (N_2467,N_2257,N_2323);
nand U2468 (N_2468,N_2305,N_2343);
nand U2469 (N_2469,N_2354,N_2236);
nor U2470 (N_2470,N_2322,N_2359);
nand U2471 (N_2471,N_2210,N_2302);
nor U2472 (N_2472,N_2358,N_2258);
nand U2473 (N_2473,N_2245,N_2206);
nor U2474 (N_2474,N_2387,N_2276);
or U2475 (N_2475,N_2344,N_2380);
or U2476 (N_2476,N_2273,N_2264);
or U2477 (N_2477,N_2378,N_2224);
or U2478 (N_2478,N_2336,N_2200);
or U2479 (N_2479,N_2307,N_2303);
nand U2480 (N_2480,N_2230,N_2316);
and U2481 (N_2481,N_2221,N_2219);
or U2482 (N_2482,N_2393,N_2280);
nor U2483 (N_2483,N_2252,N_2333);
xnor U2484 (N_2484,N_2211,N_2337);
nor U2485 (N_2485,N_2226,N_2213);
nand U2486 (N_2486,N_2364,N_2330);
and U2487 (N_2487,N_2218,N_2240);
and U2488 (N_2488,N_2355,N_2319);
nand U2489 (N_2489,N_2318,N_2361);
nand U2490 (N_2490,N_2335,N_2341);
nor U2491 (N_2491,N_2338,N_2296);
nand U2492 (N_2492,N_2250,N_2324);
or U2493 (N_2493,N_2242,N_2379);
nand U2494 (N_2494,N_2332,N_2293);
and U2495 (N_2495,N_2294,N_2256);
nor U2496 (N_2496,N_2217,N_2270);
or U2497 (N_2497,N_2228,N_2292);
nor U2498 (N_2498,N_2251,N_2300);
or U2499 (N_2499,N_2244,N_2365);
or U2500 (N_2500,N_2276,N_2220);
nor U2501 (N_2501,N_2239,N_2338);
nor U2502 (N_2502,N_2290,N_2259);
nor U2503 (N_2503,N_2285,N_2294);
or U2504 (N_2504,N_2251,N_2345);
nand U2505 (N_2505,N_2290,N_2215);
and U2506 (N_2506,N_2276,N_2200);
nor U2507 (N_2507,N_2278,N_2221);
nor U2508 (N_2508,N_2384,N_2370);
nand U2509 (N_2509,N_2246,N_2320);
nor U2510 (N_2510,N_2248,N_2344);
or U2511 (N_2511,N_2299,N_2203);
and U2512 (N_2512,N_2241,N_2327);
nor U2513 (N_2513,N_2325,N_2299);
nand U2514 (N_2514,N_2282,N_2261);
or U2515 (N_2515,N_2359,N_2302);
or U2516 (N_2516,N_2250,N_2207);
nor U2517 (N_2517,N_2349,N_2374);
nand U2518 (N_2518,N_2399,N_2348);
nor U2519 (N_2519,N_2292,N_2340);
xnor U2520 (N_2520,N_2346,N_2201);
or U2521 (N_2521,N_2300,N_2379);
nor U2522 (N_2522,N_2214,N_2224);
and U2523 (N_2523,N_2284,N_2216);
or U2524 (N_2524,N_2326,N_2344);
nor U2525 (N_2525,N_2231,N_2344);
nor U2526 (N_2526,N_2224,N_2390);
or U2527 (N_2527,N_2325,N_2351);
and U2528 (N_2528,N_2375,N_2274);
or U2529 (N_2529,N_2315,N_2281);
and U2530 (N_2530,N_2341,N_2392);
nor U2531 (N_2531,N_2328,N_2340);
and U2532 (N_2532,N_2373,N_2255);
nand U2533 (N_2533,N_2276,N_2368);
nand U2534 (N_2534,N_2331,N_2320);
and U2535 (N_2535,N_2311,N_2278);
nor U2536 (N_2536,N_2382,N_2295);
and U2537 (N_2537,N_2282,N_2215);
nand U2538 (N_2538,N_2311,N_2390);
nand U2539 (N_2539,N_2252,N_2308);
and U2540 (N_2540,N_2338,N_2373);
and U2541 (N_2541,N_2398,N_2281);
nand U2542 (N_2542,N_2263,N_2361);
or U2543 (N_2543,N_2295,N_2350);
nor U2544 (N_2544,N_2226,N_2239);
or U2545 (N_2545,N_2340,N_2251);
or U2546 (N_2546,N_2331,N_2288);
and U2547 (N_2547,N_2215,N_2249);
nand U2548 (N_2548,N_2395,N_2385);
and U2549 (N_2549,N_2373,N_2319);
nor U2550 (N_2550,N_2225,N_2267);
nand U2551 (N_2551,N_2231,N_2311);
or U2552 (N_2552,N_2209,N_2392);
and U2553 (N_2553,N_2214,N_2319);
and U2554 (N_2554,N_2286,N_2226);
and U2555 (N_2555,N_2358,N_2333);
nor U2556 (N_2556,N_2214,N_2337);
or U2557 (N_2557,N_2238,N_2394);
and U2558 (N_2558,N_2293,N_2247);
nand U2559 (N_2559,N_2331,N_2363);
nor U2560 (N_2560,N_2392,N_2380);
and U2561 (N_2561,N_2219,N_2396);
nand U2562 (N_2562,N_2290,N_2292);
nand U2563 (N_2563,N_2321,N_2376);
nor U2564 (N_2564,N_2213,N_2216);
nand U2565 (N_2565,N_2399,N_2286);
nor U2566 (N_2566,N_2205,N_2240);
and U2567 (N_2567,N_2246,N_2305);
and U2568 (N_2568,N_2314,N_2322);
and U2569 (N_2569,N_2244,N_2223);
nand U2570 (N_2570,N_2259,N_2268);
nand U2571 (N_2571,N_2211,N_2315);
nand U2572 (N_2572,N_2343,N_2312);
nand U2573 (N_2573,N_2278,N_2379);
nor U2574 (N_2574,N_2223,N_2294);
nand U2575 (N_2575,N_2239,N_2297);
or U2576 (N_2576,N_2312,N_2378);
and U2577 (N_2577,N_2212,N_2391);
nor U2578 (N_2578,N_2252,N_2339);
nand U2579 (N_2579,N_2303,N_2355);
nor U2580 (N_2580,N_2369,N_2381);
or U2581 (N_2581,N_2374,N_2318);
or U2582 (N_2582,N_2264,N_2364);
nor U2583 (N_2583,N_2210,N_2351);
nor U2584 (N_2584,N_2261,N_2251);
or U2585 (N_2585,N_2398,N_2289);
and U2586 (N_2586,N_2249,N_2368);
and U2587 (N_2587,N_2354,N_2275);
and U2588 (N_2588,N_2326,N_2257);
nand U2589 (N_2589,N_2291,N_2273);
xnor U2590 (N_2590,N_2267,N_2218);
or U2591 (N_2591,N_2389,N_2363);
or U2592 (N_2592,N_2397,N_2321);
and U2593 (N_2593,N_2239,N_2255);
or U2594 (N_2594,N_2379,N_2282);
and U2595 (N_2595,N_2247,N_2380);
nor U2596 (N_2596,N_2277,N_2379);
nand U2597 (N_2597,N_2333,N_2212);
and U2598 (N_2598,N_2338,N_2230);
nor U2599 (N_2599,N_2262,N_2319);
nor U2600 (N_2600,N_2578,N_2554);
or U2601 (N_2601,N_2401,N_2425);
and U2602 (N_2602,N_2552,N_2457);
nor U2603 (N_2603,N_2531,N_2557);
nor U2604 (N_2604,N_2451,N_2454);
nor U2605 (N_2605,N_2414,N_2495);
nand U2606 (N_2606,N_2408,N_2573);
or U2607 (N_2607,N_2527,N_2585);
and U2608 (N_2608,N_2506,N_2536);
or U2609 (N_2609,N_2515,N_2511);
nand U2610 (N_2610,N_2418,N_2519);
and U2611 (N_2611,N_2522,N_2470);
nor U2612 (N_2612,N_2491,N_2586);
nor U2613 (N_2613,N_2464,N_2494);
and U2614 (N_2614,N_2526,N_2404);
and U2615 (N_2615,N_2503,N_2444);
nor U2616 (N_2616,N_2489,N_2547);
nor U2617 (N_2617,N_2566,N_2529);
nand U2618 (N_2618,N_2535,N_2540);
and U2619 (N_2619,N_2591,N_2570);
nand U2620 (N_2620,N_2471,N_2400);
nand U2621 (N_2621,N_2473,N_2508);
nand U2622 (N_2622,N_2475,N_2423);
and U2623 (N_2623,N_2550,N_2556);
nor U2624 (N_2624,N_2460,N_2448);
nor U2625 (N_2625,N_2525,N_2458);
xor U2626 (N_2626,N_2504,N_2434);
or U2627 (N_2627,N_2483,N_2590);
nor U2628 (N_2628,N_2545,N_2539);
and U2629 (N_2629,N_2598,N_2538);
nor U2630 (N_2630,N_2524,N_2509);
nand U2631 (N_2631,N_2426,N_2542);
or U2632 (N_2632,N_2594,N_2463);
or U2633 (N_2633,N_2592,N_2498);
or U2634 (N_2634,N_2450,N_2493);
nand U2635 (N_2635,N_2518,N_2419);
and U2636 (N_2636,N_2486,N_2572);
nand U2637 (N_2637,N_2429,N_2565);
and U2638 (N_2638,N_2459,N_2422);
nand U2639 (N_2639,N_2530,N_2569);
and U2640 (N_2640,N_2523,N_2580);
and U2641 (N_2641,N_2582,N_2480);
nand U2642 (N_2642,N_2555,N_2497);
nor U2643 (N_2643,N_2479,N_2558);
nor U2644 (N_2644,N_2517,N_2412);
and U2645 (N_2645,N_2577,N_2544);
or U2646 (N_2646,N_2443,N_2501);
or U2647 (N_2647,N_2561,N_2512);
nand U2648 (N_2648,N_2488,N_2467);
nor U2649 (N_2649,N_2462,N_2417);
and U2650 (N_2650,N_2532,N_2560);
or U2651 (N_2651,N_2553,N_2407);
or U2652 (N_2652,N_2430,N_2469);
or U2653 (N_2653,N_2563,N_2411);
or U2654 (N_2654,N_2507,N_2571);
xnor U2655 (N_2655,N_2514,N_2421);
nand U2656 (N_2656,N_2496,N_2499);
nand U2657 (N_2657,N_2445,N_2477);
xor U2658 (N_2658,N_2431,N_2505);
nand U2659 (N_2659,N_2437,N_2597);
or U2660 (N_2660,N_2564,N_2482);
nand U2661 (N_2661,N_2438,N_2510);
nand U2662 (N_2662,N_2428,N_2435);
or U2663 (N_2663,N_2520,N_2551);
and U2664 (N_2664,N_2452,N_2568);
and U2665 (N_2665,N_2490,N_2413);
and U2666 (N_2666,N_2567,N_2456);
nand U2667 (N_2667,N_2574,N_2581);
nor U2668 (N_2668,N_2593,N_2521);
nor U2669 (N_2669,N_2442,N_2472);
and U2670 (N_2670,N_2576,N_2583);
or U2671 (N_2671,N_2453,N_2466);
or U2672 (N_2672,N_2546,N_2405);
nor U2673 (N_2673,N_2402,N_2433);
nor U2674 (N_2674,N_2549,N_2432);
or U2675 (N_2675,N_2492,N_2579);
or U2676 (N_2676,N_2589,N_2409);
nand U2677 (N_2677,N_2502,N_2485);
nor U2678 (N_2678,N_2500,N_2416);
and U2679 (N_2679,N_2587,N_2588);
nand U2680 (N_2680,N_2533,N_2534);
nand U2681 (N_2681,N_2455,N_2562);
or U2682 (N_2682,N_2487,N_2449);
or U2683 (N_2683,N_2446,N_2575);
and U2684 (N_2684,N_2420,N_2541);
or U2685 (N_2685,N_2595,N_2427);
nand U2686 (N_2686,N_2403,N_2584);
nor U2687 (N_2687,N_2415,N_2599);
and U2688 (N_2688,N_2440,N_2406);
and U2689 (N_2689,N_2447,N_2410);
or U2690 (N_2690,N_2424,N_2528);
nand U2691 (N_2691,N_2548,N_2436);
or U2692 (N_2692,N_2537,N_2441);
nor U2693 (N_2693,N_2474,N_2465);
or U2694 (N_2694,N_2516,N_2513);
nor U2695 (N_2695,N_2478,N_2481);
or U2696 (N_2696,N_2543,N_2476);
nand U2697 (N_2697,N_2461,N_2596);
nand U2698 (N_2698,N_2484,N_2439);
nor U2699 (N_2699,N_2559,N_2468);
nor U2700 (N_2700,N_2510,N_2561);
nand U2701 (N_2701,N_2587,N_2565);
nor U2702 (N_2702,N_2589,N_2531);
and U2703 (N_2703,N_2526,N_2531);
nand U2704 (N_2704,N_2426,N_2517);
nor U2705 (N_2705,N_2440,N_2584);
nor U2706 (N_2706,N_2411,N_2559);
nand U2707 (N_2707,N_2588,N_2582);
nor U2708 (N_2708,N_2465,N_2562);
nand U2709 (N_2709,N_2424,N_2549);
and U2710 (N_2710,N_2514,N_2403);
nand U2711 (N_2711,N_2450,N_2542);
or U2712 (N_2712,N_2461,N_2415);
nor U2713 (N_2713,N_2449,N_2431);
or U2714 (N_2714,N_2462,N_2588);
nor U2715 (N_2715,N_2404,N_2562);
and U2716 (N_2716,N_2492,N_2408);
and U2717 (N_2717,N_2585,N_2557);
nand U2718 (N_2718,N_2584,N_2516);
or U2719 (N_2719,N_2406,N_2479);
nor U2720 (N_2720,N_2411,N_2556);
or U2721 (N_2721,N_2429,N_2477);
or U2722 (N_2722,N_2529,N_2520);
and U2723 (N_2723,N_2500,N_2493);
nand U2724 (N_2724,N_2499,N_2560);
nor U2725 (N_2725,N_2474,N_2539);
nand U2726 (N_2726,N_2588,N_2520);
and U2727 (N_2727,N_2406,N_2482);
or U2728 (N_2728,N_2513,N_2405);
nand U2729 (N_2729,N_2546,N_2416);
nand U2730 (N_2730,N_2516,N_2504);
and U2731 (N_2731,N_2563,N_2567);
xnor U2732 (N_2732,N_2467,N_2453);
nand U2733 (N_2733,N_2552,N_2401);
nand U2734 (N_2734,N_2402,N_2449);
and U2735 (N_2735,N_2443,N_2402);
nor U2736 (N_2736,N_2581,N_2584);
nor U2737 (N_2737,N_2581,N_2547);
and U2738 (N_2738,N_2578,N_2599);
nand U2739 (N_2739,N_2540,N_2555);
nand U2740 (N_2740,N_2583,N_2574);
or U2741 (N_2741,N_2447,N_2580);
or U2742 (N_2742,N_2423,N_2477);
nor U2743 (N_2743,N_2403,N_2597);
or U2744 (N_2744,N_2493,N_2522);
or U2745 (N_2745,N_2411,N_2506);
and U2746 (N_2746,N_2464,N_2448);
nand U2747 (N_2747,N_2457,N_2526);
nand U2748 (N_2748,N_2430,N_2592);
or U2749 (N_2749,N_2528,N_2513);
xor U2750 (N_2750,N_2511,N_2493);
and U2751 (N_2751,N_2447,N_2438);
and U2752 (N_2752,N_2419,N_2467);
or U2753 (N_2753,N_2528,N_2558);
and U2754 (N_2754,N_2489,N_2473);
nor U2755 (N_2755,N_2485,N_2493);
and U2756 (N_2756,N_2439,N_2465);
and U2757 (N_2757,N_2560,N_2403);
nor U2758 (N_2758,N_2455,N_2563);
or U2759 (N_2759,N_2556,N_2440);
or U2760 (N_2760,N_2577,N_2454);
and U2761 (N_2761,N_2411,N_2486);
nand U2762 (N_2762,N_2553,N_2531);
nor U2763 (N_2763,N_2572,N_2439);
and U2764 (N_2764,N_2561,N_2489);
or U2765 (N_2765,N_2523,N_2517);
or U2766 (N_2766,N_2504,N_2486);
or U2767 (N_2767,N_2512,N_2586);
or U2768 (N_2768,N_2462,N_2472);
and U2769 (N_2769,N_2475,N_2590);
and U2770 (N_2770,N_2499,N_2504);
or U2771 (N_2771,N_2456,N_2501);
or U2772 (N_2772,N_2539,N_2521);
or U2773 (N_2773,N_2526,N_2494);
and U2774 (N_2774,N_2563,N_2550);
nor U2775 (N_2775,N_2535,N_2525);
or U2776 (N_2776,N_2529,N_2435);
and U2777 (N_2777,N_2410,N_2441);
nand U2778 (N_2778,N_2567,N_2552);
xnor U2779 (N_2779,N_2560,N_2468);
nor U2780 (N_2780,N_2464,N_2546);
nor U2781 (N_2781,N_2486,N_2402);
nand U2782 (N_2782,N_2518,N_2566);
nand U2783 (N_2783,N_2503,N_2415);
and U2784 (N_2784,N_2557,N_2415);
and U2785 (N_2785,N_2571,N_2428);
or U2786 (N_2786,N_2416,N_2497);
nand U2787 (N_2787,N_2474,N_2457);
or U2788 (N_2788,N_2574,N_2431);
nor U2789 (N_2789,N_2526,N_2429);
nand U2790 (N_2790,N_2585,N_2551);
and U2791 (N_2791,N_2414,N_2598);
nor U2792 (N_2792,N_2527,N_2553);
or U2793 (N_2793,N_2552,N_2581);
or U2794 (N_2794,N_2445,N_2588);
or U2795 (N_2795,N_2550,N_2529);
and U2796 (N_2796,N_2531,N_2570);
nor U2797 (N_2797,N_2411,N_2455);
and U2798 (N_2798,N_2560,N_2446);
nand U2799 (N_2799,N_2542,N_2452);
nor U2800 (N_2800,N_2726,N_2722);
nand U2801 (N_2801,N_2641,N_2648);
or U2802 (N_2802,N_2606,N_2600);
and U2803 (N_2803,N_2655,N_2786);
or U2804 (N_2804,N_2628,N_2669);
nand U2805 (N_2805,N_2728,N_2663);
and U2806 (N_2806,N_2686,N_2601);
nand U2807 (N_2807,N_2671,N_2721);
nor U2808 (N_2808,N_2703,N_2610);
nor U2809 (N_2809,N_2715,N_2675);
and U2810 (N_2810,N_2734,N_2690);
nor U2811 (N_2811,N_2615,N_2616);
nor U2812 (N_2812,N_2749,N_2634);
nor U2813 (N_2813,N_2602,N_2797);
nand U2814 (N_2814,N_2798,N_2767);
xnor U2815 (N_2815,N_2765,N_2658);
nor U2816 (N_2816,N_2691,N_2605);
nor U2817 (N_2817,N_2753,N_2617);
and U2818 (N_2818,N_2704,N_2632);
xor U2819 (N_2819,N_2707,N_2727);
nand U2820 (N_2820,N_2699,N_2619);
and U2821 (N_2821,N_2621,N_2693);
nand U2822 (N_2822,N_2756,N_2731);
and U2823 (N_2823,N_2656,N_2766);
nor U2824 (N_2824,N_2687,N_2636);
or U2825 (N_2825,N_2633,N_2740);
nor U2826 (N_2826,N_2739,N_2737);
or U2827 (N_2827,N_2657,N_2670);
nor U2828 (N_2828,N_2682,N_2735);
nor U2829 (N_2829,N_2757,N_2781);
nor U2830 (N_2830,N_2794,N_2762);
or U2831 (N_2831,N_2697,N_2775);
nand U2832 (N_2832,N_2607,N_2709);
and U2833 (N_2833,N_2755,N_2776);
or U2834 (N_2834,N_2647,N_2666);
and U2835 (N_2835,N_2646,N_2723);
or U2836 (N_2836,N_2629,N_2718);
nor U2837 (N_2837,N_2638,N_2623);
or U2838 (N_2838,N_2788,N_2660);
nand U2839 (N_2839,N_2613,N_2712);
and U2840 (N_2840,N_2680,N_2787);
xor U2841 (N_2841,N_2716,N_2685);
or U2842 (N_2842,N_2732,N_2618);
or U2843 (N_2843,N_2791,N_2665);
nor U2844 (N_2844,N_2729,N_2745);
nor U2845 (N_2845,N_2758,N_2688);
or U2846 (N_2846,N_2612,N_2741);
nor U2847 (N_2847,N_2770,N_2695);
nor U2848 (N_2848,N_2789,N_2692);
and U2849 (N_2849,N_2662,N_2677);
or U2850 (N_2850,N_2780,N_2730);
nor U2851 (N_2851,N_2774,N_2667);
or U2852 (N_2852,N_2604,N_2706);
nor U2853 (N_2853,N_2661,N_2635);
and U2854 (N_2854,N_2696,N_2773);
nand U2855 (N_2855,N_2694,N_2637);
nor U2856 (N_2856,N_2724,N_2751);
nand U2857 (N_2857,N_2793,N_2783);
and U2858 (N_2858,N_2701,N_2627);
nor U2859 (N_2859,N_2748,N_2674);
and U2860 (N_2860,N_2684,N_2673);
and U2861 (N_2861,N_2733,N_2799);
nor U2862 (N_2862,N_2643,N_2796);
nor U2863 (N_2863,N_2654,N_2760);
nand U2864 (N_2864,N_2652,N_2764);
or U2865 (N_2865,N_2743,N_2644);
or U2866 (N_2866,N_2746,N_2603);
nor U2867 (N_2867,N_2676,N_2744);
nand U2868 (N_2868,N_2725,N_2705);
nand U2869 (N_2869,N_2790,N_2747);
and U2870 (N_2870,N_2681,N_2768);
nand U2871 (N_2871,N_2710,N_2763);
nor U2872 (N_2872,N_2719,N_2738);
nand U2873 (N_2873,N_2678,N_2711);
nor U2874 (N_2874,N_2717,N_2700);
or U2875 (N_2875,N_2750,N_2713);
and U2876 (N_2876,N_2625,N_2708);
or U2877 (N_2877,N_2668,N_2650);
nand U2878 (N_2878,N_2720,N_2614);
or U2879 (N_2879,N_2626,N_2645);
or U2880 (N_2880,N_2777,N_2651);
and U2881 (N_2881,N_2611,N_2642);
nor U2882 (N_2882,N_2759,N_2653);
nand U2883 (N_2883,N_2778,N_2698);
and U2884 (N_2884,N_2784,N_2792);
nand U2885 (N_2885,N_2624,N_2782);
or U2886 (N_2886,N_2702,N_2761);
and U2887 (N_2887,N_2754,N_2622);
nand U2888 (N_2888,N_2736,N_2672);
and U2889 (N_2889,N_2608,N_2630);
and U2890 (N_2890,N_2640,N_2769);
and U2891 (N_2891,N_2779,N_2664);
nand U2892 (N_2892,N_2771,N_2649);
nor U2893 (N_2893,N_2609,N_2639);
nand U2894 (N_2894,N_2772,N_2683);
nand U2895 (N_2895,N_2752,N_2659);
and U2896 (N_2896,N_2689,N_2714);
and U2897 (N_2897,N_2742,N_2785);
and U2898 (N_2898,N_2795,N_2679);
nor U2899 (N_2899,N_2620,N_2631);
nand U2900 (N_2900,N_2677,N_2798);
or U2901 (N_2901,N_2605,N_2671);
nor U2902 (N_2902,N_2767,N_2708);
and U2903 (N_2903,N_2773,N_2759);
and U2904 (N_2904,N_2603,N_2706);
or U2905 (N_2905,N_2670,N_2789);
and U2906 (N_2906,N_2684,N_2631);
nand U2907 (N_2907,N_2751,N_2661);
nor U2908 (N_2908,N_2751,N_2647);
nand U2909 (N_2909,N_2773,N_2796);
nand U2910 (N_2910,N_2770,N_2709);
and U2911 (N_2911,N_2713,N_2670);
nor U2912 (N_2912,N_2779,N_2631);
nor U2913 (N_2913,N_2652,N_2673);
nor U2914 (N_2914,N_2603,N_2749);
or U2915 (N_2915,N_2779,N_2606);
nor U2916 (N_2916,N_2792,N_2695);
and U2917 (N_2917,N_2690,N_2682);
and U2918 (N_2918,N_2665,N_2778);
or U2919 (N_2919,N_2753,N_2782);
and U2920 (N_2920,N_2778,N_2743);
or U2921 (N_2921,N_2779,N_2653);
or U2922 (N_2922,N_2714,N_2608);
or U2923 (N_2923,N_2696,N_2791);
or U2924 (N_2924,N_2621,N_2689);
and U2925 (N_2925,N_2714,N_2668);
or U2926 (N_2926,N_2731,N_2683);
or U2927 (N_2927,N_2615,N_2607);
nor U2928 (N_2928,N_2747,N_2674);
nand U2929 (N_2929,N_2632,N_2795);
nor U2930 (N_2930,N_2693,N_2799);
or U2931 (N_2931,N_2636,N_2643);
nor U2932 (N_2932,N_2600,N_2706);
and U2933 (N_2933,N_2701,N_2736);
nand U2934 (N_2934,N_2709,N_2744);
nand U2935 (N_2935,N_2705,N_2746);
nor U2936 (N_2936,N_2656,N_2672);
and U2937 (N_2937,N_2688,N_2722);
nand U2938 (N_2938,N_2659,N_2645);
nand U2939 (N_2939,N_2714,N_2655);
nand U2940 (N_2940,N_2765,N_2681);
or U2941 (N_2941,N_2649,N_2759);
xor U2942 (N_2942,N_2730,N_2744);
nand U2943 (N_2943,N_2628,N_2720);
or U2944 (N_2944,N_2744,N_2722);
nand U2945 (N_2945,N_2747,N_2769);
nor U2946 (N_2946,N_2604,N_2689);
nor U2947 (N_2947,N_2732,N_2738);
or U2948 (N_2948,N_2741,N_2786);
and U2949 (N_2949,N_2606,N_2626);
nor U2950 (N_2950,N_2663,N_2737);
nand U2951 (N_2951,N_2601,N_2616);
nand U2952 (N_2952,N_2653,N_2755);
or U2953 (N_2953,N_2751,N_2656);
nand U2954 (N_2954,N_2602,N_2697);
nand U2955 (N_2955,N_2633,N_2732);
and U2956 (N_2956,N_2707,N_2750);
nor U2957 (N_2957,N_2683,N_2642);
and U2958 (N_2958,N_2623,N_2603);
nand U2959 (N_2959,N_2792,N_2682);
or U2960 (N_2960,N_2619,N_2684);
nand U2961 (N_2961,N_2709,N_2758);
nor U2962 (N_2962,N_2725,N_2620);
and U2963 (N_2963,N_2740,N_2770);
or U2964 (N_2964,N_2604,N_2753);
nor U2965 (N_2965,N_2606,N_2716);
and U2966 (N_2966,N_2704,N_2730);
nor U2967 (N_2967,N_2722,N_2794);
nand U2968 (N_2968,N_2666,N_2706);
or U2969 (N_2969,N_2604,N_2768);
and U2970 (N_2970,N_2717,N_2669);
nand U2971 (N_2971,N_2746,N_2654);
nor U2972 (N_2972,N_2701,N_2726);
and U2973 (N_2973,N_2682,N_2731);
or U2974 (N_2974,N_2617,N_2635);
or U2975 (N_2975,N_2690,N_2793);
nand U2976 (N_2976,N_2732,N_2756);
nor U2977 (N_2977,N_2756,N_2766);
nor U2978 (N_2978,N_2679,N_2700);
nor U2979 (N_2979,N_2767,N_2648);
nand U2980 (N_2980,N_2624,N_2668);
and U2981 (N_2981,N_2764,N_2706);
or U2982 (N_2982,N_2770,N_2604);
and U2983 (N_2983,N_2689,N_2653);
and U2984 (N_2984,N_2671,N_2711);
and U2985 (N_2985,N_2679,N_2633);
nor U2986 (N_2986,N_2652,N_2688);
nor U2987 (N_2987,N_2759,N_2752);
nand U2988 (N_2988,N_2659,N_2639);
nand U2989 (N_2989,N_2600,N_2748);
nor U2990 (N_2990,N_2632,N_2620);
and U2991 (N_2991,N_2664,N_2634);
nor U2992 (N_2992,N_2737,N_2728);
nor U2993 (N_2993,N_2631,N_2703);
or U2994 (N_2994,N_2606,N_2741);
or U2995 (N_2995,N_2673,N_2729);
nor U2996 (N_2996,N_2768,N_2642);
and U2997 (N_2997,N_2601,N_2794);
or U2998 (N_2998,N_2659,N_2722);
nor U2999 (N_2999,N_2795,N_2762);
or U3000 (N_3000,N_2840,N_2969);
or U3001 (N_3001,N_2846,N_2916);
nand U3002 (N_3002,N_2985,N_2866);
nor U3003 (N_3003,N_2820,N_2815);
nand U3004 (N_3004,N_2946,N_2897);
or U3005 (N_3005,N_2800,N_2943);
nor U3006 (N_3006,N_2966,N_2944);
or U3007 (N_3007,N_2808,N_2886);
and U3008 (N_3008,N_2898,N_2930);
nand U3009 (N_3009,N_2842,N_2857);
nand U3010 (N_3010,N_2814,N_2903);
nor U3011 (N_3011,N_2813,N_2981);
nor U3012 (N_3012,N_2934,N_2852);
and U3013 (N_3013,N_2810,N_2821);
nor U3014 (N_3014,N_2957,N_2988);
or U3015 (N_3015,N_2913,N_2824);
or U3016 (N_3016,N_2950,N_2952);
or U3017 (N_3017,N_2933,N_2971);
or U3018 (N_3018,N_2882,N_2830);
and U3019 (N_3019,N_2805,N_2844);
or U3020 (N_3020,N_2883,N_2975);
nor U3021 (N_3021,N_2861,N_2851);
nand U3022 (N_3022,N_2826,N_2809);
or U3023 (N_3023,N_2847,N_2899);
nand U3024 (N_3024,N_2850,N_2907);
and U3025 (N_3025,N_2807,N_2864);
and U3026 (N_3026,N_2994,N_2843);
nand U3027 (N_3027,N_2995,N_2962);
or U3028 (N_3028,N_2993,N_2875);
nand U3029 (N_3029,N_2858,N_2827);
nand U3030 (N_3030,N_2926,N_2914);
nor U3031 (N_3031,N_2972,N_2856);
or U3032 (N_3032,N_2910,N_2928);
nand U3033 (N_3033,N_2859,N_2956);
nor U3034 (N_3034,N_2837,N_2876);
or U3035 (N_3035,N_2991,N_2902);
nand U3036 (N_3036,N_2999,N_2948);
nand U3037 (N_3037,N_2881,N_2869);
nand U3038 (N_3038,N_2941,N_2855);
nand U3039 (N_3039,N_2945,N_2803);
and U3040 (N_3040,N_2970,N_2990);
nor U3041 (N_3041,N_2929,N_2890);
nand U3042 (N_3042,N_2908,N_2983);
nand U3043 (N_3043,N_2887,N_2918);
nor U3044 (N_3044,N_2996,N_2839);
nand U3045 (N_3045,N_2968,N_2959);
or U3046 (N_3046,N_2801,N_2901);
nand U3047 (N_3047,N_2925,N_2920);
and U3048 (N_3048,N_2896,N_2838);
nand U3049 (N_3049,N_2989,N_2919);
nand U3050 (N_3050,N_2848,N_2997);
or U3051 (N_3051,N_2818,N_2817);
nor U3052 (N_3052,N_2963,N_2806);
nor U3053 (N_3053,N_2937,N_2804);
nand U3054 (N_3054,N_2885,N_2947);
nor U3055 (N_3055,N_2825,N_2878);
nand U3056 (N_3056,N_2854,N_2976);
nand U3057 (N_3057,N_2822,N_2833);
nand U3058 (N_3058,N_2949,N_2845);
nand U3059 (N_3059,N_2982,N_2924);
nand U3060 (N_3060,N_2960,N_2867);
or U3061 (N_3061,N_2936,N_2849);
and U3062 (N_3062,N_2961,N_2954);
nor U3063 (N_3063,N_2880,N_2965);
or U3064 (N_3064,N_2868,N_2905);
nor U3065 (N_3065,N_2888,N_2955);
nand U3066 (N_3066,N_2835,N_2874);
nand U3067 (N_3067,N_2992,N_2853);
and U3068 (N_3068,N_2832,N_2931);
or U3069 (N_3069,N_2980,N_2823);
nor U3070 (N_3070,N_2872,N_2877);
nor U3071 (N_3071,N_2841,N_2974);
nor U3072 (N_3072,N_2900,N_2938);
nand U3073 (N_3073,N_2860,N_2889);
nor U3074 (N_3074,N_2923,N_2942);
or U3075 (N_3075,N_2984,N_2921);
nand U3076 (N_3076,N_2979,N_2953);
and U3077 (N_3077,N_2893,N_2951);
nor U3078 (N_3078,N_2879,N_2964);
or U3079 (N_3079,N_2927,N_2935);
or U3080 (N_3080,N_2819,N_2973);
and U3081 (N_3081,N_2894,N_2831);
nor U3082 (N_3082,N_2836,N_2884);
nor U3083 (N_3083,N_2986,N_2998);
or U3084 (N_3084,N_2828,N_2863);
and U3085 (N_3085,N_2811,N_2940);
nand U3086 (N_3086,N_2816,N_2906);
or U3087 (N_3087,N_2939,N_2909);
nor U3088 (N_3088,N_2862,N_2891);
or U3089 (N_3089,N_2917,N_2912);
and U3090 (N_3090,N_2865,N_2978);
and U3091 (N_3091,N_2802,N_2829);
and U3092 (N_3092,N_2922,N_2834);
or U3093 (N_3093,N_2892,N_2904);
or U3094 (N_3094,N_2932,N_2911);
or U3095 (N_3095,N_2915,N_2958);
and U3096 (N_3096,N_2873,N_2812);
nor U3097 (N_3097,N_2870,N_2895);
nand U3098 (N_3098,N_2871,N_2967);
nor U3099 (N_3099,N_2987,N_2977);
or U3100 (N_3100,N_2881,N_2833);
and U3101 (N_3101,N_2812,N_2965);
nor U3102 (N_3102,N_2945,N_2806);
xor U3103 (N_3103,N_2831,N_2879);
and U3104 (N_3104,N_2958,N_2949);
nand U3105 (N_3105,N_2921,N_2935);
and U3106 (N_3106,N_2842,N_2885);
and U3107 (N_3107,N_2881,N_2987);
xor U3108 (N_3108,N_2846,N_2879);
nor U3109 (N_3109,N_2965,N_2841);
and U3110 (N_3110,N_2956,N_2908);
or U3111 (N_3111,N_2888,N_2889);
nand U3112 (N_3112,N_2851,N_2847);
or U3113 (N_3113,N_2917,N_2972);
or U3114 (N_3114,N_2922,N_2868);
or U3115 (N_3115,N_2848,N_2873);
or U3116 (N_3116,N_2976,N_2856);
and U3117 (N_3117,N_2849,N_2894);
or U3118 (N_3118,N_2806,N_2903);
nand U3119 (N_3119,N_2919,N_2810);
nor U3120 (N_3120,N_2880,N_2887);
nor U3121 (N_3121,N_2863,N_2860);
nor U3122 (N_3122,N_2807,N_2804);
nand U3123 (N_3123,N_2938,N_2940);
or U3124 (N_3124,N_2869,N_2882);
or U3125 (N_3125,N_2839,N_2943);
nor U3126 (N_3126,N_2817,N_2913);
nor U3127 (N_3127,N_2896,N_2991);
and U3128 (N_3128,N_2852,N_2920);
or U3129 (N_3129,N_2933,N_2837);
nor U3130 (N_3130,N_2814,N_2882);
nor U3131 (N_3131,N_2935,N_2855);
nor U3132 (N_3132,N_2816,N_2883);
or U3133 (N_3133,N_2916,N_2900);
and U3134 (N_3134,N_2885,N_2849);
nand U3135 (N_3135,N_2971,N_2990);
and U3136 (N_3136,N_2804,N_2967);
nor U3137 (N_3137,N_2810,N_2901);
nor U3138 (N_3138,N_2842,N_2932);
nand U3139 (N_3139,N_2828,N_2852);
or U3140 (N_3140,N_2890,N_2909);
or U3141 (N_3141,N_2977,N_2994);
or U3142 (N_3142,N_2952,N_2859);
nor U3143 (N_3143,N_2859,N_2851);
nand U3144 (N_3144,N_2904,N_2821);
or U3145 (N_3145,N_2860,N_2942);
nand U3146 (N_3146,N_2846,N_2874);
or U3147 (N_3147,N_2921,N_2805);
or U3148 (N_3148,N_2894,N_2886);
or U3149 (N_3149,N_2804,N_2890);
or U3150 (N_3150,N_2806,N_2910);
or U3151 (N_3151,N_2946,N_2884);
nor U3152 (N_3152,N_2982,N_2909);
or U3153 (N_3153,N_2978,N_2919);
or U3154 (N_3154,N_2969,N_2936);
nor U3155 (N_3155,N_2925,N_2834);
nand U3156 (N_3156,N_2913,N_2844);
nor U3157 (N_3157,N_2846,N_2819);
or U3158 (N_3158,N_2959,N_2899);
nor U3159 (N_3159,N_2960,N_2915);
and U3160 (N_3160,N_2876,N_2971);
nand U3161 (N_3161,N_2887,N_2879);
and U3162 (N_3162,N_2987,N_2888);
nor U3163 (N_3163,N_2899,N_2935);
nand U3164 (N_3164,N_2913,N_2808);
nor U3165 (N_3165,N_2917,N_2811);
nand U3166 (N_3166,N_2975,N_2928);
or U3167 (N_3167,N_2883,N_2870);
nor U3168 (N_3168,N_2909,N_2831);
and U3169 (N_3169,N_2932,N_2933);
nand U3170 (N_3170,N_2838,N_2802);
or U3171 (N_3171,N_2857,N_2908);
nand U3172 (N_3172,N_2949,N_2976);
nor U3173 (N_3173,N_2948,N_2879);
nand U3174 (N_3174,N_2905,N_2965);
nand U3175 (N_3175,N_2987,N_2955);
nor U3176 (N_3176,N_2839,N_2908);
and U3177 (N_3177,N_2978,N_2931);
and U3178 (N_3178,N_2970,N_2934);
or U3179 (N_3179,N_2862,N_2985);
or U3180 (N_3180,N_2820,N_2955);
and U3181 (N_3181,N_2808,N_2989);
and U3182 (N_3182,N_2892,N_2977);
and U3183 (N_3183,N_2871,N_2964);
and U3184 (N_3184,N_2833,N_2967);
nand U3185 (N_3185,N_2826,N_2919);
or U3186 (N_3186,N_2903,N_2911);
nand U3187 (N_3187,N_2970,N_2993);
nand U3188 (N_3188,N_2998,N_2864);
nand U3189 (N_3189,N_2850,N_2820);
and U3190 (N_3190,N_2915,N_2846);
nand U3191 (N_3191,N_2967,N_2907);
nor U3192 (N_3192,N_2991,N_2818);
and U3193 (N_3193,N_2899,N_2870);
nand U3194 (N_3194,N_2956,N_2905);
and U3195 (N_3195,N_2935,N_2969);
nor U3196 (N_3196,N_2850,N_2834);
nor U3197 (N_3197,N_2874,N_2800);
and U3198 (N_3198,N_2948,N_2865);
and U3199 (N_3199,N_2828,N_2818);
and U3200 (N_3200,N_3139,N_3167);
xnor U3201 (N_3201,N_3136,N_3026);
nor U3202 (N_3202,N_3131,N_3092);
nor U3203 (N_3203,N_3186,N_3001);
xor U3204 (N_3204,N_3119,N_3076);
or U3205 (N_3205,N_3009,N_3081);
nor U3206 (N_3206,N_3097,N_3008);
and U3207 (N_3207,N_3163,N_3027);
nand U3208 (N_3208,N_3133,N_3109);
or U3209 (N_3209,N_3111,N_3180);
and U3210 (N_3210,N_3091,N_3166);
nand U3211 (N_3211,N_3158,N_3090);
nor U3212 (N_3212,N_3058,N_3066);
nor U3213 (N_3213,N_3054,N_3032);
nor U3214 (N_3214,N_3197,N_3036);
nor U3215 (N_3215,N_3017,N_3025);
or U3216 (N_3216,N_3022,N_3074);
and U3217 (N_3217,N_3103,N_3031);
and U3218 (N_3218,N_3077,N_3118);
or U3219 (N_3219,N_3037,N_3129);
nand U3220 (N_3220,N_3089,N_3095);
and U3221 (N_3221,N_3198,N_3101);
nand U3222 (N_3222,N_3137,N_3003);
nor U3223 (N_3223,N_3106,N_3080);
nor U3224 (N_3224,N_3142,N_3065);
or U3225 (N_3225,N_3178,N_3041);
or U3226 (N_3226,N_3038,N_3056);
and U3227 (N_3227,N_3039,N_3168);
nand U3228 (N_3228,N_3023,N_3173);
nor U3229 (N_3229,N_3086,N_3130);
nand U3230 (N_3230,N_3196,N_3110);
and U3231 (N_3231,N_3105,N_3070);
and U3232 (N_3232,N_3148,N_3064);
or U3233 (N_3233,N_3072,N_3071);
nand U3234 (N_3234,N_3159,N_3062);
or U3235 (N_3235,N_3011,N_3042);
nand U3236 (N_3236,N_3000,N_3108);
or U3237 (N_3237,N_3084,N_3012);
or U3238 (N_3238,N_3060,N_3195);
nand U3239 (N_3239,N_3147,N_3191);
or U3240 (N_3240,N_3132,N_3170);
nand U3241 (N_3241,N_3007,N_3115);
or U3242 (N_3242,N_3113,N_3185);
nor U3243 (N_3243,N_3184,N_3134);
or U3244 (N_3244,N_3154,N_3028);
or U3245 (N_3245,N_3157,N_3193);
or U3246 (N_3246,N_3061,N_3127);
xnor U3247 (N_3247,N_3015,N_3010);
or U3248 (N_3248,N_3112,N_3018);
or U3249 (N_3249,N_3045,N_3181);
or U3250 (N_3250,N_3050,N_3135);
and U3251 (N_3251,N_3047,N_3144);
nand U3252 (N_3252,N_3182,N_3016);
nor U3253 (N_3253,N_3052,N_3006);
or U3254 (N_3254,N_3151,N_3161);
and U3255 (N_3255,N_3165,N_3145);
or U3256 (N_3256,N_3035,N_3169);
or U3257 (N_3257,N_3073,N_3044);
nor U3258 (N_3258,N_3189,N_3153);
nand U3259 (N_3259,N_3059,N_3152);
nand U3260 (N_3260,N_3125,N_3120);
or U3261 (N_3261,N_3087,N_3083);
and U3262 (N_3262,N_3141,N_3005);
nand U3263 (N_3263,N_3075,N_3116);
and U3264 (N_3264,N_3063,N_3187);
nor U3265 (N_3265,N_3172,N_3069);
or U3266 (N_3266,N_3194,N_3099);
nand U3267 (N_3267,N_3094,N_3093);
nor U3268 (N_3268,N_3160,N_3190);
and U3269 (N_3269,N_3107,N_3174);
or U3270 (N_3270,N_3183,N_3146);
and U3271 (N_3271,N_3019,N_3171);
nand U3272 (N_3272,N_3102,N_3029);
and U3273 (N_3273,N_3155,N_3126);
nor U3274 (N_3274,N_3053,N_3088);
nor U3275 (N_3275,N_3024,N_3122);
nand U3276 (N_3276,N_3046,N_3175);
nor U3277 (N_3277,N_3096,N_3114);
nor U3278 (N_3278,N_3082,N_3079);
nand U3279 (N_3279,N_3098,N_3068);
and U3280 (N_3280,N_3140,N_3078);
and U3281 (N_3281,N_3021,N_3004);
nand U3282 (N_3282,N_3067,N_3055);
and U3283 (N_3283,N_3164,N_3043);
and U3284 (N_3284,N_3179,N_3104);
nor U3285 (N_3285,N_3143,N_3121);
and U3286 (N_3286,N_3034,N_3100);
or U3287 (N_3287,N_3057,N_3138);
nor U3288 (N_3288,N_3117,N_3123);
nand U3289 (N_3289,N_3048,N_3020);
or U3290 (N_3290,N_3014,N_3124);
nor U3291 (N_3291,N_3199,N_3051);
nand U3292 (N_3292,N_3156,N_3128);
or U3293 (N_3293,N_3030,N_3085);
and U3294 (N_3294,N_3149,N_3013);
nand U3295 (N_3295,N_3033,N_3049);
nand U3296 (N_3296,N_3002,N_3176);
and U3297 (N_3297,N_3192,N_3040);
and U3298 (N_3298,N_3150,N_3162);
nor U3299 (N_3299,N_3188,N_3177);
or U3300 (N_3300,N_3159,N_3064);
and U3301 (N_3301,N_3020,N_3085);
nor U3302 (N_3302,N_3010,N_3156);
nand U3303 (N_3303,N_3162,N_3041);
or U3304 (N_3304,N_3153,N_3185);
or U3305 (N_3305,N_3136,N_3117);
or U3306 (N_3306,N_3175,N_3062);
nand U3307 (N_3307,N_3148,N_3185);
nand U3308 (N_3308,N_3116,N_3004);
nor U3309 (N_3309,N_3082,N_3003);
or U3310 (N_3310,N_3007,N_3134);
nand U3311 (N_3311,N_3115,N_3050);
nor U3312 (N_3312,N_3099,N_3133);
nor U3313 (N_3313,N_3063,N_3051);
nand U3314 (N_3314,N_3171,N_3068);
nand U3315 (N_3315,N_3035,N_3151);
nor U3316 (N_3316,N_3075,N_3196);
nor U3317 (N_3317,N_3113,N_3037);
or U3318 (N_3318,N_3186,N_3000);
and U3319 (N_3319,N_3165,N_3020);
nor U3320 (N_3320,N_3119,N_3058);
nor U3321 (N_3321,N_3043,N_3152);
and U3322 (N_3322,N_3100,N_3118);
and U3323 (N_3323,N_3081,N_3152);
and U3324 (N_3324,N_3139,N_3081);
or U3325 (N_3325,N_3021,N_3047);
nand U3326 (N_3326,N_3131,N_3043);
and U3327 (N_3327,N_3000,N_3059);
nand U3328 (N_3328,N_3080,N_3014);
or U3329 (N_3329,N_3151,N_3078);
nand U3330 (N_3330,N_3029,N_3086);
nand U3331 (N_3331,N_3172,N_3078);
or U3332 (N_3332,N_3085,N_3084);
and U3333 (N_3333,N_3191,N_3139);
nor U3334 (N_3334,N_3120,N_3161);
nor U3335 (N_3335,N_3123,N_3196);
or U3336 (N_3336,N_3070,N_3055);
nor U3337 (N_3337,N_3013,N_3193);
nor U3338 (N_3338,N_3101,N_3089);
nand U3339 (N_3339,N_3186,N_3007);
nor U3340 (N_3340,N_3092,N_3045);
and U3341 (N_3341,N_3122,N_3020);
and U3342 (N_3342,N_3047,N_3012);
nand U3343 (N_3343,N_3074,N_3028);
and U3344 (N_3344,N_3185,N_3015);
nor U3345 (N_3345,N_3095,N_3061);
nand U3346 (N_3346,N_3000,N_3123);
nor U3347 (N_3347,N_3005,N_3008);
or U3348 (N_3348,N_3087,N_3184);
or U3349 (N_3349,N_3127,N_3057);
nand U3350 (N_3350,N_3009,N_3084);
nor U3351 (N_3351,N_3015,N_3052);
nor U3352 (N_3352,N_3189,N_3145);
nor U3353 (N_3353,N_3156,N_3095);
or U3354 (N_3354,N_3189,N_3159);
nor U3355 (N_3355,N_3046,N_3062);
nor U3356 (N_3356,N_3032,N_3196);
and U3357 (N_3357,N_3081,N_3034);
or U3358 (N_3358,N_3082,N_3066);
or U3359 (N_3359,N_3134,N_3168);
nor U3360 (N_3360,N_3021,N_3061);
and U3361 (N_3361,N_3170,N_3072);
and U3362 (N_3362,N_3184,N_3187);
nor U3363 (N_3363,N_3110,N_3163);
nand U3364 (N_3364,N_3157,N_3096);
or U3365 (N_3365,N_3038,N_3172);
nor U3366 (N_3366,N_3167,N_3034);
and U3367 (N_3367,N_3109,N_3158);
and U3368 (N_3368,N_3139,N_3005);
nor U3369 (N_3369,N_3048,N_3019);
nand U3370 (N_3370,N_3024,N_3009);
and U3371 (N_3371,N_3056,N_3117);
nand U3372 (N_3372,N_3065,N_3156);
nand U3373 (N_3373,N_3032,N_3094);
and U3374 (N_3374,N_3178,N_3167);
nor U3375 (N_3375,N_3042,N_3181);
or U3376 (N_3376,N_3160,N_3065);
nor U3377 (N_3377,N_3099,N_3142);
nor U3378 (N_3378,N_3181,N_3104);
and U3379 (N_3379,N_3017,N_3083);
nand U3380 (N_3380,N_3152,N_3173);
nor U3381 (N_3381,N_3181,N_3169);
nand U3382 (N_3382,N_3086,N_3180);
or U3383 (N_3383,N_3023,N_3004);
and U3384 (N_3384,N_3053,N_3187);
nand U3385 (N_3385,N_3087,N_3063);
and U3386 (N_3386,N_3114,N_3116);
or U3387 (N_3387,N_3133,N_3190);
or U3388 (N_3388,N_3089,N_3044);
nand U3389 (N_3389,N_3008,N_3021);
or U3390 (N_3390,N_3116,N_3051);
nor U3391 (N_3391,N_3064,N_3115);
nor U3392 (N_3392,N_3126,N_3139);
nor U3393 (N_3393,N_3036,N_3072);
nand U3394 (N_3394,N_3146,N_3101);
and U3395 (N_3395,N_3122,N_3157);
nand U3396 (N_3396,N_3022,N_3019);
nand U3397 (N_3397,N_3170,N_3015);
and U3398 (N_3398,N_3092,N_3181);
or U3399 (N_3399,N_3190,N_3062);
and U3400 (N_3400,N_3247,N_3343);
nand U3401 (N_3401,N_3207,N_3281);
and U3402 (N_3402,N_3289,N_3366);
or U3403 (N_3403,N_3228,N_3326);
nor U3404 (N_3404,N_3220,N_3230);
and U3405 (N_3405,N_3330,N_3285);
and U3406 (N_3406,N_3331,N_3306);
xnor U3407 (N_3407,N_3335,N_3292);
xnor U3408 (N_3408,N_3344,N_3268);
nor U3409 (N_3409,N_3209,N_3234);
nor U3410 (N_3410,N_3244,N_3273);
nor U3411 (N_3411,N_3338,N_3210);
and U3412 (N_3412,N_3382,N_3358);
nand U3413 (N_3413,N_3216,N_3327);
and U3414 (N_3414,N_3386,N_3368);
or U3415 (N_3415,N_3391,N_3266);
nand U3416 (N_3416,N_3373,N_3224);
or U3417 (N_3417,N_3283,N_3323);
nor U3418 (N_3418,N_3233,N_3305);
and U3419 (N_3419,N_3267,N_3262);
nand U3420 (N_3420,N_3299,N_3212);
and U3421 (N_3421,N_3282,N_3302);
nor U3422 (N_3422,N_3340,N_3387);
nor U3423 (N_3423,N_3258,N_3355);
nor U3424 (N_3424,N_3398,N_3385);
or U3425 (N_3425,N_3278,N_3201);
nor U3426 (N_3426,N_3265,N_3333);
nand U3427 (N_3427,N_3375,N_3222);
nor U3428 (N_3428,N_3249,N_3328);
or U3429 (N_3429,N_3237,N_3242);
and U3430 (N_3430,N_3360,N_3232);
nor U3431 (N_3431,N_3239,N_3378);
and U3432 (N_3432,N_3284,N_3351);
xnor U3433 (N_3433,N_3356,N_3397);
or U3434 (N_3434,N_3280,N_3269);
or U3435 (N_3435,N_3223,N_3213);
or U3436 (N_3436,N_3384,N_3322);
or U3437 (N_3437,N_3371,N_3349);
nor U3438 (N_3438,N_3245,N_3252);
or U3439 (N_3439,N_3246,N_3253);
nor U3440 (N_3440,N_3394,N_3229);
nor U3441 (N_3441,N_3240,N_3297);
or U3442 (N_3442,N_3308,N_3257);
and U3443 (N_3443,N_3298,N_3369);
nor U3444 (N_3444,N_3365,N_3286);
nor U3445 (N_3445,N_3295,N_3300);
nand U3446 (N_3446,N_3259,N_3309);
nor U3447 (N_3447,N_3337,N_3264);
nor U3448 (N_3448,N_3241,N_3321);
xor U3449 (N_3449,N_3251,N_3279);
or U3450 (N_3450,N_3270,N_3383);
nand U3451 (N_3451,N_3236,N_3315);
nor U3452 (N_3452,N_3296,N_3380);
or U3453 (N_3453,N_3332,N_3354);
and U3454 (N_3454,N_3352,N_3218);
nand U3455 (N_3455,N_3392,N_3260);
and U3456 (N_3456,N_3291,N_3334);
and U3457 (N_3457,N_3348,N_3275);
nor U3458 (N_3458,N_3219,N_3290);
or U3459 (N_3459,N_3206,N_3395);
or U3460 (N_3460,N_3362,N_3341);
or U3461 (N_3461,N_3250,N_3320);
nand U3462 (N_3462,N_3324,N_3377);
nand U3463 (N_3463,N_3339,N_3381);
nand U3464 (N_3464,N_3288,N_3347);
and U3465 (N_3465,N_3255,N_3263);
nor U3466 (N_3466,N_3346,N_3226);
nand U3467 (N_3467,N_3204,N_3271);
nand U3468 (N_3468,N_3202,N_3208);
or U3469 (N_3469,N_3256,N_3310);
or U3470 (N_3470,N_3221,N_3316);
and U3471 (N_3471,N_3248,N_3363);
nand U3472 (N_3472,N_3374,N_3238);
and U3473 (N_3473,N_3200,N_3361);
or U3474 (N_3474,N_3336,N_3376);
and U3475 (N_3475,N_3388,N_3203);
nor U3476 (N_3476,N_3307,N_3276);
and U3477 (N_3477,N_3372,N_3205);
or U3478 (N_3478,N_3301,N_3367);
nand U3479 (N_3479,N_3370,N_3311);
nor U3480 (N_3480,N_3314,N_3318);
or U3481 (N_3481,N_3293,N_3393);
nor U3482 (N_3482,N_3287,N_3225);
and U3483 (N_3483,N_3227,N_3304);
or U3484 (N_3484,N_3217,N_3231);
nor U3485 (N_3485,N_3390,N_3379);
nor U3486 (N_3486,N_3319,N_3294);
nand U3487 (N_3487,N_3312,N_3215);
nand U3488 (N_3488,N_3243,N_3353);
nor U3489 (N_3489,N_3399,N_3359);
or U3490 (N_3490,N_3317,N_3214);
nand U3491 (N_3491,N_3261,N_3235);
or U3492 (N_3492,N_3211,N_3345);
nand U3493 (N_3493,N_3254,N_3389);
nor U3494 (N_3494,N_3313,N_3329);
and U3495 (N_3495,N_3364,N_3342);
and U3496 (N_3496,N_3272,N_3350);
and U3497 (N_3497,N_3396,N_3357);
or U3498 (N_3498,N_3325,N_3303);
nand U3499 (N_3499,N_3274,N_3277);
nor U3500 (N_3500,N_3201,N_3361);
nand U3501 (N_3501,N_3203,N_3223);
nand U3502 (N_3502,N_3391,N_3270);
nor U3503 (N_3503,N_3215,N_3390);
nand U3504 (N_3504,N_3294,N_3287);
xor U3505 (N_3505,N_3329,N_3276);
and U3506 (N_3506,N_3279,N_3300);
nand U3507 (N_3507,N_3283,N_3346);
and U3508 (N_3508,N_3278,N_3220);
nor U3509 (N_3509,N_3354,N_3234);
and U3510 (N_3510,N_3397,N_3285);
nor U3511 (N_3511,N_3227,N_3318);
and U3512 (N_3512,N_3390,N_3239);
and U3513 (N_3513,N_3244,N_3307);
and U3514 (N_3514,N_3200,N_3261);
nor U3515 (N_3515,N_3328,N_3246);
or U3516 (N_3516,N_3215,N_3310);
nor U3517 (N_3517,N_3259,N_3238);
nand U3518 (N_3518,N_3227,N_3232);
nor U3519 (N_3519,N_3392,N_3280);
or U3520 (N_3520,N_3256,N_3331);
nor U3521 (N_3521,N_3240,N_3217);
nor U3522 (N_3522,N_3354,N_3385);
and U3523 (N_3523,N_3311,N_3268);
and U3524 (N_3524,N_3348,N_3394);
nor U3525 (N_3525,N_3212,N_3318);
nand U3526 (N_3526,N_3335,N_3223);
nand U3527 (N_3527,N_3355,N_3336);
or U3528 (N_3528,N_3309,N_3367);
nor U3529 (N_3529,N_3314,N_3288);
nand U3530 (N_3530,N_3365,N_3271);
nand U3531 (N_3531,N_3338,N_3375);
and U3532 (N_3532,N_3225,N_3258);
nor U3533 (N_3533,N_3336,N_3225);
nor U3534 (N_3534,N_3375,N_3304);
and U3535 (N_3535,N_3246,N_3326);
and U3536 (N_3536,N_3375,N_3207);
nand U3537 (N_3537,N_3278,N_3357);
nand U3538 (N_3538,N_3216,N_3379);
and U3539 (N_3539,N_3211,N_3339);
and U3540 (N_3540,N_3376,N_3350);
or U3541 (N_3541,N_3259,N_3357);
nand U3542 (N_3542,N_3280,N_3388);
and U3543 (N_3543,N_3354,N_3338);
and U3544 (N_3544,N_3388,N_3331);
nor U3545 (N_3545,N_3290,N_3354);
and U3546 (N_3546,N_3388,N_3231);
and U3547 (N_3547,N_3271,N_3285);
and U3548 (N_3548,N_3210,N_3310);
or U3549 (N_3549,N_3242,N_3276);
and U3550 (N_3550,N_3220,N_3248);
and U3551 (N_3551,N_3317,N_3360);
nand U3552 (N_3552,N_3233,N_3366);
nor U3553 (N_3553,N_3212,N_3204);
nand U3554 (N_3554,N_3379,N_3327);
nand U3555 (N_3555,N_3306,N_3364);
or U3556 (N_3556,N_3310,N_3255);
and U3557 (N_3557,N_3289,N_3360);
nand U3558 (N_3558,N_3271,N_3213);
and U3559 (N_3559,N_3347,N_3251);
or U3560 (N_3560,N_3314,N_3337);
nand U3561 (N_3561,N_3227,N_3317);
nor U3562 (N_3562,N_3310,N_3353);
or U3563 (N_3563,N_3324,N_3296);
and U3564 (N_3564,N_3251,N_3312);
nor U3565 (N_3565,N_3275,N_3389);
nor U3566 (N_3566,N_3304,N_3279);
or U3567 (N_3567,N_3310,N_3208);
nor U3568 (N_3568,N_3298,N_3325);
nor U3569 (N_3569,N_3387,N_3213);
or U3570 (N_3570,N_3295,N_3393);
nor U3571 (N_3571,N_3231,N_3279);
nand U3572 (N_3572,N_3227,N_3350);
nor U3573 (N_3573,N_3210,N_3277);
or U3574 (N_3574,N_3242,N_3359);
or U3575 (N_3575,N_3330,N_3244);
or U3576 (N_3576,N_3294,N_3341);
or U3577 (N_3577,N_3257,N_3200);
and U3578 (N_3578,N_3257,N_3256);
nand U3579 (N_3579,N_3202,N_3358);
nor U3580 (N_3580,N_3208,N_3268);
and U3581 (N_3581,N_3252,N_3251);
and U3582 (N_3582,N_3230,N_3354);
nand U3583 (N_3583,N_3288,N_3334);
or U3584 (N_3584,N_3348,N_3327);
nor U3585 (N_3585,N_3230,N_3216);
and U3586 (N_3586,N_3391,N_3307);
nand U3587 (N_3587,N_3221,N_3345);
and U3588 (N_3588,N_3259,N_3249);
nor U3589 (N_3589,N_3364,N_3292);
and U3590 (N_3590,N_3216,N_3345);
xor U3591 (N_3591,N_3204,N_3293);
or U3592 (N_3592,N_3284,N_3218);
or U3593 (N_3593,N_3352,N_3293);
nor U3594 (N_3594,N_3252,N_3211);
nand U3595 (N_3595,N_3313,N_3226);
or U3596 (N_3596,N_3233,N_3231);
nand U3597 (N_3597,N_3316,N_3368);
nand U3598 (N_3598,N_3322,N_3299);
nor U3599 (N_3599,N_3313,N_3307);
or U3600 (N_3600,N_3427,N_3494);
nand U3601 (N_3601,N_3462,N_3414);
nand U3602 (N_3602,N_3415,N_3450);
nor U3603 (N_3603,N_3546,N_3472);
nor U3604 (N_3604,N_3528,N_3481);
and U3605 (N_3605,N_3547,N_3422);
or U3606 (N_3606,N_3521,N_3435);
or U3607 (N_3607,N_3479,N_3585);
nand U3608 (N_3608,N_3562,N_3413);
and U3609 (N_3609,N_3556,N_3540);
and U3610 (N_3610,N_3590,N_3424);
nand U3611 (N_3611,N_3572,N_3593);
nand U3612 (N_3612,N_3488,N_3516);
nand U3613 (N_3613,N_3577,N_3430);
or U3614 (N_3614,N_3486,N_3407);
and U3615 (N_3615,N_3538,N_3477);
nand U3616 (N_3616,N_3511,N_3532);
nor U3617 (N_3617,N_3550,N_3519);
and U3618 (N_3618,N_3558,N_3594);
nand U3619 (N_3619,N_3412,N_3518);
nand U3620 (N_3620,N_3539,N_3416);
and U3621 (N_3621,N_3551,N_3581);
nand U3622 (N_3622,N_3542,N_3433);
or U3623 (N_3623,N_3478,N_3557);
or U3624 (N_3624,N_3492,N_3501);
and U3625 (N_3625,N_3440,N_3506);
nand U3626 (N_3626,N_3434,N_3460);
and U3627 (N_3627,N_3443,N_3497);
nor U3628 (N_3628,N_3476,N_3522);
xnor U3629 (N_3629,N_3564,N_3586);
nor U3630 (N_3630,N_3406,N_3510);
nand U3631 (N_3631,N_3587,N_3534);
nor U3632 (N_3632,N_3439,N_3451);
and U3633 (N_3633,N_3405,N_3583);
nand U3634 (N_3634,N_3491,N_3535);
nand U3635 (N_3635,N_3589,N_3504);
nand U3636 (N_3636,N_3468,N_3567);
or U3637 (N_3637,N_3541,N_3467);
nand U3638 (N_3638,N_3463,N_3552);
and U3639 (N_3639,N_3599,N_3520);
and U3640 (N_3640,N_3484,N_3465);
nor U3641 (N_3641,N_3489,N_3420);
nand U3642 (N_3642,N_3445,N_3570);
and U3643 (N_3643,N_3400,N_3560);
and U3644 (N_3644,N_3448,N_3455);
or U3645 (N_3645,N_3452,N_3576);
and U3646 (N_3646,N_3568,N_3513);
and U3647 (N_3647,N_3574,N_3573);
and U3648 (N_3648,N_3512,N_3490);
and U3649 (N_3649,N_3417,N_3453);
nor U3650 (N_3650,N_3480,N_3505);
or U3651 (N_3651,N_3525,N_3498);
nand U3652 (N_3652,N_3426,N_3571);
or U3653 (N_3653,N_3575,N_3553);
nand U3654 (N_3654,N_3597,N_3409);
or U3655 (N_3655,N_3471,N_3548);
nor U3656 (N_3656,N_3456,N_3565);
xor U3657 (N_3657,N_3580,N_3584);
and U3658 (N_3658,N_3444,N_3598);
and U3659 (N_3659,N_3410,N_3507);
and U3660 (N_3660,N_3531,N_3447);
nand U3661 (N_3661,N_3428,N_3537);
or U3662 (N_3662,N_3429,N_3530);
or U3663 (N_3663,N_3495,N_3543);
nor U3664 (N_3664,N_3561,N_3527);
nand U3665 (N_3665,N_3523,N_3469);
nand U3666 (N_3666,N_3544,N_3503);
nand U3667 (N_3667,N_3421,N_3437);
or U3668 (N_3668,N_3458,N_3402);
nand U3669 (N_3669,N_3419,N_3457);
and U3670 (N_3670,N_3563,N_3432);
and U3671 (N_3671,N_3485,N_3408);
nand U3672 (N_3672,N_3438,N_3517);
or U3673 (N_3673,N_3425,N_3470);
nor U3674 (N_3674,N_3588,N_3554);
nand U3675 (N_3675,N_3493,N_3526);
nand U3676 (N_3676,N_3536,N_3423);
and U3677 (N_3677,N_3403,N_3591);
nor U3678 (N_3678,N_3529,N_3592);
and U3679 (N_3679,N_3482,N_3441);
and U3680 (N_3680,N_3401,N_3533);
nor U3681 (N_3681,N_3508,N_3555);
and U3682 (N_3682,N_3496,N_3524);
and U3683 (N_3683,N_3502,N_3449);
and U3684 (N_3684,N_3475,N_3515);
nor U3685 (N_3685,N_3454,N_3431);
nand U3686 (N_3686,N_3446,N_3596);
or U3687 (N_3687,N_3582,N_3442);
nor U3688 (N_3688,N_3579,N_3500);
nor U3689 (N_3689,N_3461,N_3487);
or U3690 (N_3690,N_3509,N_3418);
nand U3691 (N_3691,N_3483,N_3473);
or U3692 (N_3692,N_3466,N_3595);
nor U3693 (N_3693,N_3514,N_3549);
nand U3694 (N_3694,N_3464,N_3436);
xnor U3695 (N_3695,N_3499,N_3578);
nor U3696 (N_3696,N_3569,N_3459);
and U3697 (N_3697,N_3411,N_3404);
nor U3698 (N_3698,N_3474,N_3559);
nor U3699 (N_3699,N_3566,N_3545);
and U3700 (N_3700,N_3488,N_3555);
nand U3701 (N_3701,N_3470,N_3400);
or U3702 (N_3702,N_3402,N_3574);
nor U3703 (N_3703,N_3505,N_3433);
and U3704 (N_3704,N_3406,N_3472);
nand U3705 (N_3705,N_3501,N_3403);
and U3706 (N_3706,N_3531,N_3438);
xnor U3707 (N_3707,N_3462,N_3483);
and U3708 (N_3708,N_3422,N_3588);
nor U3709 (N_3709,N_3507,N_3515);
and U3710 (N_3710,N_3461,N_3501);
nand U3711 (N_3711,N_3424,N_3463);
or U3712 (N_3712,N_3507,N_3577);
and U3713 (N_3713,N_3452,N_3450);
or U3714 (N_3714,N_3574,N_3533);
or U3715 (N_3715,N_3573,N_3583);
nand U3716 (N_3716,N_3490,N_3457);
and U3717 (N_3717,N_3562,N_3505);
and U3718 (N_3718,N_3551,N_3521);
nor U3719 (N_3719,N_3540,N_3440);
or U3720 (N_3720,N_3563,N_3426);
and U3721 (N_3721,N_3572,N_3503);
or U3722 (N_3722,N_3587,N_3583);
and U3723 (N_3723,N_3501,N_3566);
xnor U3724 (N_3724,N_3530,N_3558);
and U3725 (N_3725,N_3453,N_3445);
or U3726 (N_3726,N_3450,N_3431);
and U3727 (N_3727,N_3583,N_3502);
and U3728 (N_3728,N_3484,N_3486);
nor U3729 (N_3729,N_3457,N_3575);
nor U3730 (N_3730,N_3507,N_3496);
and U3731 (N_3731,N_3454,N_3435);
nor U3732 (N_3732,N_3417,N_3413);
or U3733 (N_3733,N_3579,N_3435);
nand U3734 (N_3734,N_3583,N_3464);
nor U3735 (N_3735,N_3479,N_3582);
or U3736 (N_3736,N_3570,N_3534);
or U3737 (N_3737,N_3547,N_3534);
and U3738 (N_3738,N_3506,N_3412);
nor U3739 (N_3739,N_3463,N_3412);
nor U3740 (N_3740,N_3514,N_3415);
and U3741 (N_3741,N_3542,N_3564);
nand U3742 (N_3742,N_3444,N_3484);
nand U3743 (N_3743,N_3564,N_3552);
or U3744 (N_3744,N_3523,N_3573);
and U3745 (N_3745,N_3568,N_3484);
and U3746 (N_3746,N_3426,N_3581);
and U3747 (N_3747,N_3493,N_3544);
nor U3748 (N_3748,N_3439,N_3532);
nand U3749 (N_3749,N_3571,N_3404);
nor U3750 (N_3750,N_3474,N_3542);
nand U3751 (N_3751,N_3510,N_3518);
or U3752 (N_3752,N_3415,N_3488);
or U3753 (N_3753,N_3430,N_3464);
nand U3754 (N_3754,N_3408,N_3573);
or U3755 (N_3755,N_3418,N_3486);
or U3756 (N_3756,N_3466,N_3578);
nand U3757 (N_3757,N_3552,N_3524);
or U3758 (N_3758,N_3529,N_3487);
and U3759 (N_3759,N_3542,N_3412);
or U3760 (N_3760,N_3569,N_3443);
or U3761 (N_3761,N_3416,N_3551);
or U3762 (N_3762,N_3549,N_3463);
and U3763 (N_3763,N_3493,N_3476);
or U3764 (N_3764,N_3540,N_3415);
nor U3765 (N_3765,N_3432,N_3537);
nor U3766 (N_3766,N_3550,N_3478);
and U3767 (N_3767,N_3507,N_3569);
and U3768 (N_3768,N_3501,N_3402);
nor U3769 (N_3769,N_3463,N_3583);
nand U3770 (N_3770,N_3520,N_3573);
nor U3771 (N_3771,N_3599,N_3587);
and U3772 (N_3772,N_3498,N_3452);
and U3773 (N_3773,N_3597,N_3504);
nand U3774 (N_3774,N_3512,N_3531);
nor U3775 (N_3775,N_3422,N_3423);
or U3776 (N_3776,N_3453,N_3489);
xnor U3777 (N_3777,N_3471,N_3540);
or U3778 (N_3778,N_3545,N_3540);
nand U3779 (N_3779,N_3477,N_3518);
or U3780 (N_3780,N_3518,N_3550);
or U3781 (N_3781,N_3532,N_3404);
nand U3782 (N_3782,N_3585,N_3412);
nand U3783 (N_3783,N_3416,N_3410);
or U3784 (N_3784,N_3504,N_3576);
or U3785 (N_3785,N_3520,N_3596);
nand U3786 (N_3786,N_3512,N_3454);
nand U3787 (N_3787,N_3524,N_3492);
and U3788 (N_3788,N_3558,N_3595);
or U3789 (N_3789,N_3584,N_3599);
or U3790 (N_3790,N_3515,N_3444);
nor U3791 (N_3791,N_3446,N_3485);
and U3792 (N_3792,N_3573,N_3519);
and U3793 (N_3793,N_3556,N_3569);
nor U3794 (N_3794,N_3598,N_3519);
nand U3795 (N_3795,N_3596,N_3476);
or U3796 (N_3796,N_3561,N_3466);
and U3797 (N_3797,N_3422,N_3496);
and U3798 (N_3798,N_3502,N_3537);
nor U3799 (N_3799,N_3581,N_3493);
or U3800 (N_3800,N_3778,N_3698);
nand U3801 (N_3801,N_3607,N_3630);
nand U3802 (N_3802,N_3676,N_3679);
and U3803 (N_3803,N_3635,N_3750);
or U3804 (N_3804,N_3684,N_3755);
and U3805 (N_3805,N_3798,N_3666);
or U3806 (N_3806,N_3770,N_3675);
and U3807 (N_3807,N_3754,N_3612);
nor U3808 (N_3808,N_3642,N_3620);
nand U3809 (N_3809,N_3625,N_3784);
or U3810 (N_3810,N_3711,N_3746);
and U3811 (N_3811,N_3696,N_3732);
nor U3812 (N_3812,N_3748,N_3660);
nand U3813 (N_3813,N_3777,N_3733);
and U3814 (N_3814,N_3749,N_3737);
nor U3815 (N_3815,N_3664,N_3744);
nand U3816 (N_3816,N_3624,N_3788);
nand U3817 (N_3817,N_3735,N_3787);
nand U3818 (N_3818,N_3626,N_3601);
nand U3819 (N_3819,N_3767,N_3700);
and U3820 (N_3820,N_3738,N_3614);
and U3821 (N_3821,N_3685,N_3656);
nand U3822 (N_3822,N_3715,N_3644);
nand U3823 (N_3823,N_3759,N_3793);
or U3824 (N_3824,N_3705,N_3668);
nor U3825 (N_3825,N_3795,N_3722);
or U3826 (N_3826,N_3689,N_3790);
and U3827 (N_3827,N_3670,N_3799);
or U3828 (N_3828,N_3710,N_3613);
nand U3829 (N_3829,N_3783,N_3681);
or U3830 (N_3830,N_3730,N_3712);
nand U3831 (N_3831,N_3682,N_3617);
nand U3832 (N_3832,N_3674,N_3725);
nor U3833 (N_3833,N_3604,N_3618);
or U3834 (N_3834,N_3780,N_3632);
or U3835 (N_3835,N_3693,N_3791);
or U3836 (N_3836,N_3667,N_3728);
and U3837 (N_3837,N_3694,N_3645);
or U3838 (N_3838,N_3756,N_3761);
or U3839 (N_3839,N_3794,N_3641);
nand U3840 (N_3840,N_3747,N_3707);
or U3841 (N_3841,N_3629,N_3655);
and U3842 (N_3842,N_3623,N_3622);
nor U3843 (N_3843,N_3619,N_3771);
nand U3844 (N_3844,N_3796,N_3661);
or U3845 (N_3845,N_3786,N_3669);
nor U3846 (N_3846,N_3648,N_3701);
nand U3847 (N_3847,N_3640,N_3729);
nand U3848 (N_3848,N_3602,N_3686);
nor U3849 (N_3849,N_3646,N_3683);
nor U3850 (N_3850,N_3719,N_3751);
or U3851 (N_3851,N_3727,N_3766);
or U3852 (N_3852,N_3610,N_3721);
nand U3853 (N_3853,N_3713,N_3690);
nor U3854 (N_3854,N_3647,N_3714);
nor U3855 (N_3855,N_3739,N_3758);
and U3856 (N_3856,N_3680,N_3768);
nand U3857 (N_3857,N_3717,N_3678);
nor U3858 (N_3858,N_3764,N_3774);
and U3859 (N_3859,N_3709,N_3651);
nand U3860 (N_3860,N_3621,N_3763);
and U3861 (N_3861,N_3745,N_3782);
nor U3862 (N_3862,N_3734,N_3743);
or U3863 (N_3863,N_3781,N_3703);
nand U3864 (N_3864,N_3697,N_3775);
nor U3865 (N_3865,N_3688,N_3760);
nor U3866 (N_3866,N_3662,N_3636);
nand U3867 (N_3867,N_3762,N_3776);
or U3868 (N_3868,N_3731,N_3772);
or U3869 (N_3869,N_3720,N_3627);
nand U3870 (N_3870,N_3633,N_3650);
and U3871 (N_3871,N_3658,N_3616);
nor U3872 (N_3872,N_3615,N_3718);
and U3873 (N_3873,N_3706,N_3665);
or U3874 (N_3874,N_3789,N_3652);
nor U3875 (N_3875,N_3653,N_3785);
and U3876 (N_3876,N_3692,N_3659);
nor U3877 (N_3877,N_3631,N_3638);
or U3878 (N_3878,N_3736,N_3657);
or U3879 (N_3879,N_3606,N_3649);
nand U3880 (N_3880,N_3671,N_3773);
nor U3881 (N_3881,N_3792,N_3677);
or U3882 (N_3882,N_3752,N_3726);
and U3883 (N_3883,N_3779,N_3757);
nor U3884 (N_3884,N_3742,N_3634);
nor U3885 (N_3885,N_3608,N_3704);
nor U3886 (N_3886,N_3673,N_3643);
or U3887 (N_3887,N_3702,N_3672);
and U3888 (N_3888,N_3708,N_3611);
nand U3889 (N_3889,N_3603,N_3769);
or U3890 (N_3890,N_3753,N_3723);
nand U3891 (N_3891,N_3716,N_3699);
and U3892 (N_3892,N_3609,N_3740);
or U3893 (N_3893,N_3654,N_3741);
nand U3894 (N_3894,N_3600,N_3605);
and U3895 (N_3895,N_3765,N_3687);
nand U3896 (N_3896,N_3639,N_3663);
xor U3897 (N_3897,N_3628,N_3691);
and U3898 (N_3898,N_3695,N_3724);
and U3899 (N_3899,N_3797,N_3637);
and U3900 (N_3900,N_3704,N_3664);
or U3901 (N_3901,N_3761,N_3783);
nor U3902 (N_3902,N_3636,N_3733);
or U3903 (N_3903,N_3762,N_3715);
or U3904 (N_3904,N_3767,N_3740);
xnor U3905 (N_3905,N_3661,N_3685);
or U3906 (N_3906,N_3730,N_3745);
nand U3907 (N_3907,N_3614,N_3682);
nor U3908 (N_3908,N_3730,N_3689);
nor U3909 (N_3909,N_3792,N_3682);
nand U3910 (N_3910,N_3744,N_3637);
nand U3911 (N_3911,N_3672,N_3600);
and U3912 (N_3912,N_3770,N_3642);
nand U3913 (N_3913,N_3625,N_3676);
nand U3914 (N_3914,N_3656,N_3742);
nand U3915 (N_3915,N_3649,N_3629);
nand U3916 (N_3916,N_3784,N_3776);
and U3917 (N_3917,N_3786,N_3701);
nand U3918 (N_3918,N_3785,N_3707);
nand U3919 (N_3919,N_3619,N_3763);
nand U3920 (N_3920,N_3745,N_3671);
nor U3921 (N_3921,N_3635,N_3621);
nor U3922 (N_3922,N_3763,N_3765);
nor U3923 (N_3923,N_3711,N_3797);
or U3924 (N_3924,N_3685,N_3700);
nor U3925 (N_3925,N_3638,N_3755);
nand U3926 (N_3926,N_3689,N_3711);
nand U3927 (N_3927,N_3678,N_3714);
nor U3928 (N_3928,N_3783,N_3634);
or U3929 (N_3929,N_3651,N_3697);
nor U3930 (N_3930,N_3709,N_3797);
and U3931 (N_3931,N_3704,N_3779);
or U3932 (N_3932,N_3790,N_3791);
nor U3933 (N_3933,N_3777,N_3731);
nand U3934 (N_3934,N_3766,N_3629);
nor U3935 (N_3935,N_3795,N_3660);
nor U3936 (N_3936,N_3711,N_3623);
nor U3937 (N_3937,N_3665,N_3600);
nor U3938 (N_3938,N_3728,N_3797);
or U3939 (N_3939,N_3724,N_3682);
or U3940 (N_3940,N_3620,N_3673);
or U3941 (N_3941,N_3768,N_3677);
nor U3942 (N_3942,N_3622,N_3758);
nand U3943 (N_3943,N_3733,N_3667);
or U3944 (N_3944,N_3683,N_3761);
nand U3945 (N_3945,N_3634,N_3766);
and U3946 (N_3946,N_3651,N_3609);
and U3947 (N_3947,N_3675,N_3742);
and U3948 (N_3948,N_3768,N_3688);
nor U3949 (N_3949,N_3796,N_3637);
and U3950 (N_3950,N_3694,N_3788);
and U3951 (N_3951,N_3707,N_3774);
nand U3952 (N_3952,N_3734,N_3756);
nand U3953 (N_3953,N_3748,N_3694);
xor U3954 (N_3954,N_3685,N_3669);
and U3955 (N_3955,N_3767,N_3668);
and U3956 (N_3956,N_3692,N_3780);
nand U3957 (N_3957,N_3696,N_3606);
nand U3958 (N_3958,N_3784,N_3676);
and U3959 (N_3959,N_3763,N_3713);
nand U3960 (N_3960,N_3743,N_3605);
and U3961 (N_3961,N_3619,N_3782);
or U3962 (N_3962,N_3631,N_3736);
nand U3963 (N_3963,N_3676,N_3776);
nand U3964 (N_3964,N_3757,N_3721);
nand U3965 (N_3965,N_3769,N_3708);
and U3966 (N_3966,N_3721,N_3778);
or U3967 (N_3967,N_3610,N_3705);
and U3968 (N_3968,N_3653,N_3798);
nand U3969 (N_3969,N_3658,N_3745);
nand U3970 (N_3970,N_3625,N_3793);
or U3971 (N_3971,N_3704,N_3645);
nand U3972 (N_3972,N_3650,N_3745);
nor U3973 (N_3973,N_3692,N_3726);
nor U3974 (N_3974,N_3681,N_3707);
or U3975 (N_3975,N_3683,N_3769);
or U3976 (N_3976,N_3713,N_3754);
or U3977 (N_3977,N_3628,N_3626);
and U3978 (N_3978,N_3652,N_3607);
nand U3979 (N_3979,N_3753,N_3687);
and U3980 (N_3980,N_3602,N_3725);
nor U3981 (N_3981,N_3696,N_3710);
nor U3982 (N_3982,N_3613,N_3730);
and U3983 (N_3983,N_3721,N_3652);
nand U3984 (N_3984,N_3684,N_3773);
or U3985 (N_3985,N_3618,N_3764);
and U3986 (N_3986,N_3767,N_3758);
or U3987 (N_3987,N_3702,N_3643);
and U3988 (N_3988,N_3779,N_3741);
nand U3989 (N_3989,N_3635,N_3658);
nand U3990 (N_3990,N_3734,N_3691);
nor U3991 (N_3991,N_3705,N_3687);
nand U3992 (N_3992,N_3751,N_3686);
and U3993 (N_3993,N_3794,N_3697);
or U3994 (N_3994,N_3762,N_3675);
and U3995 (N_3995,N_3792,N_3739);
and U3996 (N_3996,N_3707,N_3789);
nor U3997 (N_3997,N_3780,N_3740);
nand U3998 (N_3998,N_3659,N_3741);
or U3999 (N_3999,N_3727,N_3718);
and U4000 (N_4000,N_3856,N_3816);
nand U4001 (N_4001,N_3980,N_3973);
or U4002 (N_4002,N_3908,N_3946);
and U4003 (N_4003,N_3822,N_3817);
or U4004 (N_4004,N_3815,N_3880);
or U4005 (N_4005,N_3934,N_3972);
or U4006 (N_4006,N_3885,N_3941);
nor U4007 (N_4007,N_3826,N_3891);
and U4008 (N_4008,N_3921,N_3986);
nand U4009 (N_4009,N_3917,N_3938);
and U4010 (N_4010,N_3871,N_3944);
and U4011 (N_4011,N_3863,N_3870);
nor U4012 (N_4012,N_3926,N_3910);
and U4013 (N_4013,N_3929,N_3902);
nand U4014 (N_4014,N_3967,N_3853);
or U4015 (N_4015,N_3997,N_3834);
nand U4016 (N_4016,N_3922,N_3876);
nand U4017 (N_4017,N_3827,N_3907);
nor U4018 (N_4018,N_3982,N_3868);
or U4019 (N_4019,N_3956,N_3903);
nand U4020 (N_4020,N_3895,N_3805);
nand U4021 (N_4021,N_3989,N_3860);
nor U4022 (N_4022,N_3844,N_3915);
nor U4023 (N_4023,N_3886,N_3840);
or U4024 (N_4024,N_3909,N_3966);
or U4025 (N_4025,N_3906,N_3806);
and U4026 (N_4026,N_3800,N_3912);
xnor U4027 (N_4027,N_3983,N_3869);
nor U4028 (N_4028,N_3803,N_3862);
nand U4029 (N_4029,N_3958,N_3961);
nand U4030 (N_4030,N_3890,N_3984);
or U4031 (N_4031,N_3998,N_3810);
nor U4032 (N_4032,N_3814,N_3925);
nand U4033 (N_4033,N_3883,N_3936);
or U4034 (N_4034,N_3951,N_3935);
or U4035 (N_4035,N_3999,N_3889);
nor U4036 (N_4036,N_3959,N_3988);
nor U4037 (N_4037,N_3969,N_3964);
nor U4038 (N_4038,N_3893,N_3924);
or U4039 (N_4039,N_3847,N_3994);
and U4040 (N_4040,N_3801,N_3829);
or U4041 (N_4041,N_3884,N_3931);
nor U4042 (N_4042,N_3874,N_3887);
nor U4043 (N_4043,N_3948,N_3954);
nor U4044 (N_4044,N_3821,N_3975);
nand U4045 (N_4045,N_3963,N_3899);
nand U4046 (N_4046,N_3960,N_3804);
or U4047 (N_4047,N_3913,N_3904);
nand U4048 (N_4048,N_3828,N_3830);
and U4049 (N_4049,N_3841,N_3916);
nand U4050 (N_4050,N_3937,N_3851);
and U4051 (N_4051,N_3859,N_3819);
nand U4052 (N_4052,N_3952,N_3914);
and U4053 (N_4053,N_3993,N_3878);
nand U4054 (N_4054,N_3832,N_3968);
and U4055 (N_4055,N_3809,N_3850);
or U4056 (N_4056,N_3802,N_3962);
or U4057 (N_4057,N_3990,N_3918);
and U4058 (N_4058,N_3808,N_3930);
nor U4059 (N_4059,N_3977,N_3858);
nand U4060 (N_4060,N_3970,N_3981);
or U4061 (N_4061,N_3985,N_3807);
nor U4062 (N_4062,N_3881,N_3875);
nor U4063 (N_4063,N_3825,N_3947);
nor U4064 (N_4064,N_3901,N_3939);
and U4065 (N_4065,N_3911,N_3919);
and U4066 (N_4066,N_3965,N_3824);
nand U4067 (N_4067,N_3849,N_3971);
nand U4068 (N_4068,N_3974,N_3818);
nor U4069 (N_4069,N_3945,N_3811);
nand U4070 (N_4070,N_3976,N_3896);
nand U4071 (N_4071,N_3812,N_3866);
nor U4072 (N_4072,N_3836,N_3845);
nor U4073 (N_4073,N_3835,N_3882);
or U4074 (N_4074,N_3855,N_3894);
nand U4075 (N_4075,N_3839,N_3979);
or U4076 (N_4076,N_3987,N_3996);
nor U4077 (N_4077,N_3897,N_3932);
nand U4078 (N_4078,N_3978,N_3861);
and U4079 (N_4079,N_3838,N_3949);
nand U4080 (N_4080,N_3865,N_3831);
or U4081 (N_4081,N_3940,N_3823);
or U4082 (N_4082,N_3995,N_3848);
and U4083 (N_4083,N_3953,N_3873);
and U4084 (N_4084,N_3864,N_3852);
nand U4085 (N_4085,N_3892,N_3842);
or U4086 (N_4086,N_3837,N_3905);
nor U4087 (N_4087,N_3933,N_3833);
nand U4088 (N_4088,N_3992,N_3857);
nor U4089 (N_4089,N_3813,N_3879);
nand U4090 (N_4090,N_3927,N_3942);
nor U4091 (N_4091,N_3888,N_3877);
nand U4092 (N_4092,N_3955,N_3923);
and U4093 (N_4093,N_3991,N_3957);
or U4094 (N_4094,N_3872,N_3943);
and U4095 (N_4095,N_3843,N_3950);
nand U4096 (N_4096,N_3928,N_3854);
nor U4097 (N_4097,N_3900,N_3898);
nor U4098 (N_4098,N_3846,N_3820);
and U4099 (N_4099,N_3920,N_3867);
nor U4100 (N_4100,N_3929,N_3925);
nor U4101 (N_4101,N_3819,N_3926);
or U4102 (N_4102,N_3974,N_3899);
or U4103 (N_4103,N_3934,N_3905);
and U4104 (N_4104,N_3972,N_3833);
and U4105 (N_4105,N_3907,N_3879);
or U4106 (N_4106,N_3858,N_3830);
or U4107 (N_4107,N_3994,N_3972);
nand U4108 (N_4108,N_3863,N_3984);
or U4109 (N_4109,N_3837,N_3997);
or U4110 (N_4110,N_3892,N_3908);
nor U4111 (N_4111,N_3939,N_3805);
and U4112 (N_4112,N_3847,N_3866);
or U4113 (N_4113,N_3994,N_3825);
nand U4114 (N_4114,N_3845,N_3912);
and U4115 (N_4115,N_3937,N_3990);
or U4116 (N_4116,N_3900,N_3828);
nand U4117 (N_4117,N_3956,N_3825);
or U4118 (N_4118,N_3976,N_3877);
nor U4119 (N_4119,N_3953,N_3934);
nor U4120 (N_4120,N_3914,N_3869);
and U4121 (N_4121,N_3862,N_3875);
nor U4122 (N_4122,N_3999,N_3902);
nor U4123 (N_4123,N_3802,N_3819);
nand U4124 (N_4124,N_3991,N_3828);
nor U4125 (N_4125,N_3921,N_3804);
nor U4126 (N_4126,N_3993,N_3976);
xnor U4127 (N_4127,N_3979,N_3985);
nand U4128 (N_4128,N_3818,N_3899);
and U4129 (N_4129,N_3990,N_3913);
nand U4130 (N_4130,N_3829,N_3907);
nor U4131 (N_4131,N_3902,N_3800);
nand U4132 (N_4132,N_3895,N_3987);
nor U4133 (N_4133,N_3979,N_3855);
nor U4134 (N_4134,N_3902,N_3998);
and U4135 (N_4135,N_3943,N_3928);
nor U4136 (N_4136,N_3880,N_3898);
or U4137 (N_4137,N_3852,N_3974);
nand U4138 (N_4138,N_3972,N_3823);
nand U4139 (N_4139,N_3815,N_3905);
nand U4140 (N_4140,N_3929,N_3996);
nand U4141 (N_4141,N_3857,N_3943);
or U4142 (N_4142,N_3979,N_3944);
and U4143 (N_4143,N_3920,N_3805);
nand U4144 (N_4144,N_3843,N_3993);
or U4145 (N_4145,N_3961,N_3988);
nor U4146 (N_4146,N_3946,N_3863);
and U4147 (N_4147,N_3979,N_3802);
nor U4148 (N_4148,N_3941,N_3845);
nor U4149 (N_4149,N_3881,N_3894);
nor U4150 (N_4150,N_3817,N_3857);
and U4151 (N_4151,N_3805,N_3963);
and U4152 (N_4152,N_3902,N_3848);
or U4153 (N_4153,N_3830,N_3881);
nor U4154 (N_4154,N_3871,N_3849);
or U4155 (N_4155,N_3919,N_3958);
or U4156 (N_4156,N_3990,N_3893);
nand U4157 (N_4157,N_3810,N_3946);
and U4158 (N_4158,N_3852,N_3866);
nor U4159 (N_4159,N_3860,N_3801);
nand U4160 (N_4160,N_3878,N_3994);
nand U4161 (N_4161,N_3836,N_3920);
nor U4162 (N_4162,N_3974,N_3902);
nor U4163 (N_4163,N_3826,N_3929);
nand U4164 (N_4164,N_3857,N_3870);
and U4165 (N_4165,N_3877,N_3940);
and U4166 (N_4166,N_3818,N_3819);
or U4167 (N_4167,N_3829,N_3842);
nand U4168 (N_4168,N_3939,N_3982);
nand U4169 (N_4169,N_3912,N_3861);
nor U4170 (N_4170,N_3901,N_3993);
and U4171 (N_4171,N_3996,N_3850);
nand U4172 (N_4172,N_3906,N_3953);
or U4173 (N_4173,N_3880,N_3847);
nor U4174 (N_4174,N_3919,N_3946);
nor U4175 (N_4175,N_3829,N_3849);
and U4176 (N_4176,N_3950,N_3976);
nor U4177 (N_4177,N_3880,N_3916);
or U4178 (N_4178,N_3803,N_3882);
nand U4179 (N_4179,N_3903,N_3822);
and U4180 (N_4180,N_3998,N_3830);
nand U4181 (N_4181,N_3879,N_3930);
nor U4182 (N_4182,N_3989,N_3994);
nand U4183 (N_4183,N_3972,N_3916);
nor U4184 (N_4184,N_3859,N_3925);
nor U4185 (N_4185,N_3836,N_3966);
or U4186 (N_4186,N_3934,N_3817);
and U4187 (N_4187,N_3998,N_3814);
or U4188 (N_4188,N_3997,N_3925);
nand U4189 (N_4189,N_3961,N_3947);
and U4190 (N_4190,N_3892,N_3856);
nor U4191 (N_4191,N_3883,N_3847);
or U4192 (N_4192,N_3971,N_3864);
and U4193 (N_4193,N_3927,N_3906);
or U4194 (N_4194,N_3956,N_3953);
nand U4195 (N_4195,N_3880,N_3899);
nand U4196 (N_4196,N_3811,N_3830);
nor U4197 (N_4197,N_3957,N_3927);
or U4198 (N_4198,N_3838,N_3945);
nand U4199 (N_4199,N_3954,N_3822);
or U4200 (N_4200,N_4181,N_4019);
and U4201 (N_4201,N_4049,N_4074);
nor U4202 (N_4202,N_4128,N_4030);
and U4203 (N_4203,N_4044,N_4184);
nand U4204 (N_4204,N_4121,N_4195);
and U4205 (N_4205,N_4018,N_4084);
nor U4206 (N_4206,N_4156,N_4176);
or U4207 (N_4207,N_4015,N_4066);
nor U4208 (N_4208,N_4021,N_4114);
or U4209 (N_4209,N_4082,N_4093);
nor U4210 (N_4210,N_4078,N_4132);
and U4211 (N_4211,N_4142,N_4081);
nand U4212 (N_4212,N_4000,N_4172);
nand U4213 (N_4213,N_4163,N_4035);
nand U4214 (N_4214,N_4186,N_4061);
or U4215 (N_4215,N_4063,N_4183);
and U4216 (N_4216,N_4130,N_4103);
nand U4217 (N_4217,N_4024,N_4145);
and U4218 (N_4218,N_4110,N_4029);
nand U4219 (N_4219,N_4127,N_4146);
nand U4220 (N_4220,N_4005,N_4067);
and U4221 (N_4221,N_4158,N_4001);
or U4222 (N_4222,N_4007,N_4010);
and U4223 (N_4223,N_4152,N_4179);
nand U4224 (N_4224,N_4032,N_4149);
and U4225 (N_4225,N_4123,N_4139);
and U4226 (N_4226,N_4174,N_4173);
or U4227 (N_4227,N_4075,N_4002);
xor U4228 (N_4228,N_4124,N_4072);
and U4229 (N_4229,N_4023,N_4085);
or U4230 (N_4230,N_4009,N_4090);
nand U4231 (N_4231,N_4047,N_4046);
or U4232 (N_4232,N_4167,N_4052);
nand U4233 (N_4233,N_4017,N_4162);
and U4234 (N_4234,N_4185,N_4168);
or U4235 (N_4235,N_4095,N_4166);
nor U4236 (N_4236,N_4056,N_4079);
or U4237 (N_4237,N_4137,N_4161);
nor U4238 (N_4238,N_4060,N_4099);
nand U4239 (N_4239,N_4109,N_4054);
nand U4240 (N_4240,N_4004,N_4042);
and U4241 (N_4241,N_4020,N_4113);
or U4242 (N_4242,N_4140,N_4169);
or U4243 (N_4243,N_4198,N_4154);
and U4244 (N_4244,N_4058,N_4129);
and U4245 (N_4245,N_4189,N_4160);
nor U4246 (N_4246,N_4196,N_4094);
and U4247 (N_4247,N_4043,N_4117);
nand U4248 (N_4248,N_4153,N_4126);
or U4249 (N_4249,N_4106,N_4141);
nor U4250 (N_4250,N_4034,N_4151);
or U4251 (N_4251,N_4112,N_4026);
and U4252 (N_4252,N_4182,N_4087);
or U4253 (N_4253,N_4116,N_4008);
or U4254 (N_4254,N_4033,N_4187);
nor U4255 (N_4255,N_4003,N_4125);
or U4256 (N_4256,N_4105,N_4057);
nor U4257 (N_4257,N_4011,N_4091);
or U4258 (N_4258,N_4122,N_4092);
nand U4259 (N_4259,N_4083,N_4144);
and U4260 (N_4260,N_4136,N_4065);
and U4261 (N_4261,N_4016,N_4188);
nor U4262 (N_4262,N_4171,N_4102);
and U4263 (N_4263,N_4076,N_4097);
or U4264 (N_4264,N_4159,N_4107);
nand U4265 (N_4265,N_4088,N_4118);
or U4266 (N_4266,N_4028,N_4077);
nor U4267 (N_4267,N_4108,N_4027);
and U4268 (N_4268,N_4138,N_4073);
or U4269 (N_4269,N_4068,N_4022);
nand U4270 (N_4270,N_4006,N_4148);
nor U4271 (N_4271,N_4135,N_4098);
nand U4272 (N_4272,N_4165,N_4180);
nand U4273 (N_4273,N_4051,N_4037);
or U4274 (N_4274,N_4193,N_4155);
or U4275 (N_4275,N_4080,N_4177);
nor U4276 (N_4276,N_4100,N_4071);
nand U4277 (N_4277,N_4111,N_4040);
and U4278 (N_4278,N_4147,N_4064);
and U4279 (N_4279,N_4119,N_4143);
and U4280 (N_4280,N_4036,N_4150);
nor U4281 (N_4281,N_4059,N_4050);
nand U4282 (N_4282,N_4062,N_4175);
or U4283 (N_4283,N_4197,N_4031);
or U4284 (N_4284,N_4115,N_4089);
or U4285 (N_4285,N_4045,N_4041);
or U4286 (N_4286,N_4199,N_4178);
nor U4287 (N_4287,N_4013,N_4133);
nand U4288 (N_4288,N_4096,N_4086);
nand U4289 (N_4289,N_4039,N_4192);
nand U4290 (N_4290,N_4120,N_4012);
nor U4291 (N_4291,N_4170,N_4038);
and U4292 (N_4292,N_4101,N_4070);
nor U4293 (N_4293,N_4025,N_4134);
or U4294 (N_4294,N_4164,N_4014);
nand U4295 (N_4295,N_4131,N_4104);
nor U4296 (N_4296,N_4190,N_4191);
and U4297 (N_4297,N_4055,N_4048);
or U4298 (N_4298,N_4157,N_4053);
nand U4299 (N_4299,N_4194,N_4069);
nand U4300 (N_4300,N_4118,N_4125);
nor U4301 (N_4301,N_4169,N_4181);
nand U4302 (N_4302,N_4189,N_4143);
and U4303 (N_4303,N_4042,N_4069);
or U4304 (N_4304,N_4026,N_4022);
and U4305 (N_4305,N_4061,N_4152);
and U4306 (N_4306,N_4027,N_4068);
and U4307 (N_4307,N_4193,N_4178);
nand U4308 (N_4308,N_4174,N_4112);
or U4309 (N_4309,N_4104,N_4028);
nor U4310 (N_4310,N_4136,N_4014);
or U4311 (N_4311,N_4159,N_4066);
or U4312 (N_4312,N_4061,N_4121);
and U4313 (N_4313,N_4124,N_4163);
or U4314 (N_4314,N_4114,N_4089);
or U4315 (N_4315,N_4164,N_4171);
nand U4316 (N_4316,N_4195,N_4178);
nand U4317 (N_4317,N_4034,N_4096);
or U4318 (N_4318,N_4179,N_4053);
or U4319 (N_4319,N_4160,N_4069);
nand U4320 (N_4320,N_4013,N_4037);
nand U4321 (N_4321,N_4133,N_4026);
and U4322 (N_4322,N_4044,N_4037);
or U4323 (N_4323,N_4176,N_4118);
nor U4324 (N_4324,N_4196,N_4010);
or U4325 (N_4325,N_4074,N_4146);
nand U4326 (N_4326,N_4164,N_4026);
and U4327 (N_4327,N_4119,N_4163);
nor U4328 (N_4328,N_4053,N_4034);
and U4329 (N_4329,N_4090,N_4082);
and U4330 (N_4330,N_4195,N_4162);
nor U4331 (N_4331,N_4078,N_4186);
or U4332 (N_4332,N_4121,N_4079);
xnor U4333 (N_4333,N_4053,N_4013);
or U4334 (N_4334,N_4089,N_4183);
or U4335 (N_4335,N_4198,N_4001);
nor U4336 (N_4336,N_4169,N_4092);
and U4337 (N_4337,N_4051,N_4195);
nand U4338 (N_4338,N_4095,N_4168);
nand U4339 (N_4339,N_4138,N_4030);
nor U4340 (N_4340,N_4120,N_4006);
or U4341 (N_4341,N_4013,N_4126);
nor U4342 (N_4342,N_4019,N_4144);
nor U4343 (N_4343,N_4190,N_4100);
nand U4344 (N_4344,N_4057,N_4084);
or U4345 (N_4345,N_4039,N_4057);
and U4346 (N_4346,N_4191,N_4155);
or U4347 (N_4347,N_4189,N_4110);
and U4348 (N_4348,N_4074,N_4048);
nand U4349 (N_4349,N_4128,N_4127);
or U4350 (N_4350,N_4150,N_4017);
nand U4351 (N_4351,N_4173,N_4002);
or U4352 (N_4352,N_4198,N_4117);
and U4353 (N_4353,N_4076,N_4132);
nand U4354 (N_4354,N_4140,N_4096);
or U4355 (N_4355,N_4177,N_4100);
nand U4356 (N_4356,N_4149,N_4187);
nor U4357 (N_4357,N_4199,N_4197);
or U4358 (N_4358,N_4052,N_4049);
and U4359 (N_4359,N_4099,N_4006);
nand U4360 (N_4360,N_4011,N_4069);
xor U4361 (N_4361,N_4016,N_4148);
nor U4362 (N_4362,N_4068,N_4140);
or U4363 (N_4363,N_4199,N_4008);
and U4364 (N_4364,N_4048,N_4166);
xnor U4365 (N_4365,N_4148,N_4086);
nand U4366 (N_4366,N_4026,N_4085);
nand U4367 (N_4367,N_4144,N_4192);
nand U4368 (N_4368,N_4022,N_4015);
or U4369 (N_4369,N_4127,N_4164);
and U4370 (N_4370,N_4190,N_4165);
or U4371 (N_4371,N_4125,N_4070);
and U4372 (N_4372,N_4099,N_4091);
nand U4373 (N_4373,N_4198,N_4133);
nand U4374 (N_4374,N_4017,N_4000);
or U4375 (N_4375,N_4175,N_4130);
nor U4376 (N_4376,N_4124,N_4198);
nand U4377 (N_4377,N_4193,N_4174);
nor U4378 (N_4378,N_4006,N_4045);
or U4379 (N_4379,N_4152,N_4169);
or U4380 (N_4380,N_4198,N_4181);
nand U4381 (N_4381,N_4051,N_4103);
nand U4382 (N_4382,N_4183,N_4072);
and U4383 (N_4383,N_4196,N_4125);
nand U4384 (N_4384,N_4126,N_4029);
nand U4385 (N_4385,N_4061,N_4134);
nand U4386 (N_4386,N_4027,N_4134);
xnor U4387 (N_4387,N_4064,N_4012);
or U4388 (N_4388,N_4099,N_4165);
nand U4389 (N_4389,N_4116,N_4079);
nor U4390 (N_4390,N_4051,N_4007);
nand U4391 (N_4391,N_4053,N_4004);
or U4392 (N_4392,N_4090,N_4050);
nand U4393 (N_4393,N_4043,N_4057);
nor U4394 (N_4394,N_4127,N_4144);
nand U4395 (N_4395,N_4002,N_4121);
or U4396 (N_4396,N_4021,N_4169);
or U4397 (N_4397,N_4156,N_4151);
nor U4398 (N_4398,N_4101,N_4045);
nand U4399 (N_4399,N_4068,N_4032);
and U4400 (N_4400,N_4306,N_4287);
nor U4401 (N_4401,N_4229,N_4203);
nor U4402 (N_4402,N_4207,N_4323);
and U4403 (N_4403,N_4208,N_4277);
or U4404 (N_4404,N_4386,N_4272);
nor U4405 (N_4405,N_4397,N_4224);
nand U4406 (N_4406,N_4248,N_4374);
or U4407 (N_4407,N_4250,N_4362);
and U4408 (N_4408,N_4202,N_4241);
nor U4409 (N_4409,N_4266,N_4271);
nand U4410 (N_4410,N_4315,N_4261);
and U4411 (N_4411,N_4210,N_4331);
nand U4412 (N_4412,N_4398,N_4347);
or U4413 (N_4413,N_4392,N_4371);
and U4414 (N_4414,N_4249,N_4256);
and U4415 (N_4415,N_4201,N_4235);
nand U4416 (N_4416,N_4239,N_4304);
or U4417 (N_4417,N_4290,N_4303);
or U4418 (N_4418,N_4321,N_4291);
nand U4419 (N_4419,N_4377,N_4330);
and U4420 (N_4420,N_4262,N_4237);
and U4421 (N_4421,N_4285,N_4369);
nor U4422 (N_4422,N_4310,N_4360);
or U4423 (N_4423,N_4329,N_4276);
nand U4424 (N_4424,N_4282,N_4351);
nand U4425 (N_4425,N_4218,N_4376);
nand U4426 (N_4426,N_4288,N_4200);
or U4427 (N_4427,N_4375,N_4220);
and U4428 (N_4428,N_4343,N_4283);
nor U4429 (N_4429,N_4252,N_4251);
and U4430 (N_4430,N_4223,N_4381);
and U4431 (N_4431,N_4242,N_4278);
xnor U4432 (N_4432,N_4380,N_4348);
or U4433 (N_4433,N_4358,N_4359);
nand U4434 (N_4434,N_4316,N_4257);
and U4435 (N_4435,N_4357,N_4391);
or U4436 (N_4436,N_4260,N_4268);
nor U4437 (N_4437,N_4286,N_4246);
or U4438 (N_4438,N_4205,N_4294);
and U4439 (N_4439,N_4300,N_4390);
and U4440 (N_4440,N_4225,N_4355);
or U4441 (N_4441,N_4267,N_4314);
nand U4442 (N_4442,N_4356,N_4211);
nand U4443 (N_4443,N_4372,N_4270);
or U4444 (N_4444,N_4297,N_4245);
and U4445 (N_4445,N_4247,N_4240);
or U4446 (N_4446,N_4309,N_4346);
and U4447 (N_4447,N_4382,N_4269);
nand U4448 (N_4448,N_4335,N_4216);
or U4449 (N_4449,N_4212,N_4365);
nand U4450 (N_4450,N_4292,N_4263);
xor U4451 (N_4451,N_4339,N_4336);
or U4452 (N_4452,N_4293,N_4325);
nand U4453 (N_4453,N_4363,N_4354);
and U4454 (N_4454,N_4384,N_4228);
or U4455 (N_4455,N_4279,N_4280);
nor U4456 (N_4456,N_4222,N_4264);
and U4457 (N_4457,N_4296,N_4299);
and U4458 (N_4458,N_4319,N_4206);
and U4459 (N_4459,N_4385,N_4328);
nand U4460 (N_4460,N_4243,N_4298);
nand U4461 (N_4461,N_4253,N_4281);
and U4462 (N_4462,N_4289,N_4295);
nand U4463 (N_4463,N_4259,N_4318);
nor U4464 (N_4464,N_4204,N_4366);
nand U4465 (N_4465,N_4236,N_4396);
and U4466 (N_4466,N_4349,N_4320);
and U4467 (N_4467,N_4341,N_4244);
nor U4468 (N_4468,N_4344,N_4361);
or U4469 (N_4469,N_4227,N_4233);
nor U4470 (N_4470,N_4333,N_4234);
nand U4471 (N_4471,N_4393,N_4373);
nand U4472 (N_4472,N_4322,N_4327);
nor U4473 (N_4473,N_4345,N_4395);
and U4474 (N_4474,N_4352,N_4340);
nand U4475 (N_4475,N_4367,N_4302);
nor U4476 (N_4476,N_4238,N_4312);
or U4477 (N_4477,N_4275,N_4338);
and U4478 (N_4478,N_4274,N_4337);
nor U4479 (N_4479,N_4364,N_4326);
or U4480 (N_4480,N_4383,N_4213);
and U4481 (N_4481,N_4370,N_4209);
and U4482 (N_4482,N_4353,N_4307);
or U4483 (N_4483,N_4389,N_4214);
or U4484 (N_4484,N_4231,N_4265);
nand U4485 (N_4485,N_4368,N_4378);
or U4486 (N_4486,N_4215,N_4388);
and U4487 (N_4487,N_4379,N_4254);
and U4488 (N_4488,N_4273,N_4399);
or U4489 (N_4489,N_4394,N_4308);
and U4490 (N_4490,N_4387,N_4342);
and U4491 (N_4491,N_4334,N_4217);
and U4492 (N_4492,N_4258,N_4350);
and U4493 (N_4493,N_4324,N_4317);
nand U4494 (N_4494,N_4226,N_4305);
nor U4495 (N_4495,N_4311,N_4284);
nand U4496 (N_4496,N_4332,N_4221);
and U4497 (N_4497,N_4230,N_4219);
nand U4498 (N_4498,N_4313,N_4232);
or U4499 (N_4499,N_4301,N_4255);
or U4500 (N_4500,N_4308,N_4226);
nand U4501 (N_4501,N_4335,N_4238);
and U4502 (N_4502,N_4348,N_4320);
and U4503 (N_4503,N_4330,N_4318);
nor U4504 (N_4504,N_4282,N_4226);
nor U4505 (N_4505,N_4374,N_4238);
nor U4506 (N_4506,N_4287,N_4301);
or U4507 (N_4507,N_4335,N_4215);
nor U4508 (N_4508,N_4288,N_4316);
nor U4509 (N_4509,N_4318,N_4258);
nor U4510 (N_4510,N_4205,N_4313);
or U4511 (N_4511,N_4370,N_4211);
nor U4512 (N_4512,N_4371,N_4320);
nor U4513 (N_4513,N_4300,N_4234);
and U4514 (N_4514,N_4243,N_4341);
nor U4515 (N_4515,N_4387,N_4348);
nand U4516 (N_4516,N_4312,N_4371);
xor U4517 (N_4517,N_4324,N_4310);
and U4518 (N_4518,N_4274,N_4321);
nor U4519 (N_4519,N_4286,N_4275);
or U4520 (N_4520,N_4285,N_4220);
nand U4521 (N_4521,N_4309,N_4319);
and U4522 (N_4522,N_4373,N_4270);
or U4523 (N_4523,N_4359,N_4246);
or U4524 (N_4524,N_4314,N_4318);
and U4525 (N_4525,N_4396,N_4219);
nand U4526 (N_4526,N_4216,N_4298);
nor U4527 (N_4527,N_4223,N_4392);
or U4528 (N_4528,N_4320,N_4262);
or U4529 (N_4529,N_4273,N_4233);
nor U4530 (N_4530,N_4222,N_4256);
nand U4531 (N_4531,N_4220,N_4371);
or U4532 (N_4532,N_4252,N_4379);
nand U4533 (N_4533,N_4337,N_4391);
nand U4534 (N_4534,N_4316,N_4239);
nand U4535 (N_4535,N_4278,N_4239);
nand U4536 (N_4536,N_4229,N_4399);
or U4537 (N_4537,N_4389,N_4204);
or U4538 (N_4538,N_4309,N_4307);
or U4539 (N_4539,N_4283,N_4316);
nor U4540 (N_4540,N_4333,N_4373);
and U4541 (N_4541,N_4233,N_4339);
nand U4542 (N_4542,N_4245,N_4291);
and U4543 (N_4543,N_4382,N_4278);
and U4544 (N_4544,N_4282,N_4270);
or U4545 (N_4545,N_4301,N_4290);
nor U4546 (N_4546,N_4352,N_4299);
and U4547 (N_4547,N_4313,N_4375);
or U4548 (N_4548,N_4266,N_4321);
nand U4549 (N_4549,N_4281,N_4325);
nand U4550 (N_4550,N_4243,N_4279);
and U4551 (N_4551,N_4374,N_4223);
nor U4552 (N_4552,N_4307,N_4398);
nor U4553 (N_4553,N_4263,N_4274);
or U4554 (N_4554,N_4326,N_4315);
nor U4555 (N_4555,N_4220,N_4328);
or U4556 (N_4556,N_4244,N_4201);
or U4557 (N_4557,N_4390,N_4366);
nor U4558 (N_4558,N_4238,N_4274);
nand U4559 (N_4559,N_4366,N_4253);
nand U4560 (N_4560,N_4216,N_4340);
nand U4561 (N_4561,N_4230,N_4228);
nor U4562 (N_4562,N_4329,N_4304);
and U4563 (N_4563,N_4295,N_4221);
nand U4564 (N_4564,N_4273,N_4332);
nand U4565 (N_4565,N_4204,N_4222);
and U4566 (N_4566,N_4211,N_4392);
nor U4567 (N_4567,N_4365,N_4254);
and U4568 (N_4568,N_4321,N_4262);
or U4569 (N_4569,N_4373,N_4252);
nor U4570 (N_4570,N_4308,N_4347);
or U4571 (N_4571,N_4365,N_4302);
and U4572 (N_4572,N_4217,N_4307);
nor U4573 (N_4573,N_4328,N_4338);
nand U4574 (N_4574,N_4324,N_4244);
nor U4575 (N_4575,N_4234,N_4388);
and U4576 (N_4576,N_4239,N_4384);
nand U4577 (N_4577,N_4213,N_4390);
nor U4578 (N_4578,N_4202,N_4346);
nand U4579 (N_4579,N_4217,N_4387);
nor U4580 (N_4580,N_4224,N_4254);
or U4581 (N_4581,N_4235,N_4218);
nand U4582 (N_4582,N_4271,N_4368);
nor U4583 (N_4583,N_4360,N_4263);
nand U4584 (N_4584,N_4285,N_4248);
or U4585 (N_4585,N_4229,N_4244);
and U4586 (N_4586,N_4279,N_4251);
and U4587 (N_4587,N_4314,N_4282);
and U4588 (N_4588,N_4326,N_4207);
xor U4589 (N_4589,N_4377,N_4214);
or U4590 (N_4590,N_4368,N_4374);
or U4591 (N_4591,N_4211,N_4367);
and U4592 (N_4592,N_4322,N_4216);
and U4593 (N_4593,N_4254,N_4302);
nand U4594 (N_4594,N_4313,N_4341);
and U4595 (N_4595,N_4381,N_4263);
nor U4596 (N_4596,N_4234,N_4305);
or U4597 (N_4597,N_4324,N_4212);
and U4598 (N_4598,N_4394,N_4383);
nor U4599 (N_4599,N_4376,N_4372);
or U4600 (N_4600,N_4536,N_4596);
nor U4601 (N_4601,N_4438,N_4533);
nand U4602 (N_4602,N_4440,N_4535);
or U4603 (N_4603,N_4578,N_4503);
xor U4604 (N_4604,N_4589,N_4484);
nand U4605 (N_4605,N_4584,N_4416);
nand U4606 (N_4606,N_4467,N_4412);
and U4607 (N_4607,N_4481,N_4498);
nor U4608 (N_4608,N_4453,N_4552);
nor U4609 (N_4609,N_4555,N_4465);
or U4610 (N_4610,N_4472,N_4441);
and U4611 (N_4611,N_4486,N_4421);
and U4612 (N_4612,N_4537,N_4435);
nor U4613 (N_4613,N_4418,N_4575);
nor U4614 (N_4614,N_4424,N_4475);
nand U4615 (N_4615,N_4574,N_4415);
nand U4616 (N_4616,N_4500,N_4429);
and U4617 (N_4617,N_4591,N_4501);
nor U4618 (N_4618,N_4433,N_4420);
and U4619 (N_4619,N_4518,N_4470);
or U4620 (N_4620,N_4547,N_4557);
nand U4621 (N_4621,N_4478,N_4595);
and U4622 (N_4622,N_4431,N_4479);
nor U4623 (N_4623,N_4492,N_4567);
xnor U4624 (N_4624,N_4411,N_4570);
or U4625 (N_4625,N_4593,N_4585);
nor U4626 (N_4626,N_4491,N_4464);
and U4627 (N_4627,N_4462,N_4451);
nand U4628 (N_4628,N_4563,N_4507);
or U4629 (N_4629,N_4520,N_4597);
and U4630 (N_4630,N_4408,N_4572);
and U4631 (N_4631,N_4490,N_4587);
nor U4632 (N_4632,N_4443,N_4571);
or U4633 (N_4633,N_4410,N_4454);
and U4634 (N_4634,N_4519,N_4581);
or U4635 (N_4635,N_4532,N_4414);
nand U4636 (N_4636,N_4588,N_4471);
nor U4637 (N_4637,N_4524,N_4437);
or U4638 (N_4638,N_4599,N_4510);
nand U4639 (N_4639,N_4447,N_4526);
and U4640 (N_4640,N_4497,N_4487);
nand U4641 (N_4641,N_4564,N_4521);
nand U4642 (N_4642,N_4534,N_4566);
nor U4643 (N_4643,N_4463,N_4565);
nor U4644 (N_4644,N_4523,N_4458);
nand U4645 (N_4645,N_4460,N_4419);
nor U4646 (N_4646,N_4541,N_4577);
nor U4647 (N_4647,N_4488,N_4407);
or U4648 (N_4648,N_4530,N_4413);
or U4649 (N_4649,N_4461,N_4469);
or U4650 (N_4650,N_4556,N_4423);
nand U4651 (N_4651,N_4402,N_4540);
and U4652 (N_4652,N_4445,N_4502);
nor U4653 (N_4653,N_4442,N_4505);
or U4654 (N_4654,N_4549,N_4562);
or U4655 (N_4655,N_4425,N_4450);
and U4656 (N_4656,N_4405,N_4427);
or U4657 (N_4657,N_4456,N_4553);
or U4658 (N_4658,N_4485,N_4582);
nand U4659 (N_4659,N_4494,N_4544);
nor U4660 (N_4660,N_4531,N_4506);
or U4661 (N_4661,N_4417,N_4516);
or U4662 (N_4662,N_4558,N_4546);
nor U4663 (N_4663,N_4569,N_4576);
or U4664 (N_4664,N_4551,N_4430);
nand U4665 (N_4665,N_4493,N_4468);
nand U4666 (N_4666,N_4449,N_4439);
nor U4667 (N_4667,N_4432,N_4580);
and U4668 (N_4668,N_4592,N_4509);
or U4669 (N_4669,N_4400,N_4586);
and U4670 (N_4670,N_4543,N_4538);
or U4671 (N_4671,N_4579,N_4446);
nor U4672 (N_4672,N_4448,N_4560);
nand U4673 (N_4673,N_4550,N_4404);
nor U4674 (N_4674,N_4517,N_4426);
nor U4675 (N_4675,N_4554,N_4466);
nor U4676 (N_4676,N_4545,N_4422);
and U4677 (N_4677,N_4406,N_4511);
and U4678 (N_4678,N_4594,N_4409);
nand U4679 (N_4679,N_4434,N_4473);
or U4680 (N_4680,N_4573,N_4598);
or U4681 (N_4681,N_4444,N_4499);
nand U4682 (N_4682,N_4527,N_4496);
or U4683 (N_4683,N_4539,N_4559);
nand U4684 (N_4684,N_4568,N_4401);
nor U4685 (N_4685,N_4513,N_4590);
nor U4686 (N_4686,N_4403,N_4477);
and U4687 (N_4687,N_4480,N_4495);
and U4688 (N_4688,N_4457,N_4561);
nand U4689 (N_4689,N_4548,N_4476);
nand U4690 (N_4690,N_4528,N_4508);
or U4691 (N_4691,N_4474,N_4504);
nand U4692 (N_4692,N_4515,N_4482);
nand U4693 (N_4693,N_4512,N_4529);
or U4694 (N_4694,N_4583,N_4459);
or U4695 (N_4695,N_4522,N_4436);
or U4696 (N_4696,N_4514,N_4525);
or U4697 (N_4697,N_4455,N_4483);
nor U4698 (N_4698,N_4489,N_4452);
and U4699 (N_4699,N_4428,N_4542);
nand U4700 (N_4700,N_4512,N_4572);
nor U4701 (N_4701,N_4560,N_4557);
and U4702 (N_4702,N_4570,N_4429);
nor U4703 (N_4703,N_4476,N_4529);
or U4704 (N_4704,N_4494,N_4597);
and U4705 (N_4705,N_4538,N_4460);
nor U4706 (N_4706,N_4578,N_4439);
and U4707 (N_4707,N_4503,N_4411);
or U4708 (N_4708,N_4589,N_4428);
and U4709 (N_4709,N_4584,N_4468);
or U4710 (N_4710,N_4400,N_4585);
nor U4711 (N_4711,N_4449,N_4524);
and U4712 (N_4712,N_4469,N_4531);
nor U4713 (N_4713,N_4418,N_4450);
nand U4714 (N_4714,N_4536,N_4462);
nand U4715 (N_4715,N_4419,N_4523);
nor U4716 (N_4716,N_4447,N_4584);
nor U4717 (N_4717,N_4568,N_4436);
nand U4718 (N_4718,N_4598,N_4599);
nand U4719 (N_4719,N_4433,N_4562);
nand U4720 (N_4720,N_4548,N_4494);
and U4721 (N_4721,N_4489,N_4478);
nor U4722 (N_4722,N_4407,N_4439);
nor U4723 (N_4723,N_4482,N_4565);
nor U4724 (N_4724,N_4456,N_4439);
nor U4725 (N_4725,N_4519,N_4412);
nand U4726 (N_4726,N_4507,N_4535);
nor U4727 (N_4727,N_4540,N_4565);
and U4728 (N_4728,N_4445,N_4539);
nand U4729 (N_4729,N_4559,N_4508);
or U4730 (N_4730,N_4463,N_4505);
xnor U4731 (N_4731,N_4523,N_4405);
or U4732 (N_4732,N_4541,N_4453);
nor U4733 (N_4733,N_4540,N_4556);
or U4734 (N_4734,N_4518,N_4503);
or U4735 (N_4735,N_4527,N_4562);
or U4736 (N_4736,N_4512,N_4481);
and U4737 (N_4737,N_4513,N_4580);
and U4738 (N_4738,N_4547,N_4587);
or U4739 (N_4739,N_4589,N_4556);
or U4740 (N_4740,N_4429,N_4418);
nor U4741 (N_4741,N_4544,N_4420);
nand U4742 (N_4742,N_4506,N_4417);
xnor U4743 (N_4743,N_4479,N_4521);
or U4744 (N_4744,N_4460,N_4491);
nand U4745 (N_4745,N_4597,N_4528);
nand U4746 (N_4746,N_4534,N_4549);
and U4747 (N_4747,N_4525,N_4421);
nand U4748 (N_4748,N_4425,N_4512);
and U4749 (N_4749,N_4599,N_4497);
nand U4750 (N_4750,N_4498,N_4406);
nor U4751 (N_4751,N_4541,N_4438);
nand U4752 (N_4752,N_4571,N_4466);
or U4753 (N_4753,N_4450,N_4525);
nand U4754 (N_4754,N_4540,N_4466);
or U4755 (N_4755,N_4433,N_4530);
nor U4756 (N_4756,N_4451,N_4509);
and U4757 (N_4757,N_4485,N_4546);
or U4758 (N_4758,N_4531,N_4501);
xor U4759 (N_4759,N_4437,N_4420);
and U4760 (N_4760,N_4563,N_4453);
nand U4761 (N_4761,N_4457,N_4527);
or U4762 (N_4762,N_4446,N_4503);
or U4763 (N_4763,N_4524,N_4484);
and U4764 (N_4764,N_4441,N_4413);
or U4765 (N_4765,N_4592,N_4581);
nor U4766 (N_4766,N_4576,N_4597);
nor U4767 (N_4767,N_4463,N_4489);
nor U4768 (N_4768,N_4505,N_4467);
and U4769 (N_4769,N_4472,N_4560);
and U4770 (N_4770,N_4498,N_4457);
nor U4771 (N_4771,N_4534,N_4548);
or U4772 (N_4772,N_4533,N_4467);
nor U4773 (N_4773,N_4590,N_4534);
or U4774 (N_4774,N_4493,N_4457);
and U4775 (N_4775,N_4580,N_4504);
and U4776 (N_4776,N_4467,N_4482);
or U4777 (N_4777,N_4497,N_4414);
or U4778 (N_4778,N_4542,N_4481);
or U4779 (N_4779,N_4538,N_4427);
nor U4780 (N_4780,N_4439,N_4568);
or U4781 (N_4781,N_4455,N_4496);
or U4782 (N_4782,N_4557,N_4531);
or U4783 (N_4783,N_4589,N_4449);
or U4784 (N_4784,N_4471,N_4487);
and U4785 (N_4785,N_4444,N_4544);
nand U4786 (N_4786,N_4412,N_4457);
or U4787 (N_4787,N_4477,N_4485);
nor U4788 (N_4788,N_4479,N_4434);
nand U4789 (N_4789,N_4416,N_4526);
nor U4790 (N_4790,N_4447,N_4537);
xnor U4791 (N_4791,N_4457,N_4402);
and U4792 (N_4792,N_4553,N_4592);
nor U4793 (N_4793,N_4489,N_4566);
nand U4794 (N_4794,N_4589,N_4547);
and U4795 (N_4795,N_4527,N_4440);
nor U4796 (N_4796,N_4573,N_4580);
or U4797 (N_4797,N_4523,N_4591);
nor U4798 (N_4798,N_4584,N_4493);
nand U4799 (N_4799,N_4518,N_4560);
nor U4800 (N_4800,N_4762,N_4712);
nor U4801 (N_4801,N_4789,N_4636);
nor U4802 (N_4802,N_4691,N_4765);
and U4803 (N_4803,N_4783,N_4781);
or U4804 (N_4804,N_4787,N_4736);
or U4805 (N_4805,N_4779,N_4650);
and U4806 (N_4806,N_4686,N_4788);
or U4807 (N_4807,N_4600,N_4729);
nor U4808 (N_4808,N_4611,N_4782);
nand U4809 (N_4809,N_4606,N_4692);
nor U4810 (N_4810,N_4718,N_4746);
and U4811 (N_4811,N_4733,N_4610);
or U4812 (N_4812,N_4613,N_4726);
or U4813 (N_4813,N_4674,N_4740);
nand U4814 (N_4814,N_4696,N_4637);
nor U4815 (N_4815,N_4678,N_4688);
and U4816 (N_4816,N_4615,N_4685);
or U4817 (N_4817,N_4748,N_4679);
and U4818 (N_4818,N_4651,N_4622);
nor U4819 (N_4819,N_4794,N_4628);
and U4820 (N_4820,N_4675,N_4668);
nand U4821 (N_4821,N_4671,N_4724);
nor U4822 (N_4822,N_4723,N_4784);
nor U4823 (N_4823,N_4728,N_4609);
nor U4824 (N_4824,N_4705,N_4706);
xor U4825 (N_4825,N_4639,N_4629);
and U4826 (N_4826,N_4796,N_4632);
nor U4827 (N_4827,N_4713,N_4774);
nand U4828 (N_4828,N_4722,N_4754);
or U4829 (N_4829,N_4742,N_4658);
nor U4830 (N_4830,N_4601,N_4631);
or U4831 (N_4831,N_4730,N_4607);
or U4832 (N_4832,N_4618,N_4614);
or U4833 (N_4833,N_4743,N_4753);
and U4834 (N_4834,N_4707,N_4769);
and U4835 (N_4835,N_4654,N_4702);
or U4836 (N_4836,N_4752,N_4662);
nor U4837 (N_4837,N_4719,N_4786);
nand U4838 (N_4838,N_4776,N_4791);
or U4839 (N_4839,N_4777,N_4709);
or U4840 (N_4840,N_4683,N_4672);
nor U4841 (N_4841,N_4612,N_4626);
or U4842 (N_4842,N_4715,N_4649);
and U4843 (N_4843,N_4655,N_4701);
nor U4844 (N_4844,N_4703,N_4656);
nor U4845 (N_4845,N_4682,N_4760);
or U4846 (N_4846,N_4633,N_4623);
or U4847 (N_4847,N_4771,N_4714);
or U4848 (N_4848,N_4694,N_4697);
nor U4849 (N_4849,N_4670,N_4751);
xor U4850 (N_4850,N_4602,N_4604);
nand U4851 (N_4851,N_4745,N_4763);
nor U4852 (N_4852,N_4663,N_4664);
or U4853 (N_4853,N_4711,N_4641);
or U4854 (N_4854,N_4665,N_4620);
or U4855 (N_4855,N_4652,N_4681);
or U4856 (N_4856,N_4644,N_4687);
nand U4857 (N_4857,N_4755,N_4630);
and U4858 (N_4858,N_4608,N_4756);
and U4859 (N_4859,N_4677,N_4661);
xnor U4860 (N_4860,N_4770,N_4699);
and U4861 (N_4861,N_4780,N_4695);
nand U4862 (N_4862,N_4721,N_4739);
or U4863 (N_4863,N_4737,N_4727);
nand U4864 (N_4864,N_4792,N_4634);
nand U4865 (N_4865,N_4619,N_4627);
nand U4866 (N_4866,N_4741,N_4772);
and U4867 (N_4867,N_4605,N_4645);
or U4868 (N_4868,N_4625,N_4759);
nand U4869 (N_4869,N_4635,N_4708);
or U4870 (N_4870,N_4640,N_4775);
nand U4871 (N_4871,N_4725,N_4716);
nor U4872 (N_4872,N_4710,N_4738);
nor U4873 (N_4873,N_4747,N_4750);
or U4874 (N_4874,N_4616,N_4793);
or U4875 (N_4875,N_4698,N_4621);
nand U4876 (N_4876,N_4704,N_4660);
nand U4877 (N_4877,N_4790,N_4617);
or U4878 (N_4878,N_4744,N_4799);
nor U4879 (N_4879,N_4768,N_4732);
nand U4880 (N_4880,N_4758,N_4603);
xnor U4881 (N_4881,N_4659,N_4638);
nand U4882 (N_4882,N_4657,N_4735);
and U4883 (N_4883,N_4767,N_4643);
nand U4884 (N_4884,N_4693,N_4761);
and U4885 (N_4885,N_4720,N_4731);
and U4886 (N_4886,N_4797,N_4764);
and U4887 (N_4887,N_4773,N_4673);
or U4888 (N_4888,N_4690,N_4795);
nor U4889 (N_4889,N_4798,N_4684);
or U4890 (N_4890,N_4680,N_4666);
nor U4891 (N_4891,N_4717,N_4647);
nand U4892 (N_4892,N_4646,N_4653);
nor U4893 (N_4893,N_4667,N_4689);
nor U4894 (N_4894,N_4778,N_4757);
nor U4895 (N_4895,N_4766,N_4669);
and U4896 (N_4896,N_4642,N_4676);
nor U4897 (N_4897,N_4648,N_4624);
or U4898 (N_4898,N_4700,N_4749);
and U4899 (N_4899,N_4785,N_4734);
nor U4900 (N_4900,N_4775,N_4783);
and U4901 (N_4901,N_4714,N_4667);
or U4902 (N_4902,N_4745,N_4746);
and U4903 (N_4903,N_4651,N_4646);
or U4904 (N_4904,N_4794,N_4799);
or U4905 (N_4905,N_4733,N_4786);
nand U4906 (N_4906,N_4776,N_4603);
nand U4907 (N_4907,N_4638,N_4615);
nor U4908 (N_4908,N_4604,N_4700);
nor U4909 (N_4909,N_4622,N_4797);
nand U4910 (N_4910,N_4670,N_4722);
nand U4911 (N_4911,N_4731,N_4680);
and U4912 (N_4912,N_4774,N_4766);
nand U4913 (N_4913,N_4753,N_4769);
and U4914 (N_4914,N_4637,N_4764);
or U4915 (N_4915,N_4678,N_4797);
and U4916 (N_4916,N_4611,N_4731);
or U4917 (N_4917,N_4600,N_4618);
or U4918 (N_4918,N_4763,N_4795);
nand U4919 (N_4919,N_4689,N_4722);
nor U4920 (N_4920,N_4622,N_4703);
and U4921 (N_4921,N_4610,N_4683);
nand U4922 (N_4922,N_4778,N_4712);
or U4923 (N_4923,N_4677,N_4667);
and U4924 (N_4924,N_4755,N_4646);
or U4925 (N_4925,N_4620,N_4631);
or U4926 (N_4926,N_4650,N_4752);
and U4927 (N_4927,N_4790,N_4601);
nand U4928 (N_4928,N_4629,N_4606);
and U4929 (N_4929,N_4720,N_4642);
nand U4930 (N_4930,N_4692,N_4688);
nor U4931 (N_4931,N_4676,N_4640);
nand U4932 (N_4932,N_4647,N_4738);
nor U4933 (N_4933,N_4631,N_4713);
or U4934 (N_4934,N_4787,N_4746);
or U4935 (N_4935,N_4600,N_4662);
nand U4936 (N_4936,N_4717,N_4616);
or U4937 (N_4937,N_4648,N_4700);
nand U4938 (N_4938,N_4730,N_4761);
nor U4939 (N_4939,N_4628,N_4773);
nor U4940 (N_4940,N_4649,N_4759);
or U4941 (N_4941,N_4625,N_4624);
or U4942 (N_4942,N_4715,N_4642);
and U4943 (N_4943,N_4713,N_4764);
nand U4944 (N_4944,N_4757,N_4743);
nand U4945 (N_4945,N_4726,N_4795);
and U4946 (N_4946,N_4779,N_4682);
nor U4947 (N_4947,N_4634,N_4615);
or U4948 (N_4948,N_4660,N_4714);
nor U4949 (N_4949,N_4747,N_4781);
and U4950 (N_4950,N_4666,N_4609);
or U4951 (N_4951,N_4748,N_4623);
nor U4952 (N_4952,N_4618,N_4631);
and U4953 (N_4953,N_4780,N_4766);
and U4954 (N_4954,N_4734,N_4740);
or U4955 (N_4955,N_4664,N_4654);
or U4956 (N_4956,N_4680,N_4632);
and U4957 (N_4957,N_4650,N_4727);
nand U4958 (N_4958,N_4603,N_4684);
nand U4959 (N_4959,N_4755,N_4751);
and U4960 (N_4960,N_4763,N_4619);
nand U4961 (N_4961,N_4722,N_4668);
or U4962 (N_4962,N_4742,N_4677);
nor U4963 (N_4963,N_4799,N_4708);
nand U4964 (N_4964,N_4674,N_4698);
and U4965 (N_4965,N_4630,N_4736);
nand U4966 (N_4966,N_4671,N_4694);
xnor U4967 (N_4967,N_4606,N_4632);
nand U4968 (N_4968,N_4675,N_4759);
or U4969 (N_4969,N_4615,N_4723);
nand U4970 (N_4970,N_4755,N_4610);
nand U4971 (N_4971,N_4684,N_4682);
or U4972 (N_4972,N_4696,N_4671);
nand U4973 (N_4973,N_4764,N_4620);
and U4974 (N_4974,N_4747,N_4757);
and U4975 (N_4975,N_4740,N_4736);
nor U4976 (N_4976,N_4672,N_4692);
and U4977 (N_4977,N_4634,N_4716);
and U4978 (N_4978,N_4672,N_4746);
nand U4979 (N_4979,N_4675,N_4793);
nor U4980 (N_4980,N_4743,N_4607);
nor U4981 (N_4981,N_4772,N_4718);
nand U4982 (N_4982,N_4715,N_4764);
nor U4983 (N_4983,N_4643,N_4636);
nor U4984 (N_4984,N_4666,N_4739);
xor U4985 (N_4985,N_4774,N_4652);
or U4986 (N_4986,N_4782,N_4773);
and U4987 (N_4987,N_4742,N_4792);
and U4988 (N_4988,N_4769,N_4612);
or U4989 (N_4989,N_4622,N_4672);
and U4990 (N_4990,N_4645,N_4647);
and U4991 (N_4991,N_4710,N_4621);
or U4992 (N_4992,N_4611,N_4762);
or U4993 (N_4993,N_4796,N_4665);
nor U4994 (N_4994,N_4682,N_4743);
or U4995 (N_4995,N_4683,N_4780);
nor U4996 (N_4996,N_4792,N_4686);
or U4997 (N_4997,N_4716,N_4683);
nor U4998 (N_4998,N_4734,N_4654);
nand U4999 (N_4999,N_4787,N_4721);
xor U5000 (N_5000,N_4921,N_4967);
nand U5001 (N_5001,N_4824,N_4929);
nor U5002 (N_5002,N_4831,N_4946);
and U5003 (N_5003,N_4807,N_4907);
or U5004 (N_5004,N_4943,N_4920);
nand U5005 (N_5005,N_4965,N_4873);
or U5006 (N_5006,N_4995,N_4811);
nand U5007 (N_5007,N_4924,N_4992);
or U5008 (N_5008,N_4996,N_4903);
nand U5009 (N_5009,N_4949,N_4945);
nand U5010 (N_5010,N_4969,N_4951);
and U5011 (N_5011,N_4880,N_4874);
nand U5012 (N_5012,N_4863,N_4820);
nand U5013 (N_5013,N_4941,N_4974);
nor U5014 (N_5014,N_4970,N_4866);
nor U5015 (N_5015,N_4844,N_4812);
and U5016 (N_5016,N_4817,N_4832);
nand U5017 (N_5017,N_4876,N_4892);
nor U5018 (N_5018,N_4814,N_4872);
or U5019 (N_5019,N_4914,N_4955);
nor U5020 (N_5020,N_4890,N_4870);
and U5021 (N_5021,N_4985,N_4956);
nand U5022 (N_5022,N_4917,N_4853);
and U5023 (N_5023,N_4815,N_4854);
nor U5024 (N_5024,N_4942,N_4984);
or U5025 (N_5025,N_4954,N_4958);
and U5026 (N_5026,N_4825,N_4983);
or U5027 (N_5027,N_4861,N_4862);
nor U5028 (N_5028,N_4897,N_4804);
and U5029 (N_5029,N_4833,N_4808);
or U5030 (N_5030,N_4961,N_4912);
and U5031 (N_5031,N_4837,N_4971);
and U5032 (N_5032,N_4898,N_4911);
or U5033 (N_5033,N_4979,N_4909);
nor U5034 (N_5034,N_4968,N_4895);
nand U5035 (N_5035,N_4998,N_4926);
nor U5036 (N_5036,N_4978,N_4973);
nand U5037 (N_5037,N_4855,N_4959);
and U5038 (N_5038,N_4997,N_4972);
or U5039 (N_5039,N_4875,N_4902);
or U5040 (N_5040,N_4850,N_4852);
and U5041 (N_5041,N_4830,N_4927);
and U5042 (N_5042,N_4806,N_4802);
or U5043 (N_5043,N_4868,N_4809);
nand U5044 (N_5044,N_4883,N_4933);
and U5045 (N_5045,N_4800,N_4988);
nor U5046 (N_5046,N_4935,N_4887);
nand U5047 (N_5047,N_4847,N_4915);
or U5048 (N_5048,N_4828,N_4953);
nand U5049 (N_5049,N_4893,N_4991);
or U5050 (N_5050,N_4841,N_4950);
or U5051 (N_5051,N_4987,N_4928);
nor U5052 (N_5052,N_4981,N_4993);
and U5053 (N_5053,N_4835,N_4846);
nor U5054 (N_5054,N_4905,N_4931);
xor U5055 (N_5055,N_4816,N_4947);
and U5056 (N_5056,N_4878,N_4840);
or U5057 (N_5057,N_4843,N_4857);
nand U5058 (N_5058,N_4813,N_4869);
or U5059 (N_5059,N_4960,N_4877);
xor U5060 (N_5060,N_4856,N_4910);
and U5061 (N_5061,N_4975,N_4901);
nor U5062 (N_5062,N_4925,N_4936);
nor U5063 (N_5063,N_4989,N_4952);
nand U5064 (N_5064,N_4836,N_4966);
and U5065 (N_5065,N_4906,N_4964);
and U5066 (N_5066,N_4805,N_4999);
nand U5067 (N_5067,N_4919,N_4849);
nor U5068 (N_5068,N_4916,N_4934);
or U5069 (N_5069,N_4818,N_4839);
and U5070 (N_5070,N_4894,N_4930);
or U5071 (N_5071,N_4904,N_4858);
nand U5072 (N_5072,N_4838,N_4939);
or U5073 (N_5073,N_4881,N_4982);
nor U5074 (N_5074,N_4829,N_4994);
nand U5075 (N_5075,N_4908,N_4826);
and U5076 (N_5076,N_4848,N_4819);
nor U5077 (N_5077,N_4823,N_4922);
nor U5078 (N_5078,N_4822,N_4885);
nor U5079 (N_5079,N_4867,N_4938);
and U5080 (N_5080,N_4834,N_4860);
and U5081 (N_5081,N_4882,N_4888);
nand U5082 (N_5082,N_4963,N_4957);
nor U5083 (N_5083,N_4913,N_4821);
or U5084 (N_5084,N_4865,N_4803);
and U5085 (N_5085,N_4948,N_4864);
and U5086 (N_5086,N_4977,N_4879);
nor U5087 (N_5087,N_4801,N_4899);
nand U5088 (N_5088,N_4980,N_4962);
and U5089 (N_5089,N_4944,N_4842);
and U5090 (N_5090,N_4845,N_4827);
nor U5091 (N_5091,N_4990,N_4891);
nor U5092 (N_5092,N_4937,N_4932);
nor U5093 (N_5093,N_4900,N_4886);
and U5094 (N_5094,N_4884,N_4976);
and U5095 (N_5095,N_4851,N_4918);
or U5096 (N_5096,N_4896,N_4940);
nand U5097 (N_5097,N_4871,N_4986);
and U5098 (N_5098,N_4889,N_4810);
nand U5099 (N_5099,N_4923,N_4859);
and U5100 (N_5100,N_4822,N_4938);
nand U5101 (N_5101,N_4807,N_4924);
nand U5102 (N_5102,N_4833,N_4915);
nand U5103 (N_5103,N_4844,N_4962);
and U5104 (N_5104,N_4867,N_4823);
or U5105 (N_5105,N_4854,N_4983);
and U5106 (N_5106,N_4839,N_4802);
nor U5107 (N_5107,N_4932,N_4954);
xnor U5108 (N_5108,N_4887,N_4955);
nor U5109 (N_5109,N_4982,N_4948);
and U5110 (N_5110,N_4856,N_4923);
nor U5111 (N_5111,N_4926,N_4992);
nor U5112 (N_5112,N_4888,N_4955);
nor U5113 (N_5113,N_4941,N_4988);
nor U5114 (N_5114,N_4929,N_4943);
nor U5115 (N_5115,N_4828,N_4913);
nor U5116 (N_5116,N_4997,N_4817);
and U5117 (N_5117,N_4844,N_4972);
or U5118 (N_5118,N_4972,N_4877);
nand U5119 (N_5119,N_4905,N_4947);
and U5120 (N_5120,N_4822,N_4868);
nor U5121 (N_5121,N_4968,N_4924);
and U5122 (N_5122,N_4993,N_4957);
and U5123 (N_5123,N_4880,N_4968);
or U5124 (N_5124,N_4906,N_4883);
nand U5125 (N_5125,N_4807,N_4896);
and U5126 (N_5126,N_4901,N_4910);
nor U5127 (N_5127,N_4894,N_4876);
or U5128 (N_5128,N_4940,N_4873);
or U5129 (N_5129,N_4850,N_4882);
nor U5130 (N_5130,N_4848,N_4807);
nor U5131 (N_5131,N_4833,N_4870);
nand U5132 (N_5132,N_4841,N_4959);
nand U5133 (N_5133,N_4998,N_4968);
nand U5134 (N_5134,N_4944,N_4943);
or U5135 (N_5135,N_4865,N_4907);
or U5136 (N_5136,N_4915,N_4878);
and U5137 (N_5137,N_4917,N_4885);
nand U5138 (N_5138,N_4824,N_4809);
nor U5139 (N_5139,N_4820,N_4844);
or U5140 (N_5140,N_4882,N_4804);
and U5141 (N_5141,N_4856,N_4959);
or U5142 (N_5142,N_4873,N_4813);
nand U5143 (N_5143,N_4888,N_4831);
nand U5144 (N_5144,N_4816,N_4865);
or U5145 (N_5145,N_4987,N_4980);
or U5146 (N_5146,N_4909,N_4902);
nor U5147 (N_5147,N_4992,N_4989);
or U5148 (N_5148,N_4991,N_4947);
and U5149 (N_5149,N_4811,N_4920);
nor U5150 (N_5150,N_4806,N_4894);
and U5151 (N_5151,N_4982,N_4959);
nor U5152 (N_5152,N_4890,N_4805);
nor U5153 (N_5153,N_4979,N_4833);
and U5154 (N_5154,N_4918,N_4985);
or U5155 (N_5155,N_4868,N_4904);
nand U5156 (N_5156,N_4989,N_4836);
and U5157 (N_5157,N_4852,N_4894);
and U5158 (N_5158,N_4907,N_4876);
nand U5159 (N_5159,N_4847,N_4843);
nor U5160 (N_5160,N_4910,N_4841);
nand U5161 (N_5161,N_4883,N_4858);
nand U5162 (N_5162,N_4927,N_4811);
and U5163 (N_5163,N_4986,N_4976);
and U5164 (N_5164,N_4938,N_4834);
nor U5165 (N_5165,N_4993,N_4842);
nand U5166 (N_5166,N_4995,N_4981);
and U5167 (N_5167,N_4949,N_4893);
nor U5168 (N_5168,N_4887,N_4950);
or U5169 (N_5169,N_4801,N_4958);
nor U5170 (N_5170,N_4867,N_4831);
nor U5171 (N_5171,N_4902,N_4930);
nand U5172 (N_5172,N_4852,N_4937);
nor U5173 (N_5173,N_4996,N_4883);
and U5174 (N_5174,N_4850,N_4977);
or U5175 (N_5175,N_4926,N_4944);
nand U5176 (N_5176,N_4908,N_4993);
or U5177 (N_5177,N_4868,N_4861);
nor U5178 (N_5178,N_4983,N_4866);
nor U5179 (N_5179,N_4979,N_4946);
nor U5180 (N_5180,N_4978,N_4852);
or U5181 (N_5181,N_4963,N_4923);
nor U5182 (N_5182,N_4806,N_4926);
nor U5183 (N_5183,N_4985,N_4982);
nand U5184 (N_5184,N_4837,N_4829);
and U5185 (N_5185,N_4879,N_4903);
and U5186 (N_5186,N_4844,N_4871);
nor U5187 (N_5187,N_4954,N_4900);
and U5188 (N_5188,N_4847,N_4939);
xnor U5189 (N_5189,N_4888,N_4802);
xnor U5190 (N_5190,N_4973,N_4972);
nor U5191 (N_5191,N_4903,N_4999);
nor U5192 (N_5192,N_4964,N_4860);
or U5193 (N_5193,N_4913,N_4959);
or U5194 (N_5194,N_4849,N_4852);
xnor U5195 (N_5195,N_4989,N_4934);
nor U5196 (N_5196,N_4878,N_4990);
nand U5197 (N_5197,N_4983,N_4918);
and U5198 (N_5198,N_4901,N_4866);
nand U5199 (N_5199,N_4919,N_4838);
or U5200 (N_5200,N_5078,N_5100);
and U5201 (N_5201,N_5138,N_5081);
nand U5202 (N_5202,N_5051,N_5110);
or U5203 (N_5203,N_5159,N_5016);
or U5204 (N_5204,N_5152,N_5182);
and U5205 (N_5205,N_5009,N_5140);
and U5206 (N_5206,N_5024,N_5008);
nor U5207 (N_5207,N_5176,N_5064);
nand U5208 (N_5208,N_5005,N_5165);
nand U5209 (N_5209,N_5099,N_5124);
nand U5210 (N_5210,N_5196,N_5119);
nor U5211 (N_5211,N_5158,N_5057);
nand U5212 (N_5212,N_5084,N_5075);
and U5213 (N_5213,N_5076,N_5171);
and U5214 (N_5214,N_5067,N_5028);
or U5215 (N_5215,N_5073,N_5006);
or U5216 (N_5216,N_5166,N_5054);
or U5217 (N_5217,N_5061,N_5040);
or U5218 (N_5218,N_5122,N_5049);
or U5219 (N_5219,N_5121,N_5025);
nor U5220 (N_5220,N_5101,N_5018);
or U5221 (N_5221,N_5037,N_5163);
nor U5222 (N_5222,N_5198,N_5023);
nand U5223 (N_5223,N_5188,N_5120);
and U5224 (N_5224,N_5162,N_5150);
or U5225 (N_5225,N_5131,N_5115);
nor U5226 (N_5226,N_5157,N_5194);
or U5227 (N_5227,N_5034,N_5184);
nand U5228 (N_5228,N_5136,N_5191);
or U5229 (N_5229,N_5145,N_5039);
and U5230 (N_5230,N_5047,N_5086);
and U5231 (N_5231,N_5070,N_5161);
nand U5232 (N_5232,N_5134,N_5192);
nor U5233 (N_5233,N_5117,N_5130);
nand U5234 (N_5234,N_5015,N_5174);
and U5235 (N_5235,N_5126,N_5036);
or U5236 (N_5236,N_5010,N_5017);
and U5237 (N_5237,N_5129,N_5193);
nand U5238 (N_5238,N_5058,N_5048);
or U5239 (N_5239,N_5001,N_5095);
nor U5240 (N_5240,N_5156,N_5183);
nand U5241 (N_5241,N_5180,N_5044);
or U5242 (N_5242,N_5133,N_5170);
and U5243 (N_5243,N_5003,N_5007);
and U5244 (N_5244,N_5060,N_5032);
nand U5245 (N_5245,N_5108,N_5030);
nor U5246 (N_5246,N_5068,N_5189);
nor U5247 (N_5247,N_5022,N_5181);
nand U5248 (N_5248,N_5094,N_5063);
and U5249 (N_5249,N_5069,N_5029);
or U5250 (N_5250,N_5000,N_5045);
nor U5251 (N_5251,N_5185,N_5105);
and U5252 (N_5252,N_5109,N_5195);
or U5253 (N_5253,N_5139,N_5097);
and U5254 (N_5254,N_5096,N_5178);
nand U5255 (N_5255,N_5013,N_5087);
and U5256 (N_5256,N_5125,N_5148);
nand U5257 (N_5257,N_5079,N_5002);
or U5258 (N_5258,N_5026,N_5107);
nor U5259 (N_5259,N_5043,N_5151);
nor U5260 (N_5260,N_5190,N_5197);
and U5261 (N_5261,N_5098,N_5167);
nor U5262 (N_5262,N_5021,N_5082);
or U5263 (N_5263,N_5141,N_5142);
and U5264 (N_5264,N_5056,N_5106);
and U5265 (N_5265,N_5012,N_5088);
nand U5266 (N_5266,N_5199,N_5093);
nand U5267 (N_5267,N_5089,N_5164);
and U5268 (N_5268,N_5019,N_5111);
nand U5269 (N_5269,N_5071,N_5103);
nand U5270 (N_5270,N_5113,N_5085);
nor U5271 (N_5271,N_5114,N_5072);
and U5272 (N_5272,N_5187,N_5160);
and U5273 (N_5273,N_5186,N_5011);
or U5274 (N_5274,N_5065,N_5020);
nor U5275 (N_5275,N_5177,N_5175);
nor U5276 (N_5276,N_5168,N_5004);
and U5277 (N_5277,N_5053,N_5123);
nor U5278 (N_5278,N_5112,N_5132);
nand U5279 (N_5279,N_5143,N_5035);
nand U5280 (N_5280,N_5077,N_5059);
or U5281 (N_5281,N_5144,N_5104);
nand U5282 (N_5282,N_5050,N_5153);
nand U5283 (N_5283,N_5083,N_5080);
and U5284 (N_5284,N_5090,N_5042);
or U5285 (N_5285,N_5149,N_5116);
or U5286 (N_5286,N_5137,N_5155);
and U5287 (N_5287,N_5033,N_5074);
nand U5288 (N_5288,N_5127,N_5179);
nand U5289 (N_5289,N_5046,N_5154);
nor U5290 (N_5290,N_5091,N_5169);
and U5291 (N_5291,N_5092,N_5052);
nor U5292 (N_5292,N_5118,N_5146);
and U5293 (N_5293,N_5014,N_5128);
nor U5294 (N_5294,N_5173,N_5038);
and U5295 (N_5295,N_5147,N_5172);
nor U5296 (N_5296,N_5066,N_5135);
nor U5297 (N_5297,N_5027,N_5102);
nor U5298 (N_5298,N_5062,N_5031);
or U5299 (N_5299,N_5055,N_5041);
nand U5300 (N_5300,N_5030,N_5133);
or U5301 (N_5301,N_5111,N_5195);
or U5302 (N_5302,N_5007,N_5041);
and U5303 (N_5303,N_5077,N_5199);
nor U5304 (N_5304,N_5026,N_5179);
nor U5305 (N_5305,N_5123,N_5023);
nand U5306 (N_5306,N_5161,N_5051);
or U5307 (N_5307,N_5178,N_5175);
or U5308 (N_5308,N_5088,N_5124);
or U5309 (N_5309,N_5192,N_5087);
and U5310 (N_5310,N_5112,N_5158);
or U5311 (N_5311,N_5065,N_5119);
nor U5312 (N_5312,N_5195,N_5005);
and U5313 (N_5313,N_5190,N_5059);
nor U5314 (N_5314,N_5162,N_5111);
or U5315 (N_5315,N_5185,N_5070);
and U5316 (N_5316,N_5171,N_5176);
or U5317 (N_5317,N_5114,N_5053);
or U5318 (N_5318,N_5025,N_5096);
and U5319 (N_5319,N_5196,N_5066);
or U5320 (N_5320,N_5076,N_5018);
nand U5321 (N_5321,N_5117,N_5187);
and U5322 (N_5322,N_5078,N_5121);
and U5323 (N_5323,N_5144,N_5138);
or U5324 (N_5324,N_5040,N_5156);
nand U5325 (N_5325,N_5098,N_5162);
nand U5326 (N_5326,N_5129,N_5161);
nor U5327 (N_5327,N_5078,N_5120);
and U5328 (N_5328,N_5141,N_5069);
and U5329 (N_5329,N_5048,N_5031);
nand U5330 (N_5330,N_5115,N_5040);
nor U5331 (N_5331,N_5121,N_5116);
and U5332 (N_5332,N_5154,N_5016);
and U5333 (N_5333,N_5164,N_5188);
nor U5334 (N_5334,N_5150,N_5160);
or U5335 (N_5335,N_5082,N_5126);
nor U5336 (N_5336,N_5184,N_5107);
and U5337 (N_5337,N_5130,N_5165);
nor U5338 (N_5338,N_5121,N_5074);
nand U5339 (N_5339,N_5153,N_5136);
nor U5340 (N_5340,N_5021,N_5089);
nor U5341 (N_5341,N_5013,N_5023);
nor U5342 (N_5342,N_5089,N_5017);
or U5343 (N_5343,N_5129,N_5018);
nor U5344 (N_5344,N_5109,N_5161);
and U5345 (N_5345,N_5081,N_5177);
nor U5346 (N_5346,N_5057,N_5059);
or U5347 (N_5347,N_5092,N_5112);
xor U5348 (N_5348,N_5156,N_5011);
and U5349 (N_5349,N_5005,N_5049);
nand U5350 (N_5350,N_5116,N_5158);
nor U5351 (N_5351,N_5148,N_5145);
and U5352 (N_5352,N_5096,N_5176);
nor U5353 (N_5353,N_5056,N_5085);
or U5354 (N_5354,N_5149,N_5166);
and U5355 (N_5355,N_5093,N_5115);
or U5356 (N_5356,N_5003,N_5133);
nor U5357 (N_5357,N_5160,N_5121);
or U5358 (N_5358,N_5020,N_5088);
nand U5359 (N_5359,N_5091,N_5071);
and U5360 (N_5360,N_5159,N_5048);
nand U5361 (N_5361,N_5030,N_5014);
nand U5362 (N_5362,N_5115,N_5196);
nand U5363 (N_5363,N_5001,N_5153);
or U5364 (N_5364,N_5084,N_5093);
nor U5365 (N_5365,N_5088,N_5118);
nand U5366 (N_5366,N_5025,N_5193);
nor U5367 (N_5367,N_5156,N_5187);
nor U5368 (N_5368,N_5143,N_5105);
nand U5369 (N_5369,N_5128,N_5069);
and U5370 (N_5370,N_5128,N_5198);
nand U5371 (N_5371,N_5162,N_5107);
nand U5372 (N_5372,N_5199,N_5149);
nor U5373 (N_5373,N_5108,N_5073);
xor U5374 (N_5374,N_5197,N_5060);
nand U5375 (N_5375,N_5153,N_5060);
and U5376 (N_5376,N_5170,N_5046);
or U5377 (N_5377,N_5065,N_5199);
nor U5378 (N_5378,N_5006,N_5020);
or U5379 (N_5379,N_5028,N_5071);
nand U5380 (N_5380,N_5192,N_5151);
and U5381 (N_5381,N_5070,N_5193);
and U5382 (N_5382,N_5156,N_5167);
and U5383 (N_5383,N_5174,N_5126);
and U5384 (N_5384,N_5083,N_5152);
nor U5385 (N_5385,N_5116,N_5181);
nor U5386 (N_5386,N_5154,N_5128);
nand U5387 (N_5387,N_5144,N_5080);
nand U5388 (N_5388,N_5190,N_5141);
or U5389 (N_5389,N_5061,N_5006);
nor U5390 (N_5390,N_5086,N_5166);
nand U5391 (N_5391,N_5096,N_5006);
nor U5392 (N_5392,N_5140,N_5191);
or U5393 (N_5393,N_5073,N_5088);
and U5394 (N_5394,N_5067,N_5065);
nor U5395 (N_5395,N_5097,N_5058);
and U5396 (N_5396,N_5065,N_5191);
and U5397 (N_5397,N_5154,N_5061);
nand U5398 (N_5398,N_5112,N_5126);
or U5399 (N_5399,N_5063,N_5000);
nor U5400 (N_5400,N_5382,N_5239);
xnor U5401 (N_5401,N_5214,N_5346);
and U5402 (N_5402,N_5282,N_5389);
or U5403 (N_5403,N_5221,N_5390);
nor U5404 (N_5404,N_5355,N_5253);
or U5405 (N_5405,N_5391,N_5333);
nor U5406 (N_5406,N_5216,N_5260);
or U5407 (N_5407,N_5331,N_5236);
nor U5408 (N_5408,N_5302,N_5265);
or U5409 (N_5409,N_5245,N_5339);
nor U5410 (N_5410,N_5304,N_5257);
nor U5411 (N_5411,N_5227,N_5250);
nand U5412 (N_5412,N_5363,N_5262);
nand U5413 (N_5413,N_5207,N_5228);
and U5414 (N_5414,N_5213,N_5200);
nand U5415 (N_5415,N_5308,N_5283);
nand U5416 (N_5416,N_5392,N_5217);
nand U5417 (N_5417,N_5277,N_5337);
or U5418 (N_5418,N_5268,N_5290);
nand U5419 (N_5419,N_5320,N_5233);
or U5420 (N_5420,N_5319,N_5259);
nor U5421 (N_5421,N_5297,N_5323);
or U5422 (N_5422,N_5359,N_5209);
or U5423 (N_5423,N_5338,N_5352);
and U5424 (N_5424,N_5347,N_5332);
and U5425 (N_5425,N_5276,N_5223);
or U5426 (N_5426,N_5350,N_5327);
and U5427 (N_5427,N_5241,N_5356);
or U5428 (N_5428,N_5295,N_5314);
and U5429 (N_5429,N_5203,N_5396);
or U5430 (N_5430,N_5201,N_5397);
xor U5431 (N_5431,N_5254,N_5362);
nor U5432 (N_5432,N_5249,N_5376);
nand U5433 (N_5433,N_5393,N_5287);
nor U5434 (N_5434,N_5235,N_5354);
or U5435 (N_5435,N_5374,N_5267);
and U5436 (N_5436,N_5368,N_5274);
or U5437 (N_5437,N_5315,N_5357);
or U5438 (N_5438,N_5312,N_5300);
or U5439 (N_5439,N_5344,N_5351);
nor U5440 (N_5440,N_5345,N_5293);
or U5441 (N_5441,N_5336,N_5311);
or U5442 (N_5442,N_5296,N_5263);
or U5443 (N_5443,N_5303,N_5219);
nand U5444 (N_5444,N_5335,N_5322);
nor U5445 (N_5445,N_5281,N_5328);
nand U5446 (N_5446,N_5211,N_5298);
nor U5447 (N_5447,N_5324,N_5398);
nand U5448 (N_5448,N_5224,N_5394);
or U5449 (N_5449,N_5310,N_5387);
nand U5450 (N_5450,N_5210,N_5273);
nand U5451 (N_5451,N_5342,N_5204);
nor U5452 (N_5452,N_5215,N_5399);
nor U5453 (N_5453,N_5229,N_5206);
or U5454 (N_5454,N_5232,N_5301);
or U5455 (N_5455,N_5358,N_5309);
or U5456 (N_5456,N_5349,N_5266);
nor U5457 (N_5457,N_5377,N_5271);
nor U5458 (N_5458,N_5348,N_5225);
nand U5459 (N_5459,N_5258,N_5329);
and U5460 (N_5460,N_5388,N_5321);
and U5461 (N_5461,N_5378,N_5270);
nand U5462 (N_5462,N_5294,N_5325);
nor U5463 (N_5463,N_5386,N_5222);
and U5464 (N_5464,N_5366,N_5318);
nand U5465 (N_5465,N_5292,N_5384);
nor U5466 (N_5466,N_5237,N_5316);
nor U5467 (N_5467,N_5286,N_5272);
or U5468 (N_5468,N_5251,N_5341);
or U5469 (N_5469,N_5305,N_5252);
nor U5470 (N_5470,N_5383,N_5380);
nor U5471 (N_5471,N_5231,N_5289);
nor U5472 (N_5472,N_5220,N_5285);
nand U5473 (N_5473,N_5306,N_5242);
nand U5474 (N_5474,N_5261,N_5269);
nor U5475 (N_5475,N_5218,N_5234);
nand U5476 (N_5476,N_5202,N_5255);
nand U5477 (N_5477,N_5330,N_5361);
nand U5478 (N_5478,N_5371,N_5334);
nand U5479 (N_5479,N_5243,N_5326);
nor U5480 (N_5480,N_5244,N_5279);
nor U5481 (N_5481,N_5353,N_5369);
nor U5482 (N_5482,N_5291,N_5248);
and U5483 (N_5483,N_5256,N_5278);
nand U5484 (N_5484,N_5343,N_5372);
and U5485 (N_5485,N_5284,N_5364);
nor U5486 (N_5486,N_5230,N_5307);
or U5487 (N_5487,N_5238,N_5275);
or U5488 (N_5488,N_5395,N_5288);
xnor U5489 (N_5489,N_5365,N_5280);
nor U5490 (N_5490,N_5381,N_5360);
nand U5491 (N_5491,N_5379,N_5317);
xor U5492 (N_5492,N_5246,N_5385);
or U5493 (N_5493,N_5313,N_5299);
nand U5494 (N_5494,N_5247,N_5205);
nand U5495 (N_5495,N_5367,N_5212);
nand U5496 (N_5496,N_5340,N_5240);
and U5497 (N_5497,N_5264,N_5375);
or U5498 (N_5498,N_5373,N_5226);
nand U5499 (N_5499,N_5370,N_5208);
or U5500 (N_5500,N_5358,N_5301);
or U5501 (N_5501,N_5276,N_5216);
or U5502 (N_5502,N_5394,N_5277);
nor U5503 (N_5503,N_5386,N_5218);
nand U5504 (N_5504,N_5246,N_5201);
and U5505 (N_5505,N_5387,N_5284);
or U5506 (N_5506,N_5345,N_5251);
and U5507 (N_5507,N_5231,N_5353);
and U5508 (N_5508,N_5362,N_5358);
nor U5509 (N_5509,N_5340,N_5351);
and U5510 (N_5510,N_5279,N_5202);
or U5511 (N_5511,N_5284,N_5257);
and U5512 (N_5512,N_5353,N_5271);
nand U5513 (N_5513,N_5285,N_5226);
or U5514 (N_5514,N_5316,N_5333);
or U5515 (N_5515,N_5388,N_5214);
nand U5516 (N_5516,N_5390,N_5318);
and U5517 (N_5517,N_5362,N_5342);
nand U5518 (N_5518,N_5348,N_5399);
and U5519 (N_5519,N_5277,N_5393);
or U5520 (N_5520,N_5305,N_5303);
and U5521 (N_5521,N_5258,N_5266);
nand U5522 (N_5522,N_5224,N_5310);
nor U5523 (N_5523,N_5278,N_5282);
nor U5524 (N_5524,N_5324,N_5200);
nor U5525 (N_5525,N_5372,N_5392);
nor U5526 (N_5526,N_5202,N_5247);
and U5527 (N_5527,N_5262,N_5335);
or U5528 (N_5528,N_5288,N_5209);
nand U5529 (N_5529,N_5378,N_5393);
and U5530 (N_5530,N_5291,N_5399);
and U5531 (N_5531,N_5392,N_5382);
nand U5532 (N_5532,N_5331,N_5394);
and U5533 (N_5533,N_5389,N_5243);
nand U5534 (N_5534,N_5234,N_5388);
and U5535 (N_5535,N_5236,N_5298);
and U5536 (N_5536,N_5240,N_5382);
and U5537 (N_5537,N_5213,N_5284);
and U5538 (N_5538,N_5322,N_5217);
and U5539 (N_5539,N_5218,N_5284);
and U5540 (N_5540,N_5264,N_5263);
nand U5541 (N_5541,N_5358,N_5256);
xor U5542 (N_5542,N_5283,N_5349);
and U5543 (N_5543,N_5302,N_5318);
nand U5544 (N_5544,N_5324,N_5338);
and U5545 (N_5545,N_5239,N_5353);
nor U5546 (N_5546,N_5320,N_5375);
nand U5547 (N_5547,N_5220,N_5398);
nand U5548 (N_5548,N_5281,N_5371);
nor U5549 (N_5549,N_5356,N_5222);
nand U5550 (N_5550,N_5364,N_5303);
or U5551 (N_5551,N_5388,N_5210);
and U5552 (N_5552,N_5352,N_5390);
nor U5553 (N_5553,N_5378,N_5210);
nor U5554 (N_5554,N_5268,N_5372);
nor U5555 (N_5555,N_5368,N_5304);
or U5556 (N_5556,N_5255,N_5347);
nand U5557 (N_5557,N_5298,N_5321);
and U5558 (N_5558,N_5249,N_5309);
nor U5559 (N_5559,N_5345,N_5214);
nand U5560 (N_5560,N_5362,N_5348);
or U5561 (N_5561,N_5219,N_5224);
nand U5562 (N_5562,N_5393,N_5334);
and U5563 (N_5563,N_5247,N_5309);
nand U5564 (N_5564,N_5286,N_5202);
nand U5565 (N_5565,N_5293,N_5342);
nand U5566 (N_5566,N_5366,N_5246);
and U5567 (N_5567,N_5214,N_5269);
and U5568 (N_5568,N_5354,N_5347);
or U5569 (N_5569,N_5364,N_5216);
and U5570 (N_5570,N_5323,N_5370);
and U5571 (N_5571,N_5344,N_5318);
and U5572 (N_5572,N_5387,N_5239);
and U5573 (N_5573,N_5227,N_5319);
and U5574 (N_5574,N_5396,N_5336);
or U5575 (N_5575,N_5268,N_5208);
or U5576 (N_5576,N_5267,N_5289);
and U5577 (N_5577,N_5289,N_5247);
nand U5578 (N_5578,N_5381,N_5263);
nor U5579 (N_5579,N_5285,N_5274);
nor U5580 (N_5580,N_5298,N_5326);
or U5581 (N_5581,N_5332,N_5320);
nand U5582 (N_5582,N_5283,N_5248);
and U5583 (N_5583,N_5228,N_5237);
nand U5584 (N_5584,N_5205,N_5344);
and U5585 (N_5585,N_5289,N_5208);
nand U5586 (N_5586,N_5394,N_5309);
nand U5587 (N_5587,N_5220,N_5318);
and U5588 (N_5588,N_5383,N_5374);
xor U5589 (N_5589,N_5294,N_5236);
nor U5590 (N_5590,N_5204,N_5390);
nand U5591 (N_5591,N_5229,N_5378);
or U5592 (N_5592,N_5278,N_5391);
nand U5593 (N_5593,N_5363,N_5333);
nor U5594 (N_5594,N_5396,N_5208);
nor U5595 (N_5595,N_5242,N_5367);
nand U5596 (N_5596,N_5240,N_5357);
or U5597 (N_5597,N_5271,N_5368);
nand U5598 (N_5598,N_5216,N_5373);
and U5599 (N_5599,N_5353,N_5363);
nor U5600 (N_5600,N_5488,N_5519);
nor U5601 (N_5601,N_5523,N_5400);
nor U5602 (N_5602,N_5484,N_5422);
nand U5603 (N_5603,N_5430,N_5502);
or U5604 (N_5604,N_5421,N_5461);
or U5605 (N_5605,N_5577,N_5442);
nor U5606 (N_5606,N_5532,N_5414);
or U5607 (N_5607,N_5591,N_5474);
and U5608 (N_5608,N_5477,N_5471);
or U5609 (N_5609,N_5452,N_5548);
or U5610 (N_5610,N_5424,N_5436);
nand U5611 (N_5611,N_5538,N_5459);
nand U5612 (N_5612,N_5581,N_5566);
nand U5613 (N_5613,N_5563,N_5470);
and U5614 (N_5614,N_5570,N_5554);
and U5615 (N_5615,N_5508,N_5499);
nor U5616 (N_5616,N_5520,N_5453);
nor U5617 (N_5617,N_5460,N_5439);
or U5618 (N_5618,N_5450,N_5464);
nor U5619 (N_5619,N_5446,N_5504);
or U5620 (N_5620,N_5483,N_5408);
and U5621 (N_5621,N_5463,N_5443);
or U5622 (N_5622,N_5413,N_5480);
nand U5623 (N_5623,N_5475,N_5423);
nor U5624 (N_5624,N_5431,N_5564);
nor U5625 (N_5625,N_5466,N_5547);
and U5626 (N_5626,N_5597,N_5418);
nand U5627 (N_5627,N_5507,N_5485);
and U5628 (N_5628,N_5575,N_5513);
xnor U5629 (N_5629,N_5494,N_5425);
and U5630 (N_5630,N_5593,N_5486);
nand U5631 (N_5631,N_5412,N_5448);
nand U5632 (N_5632,N_5540,N_5567);
nor U5633 (N_5633,N_5451,N_5449);
nand U5634 (N_5634,N_5496,N_5556);
or U5635 (N_5635,N_5403,N_5510);
nand U5636 (N_5636,N_5506,N_5557);
nor U5637 (N_5637,N_5522,N_5517);
or U5638 (N_5638,N_5509,N_5573);
xnor U5639 (N_5639,N_5565,N_5571);
nand U5640 (N_5640,N_5497,N_5440);
nand U5641 (N_5641,N_5530,N_5427);
and U5642 (N_5642,N_5415,N_5587);
or U5643 (N_5643,N_5489,N_5582);
nand U5644 (N_5644,N_5405,N_5589);
or U5645 (N_5645,N_5598,N_5516);
and U5646 (N_5646,N_5553,N_5526);
nand U5647 (N_5647,N_5447,N_5482);
nand U5648 (N_5648,N_5562,N_5503);
xor U5649 (N_5649,N_5455,N_5535);
nand U5650 (N_5650,N_5402,N_5576);
or U5651 (N_5651,N_5435,N_5527);
xnor U5652 (N_5652,N_5479,N_5596);
nor U5653 (N_5653,N_5595,N_5539);
nor U5654 (N_5654,N_5438,N_5478);
nand U5655 (N_5655,N_5457,N_5492);
and U5656 (N_5656,N_5417,N_5501);
nand U5657 (N_5657,N_5444,N_5584);
nor U5658 (N_5658,N_5546,N_5433);
nor U5659 (N_5659,N_5420,N_5580);
nand U5660 (N_5660,N_5524,N_5594);
nor U5661 (N_5661,N_5531,N_5560);
or U5662 (N_5662,N_5572,N_5528);
nand U5663 (N_5663,N_5586,N_5536);
and U5664 (N_5664,N_5541,N_5518);
nand U5665 (N_5665,N_5409,N_5544);
nor U5666 (N_5666,N_5491,N_5545);
nand U5667 (N_5667,N_5411,N_5500);
nand U5668 (N_5668,N_5543,N_5515);
nand U5669 (N_5669,N_5551,N_5406);
and U5670 (N_5670,N_5579,N_5592);
nand U5671 (N_5671,N_5454,N_5549);
nand U5672 (N_5672,N_5590,N_5529);
or U5673 (N_5673,N_5469,N_5521);
nor U5674 (N_5674,N_5490,N_5583);
or U5675 (N_5675,N_5476,N_5410);
nand U5676 (N_5676,N_5441,N_5487);
nand U5677 (N_5677,N_5437,N_5585);
nor U5678 (N_5678,N_5445,N_5552);
and U5679 (N_5679,N_5419,N_5542);
nand U5680 (N_5680,N_5558,N_5473);
nand U5681 (N_5681,N_5429,N_5434);
nor U5682 (N_5682,N_5537,N_5514);
and U5683 (N_5683,N_5495,N_5505);
or U5684 (N_5684,N_5533,N_5561);
nor U5685 (N_5685,N_5512,N_5555);
or U5686 (N_5686,N_5525,N_5550);
nor U5687 (N_5687,N_5428,N_5493);
nand U5688 (N_5688,N_5481,N_5511);
or U5689 (N_5689,N_5578,N_5599);
nand U5690 (N_5690,N_5498,N_5432);
nor U5691 (N_5691,N_5456,N_5401);
or U5692 (N_5692,N_5574,N_5462);
and U5693 (N_5693,N_5426,N_5534);
and U5694 (N_5694,N_5407,N_5568);
or U5695 (N_5695,N_5468,N_5467);
or U5696 (N_5696,N_5588,N_5472);
nor U5697 (N_5697,N_5416,N_5404);
or U5698 (N_5698,N_5458,N_5559);
and U5699 (N_5699,N_5569,N_5465);
and U5700 (N_5700,N_5511,N_5462);
or U5701 (N_5701,N_5478,N_5427);
or U5702 (N_5702,N_5560,N_5436);
nand U5703 (N_5703,N_5491,N_5553);
nand U5704 (N_5704,N_5487,N_5489);
nor U5705 (N_5705,N_5572,N_5578);
nor U5706 (N_5706,N_5582,N_5530);
nand U5707 (N_5707,N_5484,N_5576);
nor U5708 (N_5708,N_5536,N_5502);
or U5709 (N_5709,N_5428,N_5491);
nor U5710 (N_5710,N_5537,N_5460);
nor U5711 (N_5711,N_5438,N_5456);
nor U5712 (N_5712,N_5595,N_5516);
or U5713 (N_5713,N_5468,N_5522);
nor U5714 (N_5714,N_5481,N_5512);
nand U5715 (N_5715,N_5446,N_5553);
nand U5716 (N_5716,N_5469,N_5460);
nor U5717 (N_5717,N_5440,N_5417);
nand U5718 (N_5718,N_5566,N_5587);
nand U5719 (N_5719,N_5529,N_5514);
and U5720 (N_5720,N_5542,N_5449);
or U5721 (N_5721,N_5523,N_5504);
nor U5722 (N_5722,N_5588,N_5581);
nand U5723 (N_5723,N_5557,N_5526);
xnor U5724 (N_5724,N_5514,N_5549);
and U5725 (N_5725,N_5482,N_5589);
nor U5726 (N_5726,N_5467,N_5440);
nand U5727 (N_5727,N_5541,N_5569);
nand U5728 (N_5728,N_5596,N_5560);
nand U5729 (N_5729,N_5469,N_5439);
or U5730 (N_5730,N_5420,N_5524);
and U5731 (N_5731,N_5570,N_5448);
nand U5732 (N_5732,N_5531,N_5528);
and U5733 (N_5733,N_5544,N_5421);
and U5734 (N_5734,N_5507,N_5474);
or U5735 (N_5735,N_5511,N_5497);
or U5736 (N_5736,N_5464,N_5529);
nor U5737 (N_5737,N_5480,N_5574);
or U5738 (N_5738,N_5455,N_5538);
nand U5739 (N_5739,N_5529,N_5500);
nand U5740 (N_5740,N_5500,N_5463);
nor U5741 (N_5741,N_5401,N_5493);
nand U5742 (N_5742,N_5571,N_5462);
or U5743 (N_5743,N_5427,N_5484);
nand U5744 (N_5744,N_5585,N_5413);
nor U5745 (N_5745,N_5400,N_5550);
and U5746 (N_5746,N_5589,N_5491);
nor U5747 (N_5747,N_5500,N_5475);
or U5748 (N_5748,N_5503,N_5435);
or U5749 (N_5749,N_5574,N_5437);
or U5750 (N_5750,N_5592,N_5491);
nor U5751 (N_5751,N_5427,N_5578);
nand U5752 (N_5752,N_5407,N_5524);
nand U5753 (N_5753,N_5490,N_5516);
nor U5754 (N_5754,N_5511,N_5504);
and U5755 (N_5755,N_5456,N_5449);
and U5756 (N_5756,N_5463,N_5423);
nand U5757 (N_5757,N_5475,N_5402);
nor U5758 (N_5758,N_5456,N_5484);
nand U5759 (N_5759,N_5476,N_5444);
or U5760 (N_5760,N_5447,N_5409);
nand U5761 (N_5761,N_5450,N_5467);
nor U5762 (N_5762,N_5450,N_5503);
nor U5763 (N_5763,N_5461,N_5418);
and U5764 (N_5764,N_5460,N_5588);
xnor U5765 (N_5765,N_5553,N_5547);
nor U5766 (N_5766,N_5549,N_5565);
nand U5767 (N_5767,N_5406,N_5412);
nor U5768 (N_5768,N_5509,N_5425);
or U5769 (N_5769,N_5475,N_5447);
or U5770 (N_5770,N_5526,N_5534);
nor U5771 (N_5771,N_5582,N_5596);
nand U5772 (N_5772,N_5455,N_5434);
nor U5773 (N_5773,N_5492,N_5518);
or U5774 (N_5774,N_5439,N_5506);
and U5775 (N_5775,N_5547,N_5530);
nor U5776 (N_5776,N_5533,N_5574);
or U5777 (N_5777,N_5535,N_5465);
or U5778 (N_5778,N_5410,N_5488);
and U5779 (N_5779,N_5497,N_5577);
nand U5780 (N_5780,N_5548,N_5536);
or U5781 (N_5781,N_5565,N_5473);
nor U5782 (N_5782,N_5537,N_5517);
nand U5783 (N_5783,N_5505,N_5400);
or U5784 (N_5784,N_5550,N_5460);
and U5785 (N_5785,N_5466,N_5582);
or U5786 (N_5786,N_5421,N_5438);
or U5787 (N_5787,N_5423,N_5435);
and U5788 (N_5788,N_5525,N_5496);
nand U5789 (N_5789,N_5483,N_5537);
nor U5790 (N_5790,N_5578,N_5555);
nor U5791 (N_5791,N_5520,N_5581);
nand U5792 (N_5792,N_5472,N_5585);
or U5793 (N_5793,N_5502,N_5443);
and U5794 (N_5794,N_5500,N_5575);
and U5795 (N_5795,N_5404,N_5422);
nor U5796 (N_5796,N_5444,N_5517);
and U5797 (N_5797,N_5597,N_5524);
nand U5798 (N_5798,N_5425,N_5505);
nor U5799 (N_5799,N_5566,N_5482);
nor U5800 (N_5800,N_5622,N_5723);
nand U5801 (N_5801,N_5717,N_5633);
nand U5802 (N_5802,N_5677,N_5678);
nor U5803 (N_5803,N_5642,N_5604);
nand U5804 (N_5804,N_5740,N_5755);
nand U5805 (N_5805,N_5735,N_5745);
nor U5806 (N_5806,N_5738,N_5646);
or U5807 (N_5807,N_5650,N_5751);
nor U5808 (N_5808,N_5785,N_5744);
and U5809 (N_5809,N_5787,N_5728);
or U5810 (N_5810,N_5747,N_5765);
or U5811 (N_5811,N_5724,N_5776);
and U5812 (N_5812,N_5764,N_5772);
and U5813 (N_5813,N_5661,N_5699);
nand U5814 (N_5814,N_5795,N_5784);
nand U5815 (N_5815,N_5609,N_5621);
or U5816 (N_5816,N_5758,N_5788);
and U5817 (N_5817,N_5783,N_5750);
or U5818 (N_5818,N_5671,N_5647);
nor U5819 (N_5819,N_5620,N_5682);
nor U5820 (N_5820,N_5666,N_5779);
nand U5821 (N_5821,N_5654,N_5658);
nand U5822 (N_5822,N_5760,N_5739);
or U5823 (N_5823,N_5681,N_5617);
nand U5824 (N_5824,N_5675,N_5632);
xor U5825 (N_5825,N_5610,N_5670);
or U5826 (N_5826,N_5746,N_5732);
and U5827 (N_5827,N_5719,N_5612);
or U5828 (N_5828,N_5718,N_5660);
and U5829 (N_5829,N_5704,N_5680);
xor U5830 (N_5830,N_5606,N_5625);
and U5831 (N_5831,N_5623,N_5708);
and U5832 (N_5832,N_5792,N_5796);
or U5833 (N_5833,N_5727,N_5641);
and U5834 (N_5834,N_5791,N_5626);
and U5835 (N_5835,N_5611,N_5798);
or U5836 (N_5836,N_5715,N_5692);
nor U5837 (N_5837,N_5733,N_5731);
and U5838 (N_5838,N_5656,N_5702);
nor U5839 (N_5839,N_5768,N_5673);
and U5840 (N_5840,N_5770,N_5655);
nor U5841 (N_5841,N_5707,N_5616);
nor U5842 (N_5842,N_5635,N_5657);
nor U5843 (N_5843,N_5722,N_5684);
or U5844 (N_5844,N_5631,N_5749);
nor U5845 (N_5845,N_5651,N_5607);
and U5846 (N_5846,N_5759,N_5696);
and U5847 (N_5847,N_5780,N_5775);
or U5848 (N_5848,N_5629,N_5648);
and U5849 (N_5849,N_5627,N_5762);
nor U5850 (N_5850,N_5608,N_5662);
nand U5851 (N_5851,N_5679,N_5725);
or U5852 (N_5852,N_5705,N_5726);
nor U5853 (N_5853,N_5634,N_5676);
or U5854 (N_5854,N_5721,N_5672);
nand U5855 (N_5855,N_5709,N_5789);
nor U5856 (N_5856,N_5754,N_5771);
or U5857 (N_5857,N_5685,N_5663);
and U5858 (N_5858,N_5630,N_5689);
nor U5859 (N_5859,N_5761,N_5763);
nand U5860 (N_5860,N_5605,N_5624);
nor U5861 (N_5861,N_5638,N_5737);
nor U5862 (N_5862,N_5777,N_5614);
xnor U5863 (N_5863,N_5652,N_5637);
or U5864 (N_5864,N_5730,N_5690);
or U5865 (N_5865,N_5734,N_5669);
or U5866 (N_5866,N_5720,N_5667);
nand U5867 (N_5867,N_5644,N_5619);
or U5868 (N_5868,N_5782,N_5603);
and U5869 (N_5869,N_5643,N_5645);
or U5870 (N_5870,N_5711,N_5649);
nand U5871 (N_5871,N_5665,N_5712);
nand U5872 (N_5872,N_5601,N_5602);
nor U5873 (N_5873,N_5686,N_5748);
nand U5874 (N_5874,N_5664,N_5613);
nand U5875 (N_5875,N_5640,N_5781);
nand U5876 (N_5876,N_5713,N_5766);
nand U5877 (N_5877,N_5706,N_5683);
nor U5878 (N_5878,N_5742,N_5756);
nand U5879 (N_5879,N_5687,N_5797);
or U5880 (N_5880,N_5743,N_5653);
xnor U5881 (N_5881,N_5636,N_5668);
nand U5882 (N_5882,N_5615,N_5753);
and U5883 (N_5883,N_5698,N_5716);
and U5884 (N_5884,N_5693,N_5700);
nor U5885 (N_5885,N_5697,N_5691);
and U5886 (N_5886,N_5639,N_5793);
nand U5887 (N_5887,N_5703,N_5659);
nand U5888 (N_5888,N_5710,N_5688);
and U5889 (N_5889,N_5736,N_5618);
nand U5890 (N_5890,N_5694,N_5790);
and U5891 (N_5891,N_5778,N_5786);
nor U5892 (N_5892,N_5714,N_5729);
or U5893 (N_5893,N_5794,N_5773);
nor U5894 (N_5894,N_5701,N_5600);
or U5895 (N_5895,N_5628,N_5799);
and U5896 (N_5896,N_5752,N_5774);
or U5897 (N_5897,N_5769,N_5695);
nand U5898 (N_5898,N_5767,N_5741);
or U5899 (N_5899,N_5674,N_5757);
nand U5900 (N_5900,N_5760,N_5791);
nor U5901 (N_5901,N_5613,N_5672);
or U5902 (N_5902,N_5698,N_5694);
nor U5903 (N_5903,N_5790,N_5757);
nand U5904 (N_5904,N_5690,N_5794);
nand U5905 (N_5905,N_5799,N_5744);
or U5906 (N_5906,N_5738,N_5687);
nand U5907 (N_5907,N_5761,N_5605);
nand U5908 (N_5908,N_5614,N_5675);
and U5909 (N_5909,N_5714,N_5681);
nand U5910 (N_5910,N_5704,N_5635);
or U5911 (N_5911,N_5684,N_5687);
and U5912 (N_5912,N_5651,N_5602);
nor U5913 (N_5913,N_5619,N_5661);
nand U5914 (N_5914,N_5782,N_5711);
or U5915 (N_5915,N_5642,N_5634);
and U5916 (N_5916,N_5719,N_5611);
nor U5917 (N_5917,N_5634,N_5732);
and U5918 (N_5918,N_5629,N_5724);
nor U5919 (N_5919,N_5686,N_5622);
and U5920 (N_5920,N_5717,N_5757);
nor U5921 (N_5921,N_5673,N_5780);
and U5922 (N_5922,N_5650,N_5733);
or U5923 (N_5923,N_5617,N_5669);
nor U5924 (N_5924,N_5772,N_5778);
nor U5925 (N_5925,N_5602,N_5783);
and U5926 (N_5926,N_5647,N_5771);
or U5927 (N_5927,N_5683,N_5680);
nor U5928 (N_5928,N_5631,N_5768);
and U5929 (N_5929,N_5684,N_5752);
and U5930 (N_5930,N_5739,N_5647);
and U5931 (N_5931,N_5763,N_5738);
nand U5932 (N_5932,N_5637,N_5624);
or U5933 (N_5933,N_5753,N_5656);
nor U5934 (N_5934,N_5670,N_5764);
or U5935 (N_5935,N_5782,N_5647);
and U5936 (N_5936,N_5798,N_5708);
and U5937 (N_5937,N_5777,N_5727);
or U5938 (N_5938,N_5713,N_5698);
and U5939 (N_5939,N_5625,N_5781);
or U5940 (N_5940,N_5670,N_5713);
nand U5941 (N_5941,N_5670,N_5709);
and U5942 (N_5942,N_5651,N_5787);
or U5943 (N_5943,N_5730,N_5705);
and U5944 (N_5944,N_5697,N_5659);
or U5945 (N_5945,N_5779,N_5614);
nand U5946 (N_5946,N_5772,N_5715);
and U5947 (N_5947,N_5633,N_5791);
nor U5948 (N_5948,N_5671,N_5754);
and U5949 (N_5949,N_5655,N_5712);
or U5950 (N_5950,N_5602,N_5622);
and U5951 (N_5951,N_5643,N_5760);
and U5952 (N_5952,N_5685,N_5705);
nand U5953 (N_5953,N_5606,N_5791);
nor U5954 (N_5954,N_5662,N_5622);
and U5955 (N_5955,N_5677,N_5612);
nand U5956 (N_5956,N_5788,N_5630);
nor U5957 (N_5957,N_5713,N_5695);
and U5958 (N_5958,N_5753,N_5713);
or U5959 (N_5959,N_5750,N_5642);
nor U5960 (N_5960,N_5708,N_5747);
nor U5961 (N_5961,N_5682,N_5645);
nand U5962 (N_5962,N_5745,N_5635);
or U5963 (N_5963,N_5754,N_5693);
or U5964 (N_5964,N_5650,N_5770);
or U5965 (N_5965,N_5657,N_5660);
and U5966 (N_5966,N_5629,N_5683);
nor U5967 (N_5967,N_5666,N_5711);
or U5968 (N_5968,N_5670,N_5691);
or U5969 (N_5969,N_5613,N_5655);
nor U5970 (N_5970,N_5735,N_5790);
or U5971 (N_5971,N_5754,N_5668);
nor U5972 (N_5972,N_5664,N_5777);
nand U5973 (N_5973,N_5697,N_5794);
nor U5974 (N_5974,N_5622,N_5786);
or U5975 (N_5975,N_5720,N_5764);
nor U5976 (N_5976,N_5756,N_5709);
and U5977 (N_5977,N_5630,N_5700);
nand U5978 (N_5978,N_5784,N_5671);
and U5979 (N_5979,N_5611,N_5692);
nor U5980 (N_5980,N_5653,N_5619);
and U5981 (N_5981,N_5671,N_5720);
nand U5982 (N_5982,N_5694,N_5650);
nand U5983 (N_5983,N_5646,N_5707);
nand U5984 (N_5984,N_5626,N_5678);
nand U5985 (N_5985,N_5760,N_5792);
nor U5986 (N_5986,N_5674,N_5798);
and U5987 (N_5987,N_5619,N_5724);
or U5988 (N_5988,N_5607,N_5622);
or U5989 (N_5989,N_5605,N_5659);
or U5990 (N_5990,N_5709,N_5633);
nand U5991 (N_5991,N_5796,N_5670);
and U5992 (N_5992,N_5618,N_5614);
nor U5993 (N_5993,N_5681,N_5656);
nand U5994 (N_5994,N_5612,N_5743);
or U5995 (N_5995,N_5786,N_5679);
and U5996 (N_5996,N_5739,N_5703);
or U5997 (N_5997,N_5798,N_5745);
and U5998 (N_5998,N_5782,N_5735);
nand U5999 (N_5999,N_5773,N_5632);
and U6000 (N_6000,N_5950,N_5946);
and U6001 (N_6001,N_5831,N_5913);
nor U6002 (N_6002,N_5916,N_5817);
nor U6003 (N_6003,N_5865,N_5927);
or U6004 (N_6004,N_5844,N_5894);
nand U6005 (N_6005,N_5814,N_5827);
nand U6006 (N_6006,N_5860,N_5834);
or U6007 (N_6007,N_5887,N_5863);
or U6008 (N_6008,N_5858,N_5838);
nor U6009 (N_6009,N_5924,N_5918);
or U6010 (N_6010,N_5902,N_5847);
and U6011 (N_6011,N_5882,N_5888);
nand U6012 (N_6012,N_5837,N_5977);
and U6013 (N_6013,N_5819,N_5984);
and U6014 (N_6014,N_5998,N_5878);
or U6015 (N_6015,N_5898,N_5921);
nor U6016 (N_6016,N_5862,N_5892);
and U6017 (N_6017,N_5936,N_5803);
or U6018 (N_6018,N_5883,N_5801);
nand U6019 (N_6019,N_5973,N_5907);
nand U6020 (N_6020,N_5939,N_5929);
and U6021 (N_6021,N_5991,N_5861);
and U6022 (N_6022,N_5864,N_5992);
nor U6023 (N_6023,N_5983,N_5877);
and U6024 (N_6024,N_5979,N_5851);
nor U6025 (N_6025,N_5830,N_5900);
nor U6026 (N_6026,N_5920,N_5962);
and U6027 (N_6027,N_5982,N_5911);
nand U6028 (N_6028,N_5909,N_5871);
and U6029 (N_6029,N_5870,N_5853);
nand U6030 (N_6030,N_5969,N_5922);
and U6031 (N_6031,N_5874,N_5896);
and U6032 (N_6032,N_5816,N_5954);
nor U6033 (N_6033,N_5800,N_5895);
or U6034 (N_6034,N_5908,N_5928);
nor U6035 (N_6035,N_5949,N_5938);
or U6036 (N_6036,N_5981,N_5825);
nand U6037 (N_6037,N_5999,N_5856);
nor U6038 (N_6038,N_5875,N_5897);
or U6039 (N_6039,N_5947,N_5906);
or U6040 (N_6040,N_5993,N_5957);
nand U6041 (N_6041,N_5812,N_5964);
nand U6042 (N_6042,N_5881,N_5869);
nor U6043 (N_6043,N_5809,N_5893);
or U6044 (N_6044,N_5805,N_5944);
or U6045 (N_6045,N_5857,N_5822);
or U6046 (N_6046,N_5975,N_5940);
nor U6047 (N_6047,N_5855,N_5959);
nand U6048 (N_6048,N_5931,N_5914);
and U6049 (N_6049,N_5833,N_5919);
nor U6050 (N_6050,N_5824,N_5876);
nand U6051 (N_6051,N_5972,N_5839);
nor U6052 (N_6052,N_5997,N_5986);
and U6053 (N_6053,N_5842,N_5845);
xnor U6054 (N_6054,N_5933,N_5852);
nor U6055 (N_6055,N_5821,N_5899);
nand U6056 (N_6056,N_5846,N_5868);
nand U6057 (N_6057,N_5873,N_5820);
or U6058 (N_6058,N_5813,N_5996);
nand U6059 (N_6059,N_5912,N_5953);
nor U6060 (N_6060,N_5811,N_5917);
or U6061 (N_6061,N_5915,N_5884);
or U6062 (N_6062,N_5818,N_5889);
and U6063 (N_6063,N_5905,N_5988);
nor U6064 (N_6064,N_5815,N_5971);
and U6065 (N_6065,N_5945,N_5836);
or U6066 (N_6066,N_5823,N_5850);
nand U6067 (N_6067,N_5943,N_5848);
or U6068 (N_6068,N_5955,N_5832);
nand U6069 (N_6069,N_5808,N_5990);
or U6070 (N_6070,N_5886,N_5935);
nand U6071 (N_6071,N_5958,N_5910);
nor U6072 (N_6072,N_5951,N_5849);
nand U6073 (N_6073,N_5967,N_5942);
nor U6074 (N_6074,N_5966,N_5807);
or U6075 (N_6075,N_5867,N_5956);
nand U6076 (N_6076,N_5948,N_5976);
nor U6077 (N_6077,N_5891,N_5989);
nor U6078 (N_6078,N_5978,N_5802);
or U6079 (N_6079,N_5970,N_5804);
or U6080 (N_6080,N_5854,N_5932);
or U6081 (N_6081,N_5923,N_5987);
or U6082 (N_6082,N_5841,N_5859);
and U6083 (N_6083,N_5994,N_5985);
nor U6084 (N_6084,N_5866,N_5872);
or U6085 (N_6085,N_5843,N_5995);
nor U6086 (N_6086,N_5840,N_5925);
or U6087 (N_6087,N_5885,N_5965);
nand U6088 (N_6088,N_5904,N_5926);
nand U6089 (N_6089,N_5828,N_5930);
nand U6090 (N_6090,N_5879,N_5835);
nand U6091 (N_6091,N_5810,N_5961);
and U6092 (N_6092,N_5960,N_5974);
and U6093 (N_6093,N_5952,N_5968);
nand U6094 (N_6094,N_5901,N_5937);
or U6095 (N_6095,N_5806,N_5880);
and U6096 (N_6096,N_5980,N_5963);
nor U6097 (N_6097,N_5934,N_5826);
and U6098 (N_6098,N_5903,N_5941);
and U6099 (N_6099,N_5890,N_5829);
or U6100 (N_6100,N_5809,N_5807);
nand U6101 (N_6101,N_5905,N_5962);
and U6102 (N_6102,N_5934,N_5897);
or U6103 (N_6103,N_5908,N_5980);
nor U6104 (N_6104,N_5834,N_5875);
nand U6105 (N_6105,N_5891,N_5812);
and U6106 (N_6106,N_5939,N_5989);
or U6107 (N_6107,N_5923,N_5827);
nor U6108 (N_6108,N_5852,N_5865);
nor U6109 (N_6109,N_5859,N_5876);
and U6110 (N_6110,N_5903,N_5943);
or U6111 (N_6111,N_5913,N_5999);
and U6112 (N_6112,N_5917,N_5943);
nand U6113 (N_6113,N_5845,N_5965);
nand U6114 (N_6114,N_5915,N_5887);
nand U6115 (N_6115,N_5900,N_5896);
nand U6116 (N_6116,N_5827,N_5854);
or U6117 (N_6117,N_5973,N_5955);
and U6118 (N_6118,N_5805,N_5951);
nand U6119 (N_6119,N_5941,N_5934);
nand U6120 (N_6120,N_5999,N_5864);
nand U6121 (N_6121,N_5952,N_5838);
nand U6122 (N_6122,N_5807,N_5881);
nand U6123 (N_6123,N_5884,N_5909);
or U6124 (N_6124,N_5879,N_5836);
and U6125 (N_6125,N_5985,N_5874);
nand U6126 (N_6126,N_5881,N_5935);
and U6127 (N_6127,N_5979,N_5948);
and U6128 (N_6128,N_5926,N_5836);
nor U6129 (N_6129,N_5917,N_5962);
or U6130 (N_6130,N_5943,N_5969);
nor U6131 (N_6131,N_5841,N_5902);
or U6132 (N_6132,N_5870,N_5963);
nand U6133 (N_6133,N_5970,N_5893);
nand U6134 (N_6134,N_5921,N_5997);
nand U6135 (N_6135,N_5960,N_5950);
and U6136 (N_6136,N_5802,N_5880);
and U6137 (N_6137,N_5987,N_5887);
nor U6138 (N_6138,N_5834,N_5827);
nor U6139 (N_6139,N_5900,N_5902);
nand U6140 (N_6140,N_5814,N_5910);
nor U6141 (N_6141,N_5906,N_5983);
nand U6142 (N_6142,N_5873,N_5992);
and U6143 (N_6143,N_5851,N_5986);
and U6144 (N_6144,N_5995,N_5985);
nand U6145 (N_6145,N_5874,N_5955);
nand U6146 (N_6146,N_5980,N_5942);
nand U6147 (N_6147,N_5817,N_5997);
and U6148 (N_6148,N_5880,N_5911);
nor U6149 (N_6149,N_5956,N_5982);
nand U6150 (N_6150,N_5984,N_5941);
nor U6151 (N_6151,N_5889,N_5865);
nand U6152 (N_6152,N_5812,N_5857);
and U6153 (N_6153,N_5987,N_5943);
or U6154 (N_6154,N_5818,N_5933);
xnor U6155 (N_6155,N_5833,N_5876);
or U6156 (N_6156,N_5886,N_5848);
nand U6157 (N_6157,N_5838,N_5816);
nor U6158 (N_6158,N_5991,N_5945);
and U6159 (N_6159,N_5952,N_5993);
nand U6160 (N_6160,N_5900,N_5886);
or U6161 (N_6161,N_5928,N_5926);
nor U6162 (N_6162,N_5865,N_5807);
or U6163 (N_6163,N_5910,N_5952);
or U6164 (N_6164,N_5956,N_5879);
or U6165 (N_6165,N_5820,N_5944);
and U6166 (N_6166,N_5955,N_5851);
or U6167 (N_6167,N_5948,N_5869);
nor U6168 (N_6168,N_5983,N_5942);
nand U6169 (N_6169,N_5854,N_5831);
nand U6170 (N_6170,N_5838,N_5831);
or U6171 (N_6171,N_5810,N_5947);
nand U6172 (N_6172,N_5828,N_5890);
or U6173 (N_6173,N_5975,N_5930);
or U6174 (N_6174,N_5834,N_5894);
nor U6175 (N_6175,N_5822,N_5874);
or U6176 (N_6176,N_5833,N_5920);
nor U6177 (N_6177,N_5856,N_5975);
nor U6178 (N_6178,N_5943,N_5860);
or U6179 (N_6179,N_5834,N_5811);
nor U6180 (N_6180,N_5901,N_5875);
nand U6181 (N_6181,N_5895,N_5805);
nor U6182 (N_6182,N_5975,N_5888);
nand U6183 (N_6183,N_5808,N_5949);
nand U6184 (N_6184,N_5980,N_5801);
and U6185 (N_6185,N_5933,N_5971);
nor U6186 (N_6186,N_5905,N_5931);
nor U6187 (N_6187,N_5993,N_5981);
and U6188 (N_6188,N_5848,N_5887);
and U6189 (N_6189,N_5836,N_5859);
or U6190 (N_6190,N_5824,N_5830);
and U6191 (N_6191,N_5841,N_5901);
nand U6192 (N_6192,N_5992,N_5955);
nand U6193 (N_6193,N_5921,N_5945);
nor U6194 (N_6194,N_5808,N_5888);
nand U6195 (N_6195,N_5967,N_5888);
and U6196 (N_6196,N_5850,N_5885);
or U6197 (N_6197,N_5914,N_5918);
and U6198 (N_6198,N_5913,N_5998);
nor U6199 (N_6199,N_5858,N_5802);
and U6200 (N_6200,N_6093,N_6152);
nor U6201 (N_6201,N_6095,N_6147);
and U6202 (N_6202,N_6016,N_6170);
or U6203 (N_6203,N_6115,N_6020);
and U6204 (N_6204,N_6172,N_6063);
nand U6205 (N_6205,N_6189,N_6180);
or U6206 (N_6206,N_6001,N_6168);
and U6207 (N_6207,N_6013,N_6046);
nand U6208 (N_6208,N_6044,N_6070);
nand U6209 (N_6209,N_6065,N_6021);
or U6210 (N_6210,N_6167,N_6188);
or U6211 (N_6211,N_6109,N_6110);
nand U6212 (N_6212,N_6127,N_6086);
or U6213 (N_6213,N_6043,N_6066);
and U6214 (N_6214,N_6184,N_6199);
and U6215 (N_6215,N_6059,N_6061);
and U6216 (N_6216,N_6062,N_6106);
nand U6217 (N_6217,N_6111,N_6009);
or U6218 (N_6218,N_6069,N_6073);
or U6219 (N_6219,N_6162,N_6154);
nand U6220 (N_6220,N_6139,N_6079);
or U6221 (N_6221,N_6174,N_6104);
and U6222 (N_6222,N_6039,N_6140);
or U6223 (N_6223,N_6071,N_6151);
nor U6224 (N_6224,N_6018,N_6072);
nor U6225 (N_6225,N_6102,N_6027);
and U6226 (N_6226,N_6198,N_6087);
nor U6227 (N_6227,N_6025,N_6196);
nor U6228 (N_6228,N_6137,N_6081);
nor U6229 (N_6229,N_6074,N_6116);
or U6230 (N_6230,N_6060,N_6058);
or U6231 (N_6231,N_6000,N_6022);
nor U6232 (N_6232,N_6068,N_6089);
nand U6233 (N_6233,N_6161,N_6177);
or U6234 (N_6234,N_6083,N_6076);
or U6235 (N_6235,N_6004,N_6100);
nor U6236 (N_6236,N_6149,N_6194);
nor U6237 (N_6237,N_6015,N_6123);
or U6238 (N_6238,N_6145,N_6164);
or U6239 (N_6239,N_6033,N_6024);
or U6240 (N_6240,N_6176,N_6088);
and U6241 (N_6241,N_6130,N_6197);
nand U6242 (N_6242,N_6148,N_6135);
nor U6243 (N_6243,N_6173,N_6160);
and U6244 (N_6244,N_6006,N_6190);
or U6245 (N_6245,N_6049,N_6091);
nor U6246 (N_6246,N_6166,N_6040);
nand U6247 (N_6247,N_6056,N_6050);
or U6248 (N_6248,N_6120,N_6126);
and U6249 (N_6249,N_6031,N_6007);
and U6250 (N_6250,N_6193,N_6008);
nor U6251 (N_6251,N_6138,N_6171);
nor U6252 (N_6252,N_6128,N_6038);
nand U6253 (N_6253,N_6084,N_6085);
and U6254 (N_6254,N_6051,N_6187);
nand U6255 (N_6255,N_6098,N_6032);
or U6256 (N_6256,N_6141,N_6041);
nand U6257 (N_6257,N_6002,N_6142);
nor U6258 (N_6258,N_6067,N_6042);
nor U6259 (N_6259,N_6003,N_6054);
or U6260 (N_6260,N_6082,N_6169);
and U6261 (N_6261,N_6057,N_6129);
and U6262 (N_6262,N_6037,N_6186);
or U6263 (N_6263,N_6026,N_6153);
nand U6264 (N_6264,N_6108,N_6119);
nor U6265 (N_6265,N_6159,N_6121);
or U6266 (N_6266,N_6113,N_6010);
or U6267 (N_6267,N_6157,N_6014);
or U6268 (N_6268,N_6143,N_6175);
nor U6269 (N_6269,N_6178,N_6090);
and U6270 (N_6270,N_6101,N_6034);
and U6271 (N_6271,N_6080,N_6185);
nor U6272 (N_6272,N_6144,N_6107);
nor U6273 (N_6273,N_6045,N_6118);
and U6274 (N_6274,N_6011,N_6012);
nor U6275 (N_6275,N_6165,N_6182);
and U6276 (N_6276,N_6125,N_6158);
nor U6277 (N_6277,N_6075,N_6112);
nand U6278 (N_6278,N_6077,N_6156);
or U6279 (N_6279,N_6183,N_6124);
and U6280 (N_6280,N_6097,N_6155);
nand U6281 (N_6281,N_6099,N_6150);
nand U6282 (N_6282,N_6019,N_6117);
or U6283 (N_6283,N_6064,N_6131);
nor U6284 (N_6284,N_6053,N_6048);
or U6285 (N_6285,N_6103,N_6163);
nand U6286 (N_6286,N_6092,N_6035);
and U6287 (N_6287,N_6005,N_6078);
and U6288 (N_6288,N_6017,N_6122);
and U6289 (N_6289,N_6096,N_6146);
and U6290 (N_6290,N_6133,N_6094);
nand U6291 (N_6291,N_6114,N_6136);
nand U6292 (N_6292,N_6055,N_6023);
nand U6293 (N_6293,N_6192,N_6134);
or U6294 (N_6294,N_6179,N_6052);
and U6295 (N_6295,N_6132,N_6036);
nand U6296 (N_6296,N_6181,N_6029);
and U6297 (N_6297,N_6047,N_6030);
nor U6298 (N_6298,N_6195,N_6028);
nor U6299 (N_6299,N_6105,N_6191);
nor U6300 (N_6300,N_6047,N_6125);
nand U6301 (N_6301,N_6164,N_6027);
and U6302 (N_6302,N_6126,N_6015);
nor U6303 (N_6303,N_6014,N_6016);
and U6304 (N_6304,N_6017,N_6177);
nand U6305 (N_6305,N_6138,N_6076);
and U6306 (N_6306,N_6050,N_6055);
nor U6307 (N_6307,N_6099,N_6199);
nand U6308 (N_6308,N_6191,N_6198);
and U6309 (N_6309,N_6176,N_6049);
nand U6310 (N_6310,N_6010,N_6069);
or U6311 (N_6311,N_6080,N_6027);
nor U6312 (N_6312,N_6139,N_6165);
nor U6313 (N_6313,N_6019,N_6146);
and U6314 (N_6314,N_6171,N_6165);
nor U6315 (N_6315,N_6089,N_6146);
nand U6316 (N_6316,N_6182,N_6185);
and U6317 (N_6317,N_6148,N_6162);
nand U6318 (N_6318,N_6134,N_6110);
and U6319 (N_6319,N_6139,N_6082);
and U6320 (N_6320,N_6026,N_6004);
and U6321 (N_6321,N_6052,N_6051);
nor U6322 (N_6322,N_6196,N_6001);
or U6323 (N_6323,N_6196,N_6103);
or U6324 (N_6324,N_6177,N_6046);
or U6325 (N_6325,N_6037,N_6112);
nor U6326 (N_6326,N_6113,N_6111);
or U6327 (N_6327,N_6021,N_6013);
nor U6328 (N_6328,N_6102,N_6166);
nor U6329 (N_6329,N_6156,N_6193);
and U6330 (N_6330,N_6193,N_6053);
nor U6331 (N_6331,N_6062,N_6010);
and U6332 (N_6332,N_6079,N_6039);
nor U6333 (N_6333,N_6176,N_6128);
or U6334 (N_6334,N_6084,N_6057);
or U6335 (N_6335,N_6032,N_6066);
nand U6336 (N_6336,N_6102,N_6008);
or U6337 (N_6337,N_6196,N_6055);
and U6338 (N_6338,N_6147,N_6123);
nor U6339 (N_6339,N_6077,N_6088);
and U6340 (N_6340,N_6176,N_6052);
or U6341 (N_6341,N_6082,N_6131);
and U6342 (N_6342,N_6021,N_6082);
and U6343 (N_6343,N_6098,N_6190);
nand U6344 (N_6344,N_6058,N_6007);
nor U6345 (N_6345,N_6050,N_6173);
nand U6346 (N_6346,N_6016,N_6069);
nand U6347 (N_6347,N_6086,N_6079);
and U6348 (N_6348,N_6159,N_6087);
nand U6349 (N_6349,N_6146,N_6012);
or U6350 (N_6350,N_6056,N_6072);
nor U6351 (N_6351,N_6173,N_6139);
and U6352 (N_6352,N_6093,N_6191);
nand U6353 (N_6353,N_6023,N_6019);
xor U6354 (N_6354,N_6059,N_6151);
or U6355 (N_6355,N_6015,N_6184);
or U6356 (N_6356,N_6017,N_6173);
nand U6357 (N_6357,N_6191,N_6057);
and U6358 (N_6358,N_6163,N_6114);
nand U6359 (N_6359,N_6195,N_6116);
and U6360 (N_6360,N_6021,N_6076);
nor U6361 (N_6361,N_6110,N_6199);
nor U6362 (N_6362,N_6114,N_6143);
or U6363 (N_6363,N_6022,N_6040);
or U6364 (N_6364,N_6043,N_6060);
nor U6365 (N_6365,N_6135,N_6115);
and U6366 (N_6366,N_6124,N_6022);
nor U6367 (N_6367,N_6136,N_6089);
or U6368 (N_6368,N_6044,N_6186);
nand U6369 (N_6369,N_6062,N_6132);
and U6370 (N_6370,N_6189,N_6107);
nand U6371 (N_6371,N_6121,N_6006);
or U6372 (N_6372,N_6126,N_6095);
nand U6373 (N_6373,N_6187,N_6170);
nor U6374 (N_6374,N_6101,N_6003);
or U6375 (N_6375,N_6029,N_6017);
and U6376 (N_6376,N_6072,N_6159);
or U6377 (N_6377,N_6126,N_6190);
or U6378 (N_6378,N_6038,N_6127);
nand U6379 (N_6379,N_6091,N_6018);
nand U6380 (N_6380,N_6180,N_6120);
or U6381 (N_6381,N_6173,N_6125);
and U6382 (N_6382,N_6010,N_6101);
and U6383 (N_6383,N_6121,N_6027);
nor U6384 (N_6384,N_6048,N_6004);
and U6385 (N_6385,N_6068,N_6085);
nand U6386 (N_6386,N_6089,N_6073);
and U6387 (N_6387,N_6015,N_6176);
and U6388 (N_6388,N_6184,N_6003);
or U6389 (N_6389,N_6157,N_6118);
nor U6390 (N_6390,N_6029,N_6137);
nand U6391 (N_6391,N_6002,N_6110);
nor U6392 (N_6392,N_6097,N_6127);
or U6393 (N_6393,N_6046,N_6005);
nand U6394 (N_6394,N_6084,N_6165);
nor U6395 (N_6395,N_6139,N_6117);
nand U6396 (N_6396,N_6144,N_6194);
and U6397 (N_6397,N_6090,N_6141);
nand U6398 (N_6398,N_6068,N_6009);
and U6399 (N_6399,N_6099,N_6011);
nand U6400 (N_6400,N_6313,N_6270);
nor U6401 (N_6401,N_6233,N_6214);
xnor U6402 (N_6402,N_6310,N_6294);
nor U6403 (N_6403,N_6221,N_6322);
nand U6404 (N_6404,N_6251,N_6392);
and U6405 (N_6405,N_6338,N_6240);
and U6406 (N_6406,N_6399,N_6295);
or U6407 (N_6407,N_6222,N_6382);
and U6408 (N_6408,N_6250,N_6277);
nor U6409 (N_6409,N_6204,N_6228);
and U6410 (N_6410,N_6298,N_6390);
or U6411 (N_6411,N_6229,N_6306);
nor U6412 (N_6412,N_6236,N_6264);
nor U6413 (N_6413,N_6260,N_6325);
or U6414 (N_6414,N_6244,N_6334);
or U6415 (N_6415,N_6211,N_6346);
nor U6416 (N_6416,N_6219,N_6351);
and U6417 (N_6417,N_6371,N_6279);
or U6418 (N_6418,N_6234,N_6318);
nor U6419 (N_6419,N_6381,N_6353);
or U6420 (N_6420,N_6223,N_6373);
nand U6421 (N_6421,N_6230,N_6385);
nor U6422 (N_6422,N_6349,N_6337);
and U6423 (N_6423,N_6342,N_6245);
or U6424 (N_6424,N_6386,N_6398);
nor U6425 (N_6425,N_6207,N_6284);
and U6426 (N_6426,N_6352,N_6269);
nand U6427 (N_6427,N_6247,N_6308);
and U6428 (N_6428,N_6215,N_6232);
or U6429 (N_6429,N_6253,N_6267);
nand U6430 (N_6430,N_6286,N_6241);
or U6431 (N_6431,N_6345,N_6374);
nand U6432 (N_6432,N_6266,N_6393);
nor U6433 (N_6433,N_6285,N_6324);
and U6434 (N_6434,N_6384,N_6344);
nor U6435 (N_6435,N_6291,N_6378);
nand U6436 (N_6436,N_6274,N_6217);
nand U6437 (N_6437,N_6327,N_6312);
or U6438 (N_6438,N_6203,N_6243);
nand U6439 (N_6439,N_6300,N_6235);
nor U6440 (N_6440,N_6305,N_6206);
nand U6441 (N_6441,N_6258,N_6273);
nor U6442 (N_6442,N_6330,N_6356);
nand U6443 (N_6443,N_6380,N_6339);
and U6444 (N_6444,N_6304,N_6303);
nand U6445 (N_6445,N_6379,N_6212);
nand U6446 (N_6446,N_6278,N_6209);
nand U6447 (N_6447,N_6281,N_6301);
nand U6448 (N_6448,N_6362,N_6259);
and U6449 (N_6449,N_6383,N_6350);
and U6450 (N_6450,N_6329,N_6358);
or U6451 (N_6451,N_6375,N_6365);
nor U6452 (N_6452,N_6395,N_6391);
and U6453 (N_6453,N_6368,N_6265);
nor U6454 (N_6454,N_6361,N_6280);
nand U6455 (N_6455,N_6314,N_6237);
or U6456 (N_6456,N_6326,N_6220);
nor U6457 (N_6457,N_6372,N_6367);
nand U6458 (N_6458,N_6311,N_6213);
or U6459 (N_6459,N_6289,N_6377);
nand U6460 (N_6460,N_6262,N_6200);
or U6461 (N_6461,N_6388,N_6299);
or U6462 (N_6462,N_6328,N_6331);
or U6463 (N_6463,N_6355,N_6323);
nand U6464 (N_6464,N_6282,N_6307);
nor U6465 (N_6465,N_6275,N_6202);
nand U6466 (N_6466,N_6319,N_6397);
or U6467 (N_6467,N_6396,N_6332);
or U6468 (N_6468,N_6268,N_6225);
or U6469 (N_6469,N_6333,N_6370);
nor U6470 (N_6470,N_6394,N_6238);
and U6471 (N_6471,N_6341,N_6248);
nand U6472 (N_6472,N_6257,N_6292);
or U6473 (N_6473,N_6343,N_6316);
and U6474 (N_6474,N_6369,N_6255);
nor U6475 (N_6475,N_6263,N_6389);
and U6476 (N_6476,N_6283,N_6256);
nor U6477 (N_6477,N_6276,N_6340);
or U6478 (N_6478,N_6315,N_6231);
nand U6479 (N_6479,N_6297,N_6302);
or U6480 (N_6480,N_6287,N_6354);
nor U6481 (N_6481,N_6218,N_6347);
nor U6482 (N_6482,N_6201,N_6366);
and U6483 (N_6483,N_6210,N_6261);
or U6484 (N_6484,N_6205,N_6272);
nand U6485 (N_6485,N_6290,N_6359);
or U6486 (N_6486,N_6336,N_6363);
or U6487 (N_6487,N_6321,N_6254);
nor U6488 (N_6488,N_6320,N_6296);
nand U6489 (N_6489,N_6246,N_6208);
or U6490 (N_6490,N_6364,N_6224);
and U6491 (N_6491,N_6216,N_6309);
nand U6492 (N_6492,N_6239,N_6335);
and U6493 (N_6493,N_6387,N_6293);
and U6494 (N_6494,N_6252,N_6288);
or U6495 (N_6495,N_6226,N_6357);
nor U6496 (N_6496,N_6317,N_6360);
or U6497 (N_6497,N_6376,N_6271);
and U6498 (N_6498,N_6348,N_6242);
nand U6499 (N_6499,N_6249,N_6227);
and U6500 (N_6500,N_6291,N_6275);
nand U6501 (N_6501,N_6264,N_6382);
or U6502 (N_6502,N_6307,N_6319);
or U6503 (N_6503,N_6213,N_6348);
and U6504 (N_6504,N_6294,N_6376);
or U6505 (N_6505,N_6347,N_6388);
nor U6506 (N_6506,N_6392,N_6241);
and U6507 (N_6507,N_6313,N_6226);
or U6508 (N_6508,N_6308,N_6386);
nor U6509 (N_6509,N_6221,N_6233);
nand U6510 (N_6510,N_6271,N_6262);
nor U6511 (N_6511,N_6297,N_6301);
or U6512 (N_6512,N_6351,N_6283);
nand U6513 (N_6513,N_6358,N_6219);
or U6514 (N_6514,N_6249,N_6395);
nand U6515 (N_6515,N_6240,N_6376);
nor U6516 (N_6516,N_6327,N_6347);
and U6517 (N_6517,N_6389,N_6318);
nor U6518 (N_6518,N_6390,N_6348);
nand U6519 (N_6519,N_6384,N_6311);
nor U6520 (N_6520,N_6381,N_6352);
or U6521 (N_6521,N_6299,N_6220);
and U6522 (N_6522,N_6396,N_6277);
nor U6523 (N_6523,N_6311,N_6202);
and U6524 (N_6524,N_6351,N_6365);
and U6525 (N_6525,N_6390,N_6366);
nor U6526 (N_6526,N_6306,N_6362);
and U6527 (N_6527,N_6371,N_6394);
nor U6528 (N_6528,N_6342,N_6218);
or U6529 (N_6529,N_6328,N_6304);
nand U6530 (N_6530,N_6370,N_6346);
nor U6531 (N_6531,N_6274,N_6244);
or U6532 (N_6532,N_6262,N_6345);
and U6533 (N_6533,N_6387,N_6329);
and U6534 (N_6534,N_6204,N_6329);
and U6535 (N_6535,N_6200,N_6316);
and U6536 (N_6536,N_6270,N_6381);
nor U6537 (N_6537,N_6203,N_6329);
xnor U6538 (N_6538,N_6256,N_6237);
and U6539 (N_6539,N_6326,N_6366);
nor U6540 (N_6540,N_6221,N_6239);
nand U6541 (N_6541,N_6200,N_6364);
and U6542 (N_6542,N_6252,N_6341);
and U6543 (N_6543,N_6380,N_6256);
or U6544 (N_6544,N_6270,N_6317);
or U6545 (N_6545,N_6261,N_6272);
nor U6546 (N_6546,N_6327,N_6313);
or U6547 (N_6547,N_6367,N_6228);
nor U6548 (N_6548,N_6389,N_6345);
xor U6549 (N_6549,N_6349,N_6232);
nor U6550 (N_6550,N_6356,N_6279);
nor U6551 (N_6551,N_6328,N_6308);
or U6552 (N_6552,N_6251,N_6366);
nor U6553 (N_6553,N_6208,N_6347);
or U6554 (N_6554,N_6242,N_6298);
or U6555 (N_6555,N_6345,N_6337);
and U6556 (N_6556,N_6278,N_6309);
nor U6557 (N_6557,N_6252,N_6343);
and U6558 (N_6558,N_6215,N_6317);
and U6559 (N_6559,N_6311,N_6291);
or U6560 (N_6560,N_6308,N_6259);
and U6561 (N_6561,N_6214,N_6280);
nand U6562 (N_6562,N_6348,N_6324);
and U6563 (N_6563,N_6239,N_6301);
nand U6564 (N_6564,N_6338,N_6373);
and U6565 (N_6565,N_6265,N_6226);
nor U6566 (N_6566,N_6395,N_6232);
and U6567 (N_6567,N_6224,N_6230);
nand U6568 (N_6568,N_6365,N_6360);
or U6569 (N_6569,N_6302,N_6282);
xor U6570 (N_6570,N_6306,N_6224);
nand U6571 (N_6571,N_6331,N_6245);
and U6572 (N_6572,N_6331,N_6286);
or U6573 (N_6573,N_6206,N_6242);
nor U6574 (N_6574,N_6282,N_6325);
and U6575 (N_6575,N_6238,N_6303);
or U6576 (N_6576,N_6375,N_6362);
nand U6577 (N_6577,N_6282,N_6294);
nand U6578 (N_6578,N_6332,N_6306);
or U6579 (N_6579,N_6302,N_6344);
or U6580 (N_6580,N_6325,N_6222);
and U6581 (N_6581,N_6230,N_6234);
or U6582 (N_6582,N_6312,N_6220);
nand U6583 (N_6583,N_6336,N_6222);
nand U6584 (N_6584,N_6209,N_6205);
nand U6585 (N_6585,N_6339,N_6342);
or U6586 (N_6586,N_6304,N_6360);
nor U6587 (N_6587,N_6290,N_6248);
nand U6588 (N_6588,N_6279,N_6245);
nand U6589 (N_6589,N_6224,N_6280);
and U6590 (N_6590,N_6354,N_6263);
or U6591 (N_6591,N_6256,N_6302);
nand U6592 (N_6592,N_6240,N_6232);
or U6593 (N_6593,N_6395,N_6215);
and U6594 (N_6594,N_6233,N_6345);
nand U6595 (N_6595,N_6253,N_6329);
nand U6596 (N_6596,N_6360,N_6281);
and U6597 (N_6597,N_6232,N_6399);
nand U6598 (N_6598,N_6273,N_6283);
nor U6599 (N_6599,N_6341,N_6276);
nor U6600 (N_6600,N_6428,N_6408);
nor U6601 (N_6601,N_6562,N_6515);
nor U6602 (N_6602,N_6445,N_6591);
nand U6603 (N_6603,N_6485,N_6461);
nand U6604 (N_6604,N_6504,N_6547);
nand U6605 (N_6605,N_6464,N_6488);
nor U6606 (N_6606,N_6435,N_6442);
and U6607 (N_6607,N_6458,N_6487);
nor U6608 (N_6608,N_6500,N_6537);
or U6609 (N_6609,N_6528,N_6462);
or U6610 (N_6610,N_6587,N_6455);
and U6611 (N_6611,N_6534,N_6543);
nand U6612 (N_6612,N_6409,N_6482);
or U6613 (N_6613,N_6539,N_6422);
or U6614 (N_6614,N_6434,N_6484);
nor U6615 (N_6615,N_6437,N_6596);
or U6616 (N_6616,N_6465,N_6536);
or U6617 (N_6617,N_6470,N_6452);
and U6618 (N_6618,N_6598,N_6541);
or U6619 (N_6619,N_6498,N_6516);
or U6620 (N_6620,N_6432,N_6508);
or U6621 (N_6621,N_6593,N_6425);
nand U6622 (N_6622,N_6492,N_6599);
and U6623 (N_6623,N_6407,N_6479);
nor U6624 (N_6624,N_6557,N_6575);
or U6625 (N_6625,N_6467,N_6440);
nand U6626 (N_6626,N_6438,N_6589);
nand U6627 (N_6627,N_6491,N_6477);
nand U6628 (N_6628,N_6405,N_6544);
nand U6629 (N_6629,N_6566,N_6563);
or U6630 (N_6630,N_6489,N_6551);
or U6631 (N_6631,N_6414,N_6585);
nand U6632 (N_6632,N_6471,N_6548);
or U6633 (N_6633,N_6597,N_6588);
nor U6634 (N_6634,N_6431,N_6573);
xnor U6635 (N_6635,N_6542,N_6506);
nor U6636 (N_6636,N_6439,N_6501);
nand U6637 (N_6637,N_6503,N_6540);
nor U6638 (N_6638,N_6524,N_6572);
or U6639 (N_6639,N_6411,N_6586);
nor U6640 (N_6640,N_6570,N_6552);
nand U6641 (N_6641,N_6520,N_6571);
and U6642 (N_6642,N_6531,N_6430);
or U6643 (N_6643,N_6460,N_6521);
and U6644 (N_6644,N_6519,N_6433);
nand U6645 (N_6645,N_6502,N_6554);
or U6646 (N_6646,N_6436,N_6402);
or U6647 (N_6647,N_6403,N_6463);
nand U6648 (N_6648,N_6561,N_6568);
or U6649 (N_6649,N_6584,N_6416);
and U6650 (N_6650,N_6595,N_6410);
and U6651 (N_6651,N_6509,N_6449);
and U6652 (N_6652,N_6514,N_6530);
or U6653 (N_6653,N_6494,N_6472);
nor U6654 (N_6654,N_6427,N_6444);
and U6655 (N_6655,N_6486,N_6419);
nor U6656 (N_6656,N_6576,N_6406);
and U6657 (N_6657,N_6594,N_6592);
and U6658 (N_6658,N_6532,N_6418);
nor U6659 (N_6659,N_6522,N_6443);
and U6660 (N_6660,N_6527,N_6424);
or U6661 (N_6661,N_6569,N_6555);
and U6662 (N_6662,N_6490,N_6469);
nand U6663 (N_6663,N_6564,N_6483);
nor U6664 (N_6664,N_6518,N_6478);
or U6665 (N_6665,N_6404,N_6580);
and U6666 (N_6666,N_6493,N_6533);
nand U6667 (N_6667,N_6511,N_6578);
and U6668 (N_6668,N_6579,N_6447);
nor U6669 (N_6669,N_6441,N_6421);
or U6670 (N_6670,N_6525,N_6423);
or U6671 (N_6671,N_6401,N_6412);
nand U6672 (N_6672,N_6558,N_6400);
nand U6673 (N_6673,N_6512,N_6590);
nand U6674 (N_6674,N_6523,N_6497);
and U6675 (N_6675,N_6453,N_6560);
nor U6676 (N_6676,N_6526,N_6415);
nand U6677 (N_6677,N_6577,N_6475);
nor U6678 (N_6678,N_6420,N_6499);
nand U6679 (N_6679,N_6454,N_6535);
and U6680 (N_6680,N_6456,N_6413);
and U6681 (N_6681,N_6474,N_6507);
nor U6682 (N_6682,N_6450,N_6559);
and U6683 (N_6683,N_6549,N_6459);
and U6684 (N_6684,N_6582,N_6466);
nand U6685 (N_6685,N_6505,N_6496);
nand U6686 (N_6686,N_6426,N_6446);
and U6687 (N_6687,N_6510,N_6468);
nand U6688 (N_6688,N_6583,N_6545);
nand U6689 (N_6689,N_6480,N_6457);
nand U6690 (N_6690,N_6553,N_6565);
and U6691 (N_6691,N_6473,N_6513);
nand U6692 (N_6692,N_6451,N_6417);
nand U6693 (N_6693,N_6495,N_6538);
or U6694 (N_6694,N_6581,N_6567);
nor U6695 (N_6695,N_6448,N_6556);
nor U6696 (N_6696,N_6546,N_6550);
nor U6697 (N_6697,N_6476,N_6517);
nor U6698 (N_6698,N_6574,N_6481);
nor U6699 (N_6699,N_6429,N_6529);
nor U6700 (N_6700,N_6543,N_6488);
nand U6701 (N_6701,N_6492,N_6463);
or U6702 (N_6702,N_6510,N_6519);
nand U6703 (N_6703,N_6536,N_6409);
nand U6704 (N_6704,N_6490,N_6431);
nand U6705 (N_6705,N_6449,N_6445);
nand U6706 (N_6706,N_6442,N_6492);
or U6707 (N_6707,N_6405,N_6540);
nor U6708 (N_6708,N_6569,N_6512);
and U6709 (N_6709,N_6504,N_6572);
nand U6710 (N_6710,N_6566,N_6498);
and U6711 (N_6711,N_6570,N_6588);
and U6712 (N_6712,N_6581,N_6596);
nand U6713 (N_6713,N_6416,N_6520);
nand U6714 (N_6714,N_6458,N_6424);
nor U6715 (N_6715,N_6428,N_6403);
nand U6716 (N_6716,N_6548,N_6543);
or U6717 (N_6717,N_6473,N_6521);
and U6718 (N_6718,N_6593,N_6562);
nand U6719 (N_6719,N_6487,N_6574);
or U6720 (N_6720,N_6544,N_6440);
and U6721 (N_6721,N_6473,N_6490);
nand U6722 (N_6722,N_6421,N_6588);
or U6723 (N_6723,N_6579,N_6585);
and U6724 (N_6724,N_6474,N_6468);
nor U6725 (N_6725,N_6550,N_6503);
nor U6726 (N_6726,N_6421,N_6581);
nor U6727 (N_6727,N_6419,N_6565);
and U6728 (N_6728,N_6442,N_6456);
and U6729 (N_6729,N_6580,N_6437);
nand U6730 (N_6730,N_6400,N_6470);
or U6731 (N_6731,N_6483,N_6559);
nand U6732 (N_6732,N_6465,N_6446);
nor U6733 (N_6733,N_6514,N_6403);
or U6734 (N_6734,N_6451,N_6413);
and U6735 (N_6735,N_6415,N_6502);
and U6736 (N_6736,N_6430,N_6524);
and U6737 (N_6737,N_6500,N_6451);
or U6738 (N_6738,N_6595,N_6592);
nand U6739 (N_6739,N_6503,N_6516);
or U6740 (N_6740,N_6513,N_6504);
nor U6741 (N_6741,N_6593,N_6553);
and U6742 (N_6742,N_6533,N_6555);
or U6743 (N_6743,N_6515,N_6531);
and U6744 (N_6744,N_6506,N_6586);
or U6745 (N_6745,N_6524,N_6446);
or U6746 (N_6746,N_6553,N_6427);
nand U6747 (N_6747,N_6508,N_6490);
xnor U6748 (N_6748,N_6456,N_6440);
and U6749 (N_6749,N_6595,N_6439);
or U6750 (N_6750,N_6493,N_6525);
nand U6751 (N_6751,N_6480,N_6523);
nand U6752 (N_6752,N_6493,N_6536);
nand U6753 (N_6753,N_6487,N_6488);
nor U6754 (N_6754,N_6513,N_6584);
and U6755 (N_6755,N_6575,N_6406);
nor U6756 (N_6756,N_6551,N_6508);
nor U6757 (N_6757,N_6420,N_6545);
or U6758 (N_6758,N_6404,N_6452);
or U6759 (N_6759,N_6562,N_6577);
and U6760 (N_6760,N_6537,N_6561);
and U6761 (N_6761,N_6486,N_6472);
nand U6762 (N_6762,N_6429,N_6459);
nand U6763 (N_6763,N_6560,N_6419);
or U6764 (N_6764,N_6577,N_6512);
and U6765 (N_6765,N_6467,N_6401);
or U6766 (N_6766,N_6466,N_6426);
xnor U6767 (N_6767,N_6452,N_6479);
nor U6768 (N_6768,N_6483,N_6507);
and U6769 (N_6769,N_6547,N_6594);
or U6770 (N_6770,N_6489,N_6536);
or U6771 (N_6771,N_6498,N_6537);
and U6772 (N_6772,N_6455,N_6470);
nand U6773 (N_6773,N_6478,N_6555);
or U6774 (N_6774,N_6537,N_6471);
or U6775 (N_6775,N_6576,N_6579);
and U6776 (N_6776,N_6561,N_6583);
nand U6777 (N_6777,N_6585,N_6560);
or U6778 (N_6778,N_6593,N_6415);
and U6779 (N_6779,N_6537,N_6512);
and U6780 (N_6780,N_6462,N_6484);
nor U6781 (N_6781,N_6400,N_6423);
and U6782 (N_6782,N_6591,N_6418);
nand U6783 (N_6783,N_6580,N_6563);
or U6784 (N_6784,N_6474,N_6462);
nor U6785 (N_6785,N_6446,N_6563);
or U6786 (N_6786,N_6402,N_6420);
nand U6787 (N_6787,N_6526,N_6457);
nand U6788 (N_6788,N_6553,N_6496);
nor U6789 (N_6789,N_6577,N_6478);
and U6790 (N_6790,N_6400,N_6564);
nor U6791 (N_6791,N_6522,N_6488);
or U6792 (N_6792,N_6583,N_6438);
or U6793 (N_6793,N_6585,N_6545);
or U6794 (N_6794,N_6467,N_6415);
or U6795 (N_6795,N_6486,N_6444);
and U6796 (N_6796,N_6412,N_6433);
or U6797 (N_6797,N_6594,N_6554);
nand U6798 (N_6798,N_6422,N_6459);
nand U6799 (N_6799,N_6437,N_6459);
and U6800 (N_6800,N_6705,N_6687);
and U6801 (N_6801,N_6792,N_6730);
or U6802 (N_6802,N_6748,N_6601);
and U6803 (N_6803,N_6750,N_6723);
xor U6804 (N_6804,N_6630,N_6793);
or U6805 (N_6805,N_6778,N_6653);
nand U6806 (N_6806,N_6627,N_6620);
nand U6807 (N_6807,N_6798,N_6649);
or U6808 (N_6808,N_6711,N_6737);
or U6809 (N_6809,N_6741,N_6739);
and U6810 (N_6810,N_6673,N_6699);
and U6811 (N_6811,N_6787,N_6765);
and U6812 (N_6812,N_6661,N_6727);
nor U6813 (N_6813,N_6663,N_6755);
nand U6814 (N_6814,N_6635,N_6701);
nor U6815 (N_6815,N_6771,N_6725);
and U6816 (N_6816,N_6784,N_6761);
or U6817 (N_6817,N_6762,N_6652);
nor U6818 (N_6818,N_6703,N_6657);
nand U6819 (N_6819,N_6733,N_6734);
nor U6820 (N_6820,N_6641,N_6618);
and U6821 (N_6821,N_6639,N_6631);
nor U6822 (N_6822,N_6735,N_6607);
nand U6823 (N_6823,N_6722,N_6685);
or U6824 (N_6824,N_6717,N_6697);
nor U6825 (N_6825,N_6622,N_6719);
and U6826 (N_6826,N_6745,N_6772);
or U6827 (N_6827,N_6647,N_6724);
or U6828 (N_6828,N_6783,N_6769);
and U6829 (N_6829,N_6691,N_6744);
or U6830 (N_6830,N_6726,N_6752);
nand U6831 (N_6831,N_6671,N_6796);
and U6832 (N_6832,N_6742,N_6781);
or U6833 (N_6833,N_6682,N_6789);
nor U6834 (N_6834,N_6642,N_6731);
nor U6835 (N_6835,N_6776,N_6611);
nor U6836 (N_6836,N_6760,N_6614);
or U6837 (N_6837,N_6626,N_6638);
nand U6838 (N_6838,N_6788,N_6616);
and U6839 (N_6839,N_6628,N_6672);
nand U6840 (N_6840,N_6621,N_6624);
nand U6841 (N_6841,N_6651,N_6766);
and U6842 (N_6842,N_6600,N_6729);
nand U6843 (N_6843,N_6680,N_6637);
or U6844 (N_6844,N_6782,N_6692);
nor U6845 (N_6845,N_6683,N_6790);
nor U6846 (N_6846,N_6718,N_6797);
nand U6847 (N_6847,N_6674,N_6704);
nand U6848 (N_6848,N_6603,N_6708);
nor U6849 (N_6849,N_6646,N_6780);
or U6850 (N_6850,N_6754,N_6791);
and U6851 (N_6851,N_6665,N_6644);
or U6852 (N_6852,N_6656,N_6640);
nand U6853 (N_6853,N_6702,N_6688);
nand U6854 (N_6854,N_6746,N_6785);
and U6855 (N_6855,N_6707,N_6655);
or U6856 (N_6856,N_6720,N_6698);
and U6857 (N_6857,N_6695,N_6700);
nor U6858 (N_6858,N_6645,N_6795);
nand U6859 (N_6859,N_6786,N_6619);
and U6860 (N_6860,N_6684,N_6666);
and U6861 (N_6861,N_6670,N_6659);
and U6862 (N_6862,N_6643,N_6678);
nor U6863 (N_6863,N_6757,N_6669);
and U6864 (N_6864,N_6650,N_6779);
and U6865 (N_6865,N_6602,N_6634);
or U6866 (N_6866,N_6681,N_6612);
or U6867 (N_6867,N_6662,N_6629);
nand U6868 (N_6868,N_6721,N_6777);
or U6869 (N_6869,N_6606,N_6728);
or U6870 (N_6870,N_6654,N_6676);
and U6871 (N_6871,N_6773,N_6774);
nand U6872 (N_6872,N_6715,N_6617);
nor U6873 (N_6873,N_6709,N_6604);
nor U6874 (N_6874,N_6668,N_6605);
and U6875 (N_6875,N_6775,N_6768);
nand U6876 (N_6876,N_6756,N_6758);
nand U6877 (N_6877,N_6696,N_6732);
nor U6878 (N_6878,N_6694,N_6623);
and U6879 (N_6879,N_6743,N_6767);
or U6880 (N_6880,N_6625,N_6660);
or U6881 (N_6881,N_6794,N_6609);
nor U6882 (N_6882,N_6658,N_6738);
and U6883 (N_6883,N_6648,N_6690);
nand U6884 (N_6884,N_6675,N_6706);
or U6885 (N_6885,N_6740,N_6633);
nor U6886 (N_6886,N_6763,N_6664);
nand U6887 (N_6887,N_6636,N_6736);
nor U6888 (N_6888,N_6677,N_6632);
and U6889 (N_6889,N_6716,N_6686);
nor U6890 (N_6890,N_6799,N_6713);
and U6891 (N_6891,N_6714,N_6747);
and U6892 (N_6892,N_6764,N_6751);
nor U6893 (N_6893,N_6679,N_6753);
and U6894 (N_6894,N_6689,N_6693);
nor U6895 (N_6895,N_6770,N_6615);
nor U6896 (N_6896,N_6613,N_6712);
and U6897 (N_6897,N_6608,N_6610);
nand U6898 (N_6898,N_6759,N_6710);
and U6899 (N_6899,N_6667,N_6749);
nor U6900 (N_6900,N_6609,N_6771);
or U6901 (N_6901,N_6655,N_6709);
nand U6902 (N_6902,N_6751,N_6664);
or U6903 (N_6903,N_6623,N_6796);
or U6904 (N_6904,N_6778,N_6640);
nor U6905 (N_6905,N_6671,N_6659);
nor U6906 (N_6906,N_6754,N_6640);
nor U6907 (N_6907,N_6736,N_6647);
nor U6908 (N_6908,N_6650,N_6656);
or U6909 (N_6909,N_6783,N_6696);
nand U6910 (N_6910,N_6719,N_6740);
or U6911 (N_6911,N_6785,N_6781);
and U6912 (N_6912,N_6685,N_6696);
nor U6913 (N_6913,N_6637,N_6787);
or U6914 (N_6914,N_6750,N_6619);
nand U6915 (N_6915,N_6778,N_6643);
nor U6916 (N_6916,N_6759,N_6610);
nand U6917 (N_6917,N_6777,N_6617);
nor U6918 (N_6918,N_6710,N_6602);
and U6919 (N_6919,N_6716,N_6690);
nand U6920 (N_6920,N_6606,N_6633);
nand U6921 (N_6921,N_6745,N_6603);
and U6922 (N_6922,N_6647,N_6699);
nor U6923 (N_6923,N_6648,N_6667);
or U6924 (N_6924,N_6777,N_6726);
and U6925 (N_6925,N_6788,N_6618);
nor U6926 (N_6926,N_6775,N_6655);
nand U6927 (N_6927,N_6788,N_6629);
and U6928 (N_6928,N_6701,N_6755);
and U6929 (N_6929,N_6748,N_6680);
nor U6930 (N_6930,N_6630,N_6722);
and U6931 (N_6931,N_6729,N_6631);
and U6932 (N_6932,N_6677,N_6627);
and U6933 (N_6933,N_6683,N_6797);
and U6934 (N_6934,N_6656,N_6768);
nor U6935 (N_6935,N_6692,N_6631);
and U6936 (N_6936,N_6785,N_6692);
nor U6937 (N_6937,N_6608,N_6686);
or U6938 (N_6938,N_6616,N_6674);
nand U6939 (N_6939,N_6702,N_6627);
nor U6940 (N_6940,N_6688,N_6636);
or U6941 (N_6941,N_6689,N_6720);
nor U6942 (N_6942,N_6638,N_6721);
nor U6943 (N_6943,N_6694,N_6692);
nand U6944 (N_6944,N_6717,N_6718);
and U6945 (N_6945,N_6655,N_6602);
and U6946 (N_6946,N_6633,N_6619);
or U6947 (N_6947,N_6609,N_6662);
nand U6948 (N_6948,N_6623,N_6684);
or U6949 (N_6949,N_6667,N_6710);
and U6950 (N_6950,N_6760,N_6781);
nand U6951 (N_6951,N_6709,N_6702);
or U6952 (N_6952,N_6793,N_6702);
and U6953 (N_6953,N_6635,N_6616);
nor U6954 (N_6954,N_6715,N_6708);
nand U6955 (N_6955,N_6628,N_6623);
nand U6956 (N_6956,N_6600,N_6784);
or U6957 (N_6957,N_6797,N_6785);
and U6958 (N_6958,N_6629,N_6699);
nor U6959 (N_6959,N_6693,N_6739);
or U6960 (N_6960,N_6793,N_6735);
nand U6961 (N_6961,N_6610,N_6672);
nor U6962 (N_6962,N_6734,N_6711);
nand U6963 (N_6963,N_6651,N_6729);
nor U6964 (N_6964,N_6669,N_6791);
and U6965 (N_6965,N_6685,N_6683);
and U6966 (N_6966,N_6652,N_6727);
nand U6967 (N_6967,N_6692,N_6786);
nand U6968 (N_6968,N_6752,N_6636);
nor U6969 (N_6969,N_6786,N_6714);
and U6970 (N_6970,N_6696,N_6703);
nand U6971 (N_6971,N_6730,N_6642);
nand U6972 (N_6972,N_6634,N_6600);
nor U6973 (N_6973,N_6770,N_6629);
or U6974 (N_6974,N_6760,N_6794);
nand U6975 (N_6975,N_6772,N_6630);
and U6976 (N_6976,N_6751,N_6683);
and U6977 (N_6977,N_6607,N_6622);
and U6978 (N_6978,N_6623,N_6769);
or U6979 (N_6979,N_6691,N_6698);
and U6980 (N_6980,N_6650,N_6712);
nand U6981 (N_6981,N_6779,N_6670);
nand U6982 (N_6982,N_6769,N_6613);
or U6983 (N_6983,N_6659,N_6732);
nand U6984 (N_6984,N_6653,N_6739);
nand U6985 (N_6985,N_6773,N_6753);
or U6986 (N_6986,N_6795,N_6770);
and U6987 (N_6987,N_6719,N_6608);
and U6988 (N_6988,N_6627,N_6610);
nor U6989 (N_6989,N_6690,N_6763);
nor U6990 (N_6990,N_6702,N_6785);
and U6991 (N_6991,N_6723,N_6661);
or U6992 (N_6992,N_6719,N_6791);
nand U6993 (N_6993,N_6785,N_6783);
nor U6994 (N_6994,N_6607,N_6731);
nand U6995 (N_6995,N_6681,N_6715);
and U6996 (N_6996,N_6671,N_6648);
nand U6997 (N_6997,N_6744,N_6685);
or U6998 (N_6998,N_6724,N_6787);
and U6999 (N_6999,N_6688,N_6653);
xnor U7000 (N_7000,N_6845,N_6988);
and U7001 (N_7001,N_6837,N_6867);
and U7002 (N_7002,N_6854,N_6972);
nand U7003 (N_7003,N_6931,N_6907);
nand U7004 (N_7004,N_6834,N_6820);
nor U7005 (N_7005,N_6817,N_6840);
and U7006 (N_7006,N_6804,N_6904);
nor U7007 (N_7007,N_6992,N_6902);
and U7008 (N_7008,N_6938,N_6801);
nand U7009 (N_7009,N_6848,N_6901);
and U7010 (N_7010,N_6940,N_6958);
nor U7011 (N_7011,N_6849,N_6893);
nor U7012 (N_7012,N_6882,N_6960);
or U7013 (N_7013,N_6895,N_6917);
nor U7014 (N_7014,N_6870,N_6855);
or U7015 (N_7015,N_6891,N_6868);
xnor U7016 (N_7016,N_6920,N_6941);
and U7017 (N_7017,N_6825,N_6857);
and U7018 (N_7018,N_6878,N_6873);
nor U7019 (N_7019,N_6957,N_6906);
and U7020 (N_7020,N_6979,N_6853);
and U7021 (N_7021,N_6962,N_6897);
nand U7022 (N_7022,N_6809,N_6954);
or U7023 (N_7023,N_6991,N_6832);
nor U7024 (N_7024,N_6909,N_6952);
or U7025 (N_7025,N_6829,N_6803);
nand U7026 (N_7026,N_6862,N_6885);
nor U7027 (N_7027,N_6861,N_6908);
and U7028 (N_7028,N_6838,N_6926);
xnor U7029 (N_7029,N_6985,N_6919);
nand U7030 (N_7030,N_6953,N_6922);
nand U7031 (N_7031,N_6866,N_6808);
or U7032 (N_7032,N_6852,N_6871);
and U7033 (N_7033,N_6928,N_6971);
nand U7034 (N_7034,N_6977,N_6935);
nand U7035 (N_7035,N_6886,N_6983);
nor U7036 (N_7036,N_6937,N_6943);
nor U7037 (N_7037,N_6858,N_6814);
or U7038 (N_7038,N_6851,N_6823);
xnor U7039 (N_7039,N_6968,N_6948);
nor U7040 (N_7040,N_6827,N_6969);
nand U7041 (N_7041,N_6877,N_6965);
xor U7042 (N_7042,N_6880,N_6973);
nand U7043 (N_7043,N_6869,N_6836);
and U7044 (N_7044,N_6950,N_6815);
nand U7045 (N_7045,N_6876,N_6949);
and U7046 (N_7046,N_6932,N_6924);
nor U7047 (N_7047,N_6864,N_6850);
nor U7048 (N_7048,N_6914,N_6860);
nand U7049 (N_7049,N_6936,N_6989);
or U7050 (N_7050,N_6844,N_6910);
nor U7051 (N_7051,N_6942,N_6822);
nand U7052 (N_7052,N_6955,N_6802);
nor U7053 (N_7053,N_6888,N_6951);
and U7054 (N_7054,N_6974,N_6821);
or U7055 (N_7055,N_6925,N_6806);
nand U7056 (N_7056,N_6921,N_6939);
nor U7057 (N_7057,N_6875,N_6986);
nand U7058 (N_7058,N_6987,N_6903);
nor U7059 (N_7059,N_6830,N_6816);
nand U7060 (N_7060,N_6846,N_6824);
nor U7061 (N_7061,N_6835,N_6923);
and U7062 (N_7062,N_6884,N_6929);
nor U7063 (N_7063,N_6999,N_6915);
nor U7064 (N_7064,N_6982,N_6981);
and U7065 (N_7065,N_6959,N_6990);
nand U7066 (N_7066,N_6847,N_6800);
nand U7067 (N_7067,N_6894,N_6856);
nor U7068 (N_7068,N_6843,N_6934);
and U7069 (N_7069,N_6841,N_6967);
or U7070 (N_7070,N_6899,N_6833);
or U7071 (N_7071,N_6883,N_6993);
or U7072 (N_7072,N_6961,N_6964);
or U7073 (N_7073,N_6811,N_6998);
nor U7074 (N_7074,N_6896,N_6898);
nand U7075 (N_7075,N_6859,N_6912);
or U7076 (N_7076,N_6826,N_6980);
nor U7077 (N_7077,N_6975,N_6916);
or U7078 (N_7078,N_6842,N_6892);
nand U7079 (N_7079,N_6997,N_6887);
and U7080 (N_7080,N_6930,N_6970);
nor U7081 (N_7081,N_6996,N_6818);
or U7082 (N_7082,N_6918,N_6807);
nand U7083 (N_7083,N_6831,N_6881);
or U7084 (N_7084,N_6839,N_6995);
nand U7085 (N_7085,N_6944,N_6865);
or U7086 (N_7086,N_6819,N_6812);
and U7087 (N_7087,N_6805,N_6900);
nand U7088 (N_7088,N_6946,N_6945);
or U7089 (N_7089,N_6984,N_6966);
and U7090 (N_7090,N_6874,N_6994);
and U7091 (N_7091,N_6976,N_6911);
or U7092 (N_7092,N_6890,N_6879);
nor U7093 (N_7093,N_6963,N_6913);
and U7094 (N_7094,N_6947,N_6828);
nor U7095 (N_7095,N_6933,N_6956);
or U7096 (N_7096,N_6889,N_6872);
nand U7097 (N_7097,N_6978,N_6863);
or U7098 (N_7098,N_6813,N_6927);
nor U7099 (N_7099,N_6810,N_6905);
nand U7100 (N_7100,N_6850,N_6997);
and U7101 (N_7101,N_6862,N_6873);
or U7102 (N_7102,N_6853,N_6922);
nand U7103 (N_7103,N_6809,N_6819);
or U7104 (N_7104,N_6826,N_6891);
nor U7105 (N_7105,N_6961,N_6867);
and U7106 (N_7106,N_6898,N_6967);
or U7107 (N_7107,N_6827,N_6980);
nand U7108 (N_7108,N_6933,N_6911);
nor U7109 (N_7109,N_6839,N_6925);
and U7110 (N_7110,N_6958,N_6813);
nor U7111 (N_7111,N_6952,N_6980);
nand U7112 (N_7112,N_6904,N_6823);
and U7113 (N_7113,N_6865,N_6823);
nand U7114 (N_7114,N_6954,N_6870);
or U7115 (N_7115,N_6827,N_6847);
or U7116 (N_7116,N_6834,N_6961);
nor U7117 (N_7117,N_6872,N_6808);
and U7118 (N_7118,N_6954,N_6803);
or U7119 (N_7119,N_6915,N_6880);
and U7120 (N_7120,N_6911,N_6827);
and U7121 (N_7121,N_6802,N_6913);
or U7122 (N_7122,N_6951,N_6880);
nand U7123 (N_7123,N_6925,N_6828);
nor U7124 (N_7124,N_6972,N_6943);
nor U7125 (N_7125,N_6850,N_6936);
and U7126 (N_7126,N_6938,N_6941);
and U7127 (N_7127,N_6920,N_6968);
and U7128 (N_7128,N_6929,N_6994);
and U7129 (N_7129,N_6964,N_6802);
nand U7130 (N_7130,N_6876,N_6861);
nand U7131 (N_7131,N_6852,N_6913);
nor U7132 (N_7132,N_6815,N_6819);
and U7133 (N_7133,N_6837,N_6810);
nor U7134 (N_7134,N_6946,N_6996);
nand U7135 (N_7135,N_6867,N_6809);
nand U7136 (N_7136,N_6834,N_6880);
nand U7137 (N_7137,N_6831,N_6875);
nand U7138 (N_7138,N_6832,N_6911);
nand U7139 (N_7139,N_6955,N_6940);
nor U7140 (N_7140,N_6833,N_6823);
xor U7141 (N_7141,N_6920,N_6966);
nor U7142 (N_7142,N_6864,N_6888);
and U7143 (N_7143,N_6861,N_6824);
and U7144 (N_7144,N_6972,N_6890);
and U7145 (N_7145,N_6938,N_6951);
and U7146 (N_7146,N_6927,N_6984);
or U7147 (N_7147,N_6880,N_6921);
or U7148 (N_7148,N_6807,N_6835);
or U7149 (N_7149,N_6871,N_6961);
nand U7150 (N_7150,N_6830,N_6805);
or U7151 (N_7151,N_6978,N_6911);
or U7152 (N_7152,N_6881,N_6989);
or U7153 (N_7153,N_6904,N_6898);
nand U7154 (N_7154,N_6822,N_6862);
or U7155 (N_7155,N_6995,N_6937);
nand U7156 (N_7156,N_6891,N_6807);
and U7157 (N_7157,N_6851,N_6809);
and U7158 (N_7158,N_6803,N_6889);
or U7159 (N_7159,N_6879,N_6888);
and U7160 (N_7160,N_6812,N_6843);
nand U7161 (N_7161,N_6957,N_6845);
and U7162 (N_7162,N_6977,N_6805);
and U7163 (N_7163,N_6956,N_6934);
or U7164 (N_7164,N_6841,N_6950);
or U7165 (N_7165,N_6966,N_6811);
nand U7166 (N_7166,N_6857,N_6972);
nor U7167 (N_7167,N_6816,N_6823);
or U7168 (N_7168,N_6999,N_6847);
and U7169 (N_7169,N_6885,N_6931);
nand U7170 (N_7170,N_6887,N_6935);
nor U7171 (N_7171,N_6860,N_6807);
nor U7172 (N_7172,N_6878,N_6916);
and U7173 (N_7173,N_6985,N_6969);
nand U7174 (N_7174,N_6845,N_6856);
or U7175 (N_7175,N_6834,N_6948);
nand U7176 (N_7176,N_6916,N_6803);
nand U7177 (N_7177,N_6841,N_6846);
or U7178 (N_7178,N_6915,N_6983);
nor U7179 (N_7179,N_6939,N_6948);
nor U7180 (N_7180,N_6903,N_6939);
and U7181 (N_7181,N_6834,N_6908);
nand U7182 (N_7182,N_6869,N_6948);
nor U7183 (N_7183,N_6857,N_6957);
and U7184 (N_7184,N_6859,N_6928);
and U7185 (N_7185,N_6902,N_6846);
nor U7186 (N_7186,N_6972,N_6856);
nor U7187 (N_7187,N_6828,N_6847);
nand U7188 (N_7188,N_6958,N_6863);
nand U7189 (N_7189,N_6983,N_6830);
nand U7190 (N_7190,N_6900,N_6884);
nor U7191 (N_7191,N_6914,N_6876);
or U7192 (N_7192,N_6893,N_6861);
or U7193 (N_7193,N_6891,N_6984);
or U7194 (N_7194,N_6945,N_6892);
nor U7195 (N_7195,N_6804,N_6802);
or U7196 (N_7196,N_6982,N_6853);
nand U7197 (N_7197,N_6808,N_6827);
xnor U7198 (N_7198,N_6878,N_6818);
and U7199 (N_7199,N_6905,N_6968);
nand U7200 (N_7200,N_7011,N_7147);
nand U7201 (N_7201,N_7197,N_7117);
and U7202 (N_7202,N_7158,N_7019);
nor U7203 (N_7203,N_7068,N_7020);
nand U7204 (N_7204,N_7045,N_7107);
nor U7205 (N_7205,N_7066,N_7067);
or U7206 (N_7206,N_7172,N_7128);
and U7207 (N_7207,N_7086,N_7195);
nor U7208 (N_7208,N_7120,N_7054);
and U7209 (N_7209,N_7143,N_7137);
and U7210 (N_7210,N_7126,N_7094);
nor U7211 (N_7211,N_7159,N_7015);
or U7212 (N_7212,N_7056,N_7186);
or U7213 (N_7213,N_7070,N_7014);
and U7214 (N_7214,N_7129,N_7028);
and U7215 (N_7215,N_7076,N_7050);
nand U7216 (N_7216,N_7079,N_7161);
nor U7217 (N_7217,N_7150,N_7156);
nor U7218 (N_7218,N_7123,N_7182);
and U7219 (N_7219,N_7059,N_7152);
and U7220 (N_7220,N_7113,N_7115);
and U7221 (N_7221,N_7169,N_7187);
and U7222 (N_7222,N_7053,N_7171);
nor U7223 (N_7223,N_7133,N_7101);
xor U7224 (N_7224,N_7127,N_7100);
xnor U7225 (N_7225,N_7191,N_7074);
and U7226 (N_7226,N_7004,N_7151);
and U7227 (N_7227,N_7078,N_7012);
nand U7228 (N_7228,N_7081,N_7130);
nor U7229 (N_7229,N_7092,N_7157);
and U7230 (N_7230,N_7185,N_7052);
nand U7231 (N_7231,N_7064,N_7062);
nor U7232 (N_7232,N_7058,N_7034);
nor U7233 (N_7233,N_7072,N_7088);
or U7234 (N_7234,N_7009,N_7170);
or U7235 (N_7235,N_7047,N_7192);
nand U7236 (N_7236,N_7043,N_7122);
and U7237 (N_7237,N_7046,N_7087);
xor U7238 (N_7238,N_7027,N_7110);
and U7239 (N_7239,N_7167,N_7093);
or U7240 (N_7240,N_7037,N_7132);
or U7241 (N_7241,N_7031,N_7138);
or U7242 (N_7242,N_7099,N_7060);
and U7243 (N_7243,N_7146,N_7044);
nand U7244 (N_7244,N_7173,N_7091);
or U7245 (N_7245,N_7061,N_7085);
or U7246 (N_7246,N_7040,N_7121);
nand U7247 (N_7247,N_7026,N_7109);
nand U7248 (N_7248,N_7055,N_7175);
nand U7249 (N_7249,N_7112,N_7057);
nor U7250 (N_7250,N_7084,N_7154);
nand U7251 (N_7251,N_7160,N_7017);
nand U7252 (N_7252,N_7166,N_7136);
and U7253 (N_7253,N_7089,N_7035);
nor U7254 (N_7254,N_7118,N_7003);
nand U7255 (N_7255,N_7111,N_7025);
nand U7256 (N_7256,N_7139,N_7069);
nand U7257 (N_7257,N_7194,N_7001);
nand U7258 (N_7258,N_7134,N_7010);
or U7259 (N_7259,N_7108,N_7131);
and U7260 (N_7260,N_7071,N_7005);
or U7261 (N_7261,N_7145,N_7181);
nor U7262 (N_7262,N_7022,N_7164);
nand U7263 (N_7263,N_7021,N_7163);
or U7264 (N_7264,N_7080,N_7180);
or U7265 (N_7265,N_7174,N_7189);
and U7266 (N_7266,N_7063,N_7188);
nand U7267 (N_7267,N_7153,N_7165);
nand U7268 (N_7268,N_7105,N_7168);
nor U7269 (N_7269,N_7075,N_7190);
nor U7270 (N_7270,N_7024,N_7162);
xnor U7271 (N_7271,N_7032,N_7103);
and U7272 (N_7272,N_7023,N_7178);
or U7273 (N_7273,N_7007,N_7198);
nor U7274 (N_7274,N_7102,N_7048);
or U7275 (N_7275,N_7140,N_7098);
and U7276 (N_7276,N_7038,N_7016);
nor U7277 (N_7277,N_7142,N_7196);
or U7278 (N_7278,N_7090,N_7013);
and U7279 (N_7279,N_7051,N_7018);
nor U7280 (N_7280,N_7155,N_7199);
and U7281 (N_7281,N_7116,N_7030);
xnor U7282 (N_7282,N_7124,N_7049);
nor U7283 (N_7283,N_7095,N_7036);
and U7284 (N_7284,N_7082,N_7135);
nand U7285 (N_7285,N_7119,N_7097);
and U7286 (N_7286,N_7104,N_7183);
nor U7287 (N_7287,N_7125,N_7073);
nand U7288 (N_7288,N_7065,N_7106);
and U7289 (N_7289,N_7008,N_7149);
and U7290 (N_7290,N_7077,N_7141);
and U7291 (N_7291,N_7148,N_7083);
nor U7292 (N_7292,N_7096,N_7184);
or U7293 (N_7293,N_7006,N_7144);
nor U7294 (N_7294,N_7179,N_7029);
nor U7295 (N_7295,N_7000,N_7039);
nor U7296 (N_7296,N_7176,N_7033);
nand U7297 (N_7297,N_7002,N_7177);
and U7298 (N_7298,N_7041,N_7114);
or U7299 (N_7299,N_7042,N_7193);
nor U7300 (N_7300,N_7034,N_7002);
nand U7301 (N_7301,N_7019,N_7151);
nor U7302 (N_7302,N_7174,N_7159);
or U7303 (N_7303,N_7097,N_7152);
nand U7304 (N_7304,N_7000,N_7038);
nor U7305 (N_7305,N_7153,N_7191);
nand U7306 (N_7306,N_7044,N_7096);
nand U7307 (N_7307,N_7118,N_7039);
nand U7308 (N_7308,N_7031,N_7130);
and U7309 (N_7309,N_7161,N_7018);
nor U7310 (N_7310,N_7102,N_7148);
nor U7311 (N_7311,N_7061,N_7052);
nand U7312 (N_7312,N_7029,N_7149);
and U7313 (N_7313,N_7123,N_7025);
or U7314 (N_7314,N_7037,N_7171);
or U7315 (N_7315,N_7085,N_7033);
or U7316 (N_7316,N_7141,N_7109);
nand U7317 (N_7317,N_7091,N_7031);
nor U7318 (N_7318,N_7031,N_7089);
nor U7319 (N_7319,N_7118,N_7052);
or U7320 (N_7320,N_7118,N_7037);
nand U7321 (N_7321,N_7061,N_7089);
or U7322 (N_7322,N_7027,N_7017);
or U7323 (N_7323,N_7138,N_7114);
and U7324 (N_7324,N_7185,N_7159);
nor U7325 (N_7325,N_7109,N_7025);
nand U7326 (N_7326,N_7061,N_7110);
and U7327 (N_7327,N_7150,N_7023);
or U7328 (N_7328,N_7137,N_7123);
or U7329 (N_7329,N_7062,N_7138);
nand U7330 (N_7330,N_7197,N_7198);
and U7331 (N_7331,N_7141,N_7139);
nand U7332 (N_7332,N_7128,N_7174);
or U7333 (N_7333,N_7196,N_7192);
or U7334 (N_7334,N_7073,N_7184);
or U7335 (N_7335,N_7017,N_7134);
nor U7336 (N_7336,N_7000,N_7027);
and U7337 (N_7337,N_7154,N_7166);
nand U7338 (N_7338,N_7189,N_7034);
nand U7339 (N_7339,N_7124,N_7043);
and U7340 (N_7340,N_7073,N_7180);
nand U7341 (N_7341,N_7099,N_7190);
and U7342 (N_7342,N_7063,N_7038);
or U7343 (N_7343,N_7134,N_7008);
and U7344 (N_7344,N_7069,N_7050);
and U7345 (N_7345,N_7143,N_7103);
or U7346 (N_7346,N_7038,N_7012);
nand U7347 (N_7347,N_7024,N_7173);
nand U7348 (N_7348,N_7199,N_7106);
nand U7349 (N_7349,N_7082,N_7168);
or U7350 (N_7350,N_7162,N_7080);
nand U7351 (N_7351,N_7109,N_7042);
nor U7352 (N_7352,N_7120,N_7142);
nor U7353 (N_7353,N_7061,N_7088);
nand U7354 (N_7354,N_7105,N_7145);
nand U7355 (N_7355,N_7185,N_7069);
or U7356 (N_7356,N_7014,N_7137);
or U7357 (N_7357,N_7097,N_7189);
nand U7358 (N_7358,N_7122,N_7132);
or U7359 (N_7359,N_7193,N_7060);
and U7360 (N_7360,N_7121,N_7080);
nand U7361 (N_7361,N_7114,N_7053);
nand U7362 (N_7362,N_7057,N_7161);
and U7363 (N_7363,N_7102,N_7138);
nand U7364 (N_7364,N_7054,N_7086);
or U7365 (N_7365,N_7045,N_7168);
nand U7366 (N_7366,N_7046,N_7101);
nor U7367 (N_7367,N_7122,N_7098);
nand U7368 (N_7368,N_7033,N_7045);
or U7369 (N_7369,N_7037,N_7060);
and U7370 (N_7370,N_7180,N_7054);
or U7371 (N_7371,N_7015,N_7120);
nor U7372 (N_7372,N_7191,N_7131);
or U7373 (N_7373,N_7139,N_7042);
nand U7374 (N_7374,N_7147,N_7191);
or U7375 (N_7375,N_7031,N_7129);
and U7376 (N_7376,N_7046,N_7157);
and U7377 (N_7377,N_7094,N_7011);
and U7378 (N_7378,N_7132,N_7098);
nand U7379 (N_7379,N_7009,N_7162);
and U7380 (N_7380,N_7138,N_7016);
nor U7381 (N_7381,N_7121,N_7056);
or U7382 (N_7382,N_7026,N_7113);
nor U7383 (N_7383,N_7133,N_7151);
or U7384 (N_7384,N_7166,N_7193);
and U7385 (N_7385,N_7139,N_7006);
or U7386 (N_7386,N_7018,N_7169);
and U7387 (N_7387,N_7168,N_7187);
and U7388 (N_7388,N_7007,N_7062);
nand U7389 (N_7389,N_7131,N_7126);
nand U7390 (N_7390,N_7184,N_7105);
nor U7391 (N_7391,N_7054,N_7134);
nand U7392 (N_7392,N_7062,N_7123);
nor U7393 (N_7393,N_7101,N_7165);
and U7394 (N_7394,N_7092,N_7082);
or U7395 (N_7395,N_7019,N_7199);
and U7396 (N_7396,N_7004,N_7024);
or U7397 (N_7397,N_7107,N_7197);
nand U7398 (N_7398,N_7013,N_7124);
nand U7399 (N_7399,N_7054,N_7179);
nor U7400 (N_7400,N_7202,N_7362);
nand U7401 (N_7401,N_7216,N_7353);
or U7402 (N_7402,N_7336,N_7373);
nand U7403 (N_7403,N_7225,N_7276);
nor U7404 (N_7404,N_7301,N_7339);
nor U7405 (N_7405,N_7283,N_7228);
or U7406 (N_7406,N_7309,N_7382);
nand U7407 (N_7407,N_7314,N_7331);
nor U7408 (N_7408,N_7380,N_7335);
or U7409 (N_7409,N_7308,N_7247);
nand U7410 (N_7410,N_7281,N_7233);
or U7411 (N_7411,N_7295,N_7240);
or U7412 (N_7412,N_7359,N_7347);
nor U7413 (N_7413,N_7213,N_7252);
nor U7414 (N_7414,N_7393,N_7268);
nand U7415 (N_7415,N_7291,N_7368);
and U7416 (N_7416,N_7248,N_7200);
or U7417 (N_7417,N_7263,N_7348);
or U7418 (N_7418,N_7260,N_7390);
and U7419 (N_7419,N_7386,N_7311);
nand U7420 (N_7420,N_7246,N_7285);
nor U7421 (N_7421,N_7304,N_7303);
nand U7422 (N_7422,N_7375,N_7284);
or U7423 (N_7423,N_7215,N_7273);
and U7424 (N_7424,N_7383,N_7267);
or U7425 (N_7425,N_7385,N_7349);
nand U7426 (N_7426,N_7312,N_7324);
and U7427 (N_7427,N_7230,N_7365);
or U7428 (N_7428,N_7346,N_7381);
nand U7429 (N_7429,N_7224,N_7302);
or U7430 (N_7430,N_7351,N_7364);
or U7431 (N_7431,N_7379,N_7210);
or U7432 (N_7432,N_7376,N_7222);
nor U7433 (N_7433,N_7374,N_7259);
nor U7434 (N_7434,N_7395,N_7378);
nand U7435 (N_7435,N_7398,N_7234);
and U7436 (N_7436,N_7226,N_7323);
nand U7437 (N_7437,N_7341,N_7297);
nor U7438 (N_7438,N_7372,N_7358);
nand U7439 (N_7439,N_7371,N_7271);
or U7440 (N_7440,N_7287,N_7206);
xnor U7441 (N_7441,N_7217,N_7275);
or U7442 (N_7442,N_7277,N_7214);
nor U7443 (N_7443,N_7329,N_7249);
nor U7444 (N_7444,N_7211,N_7239);
nand U7445 (N_7445,N_7265,N_7257);
or U7446 (N_7446,N_7310,N_7299);
nor U7447 (N_7447,N_7332,N_7356);
and U7448 (N_7448,N_7327,N_7369);
nand U7449 (N_7449,N_7363,N_7366);
xnor U7450 (N_7450,N_7212,N_7337);
or U7451 (N_7451,N_7218,N_7318);
and U7452 (N_7452,N_7392,N_7333);
nor U7453 (N_7453,N_7242,N_7231);
or U7454 (N_7454,N_7221,N_7288);
nor U7455 (N_7455,N_7223,N_7317);
and U7456 (N_7456,N_7296,N_7399);
and U7457 (N_7457,N_7269,N_7328);
or U7458 (N_7458,N_7290,N_7227);
and U7459 (N_7459,N_7289,N_7278);
nand U7460 (N_7460,N_7298,N_7326);
nor U7461 (N_7461,N_7229,N_7321);
nor U7462 (N_7462,N_7220,N_7342);
or U7463 (N_7463,N_7207,N_7274);
nand U7464 (N_7464,N_7319,N_7305);
and U7465 (N_7465,N_7261,N_7262);
nor U7466 (N_7466,N_7243,N_7258);
nor U7467 (N_7467,N_7279,N_7235);
xor U7468 (N_7468,N_7397,N_7241);
and U7469 (N_7469,N_7357,N_7270);
nand U7470 (N_7470,N_7345,N_7264);
nand U7471 (N_7471,N_7313,N_7388);
or U7472 (N_7472,N_7354,N_7244);
nor U7473 (N_7473,N_7236,N_7316);
and U7474 (N_7474,N_7255,N_7350);
or U7475 (N_7475,N_7306,N_7237);
and U7476 (N_7476,N_7389,N_7338);
nor U7477 (N_7477,N_7394,N_7387);
or U7478 (N_7478,N_7343,N_7396);
and U7479 (N_7479,N_7293,N_7219);
nand U7480 (N_7480,N_7204,N_7292);
nor U7481 (N_7481,N_7205,N_7251);
nor U7482 (N_7482,N_7370,N_7209);
and U7483 (N_7483,N_7377,N_7232);
nand U7484 (N_7484,N_7360,N_7344);
nor U7485 (N_7485,N_7245,N_7367);
nand U7486 (N_7486,N_7325,N_7361);
or U7487 (N_7487,N_7280,N_7355);
or U7488 (N_7488,N_7334,N_7256);
and U7489 (N_7489,N_7208,N_7286);
nand U7490 (N_7490,N_7266,N_7315);
nand U7491 (N_7491,N_7201,N_7391);
nor U7492 (N_7492,N_7352,N_7282);
nor U7493 (N_7493,N_7253,N_7320);
and U7494 (N_7494,N_7238,N_7330);
nor U7495 (N_7495,N_7384,N_7203);
nand U7496 (N_7496,N_7254,N_7250);
or U7497 (N_7497,N_7340,N_7322);
nand U7498 (N_7498,N_7294,N_7272);
nand U7499 (N_7499,N_7300,N_7307);
and U7500 (N_7500,N_7395,N_7379);
or U7501 (N_7501,N_7340,N_7215);
nor U7502 (N_7502,N_7391,N_7266);
nand U7503 (N_7503,N_7381,N_7280);
or U7504 (N_7504,N_7394,N_7291);
and U7505 (N_7505,N_7229,N_7349);
nor U7506 (N_7506,N_7204,N_7227);
and U7507 (N_7507,N_7342,N_7242);
or U7508 (N_7508,N_7378,N_7384);
nor U7509 (N_7509,N_7296,N_7298);
and U7510 (N_7510,N_7397,N_7295);
nor U7511 (N_7511,N_7277,N_7335);
nand U7512 (N_7512,N_7260,N_7234);
and U7513 (N_7513,N_7275,N_7350);
and U7514 (N_7514,N_7271,N_7384);
or U7515 (N_7515,N_7379,N_7399);
nor U7516 (N_7516,N_7396,N_7276);
and U7517 (N_7517,N_7358,N_7320);
nor U7518 (N_7518,N_7313,N_7302);
or U7519 (N_7519,N_7349,N_7364);
or U7520 (N_7520,N_7345,N_7218);
and U7521 (N_7521,N_7399,N_7277);
and U7522 (N_7522,N_7211,N_7380);
or U7523 (N_7523,N_7343,N_7313);
nand U7524 (N_7524,N_7219,N_7201);
or U7525 (N_7525,N_7219,N_7262);
nand U7526 (N_7526,N_7237,N_7256);
nor U7527 (N_7527,N_7386,N_7383);
or U7528 (N_7528,N_7203,N_7207);
nand U7529 (N_7529,N_7271,N_7219);
and U7530 (N_7530,N_7334,N_7394);
nor U7531 (N_7531,N_7300,N_7345);
xor U7532 (N_7532,N_7239,N_7339);
or U7533 (N_7533,N_7254,N_7223);
or U7534 (N_7534,N_7307,N_7380);
or U7535 (N_7535,N_7244,N_7376);
or U7536 (N_7536,N_7368,N_7369);
and U7537 (N_7537,N_7397,N_7237);
or U7538 (N_7538,N_7320,N_7237);
nor U7539 (N_7539,N_7329,N_7256);
nand U7540 (N_7540,N_7250,N_7209);
or U7541 (N_7541,N_7356,N_7213);
or U7542 (N_7542,N_7203,N_7302);
or U7543 (N_7543,N_7301,N_7246);
xor U7544 (N_7544,N_7322,N_7235);
nor U7545 (N_7545,N_7286,N_7260);
or U7546 (N_7546,N_7261,N_7371);
nor U7547 (N_7547,N_7352,N_7244);
or U7548 (N_7548,N_7325,N_7249);
and U7549 (N_7549,N_7399,N_7249);
nor U7550 (N_7550,N_7249,N_7264);
and U7551 (N_7551,N_7219,N_7291);
nor U7552 (N_7552,N_7305,N_7257);
or U7553 (N_7553,N_7200,N_7297);
nor U7554 (N_7554,N_7344,N_7353);
nor U7555 (N_7555,N_7376,N_7299);
and U7556 (N_7556,N_7289,N_7223);
nand U7557 (N_7557,N_7314,N_7225);
or U7558 (N_7558,N_7235,N_7282);
nand U7559 (N_7559,N_7376,N_7214);
nand U7560 (N_7560,N_7235,N_7396);
and U7561 (N_7561,N_7385,N_7201);
nor U7562 (N_7562,N_7344,N_7202);
and U7563 (N_7563,N_7277,N_7269);
nand U7564 (N_7564,N_7317,N_7307);
and U7565 (N_7565,N_7205,N_7336);
and U7566 (N_7566,N_7260,N_7268);
or U7567 (N_7567,N_7260,N_7211);
or U7568 (N_7568,N_7264,N_7323);
nor U7569 (N_7569,N_7260,N_7389);
and U7570 (N_7570,N_7330,N_7365);
nor U7571 (N_7571,N_7257,N_7208);
nand U7572 (N_7572,N_7315,N_7323);
or U7573 (N_7573,N_7258,N_7223);
or U7574 (N_7574,N_7330,N_7350);
nand U7575 (N_7575,N_7331,N_7340);
xnor U7576 (N_7576,N_7363,N_7238);
and U7577 (N_7577,N_7386,N_7325);
or U7578 (N_7578,N_7230,N_7213);
nor U7579 (N_7579,N_7378,N_7370);
and U7580 (N_7580,N_7337,N_7265);
nand U7581 (N_7581,N_7398,N_7253);
nor U7582 (N_7582,N_7233,N_7226);
nand U7583 (N_7583,N_7281,N_7204);
or U7584 (N_7584,N_7388,N_7253);
and U7585 (N_7585,N_7274,N_7303);
nor U7586 (N_7586,N_7203,N_7296);
and U7587 (N_7587,N_7356,N_7339);
nand U7588 (N_7588,N_7292,N_7250);
nor U7589 (N_7589,N_7247,N_7217);
nor U7590 (N_7590,N_7241,N_7381);
and U7591 (N_7591,N_7216,N_7376);
nand U7592 (N_7592,N_7344,N_7204);
xnor U7593 (N_7593,N_7245,N_7279);
nand U7594 (N_7594,N_7312,N_7392);
and U7595 (N_7595,N_7349,N_7218);
nor U7596 (N_7596,N_7348,N_7362);
nand U7597 (N_7597,N_7304,N_7258);
nor U7598 (N_7598,N_7228,N_7328);
or U7599 (N_7599,N_7393,N_7399);
nor U7600 (N_7600,N_7400,N_7416);
nor U7601 (N_7601,N_7485,N_7508);
or U7602 (N_7602,N_7598,N_7596);
nor U7603 (N_7603,N_7501,N_7449);
and U7604 (N_7604,N_7479,N_7504);
and U7605 (N_7605,N_7424,N_7438);
nand U7606 (N_7606,N_7537,N_7455);
or U7607 (N_7607,N_7489,N_7505);
and U7608 (N_7608,N_7588,N_7576);
nand U7609 (N_7609,N_7522,N_7413);
and U7610 (N_7610,N_7402,N_7597);
nor U7611 (N_7611,N_7414,N_7519);
or U7612 (N_7612,N_7443,N_7446);
and U7613 (N_7613,N_7401,N_7442);
nand U7614 (N_7614,N_7492,N_7549);
or U7615 (N_7615,N_7439,N_7408);
and U7616 (N_7616,N_7564,N_7570);
nand U7617 (N_7617,N_7429,N_7534);
and U7618 (N_7618,N_7499,N_7465);
or U7619 (N_7619,N_7419,N_7430);
nand U7620 (N_7620,N_7454,N_7582);
nor U7621 (N_7621,N_7587,N_7433);
or U7622 (N_7622,N_7517,N_7420);
nor U7623 (N_7623,N_7553,N_7432);
nand U7624 (N_7624,N_7525,N_7556);
or U7625 (N_7625,N_7417,N_7536);
nand U7626 (N_7626,N_7487,N_7476);
nand U7627 (N_7627,N_7464,N_7494);
or U7628 (N_7628,N_7579,N_7410);
or U7629 (N_7629,N_7589,N_7561);
nor U7630 (N_7630,N_7523,N_7569);
xor U7631 (N_7631,N_7542,N_7510);
nand U7632 (N_7632,N_7447,N_7486);
nand U7633 (N_7633,N_7571,N_7456);
and U7634 (N_7634,N_7593,N_7546);
nor U7635 (N_7635,N_7541,N_7547);
nand U7636 (N_7636,N_7452,N_7490);
nor U7637 (N_7637,N_7488,N_7491);
or U7638 (N_7638,N_7484,N_7471);
and U7639 (N_7639,N_7509,N_7441);
nand U7640 (N_7640,N_7535,N_7544);
and U7641 (N_7641,N_7437,N_7466);
nand U7642 (N_7642,N_7403,N_7532);
nor U7643 (N_7643,N_7468,N_7451);
nor U7644 (N_7644,N_7574,N_7426);
and U7645 (N_7645,N_7469,N_7462);
or U7646 (N_7646,N_7592,N_7458);
or U7647 (N_7647,N_7473,N_7467);
nor U7648 (N_7648,N_7533,N_7497);
and U7649 (N_7649,N_7436,N_7459);
and U7650 (N_7650,N_7415,N_7503);
or U7651 (N_7651,N_7545,N_7568);
and U7652 (N_7652,N_7445,N_7538);
and U7653 (N_7653,N_7552,N_7453);
nand U7654 (N_7654,N_7421,N_7422);
and U7655 (N_7655,N_7411,N_7590);
nand U7656 (N_7656,N_7506,N_7515);
nand U7657 (N_7657,N_7493,N_7512);
nand U7658 (N_7658,N_7483,N_7584);
and U7659 (N_7659,N_7594,N_7527);
and U7660 (N_7660,N_7528,N_7550);
nor U7661 (N_7661,N_7435,N_7406);
nor U7662 (N_7662,N_7502,N_7412);
nand U7663 (N_7663,N_7575,N_7585);
nor U7664 (N_7664,N_7562,N_7511);
nand U7665 (N_7665,N_7434,N_7428);
and U7666 (N_7666,N_7591,N_7521);
nor U7667 (N_7667,N_7495,N_7478);
nand U7668 (N_7668,N_7470,N_7480);
and U7669 (N_7669,N_7477,N_7460);
or U7670 (N_7670,N_7516,N_7539);
nor U7671 (N_7671,N_7404,N_7444);
or U7672 (N_7672,N_7496,N_7405);
or U7673 (N_7673,N_7457,N_7448);
nand U7674 (N_7674,N_7431,N_7409);
nor U7675 (N_7675,N_7572,N_7578);
or U7676 (N_7676,N_7583,N_7560);
or U7677 (N_7677,N_7530,N_7599);
nand U7678 (N_7678,N_7543,N_7540);
and U7679 (N_7679,N_7440,N_7472);
and U7680 (N_7680,N_7461,N_7595);
nor U7681 (N_7681,N_7463,N_7520);
nor U7682 (N_7682,N_7555,N_7482);
and U7683 (N_7683,N_7567,N_7514);
and U7684 (N_7684,N_7425,N_7551);
and U7685 (N_7685,N_7581,N_7481);
nand U7686 (N_7686,N_7548,N_7475);
nand U7687 (N_7687,N_7498,N_7531);
nor U7688 (N_7688,N_7580,N_7423);
nor U7689 (N_7689,N_7577,N_7565);
nor U7690 (N_7690,N_7558,N_7586);
nand U7691 (N_7691,N_7524,N_7474);
or U7692 (N_7692,N_7559,N_7529);
nor U7693 (N_7693,N_7518,N_7407);
nor U7694 (N_7694,N_7500,N_7554);
nand U7695 (N_7695,N_7507,N_7563);
or U7696 (N_7696,N_7526,N_7513);
nand U7697 (N_7697,N_7418,N_7557);
nor U7698 (N_7698,N_7566,N_7427);
and U7699 (N_7699,N_7573,N_7450);
and U7700 (N_7700,N_7473,N_7417);
or U7701 (N_7701,N_7430,N_7467);
and U7702 (N_7702,N_7533,N_7578);
or U7703 (N_7703,N_7518,N_7553);
nor U7704 (N_7704,N_7427,N_7449);
nand U7705 (N_7705,N_7465,N_7464);
or U7706 (N_7706,N_7407,N_7415);
and U7707 (N_7707,N_7502,N_7526);
nand U7708 (N_7708,N_7548,N_7420);
or U7709 (N_7709,N_7452,N_7492);
or U7710 (N_7710,N_7575,N_7441);
nand U7711 (N_7711,N_7401,N_7597);
nor U7712 (N_7712,N_7481,N_7573);
nand U7713 (N_7713,N_7416,N_7415);
nor U7714 (N_7714,N_7526,N_7444);
or U7715 (N_7715,N_7470,N_7599);
and U7716 (N_7716,N_7482,N_7417);
and U7717 (N_7717,N_7503,N_7495);
and U7718 (N_7718,N_7448,N_7507);
nand U7719 (N_7719,N_7415,N_7540);
nor U7720 (N_7720,N_7464,N_7507);
and U7721 (N_7721,N_7544,N_7522);
nand U7722 (N_7722,N_7574,N_7440);
or U7723 (N_7723,N_7524,N_7407);
nor U7724 (N_7724,N_7557,N_7452);
and U7725 (N_7725,N_7449,N_7490);
nand U7726 (N_7726,N_7528,N_7515);
nand U7727 (N_7727,N_7577,N_7423);
nand U7728 (N_7728,N_7585,N_7593);
or U7729 (N_7729,N_7513,N_7520);
nor U7730 (N_7730,N_7507,N_7402);
nand U7731 (N_7731,N_7543,N_7437);
and U7732 (N_7732,N_7566,N_7525);
nor U7733 (N_7733,N_7484,N_7404);
and U7734 (N_7734,N_7581,N_7559);
nor U7735 (N_7735,N_7489,N_7439);
nand U7736 (N_7736,N_7559,N_7572);
and U7737 (N_7737,N_7427,N_7435);
and U7738 (N_7738,N_7448,N_7464);
nor U7739 (N_7739,N_7591,N_7425);
or U7740 (N_7740,N_7561,N_7513);
or U7741 (N_7741,N_7407,N_7564);
or U7742 (N_7742,N_7490,N_7539);
nand U7743 (N_7743,N_7458,N_7594);
nand U7744 (N_7744,N_7473,N_7498);
and U7745 (N_7745,N_7546,N_7523);
nor U7746 (N_7746,N_7451,N_7599);
nand U7747 (N_7747,N_7431,N_7530);
and U7748 (N_7748,N_7445,N_7401);
xor U7749 (N_7749,N_7493,N_7449);
and U7750 (N_7750,N_7528,N_7541);
or U7751 (N_7751,N_7475,N_7447);
and U7752 (N_7752,N_7479,N_7550);
nor U7753 (N_7753,N_7458,N_7508);
nor U7754 (N_7754,N_7458,N_7507);
xnor U7755 (N_7755,N_7538,N_7585);
or U7756 (N_7756,N_7531,N_7522);
and U7757 (N_7757,N_7557,N_7571);
or U7758 (N_7758,N_7586,N_7428);
or U7759 (N_7759,N_7507,N_7574);
nor U7760 (N_7760,N_7558,N_7543);
nand U7761 (N_7761,N_7435,N_7544);
nand U7762 (N_7762,N_7402,N_7541);
nand U7763 (N_7763,N_7401,N_7499);
nand U7764 (N_7764,N_7400,N_7422);
nor U7765 (N_7765,N_7592,N_7566);
or U7766 (N_7766,N_7483,N_7490);
nand U7767 (N_7767,N_7579,N_7586);
or U7768 (N_7768,N_7515,N_7465);
nor U7769 (N_7769,N_7553,N_7573);
nor U7770 (N_7770,N_7565,N_7544);
nand U7771 (N_7771,N_7539,N_7521);
or U7772 (N_7772,N_7567,N_7590);
nor U7773 (N_7773,N_7494,N_7590);
nor U7774 (N_7774,N_7453,N_7486);
nand U7775 (N_7775,N_7563,N_7424);
nor U7776 (N_7776,N_7426,N_7443);
nor U7777 (N_7777,N_7579,N_7447);
nand U7778 (N_7778,N_7425,N_7568);
or U7779 (N_7779,N_7517,N_7486);
nor U7780 (N_7780,N_7580,N_7449);
nand U7781 (N_7781,N_7564,N_7424);
and U7782 (N_7782,N_7448,N_7499);
nor U7783 (N_7783,N_7460,N_7433);
nand U7784 (N_7784,N_7487,N_7496);
or U7785 (N_7785,N_7555,N_7556);
nor U7786 (N_7786,N_7556,N_7539);
nor U7787 (N_7787,N_7519,N_7596);
nand U7788 (N_7788,N_7514,N_7484);
and U7789 (N_7789,N_7420,N_7594);
or U7790 (N_7790,N_7575,N_7517);
nor U7791 (N_7791,N_7495,N_7538);
or U7792 (N_7792,N_7425,N_7497);
and U7793 (N_7793,N_7428,N_7499);
and U7794 (N_7794,N_7404,N_7424);
or U7795 (N_7795,N_7440,N_7534);
nor U7796 (N_7796,N_7400,N_7473);
nor U7797 (N_7797,N_7511,N_7587);
nor U7798 (N_7798,N_7583,N_7588);
or U7799 (N_7799,N_7583,N_7547);
nor U7800 (N_7800,N_7701,N_7763);
nand U7801 (N_7801,N_7618,N_7705);
nand U7802 (N_7802,N_7648,N_7706);
or U7803 (N_7803,N_7780,N_7777);
nand U7804 (N_7804,N_7622,N_7770);
and U7805 (N_7805,N_7782,N_7781);
or U7806 (N_7806,N_7792,N_7734);
and U7807 (N_7807,N_7634,N_7649);
or U7808 (N_7808,N_7604,N_7756);
nand U7809 (N_7809,N_7656,N_7657);
nand U7810 (N_7810,N_7779,N_7762);
nand U7811 (N_7811,N_7717,N_7644);
or U7812 (N_7812,N_7747,N_7632);
nor U7813 (N_7813,N_7676,N_7776);
nor U7814 (N_7814,N_7736,N_7645);
and U7815 (N_7815,N_7744,N_7673);
or U7816 (N_7816,N_7708,N_7670);
and U7817 (N_7817,N_7628,N_7797);
or U7818 (N_7818,N_7669,N_7684);
nor U7819 (N_7819,N_7752,N_7601);
nor U7820 (N_7820,N_7778,N_7619);
or U7821 (N_7821,N_7691,N_7715);
nor U7822 (N_7822,N_7603,N_7758);
and U7823 (N_7823,N_7681,N_7600);
and U7824 (N_7824,N_7652,N_7639);
or U7825 (N_7825,N_7612,N_7726);
nand U7826 (N_7826,N_7703,N_7740);
and U7827 (N_7827,N_7650,N_7651);
nor U7828 (N_7828,N_7727,N_7694);
nand U7829 (N_7829,N_7700,N_7606);
nor U7830 (N_7830,N_7718,N_7682);
nand U7831 (N_7831,N_7624,N_7610);
nor U7832 (N_7832,N_7794,N_7766);
or U7833 (N_7833,N_7623,N_7605);
nand U7834 (N_7834,N_7641,N_7668);
or U7835 (N_7835,N_7689,N_7754);
or U7836 (N_7836,N_7633,N_7637);
or U7837 (N_7837,N_7602,N_7755);
and U7838 (N_7838,N_7742,N_7661);
xor U7839 (N_7839,N_7768,N_7646);
nand U7840 (N_7840,N_7728,N_7743);
nand U7841 (N_7841,N_7765,N_7720);
nor U7842 (N_7842,N_7731,N_7749);
or U7843 (N_7843,N_7722,N_7757);
and U7844 (N_7844,N_7616,N_7741);
or U7845 (N_7845,N_7738,N_7793);
or U7846 (N_7846,N_7611,N_7786);
nor U7847 (N_7847,N_7729,N_7721);
and U7848 (N_7848,N_7697,N_7658);
and U7849 (N_7849,N_7638,N_7745);
nor U7850 (N_7850,N_7693,N_7685);
or U7851 (N_7851,N_7635,N_7653);
nand U7852 (N_7852,N_7680,N_7699);
nor U7853 (N_7853,N_7716,N_7774);
nand U7854 (N_7854,N_7772,N_7615);
nor U7855 (N_7855,N_7631,N_7704);
or U7856 (N_7856,N_7698,N_7788);
nor U7857 (N_7857,N_7709,N_7679);
or U7858 (N_7858,N_7664,N_7674);
nor U7859 (N_7859,N_7724,N_7672);
nand U7860 (N_7860,N_7712,N_7753);
and U7861 (N_7861,N_7733,N_7764);
and U7862 (N_7862,N_7710,N_7723);
nand U7863 (N_7863,N_7789,N_7769);
nor U7864 (N_7864,N_7730,N_7785);
nand U7865 (N_7865,N_7771,N_7750);
nand U7866 (N_7866,N_7714,N_7751);
nor U7867 (N_7867,N_7671,N_7795);
or U7868 (N_7868,N_7799,N_7692);
nand U7869 (N_7869,N_7607,N_7688);
nor U7870 (N_7870,N_7783,N_7663);
nor U7871 (N_7871,N_7640,N_7630);
or U7872 (N_7872,N_7767,N_7735);
and U7873 (N_7873,N_7614,N_7654);
or U7874 (N_7874,N_7719,N_7609);
xnor U7875 (N_7875,N_7761,N_7675);
and U7876 (N_7876,N_7713,N_7647);
nor U7877 (N_7877,N_7690,N_7760);
nor U7878 (N_7878,N_7711,N_7620);
and U7879 (N_7879,N_7791,N_7642);
or U7880 (N_7880,N_7798,N_7655);
and U7881 (N_7881,N_7683,N_7626);
or U7882 (N_7882,N_7790,N_7696);
and U7883 (N_7883,N_7737,N_7677);
and U7884 (N_7884,N_7643,N_7732);
and U7885 (N_7885,N_7667,N_7666);
and U7886 (N_7886,N_7659,N_7787);
and U7887 (N_7887,N_7739,N_7707);
or U7888 (N_7888,N_7678,N_7759);
or U7889 (N_7889,N_7660,N_7746);
nand U7890 (N_7890,N_7662,N_7686);
or U7891 (N_7891,N_7625,N_7627);
nand U7892 (N_7892,N_7784,N_7725);
xor U7893 (N_7893,N_7613,N_7621);
and U7894 (N_7894,N_7796,N_7636);
or U7895 (N_7895,N_7608,N_7687);
or U7896 (N_7896,N_7773,N_7702);
nand U7897 (N_7897,N_7748,N_7695);
or U7898 (N_7898,N_7629,N_7665);
nor U7899 (N_7899,N_7617,N_7775);
nor U7900 (N_7900,N_7627,N_7692);
nor U7901 (N_7901,N_7759,N_7790);
nand U7902 (N_7902,N_7643,N_7668);
and U7903 (N_7903,N_7680,N_7738);
or U7904 (N_7904,N_7619,N_7787);
nand U7905 (N_7905,N_7626,N_7718);
or U7906 (N_7906,N_7790,N_7633);
nand U7907 (N_7907,N_7662,N_7621);
nor U7908 (N_7908,N_7658,N_7770);
nor U7909 (N_7909,N_7604,N_7667);
nor U7910 (N_7910,N_7685,N_7730);
and U7911 (N_7911,N_7733,N_7648);
nand U7912 (N_7912,N_7695,N_7715);
nand U7913 (N_7913,N_7695,N_7620);
and U7914 (N_7914,N_7601,N_7715);
or U7915 (N_7915,N_7679,N_7770);
nand U7916 (N_7916,N_7695,N_7691);
nand U7917 (N_7917,N_7675,N_7606);
and U7918 (N_7918,N_7643,N_7663);
or U7919 (N_7919,N_7617,N_7613);
nand U7920 (N_7920,N_7748,N_7664);
or U7921 (N_7921,N_7602,N_7779);
nor U7922 (N_7922,N_7715,N_7676);
nand U7923 (N_7923,N_7619,N_7729);
and U7924 (N_7924,N_7653,N_7683);
and U7925 (N_7925,N_7713,N_7620);
or U7926 (N_7926,N_7776,N_7649);
nand U7927 (N_7927,N_7610,N_7621);
nor U7928 (N_7928,N_7711,N_7772);
or U7929 (N_7929,N_7779,N_7721);
and U7930 (N_7930,N_7669,N_7679);
and U7931 (N_7931,N_7798,N_7635);
or U7932 (N_7932,N_7752,N_7715);
and U7933 (N_7933,N_7700,N_7747);
nand U7934 (N_7934,N_7645,N_7676);
nand U7935 (N_7935,N_7705,N_7658);
or U7936 (N_7936,N_7709,N_7790);
nand U7937 (N_7937,N_7755,N_7626);
and U7938 (N_7938,N_7772,N_7682);
or U7939 (N_7939,N_7633,N_7777);
nor U7940 (N_7940,N_7629,N_7650);
nor U7941 (N_7941,N_7742,N_7669);
nor U7942 (N_7942,N_7775,N_7703);
nand U7943 (N_7943,N_7746,N_7796);
or U7944 (N_7944,N_7689,N_7731);
and U7945 (N_7945,N_7748,N_7675);
nor U7946 (N_7946,N_7691,N_7701);
or U7947 (N_7947,N_7796,N_7663);
nor U7948 (N_7948,N_7667,N_7707);
and U7949 (N_7949,N_7604,N_7645);
nand U7950 (N_7950,N_7791,N_7785);
nor U7951 (N_7951,N_7757,N_7799);
nand U7952 (N_7952,N_7675,N_7714);
nor U7953 (N_7953,N_7759,N_7696);
and U7954 (N_7954,N_7651,N_7769);
nor U7955 (N_7955,N_7724,N_7749);
and U7956 (N_7956,N_7606,N_7734);
and U7957 (N_7957,N_7774,N_7673);
nand U7958 (N_7958,N_7697,N_7706);
or U7959 (N_7959,N_7771,N_7749);
and U7960 (N_7960,N_7765,N_7725);
nand U7961 (N_7961,N_7759,N_7649);
nand U7962 (N_7962,N_7636,N_7690);
nand U7963 (N_7963,N_7709,N_7614);
nor U7964 (N_7964,N_7656,N_7742);
nor U7965 (N_7965,N_7654,N_7707);
nand U7966 (N_7966,N_7684,N_7616);
or U7967 (N_7967,N_7768,N_7760);
nand U7968 (N_7968,N_7641,N_7761);
and U7969 (N_7969,N_7793,N_7673);
or U7970 (N_7970,N_7767,N_7742);
and U7971 (N_7971,N_7746,N_7679);
or U7972 (N_7972,N_7796,N_7737);
nor U7973 (N_7973,N_7719,N_7671);
or U7974 (N_7974,N_7744,N_7777);
nand U7975 (N_7975,N_7719,N_7789);
nor U7976 (N_7976,N_7706,N_7656);
or U7977 (N_7977,N_7716,N_7714);
or U7978 (N_7978,N_7772,N_7639);
and U7979 (N_7979,N_7724,N_7708);
nand U7980 (N_7980,N_7730,N_7628);
nor U7981 (N_7981,N_7702,N_7602);
or U7982 (N_7982,N_7631,N_7627);
or U7983 (N_7983,N_7715,N_7633);
nand U7984 (N_7984,N_7613,N_7748);
nand U7985 (N_7985,N_7729,N_7775);
nand U7986 (N_7986,N_7755,N_7634);
nand U7987 (N_7987,N_7673,N_7729);
or U7988 (N_7988,N_7612,N_7735);
nor U7989 (N_7989,N_7625,N_7747);
and U7990 (N_7990,N_7680,N_7774);
or U7991 (N_7991,N_7663,N_7735);
and U7992 (N_7992,N_7675,N_7645);
nor U7993 (N_7993,N_7725,N_7756);
xor U7994 (N_7994,N_7684,N_7621);
nor U7995 (N_7995,N_7768,N_7718);
and U7996 (N_7996,N_7776,N_7690);
nor U7997 (N_7997,N_7611,N_7648);
xor U7998 (N_7998,N_7642,N_7739);
and U7999 (N_7999,N_7747,N_7742);
and U8000 (N_8000,N_7982,N_7832);
and U8001 (N_8001,N_7936,N_7957);
nand U8002 (N_8002,N_7917,N_7921);
or U8003 (N_8003,N_7891,N_7986);
nand U8004 (N_8004,N_7985,N_7870);
nor U8005 (N_8005,N_7941,N_7900);
nand U8006 (N_8006,N_7833,N_7823);
and U8007 (N_8007,N_7830,N_7945);
nor U8008 (N_8008,N_7866,N_7812);
and U8009 (N_8009,N_7886,N_7913);
and U8010 (N_8010,N_7804,N_7839);
or U8011 (N_8011,N_7828,N_7869);
and U8012 (N_8012,N_7905,N_7808);
and U8013 (N_8013,N_7883,N_7931);
nor U8014 (N_8014,N_7923,N_7852);
or U8015 (N_8015,N_7879,N_7893);
nand U8016 (N_8016,N_7890,N_7959);
or U8017 (N_8017,N_7930,N_7916);
or U8018 (N_8018,N_7840,N_7861);
xnor U8019 (N_8019,N_7807,N_7826);
nand U8020 (N_8020,N_7805,N_7819);
or U8021 (N_8021,N_7860,N_7984);
nor U8022 (N_8022,N_7909,N_7868);
nand U8023 (N_8023,N_7952,N_7845);
nand U8024 (N_8024,N_7871,N_7859);
or U8025 (N_8025,N_7932,N_7961);
nand U8026 (N_8026,N_7971,N_7875);
or U8027 (N_8027,N_7838,N_7981);
or U8028 (N_8028,N_7882,N_7876);
nor U8029 (N_8029,N_7865,N_7946);
nand U8030 (N_8030,N_7806,N_7847);
nand U8031 (N_8031,N_7851,N_7873);
nand U8032 (N_8032,N_7885,N_7996);
or U8033 (N_8033,N_7944,N_7906);
xnor U8034 (N_8034,N_7953,N_7935);
or U8035 (N_8035,N_7822,N_7902);
and U8036 (N_8036,N_7979,N_7827);
and U8037 (N_8037,N_7801,N_7993);
nor U8038 (N_8038,N_7948,N_7815);
and U8039 (N_8039,N_7898,N_7825);
and U8040 (N_8040,N_7991,N_7872);
or U8041 (N_8041,N_7968,N_7999);
xor U8042 (N_8042,N_7889,N_7926);
and U8043 (N_8043,N_7943,N_7934);
nand U8044 (N_8044,N_7973,N_7818);
nand U8045 (N_8045,N_7835,N_7858);
and U8046 (N_8046,N_7951,N_7834);
or U8047 (N_8047,N_7849,N_7987);
and U8048 (N_8048,N_7842,N_7896);
or U8049 (N_8049,N_7848,N_7844);
nor U8050 (N_8050,N_7992,N_7978);
nor U8051 (N_8051,N_7908,N_7862);
nor U8052 (N_8052,N_7837,N_7942);
or U8053 (N_8053,N_7924,N_7950);
nor U8054 (N_8054,N_7910,N_7867);
nor U8055 (N_8055,N_7878,N_7892);
or U8056 (N_8056,N_7956,N_7937);
or U8057 (N_8057,N_7811,N_7966);
or U8058 (N_8058,N_7977,N_7997);
or U8059 (N_8059,N_7850,N_7960);
nand U8060 (N_8060,N_7824,N_7955);
nand U8061 (N_8061,N_7816,N_7853);
nand U8062 (N_8062,N_7964,N_7970);
and U8063 (N_8063,N_7962,N_7933);
and U8064 (N_8064,N_7928,N_7949);
and U8065 (N_8065,N_7820,N_7969);
or U8066 (N_8066,N_7920,N_7809);
or U8067 (N_8067,N_7903,N_7854);
nor U8068 (N_8068,N_7888,N_7915);
nor U8069 (N_8069,N_7958,N_7831);
or U8070 (N_8070,N_7884,N_7874);
or U8071 (N_8071,N_7919,N_7963);
nor U8072 (N_8072,N_7972,N_7803);
or U8073 (N_8073,N_7855,N_7975);
nand U8074 (N_8074,N_7990,N_7857);
nand U8075 (N_8075,N_7894,N_7904);
and U8076 (N_8076,N_7912,N_7800);
and U8077 (N_8077,N_7899,N_7974);
nand U8078 (N_8078,N_7856,N_7843);
nor U8079 (N_8079,N_7841,N_7817);
nor U8080 (N_8080,N_7954,N_7821);
and U8081 (N_8081,N_7939,N_7901);
or U8082 (N_8082,N_7877,N_7846);
nand U8083 (N_8083,N_7863,N_7813);
nand U8084 (N_8084,N_7995,N_7895);
and U8085 (N_8085,N_7967,N_7980);
nor U8086 (N_8086,N_7922,N_7918);
or U8087 (N_8087,N_7965,N_7914);
nand U8088 (N_8088,N_7814,N_7983);
nand U8089 (N_8089,N_7994,N_7897);
and U8090 (N_8090,N_7829,N_7810);
or U8091 (N_8091,N_7947,N_7911);
nand U8092 (N_8092,N_7998,N_7864);
nor U8093 (N_8093,N_7907,N_7881);
or U8094 (N_8094,N_7887,N_7836);
xor U8095 (N_8095,N_7988,N_7927);
and U8096 (N_8096,N_7880,N_7989);
nor U8097 (N_8097,N_7929,N_7976);
nand U8098 (N_8098,N_7940,N_7802);
nand U8099 (N_8099,N_7938,N_7925);
nor U8100 (N_8100,N_7976,N_7825);
nand U8101 (N_8101,N_7842,N_7963);
and U8102 (N_8102,N_7862,N_7954);
and U8103 (N_8103,N_7850,N_7911);
nor U8104 (N_8104,N_7934,N_7982);
or U8105 (N_8105,N_7900,N_7915);
nor U8106 (N_8106,N_7896,N_7997);
nor U8107 (N_8107,N_7857,N_7979);
nand U8108 (N_8108,N_7939,N_7979);
and U8109 (N_8109,N_7865,N_7892);
or U8110 (N_8110,N_7907,N_7960);
and U8111 (N_8111,N_7903,N_7984);
nand U8112 (N_8112,N_7894,N_7859);
and U8113 (N_8113,N_7844,N_7831);
nand U8114 (N_8114,N_7813,N_7875);
nor U8115 (N_8115,N_7962,N_7813);
xnor U8116 (N_8116,N_7874,N_7949);
nand U8117 (N_8117,N_7977,N_7988);
nand U8118 (N_8118,N_7963,N_7946);
nor U8119 (N_8119,N_7951,N_7909);
nand U8120 (N_8120,N_7983,N_7849);
nand U8121 (N_8121,N_7987,N_7829);
or U8122 (N_8122,N_7806,N_7966);
and U8123 (N_8123,N_7832,N_7898);
or U8124 (N_8124,N_7875,N_7916);
nand U8125 (N_8125,N_7946,N_7934);
nand U8126 (N_8126,N_7927,N_7916);
or U8127 (N_8127,N_7967,N_7973);
nor U8128 (N_8128,N_7938,N_7803);
and U8129 (N_8129,N_7843,N_7817);
nor U8130 (N_8130,N_7977,N_7825);
nand U8131 (N_8131,N_7817,N_7954);
nor U8132 (N_8132,N_7905,N_7833);
nand U8133 (N_8133,N_7926,N_7974);
nand U8134 (N_8134,N_7870,N_7980);
or U8135 (N_8135,N_7959,N_7822);
or U8136 (N_8136,N_7829,N_7943);
or U8137 (N_8137,N_7839,N_7817);
or U8138 (N_8138,N_7807,N_7855);
and U8139 (N_8139,N_7890,N_7871);
and U8140 (N_8140,N_7942,N_7818);
xor U8141 (N_8141,N_7933,N_7870);
and U8142 (N_8142,N_7836,N_7898);
nor U8143 (N_8143,N_7993,N_7850);
nor U8144 (N_8144,N_7814,N_7868);
or U8145 (N_8145,N_7814,N_7818);
nor U8146 (N_8146,N_7945,N_7910);
or U8147 (N_8147,N_7984,N_7826);
nor U8148 (N_8148,N_7930,N_7847);
and U8149 (N_8149,N_7810,N_7879);
and U8150 (N_8150,N_7944,N_7868);
and U8151 (N_8151,N_7820,N_7838);
nand U8152 (N_8152,N_7816,N_7995);
nand U8153 (N_8153,N_7900,N_7990);
and U8154 (N_8154,N_7992,N_7967);
nand U8155 (N_8155,N_7885,N_7881);
or U8156 (N_8156,N_7924,N_7942);
nand U8157 (N_8157,N_7998,N_7986);
nor U8158 (N_8158,N_7925,N_7806);
nor U8159 (N_8159,N_7934,N_7944);
nor U8160 (N_8160,N_7958,N_7803);
nand U8161 (N_8161,N_7849,N_7817);
nand U8162 (N_8162,N_7847,N_7987);
nor U8163 (N_8163,N_7826,N_7933);
nor U8164 (N_8164,N_7929,N_7907);
nor U8165 (N_8165,N_7969,N_7808);
nor U8166 (N_8166,N_7944,N_7822);
and U8167 (N_8167,N_7978,N_7803);
nand U8168 (N_8168,N_7964,N_7816);
or U8169 (N_8169,N_7881,N_7927);
nor U8170 (N_8170,N_7934,N_7910);
and U8171 (N_8171,N_7950,N_7807);
and U8172 (N_8172,N_7963,N_7838);
nor U8173 (N_8173,N_7892,N_7988);
and U8174 (N_8174,N_7929,N_7845);
nor U8175 (N_8175,N_7859,N_7885);
nand U8176 (N_8176,N_7819,N_7890);
or U8177 (N_8177,N_7998,N_7886);
nor U8178 (N_8178,N_7867,N_7889);
nand U8179 (N_8179,N_7832,N_7988);
nor U8180 (N_8180,N_7853,N_7889);
nor U8181 (N_8181,N_7866,N_7842);
and U8182 (N_8182,N_7938,N_7884);
nor U8183 (N_8183,N_7849,N_7925);
nor U8184 (N_8184,N_7896,N_7888);
nor U8185 (N_8185,N_7918,N_7974);
nor U8186 (N_8186,N_7837,N_7821);
and U8187 (N_8187,N_7907,N_7922);
and U8188 (N_8188,N_7901,N_7812);
xnor U8189 (N_8189,N_7813,N_7898);
nand U8190 (N_8190,N_7884,N_7809);
nor U8191 (N_8191,N_7862,N_7963);
or U8192 (N_8192,N_7837,N_7846);
nor U8193 (N_8193,N_7878,N_7977);
or U8194 (N_8194,N_7995,N_7820);
and U8195 (N_8195,N_7923,N_7975);
and U8196 (N_8196,N_7966,N_7977);
nor U8197 (N_8197,N_7952,N_7834);
or U8198 (N_8198,N_7851,N_7833);
or U8199 (N_8199,N_7870,N_7969);
nand U8200 (N_8200,N_8042,N_8072);
or U8201 (N_8201,N_8086,N_8045);
nand U8202 (N_8202,N_8061,N_8055);
xnor U8203 (N_8203,N_8067,N_8001);
or U8204 (N_8204,N_8174,N_8176);
nand U8205 (N_8205,N_8081,N_8126);
nor U8206 (N_8206,N_8106,N_8150);
nor U8207 (N_8207,N_8037,N_8164);
nor U8208 (N_8208,N_8108,N_8119);
or U8209 (N_8209,N_8073,N_8123);
nor U8210 (N_8210,N_8191,N_8057);
and U8211 (N_8211,N_8082,N_8140);
nor U8212 (N_8212,N_8133,N_8146);
or U8213 (N_8213,N_8098,N_8135);
nand U8214 (N_8214,N_8091,N_8104);
and U8215 (N_8215,N_8148,N_8010);
and U8216 (N_8216,N_8145,N_8169);
or U8217 (N_8217,N_8110,N_8136);
nand U8218 (N_8218,N_8161,N_8163);
or U8219 (N_8219,N_8012,N_8141);
nor U8220 (N_8220,N_8155,N_8075);
and U8221 (N_8221,N_8187,N_8197);
nand U8222 (N_8222,N_8180,N_8114);
or U8223 (N_8223,N_8181,N_8051);
and U8224 (N_8224,N_8017,N_8031);
and U8225 (N_8225,N_8142,N_8097);
or U8226 (N_8226,N_8194,N_8183);
and U8227 (N_8227,N_8027,N_8168);
nand U8228 (N_8228,N_8127,N_8166);
or U8229 (N_8229,N_8059,N_8118);
nor U8230 (N_8230,N_8100,N_8087);
and U8231 (N_8231,N_8002,N_8043);
nand U8232 (N_8232,N_8056,N_8151);
and U8233 (N_8233,N_8048,N_8144);
and U8234 (N_8234,N_8109,N_8038);
and U8235 (N_8235,N_8156,N_8034);
nor U8236 (N_8236,N_8049,N_8112);
nand U8237 (N_8237,N_8005,N_8193);
nand U8238 (N_8238,N_8186,N_8095);
nand U8239 (N_8239,N_8154,N_8153);
or U8240 (N_8240,N_8060,N_8089);
and U8241 (N_8241,N_8117,N_8063);
and U8242 (N_8242,N_8015,N_8068);
nand U8243 (N_8243,N_8147,N_8022);
and U8244 (N_8244,N_8129,N_8058);
nand U8245 (N_8245,N_8115,N_8111);
and U8246 (N_8246,N_8040,N_8029);
nor U8247 (N_8247,N_8101,N_8132);
nor U8248 (N_8248,N_8125,N_8152);
and U8249 (N_8249,N_8192,N_8007);
or U8250 (N_8250,N_8088,N_8116);
nor U8251 (N_8251,N_8134,N_8046);
nor U8252 (N_8252,N_8032,N_8196);
nor U8253 (N_8253,N_8096,N_8071);
nand U8254 (N_8254,N_8175,N_8178);
nand U8255 (N_8255,N_8138,N_8172);
and U8256 (N_8256,N_8139,N_8011);
nand U8257 (N_8257,N_8099,N_8177);
nor U8258 (N_8258,N_8198,N_8107);
and U8259 (N_8259,N_8021,N_8185);
nand U8260 (N_8260,N_8105,N_8028);
or U8261 (N_8261,N_8062,N_8189);
and U8262 (N_8262,N_8120,N_8137);
nor U8263 (N_8263,N_8170,N_8016);
and U8264 (N_8264,N_8094,N_8084);
nor U8265 (N_8265,N_8023,N_8065);
nand U8266 (N_8266,N_8128,N_8026);
and U8267 (N_8267,N_8074,N_8158);
nand U8268 (N_8268,N_8064,N_8009);
nor U8269 (N_8269,N_8020,N_8008);
nand U8270 (N_8270,N_8167,N_8013);
and U8271 (N_8271,N_8157,N_8173);
nand U8272 (N_8272,N_8069,N_8149);
or U8273 (N_8273,N_8122,N_8036);
and U8274 (N_8274,N_8171,N_8006);
nor U8275 (N_8275,N_8033,N_8184);
xor U8276 (N_8276,N_8000,N_8039);
nor U8277 (N_8277,N_8085,N_8083);
or U8278 (N_8278,N_8103,N_8090);
and U8279 (N_8279,N_8077,N_8143);
or U8280 (N_8280,N_8113,N_8030);
nor U8281 (N_8281,N_8092,N_8162);
nand U8282 (N_8282,N_8165,N_8003);
nand U8283 (N_8283,N_8054,N_8050);
nand U8284 (N_8284,N_8121,N_8130);
nor U8285 (N_8285,N_8052,N_8179);
nor U8286 (N_8286,N_8025,N_8190);
or U8287 (N_8287,N_8004,N_8182);
and U8288 (N_8288,N_8093,N_8188);
and U8289 (N_8289,N_8035,N_8076);
nor U8290 (N_8290,N_8024,N_8079);
nand U8291 (N_8291,N_8041,N_8070);
and U8292 (N_8292,N_8080,N_8018);
or U8293 (N_8293,N_8014,N_8199);
or U8294 (N_8294,N_8019,N_8044);
or U8295 (N_8295,N_8131,N_8047);
and U8296 (N_8296,N_8160,N_8102);
and U8297 (N_8297,N_8078,N_8124);
nor U8298 (N_8298,N_8195,N_8053);
and U8299 (N_8299,N_8159,N_8066);
nand U8300 (N_8300,N_8080,N_8126);
nand U8301 (N_8301,N_8149,N_8081);
or U8302 (N_8302,N_8017,N_8005);
nand U8303 (N_8303,N_8019,N_8090);
nand U8304 (N_8304,N_8199,N_8093);
and U8305 (N_8305,N_8081,N_8010);
or U8306 (N_8306,N_8069,N_8137);
nor U8307 (N_8307,N_8100,N_8021);
nor U8308 (N_8308,N_8031,N_8121);
nand U8309 (N_8309,N_8144,N_8011);
nor U8310 (N_8310,N_8140,N_8103);
or U8311 (N_8311,N_8115,N_8011);
and U8312 (N_8312,N_8063,N_8171);
or U8313 (N_8313,N_8151,N_8008);
nand U8314 (N_8314,N_8083,N_8116);
and U8315 (N_8315,N_8126,N_8177);
and U8316 (N_8316,N_8140,N_8132);
xnor U8317 (N_8317,N_8123,N_8173);
or U8318 (N_8318,N_8129,N_8156);
and U8319 (N_8319,N_8165,N_8020);
nand U8320 (N_8320,N_8017,N_8077);
nor U8321 (N_8321,N_8003,N_8063);
or U8322 (N_8322,N_8027,N_8169);
nand U8323 (N_8323,N_8035,N_8006);
nand U8324 (N_8324,N_8122,N_8139);
nor U8325 (N_8325,N_8197,N_8013);
nand U8326 (N_8326,N_8001,N_8093);
nand U8327 (N_8327,N_8040,N_8071);
nand U8328 (N_8328,N_8049,N_8010);
and U8329 (N_8329,N_8143,N_8188);
nor U8330 (N_8330,N_8016,N_8109);
or U8331 (N_8331,N_8118,N_8194);
nand U8332 (N_8332,N_8166,N_8101);
or U8333 (N_8333,N_8038,N_8074);
nand U8334 (N_8334,N_8038,N_8009);
nor U8335 (N_8335,N_8068,N_8101);
nand U8336 (N_8336,N_8198,N_8180);
nand U8337 (N_8337,N_8097,N_8021);
or U8338 (N_8338,N_8115,N_8133);
nand U8339 (N_8339,N_8026,N_8074);
and U8340 (N_8340,N_8159,N_8014);
nor U8341 (N_8341,N_8190,N_8148);
or U8342 (N_8342,N_8079,N_8066);
nor U8343 (N_8343,N_8108,N_8183);
or U8344 (N_8344,N_8033,N_8156);
and U8345 (N_8345,N_8105,N_8161);
nand U8346 (N_8346,N_8010,N_8168);
nor U8347 (N_8347,N_8172,N_8135);
nand U8348 (N_8348,N_8108,N_8003);
and U8349 (N_8349,N_8142,N_8013);
and U8350 (N_8350,N_8135,N_8068);
and U8351 (N_8351,N_8009,N_8162);
and U8352 (N_8352,N_8106,N_8183);
and U8353 (N_8353,N_8076,N_8113);
and U8354 (N_8354,N_8001,N_8119);
or U8355 (N_8355,N_8028,N_8068);
nand U8356 (N_8356,N_8082,N_8049);
and U8357 (N_8357,N_8119,N_8128);
nand U8358 (N_8358,N_8173,N_8041);
or U8359 (N_8359,N_8103,N_8198);
nand U8360 (N_8360,N_8077,N_8110);
nand U8361 (N_8361,N_8052,N_8043);
and U8362 (N_8362,N_8150,N_8077);
or U8363 (N_8363,N_8040,N_8137);
and U8364 (N_8364,N_8061,N_8072);
or U8365 (N_8365,N_8077,N_8158);
or U8366 (N_8366,N_8088,N_8141);
and U8367 (N_8367,N_8061,N_8150);
and U8368 (N_8368,N_8121,N_8015);
nor U8369 (N_8369,N_8003,N_8193);
and U8370 (N_8370,N_8129,N_8191);
and U8371 (N_8371,N_8176,N_8073);
and U8372 (N_8372,N_8063,N_8072);
or U8373 (N_8373,N_8043,N_8173);
or U8374 (N_8374,N_8199,N_8062);
nor U8375 (N_8375,N_8182,N_8032);
or U8376 (N_8376,N_8199,N_8139);
nand U8377 (N_8377,N_8024,N_8162);
nand U8378 (N_8378,N_8058,N_8000);
nor U8379 (N_8379,N_8047,N_8160);
or U8380 (N_8380,N_8130,N_8193);
and U8381 (N_8381,N_8114,N_8164);
nor U8382 (N_8382,N_8033,N_8198);
and U8383 (N_8383,N_8075,N_8132);
nand U8384 (N_8384,N_8164,N_8143);
nor U8385 (N_8385,N_8149,N_8021);
xor U8386 (N_8386,N_8117,N_8082);
nor U8387 (N_8387,N_8020,N_8194);
nand U8388 (N_8388,N_8004,N_8161);
nand U8389 (N_8389,N_8095,N_8096);
and U8390 (N_8390,N_8039,N_8100);
nor U8391 (N_8391,N_8140,N_8030);
nor U8392 (N_8392,N_8107,N_8148);
nand U8393 (N_8393,N_8036,N_8197);
nor U8394 (N_8394,N_8115,N_8083);
or U8395 (N_8395,N_8125,N_8181);
nand U8396 (N_8396,N_8074,N_8049);
nand U8397 (N_8397,N_8041,N_8108);
or U8398 (N_8398,N_8067,N_8080);
and U8399 (N_8399,N_8012,N_8004);
or U8400 (N_8400,N_8309,N_8355);
nand U8401 (N_8401,N_8229,N_8264);
nor U8402 (N_8402,N_8391,N_8226);
nor U8403 (N_8403,N_8313,N_8288);
or U8404 (N_8404,N_8270,N_8281);
and U8405 (N_8405,N_8344,N_8316);
nor U8406 (N_8406,N_8279,N_8219);
nand U8407 (N_8407,N_8342,N_8381);
or U8408 (N_8408,N_8374,N_8203);
and U8409 (N_8409,N_8283,N_8236);
nand U8410 (N_8410,N_8248,N_8246);
and U8411 (N_8411,N_8321,N_8209);
or U8412 (N_8412,N_8276,N_8349);
and U8413 (N_8413,N_8335,N_8261);
nand U8414 (N_8414,N_8322,N_8388);
and U8415 (N_8415,N_8385,N_8341);
or U8416 (N_8416,N_8319,N_8232);
nand U8417 (N_8417,N_8206,N_8234);
and U8418 (N_8418,N_8375,N_8367);
nor U8419 (N_8419,N_8253,N_8207);
nand U8420 (N_8420,N_8259,N_8320);
nor U8421 (N_8421,N_8312,N_8364);
nand U8422 (N_8422,N_8244,N_8386);
or U8423 (N_8423,N_8373,N_8363);
nor U8424 (N_8424,N_8208,N_8360);
and U8425 (N_8425,N_8269,N_8224);
nor U8426 (N_8426,N_8387,N_8358);
nand U8427 (N_8427,N_8324,N_8222);
or U8428 (N_8428,N_8353,N_8352);
nor U8429 (N_8429,N_8299,N_8250);
nor U8430 (N_8430,N_8325,N_8327);
or U8431 (N_8431,N_8204,N_8225);
nand U8432 (N_8432,N_8376,N_8392);
nor U8433 (N_8433,N_8223,N_8240);
or U8434 (N_8434,N_8368,N_8365);
nor U8435 (N_8435,N_8297,N_8267);
and U8436 (N_8436,N_8359,N_8336);
nor U8437 (N_8437,N_8295,N_8256);
or U8438 (N_8438,N_8286,N_8252);
nor U8439 (N_8439,N_8379,N_8380);
or U8440 (N_8440,N_8307,N_8356);
nand U8441 (N_8441,N_8318,N_8306);
nand U8442 (N_8442,N_8287,N_8315);
or U8443 (N_8443,N_8378,N_8289);
nand U8444 (N_8444,N_8370,N_8280);
or U8445 (N_8445,N_8348,N_8372);
nor U8446 (N_8446,N_8228,N_8333);
or U8447 (N_8447,N_8218,N_8255);
and U8448 (N_8448,N_8357,N_8243);
nand U8449 (N_8449,N_8214,N_8314);
nor U8450 (N_8450,N_8258,N_8210);
and U8451 (N_8451,N_8294,N_8266);
nor U8452 (N_8452,N_8260,N_8369);
or U8453 (N_8453,N_8371,N_8201);
and U8454 (N_8454,N_8346,N_8384);
nor U8455 (N_8455,N_8323,N_8254);
or U8456 (N_8456,N_8278,N_8302);
xor U8457 (N_8457,N_8310,N_8383);
nand U8458 (N_8458,N_8257,N_8247);
nand U8459 (N_8459,N_8397,N_8398);
nand U8460 (N_8460,N_8202,N_8275);
or U8461 (N_8461,N_8317,N_8227);
or U8462 (N_8462,N_8235,N_8361);
or U8463 (N_8463,N_8330,N_8331);
or U8464 (N_8464,N_8211,N_8268);
nand U8465 (N_8465,N_8262,N_8212);
nor U8466 (N_8466,N_8200,N_8389);
and U8467 (N_8467,N_8350,N_8311);
and U8468 (N_8468,N_8366,N_8274);
nor U8469 (N_8469,N_8277,N_8345);
or U8470 (N_8470,N_8242,N_8233);
and U8471 (N_8471,N_8220,N_8272);
nand U8472 (N_8472,N_8339,N_8354);
nand U8473 (N_8473,N_8290,N_8304);
and U8474 (N_8474,N_8305,N_8239);
or U8475 (N_8475,N_8251,N_8282);
nand U8476 (N_8476,N_8230,N_8326);
or U8477 (N_8477,N_8238,N_8394);
nand U8478 (N_8478,N_8340,N_8377);
and U8479 (N_8479,N_8245,N_8337);
nor U8480 (N_8480,N_8216,N_8241);
or U8481 (N_8481,N_8347,N_8298);
and U8482 (N_8482,N_8273,N_8271);
and U8483 (N_8483,N_8351,N_8231);
nor U8484 (N_8484,N_8328,N_8334);
nand U8485 (N_8485,N_8303,N_8329);
or U8486 (N_8486,N_8249,N_8265);
nor U8487 (N_8487,N_8395,N_8308);
nor U8488 (N_8488,N_8215,N_8390);
or U8489 (N_8489,N_8301,N_8285);
or U8490 (N_8490,N_8221,N_8217);
and U8491 (N_8491,N_8338,N_8332);
nand U8492 (N_8492,N_8382,N_8263);
or U8493 (N_8493,N_8296,N_8291);
or U8494 (N_8494,N_8292,N_8293);
nor U8495 (N_8495,N_8205,N_8300);
nand U8496 (N_8496,N_8393,N_8213);
or U8497 (N_8497,N_8284,N_8399);
nor U8498 (N_8498,N_8343,N_8237);
or U8499 (N_8499,N_8396,N_8362);
and U8500 (N_8500,N_8264,N_8393);
nand U8501 (N_8501,N_8229,N_8276);
or U8502 (N_8502,N_8252,N_8276);
nand U8503 (N_8503,N_8322,N_8295);
nand U8504 (N_8504,N_8368,N_8318);
nor U8505 (N_8505,N_8351,N_8302);
or U8506 (N_8506,N_8271,N_8361);
and U8507 (N_8507,N_8379,N_8276);
or U8508 (N_8508,N_8209,N_8203);
or U8509 (N_8509,N_8212,N_8264);
and U8510 (N_8510,N_8326,N_8283);
or U8511 (N_8511,N_8394,N_8371);
nor U8512 (N_8512,N_8226,N_8344);
nand U8513 (N_8513,N_8387,N_8254);
and U8514 (N_8514,N_8315,N_8394);
and U8515 (N_8515,N_8371,N_8209);
nand U8516 (N_8516,N_8243,N_8387);
and U8517 (N_8517,N_8394,N_8261);
nand U8518 (N_8518,N_8328,N_8274);
and U8519 (N_8519,N_8395,N_8337);
and U8520 (N_8520,N_8317,N_8210);
and U8521 (N_8521,N_8369,N_8343);
nand U8522 (N_8522,N_8317,N_8244);
nand U8523 (N_8523,N_8293,N_8357);
or U8524 (N_8524,N_8257,N_8330);
and U8525 (N_8525,N_8231,N_8246);
xor U8526 (N_8526,N_8220,N_8363);
or U8527 (N_8527,N_8353,N_8212);
nor U8528 (N_8528,N_8272,N_8346);
and U8529 (N_8529,N_8327,N_8354);
and U8530 (N_8530,N_8251,N_8384);
nand U8531 (N_8531,N_8284,N_8244);
and U8532 (N_8532,N_8218,N_8287);
nand U8533 (N_8533,N_8310,N_8329);
nor U8534 (N_8534,N_8269,N_8381);
or U8535 (N_8535,N_8325,N_8217);
or U8536 (N_8536,N_8210,N_8375);
and U8537 (N_8537,N_8323,N_8378);
or U8538 (N_8538,N_8314,N_8385);
nand U8539 (N_8539,N_8332,N_8352);
nand U8540 (N_8540,N_8372,N_8236);
nand U8541 (N_8541,N_8296,N_8248);
and U8542 (N_8542,N_8299,N_8290);
and U8543 (N_8543,N_8372,N_8365);
nand U8544 (N_8544,N_8377,N_8262);
nor U8545 (N_8545,N_8218,N_8361);
nand U8546 (N_8546,N_8272,N_8356);
nand U8547 (N_8547,N_8230,N_8261);
and U8548 (N_8548,N_8370,N_8305);
and U8549 (N_8549,N_8353,N_8310);
nand U8550 (N_8550,N_8256,N_8312);
nand U8551 (N_8551,N_8389,N_8364);
and U8552 (N_8552,N_8263,N_8215);
and U8553 (N_8553,N_8314,N_8288);
nor U8554 (N_8554,N_8315,N_8239);
nand U8555 (N_8555,N_8387,N_8218);
nand U8556 (N_8556,N_8386,N_8206);
nand U8557 (N_8557,N_8216,N_8261);
and U8558 (N_8558,N_8313,N_8342);
nand U8559 (N_8559,N_8233,N_8335);
nor U8560 (N_8560,N_8214,N_8230);
nand U8561 (N_8561,N_8285,N_8382);
nand U8562 (N_8562,N_8245,N_8385);
nor U8563 (N_8563,N_8208,N_8348);
nor U8564 (N_8564,N_8312,N_8252);
nor U8565 (N_8565,N_8333,N_8303);
nor U8566 (N_8566,N_8261,N_8315);
nor U8567 (N_8567,N_8272,N_8251);
nor U8568 (N_8568,N_8235,N_8212);
and U8569 (N_8569,N_8352,N_8363);
nand U8570 (N_8570,N_8276,N_8389);
and U8571 (N_8571,N_8336,N_8385);
nand U8572 (N_8572,N_8249,N_8370);
and U8573 (N_8573,N_8291,N_8219);
or U8574 (N_8574,N_8388,N_8221);
and U8575 (N_8575,N_8279,N_8375);
nor U8576 (N_8576,N_8208,N_8389);
nor U8577 (N_8577,N_8206,N_8280);
nor U8578 (N_8578,N_8356,N_8304);
nand U8579 (N_8579,N_8248,N_8317);
and U8580 (N_8580,N_8208,N_8362);
xnor U8581 (N_8581,N_8399,N_8349);
nor U8582 (N_8582,N_8377,N_8288);
nor U8583 (N_8583,N_8348,N_8259);
and U8584 (N_8584,N_8319,N_8376);
or U8585 (N_8585,N_8323,N_8387);
or U8586 (N_8586,N_8210,N_8236);
nand U8587 (N_8587,N_8356,N_8231);
nand U8588 (N_8588,N_8216,N_8286);
nor U8589 (N_8589,N_8213,N_8307);
or U8590 (N_8590,N_8398,N_8344);
nand U8591 (N_8591,N_8305,N_8300);
nor U8592 (N_8592,N_8238,N_8322);
nor U8593 (N_8593,N_8317,N_8392);
nor U8594 (N_8594,N_8278,N_8369);
nand U8595 (N_8595,N_8312,N_8286);
nor U8596 (N_8596,N_8371,N_8315);
and U8597 (N_8597,N_8315,N_8269);
nor U8598 (N_8598,N_8311,N_8316);
and U8599 (N_8599,N_8272,N_8237);
nor U8600 (N_8600,N_8400,N_8595);
and U8601 (N_8601,N_8577,N_8536);
or U8602 (N_8602,N_8598,N_8421);
or U8603 (N_8603,N_8593,N_8544);
or U8604 (N_8604,N_8546,N_8542);
and U8605 (N_8605,N_8427,N_8440);
nor U8606 (N_8606,N_8460,N_8465);
nand U8607 (N_8607,N_8489,N_8420);
or U8608 (N_8608,N_8446,N_8579);
or U8609 (N_8609,N_8584,N_8521);
nand U8610 (N_8610,N_8447,N_8423);
or U8611 (N_8611,N_8478,N_8456);
or U8612 (N_8612,N_8473,N_8592);
or U8613 (N_8613,N_8506,N_8588);
and U8614 (N_8614,N_8591,N_8484);
or U8615 (N_8615,N_8550,N_8408);
or U8616 (N_8616,N_8437,N_8475);
nand U8617 (N_8617,N_8479,N_8454);
nor U8618 (N_8618,N_8496,N_8486);
nor U8619 (N_8619,N_8438,N_8426);
or U8620 (N_8620,N_8540,N_8406);
and U8621 (N_8621,N_8562,N_8582);
nor U8622 (N_8622,N_8590,N_8512);
and U8623 (N_8623,N_8573,N_8411);
or U8624 (N_8624,N_8409,N_8463);
nor U8625 (N_8625,N_8466,N_8439);
nor U8626 (N_8626,N_8572,N_8509);
nand U8627 (N_8627,N_8514,N_8574);
nand U8628 (N_8628,N_8494,N_8442);
or U8629 (N_8629,N_8445,N_8545);
nand U8630 (N_8630,N_8414,N_8425);
and U8631 (N_8631,N_8461,N_8551);
nor U8632 (N_8632,N_8534,N_8441);
and U8633 (N_8633,N_8524,N_8527);
or U8634 (N_8634,N_8531,N_8568);
or U8635 (N_8635,N_8499,N_8468);
and U8636 (N_8636,N_8529,N_8552);
or U8637 (N_8637,N_8462,N_8515);
nand U8638 (N_8638,N_8508,N_8500);
and U8639 (N_8639,N_8491,N_8434);
and U8640 (N_8640,N_8516,N_8513);
or U8641 (N_8641,N_8424,N_8578);
nor U8642 (N_8642,N_8498,N_8548);
nand U8643 (N_8643,N_8549,N_8449);
nor U8644 (N_8644,N_8430,N_8415);
or U8645 (N_8645,N_8448,N_8416);
nor U8646 (N_8646,N_8556,N_8472);
nor U8647 (N_8647,N_8526,N_8530);
nor U8648 (N_8648,N_8528,N_8537);
or U8649 (N_8649,N_8453,N_8410);
nor U8650 (N_8650,N_8589,N_8597);
nand U8651 (N_8651,N_8443,N_8429);
and U8652 (N_8652,N_8532,N_8518);
or U8653 (N_8653,N_8422,N_8431);
or U8654 (N_8654,N_8560,N_8523);
and U8655 (N_8655,N_8407,N_8404);
or U8656 (N_8656,N_8554,N_8569);
nand U8657 (N_8657,N_8464,N_8567);
and U8658 (N_8658,N_8547,N_8482);
nand U8659 (N_8659,N_8561,N_8511);
nor U8660 (N_8660,N_8580,N_8522);
nor U8661 (N_8661,N_8559,N_8481);
nor U8662 (N_8662,N_8488,N_8510);
or U8663 (N_8663,N_8570,N_8503);
nand U8664 (N_8664,N_8576,N_8432);
nand U8665 (N_8665,N_8507,N_8519);
nor U8666 (N_8666,N_8470,N_8413);
nand U8667 (N_8667,N_8555,N_8557);
or U8668 (N_8668,N_8586,N_8435);
or U8669 (N_8669,N_8596,N_8585);
nand U8670 (N_8670,N_8452,N_8467);
and U8671 (N_8671,N_8517,N_8520);
nand U8672 (N_8672,N_8539,N_8455);
nand U8673 (N_8673,N_8495,N_8474);
or U8674 (N_8674,N_8571,N_8497);
and U8675 (N_8675,N_8459,N_8418);
nor U8676 (N_8676,N_8403,N_8505);
and U8677 (N_8677,N_8587,N_8402);
and U8678 (N_8678,N_8405,N_8525);
nand U8679 (N_8679,N_8487,N_8594);
or U8680 (N_8680,N_8492,N_8476);
and U8681 (N_8681,N_8533,N_8504);
or U8682 (N_8682,N_8541,N_8599);
or U8683 (N_8683,N_8419,N_8564);
nand U8684 (N_8684,N_8583,N_8469);
nor U8685 (N_8685,N_8433,N_8483);
nand U8686 (N_8686,N_8566,N_8581);
and U8687 (N_8687,N_8401,N_8480);
or U8688 (N_8688,N_8501,N_8451);
or U8689 (N_8689,N_8417,N_8565);
and U8690 (N_8690,N_8428,N_8436);
nor U8691 (N_8691,N_8412,N_8471);
and U8692 (N_8692,N_8493,N_8575);
nor U8693 (N_8693,N_8457,N_8558);
nand U8694 (N_8694,N_8477,N_8543);
nor U8695 (N_8695,N_8538,N_8450);
or U8696 (N_8696,N_8490,N_8563);
nand U8697 (N_8697,N_8502,N_8458);
nand U8698 (N_8698,N_8444,N_8485);
nand U8699 (N_8699,N_8553,N_8535);
nand U8700 (N_8700,N_8470,N_8560);
or U8701 (N_8701,N_8514,N_8598);
nor U8702 (N_8702,N_8533,N_8581);
and U8703 (N_8703,N_8408,N_8527);
nand U8704 (N_8704,N_8407,N_8495);
and U8705 (N_8705,N_8406,N_8413);
or U8706 (N_8706,N_8533,N_8526);
nor U8707 (N_8707,N_8503,N_8484);
or U8708 (N_8708,N_8481,N_8418);
nor U8709 (N_8709,N_8567,N_8544);
nand U8710 (N_8710,N_8510,N_8509);
nor U8711 (N_8711,N_8560,N_8595);
nand U8712 (N_8712,N_8546,N_8504);
nor U8713 (N_8713,N_8515,N_8593);
or U8714 (N_8714,N_8464,N_8547);
or U8715 (N_8715,N_8532,N_8588);
nor U8716 (N_8716,N_8432,N_8520);
and U8717 (N_8717,N_8599,N_8435);
nor U8718 (N_8718,N_8501,N_8584);
or U8719 (N_8719,N_8467,N_8492);
or U8720 (N_8720,N_8577,N_8422);
nor U8721 (N_8721,N_8571,N_8481);
nor U8722 (N_8722,N_8467,N_8445);
nand U8723 (N_8723,N_8443,N_8486);
or U8724 (N_8724,N_8538,N_8454);
or U8725 (N_8725,N_8469,N_8464);
nand U8726 (N_8726,N_8517,N_8532);
nand U8727 (N_8727,N_8423,N_8503);
nand U8728 (N_8728,N_8536,N_8525);
nand U8729 (N_8729,N_8509,N_8419);
nand U8730 (N_8730,N_8583,N_8501);
and U8731 (N_8731,N_8410,N_8406);
or U8732 (N_8732,N_8449,N_8424);
or U8733 (N_8733,N_8523,N_8522);
or U8734 (N_8734,N_8556,N_8420);
xor U8735 (N_8735,N_8480,N_8591);
or U8736 (N_8736,N_8526,N_8451);
or U8737 (N_8737,N_8533,N_8572);
nor U8738 (N_8738,N_8441,N_8424);
nand U8739 (N_8739,N_8542,N_8464);
nor U8740 (N_8740,N_8460,N_8568);
nand U8741 (N_8741,N_8453,N_8429);
and U8742 (N_8742,N_8421,N_8492);
and U8743 (N_8743,N_8416,N_8431);
nor U8744 (N_8744,N_8480,N_8529);
and U8745 (N_8745,N_8491,N_8419);
nor U8746 (N_8746,N_8491,N_8497);
nand U8747 (N_8747,N_8484,N_8470);
and U8748 (N_8748,N_8560,N_8518);
or U8749 (N_8749,N_8490,N_8553);
nand U8750 (N_8750,N_8462,N_8445);
nand U8751 (N_8751,N_8438,N_8419);
and U8752 (N_8752,N_8484,N_8539);
nor U8753 (N_8753,N_8451,N_8521);
and U8754 (N_8754,N_8478,N_8457);
and U8755 (N_8755,N_8500,N_8411);
xnor U8756 (N_8756,N_8453,N_8422);
and U8757 (N_8757,N_8409,N_8527);
or U8758 (N_8758,N_8532,N_8453);
or U8759 (N_8759,N_8405,N_8404);
and U8760 (N_8760,N_8489,N_8582);
nor U8761 (N_8761,N_8548,N_8506);
or U8762 (N_8762,N_8544,N_8547);
nor U8763 (N_8763,N_8465,N_8488);
and U8764 (N_8764,N_8465,N_8406);
or U8765 (N_8765,N_8442,N_8439);
or U8766 (N_8766,N_8407,N_8429);
or U8767 (N_8767,N_8586,N_8564);
or U8768 (N_8768,N_8571,N_8536);
and U8769 (N_8769,N_8449,N_8586);
and U8770 (N_8770,N_8513,N_8464);
nand U8771 (N_8771,N_8435,N_8534);
and U8772 (N_8772,N_8534,N_8492);
or U8773 (N_8773,N_8599,N_8434);
and U8774 (N_8774,N_8440,N_8477);
and U8775 (N_8775,N_8590,N_8530);
and U8776 (N_8776,N_8479,N_8441);
nor U8777 (N_8777,N_8575,N_8474);
or U8778 (N_8778,N_8445,N_8423);
or U8779 (N_8779,N_8532,N_8560);
or U8780 (N_8780,N_8502,N_8529);
and U8781 (N_8781,N_8477,N_8562);
nand U8782 (N_8782,N_8466,N_8475);
or U8783 (N_8783,N_8500,N_8468);
and U8784 (N_8784,N_8551,N_8411);
and U8785 (N_8785,N_8487,N_8514);
and U8786 (N_8786,N_8435,N_8523);
or U8787 (N_8787,N_8414,N_8572);
or U8788 (N_8788,N_8549,N_8596);
and U8789 (N_8789,N_8529,N_8595);
nand U8790 (N_8790,N_8401,N_8523);
nand U8791 (N_8791,N_8570,N_8512);
or U8792 (N_8792,N_8590,N_8500);
and U8793 (N_8793,N_8555,N_8400);
and U8794 (N_8794,N_8467,N_8474);
nor U8795 (N_8795,N_8405,N_8521);
nand U8796 (N_8796,N_8550,N_8543);
and U8797 (N_8797,N_8455,N_8573);
or U8798 (N_8798,N_8441,N_8519);
nand U8799 (N_8799,N_8539,N_8532);
or U8800 (N_8800,N_8709,N_8644);
nor U8801 (N_8801,N_8681,N_8765);
nor U8802 (N_8802,N_8747,N_8686);
nor U8803 (N_8803,N_8653,N_8612);
nor U8804 (N_8804,N_8734,N_8691);
or U8805 (N_8805,N_8677,N_8659);
and U8806 (N_8806,N_8760,N_8702);
nor U8807 (N_8807,N_8725,N_8637);
or U8808 (N_8808,N_8689,N_8754);
nor U8809 (N_8809,N_8678,N_8640);
nor U8810 (N_8810,N_8753,N_8737);
nor U8811 (N_8811,N_8776,N_8665);
nor U8812 (N_8812,N_8626,N_8791);
nand U8813 (N_8813,N_8668,N_8704);
nor U8814 (N_8814,N_8770,N_8625);
or U8815 (N_8815,N_8690,N_8620);
nor U8816 (N_8816,N_8797,N_8636);
nor U8817 (N_8817,N_8731,N_8706);
or U8818 (N_8818,N_8750,N_8696);
nand U8819 (N_8819,N_8680,N_8749);
nand U8820 (N_8820,N_8628,N_8738);
nand U8821 (N_8821,N_8735,N_8710);
nand U8822 (N_8822,N_8707,N_8671);
and U8823 (N_8823,N_8605,N_8661);
or U8824 (N_8824,N_8601,N_8660);
nor U8825 (N_8825,N_8729,N_8715);
nor U8826 (N_8826,N_8792,N_8795);
nand U8827 (N_8827,N_8751,N_8767);
and U8828 (N_8828,N_8774,N_8647);
nand U8829 (N_8829,N_8787,N_8627);
and U8830 (N_8830,N_8739,N_8728);
nand U8831 (N_8831,N_8693,N_8727);
and U8832 (N_8832,N_8632,N_8759);
or U8833 (N_8833,N_8676,N_8799);
and U8834 (N_8834,N_8736,N_8633);
nand U8835 (N_8835,N_8764,N_8788);
and U8836 (N_8836,N_8651,N_8744);
xnor U8837 (N_8837,N_8624,N_8786);
and U8838 (N_8838,N_8723,N_8679);
and U8839 (N_8839,N_8635,N_8666);
and U8840 (N_8840,N_8656,N_8746);
nor U8841 (N_8841,N_8748,N_8609);
or U8842 (N_8842,N_8782,N_8768);
nor U8843 (N_8843,N_8726,N_8649);
or U8844 (N_8844,N_8694,N_8667);
and U8845 (N_8845,N_8663,N_8712);
and U8846 (N_8846,N_8745,N_8621);
nor U8847 (N_8847,N_8670,N_8692);
or U8848 (N_8848,N_8714,N_8718);
or U8849 (N_8849,N_8793,N_8648);
nor U8850 (N_8850,N_8672,N_8711);
and U8851 (N_8851,N_8716,N_8783);
nor U8852 (N_8852,N_8699,N_8766);
and U8853 (N_8853,N_8600,N_8683);
and U8854 (N_8854,N_8616,N_8602);
nand U8855 (N_8855,N_8763,N_8769);
and U8856 (N_8856,N_8733,N_8789);
or U8857 (N_8857,N_8752,N_8743);
or U8858 (N_8858,N_8794,N_8761);
and U8859 (N_8859,N_8701,N_8675);
nor U8860 (N_8860,N_8720,N_8664);
and U8861 (N_8861,N_8777,N_8781);
nand U8862 (N_8862,N_8604,N_8708);
nand U8863 (N_8863,N_8703,N_8643);
nand U8864 (N_8864,N_8742,N_8619);
and U8865 (N_8865,N_8611,N_8730);
nor U8866 (N_8866,N_8790,N_8682);
and U8867 (N_8867,N_8719,N_8614);
nor U8868 (N_8868,N_8608,N_8740);
and U8869 (N_8869,N_8772,N_8606);
nor U8870 (N_8870,N_8629,N_8631);
nor U8871 (N_8871,N_8658,N_8654);
and U8872 (N_8872,N_8673,N_8721);
nand U8873 (N_8873,N_8652,N_8655);
or U8874 (N_8874,N_8757,N_8758);
nor U8875 (N_8875,N_8779,N_8617);
or U8876 (N_8876,N_8775,N_8695);
and U8877 (N_8877,N_8642,N_8646);
and U8878 (N_8878,N_8756,N_8634);
and U8879 (N_8879,N_8773,N_8717);
nor U8880 (N_8880,N_8639,N_8771);
or U8881 (N_8881,N_8798,N_8630);
nand U8882 (N_8882,N_8623,N_8796);
xor U8883 (N_8883,N_8784,N_8662);
nor U8884 (N_8884,N_8778,N_8724);
and U8885 (N_8885,N_8684,N_8615);
or U8886 (N_8886,N_8618,N_8650);
nand U8887 (N_8887,N_8674,N_8645);
or U8888 (N_8888,N_8780,N_8613);
nand U8889 (N_8889,N_8638,N_8697);
and U8890 (N_8890,N_8603,N_8741);
and U8891 (N_8891,N_8669,N_8785);
and U8892 (N_8892,N_8755,N_8610);
nor U8893 (N_8893,N_8641,N_8698);
nand U8894 (N_8894,N_8688,N_8687);
or U8895 (N_8895,N_8622,N_8713);
and U8896 (N_8896,N_8685,N_8722);
and U8897 (N_8897,N_8732,N_8762);
nand U8898 (N_8898,N_8700,N_8657);
and U8899 (N_8899,N_8705,N_8607);
nand U8900 (N_8900,N_8692,N_8792);
nand U8901 (N_8901,N_8783,N_8726);
xnor U8902 (N_8902,N_8764,N_8676);
or U8903 (N_8903,N_8716,N_8613);
nor U8904 (N_8904,N_8703,N_8721);
and U8905 (N_8905,N_8653,N_8731);
and U8906 (N_8906,N_8617,N_8791);
and U8907 (N_8907,N_8644,N_8710);
nand U8908 (N_8908,N_8764,N_8677);
or U8909 (N_8909,N_8624,N_8749);
and U8910 (N_8910,N_8776,N_8682);
or U8911 (N_8911,N_8679,N_8668);
nand U8912 (N_8912,N_8752,N_8728);
nor U8913 (N_8913,N_8711,N_8706);
nand U8914 (N_8914,N_8739,N_8611);
nor U8915 (N_8915,N_8748,N_8794);
and U8916 (N_8916,N_8753,N_8671);
or U8917 (N_8917,N_8653,N_8683);
or U8918 (N_8918,N_8691,N_8669);
and U8919 (N_8919,N_8648,N_8654);
nor U8920 (N_8920,N_8700,N_8611);
nor U8921 (N_8921,N_8619,N_8719);
and U8922 (N_8922,N_8763,N_8626);
nand U8923 (N_8923,N_8616,N_8703);
or U8924 (N_8924,N_8755,N_8620);
nor U8925 (N_8925,N_8688,N_8609);
nand U8926 (N_8926,N_8632,N_8623);
and U8927 (N_8927,N_8729,N_8782);
nor U8928 (N_8928,N_8624,N_8766);
and U8929 (N_8929,N_8654,N_8719);
and U8930 (N_8930,N_8746,N_8655);
nor U8931 (N_8931,N_8745,N_8768);
nand U8932 (N_8932,N_8711,N_8628);
and U8933 (N_8933,N_8764,N_8678);
and U8934 (N_8934,N_8689,N_8720);
and U8935 (N_8935,N_8710,N_8754);
and U8936 (N_8936,N_8664,N_8638);
or U8937 (N_8937,N_8766,N_8622);
nand U8938 (N_8938,N_8749,N_8620);
or U8939 (N_8939,N_8797,N_8790);
or U8940 (N_8940,N_8642,N_8622);
nor U8941 (N_8941,N_8797,N_8696);
or U8942 (N_8942,N_8741,N_8619);
or U8943 (N_8943,N_8685,N_8652);
nor U8944 (N_8944,N_8727,N_8630);
nor U8945 (N_8945,N_8652,N_8670);
nor U8946 (N_8946,N_8713,N_8685);
nor U8947 (N_8947,N_8788,N_8701);
and U8948 (N_8948,N_8787,N_8676);
or U8949 (N_8949,N_8728,N_8673);
nand U8950 (N_8950,N_8787,N_8777);
and U8951 (N_8951,N_8650,N_8674);
or U8952 (N_8952,N_8671,N_8770);
nor U8953 (N_8953,N_8613,N_8773);
nand U8954 (N_8954,N_8733,N_8683);
and U8955 (N_8955,N_8625,N_8709);
or U8956 (N_8956,N_8657,N_8631);
and U8957 (N_8957,N_8615,N_8781);
and U8958 (N_8958,N_8724,N_8633);
nor U8959 (N_8959,N_8776,N_8610);
nand U8960 (N_8960,N_8616,N_8627);
nand U8961 (N_8961,N_8614,N_8771);
nor U8962 (N_8962,N_8733,N_8703);
xor U8963 (N_8963,N_8742,N_8797);
or U8964 (N_8964,N_8752,N_8651);
nand U8965 (N_8965,N_8712,N_8719);
and U8966 (N_8966,N_8686,N_8652);
and U8967 (N_8967,N_8710,N_8635);
nand U8968 (N_8968,N_8614,N_8605);
and U8969 (N_8969,N_8666,N_8671);
and U8970 (N_8970,N_8762,N_8679);
nand U8971 (N_8971,N_8762,N_8729);
or U8972 (N_8972,N_8631,N_8701);
nor U8973 (N_8973,N_8650,N_8692);
nor U8974 (N_8974,N_8668,N_8744);
or U8975 (N_8975,N_8672,N_8690);
nor U8976 (N_8976,N_8797,N_8746);
nand U8977 (N_8977,N_8744,N_8672);
nand U8978 (N_8978,N_8749,N_8618);
nand U8979 (N_8979,N_8716,N_8768);
or U8980 (N_8980,N_8663,N_8693);
nor U8981 (N_8981,N_8651,N_8624);
nand U8982 (N_8982,N_8681,N_8705);
nand U8983 (N_8983,N_8772,N_8750);
or U8984 (N_8984,N_8782,N_8674);
and U8985 (N_8985,N_8709,N_8736);
nand U8986 (N_8986,N_8658,N_8701);
nand U8987 (N_8987,N_8607,N_8708);
and U8988 (N_8988,N_8616,N_8772);
or U8989 (N_8989,N_8602,N_8658);
nand U8990 (N_8990,N_8780,N_8603);
or U8991 (N_8991,N_8650,N_8655);
or U8992 (N_8992,N_8683,N_8798);
or U8993 (N_8993,N_8676,N_8601);
nand U8994 (N_8994,N_8789,N_8709);
or U8995 (N_8995,N_8739,N_8755);
nand U8996 (N_8996,N_8770,N_8786);
nor U8997 (N_8997,N_8600,N_8707);
nand U8998 (N_8998,N_8709,N_8730);
nor U8999 (N_8999,N_8654,N_8717);
nand U9000 (N_9000,N_8823,N_8946);
nor U9001 (N_9001,N_8886,N_8935);
nor U9002 (N_9002,N_8862,N_8852);
nor U9003 (N_9003,N_8909,N_8937);
nand U9004 (N_9004,N_8825,N_8982);
or U9005 (N_9005,N_8840,N_8861);
nor U9006 (N_9006,N_8865,N_8815);
or U9007 (N_9007,N_8959,N_8822);
nor U9008 (N_9008,N_8806,N_8858);
or U9009 (N_9009,N_8938,N_8870);
or U9010 (N_9010,N_8936,N_8878);
and U9011 (N_9011,N_8873,N_8820);
nand U9012 (N_9012,N_8836,N_8996);
or U9013 (N_9013,N_8955,N_8966);
nand U9014 (N_9014,N_8802,N_8818);
or U9015 (N_9015,N_8869,N_8835);
nand U9016 (N_9016,N_8892,N_8979);
and U9017 (N_9017,N_8898,N_8880);
and U9018 (N_9018,N_8863,N_8964);
nor U9019 (N_9019,N_8953,N_8987);
or U9020 (N_9020,N_8977,N_8881);
or U9021 (N_9021,N_8947,N_8970);
and U9022 (N_9022,N_8847,N_8916);
nor U9023 (N_9023,N_8969,N_8997);
or U9024 (N_9024,N_8976,N_8853);
nand U9025 (N_9025,N_8911,N_8854);
nand U9026 (N_9026,N_8828,N_8926);
or U9027 (N_9027,N_8950,N_8952);
and U9028 (N_9028,N_8986,N_8967);
or U9029 (N_9029,N_8837,N_8894);
nand U9030 (N_9030,N_8891,N_8963);
nand U9031 (N_9031,N_8857,N_8920);
nand U9032 (N_9032,N_8887,N_8958);
nor U9033 (N_9033,N_8921,N_8819);
or U9034 (N_9034,N_8949,N_8848);
nor U9035 (N_9035,N_8992,N_8877);
or U9036 (N_9036,N_8808,N_8838);
nor U9037 (N_9037,N_8991,N_8804);
and U9038 (N_9038,N_8839,N_8951);
or U9039 (N_9039,N_8994,N_8905);
and U9040 (N_9040,N_8812,N_8895);
nor U9041 (N_9041,N_8919,N_8929);
nand U9042 (N_9042,N_8914,N_8980);
or U9043 (N_9043,N_8875,N_8957);
nand U9044 (N_9044,N_8830,N_8805);
nand U9045 (N_9045,N_8908,N_8864);
nor U9046 (N_9046,N_8826,N_8810);
nand U9047 (N_9047,N_8912,N_8884);
or U9048 (N_9048,N_8910,N_8934);
nand U9049 (N_9049,N_8915,N_8829);
nand U9050 (N_9050,N_8813,N_8859);
and U9051 (N_9051,N_8849,N_8893);
nor U9052 (N_9052,N_8917,N_8948);
or U9053 (N_9053,N_8883,N_8931);
or U9054 (N_9054,N_8956,N_8999);
or U9055 (N_9055,N_8906,N_8845);
nor U9056 (N_9056,N_8960,N_8855);
nand U9057 (N_9057,N_8834,N_8885);
nor U9058 (N_9058,N_8843,N_8942);
and U9059 (N_9059,N_8868,N_8896);
and U9060 (N_9060,N_8965,N_8872);
nand U9061 (N_9061,N_8962,N_8882);
nor U9062 (N_9062,N_8814,N_8945);
and U9063 (N_9063,N_8890,N_8972);
and U9064 (N_9064,N_8803,N_8832);
or U9065 (N_9065,N_8831,N_8807);
and U9066 (N_9066,N_8833,N_8867);
nand U9067 (N_9067,N_8827,N_8924);
and U9068 (N_9068,N_8866,N_8801);
nand U9069 (N_9069,N_8809,N_8922);
xor U9070 (N_9070,N_8816,N_8876);
or U9071 (N_9071,N_8940,N_8904);
or U9072 (N_9072,N_8817,N_8998);
nand U9073 (N_9073,N_8933,N_8971);
and U9074 (N_9074,N_8974,N_8901);
or U9075 (N_9075,N_8811,N_8918);
nand U9076 (N_9076,N_8984,N_8850);
or U9077 (N_9077,N_8871,N_8897);
nor U9078 (N_9078,N_8932,N_8989);
and U9079 (N_9079,N_8939,N_8928);
and U9080 (N_9080,N_8930,N_8923);
nand U9081 (N_9081,N_8841,N_8824);
nor U9082 (N_9082,N_8889,N_8978);
or U9083 (N_9083,N_8903,N_8851);
nand U9084 (N_9084,N_8925,N_8913);
nand U9085 (N_9085,N_8988,N_8860);
or U9086 (N_9086,N_8995,N_8900);
and U9087 (N_9087,N_8821,N_8842);
nor U9088 (N_9088,N_8944,N_8993);
nand U9089 (N_9089,N_8990,N_8800);
nand U9090 (N_9090,N_8899,N_8985);
nand U9091 (N_9091,N_8941,N_8961);
and U9092 (N_9092,N_8844,N_8981);
nor U9093 (N_9093,N_8927,N_8846);
nor U9094 (N_9094,N_8975,N_8954);
nor U9095 (N_9095,N_8973,N_8907);
nor U9096 (N_9096,N_8943,N_8856);
or U9097 (N_9097,N_8874,N_8879);
nand U9098 (N_9098,N_8983,N_8902);
nand U9099 (N_9099,N_8888,N_8968);
nor U9100 (N_9100,N_8972,N_8968);
nand U9101 (N_9101,N_8906,N_8853);
nand U9102 (N_9102,N_8817,N_8851);
nand U9103 (N_9103,N_8889,N_8832);
nand U9104 (N_9104,N_8980,N_8966);
and U9105 (N_9105,N_8895,N_8931);
nand U9106 (N_9106,N_8892,N_8835);
nand U9107 (N_9107,N_8838,N_8821);
or U9108 (N_9108,N_8827,N_8940);
nor U9109 (N_9109,N_8852,N_8945);
nand U9110 (N_9110,N_8912,N_8825);
nor U9111 (N_9111,N_8887,N_8860);
and U9112 (N_9112,N_8936,N_8985);
or U9113 (N_9113,N_8872,N_8828);
nand U9114 (N_9114,N_8881,N_8821);
and U9115 (N_9115,N_8900,N_8901);
and U9116 (N_9116,N_8818,N_8842);
and U9117 (N_9117,N_8843,N_8826);
or U9118 (N_9118,N_8811,N_8844);
nor U9119 (N_9119,N_8877,N_8876);
nand U9120 (N_9120,N_8827,N_8808);
nand U9121 (N_9121,N_8830,N_8867);
or U9122 (N_9122,N_8847,N_8851);
nor U9123 (N_9123,N_8899,N_8996);
and U9124 (N_9124,N_8964,N_8982);
nor U9125 (N_9125,N_8979,N_8967);
nand U9126 (N_9126,N_8984,N_8818);
or U9127 (N_9127,N_8991,N_8829);
xnor U9128 (N_9128,N_8832,N_8883);
nand U9129 (N_9129,N_8863,N_8937);
and U9130 (N_9130,N_8993,N_8804);
and U9131 (N_9131,N_8904,N_8898);
nor U9132 (N_9132,N_8820,N_8979);
nor U9133 (N_9133,N_8931,N_8891);
and U9134 (N_9134,N_8924,N_8991);
or U9135 (N_9135,N_8844,N_8907);
and U9136 (N_9136,N_8965,N_8909);
and U9137 (N_9137,N_8896,N_8840);
nand U9138 (N_9138,N_8872,N_8928);
nor U9139 (N_9139,N_8995,N_8888);
nand U9140 (N_9140,N_8991,N_8987);
and U9141 (N_9141,N_8835,N_8933);
nand U9142 (N_9142,N_8891,N_8897);
and U9143 (N_9143,N_8897,N_8853);
nor U9144 (N_9144,N_8905,N_8847);
or U9145 (N_9145,N_8821,N_8986);
and U9146 (N_9146,N_8844,N_8975);
or U9147 (N_9147,N_8887,N_8975);
nor U9148 (N_9148,N_8809,N_8891);
and U9149 (N_9149,N_8822,N_8863);
nor U9150 (N_9150,N_8879,N_8901);
and U9151 (N_9151,N_8917,N_8820);
nor U9152 (N_9152,N_8852,N_8941);
nor U9153 (N_9153,N_8816,N_8889);
nand U9154 (N_9154,N_8950,N_8991);
and U9155 (N_9155,N_8835,N_8919);
nand U9156 (N_9156,N_8824,N_8977);
nor U9157 (N_9157,N_8887,N_8968);
and U9158 (N_9158,N_8978,N_8885);
and U9159 (N_9159,N_8821,N_8925);
nor U9160 (N_9160,N_8938,N_8842);
or U9161 (N_9161,N_8875,N_8892);
or U9162 (N_9162,N_8873,N_8901);
and U9163 (N_9163,N_8839,N_8939);
nand U9164 (N_9164,N_8952,N_8818);
nor U9165 (N_9165,N_8907,N_8824);
or U9166 (N_9166,N_8895,N_8941);
and U9167 (N_9167,N_8972,N_8832);
or U9168 (N_9168,N_8823,N_8833);
or U9169 (N_9169,N_8883,N_8878);
nand U9170 (N_9170,N_8962,N_8958);
nor U9171 (N_9171,N_8835,N_8844);
and U9172 (N_9172,N_8881,N_8844);
nand U9173 (N_9173,N_8870,N_8968);
nor U9174 (N_9174,N_8898,N_8970);
nor U9175 (N_9175,N_8989,N_8815);
xnor U9176 (N_9176,N_8906,N_8867);
or U9177 (N_9177,N_8810,N_8860);
nand U9178 (N_9178,N_8922,N_8839);
or U9179 (N_9179,N_8939,N_8941);
or U9180 (N_9180,N_8820,N_8932);
and U9181 (N_9181,N_8806,N_8847);
nor U9182 (N_9182,N_8992,N_8976);
and U9183 (N_9183,N_8983,N_8904);
and U9184 (N_9184,N_8978,N_8936);
and U9185 (N_9185,N_8944,N_8915);
and U9186 (N_9186,N_8905,N_8804);
nand U9187 (N_9187,N_8935,N_8802);
nand U9188 (N_9188,N_8928,N_8820);
and U9189 (N_9189,N_8863,N_8801);
and U9190 (N_9190,N_8822,N_8975);
nor U9191 (N_9191,N_8860,N_8978);
nand U9192 (N_9192,N_8893,N_8853);
or U9193 (N_9193,N_8869,N_8897);
nand U9194 (N_9194,N_8971,N_8824);
or U9195 (N_9195,N_8909,N_8913);
and U9196 (N_9196,N_8824,N_8924);
and U9197 (N_9197,N_8859,N_8819);
nand U9198 (N_9198,N_8824,N_8837);
nor U9199 (N_9199,N_8979,N_8897);
or U9200 (N_9200,N_9044,N_9052);
nand U9201 (N_9201,N_9089,N_9090);
nand U9202 (N_9202,N_9159,N_9108);
nand U9203 (N_9203,N_9135,N_9158);
or U9204 (N_9204,N_9098,N_9039);
nand U9205 (N_9205,N_9035,N_9000);
and U9206 (N_9206,N_9173,N_9130);
nor U9207 (N_9207,N_9085,N_9147);
or U9208 (N_9208,N_9177,N_9183);
and U9209 (N_9209,N_9049,N_9061);
xnor U9210 (N_9210,N_9124,N_9042);
and U9211 (N_9211,N_9146,N_9080);
nand U9212 (N_9212,N_9003,N_9104);
and U9213 (N_9213,N_9005,N_9015);
and U9214 (N_9214,N_9144,N_9188);
and U9215 (N_9215,N_9161,N_9165);
nand U9216 (N_9216,N_9132,N_9154);
nor U9217 (N_9217,N_9068,N_9156);
and U9218 (N_9218,N_9100,N_9187);
xor U9219 (N_9219,N_9181,N_9055);
nand U9220 (N_9220,N_9109,N_9025);
or U9221 (N_9221,N_9081,N_9167);
and U9222 (N_9222,N_9024,N_9107);
nor U9223 (N_9223,N_9071,N_9134);
nand U9224 (N_9224,N_9149,N_9190);
nand U9225 (N_9225,N_9191,N_9194);
or U9226 (N_9226,N_9155,N_9007);
nor U9227 (N_9227,N_9133,N_9150);
and U9228 (N_9228,N_9182,N_9162);
nor U9229 (N_9229,N_9066,N_9057);
and U9230 (N_9230,N_9063,N_9004);
nand U9231 (N_9231,N_9119,N_9088);
nor U9232 (N_9232,N_9112,N_9127);
or U9233 (N_9233,N_9169,N_9197);
nand U9234 (N_9234,N_9062,N_9185);
nand U9235 (N_9235,N_9117,N_9189);
nor U9236 (N_9236,N_9184,N_9067);
or U9237 (N_9237,N_9125,N_9170);
and U9238 (N_9238,N_9145,N_9141);
nor U9239 (N_9239,N_9199,N_9139);
or U9240 (N_9240,N_9102,N_9023);
nor U9241 (N_9241,N_9010,N_9195);
and U9242 (N_9242,N_9020,N_9048);
or U9243 (N_9243,N_9163,N_9040);
or U9244 (N_9244,N_9050,N_9019);
and U9245 (N_9245,N_9120,N_9175);
nor U9246 (N_9246,N_9017,N_9101);
or U9247 (N_9247,N_9051,N_9069);
nor U9248 (N_9248,N_9168,N_9002);
nand U9249 (N_9249,N_9001,N_9128);
nand U9250 (N_9250,N_9093,N_9111);
nor U9251 (N_9251,N_9045,N_9014);
and U9252 (N_9252,N_9073,N_9129);
or U9253 (N_9253,N_9043,N_9118);
or U9254 (N_9254,N_9131,N_9065);
nand U9255 (N_9255,N_9114,N_9030);
or U9256 (N_9256,N_9011,N_9008);
and U9257 (N_9257,N_9026,N_9121);
and U9258 (N_9258,N_9196,N_9126);
or U9259 (N_9259,N_9054,N_9157);
and U9260 (N_9260,N_9099,N_9013);
nand U9261 (N_9261,N_9077,N_9031);
or U9262 (N_9262,N_9174,N_9105);
nand U9263 (N_9263,N_9009,N_9122);
nor U9264 (N_9264,N_9038,N_9072);
nor U9265 (N_9265,N_9036,N_9091);
nand U9266 (N_9266,N_9138,N_9016);
and U9267 (N_9267,N_9106,N_9083);
nor U9268 (N_9268,N_9171,N_9164);
nor U9269 (N_9269,N_9092,N_9074);
nand U9270 (N_9270,N_9041,N_9153);
and U9271 (N_9271,N_9186,N_9053);
and U9272 (N_9272,N_9151,N_9059);
nand U9273 (N_9273,N_9137,N_9070);
and U9274 (N_9274,N_9096,N_9198);
and U9275 (N_9275,N_9027,N_9094);
nor U9276 (N_9276,N_9113,N_9136);
nor U9277 (N_9277,N_9082,N_9116);
or U9278 (N_9278,N_9152,N_9103);
nor U9279 (N_9279,N_9058,N_9097);
nor U9280 (N_9280,N_9032,N_9047);
nand U9281 (N_9281,N_9148,N_9084);
nand U9282 (N_9282,N_9095,N_9078);
and U9283 (N_9283,N_9110,N_9076);
nand U9284 (N_9284,N_9123,N_9022);
nand U9285 (N_9285,N_9018,N_9086);
nand U9286 (N_9286,N_9115,N_9046);
nand U9287 (N_9287,N_9006,N_9142);
nor U9288 (N_9288,N_9021,N_9075);
nand U9289 (N_9289,N_9160,N_9192);
or U9290 (N_9290,N_9179,N_9178);
or U9291 (N_9291,N_9176,N_9033);
nand U9292 (N_9292,N_9029,N_9166);
or U9293 (N_9293,N_9064,N_9172);
nand U9294 (N_9294,N_9028,N_9060);
and U9295 (N_9295,N_9012,N_9079);
nand U9296 (N_9296,N_9193,N_9087);
or U9297 (N_9297,N_9037,N_9143);
and U9298 (N_9298,N_9056,N_9180);
nand U9299 (N_9299,N_9034,N_9140);
nor U9300 (N_9300,N_9106,N_9003);
and U9301 (N_9301,N_9065,N_9174);
nand U9302 (N_9302,N_9103,N_9120);
or U9303 (N_9303,N_9093,N_9006);
nor U9304 (N_9304,N_9129,N_9001);
nand U9305 (N_9305,N_9086,N_9155);
nor U9306 (N_9306,N_9034,N_9188);
nor U9307 (N_9307,N_9196,N_9121);
or U9308 (N_9308,N_9103,N_9141);
nand U9309 (N_9309,N_9086,N_9157);
and U9310 (N_9310,N_9024,N_9121);
or U9311 (N_9311,N_9198,N_9080);
or U9312 (N_9312,N_9041,N_9005);
or U9313 (N_9313,N_9136,N_9142);
nand U9314 (N_9314,N_9142,N_9108);
and U9315 (N_9315,N_9138,N_9169);
nand U9316 (N_9316,N_9071,N_9179);
nor U9317 (N_9317,N_9158,N_9076);
nor U9318 (N_9318,N_9168,N_9142);
nor U9319 (N_9319,N_9185,N_9194);
or U9320 (N_9320,N_9066,N_9027);
nand U9321 (N_9321,N_9185,N_9187);
or U9322 (N_9322,N_9035,N_9091);
or U9323 (N_9323,N_9187,N_9021);
and U9324 (N_9324,N_9079,N_9042);
nand U9325 (N_9325,N_9078,N_9136);
nor U9326 (N_9326,N_9120,N_9110);
nand U9327 (N_9327,N_9050,N_9023);
xnor U9328 (N_9328,N_9104,N_9172);
or U9329 (N_9329,N_9077,N_9022);
or U9330 (N_9330,N_9047,N_9187);
nor U9331 (N_9331,N_9022,N_9031);
nand U9332 (N_9332,N_9041,N_9118);
or U9333 (N_9333,N_9017,N_9119);
nand U9334 (N_9334,N_9140,N_9129);
nor U9335 (N_9335,N_9081,N_9109);
and U9336 (N_9336,N_9022,N_9191);
and U9337 (N_9337,N_9143,N_9115);
and U9338 (N_9338,N_9153,N_9117);
nor U9339 (N_9339,N_9024,N_9012);
nand U9340 (N_9340,N_9093,N_9041);
or U9341 (N_9341,N_9051,N_9086);
nand U9342 (N_9342,N_9015,N_9094);
xnor U9343 (N_9343,N_9158,N_9117);
and U9344 (N_9344,N_9092,N_9100);
or U9345 (N_9345,N_9138,N_9050);
nand U9346 (N_9346,N_9096,N_9132);
nand U9347 (N_9347,N_9140,N_9008);
nand U9348 (N_9348,N_9025,N_9090);
nand U9349 (N_9349,N_9163,N_9089);
nor U9350 (N_9350,N_9052,N_9091);
and U9351 (N_9351,N_9182,N_9049);
nor U9352 (N_9352,N_9086,N_9139);
nand U9353 (N_9353,N_9024,N_9074);
nand U9354 (N_9354,N_9129,N_9053);
nand U9355 (N_9355,N_9077,N_9089);
and U9356 (N_9356,N_9144,N_9056);
or U9357 (N_9357,N_9051,N_9095);
nand U9358 (N_9358,N_9013,N_9171);
or U9359 (N_9359,N_9087,N_9003);
nor U9360 (N_9360,N_9097,N_9053);
nand U9361 (N_9361,N_9057,N_9049);
and U9362 (N_9362,N_9196,N_9164);
nor U9363 (N_9363,N_9090,N_9092);
nand U9364 (N_9364,N_9177,N_9106);
nand U9365 (N_9365,N_9092,N_9197);
or U9366 (N_9366,N_9191,N_9079);
and U9367 (N_9367,N_9030,N_9016);
and U9368 (N_9368,N_9197,N_9053);
nand U9369 (N_9369,N_9124,N_9118);
or U9370 (N_9370,N_9058,N_9069);
and U9371 (N_9371,N_9158,N_9010);
nor U9372 (N_9372,N_9184,N_9135);
or U9373 (N_9373,N_9022,N_9089);
or U9374 (N_9374,N_9162,N_9049);
and U9375 (N_9375,N_9176,N_9029);
nor U9376 (N_9376,N_9137,N_9076);
nand U9377 (N_9377,N_9133,N_9152);
nor U9378 (N_9378,N_9032,N_9190);
or U9379 (N_9379,N_9035,N_9171);
nor U9380 (N_9380,N_9186,N_9119);
and U9381 (N_9381,N_9068,N_9155);
nand U9382 (N_9382,N_9190,N_9151);
and U9383 (N_9383,N_9128,N_9106);
nor U9384 (N_9384,N_9057,N_9040);
and U9385 (N_9385,N_9072,N_9181);
and U9386 (N_9386,N_9016,N_9089);
or U9387 (N_9387,N_9065,N_9004);
or U9388 (N_9388,N_9129,N_9064);
and U9389 (N_9389,N_9162,N_9186);
or U9390 (N_9390,N_9062,N_9134);
nor U9391 (N_9391,N_9042,N_9088);
or U9392 (N_9392,N_9158,N_9163);
nor U9393 (N_9393,N_9124,N_9166);
nand U9394 (N_9394,N_9125,N_9054);
nand U9395 (N_9395,N_9026,N_9188);
or U9396 (N_9396,N_9197,N_9029);
or U9397 (N_9397,N_9118,N_9113);
nand U9398 (N_9398,N_9199,N_9179);
or U9399 (N_9399,N_9175,N_9075);
and U9400 (N_9400,N_9252,N_9399);
or U9401 (N_9401,N_9356,N_9218);
nor U9402 (N_9402,N_9326,N_9306);
nor U9403 (N_9403,N_9290,N_9340);
nor U9404 (N_9404,N_9271,N_9219);
nor U9405 (N_9405,N_9257,N_9342);
or U9406 (N_9406,N_9328,N_9231);
nand U9407 (N_9407,N_9253,N_9280);
and U9408 (N_9408,N_9311,N_9343);
nand U9409 (N_9409,N_9386,N_9235);
or U9410 (N_9410,N_9313,N_9350);
and U9411 (N_9411,N_9293,N_9322);
nor U9412 (N_9412,N_9375,N_9250);
or U9413 (N_9413,N_9345,N_9241);
or U9414 (N_9414,N_9330,N_9384);
or U9415 (N_9415,N_9365,N_9292);
nor U9416 (N_9416,N_9381,N_9305);
nor U9417 (N_9417,N_9207,N_9315);
or U9418 (N_9418,N_9352,N_9244);
nand U9419 (N_9419,N_9216,N_9211);
nor U9420 (N_9420,N_9301,N_9310);
nand U9421 (N_9421,N_9254,N_9300);
nand U9422 (N_9422,N_9243,N_9391);
and U9423 (N_9423,N_9288,N_9261);
and U9424 (N_9424,N_9388,N_9284);
nand U9425 (N_9425,N_9298,N_9251);
or U9426 (N_9426,N_9237,N_9378);
xnor U9427 (N_9427,N_9291,N_9377);
and U9428 (N_9428,N_9239,N_9255);
or U9429 (N_9429,N_9323,N_9361);
nor U9430 (N_9430,N_9238,N_9389);
and U9431 (N_9431,N_9351,N_9396);
nand U9432 (N_9432,N_9325,N_9287);
or U9433 (N_9433,N_9208,N_9312);
nor U9434 (N_9434,N_9303,N_9392);
and U9435 (N_9435,N_9339,N_9282);
nand U9436 (N_9436,N_9379,N_9265);
and U9437 (N_9437,N_9225,N_9245);
nor U9438 (N_9438,N_9358,N_9240);
nor U9439 (N_9439,N_9316,N_9318);
or U9440 (N_9440,N_9324,N_9349);
nand U9441 (N_9441,N_9275,N_9363);
nor U9442 (N_9442,N_9354,N_9299);
or U9443 (N_9443,N_9232,N_9209);
nor U9444 (N_9444,N_9314,N_9387);
nor U9445 (N_9445,N_9226,N_9228);
and U9446 (N_9446,N_9248,N_9360);
nand U9447 (N_9447,N_9395,N_9373);
nand U9448 (N_9448,N_9344,N_9274);
and U9449 (N_9449,N_9327,N_9269);
nor U9450 (N_9450,N_9286,N_9260);
or U9451 (N_9451,N_9385,N_9236);
or U9452 (N_9452,N_9304,N_9266);
or U9453 (N_9453,N_9234,N_9337);
or U9454 (N_9454,N_9294,N_9206);
and U9455 (N_9455,N_9268,N_9202);
nor U9456 (N_9456,N_9222,N_9224);
or U9457 (N_9457,N_9347,N_9259);
and U9458 (N_9458,N_9215,N_9364);
nand U9459 (N_9459,N_9263,N_9267);
nand U9460 (N_9460,N_9247,N_9217);
and U9461 (N_9461,N_9276,N_9397);
and U9462 (N_9462,N_9264,N_9338);
and U9463 (N_9463,N_9331,N_9212);
nor U9464 (N_9464,N_9332,N_9289);
and U9465 (N_9465,N_9201,N_9205);
or U9466 (N_9466,N_9355,N_9213);
nor U9467 (N_9467,N_9273,N_9229);
nand U9468 (N_9468,N_9204,N_9302);
nor U9469 (N_9469,N_9249,N_9336);
and U9470 (N_9470,N_9262,N_9348);
nor U9471 (N_9471,N_9281,N_9285);
and U9472 (N_9472,N_9200,N_9320);
nor U9473 (N_9473,N_9221,N_9278);
and U9474 (N_9474,N_9359,N_9321);
and U9475 (N_9475,N_9214,N_9370);
and U9476 (N_9476,N_9242,N_9258);
nand U9477 (N_9477,N_9296,N_9371);
and U9478 (N_9478,N_9367,N_9279);
nor U9479 (N_9479,N_9390,N_9246);
xnor U9480 (N_9480,N_9256,N_9334);
and U9481 (N_9481,N_9295,N_9307);
or U9482 (N_9482,N_9394,N_9227);
nand U9483 (N_9483,N_9357,N_9270);
or U9484 (N_9484,N_9335,N_9398);
nand U9485 (N_9485,N_9346,N_9210);
nor U9486 (N_9486,N_9297,N_9376);
or U9487 (N_9487,N_9341,N_9308);
nor U9488 (N_9488,N_9372,N_9380);
or U9489 (N_9489,N_9309,N_9283);
and U9490 (N_9490,N_9220,N_9317);
nor U9491 (N_9491,N_9223,N_9329);
and U9492 (N_9492,N_9362,N_9277);
nor U9493 (N_9493,N_9374,N_9369);
nand U9494 (N_9494,N_9272,N_9366);
nand U9495 (N_9495,N_9353,N_9319);
or U9496 (N_9496,N_9230,N_9383);
nor U9497 (N_9497,N_9393,N_9203);
nor U9498 (N_9498,N_9368,N_9333);
nand U9499 (N_9499,N_9382,N_9233);
or U9500 (N_9500,N_9345,N_9325);
nor U9501 (N_9501,N_9361,N_9299);
and U9502 (N_9502,N_9285,N_9311);
nand U9503 (N_9503,N_9224,N_9207);
or U9504 (N_9504,N_9220,N_9319);
nor U9505 (N_9505,N_9283,N_9302);
nand U9506 (N_9506,N_9237,N_9245);
and U9507 (N_9507,N_9349,N_9331);
nor U9508 (N_9508,N_9217,N_9320);
and U9509 (N_9509,N_9208,N_9214);
or U9510 (N_9510,N_9384,N_9297);
or U9511 (N_9511,N_9323,N_9246);
and U9512 (N_9512,N_9398,N_9298);
and U9513 (N_9513,N_9258,N_9212);
nand U9514 (N_9514,N_9261,N_9212);
and U9515 (N_9515,N_9211,N_9373);
and U9516 (N_9516,N_9292,N_9256);
or U9517 (N_9517,N_9343,N_9338);
and U9518 (N_9518,N_9215,N_9207);
nor U9519 (N_9519,N_9249,N_9384);
nor U9520 (N_9520,N_9286,N_9282);
or U9521 (N_9521,N_9356,N_9393);
nor U9522 (N_9522,N_9242,N_9298);
nand U9523 (N_9523,N_9362,N_9273);
and U9524 (N_9524,N_9364,N_9311);
or U9525 (N_9525,N_9245,N_9296);
or U9526 (N_9526,N_9220,N_9235);
nand U9527 (N_9527,N_9300,N_9362);
or U9528 (N_9528,N_9223,N_9396);
or U9529 (N_9529,N_9324,N_9354);
or U9530 (N_9530,N_9339,N_9338);
nand U9531 (N_9531,N_9225,N_9256);
or U9532 (N_9532,N_9243,N_9221);
nand U9533 (N_9533,N_9202,N_9326);
nor U9534 (N_9534,N_9393,N_9270);
or U9535 (N_9535,N_9209,N_9379);
and U9536 (N_9536,N_9220,N_9329);
or U9537 (N_9537,N_9238,N_9314);
or U9538 (N_9538,N_9333,N_9226);
and U9539 (N_9539,N_9201,N_9274);
nand U9540 (N_9540,N_9269,N_9257);
and U9541 (N_9541,N_9222,N_9277);
nand U9542 (N_9542,N_9284,N_9270);
nor U9543 (N_9543,N_9337,N_9306);
nor U9544 (N_9544,N_9213,N_9325);
or U9545 (N_9545,N_9265,N_9380);
and U9546 (N_9546,N_9380,N_9261);
nor U9547 (N_9547,N_9265,N_9285);
or U9548 (N_9548,N_9338,N_9279);
nor U9549 (N_9549,N_9361,N_9392);
nor U9550 (N_9550,N_9330,N_9275);
nor U9551 (N_9551,N_9282,N_9398);
and U9552 (N_9552,N_9389,N_9231);
or U9553 (N_9553,N_9307,N_9288);
nor U9554 (N_9554,N_9290,N_9276);
or U9555 (N_9555,N_9251,N_9379);
nand U9556 (N_9556,N_9366,N_9204);
and U9557 (N_9557,N_9206,N_9398);
or U9558 (N_9558,N_9287,N_9227);
or U9559 (N_9559,N_9250,N_9243);
or U9560 (N_9560,N_9293,N_9287);
and U9561 (N_9561,N_9343,N_9367);
or U9562 (N_9562,N_9233,N_9311);
and U9563 (N_9563,N_9314,N_9375);
nand U9564 (N_9564,N_9321,N_9238);
nand U9565 (N_9565,N_9312,N_9212);
nand U9566 (N_9566,N_9326,N_9393);
nor U9567 (N_9567,N_9340,N_9356);
nor U9568 (N_9568,N_9387,N_9201);
and U9569 (N_9569,N_9335,N_9372);
nor U9570 (N_9570,N_9373,N_9252);
or U9571 (N_9571,N_9285,N_9372);
and U9572 (N_9572,N_9325,N_9310);
or U9573 (N_9573,N_9277,N_9256);
nand U9574 (N_9574,N_9379,N_9271);
nor U9575 (N_9575,N_9249,N_9374);
nand U9576 (N_9576,N_9386,N_9224);
and U9577 (N_9577,N_9211,N_9329);
xnor U9578 (N_9578,N_9291,N_9218);
nand U9579 (N_9579,N_9265,N_9309);
or U9580 (N_9580,N_9349,N_9308);
and U9581 (N_9581,N_9288,N_9227);
or U9582 (N_9582,N_9209,N_9352);
or U9583 (N_9583,N_9201,N_9209);
or U9584 (N_9584,N_9249,N_9223);
and U9585 (N_9585,N_9228,N_9206);
nand U9586 (N_9586,N_9206,N_9263);
and U9587 (N_9587,N_9281,N_9392);
nand U9588 (N_9588,N_9310,N_9233);
nand U9589 (N_9589,N_9339,N_9279);
nor U9590 (N_9590,N_9264,N_9310);
nand U9591 (N_9591,N_9214,N_9243);
nor U9592 (N_9592,N_9204,N_9251);
and U9593 (N_9593,N_9285,N_9262);
nand U9594 (N_9594,N_9227,N_9387);
or U9595 (N_9595,N_9354,N_9338);
nor U9596 (N_9596,N_9320,N_9230);
and U9597 (N_9597,N_9222,N_9241);
nor U9598 (N_9598,N_9398,N_9255);
nor U9599 (N_9599,N_9257,N_9365);
nor U9600 (N_9600,N_9430,N_9426);
or U9601 (N_9601,N_9586,N_9570);
and U9602 (N_9602,N_9551,N_9478);
or U9603 (N_9603,N_9501,N_9591);
and U9604 (N_9604,N_9552,N_9406);
nor U9605 (N_9605,N_9487,N_9491);
or U9606 (N_9606,N_9483,N_9416);
and U9607 (N_9607,N_9454,N_9549);
nand U9608 (N_9608,N_9543,N_9578);
nor U9609 (N_9609,N_9488,N_9444);
and U9610 (N_9610,N_9503,N_9525);
or U9611 (N_9611,N_9489,N_9598);
and U9612 (N_9612,N_9412,N_9485);
and U9613 (N_9613,N_9472,N_9481);
or U9614 (N_9614,N_9475,N_9474);
nand U9615 (N_9615,N_9523,N_9568);
or U9616 (N_9616,N_9431,N_9419);
nand U9617 (N_9617,N_9470,N_9415);
nand U9618 (N_9618,N_9544,N_9413);
and U9619 (N_9619,N_9467,N_9546);
nor U9620 (N_9620,N_9461,N_9471);
nand U9621 (N_9621,N_9443,N_9548);
or U9622 (N_9622,N_9580,N_9417);
nor U9623 (N_9623,N_9505,N_9533);
xnor U9624 (N_9624,N_9411,N_9482);
or U9625 (N_9625,N_9421,N_9409);
nor U9626 (N_9626,N_9433,N_9539);
and U9627 (N_9627,N_9537,N_9404);
nor U9628 (N_9628,N_9418,N_9506);
nand U9629 (N_9629,N_9561,N_9439);
nand U9630 (N_9630,N_9516,N_9555);
and U9631 (N_9631,N_9550,N_9473);
or U9632 (N_9632,N_9596,N_9542);
and U9633 (N_9633,N_9521,N_9587);
nor U9634 (N_9634,N_9447,N_9502);
xor U9635 (N_9635,N_9480,N_9595);
or U9636 (N_9636,N_9508,N_9532);
nor U9637 (N_9637,N_9520,N_9469);
or U9638 (N_9638,N_9420,N_9466);
nand U9639 (N_9639,N_9517,N_9510);
or U9640 (N_9640,N_9524,N_9445);
nand U9641 (N_9641,N_9424,N_9455);
nor U9642 (N_9642,N_9526,N_9559);
nor U9643 (N_9643,N_9460,N_9400);
nand U9644 (N_9644,N_9541,N_9574);
nand U9645 (N_9645,N_9442,N_9512);
and U9646 (N_9646,N_9435,N_9434);
nand U9647 (N_9647,N_9545,N_9499);
and U9648 (N_9648,N_9402,N_9518);
and U9649 (N_9649,N_9438,N_9407);
or U9650 (N_9650,N_9590,N_9448);
or U9651 (N_9651,N_9450,N_9437);
or U9652 (N_9652,N_9563,N_9515);
nand U9653 (N_9653,N_9408,N_9560);
nand U9654 (N_9654,N_9441,N_9527);
nand U9655 (N_9655,N_9522,N_9562);
nand U9656 (N_9656,N_9565,N_9556);
and U9657 (N_9657,N_9540,N_9584);
nor U9658 (N_9658,N_9476,N_9456);
or U9659 (N_9659,N_9405,N_9597);
nor U9660 (N_9660,N_9534,N_9449);
and U9661 (N_9661,N_9509,N_9589);
or U9662 (N_9662,N_9464,N_9423);
or U9663 (N_9663,N_9538,N_9484);
nor U9664 (N_9664,N_9529,N_9576);
nand U9665 (N_9665,N_9494,N_9429);
nor U9666 (N_9666,N_9414,N_9566);
nand U9667 (N_9667,N_9577,N_9585);
or U9668 (N_9668,N_9492,N_9453);
nand U9669 (N_9669,N_9468,N_9452);
nand U9670 (N_9670,N_9451,N_9536);
nand U9671 (N_9671,N_9582,N_9401);
nor U9672 (N_9672,N_9519,N_9479);
and U9673 (N_9673,N_9462,N_9547);
or U9674 (N_9674,N_9496,N_9528);
and U9675 (N_9675,N_9511,N_9531);
nand U9676 (N_9676,N_9514,N_9436);
nor U9677 (N_9677,N_9463,N_9573);
nor U9678 (N_9678,N_9507,N_9572);
and U9679 (N_9679,N_9567,N_9569);
or U9680 (N_9680,N_9457,N_9497);
nor U9681 (N_9681,N_9459,N_9465);
or U9682 (N_9682,N_9490,N_9403);
nand U9683 (N_9683,N_9557,N_9535);
nor U9684 (N_9684,N_9422,N_9493);
nand U9685 (N_9685,N_9575,N_9440);
xnor U9686 (N_9686,N_9504,N_9583);
nor U9687 (N_9687,N_9599,N_9458);
or U9688 (N_9688,N_9410,N_9593);
nand U9689 (N_9689,N_9500,N_9495);
and U9690 (N_9690,N_9594,N_9432);
and U9691 (N_9691,N_9428,N_9498);
and U9692 (N_9692,N_9427,N_9530);
and U9693 (N_9693,N_9446,N_9588);
and U9694 (N_9694,N_9513,N_9579);
nor U9695 (N_9695,N_9564,N_9554);
and U9696 (N_9696,N_9581,N_9571);
nor U9697 (N_9697,N_9486,N_9425);
nor U9698 (N_9698,N_9592,N_9558);
nand U9699 (N_9699,N_9477,N_9553);
nor U9700 (N_9700,N_9583,N_9459);
nand U9701 (N_9701,N_9507,N_9433);
nand U9702 (N_9702,N_9446,N_9438);
nor U9703 (N_9703,N_9567,N_9596);
nand U9704 (N_9704,N_9543,N_9437);
nor U9705 (N_9705,N_9585,N_9473);
nor U9706 (N_9706,N_9435,N_9403);
nor U9707 (N_9707,N_9532,N_9538);
and U9708 (N_9708,N_9436,N_9528);
and U9709 (N_9709,N_9536,N_9503);
and U9710 (N_9710,N_9446,N_9454);
nand U9711 (N_9711,N_9510,N_9541);
and U9712 (N_9712,N_9432,N_9512);
nand U9713 (N_9713,N_9407,N_9481);
nand U9714 (N_9714,N_9471,N_9424);
and U9715 (N_9715,N_9569,N_9556);
nand U9716 (N_9716,N_9563,N_9481);
and U9717 (N_9717,N_9514,N_9494);
or U9718 (N_9718,N_9469,N_9521);
and U9719 (N_9719,N_9592,N_9419);
nor U9720 (N_9720,N_9530,N_9456);
or U9721 (N_9721,N_9437,N_9418);
nand U9722 (N_9722,N_9545,N_9403);
and U9723 (N_9723,N_9452,N_9587);
nor U9724 (N_9724,N_9556,N_9511);
and U9725 (N_9725,N_9413,N_9560);
nor U9726 (N_9726,N_9591,N_9441);
nor U9727 (N_9727,N_9543,N_9550);
and U9728 (N_9728,N_9408,N_9467);
and U9729 (N_9729,N_9549,N_9515);
or U9730 (N_9730,N_9491,N_9572);
nand U9731 (N_9731,N_9405,N_9509);
nand U9732 (N_9732,N_9536,N_9457);
and U9733 (N_9733,N_9417,N_9491);
xor U9734 (N_9734,N_9409,N_9552);
nor U9735 (N_9735,N_9531,N_9427);
and U9736 (N_9736,N_9556,N_9552);
nand U9737 (N_9737,N_9438,N_9595);
xnor U9738 (N_9738,N_9530,N_9509);
nand U9739 (N_9739,N_9485,N_9425);
and U9740 (N_9740,N_9428,N_9431);
or U9741 (N_9741,N_9402,N_9468);
or U9742 (N_9742,N_9410,N_9543);
nor U9743 (N_9743,N_9553,N_9459);
nor U9744 (N_9744,N_9462,N_9430);
nor U9745 (N_9745,N_9468,N_9472);
or U9746 (N_9746,N_9523,N_9483);
or U9747 (N_9747,N_9481,N_9566);
nor U9748 (N_9748,N_9505,N_9446);
and U9749 (N_9749,N_9521,N_9502);
nand U9750 (N_9750,N_9593,N_9527);
or U9751 (N_9751,N_9523,N_9484);
nand U9752 (N_9752,N_9532,N_9456);
or U9753 (N_9753,N_9512,N_9447);
or U9754 (N_9754,N_9504,N_9425);
nor U9755 (N_9755,N_9527,N_9508);
and U9756 (N_9756,N_9491,N_9482);
nor U9757 (N_9757,N_9573,N_9587);
nor U9758 (N_9758,N_9525,N_9411);
nand U9759 (N_9759,N_9403,N_9462);
nand U9760 (N_9760,N_9537,N_9540);
or U9761 (N_9761,N_9499,N_9451);
nor U9762 (N_9762,N_9426,N_9503);
nor U9763 (N_9763,N_9503,N_9512);
or U9764 (N_9764,N_9517,N_9456);
and U9765 (N_9765,N_9476,N_9566);
or U9766 (N_9766,N_9579,N_9458);
or U9767 (N_9767,N_9422,N_9547);
nand U9768 (N_9768,N_9458,N_9517);
or U9769 (N_9769,N_9424,N_9420);
and U9770 (N_9770,N_9540,N_9535);
or U9771 (N_9771,N_9481,N_9519);
nor U9772 (N_9772,N_9500,N_9508);
and U9773 (N_9773,N_9415,N_9546);
and U9774 (N_9774,N_9515,N_9577);
or U9775 (N_9775,N_9428,N_9494);
or U9776 (N_9776,N_9437,N_9596);
and U9777 (N_9777,N_9404,N_9499);
nand U9778 (N_9778,N_9412,N_9556);
or U9779 (N_9779,N_9529,N_9515);
and U9780 (N_9780,N_9526,N_9463);
nor U9781 (N_9781,N_9468,N_9540);
nor U9782 (N_9782,N_9547,N_9581);
or U9783 (N_9783,N_9428,N_9416);
and U9784 (N_9784,N_9440,N_9503);
or U9785 (N_9785,N_9485,N_9530);
or U9786 (N_9786,N_9537,N_9592);
or U9787 (N_9787,N_9483,N_9575);
or U9788 (N_9788,N_9550,N_9422);
nand U9789 (N_9789,N_9517,N_9489);
nand U9790 (N_9790,N_9596,N_9455);
and U9791 (N_9791,N_9411,N_9486);
and U9792 (N_9792,N_9448,N_9469);
nor U9793 (N_9793,N_9433,N_9523);
and U9794 (N_9794,N_9476,N_9409);
or U9795 (N_9795,N_9453,N_9598);
nor U9796 (N_9796,N_9531,N_9450);
and U9797 (N_9797,N_9415,N_9439);
or U9798 (N_9798,N_9557,N_9571);
nor U9799 (N_9799,N_9577,N_9573);
or U9800 (N_9800,N_9714,N_9782);
or U9801 (N_9801,N_9632,N_9662);
or U9802 (N_9802,N_9787,N_9688);
or U9803 (N_9803,N_9701,N_9677);
and U9804 (N_9804,N_9682,N_9678);
or U9805 (N_9805,N_9692,N_9654);
and U9806 (N_9806,N_9746,N_9699);
nor U9807 (N_9807,N_9736,N_9656);
or U9808 (N_9808,N_9653,N_9716);
or U9809 (N_9809,N_9764,N_9695);
nor U9810 (N_9810,N_9633,N_9747);
or U9811 (N_9811,N_9786,N_9655);
nand U9812 (N_9812,N_9759,N_9603);
nand U9813 (N_9813,N_9608,N_9720);
nor U9814 (N_9814,N_9730,N_9700);
nor U9815 (N_9815,N_9740,N_9733);
nor U9816 (N_9816,N_9774,N_9789);
or U9817 (N_9817,N_9694,N_9673);
and U9818 (N_9818,N_9659,N_9643);
nor U9819 (N_9819,N_9609,N_9616);
or U9820 (N_9820,N_9766,N_9696);
nand U9821 (N_9821,N_9621,N_9624);
nand U9822 (N_9822,N_9638,N_9640);
nor U9823 (N_9823,N_9614,N_9718);
or U9824 (N_9824,N_9630,N_9672);
and U9825 (N_9825,N_9618,N_9732);
and U9826 (N_9826,N_9708,N_9785);
nor U9827 (N_9827,N_9623,N_9619);
or U9828 (N_9828,N_9681,N_9639);
and U9829 (N_9829,N_9757,N_9684);
nand U9830 (N_9830,N_9778,N_9601);
or U9831 (N_9831,N_9652,N_9791);
or U9832 (N_9832,N_9669,N_9602);
nor U9833 (N_9833,N_9750,N_9650);
nand U9834 (N_9834,N_9731,N_9600);
nand U9835 (N_9835,N_9610,N_9768);
or U9836 (N_9836,N_9749,N_9751);
and U9837 (N_9837,N_9710,N_9685);
nor U9838 (N_9838,N_9691,N_9664);
nand U9839 (N_9839,N_9668,N_9661);
and U9840 (N_9840,N_9741,N_9698);
nand U9841 (N_9841,N_9707,N_9671);
nand U9842 (N_9842,N_9713,N_9617);
nand U9843 (N_9843,N_9753,N_9756);
nor U9844 (N_9844,N_9611,N_9796);
and U9845 (N_9845,N_9667,N_9663);
nand U9846 (N_9846,N_9739,N_9779);
nor U9847 (N_9847,N_9674,N_9675);
nand U9848 (N_9848,N_9792,N_9709);
and U9849 (N_9849,N_9666,N_9765);
nor U9850 (N_9850,N_9615,N_9712);
nand U9851 (N_9851,N_9752,N_9689);
nor U9852 (N_9852,N_9795,N_9705);
nand U9853 (N_9853,N_9797,N_9637);
or U9854 (N_9854,N_9612,N_9729);
or U9855 (N_9855,N_9620,N_9651);
and U9856 (N_9856,N_9613,N_9735);
nand U9857 (N_9857,N_9636,N_9683);
or U9858 (N_9858,N_9760,N_9676);
and U9859 (N_9859,N_9743,N_9706);
nand U9860 (N_9860,N_9755,N_9727);
nor U9861 (N_9861,N_9771,N_9649);
or U9862 (N_9862,N_9780,N_9728);
and U9863 (N_9863,N_9784,N_9629);
nor U9864 (N_9864,N_9723,N_9690);
nand U9865 (N_9865,N_9607,N_9679);
nor U9866 (N_9866,N_9622,N_9634);
nor U9867 (N_9867,N_9646,N_9758);
nand U9868 (N_9868,N_9790,N_9604);
nor U9869 (N_9869,N_9631,N_9793);
nand U9870 (N_9870,N_9773,N_9658);
and U9871 (N_9871,N_9697,N_9794);
nor U9872 (N_9872,N_9719,N_9722);
or U9873 (N_9873,N_9703,N_9648);
nor U9874 (N_9874,N_9645,N_9738);
nor U9875 (N_9875,N_9744,N_9776);
or U9876 (N_9876,N_9641,N_9721);
or U9877 (N_9877,N_9665,N_9625);
nor U9878 (N_9878,N_9702,N_9783);
and U9879 (N_9879,N_9627,N_9660);
or U9880 (N_9880,N_9670,N_9686);
or U9881 (N_9881,N_9724,N_9788);
nand U9882 (N_9882,N_9799,N_9777);
or U9883 (N_9883,N_9606,N_9647);
or U9884 (N_9884,N_9769,N_9711);
and U9885 (N_9885,N_9715,N_9680);
nor U9886 (N_9886,N_9772,N_9642);
and U9887 (N_9887,N_9754,N_9767);
nor U9888 (N_9888,N_9770,N_9635);
and U9889 (N_9889,N_9762,N_9693);
nor U9890 (N_9890,N_9605,N_9644);
nand U9891 (N_9891,N_9781,N_9726);
nand U9892 (N_9892,N_9725,N_9737);
or U9893 (N_9893,N_9657,N_9687);
nor U9894 (N_9894,N_9734,N_9745);
and U9895 (N_9895,N_9628,N_9704);
or U9896 (N_9896,N_9775,N_9626);
and U9897 (N_9897,N_9761,N_9748);
xor U9898 (N_9898,N_9717,N_9742);
xnor U9899 (N_9899,N_9763,N_9798);
and U9900 (N_9900,N_9750,N_9764);
or U9901 (N_9901,N_9738,N_9772);
and U9902 (N_9902,N_9649,N_9619);
and U9903 (N_9903,N_9678,N_9778);
nor U9904 (N_9904,N_9735,N_9648);
and U9905 (N_9905,N_9762,N_9615);
and U9906 (N_9906,N_9699,N_9666);
or U9907 (N_9907,N_9648,N_9644);
nand U9908 (N_9908,N_9621,N_9607);
and U9909 (N_9909,N_9768,N_9643);
and U9910 (N_9910,N_9604,N_9728);
nand U9911 (N_9911,N_9791,N_9688);
or U9912 (N_9912,N_9622,N_9620);
nor U9913 (N_9913,N_9765,N_9777);
nand U9914 (N_9914,N_9704,N_9724);
nand U9915 (N_9915,N_9711,N_9662);
nand U9916 (N_9916,N_9775,N_9792);
and U9917 (N_9917,N_9780,N_9754);
and U9918 (N_9918,N_9701,N_9645);
or U9919 (N_9919,N_9691,N_9754);
nor U9920 (N_9920,N_9630,N_9792);
nand U9921 (N_9921,N_9695,N_9704);
and U9922 (N_9922,N_9749,N_9666);
or U9923 (N_9923,N_9735,N_9622);
and U9924 (N_9924,N_9670,N_9790);
nand U9925 (N_9925,N_9630,N_9720);
or U9926 (N_9926,N_9674,N_9667);
or U9927 (N_9927,N_9698,N_9683);
or U9928 (N_9928,N_9636,N_9708);
or U9929 (N_9929,N_9788,N_9630);
nand U9930 (N_9930,N_9634,N_9678);
or U9931 (N_9931,N_9751,N_9797);
nand U9932 (N_9932,N_9680,N_9791);
nor U9933 (N_9933,N_9646,N_9715);
or U9934 (N_9934,N_9711,N_9788);
and U9935 (N_9935,N_9606,N_9619);
nor U9936 (N_9936,N_9772,N_9638);
or U9937 (N_9937,N_9780,N_9750);
or U9938 (N_9938,N_9658,N_9653);
nand U9939 (N_9939,N_9647,N_9625);
nor U9940 (N_9940,N_9782,N_9698);
or U9941 (N_9941,N_9670,N_9663);
nand U9942 (N_9942,N_9751,N_9793);
nor U9943 (N_9943,N_9772,N_9712);
nand U9944 (N_9944,N_9761,N_9658);
or U9945 (N_9945,N_9633,N_9674);
nor U9946 (N_9946,N_9774,N_9713);
nor U9947 (N_9947,N_9715,N_9614);
or U9948 (N_9948,N_9636,N_9670);
and U9949 (N_9949,N_9775,N_9746);
and U9950 (N_9950,N_9719,N_9626);
nor U9951 (N_9951,N_9770,N_9767);
nor U9952 (N_9952,N_9626,N_9623);
nand U9953 (N_9953,N_9667,N_9698);
or U9954 (N_9954,N_9622,N_9784);
nand U9955 (N_9955,N_9675,N_9741);
or U9956 (N_9956,N_9795,N_9761);
nand U9957 (N_9957,N_9777,N_9723);
or U9958 (N_9958,N_9636,N_9760);
nor U9959 (N_9959,N_9789,N_9632);
nor U9960 (N_9960,N_9744,N_9766);
and U9961 (N_9961,N_9659,N_9769);
nand U9962 (N_9962,N_9780,N_9760);
and U9963 (N_9963,N_9606,N_9796);
nand U9964 (N_9964,N_9701,N_9612);
nor U9965 (N_9965,N_9778,N_9775);
or U9966 (N_9966,N_9763,N_9787);
or U9967 (N_9967,N_9681,N_9677);
or U9968 (N_9968,N_9671,N_9755);
nor U9969 (N_9969,N_9729,N_9789);
or U9970 (N_9970,N_9725,N_9685);
nand U9971 (N_9971,N_9619,N_9650);
nor U9972 (N_9972,N_9742,N_9774);
and U9973 (N_9973,N_9654,N_9649);
nor U9974 (N_9974,N_9607,N_9797);
nand U9975 (N_9975,N_9746,N_9714);
nor U9976 (N_9976,N_9799,N_9724);
nor U9977 (N_9977,N_9620,N_9774);
and U9978 (N_9978,N_9770,N_9748);
or U9979 (N_9979,N_9782,N_9690);
nor U9980 (N_9980,N_9737,N_9792);
nand U9981 (N_9981,N_9694,N_9722);
and U9982 (N_9982,N_9774,N_9788);
nor U9983 (N_9983,N_9777,N_9747);
nand U9984 (N_9984,N_9739,N_9799);
or U9985 (N_9985,N_9796,N_9685);
or U9986 (N_9986,N_9721,N_9738);
nand U9987 (N_9987,N_9729,N_9613);
nand U9988 (N_9988,N_9651,N_9618);
or U9989 (N_9989,N_9619,N_9786);
nor U9990 (N_9990,N_9732,N_9647);
nand U9991 (N_9991,N_9788,N_9772);
nand U9992 (N_9992,N_9654,N_9733);
or U9993 (N_9993,N_9657,N_9658);
nand U9994 (N_9994,N_9698,N_9663);
nor U9995 (N_9995,N_9716,N_9751);
and U9996 (N_9996,N_9685,N_9686);
or U9997 (N_9997,N_9724,N_9654);
nand U9998 (N_9998,N_9693,N_9605);
nor U9999 (N_9999,N_9668,N_9714);
nor U10000 (N_10000,N_9920,N_9893);
or U10001 (N_10001,N_9870,N_9801);
and U10002 (N_10002,N_9880,N_9950);
or U10003 (N_10003,N_9864,N_9899);
or U10004 (N_10004,N_9878,N_9811);
nand U10005 (N_10005,N_9934,N_9919);
or U10006 (N_10006,N_9925,N_9944);
nand U10007 (N_10007,N_9975,N_9904);
nor U10008 (N_10008,N_9986,N_9884);
and U10009 (N_10009,N_9957,N_9971);
nand U10010 (N_10010,N_9809,N_9976);
and U10011 (N_10011,N_9990,N_9860);
or U10012 (N_10012,N_9964,N_9928);
or U10013 (N_10013,N_9840,N_9933);
or U10014 (N_10014,N_9952,N_9824);
nand U10015 (N_10015,N_9865,N_9815);
nor U10016 (N_10016,N_9953,N_9965);
nor U10017 (N_10017,N_9841,N_9836);
or U10018 (N_10018,N_9888,N_9974);
and U10019 (N_10019,N_9803,N_9851);
and U10020 (N_10020,N_9983,N_9979);
or U10021 (N_10021,N_9854,N_9827);
or U10022 (N_10022,N_9821,N_9923);
and U10023 (N_10023,N_9882,N_9984);
and U10024 (N_10024,N_9962,N_9945);
nand U10025 (N_10025,N_9881,N_9946);
nor U10026 (N_10026,N_9829,N_9929);
or U10027 (N_10027,N_9875,N_9958);
and U10028 (N_10028,N_9856,N_9847);
or U10029 (N_10029,N_9995,N_9871);
and U10030 (N_10030,N_9895,N_9901);
or U10031 (N_10031,N_9850,N_9940);
or U10032 (N_10032,N_9802,N_9857);
or U10033 (N_10033,N_9885,N_9999);
nor U10034 (N_10034,N_9843,N_9973);
nand U10035 (N_10035,N_9879,N_9839);
and U10036 (N_10036,N_9900,N_9867);
nor U10037 (N_10037,N_9804,N_9921);
or U10038 (N_10038,N_9806,N_9993);
nand U10039 (N_10039,N_9833,N_9859);
or U10040 (N_10040,N_9931,N_9862);
nor U10041 (N_10041,N_9820,N_9902);
nor U10042 (N_10042,N_9826,N_9819);
and U10043 (N_10043,N_9936,N_9830);
nand U10044 (N_10044,N_9918,N_9810);
or U10045 (N_10045,N_9994,N_9996);
nand U10046 (N_10046,N_9991,N_9838);
nor U10047 (N_10047,N_9926,N_9968);
or U10048 (N_10048,N_9992,N_9892);
nand U10049 (N_10049,N_9861,N_9998);
or U10050 (N_10050,N_9906,N_9907);
and U10051 (N_10051,N_9914,N_9935);
nand U10052 (N_10052,N_9985,N_9825);
or U10053 (N_10053,N_9886,N_9989);
and U10054 (N_10054,N_9932,N_9938);
or U10055 (N_10055,N_9948,N_9890);
or U10056 (N_10056,N_9845,N_9942);
or U10057 (N_10057,N_9988,N_9831);
and U10058 (N_10058,N_9949,N_9908);
and U10059 (N_10059,N_9951,N_9987);
or U10060 (N_10060,N_9896,N_9818);
and U10061 (N_10061,N_9980,N_9954);
nand U10062 (N_10062,N_9910,N_9813);
and U10063 (N_10063,N_9972,N_9855);
and U10064 (N_10064,N_9828,N_9916);
nand U10065 (N_10065,N_9959,N_9963);
and U10066 (N_10066,N_9977,N_9808);
nand U10067 (N_10067,N_9853,N_9947);
nor U10068 (N_10068,N_9930,N_9911);
or U10069 (N_10069,N_9967,N_9842);
nor U10070 (N_10070,N_9816,N_9922);
and U10071 (N_10071,N_9939,N_9863);
nand U10072 (N_10072,N_9869,N_9978);
xor U10073 (N_10073,N_9898,N_9956);
nor U10074 (N_10074,N_9874,N_9858);
or U10075 (N_10075,N_9805,N_9917);
or U10076 (N_10076,N_9866,N_9981);
nand U10077 (N_10077,N_9837,N_9834);
nand U10078 (N_10078,N_9960,N_9844);
and U10079 (N_10079,N_9887,N_9846);
and U10080 (N_10080,N_9909,N_9852);
nor U10081 (N_10081,N_9848,N_9894);
and U10082 (N_10082,N_9903,N_9961);
or U10083 (N_10083,N_9924,N_9889);
and U10084 (N_10084,N_9868,N_9969);
nand U10085 (N_10085,N_9822,N_9877);
nand U10086 (N_10086,N_9913,N_9812);
and U10087 (N_10087,N_9915,N_9997);
and U10088 (N_10088,N_9873,N_9817);
or U10089 (N_10089,N_9835,N_9832);
or U10090 (N_10090,N_9800,N_9883);
nand U10091 (N_10091,N_9876,N_9982);
nand U10092 (N_10092,N_9966,N_9937);
or U10093 (N_10093,N_9891,N_9943);
nor U10094 (N_10094,N_9814,N_9872);
nor U10095 (N_10095,N_9955,N_9905);
nand U10096 (N_10096,N_9897,N_9823);
nor U10097 (N_10097,N_9807,N_9941);
and U10098 (N_10098,N_9912,N_9927);
or U10099 (N_10099,N_9970,N_9849);
or U10100 (N_10100,N_9862,N_9868);
nor U10101 (N_10101,N_9804,N_9855);
xnor U10102 (N_10102,N_9805,N_9958);
nor U10103 (N_10103,N_9816,N_9915);
nor U10104 (N_10104,N_9916,N_9800);
or U10105 (N_10105,N_9995,N_9907);
nor U10106 (N_10106,N_9888,N_9959);
or U10107 (N_10107,N_9953,N_9862);
nand U10108 (N_10108,N_9964,N_9847);
and U10109 (N_10109,N_9810,N_9851);
nand U10110 (N_10110,N_9851,N_9958);
or U10111 (N_10111,N_9908,N_9974);
and U10112 (N_10112,N_9865,N_9809);
nor U10113 (N_10113,N_9996,N_9888);
nor U10114 (N_10114,N_9878,N_9992);
or U10115 (N_10115,N_9994,N_9960);
xnor U10116 (N_10116,N_9853,N_9997);
or U10117 (N_10117,N_9924,N_9805);
nand U10118 (N_10118,N_9901,N_9939);
nand U10119 (N_10119,N_9838,N_9873);
nor U10120 (N_10120,N_9969,N_9859);
nand U10121 (N_10121,N_9833,N_9921);
or U10122 (N_10122,N_9866,N_9898);
or U10123 (N_10123,N_9862,N_9870);
nor U10124 (N_10124,N_9822,N_9874);
or U10125 (N_10125,N_9948,N_9923);
nor U10126 (N_10126,N_9942,N_9872);
or U10127 (N_10127,N_9915,N_9957);
or U10128 (N_10128,N_9816,N_9805);
nand U10129 (N_10129,N_9950,N_9896);
or U10130 (N_10130,N_9894,N_9936);
nand U10131 (N_10131,N_9905,N_9923);
or U10132 (N_10132,N_9970,N_9997);
and U10133 (N_10133,N_9989,N_9939);
nor U10134 (N_10134,N_9922,N_9863);
nor U10135 (N_10135,N_9866,N_9998);
or U10136 (N_10136,N_9899,N_9949);
nor U10137 (N_10137,N_9970,N_9936);
nand U10138 (N_10138,N_9955,N_9846);
nor U10139 (N_10139,N_9902,N_9807);
nand U10140 (N_10140,N_9973,N_9933);
nand U10141 (N_10141,N_9846,N_9863);
or U10142 (N_10142,N_9893,N_9958);
nand U10143 (N_10143,N_9975,N_9984);
or U10144 (N_10144,N_9891,N_9983);
and U10145 (N_10145,N_9892,N_9956);
nor U10146 (N_10146,N_9891,N_9940);
and U10147 (N_10147,N_9885,N_9837);
and U10148 (N_10148,N_9800,N_9845);
nor U10149 (N_10149,N_9860,N_9875);
nand U10150 (N_10150,N_9983,N_9857);
nor U10151 (N_10151,N_9963,N_9802);
or U10152 (N_10152,N_9837,N_9983);
nor U10153 (N_10153,N_9955,N_9950);
nand U10154 (N_10154,N_9831,N_9811);
nor U10155 (N_10155,N_9812,N_9857);
or U10156 (N_10156,N_9921,N_9882);
nor U10157 (N_10157,N_9929,N_9865);
or U10158 (N_10158,N_9857,N_9891);
or U10159 (N_10159,N_9995,N_9997);
or U10160 (N_10160,N_9805,N_9822);
or U10161 (N_10161,N_9859,N_9958);
and U10162 (N_10162,N_9872,N_9938);
nor U10163 (N_10163,N_9892,N_9809);
nor U10164 (N_10164,N_9862,N_9905);
nand U10165 (N_10165,N_9978,N_9970);
or U10166 (N_10166,N_9981,N_9915);
and U10167 (N_10167,N_9919,N_9954);
and U10168 (N_10168,N_9962,N_9916);
or U10169 (N_10169,N_9929,N_9880);
or U10170 (N_10170,N_9915,N_9958);
nand U10171 (N_10171,N_9953,N_9853);
and U10172 (N_10172,N_9901,N_9801);
nor U10173 (N_10173,N_9824,N_9808);
and U10174 (N_10174,N_9923,N_9882);
or U10175 (N_10175,N_9980,N_9993);
and U10176 (N_10176,N_9814,N_9898);
and U10177 (N_10177,N_9912,N_9816);
and U10178 (N_10178,N_9915,N_9909);
or U10179 (N_10179,N_9916,N_9992);
or U10180 (N_10180,N_9939,N_9802);
nand U10181 (N_10181,N_9916,N_9968);
and U10182 (N_10182,N_9884,N_9873);
and U10183 (N_10183,N_9852,N_9992);
or U10184 (N_10184,N_9960,N_9939);
nor U10185 (N_10185,N_9935,N_9903);
nor U10186 (N_10186,N_9955,N_9958);
or U10187 (N_10187,N_9941,N_9822);
nand U10188 (N_10188,N_9952,N_9916);
or U10189 (N_10189,N_9890,N_9815);
or U10190 (N_10190,N_9959,N_9869);
nand U10191 (N_10191,N_9860,N_9809);
nand U10192 (N_10192,N_9940,N_9935);
or U10193 (N_10193,N_9818,N_9801);
and U10194 (N_10194,N_9838,N_9953);
nor U10195 (N_10195,N_9988,N_9868);
or U10196 (N_10196,N_9808,N_9876);
and U10197 (N_10197,N_9861,N_9910);
and U10198 (N_10198,N_9815,N_9817);
nand U10199 (N_10199,N_9966,N_9818);
nand U10200 (N_10200,N_10040,N_10077);
nor U10201 (N_10201,N_10094,N_10047);
and U10202 (N_10202,N_10139,N_10191);
and U10203 (N_10203,N_10142,N_10025);
or U10204 (N_10204,N_10118,N_10081);
nand U10205 (N_10205,N_10003,N_10024);
nor U10206 (N_10206,N_10145,N_10074);
nor U10207 (N_10207,N_10057,N_10158);
and U10208 (N_10208,N_10138,N_10190);
nand U10209 (N_10209,N_10110,N_10187);
nor U10210 (N_10210,N_10133,N_10028);
and U10211 (N_10211,N_10186,N_10175);
or U10212 (N_10212,N_10056,N_10012);
nand U10213 (N_10213,N_10103,N_10100);
and U10214 (N_10214,N_10073,N_10184);
nand U10215 (N_10215,N_10123,N_10048);
and U10216 (N_10216,N_10041,N_10078);
and U10217 (N_10217,N_10196,N_10069);
nand U10218 (N_10218,N_10082,N_10031);
and U10219 (N_10219,N_10049,N_10044);
nand U10220 (N_10220,N_10091,N_10146);
and U10221 (N_10221,N_10068,N_10092);
nand U10222 (N_10222,N_10052,N_10021);
or U10223 (N_10223,N_10086,N_10119);
and U10224 (N_10224,N_10071,N_10065);
nor U10225 (N_10225,N_10037,N_10181);
or U10226 (N_10226,N_10140,N_10015);
and U10227 (N_10227,N_10029,N_10008);
nor U10228 (N_10228,N_10155,N_10107);
or U10229 (N_10229,N_10087,N_10157);
and U10230 (N_10230,N_10173,N_10160);
nor U10231 (N_10231,N_10050,N_10112);
nand U10232 (N_10232,N_10114,N_10095);
or U10233 (N_10233,N_10055,N_10034);
nand U10234 (N_10234,N_10166,N_10013);
nand U10235 (N_10235,N_10168,N_10000);
and U10236 (N_10236,N_10002,N_10135);
and U10237 (N_10237,N_10122,N_10197);
or U10238 (N_10238,N_10007,N_10098);
and U10239 (N_10239,N_10062,N_10060);
nor U10240 (N_10240,N_10179,N_10177);
nand U10241 (N_10241,N_10009,N_10120);
or U10242 (N_10242,N_10035,N_10001);
or U10243 (N_10243,N_10165,N_10144);
and U10244 (N_10244,N_10017,N_10032);
nor U10245 (N_10245,N_10020,N_10115);
nor U10246 (N_10246,N_10036,N_10083);
or U10247 (N_10247,N_10075,N_10054);
and U10248 (N_10248,N_10059,N_10051);
and U10249 (N_10249,N_10180,N_10006);
and U10250 (N_10250,N_10038,N_10163);
or U10251 (N_10251,N_10010,N_10005);
nor U10252 (N_10252,N_10080,N_10189);
nor U10253 (N_10253,N_10104,N_10113);
nor U10254 (N_10254,N_10164,N_10064);
and U10255 (N_10255,N_10088,N_10063);
nand U10256 (N_10256,N_10131,N_10170);
nand U10257 (N_10257,N_10148,N_10090);
or U10258 (N_10258,N_10195,N_10079);
or U10259 (N_10259,N_10162,N_10117);
or U10260 (N_10260,N_10085,N_10106);
nand U10261 (N_10261,N_10102,N_10198);
and U10262 (N_10262,N_10188,N_10101);
nand U10263 (N_10263,N_10169,N_10150);
nand U10264 (N_10264,N_10105,N_10194);
and U10265 (N_10265,N_10137,N_10124);
nor U10266 (N_10266,N_10152,N_10159);
nor U10267 (N_10267,N_10066,N_10116);
nand U10268 (N_10268,N_10171,N_10134);
and U10269 (N_10269,N_10072,N_10033);
nor U10270 (N_10270,N_10185,N_10027);
nor U10271 (N_10271,N_10046,N_10111);
nor U10272 (N_10272,N_10149,N_10174);
or U10273 (N_10273,N_10127,N_10128);
nand U10274 (N_10274,N_10023,N_10070);
nand U10275 (N_10275,N_10121,N_10076);
nand U10276 (N_10276,N_10161,N_10192);
or U10277 (N_10277,N_10147,N_10130);
or U10278 (N_10278,N_10058,N_10132);
or U10279 (N_10279,N_10199,N_10026);
or U10280 (N_10280,N_10061,N_10156);
nor U10281 (N_10281,N_10016,N_10022);
nand U10282 (N_10282,N_10045,N_10178);
nor U10283 (N_10283,N_10182,N_10176);
nor U10284 (N_10284,N_10039,N_10004);
and U10285 (N_10285,N_10154,N_10011);
and U10286 (N_10286,N_10172,N_10109);
nand U10287 (N_10287,N_10042,N_10141);
nor U10288 (N_10288,N_10136,N_10099);
and U10289 (N_10289,N_10193,N_10043);
and U10290 (N_10290,N_10129,N_10151);
nor U10291 (N_10291,N_10019,N_10097);
or U10292 (N_10292,N_10030,N_10067);
nand U10293 (N_10293,N_10018,N_10096);
nor U10294 (N_10294,N_10014,N_10153);
and U10295 (N_10295,N_10053,N_10093);
nor U10296 (N_10296,N_10108,N_10125);
or U10297 (N_10297,N_10167,N_10143);
nand U10298 (N_10298,N_10183,N_10126);
nor U10299 (N_10299,N_10089,N_10084);
nor U10300 (N_10300,N_10157,N_10103);
nor U10301 (N_10301,N_10191,N_10144);
and U10302 (N_10302,N_10029,N_10156);
or U10303 (N_10303,N_10089,N_10137);
nand U10304 (N_10304,N_10078,N_10106);
or U10305 (N_10305,N_10156,N_10006);
nor U10306 (N_10306,N_10167,N_10184);
or U10307 (N_10307,N_10079,N_10107);
nor U10308 (N_10308,N_10155,N_10066);
nor U10309 (N_10309,N_10058,N_10064);
and U10310 (N_10310,N_10196,N_10115);
nor U10311 (N_10311,N_10103,N_10083);
or U10312 (N_10312,N_10086,N_10165);
nor U10313 (N_10313,N_10141,N_10061);
and U10314 (N_10314,N_10013,N_10126);
or U10315 (N_10315,N_10078,N_10149);
and U10316 (N_10316,N_10197,N_10172);
nor U10317 (N_10317,N_10008,N_10091);
nand U10318 (N_10318,N_10160,N_10132);
nand U10319 (N_10319,N_10069,N_10064);
nand U10320 (N_10320,N_10148,N_10169);
nor U10321 (N_10321,N_10167,N_10082);
and U10322 (N_10322,N_10061,N_10031);
or U10323 (N_10323,N_10195,N_10186);
nor U10324 (N_10324,N_10089,N_10010);
nor U10325 (N_10325,N_10069,N_10001);
and U10326 (N_10326,N_10104,N_10055);
nand U10327 (N_10327,N_10085,N_10097);
and U10328 (N_10328,N_10129,N_10004);
nand U10329 (N_10329,N_10003,N_10164);
and U10330 (N_10330,N_10010,N_10062);
nand U10331 (N_10331,N_10120,N_10135);
and U10332 (N_10332,N_10110,N_10071);
and U10333 (N_10333,N_10141,N_10129);
nand U10334 (N_10334,N_10135,N_10191);
nor U10335 (N_10335,N_10044,N_10125);
and U10336 (N_10336,N_10186,N_10012);
and U10337 (N_10337,N_10042,N_10075);
nand U10338 (N_10338,N_10187,N_10013);
nor U10339 (N_10339,N_10134,N_10027);
nor U10340 (N_10340,N_10165,N_10188);
or U10341 (N_10341,N_10078,N_10094);
nand U10342 (N_10342,N_10161,N_10165);
nand U10343 (N_10343,N_10094,N_10004);
nor U10344 (N_10344,N_10037,N_10116);
nor U10345 (N_10345,N_10181,N_10108);
nand U10346 (N_10346,N_10142,N_10118);
nand U10347 (N_10347,N_10074,N_10177);
and U10348 (N_10348,N_10040,N_10198);
nand U10349 (N_10349,N_10070,N_10170);
and U10350 (N_10350,N_10093,N_10158);
and U10351 (N_10351,N_10066,N_10196);
and U10352 (N_10352,N_10156,N_10135);
nor U10353 (N_10353,N_10008,N_10009);
nand U10354 (N_10354,N_10129,N_10191);
or U10355 (N_10355,N_10194,N_10142);
nand U10356 (N_10356,N_10009,N_10014);
nand U10357 (N_10357,N_10127,N_10169);
nor U10358 (N_10358,N_10154,N_10057);
or U10359 (N_10359,N_10011,N_10148);
and U10360 (N_10360,N_10007,N_10162);
nor U10361 (N_10361,N_10139,N_10065);
nor U10362 (N_10362,N_10092,N_10144);
nor U10363 (N_10363,N_10166,N_10073);
and U10364 (N_10364,N_10123,N_10190);
nor U10365 (N_10365,N_10152,N_10103);
and U10366 (N_10366,N_10143,N_10158);
and U10367 (N_10367,N_10032,N_10053);
or U10368 (N_10368,N_10125,N_10175);
nor U10369 (N_10369,N_10096,N_10161);
and U10370 (N_10370,N_10198,N_10005);
or U10371 (N_10371,N_10124,N_10054);
nor U10372 (N_10372,N_10050,N_10141);
and U10373 (N_10373,N_10165,N_10049);
or U10374 (N_10374,N_10057,N_10032);
nor U10375 (N_10375,N_10014,N_10102);
and U10376 (N_10376,N_10151,N_10093);
nand U10377 (N_10377,N_10023,N_10061);
nand U10378 (N_10378,N_10002,N_10037);
nor U10379 (N_10379,N_10094,N_10031);
nor U10380 (N_10380,N_10060,N_10001);
xor U10381 (N_10381,N_10097,N_10023);
nor U10382 (N_10382,N_10027,N_10004);
and U10383 (N_10383,N_10147,N_10102);
and U10384 (N_10384,N_10168,N_10048);
and U10385 (N_10385,N_10190,N_10137);
nor U10386 (N_10386,N_10124,N_10149);
and U10387 (N_10387,N_10122,N_10084);
or U10388 (N_10388,N_10086,N_10046);
or U10389 (N_10389,N_10041,N_10186);
or U10390 (N_10390,N_10056,N_10117);
and U10391 (N_10391,N_10090,N_10124);
or U10392 (N_10392,N_10055,N_10153);
and U10393 (N_10393,N_10010,N_10058);
and U10394 (N_10394,N_10165,N_10089);
nor U10395 (N_10395,N_10157,N_10067);
and U10396 (N_10396,N_10185,N_10104);
and U10397 (N_10397,N_10189,N_10170);
nand U10398 (N_10398,N_10012,N_10174);
nor U10399 (N_10399,N_10123,N_10080);
or U10400 (N_10400,N_10288,N_10338);
nor U10401 (N_10401,N_10390,N_10282);
nor U10402 (N_10402,N_10235,N_10203);
nand U10403 (N_10403,N_10334,N_10398);
or U10404 (N_10404,N_10388,N_10290);
nand U10405 (N_10405,N_10232,N_10377);
nand U10406 (N_10406,N_10253,N_10245);
nor U10407 (N_10407,N_10254,N_10383);
and U10408 (N_10408,N_10387,N_10226);
and U10409 (N_10409,N_10242,N_10228);
and U10410 (N_10410,N_10375,N_10366);
nand U10411 (N_10411,N_10259,N_10295);
and U10412 (N_10412,N_10372,N_10252);
nand U10413 (N_10413,N_10393,N_10329);
and U10414 (N_10414,N_10307,N_10371);
or U10415 (N_10415,N_10362,N_10359);
nor U10416 (N_10416,N_10279,N_10317);
nor U10417 (N_10417,N_10328,N_10268);
nand U10418 (N_10418,N_10283,N_10353);
or U10419 (N_10419,N_10357,N_10231);
and U10420 (N_10420,N_10222,N_10323);
and U10421 (N_10421,N_10369,N_10325);
nor U10422 (N_10422,N_10356,N_10297);
or U10423 (N_10423,N_10292,N_10301);
nor U10424 (N_10424,N_10233,N_10237);
nor U10425 (N_10425,N_10281,N_10251);
nand U10426 (N_10426,N_10376,N_10221);
nand U10427 (N_10427,N_10285,N_10343);
nor U10428 (N_10428,N_10315,N_10225);
and U10429 (N_10429,N_10223,N_10263);
and U10430 (N_10430,N_10379,N_10370);
or U10431 (N_10431,N_10274,N_10354);
nor U10432 (N_10432,N_10286,N_10346);
and U10433 (N_10433,N_10219,N_10305);
and U10434 (N_10434,N_10358,N_10244);
nor U10435 (N_10435,N_10255,N_10350);
and U10436 (N_10436,N_10342,N_10257);
and U10437 (N_10437,N_10275,N_10368);
nand U10438 (N_10438,N_10215,N_10316);
or U10439 (N_10439,N_10239,N_10310);
or U10440 (N_10440,N_10332,N_10363);
nand U10441 (N_10441,N_10336,N_10318);
nor U10442 (N_10442,N_10200,N_10355);
or U10443 (N_10443,N_10384,N_10381);
or U10444 (N_10444,N_10210,N_10211);
nand U10445 (N_10445,N_10280,N_10227);
and U10446 (N_10446,N_10392,N_10367);
or U10447 (N_10447,N_10265,N_10208);
and U10448 (N_10448,N_10333,N_10380);
and U10449 (N_10449,N_10272,N_10246);
and U10450 (N_10450,N_10269,N_10287);
nor U10451 (N_10451,N_10261,N_10296);
or U10452 (N_10452,N_10293,N_10320);
or U10453 (N_10453,N_10243,N_10205);
nor U10454 (N_10454,N_10224,N_10230);
nor U10455 (N_10455,N_10277,N_10399);
nor U10456 (N_10456,N_10212,N_10351);
nor U10457 (N_10457,N_10308,N_10340);
nor U10458 (N_10458,N_10335,N_10213);
nand U10459 (N_10459,N_10349,N_10247);
or U10460 (N_10460,N_10266,N_10256);
or U10461 (N_10461,N_10339,N_10322);
or U10462 (N_10462,N_10396,N_10229);
and U10463 (N_10463,N_10391,N_10386);
nand U10464 (N_10464,N_10300,N_10344);
nand U10465 (N_10465,N_10278,N_10394);
nand U10466 (N_10466,N_10291,N_10250);
nand U10467 (N_10467,N_10309,N_10321);
nor U10468 (N_10468,N_10313,N_10330);
and U10469 (N_10469,N_10382,N_10214);
or U10470 (N_10470,N_10352,N_10209);
and U10471 (N_10471,N_10206,N_10289);
or U10472 (N_10472,N_10267,N_10238);
nor U10473 (N_10473,N_10364,N_10324);
and U10474 (N_10474,N_10236,N_10299);
nand U10475 (N_10475,N_10395,N_10312);
nand U10476 (N_10476,N_10326,N_10258);
and U10477 (N_10477,N_10202,N_10216);
and U10478 (N_10478,N_10234,N_10306);
or U10479 (N_10479,N_10378,N_10389);
nor U10480 (N_10480,N_10302,N_10341);
nor U10481 (N_10481,N_10271,N_10262);
xor U10482 (N_10482,N_10373,N_10348);
nand U10483 (N_10483,N_10304,N_10374);
nand U10484 (N_10484,N_10270,N_10201);
nor U10485 (N_10485,N_10217,N_10260);
or U10486 (N_10486,N_10207,N_10249);
and U10487 (N_10487,N_10319,N_10311);
and U10488 (N_10488,N_10264,N_10220);
or U10489 (N_10489,N_10337,N_10347);
or U10490 (N_10490,N_10294,N_10365);
nor U10491 (N_10491,N_10273,N_10314);
and U10492 (N_10492,N_10204,N_10397);
nand U10493 (N_10493,N_10240,N_10298);
and U10494 (N_10494,N_10327,N_10248);
nor U10495 (N_10495,N_10241,N_10385);
nor U10496 (N_10496,N_10284,N_10276);
nor U10497 (N_10497,N_10360,N_10345);
nor U10498 (N_10498,N_10331,N_10218);
nand U10499 (N_10499,N_10303,N_10361);
and U10500 (N_10500,N_10396,N_10205);
and U10501 (N_10501,N_10254,N_10321);
or U10502 (N_10502,N_10305,N_10204);
nand U10503 (N_10503,N_10384,N_10390);
nand U10504 (N_10504,N_10328,N_10279);
and U10505 (N_10505,N_10275,N_10366);
nand U10506 (N_10506,N_10293,N_10394);
xor U10507 (N_10507,N_10311,N_10346);
nor U10508 (N_10508,N_10331,N_10268);
and U10509 (N_10509,N_10383,N_10329);
nand U10510 (N_10510,N_10375,N_10311);
or U10511 (N_10511,N_10246,N_10236);
nand U10512 (N_10512,N_10381,N_10201);
nand U10513 (N_10513,N_10385,N_10376);
nor U10514 (N_10514,N_10341,N_10319);
nor U10515 (N_10515,N_10335,N_10268);
or U10516 (N_10516,N_10227,N_10373);
nor U10517 (N_10517,N_10350,N_10386);
nand U10518 (N_10518,N_10324,N_10264);
nor U10519 (N_10519,N_10247,N_10285);
and U10520 (N_10520,N_10328,N_10311);
nor U10521 (N_10521,N_10280,N_10213);
or U10522 (N_10522,N_10202,N_10212);
or U10523 (N_10523,N_10340,N_10311);
or U10524 (N_10524,N_10321,N_10354);
nor U10525 (N_10525,N_10352,N_10371);
nor U10526 (N_10526,N_10279,N_10397);
or U10527 (N_10527,N_10214,N_10241);
or U10528 (N_10528,N_10286,N_10383);
nor U10529 (N_10529,N_10323,N_10281);
and U10530 (N_10530,N_10206,N_10261);
nor U10531 (N_10531,N_10333,N_10288);
nand U10532 (N_10532,N_10351,N_10300);
or U10533 (N_10533,N_10202,N_10382);
nor U10534 (N_10534,N_10335,N_10276);
and U10535 (N_10535,N_10372,N_10258);
or U10536 (N_10536,N_10356,N_10239);
or U10537 (N_10537,N_10336,N_10328);
or U10538 (N_10538,N_10256,N_10390);
and U10539 (N_10539,N_10360,N_10221);
nand U10540 (N_10540,N_10282,N_10249);
or U10541 (N_10541,N_10242,N_10262);
or U10542 (N_10542,N_10327,N_10233);
and U10543 (N_10543,N_10381,N_10222);
or U10544 (N_10544,N_10200,N_10374);
nor U10545 (N_10545,N_10377,N_10230);
nor U10546 (N_10546,N_10279,N_10314);
or U10547 (N_10547,N_10203,N_10350);
nand U10548 (N_10548,N_10380,N_10262);
nand U10549 (N_10549,N_10262,N_10227);
and U10550 (N_10550,N_10278,N_10297);
and U10551 (N_10551,N_10256,N_10254);
nand U10552 (N_10552,N_10233,N_10220);
nor U10553 (N_10553,N_10340,N_10366);
nand U10554 (N_10554,N_10365,N_10349);
nor U10555 (N_10555,N_10219,N_10323);
and U10556 (N_10556,N_10317,N_10230);
and U10557 (N_10557,N_10273,N_10369);
nor U10558 (N_10558,N_10330,N_10326);
and U10559 (N_10559,N_10259,N_10345);
and U10560 (N_10560,N_10272,N_10319);
xor U10561 (N_10561,N_10344,N_10386);
nor U10562 (N_10562,N_10343,N_10367);
nor U10563 (N_10563,N_10310,N_10232);
nand U10564 (N_10564,N_10292,N_10352);
and U10565 (N_10565,N_10334,N_10289);
nor U10566 (N_10566,N_10202,N_10299);
nand U10567 (N_10567,N_10261,N_10259);
nand U10568 (N_10568,N_10387,N_10275);
and U10569 (N_10569,N_10373,N_10293);
and U10570 (N_10570,N_10348,N_10387);
and U10571 (N_10571,N_10263,N_10353);
or U10572 (N_10572,N_10283,N_10211);
nand U10573 (N_10573,N_10204,N_10213);
or U10574 (N_10574,N_10301,N_10350);
or U10575 (N_10575,N_10260,N_10238);
nand U10576 (N_10576,N_10215,N_10253);
and U10577 (N_10577,N_10273,N_10239);
nor U10578 (N_10578,N_10314,N_10350);
or U10579 (N_10579,N_10217,N_10279);
nand U10580 (N_10580,N_10323,N_10292);
nand U10581 (N_10581,N_10287,N_10350);
nor U10582 (N_10582,N_10392,N_10385);
or U10583 (N_10583,N_10370,N_10378);
and U10584 (N_10584,N_10217,N_10296);
and U10585 (N_10585,N_10262,N_10269);
and U10586 (N_10586,N_10224,N_10376);
or U10587 (N_10587,N_10376,N_10205);
nand U10588 (N_10588,N_10306,N_10314);
nor U10589 (N_10589,N_10274,N_10371);
and U10590 (N_10590,N_10372,N_10211);
or U10591 (N_10591,N_10228,N_10201);
nor U10592 (N_10592,N_10397,N_10222);
nand U10593 (N_10593,N_10294,N_10383);
and U10594 (N_10594,N_10369,N_10230);
or U10595 (N_10595,N_10355,N_10317);
nand U10596 (N_10596,N_10352,N_10357);
nor U10597 (N_10597,N_10243,N_10354);
or U10598 (N_10598,N_10377,N_10371);
and U10599 (N_10599,N_10211,N_10254);
nor U10600 (N_10600,N_10515,N_10407);
nor U10601 (N_10601,N_10536,N_10502);
nand U10602 (N_10602,N_10518,N_10447);
nand U10603 (N_10603,N_10471,N_10492);
nand U10604 (N_10604,N_10481,N_10423);
nand U10605 (N_10605,N_10563,N_10528);
nor U10606 (N_10606,N_10504,N_10573);
nand U10607 (N_10607,N_10433,N_10538);
or U10608 (N_10608,N_10400,N_10449);
nand U10609 (N_10609,N_10559,N_10495);
nor U10610 (N_10610,N_10470,N_10439);
and U10611 (N_10611,N_10417,N_10461);
and U10612 (N_10612,N_10462,N_10452);
nand U10613 (N_10613,N_10507,N_10485);
and U10614 (N_10614,N_10429,N_10413);
and U10615 (N_10615,N_10503,N_10565);
or U10616 (N_10616,N_10476,N_10488);
nor U10617 (N_10617,N_10522,N_10438);
nor U10618 (N_10618,N_10500,N_10548);
nor U10619 (N_10619,N_10555,N_10463);
and U10620 (N_10620,N_10520,N_10435);
nor U10621 (N_10621,N_10570,N_10456);
and U10622 (N_10622,N_10594,N_10531);
and U10623 (N_10623,N_10479,N_10458);
nand U10624 (N_10624,N_10491,N_10455);
nand U10625 (N_10625,N_10525,N_10547);
and U10626 (N_10626,N_10478,N_10450);
and U10627 (N_10627,N_10501,N_10475);
or U10628 (N_10628,N_10505,N_10446);
nand U10629 (N_10629,N_10402,N_10483);
and U10630 (N_10630,N_10514,N_10541);
nand U10631 (N_10631,N_10437,N_10572);
nor U10632 (N_10632,N_10568,N_10482);
nor U10633 (N_10633,N_10408,N_10409);
nor U10634 (N_10634,N_10587,N_10445);
or U10635 (N_10635,N_10578,N_10591);
or U10636 (N_10636,N_10421,N_10532);
nand U10637 (N_10637,N_10596,N_10526);
nor U10638 (N_10638,N_10549,N_10472);
and U10639 (N_10639,N_10403,N_10410);
nor U10640 (N_10640,N_10561,N_10582);
nor U10641 (N_10641,N_10506,N_10422);
and U10642 (N_10642,N_10551,N_10477);
nand U10643 (N_10643,N_10431,N_10566);
nor U10644 (N_10644,N_10489,N_10552);
nor U10645 (N_10645,N_10508,N_10599);
nand U10646 (N_10646,N_10484,N_10442);
nand U10647 (N_10647,N_10537,N_10467);
nand U10648 (N_10648,N_10436,N_10516);
nor U10649 (N_10649,N_10590,N_10598);
or U10650 (N_10650,N_10546,N_10564);
and U10651 (N_10651,N_10513,N_10441);
nor U10652 (N_10652,N_10579,N_10576);
or U10653 (N_10653,N_10597,N_10524);
nor U10654 (N_10654,N_10530,N_10490);
xor U10655 (N_10655,N_10440,N_10404);
nand U10656 (N_10656,N_10499,N_10560);
nor U10657 (N_10657,N_10406,N_10527);
and U10658 (N_10658,N_10412,N_10593);
nor U10659 (N_10659,N_10535,N_10567);
nor U10660 (N_10660,N_10543,N_10468);
and U10661 (N_10661,N_10512,N_10496);
nor U10662 (N_10662,N_10592,N_10554);
nor U10663 (N_10663,N_10511,N_10428);
nor U10664 (N_10664,N_10517,N_10588);
nand U10665 (N_10665,N_10464,N_10448);
nand U10666 (N_10666,N_10562,N_10411);
nor U10667 (N_10667,N_10589,N_10533);
or U10668 (N_10668,N_10498,N_10584);
nor U10669 (N_10669,N_10473,N_10466);
nand U10670 (N_10670,N_10443,N_10469);
nor U10671 (N_10671,N_10540,N_10427);
and U10672 (N_10672,N_10557,N_10414);
nor U10673 (N_10673,N_10486,N_10558);
and U10674 (N_10674,N_10577,N_10453);
nand U10675 (N_10675,N_10424,N_10460);
nor U10676 (N_10676,N_10542,N_10419);
nor U10677 (N_10677,N_10426,N_10425);
or U10678 (N_10678,N_10509,N_10474);
nand U10679 (N_10679,N_10401,N_10529);
and U10680 (N_10680,N_10432,N_10521);
nand U10681 (N_10681,N_10444,N_10569);
and U10682 (N_10682,N_10556,N_10583);
nor U10683 (N_10683,N_10415,N_10497);
nor U10684 (N_10684,N_10571,N_10534);
nand U10685 (N_10685,N_10480,N_10459);
nor U10686 (N_10686,N_10493,N_10595);
or U10687 (N_10687,N_10545,N_10420);
or U10688 (N_10688,N_10451,N_10430);
or U10689 (N_10689,N_10550,N_10580);
nor U10690 (N_10690,N_10544,N_10434);
nor U10691 (N_10691,N_10510,N_10585);
or U10692 (N_10692,N_10574,N_10519);
nor U10693 (N_10693,N_10487,N_10405);
and U10694 (N_10694,N_10575,N_10581);
or U10695 (N_10695,N_10586,N_10494);
and U10696 (N_10696,N_10539,N_10416);
or U10697 (N_10697,N_10523,N_10457);
nand U10698 (N_10698,N_10418,N_10454);
nand U10699 (N_10699,N_10553,N_10465);
nand U10700 (N_10700,N_10423,N_10524);
xor U10701 (N_10701,N_10536,N_10599);
nor U10702 (N_10702,N_10421,N_10510);
nor U10703 (N_10703,N_10444,N_10558);
nand U10704 (N_10704,N_10471,N_10417);
nand U10705 (N_10705,N_10596,N_10434);
or U10706 (N_10706,N_10570,N_10563);
nand U10707 (N_10707,N_10495,N_10586);
and U10708 (N_10708,N_10533,N_10451);
or U10709 (N_10709,N_10458,N_10589);
nand U10710 (N_10710,N_10599,N_10570);
nand U10711 (N_10711,N_10450,N_10518);
nor U10712 (N_10712,N_10560,N_10520);
nor U10713 (N_10713,N_10412,N_10426);
and U10714 (N_10714,N_10431,N_10437);
nor U10715 (N_10715,N_10594,N_10555);
and U10716 (N_10716,N_10546,N_10480);
nand U10717 (N_10717,N_10541,N_10425);
nor U10718 (N_10718,N_10555,N_10592);
or U10719 (N_10719,N_10557,N_10515);
nand U10720 (N_10720,N_10495,N_10524);
nand U10721 (N_10721,N_10554,N_10555);
nand U10722 (N_10722,N_10530,N_10463);
and U10723 (N_10723,N_10424,N_10422);
or U10724 (N_10724,N_10400,N_10453);
or U10725 (N_10725,N_10515,N_10456);
and U10726 (N_10726,N_10450,N_10401);
nor U10727 (N_10727,N_10573,N_10482);
nand U10728 (N_10728,N_10523,N_10553);
and U10729 (N_10729,N_10557,N_10451);
or U10730 (N_10730,N_10597,N_10483);
or U10731 (N_10731,N_10421,N_10520);
nor U10732 (N_10732,N_10587,N_10588);
nor U10733 (N_10733,N_10417,N_10418);
nor U10734 (N_10734,N_10564,N_10430);
and U10735 (N_10735,N_10518,N_10493);
and U10736 (N_10736,N_10461,N_10471);
or U10737 (N_10737,N_10435,N_10405);
or U10738 (N_10738,N_10412,N_10565);
nand U10739 (N_10739,N_10421,N_10443);
nand U10740 (N_10740,N_10477,N_10401);
nand U10741 (N_10741,N_10595,N_10567);
nand U10742 (N_10742,N_10426,N_10455);
nor U10743 (N_10743,N_10550,N_10555);
and U10744 (N_10744,N_10585,N_10576);
nor U10745 (N_10745,N_10445,N_10497);
nor U10746 (N_10746,N_10515,N_10577);
nand U10747 (N_10747,N_10426,N_10591);
or U10748 (N_10748,N_10455,N_10555);
nand U10749 (N_10749,N_10568,N_10545);
and U10750 (N_10750,N_10532,N_10485);
nand U10751 (N_10751,N_10407,N_10441);
or U10752 (N_10752,N_10447,N_10427);
and U10753 (N_10753,N_10557,N_10508);
nor U10754 (N_10754,N_10430,N_10557);
nor U10755 (N_10755,N_10461,N_10550);
nand U10756 (N_10756,N_10408,N_10548);
and U10757 (N_10757,N_10425,N_10583);
nand U10758 (N_10758,N_10586,N_10588);
nor U10759 (N_10759,N_10539,N_10573);
or U10760 (N_10760,N_10427,N_10551);
nor U10761 (N_10761,N_10534,N_10597);
and U10762 (N_10762,N_10577,N_10531);
nand U10763 (N_10763,N_10462,N_10428);
nand U10764 (N_10764,N_10580,N_10532);
and U10765 (N_10765,N_10480,N_10536);
nor U10766 (N_10766,N_10572,N_10473);
nor U10767 (N_10767,N_10562,N_10547);
nand U10768 (N_10768,N_10550,N_10402);
or U10769 (N_10769,N_10445,N_10447);
or U10770 (N_10770,N_10414,N_10460);
and U10771 (N_10771,N_10496,N_10433);
and U10772 (N_10772,N_10591,N_10410);
nor U10773 (N_10773,N_10443,N_10585);
or U10774 (N_10774,N_10581,N_10567);
nor U10775 (N_10775,N_10543,N_10445);
xnor U10776 (N_10776,N_10431,N_10533);
or U10777 (N_10777,N_10558,N_10427);
nor U10778 (N_10778,N_10461,N_10589);
or U10779 (N_10779,N_10565,N_10427);
and U10780 (N_10780,N_10518,N_10418);
and U10781 (N_10781,N_10524,N_10554);
or U10782 (N_10782,N_10520,N_10417);
nor U10783 (N_10783,N_10444,N_10467);
nor U10784 (N_10784,N_10421,N_10412);
or U10785 (N_10785,N_10589,N_10450);
nand U10786 (N_10786,N_10494,N_10515);
or U10787 (N_10787,N_10411,N_10406);
or U10788 (N_10788,N_10480,N_10412);
and U10789 (N_10789,N_10494,N_10565);
nor U10790 (N_10790,N_10508,N_10523);
nand U10791 (N_10791,N_10542,N_10470);
and U10792 (N_10792,N_10584,N_10540);
or U10793 (N_10793,N_10431,N_10570);
xnor U10794 (N_10794,N_10590,N_10473);
nand U10795 (N_10795,N_10404,N_10538);
nor U10796 (N_10796,N_10554,N_10589);
nand U10797 (N_10797,N_10525,N_10487);
and U10798 (N_10798,N_10458,N_10560);
nand U10799 (N_10799,N_10587,N_10526);
nor U10800 (N_10800,N_10648,N_10664);
nor U10801 (N_10801,N_10689,N_10683);
and U10802 (N_10802,N_10742,N_10791);
nand U10803 (N_10803,N_10619,N_10758);
and U10804 (N_10804,N_10681,N_10734);
nor U10805 (N_10805,N_10631,N_10719);
or U10806 (N_10806,N_10700,N_10751);
nand U10807 (N_10807,N_10729,N_10602);
nand U10808 (N_10808,N_10653,N_10651);
nor U10809 (N_10809,N_10647,N_10748);
and U10810 (N_10810,N_10665,N_10762);
or U10811 (N_10811,N_10600,N_10777);
nand U10812 (N_10812,N_10636,N_10660);
or U10813 (N_10813,N_10711,N_10629);
or U10814 (N_10814,N_10769,N_10644);
or U10815 (N_10815,N_10618,N_10639);
nor U10816 (N_10816,N_10690,N_10720);
nand U10817 (N_10817,N_10684,N_10753);
nand U10818 (N_10818,N_10642,N_10691);
and U10819 (N_10819,N_10735,N_10756);
nor U10820 (N_10820,N_10633,N_10725);
or U10821 (N_10821,N_10780,N_10792);
and U10822 (N_10822,N_10652,N_10787);
or U10823 (N_10823,N_10727,N_10752);
nand U10824 (N_10824,N_10718,N_10646);
nor U10825 (N_10825,N_10784,N_10692);
nand U10826 (N_10826,N_10702,N_10772);
or U10827 (N_10827,N_10715,N_10797);
nand U10828 (N_10828,N_10616,N_10697);
nor U10829 (N_10829,N_10632,N_10626);
or U10830 (N_10830,N_10782,N_10606);
nor U10831 (N_10831,N_10658,N_10678);
or U10832 (N_10832,N_10737,N_10650);
and U10833 (N_10833,N_10789,N_10793);
nand U10834 (N_10834,N_10614,N_10688);
nand U10835 (N_10835,N_10667,N_10798);
or U10836 (N_10836,N_10745,N_10649);
nand U10837 (N_10837,N_10721,N_10628);
nand U10838 (N_10838,N_10739,N_10669);
and U10839 (N_10839,N_10731,N_10637);
and U10840 (N_10840,N_10761,N_10607);
nand U10841 (N_10841,N_10736,N_10612);
nand U10842 (N_10842,N_10682,N_10638);
and U10843 (N_10843,N_10749,N_10712);
and U10844 (N_10844,N_10738,N_10645);
and U10845 (N_10845,N_10795,N_10770);
and U10846 (N_10846,N_10760,N_10617);
or U10847 (N_10847,N_10601,N_10695);
nor U10848 (N_10848,N_10754,N_10698);
nor U10849 (N_10849,N_10679,N_10701);
nor U10850 (N_10850,N_10783,N_10613);
or U10851 (N_10851,N_10705,N_10611);
nor U10852 (N_10852,N_10709,N_10670);
or U10853 (N_10853,N_10696,N_10656);
nor U10854 (N_10854,N_10620,N_10680);
nand U10855 (N_10855,N_10757,N_10746);
nor U10856 (N_10856,N_10774,N_10763);
nand U10857 (N_10857,N_10659,N_10625);
nand U10858 (N_10858,N_10661,N_10786);
or U10859 (N_10859,N_10641,N_10759);
and U10860 (N_10860,N_10766,N_10703);
nor U10861 (N_10861,N_10710,N_10730);
nor U10862 (N_10862,N_10704,N_10785);
and U10863 (N_10863,N_10741,N_10671);
nand U10864 (N_10864,N_10673,N_10716);
or U10865 (N_10865,N_10621,N_10676);
or U10866 (N_10866,N_10687,N_10672);
and U10867 (N_10867,N_10694,N_10771);
nand U10868 (N_10868,N_10765,N_10615);
and U10869 (N_10869,N_10778,N_10723);
nand U10870 (N_10870,N_10685,N_10790);
or U10871 (N_10871,N_10686,N_10609);
or U10872 (N_10872,N_10728,N_10605);
or U10873 (N_10873,N_10726,N_10717);
and U10874 (N_10874,N_10747,N_10773);
nand U10875 (N_10875,N_10714,N_10744);
and U10876 (N_10876,N_10634,N_10799);
and U10877 (N_10877,N_10767,N_10724);
and U10878 (N_10878,N_10630,N_10779);
nand U10879 (N_10879,N_10608,N_10768);
nor U10880 (N_10880,N_10677,N_10781);
or U10881 (N_10881,N_10707,N_10627);
nor U10882 (N_10882,N_10635,N_10794);
or U10883 (N_10883,N_10663,N_10713);
and U10884 (N_10884,N_10668,N_10623);
nor U10885 (N_10885,N_10655,N_10740);
or U10886 (N_10886,N_10674,N_10733);
nor U10887 (N_10887,N_10743,N_10675);
and U10888 (N_10888,N_10603,N_10775);
nand U10889 (N_10889,N_10604,N_10654);
nor U10890 (N_10890,N_10755,N_10788);
or U10891 (N_10891,N_10764,N_10708);
nand U10892 (N_10892,N_10706,N_10750);
nor U10893 (N_10893,N_10610,N_10732);
nand U10894 (N_10894,N_10643,N_10657);
or U10895 (N_10895,N_10624,N_10666);
and U10896 (N_10896,N_10640,N_10796);
nand U10897 (N_10897,N_10662,N_10699);
nor U10898 (N_10898,N_10722,N_10622);
or U10899 (N_10899,N_10776,N_10693);
nor U10900 (N_10900,N_10633,N_10751);
nor U10901 (N_10901,N_10764,N_10698);
nand U10902 (N_10902,N_10780,N_10647);
or U10903 (N_10903,N_10717,N_10687);
nand U10904 (N_10904,N_10631,N_10717);
or U10905 (N_10905,N_10780,N_10750);
nand U10906 (N_10906,N_10616,N_10618);
nand U10907 (N_10907,N_10666,N_10731);
and U10908 (N_10908,N_10768,N_10729);
nand U10909 (N_10909,N_10765,N_10691);
nand U10910 (N_10910,N_10605,N_10671);
nand U10911 (N_10911,N_10627,N_10640);
and U10912 (N_10912,N_10696,N_10703);
or U10913 (N_10913,N_10609,N_10623);
nand U10914 (N_10914,N_10601,N_10608);
or U10915 (N_10915,N_10678,N_10623);
nand U10916 (N_10916,N_10770,N_10754);
and U10917 (N_10917,N_10691,N_10639);
and U10918 (N_10918,N_10649,N_10720);
nor U10919 (N_10919,N_10659,N_10680);
or U10920 (N_10920,N_10672,N_10757);
or U10921 (N_10921,N_10610,N_10787);
nor U10922 (N_10922,N_10602,N_10770);
and U10923 (N_10923,N_10600,N_10747);
nand U10924 (N_10924,N_10661,N_10728);
nand U10925 (N_10925,N_10763,N_10714);
and U10926 (N_10926,N_10735,N_10612);
or U10927 (N_10927,N_10634,N_10768);
nor U10928 (N_10928,N_10762,N_10718);
nand U10929 (N_10929,N_10777,N_10645);
nor U10930 (N_10930,N_10611,N_10640);
nand U10931 (N_10931,N_10785,N_10649);
nor U10932 (N_10932,N_10667,N_10661);
and U10933 (N_10933,N_10676,N_10716);
nor U10934 (N_10934,N_10717,N_10713);
nor U10935 (N_10935,N_10781,N_10767);
nand U10936 (N_10936,N_10665,N_10700);
and U10937 (N_10937,N_10739,N_10747);
or U10938 (N_10938,N_10778,N_10660);
nand U10939 (N_10939,N_10657,N_10699);
or U10940 (N_10940,N_10646,N_10659);
nor U10941 (N_10941,N_10642,N_10635);
nor U10942 (N_10942,N_10629,N_10639);
nand U10943 (N_10943,N_10741,N_10735);
nor U10944 (N_10944,N_10693,N_10725);
nor U10945 (N_10945,N_10778,N_10732);
nor U10946 (N_10946,N_10771,N_10635);
nand U10947 (N_10947,N_10715,N_10760);
nand U10948 (N_10948,N_10605,N_10660);
nor U10949 (N_10949,N_10775,N_10605);
nand U10950 (N_10950,N_10690,N_10759);
nor U10951 (N_10951,N_10792,N_10767);
and U10952 (N_10952,N_10707,N_10724);
or U10953 (N_10953,N_10754,N_10729);
or U10954 (N_10954,N_10766,N_10794);
nor U10955 (N_10955,N_10602,N_10682);
and U10956 (N_10956,N_10682,N_10680);
or U10957 (N_10957,N_10726,N_10711);
or U10958 (N_10958,N_10617,N_10603);
nor U10959 (N_10959,N_10677,N_10626);
or U10960 (N_10960,N_10686,N_10683);
and U10961 (N_10961,N_10608,N_10694);
nand U10962 (N_10962,N_10677,N_10748);
nand U10963 (N_10963,N_10794,N_10733);
nand U10964 (N_10964,N_10642,N_10770);
or U10965 (N_10965,N_10689,N_10756);
nor U10966 (N_10966,N_10622,N_10726);
nor U10967 (N_10967,N_10744,N_10616);
or U10968 (N_10968,N_10759,N_10761);
or U10969 (N_10969,N_10770,N_10792);
and U10970 (N_10970,N_10673,N_10625);
nor U10971 (N_10971,N_10642,N_10776);
and U10972 (N_10972,N_10681,N_10755);
or U10973 (N_10973,N_10798,N_10695);
and U10974 (N_10974,N_10731,N_10634);
and U10975 (N_10975,N_10744,N_10772);
or U10976 (N_10976,N_10726,N_10786);
nor U10977 (N_10977,N_10616,N_10693);
or U10978 (N_10978,N_10642,N_10721);
and U10979 (N_10979,N_10782,N_10751);
nor U10980 (N_10980,N_10665,N_10660);
nand U10981 (N_10981,N_10631,N_10625);
nor U10982 (N_10982,N_10613,N_10677);
and U10983 (N_10983,N_10663,N_10681);
nor U10984 (N_10984,N_10629,N_10732);
or U10985 (N_10985,N_10672,N_10649);
or U10986 (N_10986,N_10696,N_10665);
nand U10987 (N_10987,N_10712,N_10663);
nor U10988 (N_10988,N_10776,N_10687);
nand U10989 (N_10989,N_10730,N_10677);
and U10990 (N_10990,N_10714,N_10603);
or U10991 (N_10991,N_10634,N_10669);
and U10992 (N_10992,N_10697,N_10669);
nand U10993 (N_10993,N_10751,N_10772);
or U10994 (N_10994,N_10708,N_10735);
or U10995 (N_10995,N_10701,N_10753);
and U10996 (N_10996,N_10757,N_10696);
nor U10997 (N_10997,N_10770,N_10633);
or U10998 (N_10998,N_10780,N_10710);
and U10999 (N_10999,N_10627,N_10680);
or U11000 (N_11000,N_10956,N_10830);
nor U11001 (N_11001,N_10902,N_10847);
nor U11002 (N_11002,N_10988,N_10971);
nand U11003 (N_11003,N_10961,N_10877);
or U11004 (N_11004,N_10917,N_10922);
nor U11005 (N_11005,N_10957,N_10976);
or U11006 (N_11006,N_10849,N_10974);
or U11007 (N_11007,N_10869,N_10803);
or U11008 (N_11008,N_10891,N_10814);
nor U11009 (N_11009,N_10929,N_10874);
nor U11010 (N_11010,N_10817,N_10898);
or U11011 (N_11011,N_10827,N_10811);
nor U11012 (N_11012,N_10839,N_10805);
and U11013 (N_11013,N_10861,N_10953);
and U11014 (N_11014,N_10809,N_10920);
nand U11015 (N_11015,N_10986,N_10822);
nand U11016 (N_11016,N_10975,N_10875);
nor U11017 (N_11017,N_10889,N_10904);
nand U11018 (N_11018,N_10853,N_10940);
or U11019 (N_11019,N_10866,N_10895);
or U11020 (N_11020,N_10941,N_10810);
nor U11021 (N_11021,N_10828,N_10960);
and U11022 (N_11022,N_10867,N_10980);
and U11023 (N_11023,N_10963,N_10883);
nor U11024 (N_11024,N_10862,N_10845);
and U11025 (N_11025,N_10958,N_10838);
or U11026 (N_11026,N_10854,N_10965);
and U11027 (N_11027,N_10824,N_10944);
and U11028 (N_11028,N_10892,N_10856);
and U11029 (N_11029,N_10930,N_10926);
and U11030 (N_11030,N_10816,N_10897);
nor U11031 (N_11031,N_10846,N_10914);
and U11032 (N_11032,N_10802,N_10978);
xor U11033 (N_11033,N_10977,N_10800);
or U11034 (N_11034,N_10871,N_10851);
or U11035 (N_11035,N_10959,N_10999);
nor U11036 (N_11036,N_10907,N_10969);
and U11037 (N_11037,N_10996,N_10860);
nand U11038 (N_11038,N_10865,N_10968);
nor U11039 (N_11039,N_10842,N_10807);
and U11040 (N_11040,N_10890,N_10893);
nand U11041 (N_11041,N_10880,N_10801);
or U11042 (N_11042,N_10858,N_10911);
or U11043 (N_11043,N_10912,N_10937);
nor U11044 (N_11044,N_10832,N_10910);
and U11045 (N_11045,N_10994,N_10868);
nor U11046 (N_11046,N_10964,N_10908);
nand U11047 (N_11047,N_10885,N_10825);
nor U11048 (N_11048,N_10947,N_10995);
nor U11049 (N_11049,N_10900,N_10821);
nor U11050 (N_11050,N_10924,N_10925);
and U11051 (N_11051,N_10984,N_10991);
or U11052 (N_11052,N_10967,N_10836);
nor U11053 (N_11053,N_10834,N_10921);
nor U11054 (N_11054,N_10997,N_10992);
nor U11055 (N_11055,N_10913,N_10927);
and U11056 (N_11056,N_10804,N_10990);
nor U11057 (N_11057,N_10833,N_10973);
nor U11058 (N_11058,N_10903,N_10939);
nor U11059 (N_11059,N_10955,N_10863);
nor U11060 (N_11060,N_10935,N_10837);
nor U11061 (N_11061,N_10981,N_10818);
or U11062 (N_11062,N_10870,N_10936);
or U11063 (N_11063,N_10933,N_10923);
nor U11064 (N_11064,N_10843,N_10979);
nand U11065 (N_11065,N_10873,N_10872);
nand U11066 (N_11066,N_10819,N_10848);
and U11067 (N_11067,N_10882,N_10962);
nand U11068 (N_11068,N_10951,N_10859);
and U11069 (N_11069,N_10950,N_10982);
nand U11070 (N_11070,N_10876,N_10966);
or U11071 (N_11071,N_10894,N_10983);
and U11072 (N_11072,N_10972,N_10918);
and U11073 (N_11073,N_10806,N_10948);
and U11074 (N_11074,N_10943,N_10906);
or U11075 (N_11075,N_10954,N_10915);
or U11076 (N_11076,N_10896,N_10899);
and U11077 (N_11077,N_10820,N_10998);
nor U11078 (N_11078,N_10823,N_10886);
nand U11079 (N_11079,N_10844,N_10934);
nor U11080 (N_11080,N_10829,N_10855);
nor U11081 (N_11081,N_10815,N_10881);
and U11082 (N_11082,N_10919,N_10987);
nor U11083 (N_11083,N_10808,N_10970);
or U11084 (N_11084,N_10864,N_10879);
nor U11085 (N_11085,N_10905,N_10928);
and U11086 (N_11086,N_10952,N_10841);
nand U11087 (N_11087,N_10884,N_10831);
xnor U11088 (N_11088,N_10945,N_10901);
nand U11089 (N_11089,N_10813,N_10932);
and U11090 (N_11090,N_10993,N_10812);
and U11091 (N_11091,N_10989,N_10840);
nand U11092 (N_11092,N_10942,N_10852);
nor U11093 (N_11093,N_10887,N_10938);
and U11094 (N_11094,N_10985,N_10826);
nor U11095 (N_11095,N_10931,N_10835);
nor U11096 (N_11096,N_10850,N_10949);
and U11097 (N_11097,N_10946,N_10888);
and U11098 (N_11098,N_10916,N_10878);
nor U11099 (N_11099,N_10857,N_10909);
and U11100 (N_11100,N_10930,N_10947);
and U11101 (N_11101,N_10998,N_10829);
nor U11102 (N_11102,N_10826,N_10916);
nand U11103 (N_11103,N_10874,N_10865);
or U11104 (N_11104,N_10817,N_10902);
nand U11105 (N_11105,N_10955,N_10991);
or U11106 (N_11106,N_10840,N_10967);
nor U11107 (N_11107,N_10850,N_10837);
and U11108 (N_11108,N_10880,N_10960);
and U11109 (N_11109,N_10803,N_10884);
nand U11110 (N_11110,N_10831,N_10834);
nor U11111 (N_11111,N_10832,N_10922);
nor U11112 (N_11112,N_10933,N_10993);
nand U11113 (N_11113,N_10876,N_10955);
nand U11114 (N_11114,N_10964,N_10967);
nand U11115 (N_11115,N_10947,N_10963);
and U11116 (N_11116,N_10843,N_10885);
nand U11117 (N_11117,N_10828,N_10888);
and U11118 (N_11118,N_10906,N_10836);
nor U11119 (N_11119,N_10966,N_10875);
nor U11120 (N_11120,N_10870,N_10821);
nor U11121 (N_11121,N_10900,N_10923);
or U11122 (N_11122,N_10830,N_10988);
nand U11123 (N_11123,N_10930,N_10809);
nand U11124 (N_11124,N_10971,N_10981);
and U11125 (N_11125,N_10920,N_10818);
nand U11126 (N_11126,N_10874,N_10801);
or U11127 (N_11127,N_10939,N_10865);
and U11128 (N_11128,N_10906,N_10948);
nand U11129 (N_11129,N_10837,N_10846);
or U11130 (N_11130,N_10876,N_10995);
nand U11131 (N_11131,N_10820,N_10947);
and U11132 (N_11132,N_10929,N_10804);
nand U11133 (N_11133,N_10937,N_10855);
nor U11134 (N_11134,N_10986,N_10858);
or U11135 (N_11135,N_10888,N_10935);
or U11136 (N_11136,N_10934,N_10900);
and U11137 (N_11137,N_10920,N_10821);
nand U11138 (N_11138,N_10966,N_10836);
xor U11139 (N_11139,N_10909,N_10897);
or U11140 (N_11140,N_10945,N_10816);
and U11141 (N_11141,N_10898,N_10961);
or U11142 (N_11142,N_10823,N_10895);
nand U11143 (N_11143,N_10800,N_10834);
and U11144 (N_11144,N_10838,N_10845);
or U11145 (N_11145,N_10865,N_10952);
and U11146 (N_11146,N_10828,N_10815);
xnor U11147 (N_11147,N_10905,N_10839);
nor U11148 (N_11148,N_10877,N_10912);
or U11149 (N_11149,N_10950,N_10873);
and U11150 (N_11150,N_10997,N_10850);
or U11151 (N_11151,N_10840,N_10879);
nor U11152 (N_11152,N_10933,N_10988);
nand U11153 (N_11153,N_10857,N_10841);
nor U11154 (N_11154,N_10869,N_10890);
nor U11155 (N_11155,N_10827,N_10856);
nor U11156 (N_11156,N_10926,N_10959);
nor U11157 (N_11157,N_10840,N_10925);
or U11158 (N_11158,N_10891,N_10905);
nor U11159 (N_11159,N_10929,N_10860);
nor U11160 (N_11160,N_10906,N_10875);
and U11161 (N_11161,N_10805,N_10890);
or U11162 (N_11162,N_10918,N_10845);
nor U11163 (N_11163,N_10876,N_10963);
or U11164 (N_11164,N_10900,N_10978);
or U11165 (N_11165,N_10981,N_10948);
or U11166 (N_11166,N_10900,N_10959);
nor U11167 (N_11167,N_10848,N_10827);
or U11168 (N_11168,N_10962,N_10910);
or U11169 (N_11169,N_10920,N_10919);
nand U11170 (N_11170,N_10989,N_10903);
or U11171 (N_11171,N_10879,N_10904);
nand U11172 (N_11172,N_10941,N_10961);
nor U11173 (N_11173,N_10920,N_10954);
nand U11174 (N_11174,N_10977,N_10901);
nand U11175 (N_11175,N_10988,N_10860);
or U11176 (N_11176,N_10846,N_10872);
and U11177 (N_11177,N_10898,N_10992);
and U11178 (N_11178,N_10971,N_10982);
nor U11179 (N_11179,N_10911,N_10822);
and U11180 (N_11180,N_10955,N_10853);
or U11181 (N_11181,N_10861,N_10923);
nor U11182 (N_11182,N_10991,N_10924);
nor U11183 (N_11183,N_10884,N_10811);
nand U11184 (N_11184,N_10896,N_10818);
nand U11185 (N_11185,N_10919,N_10805);
nand U11186 (N_11186,N_10829,N_10825);
nand U11187 (N_11187,N_10916,N_10849);
nor U11188 (N_11188,N_10922,N_10818);
nor U11189 (N_11189,N_10860,N_10848);
nand U11190 (N_11190,N_10965,N_10816);
and U11191 (N_11191,N_10937,N_10802);
nand U11192 (N_11192,N_10818,N_10802);
or U11193 (N_11193,N_10908,N_10830);
nor U11194 (N_11194,N_10994,N_10913);
or U11195 (N_11195,N_10966,N_10888);
nor U11196 (N_11196,N_10994,N_10978);
nor U11197 (N_11197,N_10966,N_10857);
nor U11198 (N_11198,N_10978,N_10888);
nor U11199 (N_11199,N_10920,N_10851);
nand U11200 (N_11200,N_11177,N_11184);
nand U11201 (N_11201,N_11017,N_11147);
and U11202 (N_11202,N_11118,N_11145);
nor U11203 (N_11203,N_11079,N_11014);
or U11204 (N_11204,N_11161,N_11087);
nor U11205 (N_11205,N_11039,N_11022);
and U11206 (N_11206,N_11018,N_11028);
nand U11207 (N_11207,N_11163,N_11178);
nand U11208 (N_11208,N_11174,N_11012);
nand U11209 (N_11209,N_11197,N_11053);
or U11210 (N_11210,N_11153,N_11157);
xor U11211 (N_11211,N_11007,N_11046);
xor U11212 (N_11212,N_11055,N_11054);
nand U11213 (N_11213,N_11098,N_11096);
nor U11214 (N_11214,N_11035,N_11063);
or U11215 (N_11215,N_11158,N_11193);
nor U11216 (N_11216,N_11072,N_11132);
and U11217 (N_11217,N_11070,N_11001);
and U11218 (N_11218,N_11099,N_11038);
and U11219 (N_11219,N_11150,N_11092);
nor U11220 (N_11220,N_11032,N_11069);
nor U11221 (N_11221,N_11121,N_11033);
or U11222 (N_11222,N_11059,N_11195);
or U11223 (N_11223,N_11029,N_11137);
or U11224 (N_11224,N_11142,N_11073);
nor U11225 (N_11225,N_11052,N_11122);
or U11226 (N_11226,N_11058,N_11152);
nor U11227 (N_11227,N_11000,N_11144);
and U11228 (N_11228,N_11068,N_11189);
and U11229 (N_11229,N_11196,N_11135);
nand U11230 (N_11230,N_11160,N_11107);
or U11231 (N_11231,N_11003,N_11190);
nand U11232 (N_11232,N_11192,N_11179);
nand U11233 (N_11233,N_11019,N_11175);
nor U11234 (N_11234,N_11113,N_11084);
nor U11235 (N_11235,N_11101,N_11108);
and U11236 (N_11236,N_11119,N_11047);
and U11237 (N_11237,N_11149,N_11091);
nand U11238 (N_11238,N_11106,N_11131);
and U11239 (N_11239,N_11020,N_11164);
and U11240 (N_11240,N_11146,N_11042);
and U11241 (N_11241,N_11067,N_11181);
nand U11242 (N_11242,N_11114,N_11148);
or U11243 (N_11243,N_11031,N_11102);
and U11244 (N_11244,N_11010,N_11051);
and U11245 (N_11245,N_11016,N_11186);
nor U11246 (N_11246,N_11088,N_11097);
nor U11247 (N_11247,N_11078,N_11129);
nand U11248 (N_11248,N_11095,N_11185);
and U11249 (N_11249,N_11110,N_11117);
nand U11250 (N_11250,N_11040,N_11109);
or U11251 (N_11251,N_11011,N_11116);
and U11252 (N_11252,N_11030,N_11015);
nand U11253 (N_11253,N_11100,N_11176);
nand U11254 (N_11254,N_11115,N_11009);
nor U11255 (N_11255,N_11105,N_11151);
and U11256 (N_11256,N_11075,N_11002);
nor U11257 (N_11257,N_11006,N_11198);
nand U11258 (N_11258,N_11170,N_11044);
and U11259 (N_11259,N_11036,N_11090);
and U11260 (N_11260,N_11133,N_11043);
nand U11261 (N_11261,N_11077,N_11143);
nand U11262 (N_11262,N_11050,N_11187);
nor U11263 (N_11263,N_11180,N_11080);
nand U11264 (N_11264,N_11167,N_11159);
nand U11265 (N_11265,N_11191,N_11104);
nor U11266 (N_11266,N_11013,N_11103);
or U11267 (N_11267,N_11127,N_11188);
nand U11268 (N_11268,N_11045,N_11083);
nor U11269 (N_11269,N_11156,N_11123);
and U11270 (N_11270,N_11048,N_11074);
or U11271 (N_11271,N_11111,N_11140);
and U11272 (N_11272,N_11071,N_11182);
nand U11273 (N_11273,N_11076,N_11124);
nor U11274 (N_11274,N_11008,N_11005);
or U11275 (N_11275,N_11171,N_11037);
nor U11276 (N_11276,N_11112,N_11065);
nand U11277 (N_11277,N_11120,N_11089);
or U11278 (N_11278,N_11134,N_11024);
or U11279 (N_11279,N_11130,N_11027);
and U11280 (N_11280,N_11155,N_11199);
and U11281 (N_11281,N_11049,N_11061);
and U11282 (N_11282,N_11141,N_11085);
nor U11283 (N_11283,N_11125,N_11004);
and U11284 (N_11284,N_11025,N_11168);
and U11285 (N_11285,N_11139,N_11166);
or U11286 (N_11286,N_11172,N_11082);
nor U11287 (N_11287,N_11023,N_11060);
or U11288 (N_11288,N_11126,N_11034);
nand U11289 (N_11289,N_11066,N_11081);
and U11290 (N_11290,N_11094,N_11162);
nor U11291 (N_11291,N_11138,N_11194);
or U11292 (N_11292,N_11093,N_11136);
nor U11293 (N_11293,N_11064,N_11173);
nand U11294 (N_11294,N_11169,N_11021);
and U11295 (N_11295,N_11165,N_11057);
nand U11296 (N_11296,N_11041,N_11154);
nand U11297 (N_11297,N_11183,N_11128);
and U11298 (N_11298,N_11056,N_11086);
nor U11299 (N_11299,N_11062,N_11026);
nor U11300 (N_11300,N_11194,N_11017);
nor U11301 (N_11301,N_11025,N_11004);
nand U11302 (N_11302,N_11197,N_11163);
and U11303 (N_11303,N_11163,N_11062);
or U11304 (N_11304,N_11109,N_11135);
and U11305 (N_11305,N_11121,N_11013);
nand U11306 (N_11306,N_11199,N_11178);
nor U11307 (N_11307,N_11063,N_11107);
and U11308 (N_11308,N_11037,N_11112);
nor U11309 (N_11309,N_11047,N_11054);
nor U11310 (N_11310,N_11014,N_11086);
xnor U11311 (N_11311,N_11159,N_11101);
nand U11312 (N_11312,N_11132,N_11041);
and U11313 (N_11313,N_11060,N_11076);
and U11314 (N_11314,N_11111,N_11065);
nor U11315 (N_11315,N_11030,N_11027);
nor U11316 (N_11316,N_11112,N_11093);
and U11317 (N_11317,N_11154,N_11023);
nand U11318 (N_11318,N_11013,N_11021);
and U11319 (N_11319,N_11128,N_11077);
and U11320 (N_11320,N_11141,N_11008);
nor U11321 (N_11321,N_11131,N_11103);
nor U11322 (N_11322,N_11006,N_11100);
or U11323 (N_11323,N_11015,N_11088);
and U11324 (N_11324,N_11134,N_11198);
and U11325 (N_11325,N_11023,N_11188);
nor U11326 (N_11326,N_11122,N_11053);
and U11327 (N_11327,N_11145,N_11182);
nor U11328 (N_11328,N_11083,N_11031);
and U11329 (N_11329,N_11108,N_11162);
nor U11330 (N_11330,N_11013,N_11105);
nand U11331 (N_11331,N_11070,N_11135);
and U11332 (N_11332,N_11177,N_11118);
or U11333 (N_11333,N_11085,N_11110);
and U11334 (N_11334,N_11098,N_11177);
and U11335 (N_11335,N_11028,N_11121);
and U11336 (N_11336,N_11019,N_11018);
and U11337 (N_11337,N_11000,N_11155);
nor U11338 (N_11338,N_11077,N_11070);
nor U11339 (N_11339,N_11072,N_11009);
nor U11340 (N_11340,N_11066,N_11161);
nor U11341 (N_11341,N_11134,N_11127);
or U11342 (N_11342,N_11105,N_11132);
nor U11343 (N_11343,N_11029,N_11008);
or U11344 (N_11344,N_11155,N_11029);
and U11345 (N_11345,N_11109,N_11151);
and U11346 (N_11346,N_11130,N_11106);
and U11347 (N_11347,N_11158,N_11116);
and U11348 (N_11348,N_11150,N_11187);
or U11349 (N_11349,N_11120,N_11048);
or U11350 (N_11350,N_11066,N_11125);
nor U11351 (N_11351,N_11065,N_11130);
nor U11352 (N_11352,N_11085,N_11036);
and U11353 (N_11353,N_11164,N_11133);
or U11354 (N_11354,N_11159,N_11008);
or U11355 (N_11355,N_11088,N_11010);
nor U11356 (N_11356,N_11118,N_11037);
or U11357 (N_11357,N_11137,N_11040);
xor U11358 (N_11358,N_11125,N_11019);
nor U11359 (N_11359,N_11072,N_11088);
or U11360 (N_11360,N_11027,N_11171);
or U11361 (N_11361,N_11037,N_11109);
nor U11362 (N_11362,N_11144,N_11123);
or U11363 (N_11363,N_11109,N_11108);
and U11364 (N_11364,N_11152,N_11074);
nor U11365 (N_11365,N_11061,N_11103);
nand U11366 (N_11366,N_11134,N_11155);
or U11367 (N_11367,N_11061,N_11117);
or U11368 (N_11368,N_11070,N_11011);
nand U11369 (N_11369,N_11150,N_11170);
nand U11370 (N_11370,N_11031,N_11003);
or U11371 (N_11371,N_11192,N_11175);
or U11372 (N_11372,N_11015,N_11017);
and U11373 (N_11373,N_11093,N_11194);
or U11374 (N_11374,N_11062,N_11079);
or U11375 (N_11375,N_11043,N_11087);
nor U11376 (N_11376,N_11047,N_11148);
or U11377 (N_11377,N_11026,N_11121);
nand U11378 (N_11378,N_11130,N_11013);
or U11379 (N_11379,N_11154,N_11169);
or U11380 (N_11380,N_11197,N_11054);
nor U11381 (N_11381,N_11072,N_11011);
nand U11382 (N_11382,N_11148,N_11098);
and U11383 (N_11383,N_11050,N_11083);
or U11384 (N_11384,N_11117,N_11124);
xnor U11385 (N_11385,N_11123,N_11185);
and U11386 (N_11386,N_11088,N_11050);
and U11387 (N_11387,N_11190,N_11103);
and U11388 (N_11388,N_11174,N_11146);
nand U11389 (N_11389,N_11050,N_11151);
nand U11390 (N_11390,N_11077,N_11027);
or U11391 (N_11391,N_11144,N_11092);
and U11392 (N_11392,N_11192,N_11199);
and U11393 (N_11393,N_11147,N_11105);
nand U11394 (N_11394,N_11125,N_11122);
or U11395 (N_11395,N_11075,N_11057);
nor U11396 (N_11396,N_11067,N_11147);
nor U11397 (N_11397,N_11013,N_11162);
nor U11398 (N_11398,N_11040,N_11175);
or U11399 (N_11399,N_11012,N_11091);
or U11400 (N_11400,N_11207,N_11339);
nor U11401 (N_11401,N_11210,N_11319);
and U11402 (N_11402,N_11272,N_11204);
and U11403 (N_11403,N_11393,N_11373);
or U11404 (N_11404,N_11254,N_11318);
or U11405 (N_11405,N_11300,N_11322);
and U11406 (N_11406,N_11276,N_11290);
nor U11407 (N_11407,N_11231,N_11235);
and U11408 (N_11408,N_11252,N_11321);
and U11409 (N_11409,N_11262,N_11338);
nor U11410 (N_11410,N_11333,N_11245);
nor U11411 (N_11411,N_11381,N_11372);
nor U11412 (N_11412,N_11340,N_11326);
and U11413 (N_11413,N_11253,N_11361);
nand U11414 (N_11414,N_11396,N_11221);
and U11415 (N_11415,N_11232,N_11279);
nor U11416 (N_11416,N_11224,N_11266);
nand U11417 (N_11417,N_11310,N_11330);
nor U11418 (N_11418,N_11202,N_11269);
or U11419 (N_11419,N_11256,N_11246);
nand U11420 (N_11420,N_11286,N_11385);
or U11421 (N_11421,N_11359,N_11309);
nand U11422 (N_11422,N_11360,N_11354);
nand U11423 (N_11423,N_11352,N_11299);
or U11424 (N_11424,N_11314,N_11275);
nand U11425 (N_11425,N_11344,N_11257);
nand U11426 (N_11426,N_11305,N_11291);
or U11427 (N_11427,N_11260,N_11205);
nand U11428 (N_11428,N_11302,N_11342);
and U11429 (N_11429,N_11311,N_11374);
and U11430 (N_11430,N_11270,N_11239);
and U11431 (N_11431,N_11297,N_11357);
nor U11432 (N_11432,N_11308,N_11370);
nor U11433 (N_11433,N_11241,N_11386);
and U11434 (N_11434,N_11278,N_11325);
nand U11435 (N_11435,N_11225,N_11250);
or U11436 (N_11436,N_11345,N_11394);
or U11437 (N_11437,N_11350,N_11209);
nand U11438 (N_11438,N_11217,N_11214);
or U11439 (N_11439,N_11371,N_11288);
nand U11440 (N_11440,N_11380,N_11324);
xor U11441 (N_11441,N_11289,N_11242);
nand U11442 (N_11442,N_11383,N_11200);
nor U11443 (N_11443,N_11397,N_11218);
or U11444 (N_11444,N_11295,N_11389);
nand U11445 (N_11445,N_11346,N_11395);
nor U11446 (N_11446,N_11223,N_11208);
and U11447 (N_11447,N_11284,N_11366);
or U11448 (N_11448,N_11343,N_11247);
nor U11449 (N_11449,N_11203,N_11329);
nand U11450 (N_11450,N_11331,N_11237);
and U11451 (N_11451,N_11229,N_11391);
and U11452 (N_11452,N_11320,N_11287);
or U11453 (N_11453,N_11244,N_11292);
or U11454 (N_11454,N_11337,N_11296);
nand U11455 (N_11455,N_11271,N_11298);
nand U11456 (N_11456,N_11238,N_11315);
or U11457 (N_11457,N_11390,N_11228);
nor U11458 (N_11458,N_11215,N_11316);
nor U11459 (N_11459,N_11317,N_11261);
and U11460 (N_11460,N_11274,N_11382);
nor U11461 (N_11461,N_11280,N_11376);
or U11462 (N_11462,N_11323,N_11216);
and U11463 (N_11463,N_11334,N_11356);
or U11464 (N_11464,N_11328,N_11236);
nor U11465 (N_11465,N_11358,N_11230);
and U11466 (N_11466,N_11222,N_11384);
and U11467 (N_11467,N_11304,N_11264);
or U11468 (N_11468,N_11303,N_11336);
or U11469 (N_11469,N_11255,N_11277);
or U11470 (N_11470,N_11312,N_11226);
or U11471 (N_11471,N_11377,N_11259);
nor U11472 (N_11472,N_11307,N_11301);
and U11473 (N_11473,N_11349,N_11335);
and U11474 (N_11474,N_11201,N_11392);
nand U11475 (N_11475,N_11398,N_11251);
and U11476 (N_11476,N_11375,N_11353);
or U11477 (N_11477,N_11240,N_11399);
and U11478 (N_11478,N_11362,N_11327);
and U11479 (N_11479,N_11347,N_11234);
nand U11480 (N_11480,N_11294,N_11313);
and U11481 (N_11481,N_11365,N_11378);
and U11482 (N_11482,N_11387,N_11281);
and U11483 (N_11483,N_11364,N_11243);
or U11484 (N_11484,N_11267,N_11282);
nor U11485 (N_11485,N_11388,N_11348);
or U11486 (N_11486,N_11363,N_11268);
and U11487 (N_11487,N_11258,N_11220);
nor U11488 (N_11488,N_11248,N_11283);
or U11489 (N_11489,N_11351,N_11211);
or U11490 (N_11490,N_11293,N_11379);
and U11491 (N_11491,N_11265,N_11367);
nor U11492 (N_11492,N_11233,N_11306);
nand U11493 (N_11493,N_11263,N_11341);
or U11494 (N_11494,N_11368,N_11285);
or U11495 (N_11495,N_11213,N_11206);
and U11496 (N_11496,N_11273,N_11355);
or U11497 (N_11497,N_11332,N_11249);
nor U11498 (N_11498,N_11227,N_11212);
nor U11499 (N_11499,N_11369,N_11219);
nand U11500 (N_11500,N_11284,N_11361);
nand U11501 (N_11501,N_11301,N_11377);
or U11502 (N_11502,N_11203,N_11334);
nor U11503 (N_11503,N_11227,N_11230);
nor U11504 (N_11504,N_11363,N_11239);
nor U11505 (N_11505,N_11260,N_11246);
nor U11506 (N_11506,N_11308,N_11279);
nor U11507 (N_11507,N_11355,N_11347);
nand U11508 (N_11508,N_11261,N_11287);
nand U11509 (N_11509,N_11366,N_11303);
nor U11510 (N_11510,N_11281,N_11256);
nand U11511 (N_11511,N_11290,N_11233);
or U11512 (N_11512,N_11394,N_11358);
nor U11513 (N_11513,N_11295,N_11315);
and U11514 (N_11514,N_11368,N_11340);
or U11515 (N_11515,N_11301,N_11309);
or U11516 (N_11516,N_11390,N_11331);
nand U11517 (N_11517,N_11375,N_11381);
or U11518 (N_11518,N_11371,N_11273);
nand U11519 (N_11519,N_11306,N_11398);
and U11520 (N_11520,N_11387,N_11361);
or U11521 (N_11521,N_11242,N_11221);
nor U11522 (N_11522,N_11222,N_11312);
nand U11523 (N_11523,N_11399,N_11267);
nor U11524 (N_11524,N_11371,N_11305);
and U11525 (N_11525,N_11239,N_11323);
xor U11526 (N_11526,N_11207,N_11262);
nand U11527 (N_11527,N_11351,N_11242);
or U11528 (N_11528,N_11312,N_11254);
or U11529 (N_11529,N_11350,N_11270);
and U11530 (N_11530,N_11327,N_11217);
nand U11531 (N_11531,N_11261,N_11209);
nand U11532 (N_11532,N_11330,N_11309);
or U11533 (N_11533,N_11391,N_11269);
or U11534 (N_11534,N_11392,N_11312);
nand U11535 (N_11535,N_11215,N_11280);
nor U11536 (N_11536,N_11209,N_11342);
nor U11537 (N_11537,N_11292,N_11322);
and U11538 (N_11538,N_11279,N_11228);
nor U11539 (N_11539,N_11210,N_11213);
nand U11540 (N_11540,N_11295,N_11217);
nand U11541 (N_11541,N_11374,N_11369);
or U11542 (N_11542,N_11384,N_11315);
nor U11543 (N_11543,N_11397,N_11330);
or U11544 (N_11544,N_11261,N_11245);
nand U11545 (N_11545,N_11205,N_11263);
and U11546 (N_11546,N_11269,N_11240);
or U11547 (N_11547,N_11362,N_11302);
nand U11548 (N_11548,N_11314,N_11250);
and U11549 (N_11549,N_11388,N_11389);
or U11550 (N_11550,N_11223,N_11374);
or U11551 (N_11551,N_11249,N_11349);
nor U11552 (N_11552,N_11351,N_11245);
and U11553 (N_11553,N_11384,N_11212);
and U11554 (N_11554,N_11294,N_11231);
or U11555 (N_11555,N_11275,N_11204);
nor U11556 (N_11556,N_11341,N_11345);
nor U11557 (N_11557,N_11256,N_11290);
nor U11558 (N_11558,N_11368,N_11326);
and U11559 (N_11559,N_11388,N_11263);
nor U11560 (N_11560,N_11297,N_11362);
or U11561 (N_11561,N_11241,N_11225);
or U11562 (N_11562,N_11295,N_11383);
nor U11563 (N_11563,N_11253,N_11292);
nand U11564 (N_11564,N_11216,N_11202);
nand U11565 (N_11565,N_11365,N_11276);
or U11566 (N_11566,N_11385,N_11283);
and U11567 (N_11567,N_11353,N_11213);
nor U11568 (N_11568,N_11206,N_11287);
nand U11569 (N_11569,N_11242,N_11366);
nand U11570 (N_11570,N_11380,N_11388);
nor U11571 (N_11571,N_11292,N_11355);
and U11572 (N_11572,N_11315,N_11318);
or U11573 (N_11573,N_11382,N_11218);
or U11574 (N_11574,N_11228,N_11328);
nor U11575 (N_11575,N_11260,N_11316);
nor U11576 (N_11576,N_11390,N_11362);
and U11577 (N_11577,N_11380,N_11228);
and U11578 (N_11578,N_11288,N_11264);
nand U11579 (N_11579,N_11232,N_11363);
or U11580 (N_11580,N_11366,N_11328);
and U11581 (N_11581,N_11281,N_11225);
and U11582 (N_11582,N_11297,N_11330);
and U11583 (N_11583,N_11283,N_11326);
nor U11584 (N_11584,N_11344,N_11294);
nor U11585 (N_11585,N_11276,N_11233);
nor U11586 (N_11586,N_11342,N_11283);
and U11587 (N_11587,N_11369,N_11363);
or U11588 (N_11588,N_11373,N_11358);
nand U11589 (N_11589,N_11298,N_11342);
and U11590 (N_11590,N_11385,N_11304);
or U11591 (N_11591,N_11242,N_11258);
and U11592 (N_11592,N_11249,N_11396);
nor U11593 (N_11593,N_11291,N_11361);
or U11594 (N_11594,N_11246,N_11337);
nand U11595 (N_11595,N_11238,N_11242);
and U11596 (N_11596,N_11398,N_11388);
and U11597 (N_11597,N_11293,N_11266);
and U11598 (N_11598,N_11315,N_11327);
and U11599 (N_11599,N_11204,N_11393);
nor U11600 (N_11600,N_11503,N_11449);
or U11601 (N_11601,N_11526,N_11484);
or U11602 (N_11602,N_11438,N_11505);
nand U11603 (N_11603,N_11400,N_11537);
and U11604 (N_11604,N_11508,N_11498);
nand U11605 (N_11605,N_11448,N_11516);
and U11606 (N_11606,N_11429,N_11542);
nor U11607 (N_11607,N_11565,N_11404);
and U11608 (N_11608,N_11468,N_11403);
and U11609 (N_11609,N_11453,N_11479);
nand U11610 (N_11610,N_11599,N_11444);
or U11611 (N_11611,N_11500,N_11519);
nor U11612 (N_11612,N_11591,N_11474);
nor U11613 (N_11613,N_11598,N_11501);
and U11614 (N_11614,N_11483,N_11408);
nor U11615 (N_11615,N_11487,N_11535);
nor U11616 (N_11616,N_11411,N_11545);
and U11617 (N_11617,N_11442,N_11469);
and U11618 (N_11618,N_11549,N_11578);
or U11619 (N_11619,N_11495,N_11527);
nand U11620 (N_11620,N_11424,N_11402);
nor U11621 (N_11621,N_11509,N_11543);
nor U11622 (N_11622,N_11588,N_11513);
nor U11623 (N_11623,N_11546,N_11446);
nor U11624 (N_11624,N_11560,N_11571);
nand U11625 (N_11625,N_11564,N_11557);
nand U11626 (N_11626,N_11412,N_11566);
or U11627 (N_11627,N_11593,N_11428);
nor U11628 (N_11628,N_11451,N_11529);
or U11629 (N_11629,N_11458,N_11540);
nand U11630 (N_11630,N_11491,N_11524);
or U11631 (N_11631,N_11561,N_11525);
nand U11632 (N_11632,N_11471,N_11481);
and U11633 (N_11633,N_11520,N_11413);
nand U11634 (N_11634,N_11436,N_11575);
and U11635 (N_11635,N_11595,N_11430);
nand U11636 (N_11636,N_11559,N_11510);
nand U11637 (N_11637,N_11504,N_11457);
and U11638 (N_11638,N_11531,N_11499);
and U11639 (N_11639,N_11410,N_11415);
and U11640 (N_11640,N_11517,N_11553);
nor U11641 (N_11641,N_11427,N_11550);
nand U11642 (N_11642,N_11456,N_11555);
nand U11643 (N_11643,N_11490,N_11472);
and U11644 (N_11644,N_11482,N_11460);
or U11645 (N_11645,N_11552,N_11554);
nand U11646 (N_11646,N_11434,N_11597);
nand U11647 (N_11647,N_11569,N_11437);
and U11648 (N_11648,N_11574,N_11488);
nand U11649 (N_11649,N_11419,N_11414);
or U11650 (N_11650,N_11558,N_11583);
nand U11651 (N_11651,N_11563,N_11551);
nor U11652 (N_11652,N_11533,N_11450);
or U11653 (N_11653,N_11512,N_11567);
and U11654 (N_11654,N_11594,N_11432);
nand U11655 (N_11655,N_11532,N_11420);
or U11656 (N_11656,N_11506,N_11568);
nor U11657 (N_11657,N_11416,N_11443);
nor U11658 (N_11658,N_11470,N_11476);
and U11659 (N_11659,N_11473,N_11580);
or U11660 (N_11660,N_11492,N_11439);
and U11661 (N_11661,N_11536,N_11480);
nor U11662 (N_11662,N_11461,N_11538);
nand U11663 (N_11663,N_11423,N_11587);
nor U11664 (N_11664,N_11425,N_11507);
nand U11665 (N_11665,N_11530,N_11466);
or U11666 (N_11666,N_11548,N_11445);
or U11667 (N_11667,N_11462,N_11497);
and U11668 (N_11668,N_11447,N_11584);
nand U11669 (N_11669,N_11418,N_11441);
or U11670 (N_11670,N_11486,N_11589);
or U11671 (N_11671,N_11401,N_11477);
nor U11672 (N_11672,N_11539,N_11435);
nand U11673 (N_11673,N_11518,N_11528);
nand U11674 (N_11674,N_11421,N_11586);
nor U11675 (N_11675,N_11455,N_11405);
nand U11676 (N_11676,N_11514,N_11452);
nand U11677 (N_11677,N_11534,N_11464);
nand U11678 (N_11678,N_11478,N_11431);
or U11679 (N_11679,N_11541,N_11422);
nor U11680 (N_11680,N_11544,N_11522);
and U11681 (N_11681,N_11406,N_11485);
or U11682 (N_11682,N_11596,N_11547);
nor U11683 (N_11683,N_11440,N_11459);
and U11684 (N_11684,N_11570,N_11417);
and U11685 (N_11685,N_11523,N_11582);
nor U11686 (N_11686,N_11577,N_11572);
nor U11687 (N_11687,N_11579,N_11511);
or U11688 (N_11688,N_11409,N_11454);
nand U11689 (N_11689,N_11585,N_11496);
nor U11690 (N_11690,N_11590,N_11576);
or U11691 (N_11691,N_11581,N_11592);
or U11692 (N_11692,N_11467,N_11573);
nor U11693 (N_11693,N_11494,N_11433);
xnor U11694 (N_11694,N_11463,N_11493);
nor U11695 (N_11695,N_11562,N_11407);
and U11696 (N_11696,N_11489,N_11502);
nor U11697 (N_11697,N_11475,N_11521);
nand U11698 (N_11698,N_11426,N_11556);
or U11699 (N_11699,N_11465,N_11515);
nand U11700 (N_11700,N_11566,N_11453);
nand U11701 (N_11701,N_11596,N_11556);
or U11702 (N_11702,N_11564,N_11472);
and U11703 (N_11703,N_11544,N_11480);
and U11704 (N_11704,N_11490,N_11403);
and U11705 (N_11705,N_11561,N_11486);
and U11706 (N_11706,N_11481,N_11494);
or U11707 (N_11707,N_11458,N_11598);
or U11708 (N_11708,N_11471,N_11448);
nand U11709 (N_11709,N_11455,N_11565);
or U11710 (N_11710,N_11598,N_11596);
or U11711 (N_11711,N_11463,N_11436);
nor U11712 (N_11712,N_11483,N_11511);
or U11713 (N_11713,N_11574,N_11530);
nand U11714 (N_11714,N_11524,N_11517);
and U11715 (N_11715,N_11440,N_11497);
or U11716 (N_11716,N_11552,N_11495);
nor U11717 (N_11717,N_11456,N_11576);
or U11718 (N_11718,N_11499,N_11438);
nor U11719 (N_11719,N_11478,N_11430);
nand U11720 (N_11720,N_11523,N_11581);
or U11721 (N_11721,N_11567,N_11401);
nor U11722 (N_11722,N_11419,N_11590);
and U11723 (N_11723,N_11559,N_11504);
or U11724 (N_11724,N_11546,N_11522);
and U11725 (N_11725,N_11509,N_11433);
or U11726 (N_11726,N_11524,N_11433);
nor U11727 (N_11727,N_11429,N_11415);
or U11728 (N_11728,N_11404,N_11499);
or U11729 (N_11729,N_11512,N_11513);
nor U11730 (N_11730,N_11448,N_11489);
or U11731 (N_11731,N_11595,N_11466);
nand U11732 (N_11732,N_11415,N_11501);
xor U11733 (N_11733,N_11470,N_11492);
and U11734 (N_11734,N_11454,N_11453);
or U11735 (N_11735,N_11511,N_11468);
and U11736 (N_11736,N_11502,N_11596);
and U11737 (N_11737,N_11569,N_11581);
and U11738 (N_11738,N_11504,N_11446);
or U11739 (N_11739,N_11589,N_11520);
nor U11740 (N_11740,N_11487,N_11455);
or U11741 (N_11741,N_11573,N_11538);
nand U11742 (N_11742,N_11411,N_11472);
nor U11743 (N_11743,N_11403,N_11574);
nand U11744 (N_11744,N_11560,N_11582);
nor U11745 (N_11745,N_11532,N_11564);
nand U11746 (N_11746,N_11530,N_11435);
nor U11747 (N_11747,N_11493,N_11422);
or U11748 (N_11748,N_11460,N_11525);
nand U11749 (N_11749,N_11576,N_11455);
nor U11750 (N_11750,N_11515,N_11510);
nor U11751 (N_11751,N_11529,N_11577);
and U11752 (N_11752,N_11516,N_11529);
nor U11753 (N_11753,N_11561,N_11571);
or U11754 (N_11754,N_11510,N_11540);
or U11755 (N_11755,N_11513,N_11519);
nand U11756 (N_11756,N_11547,N_11471);
nor U11757 (N_11757,N_11562,N_11590);
xor U11758 (N_11758,N_11527,N_11548);
and U11759 (N_11759,N_11421,N_11464);
or U11760 (N_11760,N_11591,N_11553);
nor U11761 (N_11761,N_11558,N_11448);
nor U11762 (N_11762,N_11517,N_11541);
nand U11763 (N_11763,N_11528,N_11578);
and U11764 (N_11764,N_11475,N_11442);
nand U11765 (N_11765,N_11437,N_11406);
xor U11766 (N_11766,N_11470,N_11430);
nor U11767 (N_11767,N_11577,N_11450);
nand U11768 (N_11768,N_11431,N_11469);
and U11769 (N_11769,N_11506,N_11457);
and U11770 (N_11770,N_11450,N_11576);
nand U11771 (N_11771,N_11406,N_11477);
and U11772 (N_11772,N_11584,N_11520);
or U11773 (N_11773,N_11588,N_11481);
nor U11774 (N_11774,N_11458,N_11485);
and U11775 (N_11775,N_11424,N_11505);
nand U11776 (N_11776,N_11440,N_11506);
and U11777 (N_11777,N_11527,N_11453);
nand U11778 (N_11778,N_11525,N_11430);
or U11779 (N_11779,N_11526,N_11446);
nor U11780 (N_11780,N_11422,N_11518);
nand U11781 (N_11781,N_11442,N_11572);
and U11782 (N_11782,N_11448,N_11592);
or U11783 (N_11783,N_11401,N_11476);
and U11784 (N_11784,N_11576,N_11447);
and U11785 (N_11785,N_11576,N_11436);
nand U11786 (N_11786,N_11536,N_11479);
nor U11787 (N_11787,N_11597,N_11516);
nand U11788 (N_11788,N_11494,N_11403);
and U11789 (N_11789,N_11470,N_11584);
and U11790 (N_11790,N_11457,N_11560);
and U11791 (N_11791,N_11583,N_11569);
or U11792 (N_11792,N_11520,N_11509);
or U11793 (N_11793,N_11547,N_11417);
nand U11794 (N_11794,N_11517,N_11593);
nand U11795 (N_11795,N_11515,N_11517);
xnor U11796 (N_11796,N_11505,N_11443);
and U11797 (N_11797,N_11555,N_11490);
or U11798 (N_11798,N_11480,N_11577);
or U11799 (N_11799,N_11518,N_11579);
and U11800 (N_11800,N_11668,N_11787);
or U11801 (N_11801,N_11645,N_11656);
nand U11802 (N_11802,N_11763,N_11608);
nor U11803 (N_11803,N_11664,N_11719);
nand U11804 (N_11804,N_11677,N_11685);
nand U11805 (N_11805,N_11747,N_11646);
and U11806 (N_11806,N_11799,N_11696);
nor U11807 (N_11807,N_11647,N_11607);
or U11808 (N_11808,N_11637,N_11779);
xnor U11809 (N_11809,N_11606,N_11609);
nand U11810 (N_11810,N_11669,N_11644);
nand U11811 (N_11811,N_11755,N_11758);
nor U11812 (N_11812,N_11707,N_11636);
nand U11813 (N_11813,N_11641,N_11643);
or U11814 (N_11814,N_11671,N_11736);
xor U11815 (N_11815,N_11695,N_11732);
nand U11816 (N_11816,N_11735,N_11778);
and U11817 (N_11817,N_11687,N_11675);
or U11818 (N_11818,N_11728,N_11774);
and U11819 (N_11819,N_11704,N_11796);
or U11820 (N_11820,N_11749,N_11793);
nor U11821 (N_11821,N_11753,N_11721);
and U11822 (N_11822,N_11700,N_11653);
and U11823 (N_11823,N_11725,N_11722);
and U11824 (N_11824,N_11631,N_11759);
nor U11825 (N_11825,N_11745,N_11613);
or U11826 (N_11826,N_11738,N_11709);
and U11827 (N_11827,N_11716,N_11605);
nor U11828 (N_11828,N_11640,N_11771);
nand U11829 (N_11829,N_11760,N_11726);
or U11830 (N_11830,N_11672,N_11750);
nand U11831 (N_11831,N_11618,N_11673);
nor U11832 (N_11832,N_11680,N_11619);
or U11833 (N_11833,N_11756,N_11697);
and U11834 (N_11834,N_11784,N_11649);
or U11835 (N_11835,N_11718,N_11625);
or U11836 (N_11836,N_11661,N_11688);
and U11837 (N_11837,N_11676,N_11723);
or U11838 (N_11838,N_11715,N_11648);
or U11839 (N_11839,N_11686,N_11781);
and U11840 (N_11840,N_11727,N_11757);
nor U11841 (N_11841,N_11691,N_11785);
nand U11842 (N_11842,N_11628,N_11772);
and U11843 (N_11843,N_11770,N_11702);
or U11844 (N_11844,N_11602,N_11764);
and U11845 (N_11845,N_11776,N_11737);
nor U11846 (N_11846,N_11730,N_11761);
nor U11847 (N_11847,N_11767,N_11678);
nor U11848 (N_11848,N_11679,N_11655);
nor U11849 (N_11849,N_11794,N_11651);
or U11850 (N_11850,N_11741,N_11711);
nand U11851 (N_11851,N_11751,N_11701);
or U11852 (N_11852,N_11604,N_11621);
nand U11853 (N_11853,N_11720,N_11775);
nand U11854 (N_11854,N_11733,N_11658);
and U11855 (N_11855,N_11638,N_11797);
and U11856 (N_11856,N_11717,N_11791);
nand U11857 (N_11857,N_11690,N_11652);
nand U11858 (N_11858,N_11600,N_11692);
and U11859 (N_11859,N_11780,N_11743);
and U11860 (N_11860,N_11659,N_11705);
nand U11861 (N_11861,N_11616,N_11666);
nand U11862 (N_11862,N_11734,N_11708);
and U11863 (N_11863,N_11682,N_11742);
or U11864 (N_11864,N_11657,N_11792);
or U11865 (N_11865,N_11610,N_11626);
nor U11866 (N_11866,N_11611,N_11615);
nor U11867 (N_11867,N_11773,N_11684);
nor U11868 (N_11868,N_11663,N_11689);
or U11869 (N_11869,N_11748,N_11693);
nor U11870 (N_11870,N_11667,N_11614);
and U11871 (N_11871,N_11782,N_11650);
nand U11872 (N_11872,N_11620,N_11788);
and U11873 (N_11873,N_11729,N_11683);
nor U11874 (N_11874,N_11633,N_11635);
xnor U11875 (N_11875,N_11752,N_11699);
nor U11876 (N_11876,N_11786,N_11713);
nor U11877 (N_11877,N_11739,N_11639);
and U11878 (N_11878,N_11601,N_11740);
nor U11879 (N_11879,N_11710,N_11766);
nor U11880 (N_11880,N_11629,N_11622);
nor U11881 (N_11881,N_11670,N_11762);
or U11882 (N_11882,N_11642,N_11769);
or U11883 (N_11883,N_11694,N_11634);
or U11884 (N_11884,N_11746,N_11765);
nor U11885 (N_11885,N_11706,N_11627);
nand U11886 (N_11886,N_11789,N_11703);
and U11887 (N_11887,N_11698,N_11665);
or U11888 (N_11888,N_11662,N_11783);
or U11889 (N_11889,N_11744,N_11681);
nand U11890 (N_11890,N_11674,N_11660);
and U11891 (N_11891,N_11624,N_11724);
or U11892 (N_11892,N_11714,N_11731);
and U11893 (N_11893,N_11617,N_11768);
and U11894 (N_11894,N_11612,N_11632);
nand U11895 (N_11895,N_11790,N_11630);
or U11896 (N_11896,N_11795,N_11712);
nand U11897 (N_11897,N_11798,N_11603);
nor U11898 (N_11898,N_11654,N_11777);
nand U11899 (N_11899,N_11623,N_11754);
or U11900 (N_11900,N_11698,N_11687);
nand U11901 (N_11901,N_11761,N_11741);
nor U11902 (N_11902,N_11686,N_11696);
or U11903 (N_11903,N_11671,N_11660);
or U11904 (N_11904,N_11690,N_11781);
and U11905 (N_11905,N_11627,N_11762);
nor U11906 (N_11906,N_11712,N_11677);
and U11907 (N_11907,N_11626,N_11799);
or U11908 (N_11908,N_11630,N_11679);
nor U11909 (N_11909,N_11614,N_11700);
or U11910 (N_11910,N_11617,N_11748);
nand U11911 (N_11911,N_11641,N_11781);
and U11912 (N_11912,N_11672,N_11660);
or U11913 (N_11913,N_11702,N_11773);
or U11914 (N_11914,N_11799,N_11688);
nor U11915 (N_11915,N_11765,N_11669);
nor U11916 (N_11916,N_11709,N_11623);
nor U11917 (N_11917,N_11616,N_11685);
and U11918 (N_11918,N_11634,N_11743);
xnor U11919 (N_11919,N_11799,N_11720);
or U11920 (N_11920,N_11795,N_11798);
nand U11921 (N_11921,N_11696,N_11633);
or U11922 (N_11922,N_11724,N_11759);
nand U11923 (N_11923,N_11671,N_11624);
nand U11924 (N_11924,N_11722,N_11708);
and U11925 (N_11925,N_11768,N_11694);
or U11926 (N_11926,N_11616,N_11762);
and U11927 (N_11927,N_11606,N_11723);
nand U11928 (N_11928,N_11734,N_11667);
nand U11929 (N_11929,N_11658,N_11675);
and U11930 (N_11930,N_11653,N_11705);
nor U11931 (N_11931,N_11610,N_11740);
nand U11932 (N_11932,N_11683,N_11766);
and U11933 (N_11933,N_11797,N_11611);
nand U11934 (N_11934,N_11771,N_11751);
nand U11935 (N_11935,N_11742,N_11750);
and U11936 (N_11936,N_11657,N_11624);
nor U11937 (N_11937,N_11698,N_11636);
nor U11938 (N_11938,N_11764,N_11626);
or U11939 (N_11939,N_11657,N_11618);
and U11940 (N_11940,N_11703,N_11601);
nand U11941 (N_11941,N_11738,N_11793);
and U11942 (N_11942,N_11645,N_11644);
nor U11943 (N_11943,N_11796,N_11676);
nand U11944 (N_11944,N_11638,N_11687);
and U11945 (N_11945,N_11799,N_11698);
nand U11946 (N_11946,N_11684,N_11790);
or U11947 (N_11947,N_11619,N_11753);
and U11948 (N_11948,N_11749,N_11683);
and U11949 (N_11949,N_11681,N_11732);
and U11950 (N_11950,N_11603,N_11703);
and U11951 (N_11951,N_11620,N_11732);
nor U11952 (N_11952,N_11742,N_11649);
or U11953 (N_11953,N_11664,N_11735);
or U11954 (N_11954,N_11693,N_11720);
nor U11955 (N_11955,N_11622,N_11762);
and U11956 (N_11956,N_11633,N_11767);
nand U11957 (N_11957,N_11724,N_11715);
nand U11958 (N_11958,N_11793,N_11620);
nand U11959 (N_11959,N_11737,N_11629);
xor U11960 (N_11960,N_11681,N_11609);
and U11961 (N_11961,N_11735,N_11669);
and U11962 (N_11962,N_11718,N_11722);
or U11963 (N_11963,N_11660,N_11788);
or U11964 (N_11964,N_11622,N_11776);
or U11965 (N_11965,N_11798,N_11601);
and U11966 (N_11966,N_11723,N_11669);
xnor U11967 (N_11967,N_11755,N_11767);
nand U11968 (N_11968,N_11702,N_11730);
nor U11969 (N_11969,N_11789,N_11650);
and U11970 (N_11970,N_11724,N_11660);
or U11971 (N_11971,N_11682,N_11679);
or U11972 (N_11972,N_11647,N_11602);
or U11973 (N_11973,N_11781,N_11645);
or U11974 (N_11974,N_11704,N_11688);
or U11975 (N_11975,N_11683,N_11662);
nor U11976 (N_11976,N_11746,N_11767);
or U11977 (N_11977,N_11737,N_11654);
nand U11978 (N_11978,N_11621,N_11664);
or U11979 (N_11979,N_11620,N_11607);
nor U11980 (N_11980,N_11715,N_11729);
and U11981 (N_11981,N_11685,N_11789);
nor U11982 (N_11982,N_11691,N_11675);
and U11983 (N_11983,N_11680,N_11657);
nor U11984 (N_11984,N_11792,N_11607);
or U11985 (N_11985,N_11747,N_11686);
or U11986 (N_11986,N_11788,N_11779);
nand U11987 (N_11987,N_11621,N_11730);
or U11988 (N_11988,N_11772,N_11619);
nand U11989 (N_11989,N_11615,N_11601);
and U11990 (N_11990,N_11718,N_11750);
and U11991 (N_11991,N_11725,N_11767);
and U11992 (N_11992,N_11754,N_11676);
or U11993 (N_11993,N_11701,N_11720);
or U11994 (N_11994,N_11777,N_11731);
and U11995 (N_11995,N_11718,N_11690);
or U11996 (N_11996,N_11636,N_11769);
nor U11997 (N_11997,N_11797,N_11635);
and U11998 (N_11998,N_11602,N_11796);
or U11999 (N_11999,N_11781,N_11653);
nand U12000 (N_12000,N_11899,N_11877);
nand U12001 (N_12001,N_11818,N_11919);
nand U12002 (N_12002,N_11986,N_11883);
and U12003 (N_12003,N_11849,N_11825);
nand U12004 (N_12004,N_11844,N_11816);
nor U12005 (N_12005,N_11856,N_11966);
nor U12006 (N_12006,N_11937,N_11840);
nand U12007 (N_12007,N_11851,N_11916);
and U12008 (N_12008,N_11805,N_11829);
and U12009 (N_12009,N_11869,N_11972);
or U12010 (N_12010,N_11803,N_11957);
nand U12011 (N_12011,N_11936,N_11900);
nand U12012 (N_12012,N_11804,N_11971);
nor U12013 (N_12013,N_11978,N_11962);
and U12014 (N_12014,N_11931,N_11864);
nor U12015 (N_12015,N_11817,N_11996);
nand U12016 (N_12016,N_11963,N_11858);
or U12017 (N_12017,N_11903,N_11874);
nand U12018 (N_12018,N_11905,N_11822);
or U12019 (N_12019,N_11909,N_11802);
or U12020 (N_12020,N_11800,N_11940);
nor U12021 (N_12021,N_11892,N_11912);
or U12022 (N_12022,N_11974,N_11867);
nor U12023 (N_12023,N_11923,N_11980);
nand U12024 (N_12024,N_11891,N_11847);
and U12025 (N_12025,N_11993,N_11872);
nor U12026 (N_12026,N_11941,N_11991);
and U12027 (N_12027,N_11808,N_11806);
nand U12028 (N_12028,N_11970,N_11944);
nand U12029 (N_12029,N_11914,N_11890);
and U12030 (N_12030,N_11838,N_11910);
or U12031 (N_12031,N_11913,N_11967);
and U12032 (N_12032,N_11871,N_11860);
nor U12033 (N_12033,N_11911,N_11995);
and U12034 (N_12034,N_11834,N_11807);
and U12035 (N_12035,N_11870,N_11981);
nand U12036 (N_12036,N_11956,N_11947);
nor U12037 (N_12037,N_11935,N_11875);
nor U12038 (N_12038,N_11907,N_11828);
and U12039 (N_12039,N_11975,N_11898);
or U12040 (N_12040,N_11813,N_11976);
and U12041 (N_12041,N_11921,N_11924);
and U12042 (N_12042,N_11876,N_11879);
nand U12043 (N_12043,N_11925,N_11964);
and U12044 (N_12044,N_11836,N_11953);
or U12045 (N_12045,N_11901,N_11873);
nand U12046 (N_12046,N_11987,N_11998);
nor U12047 (N_12047,N_11897,N_11843);
nand U12048 (N_12048,N_11983,N_11889);
or U12049 (N_12049,N_11908,N_11952);
or U12050 (N_12050,N_11832,N_11917);
and U12051 (N_12051,N_11853,N_11968);
nor U12052 (N_12052,N_11943,N_11933);
and U12053 (N_12053,N_11865,N_11927);
nand U12054 (N_12054,N_11812,N_11922);
nand U12055 (N_12055,N_11868,N_11918);
nor U12056 (N_12056,N_11842,N_11939);
or U12057 (N_12057,N_11824,N_11886);
nand U12058 (N_12058,N_11835,N_11882);
or U12059 (N_12059,N_11961,N_11948);
and U12060 (N_12060,N_11820,N_11887);
nor U12061 (N_12061,N_11814,N_11997);
nor U12062 (N_12062,N_11945,N_11878);
and U12063 (N_12063,N_11982,N_11973);
or U12064 (N_12064,N_11926,N_11984);
or U12065 (N_12065,N_11992,N_11809);
nand U12066 (N_12066,N_11942,N_11801);
nand U12067 (N_12067,N_11958,N_11896);
or U12068 (N_12068,N_11938,N_11920);
nand U12069 (N_12069,N_11852,N_11930);
nor U12070 (N_12070,N_11946,N_11932);
nor U12071 (N_12071,N_11960,N_11859);
nand U12072 (N_12072,N_11949,N_11977);
nand U12073 (N_12073,N_11857,N_11846);
nor U12074 (N_12074,N_11885,N_11810);
nand U12075 (N_12075,N_11934,N_11884);
nor U12076 (N_12076,N_11850,N_11950);
nor U12077 (N_12077,N_11951,N_11862);
nand U12078 (N_12078,N_11861,N_11881);
nor U12079 (N_12079,N_11830,N_11904);
nand U12080 (N_12080,N_11988,N_11831);
nor U12081 (N_12081,N_11815,N_11863);
or U12082 (N_12082,N_11839,N_11969);
and U12083 (N_12083,N_11965,N_11979);
and U12084 (N_12084,N_11894,N_11902);
or U12085 (N_12085,N_11915,N_11827);
nor U12086 (N_12086,N_11888,N_11985);
or U12087 (N_12087,N_11855,N_11841);
or U12088 (N_12088,N_11866,N_11811);
nor U12089 (N_12089,N_11928,N_11989);
or U12090 (N_12090,N_11848,N_11837);
and U12091 (N_12091,N_11906,N_11955);
nand U12092 (N_12092,N_11826,N_11895);
or U12093 (N_12093,N_11990,N_11819);
nor U12094 (N_12094,N_11954,N_11845);
nor U12095 (N_12095,N_11893,N_11959);
or U12096 (N_12096,N_11854,N_11821);
and U12097 (N_12097,N_11999,N_11823);
nand U12098 (N_12098,N_11929,N_11833);
nor U12099 (N_12099,N_11880,N_11994);
nor U12100 (N_12100,N_11803,N_11842);
or U12101 (N_12101,N_11930,N_11921);
nor U12102 (N_12102,N_11825,N_11882);
and U12103 (N_12103,N_11901,N_11911);
nand U12104 (N_12104,N_11881,N_11959);
or U12105 (N_12105,N_11855,N_11808);
or U12106 (N_12106,N_11965,N_11824);
or U12107 (N_12107,N_11964,N_11913);
and U12108 (N_12108,N_11983,N_11903);
or U12109 (N_12109,N_11965,N_11954);
nand U12110 (N_12110,N_11837,N_11802);
or U12111 (N_12111,N_11885,N_11845);
and U12112 (N_12112,N_11949,N_11966);
nand U12113 (N_12113,N_11853,N_11826);
nand U12114 (N_12114,N_11859,N_11838);
or U12115 (N_12115,N_11887,N_11808);
nand U12116 (N_12116,N_11854,N_11954);
nor U12117 (N_12117,N_11997,N_11867);
nor U12118 (N_12118,N_11918,N_11963);
nor U12119 (N_12119,N_11996,N_11836);
nand U12120 (N_12120,N_11895,N_11861);
nor U12121 (N_12121,N_11834,N_11983);
or U12122 (N_12122,N_11833,N_11850);
and U12123 (N_12123,N_11908,N_11898);
and U12124 (N_12124,N_11800,N_11888);
and U12125 (N_12125,N_11939,N_11941);
nand U12126 (N_12126,N_11941,N_11972);
nor U12127 (N_12127,N_11948,N_11835);
nor U12128 (N_12128,N_11992,N_11916);
nand U12129 (N_12129,N_11933,N_11970);
or U12130 (N_12130,N_11902,N_11931);
nor U12131 (N_12131,N_11901,N_11977);
and U12132 (N_12132,N_11993,N_11966);
nand U12133 (N_12133,N_11911,N_11875);
or U12134 (N_12134,N_11964,N_11930);
nand U12135 (N_12135,N_11806,N_11969);
nand U12136 (N_12136,N_11939,N_11873);
nor U12137 (N_12137,N_11959,N_11932);
nand U12138 (N_12138,N_11952,N_11937);
and U12139 (N_12139,N_11872,N_11844);
nand U12140 (N_12140,N_11932,N_11912);
nor U12141 (N_12141,N_11954,N_11941);
nand U12142 (N_12142,N_11893,N_11875);
nor U12143 (N_12143,N_11990,N_11982);
or U12144 (N_12144,N_11997,N_11801);
nor U12145 (N_12145,N_11894,N_11827);
and U12146 (N_12146,N_11827,N_11949);
nand U12147 (N_12147,N_11820,N_11867);
nand U12148 (N_12148,N_11924,N_11865);
nand U12149 (N_12149,N_11807,N_11931);
and U12150 (N_12150,N_11918,N_11855);
nand U12151 (N_12151,N_11869,N_11996);
or U12152 (N_12152,N_11850,N_11854);
nor U12153 (N_12153,N_11800,N_11873);
and U12154 (N_12154,N_11910,N_11861);
nor U12155 (N_12155,N_11902,N_11991);
and U12156 (N_12156,N_11908,N_11976);
and U12157 (N_12157,N_11941,N_11886);
nor U12158 (N_12158,N_11960,N_11996);
or U12159 (N_12159,N_11894,N_11955);
nand U12160 (N_12160,N_11801,N_11884);
nand U12161 (N_12161,N_11885,N_11866);
or U12162 (N_12162,N_11988,N_11930);
and U12163 (N_12163,N_11998,N_11985);
and U12164 (N_12164,N_11981,N_11942);
nand U12165 (N_12165,N_11945,N_11992);
nand U12166 (N_12166,N_11881,N_11830);
or U12167 (N_12167,N_11932,N_11858);
or U12168 (N_12168,N_11926,N_11881);
nand U12169 (N_12169,N_11832,N_11847);
or U12170 (N_12170,N_11868,N_11953);
and U12171 (N_12171,N_11976,N_11994);
nor U12172 (N_12172,N_11911,N_11824);
and U12173 (N_12173,N_11914,N_11821);
nand U12174 (N_12174,N_11944,N_11810);
nand U12175 (N_12175,N_11977,N_11945);
nand U12176 (N_12176,N_11914,N_11826);
nor U12177 (N_12177,N_11833,N_11901);
nor U12178 (N_12178,N_11901,N_11957);
nor U12179 (N_12179,N_11811,N_11991);
or U12180 (N_12180,N_11931,N_11814);
nand U12181 (N_12181,N_11836,N_11947);
nand U12182 (N_12182,N_11986,N_11992);
nor U12183 (N_12183,N_11990,N_11888);
nand U12184 (N_12184,N_11888,N_11930);
nor U12185 (N_12185,N_11982,N_11857);
or U12186 (N_12186,N_11825,N_11957);
and U12187 (N_12187,N_11926,N_11979);
nor U12188 (N_12188,N_11913,N_11997);
nor U12189 (N_12189,N_11996,N_11884);
nand U12190 (N_12190,N_11807,N_11819);
nor U12191 (N_12191,N_11816,N_11857);
nand U12192 (N_12192,N_11894,N_11948);
nand U12193 (N_12193,N_11967,N_11844);
and U12194 (N_12194,N_11831,N_11971);
and U12195 (N_12195,N_11949,N_11988);
nor U12196 (N_12196,N_11971,N_11937);
nand U12197 (N_12197,N_11988,N_11868);
or U12198 (N_12198,N_11937,N_11861);
and U12199 (N_12199,N_11944,N_11886);
or U12200 (N_12200,N_12038,N_12076);
xnor U12201 (N_12201,N_12131,N_12125);
nand U12202 (N_12202,N_12100,N_12087);
or U12203 (N_12203,N_12024,N_12023);
nor U12204 (N_12204,N_12107,N_12173);
nor U12205 (N_12205,N_12090,N_12036);
or U12206 (N_12206,N_12055,N_12190);
and U12207 (N_12207,N_12033,N_12058);
and U12208 (N_12208,N_12109,N_12150);
nor U12209 (N_12209,N_12022,N_12017);
or U12210 (N_12210,N_12050,N_12132);
or U12211 (N_12211,N_12148,N_12097);
and U12212 (N_12212,N_12045,N_12041);
nor U12213 (N_12213,N_12053,N_12069);
or U12214 (N_12214,N_12077,N_12199);
or U12215 (N_12215,N_12164,N_12152);
nor U12216 (N_12216,N_12191,N_12016);
nand U12217 (N_12217,N_12003,N_12143);
and U12218 (N_12218,N_12001,N_12151);
and U12219 (N_12219,N_12138,N_12079);
or U12220 (N_12220,N_12176,N_12096);
nor U12221 (N_12221,N_12064,N_12091);
nor U12222 (N_12222,N_12026,N_12130);
and U12223 (N_12223,N_12065,N_12184);
nand U12224 (N_12224,N_12140,N_12012);
and U12225 (N_12225,N_12000,N_12004);
nor U12226 (N_12226,N_12035,N_12052);
or U12227 (N_12227,N_12080,N_12127);
and U12228 (N_12228,N_12057,N_12128);
xnor U12229 (N_12229,N_12048,N_12155);
nor U12230 (N_12230,N_12037,N_12175);
or U12231 (N_12231,N_12161,N_12174);
nor U12232 (N_12232,N_12018,N_12020);
and U12233 (N_12233,N_12185,N_12123);
nor U12234 (N_12234,N_12154,N_12193);
nor U12235 (N_12235,N_12031,N_12168);
nor U12236 (N_12236,N_12046,N_12169);
and U12237 (N_12237,N_12039,N_12139);
or U12238 (N_12238,N_12124,N_12092);
and U12239 (N_12239,N_12089,N_12186);
or U12240 (N_12240,N_12112,N_12141);
and U12241 (N_12241,N_12074,N_12145);
nor U12242 (N_12242,N_12044,N_12054);
xnor U12243 (N_12243,N_12178,N_12059);
and U12244 (N_12244,N_12021,N_12180);
or U12245 (N_12245,N_12116,N_12095);
nand U12246 (N_12246,N_12117,N_12042);
or U12247 (N_12247,N_12113,N_12027);
or U12248 (N_12248,N_12170,N_12196);
or U12249 (N_12249,N_12149,N_12120);
or U12250 (N_12250,N_12106,N_12158);
and U12251 (N_12251,N_12034,N_12085);
xor U12252 (N_12252,N_12111,N_12072);
and U12253 (N_12253,N_12093,N_12133);
nand U12254 (N_12254,N_12002,N_12153);
or U12255 (N_12255,N_12105,N_12009);
and U12256 (N_12256,N_12011,N_12066);
nor U12257 (N_12257,N_12094,N_12115);
nor U12258 (N_12258,N_12192,N_12137);
and U12259 (N_12259,N_12010,N_12099);
nand U12260 (N_12260,N_12049,N_12081);
and U12261 (N_12261,N_12082,N_12062);
nand U12262 (N_12262,N_12068,N_12088);
nand U12263 (N_12263,N_12156,N_12135);
or U12264 (N_12264,N_12121,N_12028);
nand U12265 (N_12265,N_12056,N_12043);
nor U12266 (N_12266,N_12103,N_12104);
and U12267 (N_12267,N_12146,N_12015);
and U12268 (N_12268,N_12040,N_12070);
or U12269 (N_12269,N_12166,N_12025);
nand U12270 (N_12270,N_12014,N_12047);
and U12271 (N_12271,N_12144,N_12182);
nand U12272 (N_12272,N_12147,N_12060);
and U12273 (N_12273,N_12084,N_12063);
nand U12274 (N_12274,N_12061,N_12172);
nand U12275 (N_12275,N_12118,N_12075);
nor U12276 (N_12276,N_12013,N_12167);
or U12277 (N_12277,N_12181,N_12189);
nand U12278 (N_12278,N_12194,N_12160);
nor U12279 (N_12279,N_12171,N_12126);
nand U12280 (N_12280,N_12083,N_12198);
and U12281 (N_12281,N_12098,N_12188);
nor U12282 (N_12282,N_12162,N_12159);
and U12283 (N_12283,N_12108,N_12032);
and U12284 (N_12284,N_12163,N_12129);
or U12285 (N_12285,N_12187,N_12177);
nand U12286 (N_12286,N_12114,N_12136);
and U12287 (N_12287,N_12134,N_12197);
nor U12288 (N_12288,N_12086,N_12030);
nor U12289 (N_12289,N_12165,N_12183);
and U12290 (N_12290,N_12101,N_12005);
nand U12291 (N_12291,N_12110,N_12122);
nor U12292 (N_12292,N_12102,N_12071);
or U12293 (N_12293,N_12078,N_12195);
and U12294 (N_12294,N_12029,N_12073);
or U12295 (N_12295,N_12142,N_12006);
nor U12296 (N_12296,N_12008,N_12119);
nor U12297 (N_12297,N_12051,N_12157);
nor U12298 (N_12298,N_12019,N_12007);
nand U12299 (N_12299,N_12179,N_12067);
and U12300 (N_12300,N_12144,N_12085);
nand U12301 (N_12301,N_12138,N_12038);
and U12302 (N_12302,N_12086,N_12198);
and U12303 (N_12303,N_12056,N_12196);
or U12304 (N_12304,N_12004,N_12129);
nor U12305 (N_12305,N_12080,N_12173);
nand U12306 (N_12306,N_12103,N_12182);
or U12307 (N_12307,N_12054,N_12015);
and U12308 (N_12308,N_12183,N_12167);
or U12309 (N_12309,N_12193,N_12134);
or U12310 (N_12310,N_12131,N_12030);
and U12311 (N_12311,N_12046,N_12104);
and U12312 (N_12312,N_12026,N_12014);
nand U12313 (N_12313,N_12041,N_12173);
nand U12314 (N_12314,N_12122,N_12124);
nand U12315 (N_12315,N_12186,N_12163);
and U12316 (N_12316,N_12006,N_12117);
or U12317 (N_12317,N_12054,N_12080);
or U12318 (N_12318,N_12054,N_12066);
and U12319 (N_12319,N_12034,N_12022);
or U12320 (N_12320,N_12162,N_12120);
nor U12321 (N_12321,N_12136,N_12145);
or U12322 (N_12322,N_12116,N_12001);
xnor U12323 (N_12323,N_12173,N_12032);
or U12324 (N_12324,N_12170,N_12055);
nand U12325 (N_12325,N_12089,N_12190);
and U12326 (N_12326,N_12142,N_12181);
and U12327 (N_12327,N_12133,N_12142);
nor U12328 (N_12328,N_12127,N_12171);
nor U12329 (N_12329,N_12187,N_12097);
nor U12330 (N_12330,N_12109,N_12039);
nand U12331 (N_12331,N_12173,N_12003);
nor U12332 (N_12332,N_12010,N_12093);
and U12333 (N_12333,N_12188,N_12159);
or U12334 (N_12334,N_12035,N_12194);
or U12335 (N_12335,N_12116,N_12174);
nor U12336 (N_12336,N_12070,N_12169);
and U12337 (N_12337,N_12106,N_12136);
nor U12338 (N_12338,N_12023,N_12142);
and U12339 (N_12339,N_12187,N_12111);
or U12340 (N_12340,N_12112,N_12198);
nor U12341 (N_12341,N_12182,N_12079);
xnor U12342 (N_12342,N_12028,N_12072);
nor U12343 (N_12343,N_12140,N_12064);
nand U12344 (N_12344,N_12082,N_12075);
nand U12345 (N_12345,N_12174,N_12114);
nand U12346 (N_12346,N_12014,N_12156);
and U12347 (N_12347,N_12079,N_12185);
nor U12348 (N_12348,N_12089,N_12007);
nor U12349 (N_12349,N_12067,N_12099);
nor U12350 (N_12350,N_12030,N_12062);
or U12351 (N_12351,N_12006,N_12146);
or U12352 (N_12352,N_12123,N_12156);
nor U12353 (N_12353,N_12167,N_12106);
nand U12354 (N_12354,N_12020,N_12127);
and U12355 (N_12355,N_12188,N_12068);
nand U12356 (N_12356,N_12059,N_12092);
nor U12357 (N_12357,N_12029,N_12066);
and U12358 (N_12358,N_12037,N_12188);
nor U12359 (N_12359,N_12144,N_12186);
nor U12360 (N_12360,N_12170,N_12005);
and U12361 (N_12361,N_12144,N_12155);
and U12362 (N_12362,N_12007,N_12198);
or U12363 (N_12363,N_12016,N_12177);
or U12364 (N_12364,N_12176,N_12141);
nor U12365 (N_12365,N_12131,N_12081);
and U12366 (N_12366,N_12053,N_12073);
nand U12367 (N_12367,N_12016,N_12136);
nand U12368 (N_12368,N_12151,N_12041);
and U12369 (N_12369,N_12015,N_12040);
nand U12370 (N_12370,N_12065,N_12176);
nor U12371 (N_12371,N_12121,N_12188);
and U12372 (N_12372,N_12199,N_12184);
nand U12373 (N_12373,N_12154,N_12114);
nand U12374 (N_12374,N_12043,N_12155);
or U12375 (N_12375,N_12008,N_12073);
nor U12376 (N_12376,N_12131,N_12072);
nor U12377 (N_12377,N_12026,N_12028);
and U12378 (N_12378,N_12070,N_12097);
nand U12379 (N_12379,N_12099,N_12088);
nor U12380 (N_12380,N_12038,N_12026);
nor U12381 (N_12381,N_12022,N_12089);
and U12382 (N_12382,N_12036,N_12007);
nand U12383 (N_12383,N_12160,N_12168);
nand U12384 (N_12384,N_12062,N_12047);
or U12385 (N_12385,N_12194,N_12112);
or U12386 (N_12386,N_12103,N_12088);
or U12387 (N_12387,N_12132,N_12098);
and U12388 (N_12388,N_12175,N_12009);
or U12389 (N_12389,N_12154,N_12146);
or U12390 (N_12390,N_12028,N_12019);
and U12391 (N_12391,N_12006,N_12046);
or U12392 (N_12392,N_12086,N_12053);
and U12393 (N_12393,N_12002,N_12063);
nand U12394 (N_12394,N_12046,N_12013);
or U12395 (N_12395,N_12134,N_12028);
and U12396 (N_12396,N_12055,N_12107);
and U12397 (N_12397,N_12078,N_12016);
and U12398 (N_12398,N_12065,N_12067);
nand U12399 (N_12399,N_12120,N_12176);
and U12400 (N_12400,N_12376,N_12200);
and U12401 (N_12401,N_12352,N_12342);
or U12402 (N_12402,N_12320,N_12222);
or U12403 (N_12403,N_12284,N_12365);
nor U12404 (N_12404,N_12211,N_12242);
nor U12405 (N_12405,N_12304,N_12287);
nand U12406 (N_12406,N_12339,N_12371);
nand U12407 (N_12407,N_12384,N_12321);
nor U12408 (N_12408,N_12363,N_12368);
nor U12409 (N_12409,N_12316,N_12399);
nand U12410 (N_12410,N_12398,N_12219);
nor U12411 (N_12411,N_12341,N_12361);
or U12412 (N_12412,N_12360,N_12292);
or U12413 (N_12413,N_12250,N_12216);
nor U12414 (N_12414,N_12346,N_12370);
nor U12415 (N_12415,N_12227,N_12230);
nor U12416 (N_12416,N_12301,N_12327);
and U12417 (N_12417,N_12322,N_12273);
nand U12418 (N_12418,N_12381,N_12239);
or U12419 (N_12419,N_12336,N_12276);
and U12420 (N_12420,N_12373,N_12272);
nand U12421 (N_12421,N_12204,N_12326);
or U12422 (N_12422,N_12282,N_12274);
or U12423 (N_12423,N_12313,N_12245);
and U12424 (N_12424,N_12234,N_12331);
nand U12425 (N_12425,N_12309,N_12306);
or U12426 (N_12426,N_12201,N_12241);
nand U12427 (N_12427,N_12218,N_12357);
or U12428 (N_12428,N_12355,N_12213);
nand U12429 (N_12429,N_12302,N_12236);
nor U12430 (N_12430,N_12291,N_12344);
nand U12431 (N_12431,N_12228,N_12212);
or U12432 (N_12432,N_12244,N_12252);
xor U12433 (N_12433,N_12297,N_12369);
nand U12434 (N_12434,N_12307,N_12392);
or U12435 (N_12435,N_12268,N_12257);
and U12436 (N_12436,N_12286,N_12259);
or U12437 (N_12437,N_12329,N_12240);
and U12438 (N_12438,N_12206,N_12229);
nand U12439 (N_12439,N_12217,N_12289);
and U12440 (N_12440,N_12308,N_12378);
nand U12441 (N_12441,N_12258,N_12347);
nand U12442 (N_12442,N_12303,N_12374);
nand U12443 (N_12443,N_12299,N_12300);
nor U12444 (N_12444,N_12350,N_12295);
nand U12445 (N_12445,N_12263,N_12260);
or U12446 (N_12446,N_12251,N_12288);
and U12447 (N_12447,N_12215,N_12281);
or U12448 (N_12448,N_12262,N_12305);
or U12449 (N_12449,N_12293,N_12277);
or U12450 (N_12450,N_12235,N_12319);
and U12451 (N_12451,N_12314,N_12380);
nand U12452 (N_12452,N_12310,N_12337);
and U12453 (N_12453,N_12395,N_12279);
nand U12454 (N_12454,N_12203,N_12270);
and U12455 (N_12455,N_12285,N_12385);
and U12456 (N_12456,N_12375,N_12311);
nand U12457 (N_12457,N_12328,N_12283);
and U12458 (N_12458,N_12358,N_12233);
and U12459 (N_12459,N_12231,N_12220);
and U12460 (N_12460,N_12394,N_12296);
or U12461 (N_12461,N_12338,N_12225);
nor U12462 (N_12462,N_12208,N_12332);
nand U12463 (N_12463,N_12278,N_12366);
and U12464 (N_12464,N_12334,N_12249);
nor U12465 (N_12465,N_12367,N_12343);
or U12466 (N_12466,N_12386,N_12214);
and U12467 (N_12467,N_12391,N_12317);
and U12468 (N_12468,N_12324,N_12261);
nor U12469 (N_12469,N_12377,N_12359);
and U12470 (N_12470,N_12248,N_12271);
or U12471 (N_12471,N_12335,N_12330);
and U12472 (N_12472,N_12246,N_12362);
nor U12473 (N_12473,N_12387,N_12353);
and U12474 (N_12474,N_12390,N_12221);
and U12475 (N_12475,N_12224,N_12318);
nand U12476 (N_12476,N_12372,N_12253);
and U12477 (N_12477,N_12382,N_12243);
xnor U12478 (N_12478,N_12348,N_12210);
nor U12479 (N_12479,N_12267,N_12205);
nand U12480 (N_12480,N_12209,N_12379);
and U12481 (N_12481,N_12255,N_12333);
nor U12482 (N_12482,N_12290,N_12254);
or U12483 (N_12483,N_12354,N_12265);
and U12484 (N_12484,N_12232,N_12280);
nand U12485 (N_12485,N_12389,N_12393);
and U12486 (N_12486,N_12238,N_12323);
or U12487 (N_12487,N_12340,N_12207);
nand U12488 (N_12488,N_12298,N_12345);
or U12489 (N_12489,N_12315,N_12356);
and U12490 (N_12490,N_12266,N_12223);
and U12491 (N_12491,N_12294,N_12269);
and U12492 (N_12492,N_12256,N_12312);
nor U12493 (N_12493,N_12264,N_12349);
nand U12494 (N_12494,N_12351,N_12396);
nor U12495 (N_12495,N_12388,N_12202);
and U12496 (N_12496,N_12325,N_12397);
nand U12497 (N_12497,N_12247,N_12364);
and U12498 (N_12498,N_12383,N_12226);
and U12499 (N_12499,N_12237,N_12275);
nor U12500 (N_12500,N_12357,N_12321);
and U12501 (N_12501,N_12258,N_12311);
and U12502 (N_12502,N_12257,N_12362);
or U12503 (N_12503,N_12320,N_12332);
and U12504 (N_12504,N_12264,N_12302);
and U12505 (N_12505,N_12246,N_12351);
and U12506 (N_12506,N_12268,N_12338);
or U12507 (N_12507,N_12243,N_12383);
nor U12508 (N_12508,N_12358,N_12396);
nor U12509 (N_12509,N_12291,N_12326);
nand U12510 (N_12510,N_12218,N_12337);
nor U12511 (N_12511,N_12332,N_12260);
or U12512 (N_12512,N_12379,N_12362);
nor U12513 (N_12513,N_12349,N_12304);
xnor U12514 (N_12514,N_12254,N_12267);
and U12515 (N_12515,N_12338,N_12310);
and U12516 (N_12516,N_12363,N_12200);
nor U12517 (N_12517,N_12224,N_12337);
or U12518 (N_12518,N_12303,N_12379);
nor U12519 (N_12519,N_12354,N_12324);
and U12520 (N_12520,N_12258,N_12355);
and U12521 (N_12521,N_12297,N_12357);
nor U12522 (N_12522,N_12291,N_12246);
or U12523 (N_12523,N_12292,N_12395);
nor U12524 (N_12524,N_12356,N_12317);
nand U12525 (N_12525,N_12368,N_12289);
and U12526 (N_12526,N_12277,N_12377);
and U12527 (N_12527,N_12237,N_12244);
and U12528 (N_12528,N_12339,N_12391);
and U12529 (N_12529,N_12210,N_12315);
nor U12530 (N_12530,N_12213,N_12284);
and U12531 (N_12531,N_12300,N_12339);
and U12532 (N_12532,N_12219,N_12380);
nand U12533 (N_12533,N_12369,N_12280);
or U12534 (N_12534,N_12359,N_12331);
or U12535 (N_12535,N_12228,N_12285);
nand U12536 (N_12536,N_12370,N_12375);
nand U12537 (N_12537,N_12397,N_12381);
and U12538 (N_12538,N_12219,N_12228);
nand U12539 (N_12539,N_12382,N_12252);
nand U12540 (N_12540,N_12225,N_12213);
or U12541 (N_12541,N_12394,N_12253);
nor U12542 (N_12542,N_12269,N_12226);
or U12543 (N_12543,N_12375,N_12323);
and U12544 (N_12544,N_12252,N_12320);
or U12545 (N_12545,N_12396,N_12278);
and U12546 (N_12546,N_12311,N_12255);
nand U12547 (N_12547,N_12393,N_12331);
nor U12548 (N_12548,N_12222,N_12325);
nor U12549 (N_12549,N_12377,N_12210);
and U12550 (N_12550,N_12379,N_12276);
nor U12551 (N_12551,N_12221,N_12378);
nor U12552 (N_12552,N_12309,N_12216);
or U12553 (N_12553,N_12257,N_12343);
nand U12554 (N_12554,N_12244,N_12239);
nand U12555 (N_12555,N_12354,N_12339);
nor U12556 (N_12556,N_12307,N_12204);
nor U12557 (N_12557,N_12365,N_12213);
nor U12558 (N_12558,N_12229,N_12307);
nor U12559 (N_12559,N_12234,N_12219);
and U12560 (N_12560,N_12380,N_12215);
or U12561 (N_12561,N_12370,N_12308);
or U12562 (N_12562,N_12372,N_12369);
and U12563 (N_12563,N_12284,N_12232);
and U12564 (N_12564,N_12346,N_12369);
or U12565 (N_12565,N_12398,N_12200);
nand U12566 (N_12566,N_12258,N_12245);
nand U12567 (N_12567,N_12306,N_12245);
nand U12568 (N_12568,N_12375,N_12398);
and U12569 (N_12569,N_12227,N_12326);
nor U12570 (N_12570,N_12234,N_12264);
nand U12571 (N_12571,N_12336,N_12288);
and U12572 (N_12572,N_12351,N_12271);
nand U12573 (N_12573,N_12335,N_12217);
or U12574 (N_12574,N_12278,N_12298);
or U12575 (N_12575,N_12253,N_12304);
nand U12576 (N_12576,N_12212,N_12323);
or U12577 (N_12577,N_12279,N_12337);
or U12578 (N_12578,N_12225,N_12380);
nor U12579 (N_12579,N_12386,N_12305);
nand U12580 (N_12580,N_12377,N_12296);
or U12581 (N_12581,N_12341,N_12366);
or U12582 (N_12582,N_12384,N_12333);
nor U12583 (N_12583,N_12381,N_12309);
nor U12584 (N_12584,N_12223,N_12210);
or U12585 (N_12585,N_12370,N_12334);
nor U12586 (N_12586,N_12367,N_12385);
nor U12587 (N_12587,N_12279,N_12357);
nand U12588 (N_12588,N_12370,N_12270);
nand U12589 (N_12589,N_12312,N_12232);
and U12590 (N_12590,N_12295,N_12340);
and U12591 (N_12591,N_12358,N_12280);
or U12592 (N_12592,N_12263,N_12334);
nand U12593 (N_12593,N_12312,N_12340);
nor U12594 (N_12594,N_12200,N_12207);
or U12595 (N_12595,N_12389,N_12321);
nand U12596 (N_12596,N_12345,N_12376);
and U12597 (N_12597,N_12240,N_12334);
nor U12598 (N_12598,N_12224,N_12331);
nor U12599 (N_12599,N_12285,N_12384);
nor U12600 (N_12600,N_12578,N_12492);
and U12601 (N_12601,N_12580,N_12547);
and U12602 (N_12602,N_12466,N_12416);
and U12603 (N_12603,N_12400,N_12403);
or U12604 (N_12604,N_12455,N_12420);
or U12605 (N_12605,N_12444,N_12512);
and U12606 (N_12606,N_12405,N_12402);
nand U12607 (N_12607,N_12484,N_12513);
nor U12608 (N_12608,N_12517,N_12510);
and U12609 (N_12609,N_12429,N_12551);
nor U12610 (N_12610,N_12490,N_12496);
or U12611 (N_12611,N_12459,N_12417);
nand U12612 (N_12612,N_12414,N_12533);
or U12613 (N_12613,N_12478,N_12558);
nand U12614 (N_12614,N_12505,N_12434);
and U12615 (N_12615,N_12410,N_12452);
nand U12616 (N_12616,N_12531,N_12438);
and U12617 (N_12617,N_12524,N_12441);
nand U12618 (N_12618,N_12593,N_12457);
or U12619 (N_12619,N_12515,N_12427);
nand U12620 (N_12620,N_12463,N_12440);
and U12621 (N_12621,N_12494,N_12585);
and U12622 (N_12622,N_12552,N_12568);
and U12623 (N_12623,N_12406,N_12514);
nor U12624 (N_12624,N_12480,N_12421);
nor U12625 (N_12625,N_12520,N_12453);
or U12626 (N_12626,N_12493,N_12486);
and U12627 (N_12627,N_12556,N_12595);
and U12628 (N_12628,N_12566,N_12415);
nor U12629 (N_12629,N_12504,N_12541);
nor U12630 (N_12630,N_12565,N_12535);
and U12631 (N_12631,N_12407,N_12481);
or U12632 (N_12632,N_12584,N_12599);
nor U12633 (N_12633,N_12491,N_12590);
and U12634 (N_12634,N_12561,N_12454);
nand U12635 (N_12635,N_12469,N_12526);
and U12636 (N_12636,N_12460,N_12579);
nand U12637 (N_12637,N_12525,N_12462);
nand U12638 (N_12638,N_12522,N_12464);
nor U12639 (N_12639,N_12408,N_12472);
nand U12640 (N_12640,N_12476,N_12428);
or U12641 (N_12641,N_12422,N_12511);
nand U12642 (N_12642,N_12439,N_12508);
nor U12643 (N_12643,N_12479,N_12569);
nand U12644 (N_12644,N_12557,N_12487);
nand U12645 (N_12645,N_12448,N_12501);
nor U12646 (N_12646,N_12443,N_12560);
or U12647 (N_12647,N_12468,N_12587);
nand U12648 (N_12648,N_12530,N_12594);
or U12649 (N_12649,N_12550,N_12485);
or U12650 (N_12650,N_12586,N_12446);
or U12651 (N_12651,N_12528,N_12553);
nor U12652 (N_12652,N_12461,N_12555);
and U12653 (N_12653,N_12426,N_12497);
nor U12654 (N_12654,N_12518,N_12475);
and U12655 (N_12655,N_12499,N_12544);
or U12656 (N_12656,N_12581,N_12467);
nor U12657 (N_12657,N_12498,N_12419);
or U12658 (N_12658,N_12506,N_12564);
nand U12659 (N_12659,N_12473,N_12483);
and U12660 (N_12660,N_12529,N_12567);
or U12661 (N_12661,N_12409,N_12554);
or U12662 (N_12662,N_12534,N_12575);
and U12663 (N_12663,N_12401,N_12542);
or U12664 (N_12664,N_12532,N_12503);
nand U12665 (N_12665,N_12516,N_12500);
or U12666 (N_12666,N_12436,N_12451);
nor U12667 (N_12667,N_12482,N_12536);
or U12668 (N_12668,N_12582,N_12591);
nor U12669 (N_12669,N_12432,N_12573);
or U12670 (N_12670,N_12540,N_12539);
nor U12671 (N_12671,N_12488,N_12447);
and U12672 (N_12672,N_12430,N_12502);
or U12673 (N_12673,N_12458,N_12576);
and U12674 (N_12674,N_12456,N_12477);
nand U12675 (N_12675,N_12588,N_12570);
or U12676 (N_12676,N_12549,N_12411);
and U12677 (N_12677,N_12418,N_12465);
and U12678 (N_12678,N_12495,N_12589);
or U12679 (N_12679,N_12519,N_12538);
or U12680 (N_12680,N_12489,N_12435);
and U12681 (N_12681,N_12424,N_12425);
nor U12682 (N_12682,N_12413,N_12537);
nand U12683 (N_12683,N_12449,N_12474);
nor U12684 (N_12684,N_12592,N_12571);
and U12685 (N_12685,N_12596,N_12527);
nand U12686 (N_12686,N_12507,N_12433);
nor U12687 (N_12687,N_12598,N_12431);
nor U12688 (N_12688,N_12574,N_12521);
nor U12689 (N_12689,N_12583,N_12543);
nor U12690 (N_12690,N_12559,N_12450);
and U12691 (N_12691,N_12545,N_12597);
and U12692 (N_12692,N_12445,N_12509);
and U12693 (N_12693,N_12404,N_12562);
nand U12694 (N_12694,N_12548,N_12577);
or U12695 (N_12695,N_12572,N_12442);
nand U12696 (N_12696,N_12471,N_12563);
nor U12697 (N_12697,N_12470,N_12412);
and U12698 (N_12698,N_12546,N_12423);
nor U12699 (N_12699,N_12523,N_12437);
nor U12700 (N_12700,N_12401,N_12475);
or U12701 (N_12701,N_12530,N_12565);
nand U12702 (N_12702,N_12530,N_12592);
nor U12703 (N_12703,N_12450,N_12550);
or U12704 (N_12704,N_12580,N_12432);
and U12705 (N_12705,N_12562,N_12489);
nand U12706 (N_12706,N_12479,N_12474);
nor U12707 (N_12707,N_12407,N_12504);
nor U12708 (N_12708,N_12519,N_12436);
nor U12709 (N_12709,N_12529,N_12585);
nand U12710 (N_12710,N_12474,N_12462);
or U12711 (N_12711,N_12491,N_12423);
and U12712 (N_12712,N_12444,N_12539);
and U12713 (N_12713,N_12420,N_12597);
or U12714 (N_12714,N_12554,N_12436);
nand U12715 (N_12715,N_12550,N_12545);
and U12716 (N_12716,N_12416,N_12443);
or U12717 (N_12717,N_12466,N_12488);
nand U12718 (N_12718,N_12576,N_12590);
nand U12719 (N_12719,N_12508,N_12512);
nor U12720 (N_12720,N_12547,N_12473);
nand U12721 (N_12721,N_12475,N_12561);
or U12722 (N_12722,N_12426,N_12427);
or U12723 (N_12723,N_12534,N_12466);
and U12724 (N_12724,N_12461,N_12412);
nand U12725 (N_12725,N_12562,N_12409);
nor U12726 (N_12726,N_12527,N_12443);
or U12727 (N_12727,N_12593,N_12467);
nand U12728 (N_12728,N_12534,N_12415);
nand U12729 (N_12729,N_12486,N_12413);
or U12730 (N_12730,N_12407,N_12442);
nand U12731 (N_12731,N_12456,N_12415);
nand U12732 (N_12732,N_12487,N_12451);
or U12733 (N_12733,N_12429,N_12499);
and U12734 (N_12734,N_12526,N_12569);
nor U12735 (N_12735,N_12419,N_12482);
nand U12736 (N_12736,N_12544,N_12445);
nand U12737 (N_12737,N_12564,N_12431);
nor U12738 (N_12738,N_12538,N_12465);
or U12739 (N_12739,N_12547,N_12416);
nand U12740 (N_12740,N_12483,N_12590);
nor U12741 (N_12741,N_12444,N_12525);
and U12742 (N_12742,N_12538,N_12452);
or U12743 (N_12743,N_12517,N_12487);
and U12744 (N_12744,N_12550,N_12552);
nor U12745 (N_12745,N_12433,N_12469);
nand U12746 (N_12746,N_12464,N_12450);
and U12747 (N_12747,N_12594,N_12574);
xor U12748 (N_12748,N_12419,N_12428);
nor U12749 (N_12749,N_12430,N_12533);
or U12750 (N_12750,N_12449,N_12556);
or U12751 (N_12751,N_12465,N_12430);
nand U12752 (N_12752,N_12539,N_12505);
and U12753 (N_12753,N_12497,N_12410);
or U12754 (N_12754,N_12508,N_12523);
or U12755 (N_12755,N_12475,N_12541);
and U12756 (N_12756,N_12483,N_12563);
nand U12757 (N_12757,N_12557,N_12411);
and U12758 (N_12758,N_12433,N_12443);
nand U12759 (N_12759,N_12501,N_12531);
nor U12760 (N_12760,N_12494,N_12488);
nand U12761 (N_12761,N_12568,N_12584);
nor U12762 (N_12762,N_12403,N_12425);
or U12763 (N_12763,N_12569,N_12521);
nor U12764 (N_12764,N_12551,N_12477);
xnor U12765 (N_12765,N_12501,N_12478);
nor U12766 (N_12766,N_12565,N_12550);
nor U12767 (N_12767,N_12441,N_12478);
or U12768 (N_12768,N_12486,N_12561);
nand U12769 (N_12769,N_12539,N_12461);
nand U12770 (N_12770,N_12474,N_12549);
nor U12771 (N_12771,N_12496,N_12428);
or U12772 (N_12772,N_12580,N_12460);
nand U12773 (N_12773,N_12476,N_12539);
nor U12774 (N_12774,N_12476,N_12545);
nand U12775 (N_12775,N_12510,N_12437);
nor U12776 (N_12776,N_12430,N_12445);
nand U12777 (N_12777,N_12588,N_12497);
nand U12778 (N_12778,N_12440,N_12493);
nor U12779 (N_12779,N_12467,N_12407);
nor U12780 (N_12780,N_12517,N_12468);
and U12781 (N_12781,N_12564,N_12472);
and U12782 (N_12782,N_12419,N_12425);
and U12783 (N_12783,N_12590,N_12573);
and U12784 (N_12784,N_12475,N_12553);
nor U12785 (N_12785,N_12438,N_12473);
and U12786 (N_12786,N_12502,N_12476);
nand U12787 (N_12787,N_12411,N_12507);
and U12788 (N_12788,N_12402,N_12439);
nand U12789 (N_12789,N_12589,N_12550);
and U12790 (N_12790,N_12480,N_12496);
and U12791 (N_12791,N_12496,N_12429);
nand U12792 (N_12792,N_12561,N_12465);
nor U12793 (N_12793,N_12541,N_12486);
and U12794 (N_12794,N_12591,N_12444);
or U12795 (N_12795,N_12491,N_12439);
or U12796 (N_12796,N_12539,N_12546);
and U12797 (N_12797,N_12571,N_12436);
and U12798 (N_12798,N_12512,N_12423);
nand U12799 (N_12799,N_12503,N_12553);
and U12800 (N_12800,N_12715,N_12631);
nor U12801 (N_12801,N_12639,N_12664);
nor U12802 (N_12802,N_12628,N_12748);
nand U12803 (N_12803,N_12729,N_12653);
or U12804 (N_12804,N_12719,N_12629);
and U12805 (N_12805,N_12710,N_12633);
or U12806 (N_12806,N_12652,N_12750);
or U12807 (N_12807,N_12766,N_12742);
nand U12808 (N_12808,N_12637,N_12743);
and U12809 (N_12809,N_12609,N_12785);
nor U12810 (N_12810,N_12618,N_12615);
and U12811 (N_12811,N_12654,N_12709);
or U12812 (N_12812,N_12781,N_12706);
nor U12813 (N_12813,N_12784,N_12613);
nor U12814 (N_12814,N_12636,N_12663);
nor U12815 (N_12815,N_12707,N_12620);
nor U12816 (N_12816,N_12676,N_12641);
nand U12817 (N_12817,N_12705,N_12722);
or U12818 (N_12818,N_12662,N_12672);
nand U12819 (N_12819,N_12756,N_12773);
and U12820 (N_12820,N_12632,N_12690);
nor U12821 (N_12821,N_12683,N_12638);
nand U12822 (N_12822,N_12695,N_12603);
and U12823 (N_12823,N_12747,N_12621);
or U12824 (N_12824,N_12744,N_12627);
and U12825 (N_12825,N_12675,N_12704);
nand U12826 (N_12826,N_12778,N_12760);
nand U12827 (N_12827,N_12699,N_12795);
or U12828 (N_12828,N_12616,N_12716);
or U12829 (N_12829,N_12721,N_12777);
nor U12830 (N_12830,N_12780,N_12625);
or U12831 (N_12831,N_12712,N_12767);
and U12832 (N_12832,N_12720,N_12793);
or U12833 (N_12833,N_12749,N_12735);
and U12834 (N_12834,N_12634,N_12752);
or U12835 (N_12835,N_12684,N_12604);
nand U12836 (N_12836,N_12659,N_12799);
and U12837 (N_12837,N_12685,N_12666);
nand U12838 (N_12838,N_12758,N_12698);
nand U12839 (N_12839,N_12623,N_12728);
and U12840 (N_12840,N_12763,N_12682);
nand U12841 (N_12841,N_12601,N_12640);
nand U12842 (N_12842,N_12622,N_12726);
nand U12843 (N_12843,N_12725,N_12741);
or U12844 (N_12844,N_12770,N_12642);
and U12845 (N_12845,N_12635,N_12762);
or U12846 (N_12846,N_12746,N_12711);
and U12847 (N_12847,N_12772,N_12754);
nand U12848 (N_12848,N_12677,N_12670);
and U12849 (N_12849,N_12619,N_12786);
and U12850 (N_12850,N_12764,N_12790);
and U12851 (N_12851,N_12674,N_12791);
and U12852 (N_12852,N_12779,N_12740);
or U12853 (N_12853,N_12727,N_12724);
nand U12854 (N_12854,N_12671,N_12797);
nand U12855 (N_12855,N_12717,N_12649);
and U12856 (N_12856,N_12687,N_12776);
nor U12857 (N_12857,N_12650,N_12646);
nand U12858 (N_12858,N_12607,N_12755);
or U12859 (N_12859,N_12730,N_12678);
nand U12860 (N_12860,N_12765,N_12680);
nor U12861 (N_12861,N_12693,N_12644);
or U12862 (N_12862,N_12734,N_12768);
nand U12863 (N_12863,N_12691,N_12733);
nor U12864 (N_12864,N_12761,N_12718);
nor U12865 (N_12865,N_12771,N_12665);
and U12866 (N_12866,N_12608,N_12703);
and U12867 (N_12867,N_12751,N_12787);
nand U12868 (N_12868,N_12792,N_12739);
nand U12869 (N_12869,N_12679,N_12611);
xor U12870 (N_12870,N_12605,N_12602);
and U12871 (N_12871,N_12689,N_12713);
and U12872 (N_12872,N_12732,N_12775);
and U12873 (N_12873,N_12774,N_12697);
or U12874 (N_12874,N_12701,N_12789);
and U12875 (N_12875,N_12651,N_12658);
nor U12876 (N_12876,N_12759,N_12694);
and U12877 (N_12877,N_12630,N_12708);
or U12878 (N_12878,N_12796,N_12617);
or U12879 (N_12879,N_12714,N_12738);
and U12880 (N_12880,N_12668,N_12753);
or U12881 (N_12881,N_12626,N_12723);
or U12882 (N_12882,N_12661,N_12648);
or U12883 (N_12883,N_12757,N_12702);
nor U12884 (N_12884,N_12783,N_12645);
nor U12885 (N_12885,N_12731,N_12788);
or U12886 (N_12886,N_12686,N_12782);
nand U12887 (N_12887,N_12660,N_12737);
or U12888 (N_12888,N_12614,N_12798);
nor U12889 (N_12889,N_12643,N_12692);
or U12890 (N_12890,N_12656,N_12688);
xor U12891 (N_12891,N_12736,N_12794);
nand U12892 (N_12892,N_12681,N_12624);
nor U12893 (N_12893,N_12673,N_12696);
nor U12894 (N_12894,N_12600,N_12745);
or U12895 (N_12895,N_12647,N_12610);
nand U12896 (N_12896,N_12669,N_12700);
and U12897 (N_12897,N_12657,N_12667);
or U12898 (N_12898,N_12655,N_12606);
and U12899 (N_12899,N_12769,N_12612);
and U12900 (N_12900,N_12784,N_12704);
nor U12901 (N_12901,N_12659,N_12683);
and U12902 (N_12902,N_12627,N_12620);
nor U12903 (N_12903,N_12673,N_12601);
or U12904 (N_12904,N_12699,N_12602);
nand U12905 (N_12905,N_12789,N_12790);
nor U12906 (N_12906,N_12671,N_12632);
or U12907 (N_12907,N_12643,N_12794);
or U12908 (N_12908,N_12686,N_12689);
nor U12909 (N_12909,N_12643,N_12748);
nand U12910 (N_12910,N_12776,N_12679);
and U12911 (N_12911,N_12743,N_12776);
nor U12912 (N_12912,N_12785,N_12682);
and U12913 (N_12913,N_12629,N_12725);
or U12914 (N_12914,N_12604,N_12681);
and U12915 (N_12915,N_12692,N_12732);
nand U12916 (N_12916,N_12784,N_12743);
nand U12917 (N_12917,N_12751,N_12674);
nand U12918 (N_12918,N_12764,N_12717);
and U12919 (N_12919,N_12664,N_12634);
and U12920 (N_12920,N_12692,N_12756);
nand U12921 (N_12921,N_12615,N_12781);
and U12922 (N_12922,N_12732,N_12795);
or U12923 (N_12923,N_12749,N_12632);
or U12924 (N_12924,N_12605,N_12645);
nand U12925 (N_12925,N_12794,N_12701);
or U12926 (N_12926,N_12784,N_12789);
or U12927 (N_12927,N_12711,N_12778);
nor U12928 (N_12928,N_12654,N_12786);
or U12929 (N_12929,N_12679,N_12738);
or U12930 (N_12930,N_12789,N_12732);
nand U12931 (N_12931,N_12748,N_12739);
nand U12932 (N_12932,N_12710,N_12748);
nor U12933 (N_12933,N_12609,N_12760);
nand U12934 (N_12934,N_12715,N_12608);
and U12935 (N_12935,N_12725,N_12662);
nor U12936 (N_12936,N_12689,N_12799);
nor U12937 (N_12937,N_12696,N_12733);
nand U12938 (N_12938,N_12732,N_12618);
and U12939 (N_12939,N_12728,N_12643);
or U12940 (N_12940,N_12678,N_12705);
and U12941 (N_12941,N_12799,N_12705);
nor U12942 (N_12942,N_12720,N_12792);
or U12943 (N_12943,N_12635,N_12763);
and U12944 (N_12944,N_12765,N_12648);
and U12945 (N_12945,N_12787,N_12612);
and U12946 (N_12946,N_12620,N_12778);
nor U12947 (N_12947,N_12749,N_12705);
nor U12948 (N_12948,N_12655,N_12779);
and U12949 (N_12949,N_12618,N_12798);
nor U12950 (N_12950,N_12603,N_12707);
nand U12951 (N_12951,N_12799,N_12660);
or U12952 (N_12952,N_12756,N_12631);
nor U12953 (N_12953,N_12752,N_12764);
and U12954 (N_12954,N_12782,N_12662);
nor U12955 (N_12955,N_12639,N_12731);
xnor U12956 (N_12956,N_12727,N_12738);
and U12957 (N_12957,N_12633,N_12734);
or U12958 (N_12958,N_12782,N_12669);
nand U12959 (N_12959,N_12728,N_12672);
or U12960 (N_12960,N_12776,N_12606);
or U12961 (N_12961,N_12645,N_12693);
or U12962 (N_12962,N_12640,N_12712);
and U12963 (N_12963,N_12671,N_12775);
nand U12964 (N_12964,N_12788,N_12717);
or U12965 (N_12965,N_12657,N_12650);
nand U12966 (N_12966,N_12650,N_12615);
nand U12967 (N_12967,N_12691,N_12656);
or U12968 (N_12968,N_12630,N_12793);
or U12969 (N_12969,N_12608,N_12742);
nand U12970 (N_12970,N_12759,N_12761);
and U12971 (N_12971,N_12637,N_12629);
nand U12972 (N_12972,N_12745,N_12793);
nand U12973 (N_12973,N_12619,N_12640);
nor U12974 (N_12974,N_12761,N_12671);
or U12975 (N_12975,N_12645,N_12756);
nand U12976 (N_12976,N_12690,N_12739);
xor U12977 (N_12977,N_12685,N_12724);
or U12978 (N_12978,N_12685,N_12757);
and U12979 (N_12979,N_12741,N_12752);
and U12980 (N_12980,N_12748,N_12670);
xor U12981 (N_12981,N_12601,N_12739);
nor U12982 (N_12982,N_12658,N_12626);
nor U12983 (N_12983,N_12603,N_12727);
nand U12984 (N_12984,N_12740,N_12654);
nor U12985 (N_12985,N_12694,N_12772);
and U12986 (N_12986,N_12771,N_12690);
nand U12987 (N_12987,N_12708,N_12781);
or U12988 (N_12988,N_12642,N_12715);
nor U12989 (N_12989,N_12601,N_12773);
and U12990 (N_12990,N_12652,N_12791);
or U12991 (N_12991,N_12788,N_12626);
nor U12992 (N_12992,N_12783,N_12654);
nand U12993 (N_12993,N_12798,N_12743);
nor U12994 (N_12994,N_12773,N_12762);
nor U12995 (N_12995,N_12701,N_12670);
nand U12996 (N_12996,N_12708,N_12654);
and U12997 (N_12997,N_12720,N_12782);
nor U12998 (N_12998,N_12643,N_12732);
nand U12999 (N_12999,N_12748,N_12718);
nor U13000 (N_13000,N_12847,N_12923);
nor U13001 (N_13001,N_12959,N_12806);
nand U13002 (N_13002,N_12829,N_12906);
nor U13003 (N_13003,N_12948,N_12824);
or U13004 (N_13004,N_12823,N_12837);
and U13005 (N_13005,N_12812,N_12851);
and U13006 (N_13006,N_12865,N_12845);
or U13007 (N_13007,N_12828,N_12911);
nor U13008 (N_13008,N_12805,N_12898);
nand U13009 (N_13009,N_12884,N_12883);
nor U13010 (N_13010,N_12933,N_12920);
or U13011 (N_13011,N_12996,N_12950);
nand U13012 (N_13012,N_12893,N_12955);
nand U13013 (N_13013,N_12834,N_12924);
nand U13014 (N_13014,N_12966,N_12808);
and U13015 (N_13015,N_12861,N_12914);
or U13016 (N_13016,N_12863,N_12854);
nand U13017 (N_13017,N_12988,N_12989);
and U13018 (N_13018,N_12998,N_12822);
nor U13019 (N_13019,N_12975,N_12952);
or U13020 (N_13020,N_12846,N_12916);
or U13021 (N_13021,N_12905,N_12973);
nand U13022 (N_13022,N_12944,N_12903);
nand U13023 (N_13023,N_12977,N_12904);
or U13024 (N_13024,N_12810,N_12919);
nand U13025 (N_13025,N_12888,N_12960);
nor U13026 (N_13026,N_12964,N_12991);
nor U13027 (N_13027,N_12942,N_12860);
and U13028 (N_13028,N_12913,N_12871);
or U13029 (N_13029,N_12842,N_12885);
or U13030 (N_13030,N_12912,N_12984);
and U13031 (N_13031,N_12872,N_12907);
nand U13032 (N_13032,N_12895,N_12877);
nor U13033 (N_13033,N_12840,N_12831);
and U13034 (N_13034,N_12910,N_12813);
nand U13035 (N_13035,N_12821,N_12856);
nor U13036 (N_13036,N_12995,N_12880);
nor U13037 (N_13037,N_12848,N_12897);
and U13038 (N_13038,N_12982,N_12934);
and U13039 (N_13039,N_12953,N_12958);
nor U13040 (N_13040,N_12839,N_12804);
and U13041 (N_13041,N_12945,N_12825);
or U13042 (N_13042,N_12949,N_12838);
or U13043 (N_13043,N_12921,N_12870);
or U13044 (N_13044,N_12967,N_12807);
or U13045 (N_13045,N_12815,N_12890);
nand U13046 (N_13046,N_12935,N_12954);
nand U13047 (N_13047,N_12971,N_12855);
and U13048 (N_13048,N_12800,N_12850);
or U13049 (N_13049,N_12816,N_12994);
nand U13050 (N_13050,N_12896,N_12836);
nand U13051 (N_13051,N_12947,N_12867);
or U13052 (N_13052,N_12818,N_12915);
or U13053 (N_13053,N_12997,N_12957);
and U13054 (N_13054,N_12974,N_12802);
or U13055 (N_13055,N_12951,N_12817);
xnor U13056 (N_13056,N_12918,N_12835);
nor U13057 (N_13057,N_12961,N_12873);
and U13058 (N_13058,N_12830,N_12882);
and U13059 (N_13059,N_12956,N_12987);
nor U13060 (N_13060,N_12833,N_12841);
or U13061 (N_13061,N_12908,N_12811);
and U13062 (N_13062,N_12986,N_12827);
or U13063 (N_13063,N_12849,N_12875);
nand U13064 (N_13064,N_12843,N_12820);
and U13065 (N_13065,N_12927,N_12878);
nor U13066 (N_13066,N_12993,N_12852);
and U13067 (N_13067,N_12862,N_12853);
nand U13068 (N_13068,N_12932,N_12874);
and U13069 (N_13069,N_12801,N_12922);
or U13070 (N_13070,N_12925,N_12976);
nand U13071 (N_13071,N_12909,N_12930);
nor U13072 (N_13072,N_12809,N_12981);
nor U13073 (N_13073,N_12965,N_12999);
and U13074 (N_13074,N_12858,N_12937);
nand U13075 (N_13075,N_12868,N_12985);
and U13076 (N_13076,N_12946,N_12887);
nor U13077 (N_13077,N_12928,N_12826);
nand U13078 (N_13078,N_12859,N_12901);
and U13079 (N_13079,N_12926,N_12931);
or U13080 (N_13080,N_12938,N_12891);
nand U13081 (N_13081,N_12881,N_12992);
nor U13082 (N_13082,N_12894,N_12979);
nor U13083 (N_13083,N_12941,N_12943);
or U13084 (N_13084,N_12879,N_12814);
or U13085 (N_13085,N_12970,N_12917);
nor U13086 (N_13086,N_12864,N_12969);
nor U13087 (N_13087,N_12990,N_12844);
nor U13088 (N_13088,N_12899,N_12980);
nand U13089 (N_13089,N_12900,N_12832);
or U13090 (N_13090,N_12962,N_12963);
nor U13091 (N_13091,N_12876,N_12819);
or U13092 (N_13092,N_12978,N_12940);
nand U13093 (N_13093,N_12939,N_12902);
or U13094 (N_13094,N_12983,N_12869);
nor U13095 (N_13095,N_12936,N_12886);
or U13096 (N_13096,N_12889,N_12929);
nand U13097 (N_13097,N_12972,N_12892);
nor U13098 (N_13098,N_12803,N_12968);
nor U13099 (N_13099,N_12857,N_12866);
and U13100 (N_13100,N_12843,N_12823);
or U13101 (N_13101,N_12818,N_12806);
nand U13102 (N_13102,N_12830,N_12845);
nand U13103 (N_13103,N_12890,N_12802);
and U13104 (N_13104,N_12943,N_12993);
and U13105 (N_13105,N_12867,N_12880);
or U13106 (N_13106,N_12814,N_12829);
or U13107 (N_13107,N_12820,N_12985);
or U13108 (N_13108,N_12958,N_12842);
or U13109 (N_13109,N_12822,N_12852);
or U13110 (N_13110,N_12967,N_12873);
and U13111 (N_13111,N_12928,N_12946);
and U13112 (N_13112,N_12825,N_12800);
and U13113 (N_13113,N_12862,N_12919);
and U13114 (N_13114,N_12973,N_12868);
nor U13115 (N_13115,N_12904,N_12893);
and U13116 (N_13116,N_12857,N_12874);
or U13117 (N_13117,N_12983,N_12818);
nor U13118 (N_13118,N_12977,N_12851);
and U13119 (N_13119,N_12833,N_12893);
and U13120 (N_13120,N_12857,N_12802);
nand U13121 (N_13121,N_12945,N_12929);
or U13122 (N_13122,N_12946,N_12858);
nor U13123 (N_13123,N_12912,N_12977);
nor U13124 (N_13124,N_12896,N_12863);
nand U13125 (N_13125,N_12828,N_12818);
and U13126 (N_13126,N_12912,N_12924);
or U13127 (N_13127,N_12800,N_12847);
nor U13128 (N_13128,N_12911,N_12850);
nand U13129 (N_13129,N_12921,N_12895);
nand U13130 (N_13130,N_12809,N_12891);
or U13131 (N_13131,N_12820,N_12805);
and U13132 (N_13132,N_12895,N_12998);
nand U13133 (N_13133,N_12824,N_12860);
or U13134 (N_13134,N_12867,N_12932);
and U13135 (N_13135,N_12860,N_12864);
nand U13136 (N_13136,N_12932,N_12978);
or U13137 (N_13137,N_12839,N_12897);
nand U13138 (N_13138,N_12821,N_12975);
or U13139 (N_13139,N_12937,N_12815);
or U13140 (N_13140,N_12835,N_12872);
and U13141 (N_13141,N_12858,N_12967);
and U13142 (N_13142,N_12948,N_12811);
nand U13143 (N_13143,N_12831,N_12945);
nand U13144 (N_13144,N_12867,N_12843);
nor U13145 (N_13145,N_12825,N_12849);
or U13146 (N_13146,N_12960,N_12821);
and U13147 (N_13147,N_12817,N_12999);
or U13148 (N_13148,N_12901,N_12978);
nand U13149 (N_13149,N_12914,N_12957);
and U13150 (N_13150,N_12822,N_12951);
or U13151 (N_13151,N_12937,N_12910);
nand U13152 (N_13152,N_12982,N_12869);
nor U13153 (N_13153,N_12985,N_12993);
nand U13154 (N_13154,N_12881,N_12832);
and U13155 (N_13155,N_12909,N_12855);
nand U13156 (N_13156,N_12963,N_12947);
nor U13157 (N_13157,N_12977,N_12948);
nor U13158 (N_13158,N_12848,N_12821);
or U13159 (N_13159,N_12968,N_12960);
and U13160 (N_13160,N_12863,N_12982);
or U13161 (N_13161,N_12989,N_12950);
nand U13162 (N_13162,N_12816,N_12949);
nor U13163 (N_13163,N_12900,N_12989);
and U13164 (N_13164,N_12810,N_12824);
nor U13165 (N_13165,N_12941,N_12992);
and U13166 (N_13166,N_12822,N_12973);
and U13167 (N_13167,N_12851,N_12956);
or U13168 (N_13168,N_12891,N_12864);
and U13169 (N_13169,N_12857,N_12988);
nand U13170 (N_13170,N_12893,N_12831);
or U13171 (N_13171,N_12973,N_12976);
nand U13172 (N_13172,N_12993,N_12919);
nor U13173 (N_13173,N_12938,N_12989);
and U13174 (N_13174,N_12997,N_12801);
or U13175 (N_13175,N_12984,N_12836);
xnor U13176 (N_13176,N_12968,N_12959);
or U13177 (N_13177,N_12930,N_12857);
and U13178 (N_13178,N_12812,N_12808);
and U13179 (N_13179,N_12853,N_12918);
and U13180 (N_13180,N_12958,N_12817);
nor U13181 (N_13181,N_12805,N_12808);
nand U13182 (N_13182,N_12809,N_12818);
nand U13183 (N_13183,N_12969,N_12960);
nor U13184 (N_13184,N_12838,N_12861);
xor U13185 (N_13185,N_12909,N_12858);
nand U13186 (N_13186,N_12816,N_12953);
and U13187 (N_13187,N_12830,N_12801);
or U13188 (N_13188,N_12853,N_12994);
nor U13189 (N_13189,N_12830,N_12967);
or U13190 (N_13190,N_12814,N_12880);
nand U13191 (N_13191,N_12905,N_12883);
nand U13192 (N_13192,N_12838,N_12865);
nor U13193 (N_13193,N_12921,N_12978);
and U13194 (N_13194,N_12829,N_12821);
and U13195 (N_13195,N_12803,N_12912);
nor U13196 (N_13196,N_12968,N_12947);
or U13197 (N_13197,N_12894,N_12870);
or U13198 (N_13198,N_12841,N_12812);
nor U13199 (N_13199,N_12819,N_12971);
nand U13200 (N_13200,N_13089,N_13160);
and U13201 (N_13201,N_13028,N_13162);
nand U13202 (N_13202,N_13106,N_13052);
and U13203 (N_13203,N_13087,N_13114);
nor U13204 (N_13204,N_13058,N_13053);
nand U13205 (N_13205,N_13167,N_13144);
and U13206 (N_13206,N_13066,N_13072);
or U13207 (N_13207,N_13140,N_13004);
nor U13208 (N_13208,N_13172,N_13020);
xor U13209 (N_13209,N_13179,N_13154);
or U13210 (N_13210,N_13043,N_13169);
or U13211 (N_13211,N_13184,N_13037);
nor U13212 (N_13212,N_13161,N_13159);
and U13213 (N_13213,N_13009,N_13067);
nor U13214 (N_13214,N_13045,N_13117);
or U13215 (N_13215,N_13060,N_13068);
nor U13216 (N_13216,N_13126,N_13012);
nor U13217 (N_13217,N_13092,N_13038);
and U13218 (N_13218,N_13123,N_13081);
and U13219 (N_13219,N_13007,N_13166);
nand U13220 (N_13220,N_13024,N_13063);
or U13221 (N_13221,N_13136,N_13109);
nor U13222 (N_13222,N_13014,N_13198);
and U13223 (N_13223,N_13189,N_13168);
nand U13224 (N_13224,N_13036,N_13199);
and U13225 (N_13225,N_13061,N_13049);
and U13226 (N_13226,N_13195,N_13175);
nand U13227 (N_13227,N_13143,N_13134);
nor U13228 (N_13228,N_13054,N_13059);
and U13229 (N_13229,N_13133,N_13181);
and U13230 (N_13230,N_13086,N_13002);
and U13231 (N_13231,N_13155,N_13101);
nand U13232 (N_13232,N_13026,N_13138);
and U13233 (N_13233,N_13030,N_13149);
and U13234 (N_13234,N_13048,N_13041);
nand U13235 (N_13235,N_13115,N_13118);
and U13236 (N_13236,N_13022,N_13191);
or U13237 (N_13237,N_13122,N_13142);
and U13238 (N_13238,N_13112,N_13147);
nand U13239 (N_13239,N_13103,N_13111);
and U13240 (N_13240,N_13046,N_13124);
and U13241 (N_13241,N_13055,N_13033);
and U13242 (N_13242,N_13165,N_13015);
nand U13243 (N_13243,N_13156,N_13008);
nand U13244 (N_13244,N_13098,N_13097);
and U13245 (N_13245,N_13108,N_13150);
nand U13246 (N_13246,N_13047,N_13141);
nor U13247 (N_13247,N_13176,N_13104);
and U13248 (N_13248,N_13158,N_13027);
or U13249 (N_13249,N_13069,N_13001);
and U13250 (N_13250,N_13183,N_13197);
and U13251 (N_13251,N_13185,N_13051);
and U13252 (N_13252,N_13035,N_13075);
or U13253 (N_13253,N_13146,N_13164);
or U13254 (N_13254,N_13129,N_13107);
and U13255 (N_13255,N_13153,N_13171);
nand U13256 (N_13256,N_13186,N_13005);
nor U13257 (N_13257,N_13082,N_13096);
nand U13258 (N_13258,N_13102,N_13021);
and U13259 (N_13259,N_13019,N_13040);
or U13260 (N_13260,N_13003,N_13148);
and U13261 (N_13261,N_13032,N_13152);
xnor U13262 (N_13262,N_13110,N_13079);
and U13263 (N_13263,N_13132,N_13119);
nand U13264 (N_13264,N_13174,N_13090);
nor U13265 (N_13265,N_13177,N_13151);
nor U13266 (N_13266,N_13016,N_13180);
or U13267 (N_13267,N_13018,N_13145);
and U13268 (N_13268,N_13044,N_13139);
nor U13269 (N_13269,N_13095,N_13091);
and U13270 (N_13270,N_13157,N_13116);
and U13271 (N_13271,N_13029,N_13057);
nand U13272 (N_13272,N_13083,N_13031);
nand U13273 (N_13273,N_13128,N_13064);
nand U13274 (N_13274,N_13125,N_13135);
and U13275 (N_13275,N_13088,N_13042);
nand U13276 (N_13276,N_13130,N_13100);
nor U13277 (N_13277,N_13073,N_13011);
nand U13278 (N_13278,N_13131,N_13071);
nand U13279 (N_13279,N_13077,N_13034);
and U13280 (N_13280,N_13078,N_13094);
or U13281 (N_13281,N_13076,N_13192);
nor U13282 (N_13282,N_13173,N_13013);
nor U13283 (N_13283,N_13039,N_13050);
nor U13284 (N_13284,N_13178,N_13010);
and U13285 (N_13285,N_13000,N_13187);
and U13286 (N_13286,N_13194,N_13017);
and U13287 (N_13287,N_13062,N_13190);
and U13288 (N_13288,N_13137,N_13074);
and U13289 (N_13289,N_13105,N_13080);
nand U13290 (N_13290,N_13093,N_13188);
and U13291 (N_13291,N_13193,N_13085);
nor U13292 (N_13292,N_13065,N_13121);
nor U13293 (N_13293,N_13025,N_13084);
or U13294 (N_13294,N_13170,N_13196);
or U13295 (N_13295,N_13182,N_13070);
nor U13296 (N_13296,N_13006,N_13127);
nor U13297 (N_13297,N_13023,N_13099);
nor U13298 (N_13298,N_13163,N_13056);
nor U13299 (N_13299,N_13113,N_13120);
nand U13300 (N_13300,N_13046,N_13145);
and U13301 (N_13301,N_13150,N_13107);
or U13302 (N_13302,N_13086,N_13115);
nand U13303 (N_13303,N_13180,N_13148);
or U13304 (N_13304,N_13124,N_13179);
and U13305 (N_13305,N_13193,N_13119);
nor U13306 (N_13306,N_13089,N_13122);
and U13307 (N_13307,N_13019,N_13178);
or U13308 (N_13308,N_13002,N_13158);
and U13309 (N_13309,N_13008,N_13021);
nor U13310 (N_13310,N_13112,N_13135);
or U13311 (N_13311,N_13067,N_13033);
and U13312 (N_13312,N_13143,N_13152);
nand U13313 (N_13313,N_13114,N_13172);
or U13314 (N_13314,N_13141,N_13088);
and U13315 (N_13315,N_13067,N_13087);
or U13316 (N_13316,N_13028,N_13154);
and U13317 (N_13317,N_13030,N_13114);
nor U13318 (N_13318,N_13001,N_13088);
nand U13319 (N_13319,N_13157,N_13152);
and U13320 (N_13320,N_13196,N_13080);
and U13321 (N_13321,N_13199,N_13183);
or U13322 (N_13322,N_13183,N_13113);
and U13323 (N_13323,N_13105,N_13050);
and U13324 (N_13324,N_13008,N_13118);
or U13325 (N_13325,N_13071,N_13079);
nor U13326 (N_13326,N_13197,N_13172);
nor U13327 (N_13327,N_13154,N_13068);
nand U13328 (N_13328,N_13083,N_13060);
nand U13329 (N_13329,N_13102,N_13033);
and U13330 (N_13330,N_13066,N_13113);
and U13331 (N_13331,N_13033,N_13084);
and U13332 (N_13332,N_13196,N_13188);
and U13333 (N_13333,N_13095,N_13004);
nand U13334 (N_13334,N_13038,N_13017);
nor U13335 (N_13335,N_13036,N_13040);
or U13336 (N_13336,N_13090,N_13035);
nor U13337 (N_13337,N_13112,N_13155);
or U13338 (N_13338,N_13102,N_13028);
nor U13339 (N_13339,N_13127,N_13165);
or U13340 (N_13340,N_13014,N_13160);
and U13341 (N_13341,N_13158,N_13192);
nand U13342 (N_13342,N_13106,N_13064);
nand U13343 (N_13343,N_13071,N_13041);
nand U13344 (N_13344,N_13153,N_13111);
nand U13345 (N_13345,N_13016,N_13036);
or U13346 (N_13346,N_13003,N_13105);
nor U13347 (N_13347,N_13082,N_13047);
nand U13348 (N_13348,N_13106,N_13166);
and U13349 (N_13349,N_13181,N_13170);
or U13350 (N_13350,N_13169,N_13110);
nand U13351 (N_13351,N_13050,N_13177);
or U13352 (N_13352,N_13032,N_13105);
or U13353 (N_13353,N_13110,N_13193);
and U13354 (N_13354,N_13192,N_13199);
or U13355 (N_13355,N_13031,N_13113);
or U13356 (N_13356,N_13055,N_13133);
and U13357 (N_13357,N_13145,N_13048);
and U13358 (N_13358,N_13138,N_13044);
and U13359 (N_13359,N_13127,N_13195);
and U13360 (N_13360,N_13129,N_13029);
or U13361 (N_13361,N_13031,N_13046);
or U13362 (N_13362,N_13022,N_13107);
nand U13363 (N_13363,N_13041,N_13153);
nor U13364 (N_13364,N_13162,N_13137);
and U13365 (N_13365,N_13188,N_13053);
or U13366 (N_13366,N_13184,N_13070);
or U13367 (N_13367,N_13046,N_13152);
or U13368 (N_13368,N_13147,N_13091);
nand U13369 (N_13369,N_13104,N_13159);
nor U13370 (N_13370,N_13001,N_13045);
and U13371 (N_13371,N_13039,N_13101);
nand U13372 (N_13372,N_13044,N_13042);
nand U13373 (N_13373,N_13105,N_13044);
nor U13374 (N_13374,N_13160,N_13169);
nand U13375 (N_13375,N_13004,N_13049);
nor U13376 (N_13376,N_13080,N_13054);
nand U13377 (N_13377,N_13196,N_13136);
and U13378 (N_13378,N_13114,N_13097);
nor U13379 (N_13379,N_13094,N_13130);
and U13380 (N_13380,N_13076,N_13005);
or U13381 (N_13381,N_13164,N_13103);
or U13382 (N_13382,N_13057,N_13071);
nand U13383 (N_13383,N_13115,N_13193);
nand U13384 (N_13384,N_13108,N_13021);
nor U13385 (N_13385,N_13037,N_13190);
nand U13386 (N_13386,N_13040,N_13123);
or U13387 (N_13387,N_13199,N_13179);
nand U13388 (N_13388,N_13131,N_13104);
or U13389 (N_13389,N_13085,N_13013);
or U13390 (N_13390,N_13073,N_13193);
or U13391 (N_13391,N_13179,N_13101);
or U13392 (N_13392,N_13177,N_13124);
and U13393 (N_13393,N_13194,N_13048);
and U13394 (N_13394,N_13025,N_13122);
and U13395 (N_13395,N_13089,N_13172);
nor U13396 (N_13396,N_13003,N_13029);
and U13397 (N_13397,N_13092,N_13108);
xor U13398 (N_13398,N_13100,N_13037);
nor U13399 (N_13399,N_13092,N_13179);
nor U13400 (N_13400,N_13223,N_13230);
nand U13401 (N_13401,N_13288,N_13359);
nor U13402 (N_13402,N_13395,N_13201);
nand U13403 (N_13403,N_13337,N_13398);
or U13404 (N_13404,N_13274,N_13377);
or U13405 (N_13405,N_13277,N_13236);
or U13406 (N_13406,N_13380,N_13289);
nor U13407 (N_13407,N_13271,N_13280);
or U13408 (N_13408,N_13373,N_13365);
and U13409 (N_13409,N_13383,N_13374);
or U13410 (N_13410,N_13316,N_13234);
or U13411 (N_13411,N_13360,N_13338);
and U13412 (N_13412,N_13286,N_13253);
or U13413 (N_13413,N_13282,N_13336);
nand U13414 (N_13414,N_13366,N_13251);
nor U13415 (N_13415,N_13264,N_13296);
nor U13416 (N_13416,N_13300,N_13312);
and U13417 (N_13417,N_13320,N_13200);
nand U13418 (N_13418,N_13206,N_13212);
and U13419 (N_13419,N_13367,N_13248);
nand U13420 (N_13420,N_13325,N_13335);
nand U13421 (N_13421,N_13311,N_13244);
and U13422 (N_13422,N_13202,N_13252);
and U13423 (N_13423,N_13396,N_13235);
or U13424 (N_13424,N_13260,N_13246);
nand U13425 (N_13425,N_13275,N_13265);
nor U13426 (N_13426,N_13256,N_13306);
and U13427 (N_13427,N_13267,N_13295);
or U13428 (N_13428,N_13392,N_13220);
nand U13429 (N_13429,N_13301,N_13371);
nor U13430 (N_13430,N_13231,N_13391);
or U13431 (N_13431,N_13238,N_13389);
nor U13432 (N_13432,N_13349,N_13217);
nor U13433 (N_13433,N_13326,N_13321);
nor U13434 (N_13434,N_13283,N_13393);
nor U13435 (N_13435,N_13250,N_13378);
or U13436 (N_13436,N_13268,N_13272);
and U13437 (N_13437,N_13315,N_13384);
nor U13438 (N_13438,N_13281,N_13352);
or U13439 (N_13439,N_13386,N_13278);
nor U13440 (N_13440,N_13329,N_13328);
nand U13441 (N_13441,N_13364,N_13203);
nand U13442 (N_13442,N_13259,N_13368);
nand U13443 (N_13443,N_13342,N_13273);
nor U13444 (N_13444,N_13237,N_13339);
and U13445 (N_13445,N_13333,N_13222);
or U13446 (N_13446,N_13348,N_13345);
nor U13447 (N_13447,N_13347,N_13387);
and U13448 (N_13448,N_13362,N_13255);
and U13449 (N_13449,N_13361,N_13287);
and U13450 (N_13450,N_13350,N_13204);
or U13451 (N_13451,N_13247,N_13375);
nor U13452 (N_13452,N_13385,N_13245);
or U13453 (N_13453,N_13307,N_13284);
nor U13454 (N_13454,N_13304,N_13322);
xnor U13455 (N_13455,N_13221,N_13317);
nand U13456 (N_13456,N_13310,N_13213);
nor U13457 (N_13457,N_13292,N_13327);
or U13458 (N_13458,N_13279,N_13209);
and U13459 (N_13459,N_13344,N_13334);
or U13460 (N_13460,N_13254,N_13372);
nand U13461 (N_13461,N_13269,N_13258);
nand U13462 (N_13462,N_13382,N_13227);
nand U13463 (N_13463,N_13257,N_13318);
nor U13464 (N_13464,N_13397,N_13241);
nor U13465 (N_13465,N_13302,N_13218);
or U13466 (N_13466,N_13353,N_13331);
or U13467 (N_13467,N_13276,N_13232);
nand U13468 (N_13468,N_13207,N_13226);
or U13469 (N_13469,N_13369,N_13305);
nor U13470 (N_13470,N_13219,N_13358);
nand U13471 (N_13471,N_13210,N_13239);
or U13472 (N_13472,N_13355,N_13376);
or U13473 (N_13473,N_13215,N_13399);
nand U13474 (N_13474,N_13211,N_13249);
or U13475 (N_13475,N_13381,N_13356);
or U13476 (N_13476,N_13308,N_13290);
xnor U13477 (N_13477,N_13351,N_13388);
and U13478 (N_13478,N_13270,N_13224);
or U13479 (N_13479,N_13216,N_13319);
nor U13480 (N_13480,N_13243,N_13262);
nand U13481 (N_13481,N_13214,N_13297);
and U13482 (N_13482,N_13285,N_13309);
or U13483 (N_13483,N_13314,N_13291);
and U13484 (N_13484,N_13363,N_13225);
or U13485 (N_13485,N_13330,N_13390);
or U13486 (N_13486,N_13298,N_13263);
or U13487 (N_13487,N_13242,N_13343);
or U13488 (N_13488,N_13240,N_13205);
nor U13489 (N_13489,N_13294,N_13324);
nand U13490 (N_13490,N_13370,N_13229);
nand U13491 (N_13491,N_13233,N_13293);
nand U13492 (N_13492,N_13228,N_13357);
and U13493 (N_13493,N_13266,N_13394);
or U13494 (N_13494,N_13354,N_13332);
nor U13495 (N_13495,N_13208,N_13303);
nand U13496 (N_13496,N_13340,N_13323);
and U13497 (N_13497,N_13346,N_13341);
nand U13498 (N_13498,N_13299,N_13313);
nor U13499 (N_13499,N_13379,N_13261);
and U13500 (N_13500,N_13276,N_13249);
or U13501 (N_13501,N_13308,N_13315);
xnor U13502 (N_13502,N_13370,N_13331);
nand U13503 (N_13503,N_13209,N_13349);
nand U13504 (N_13504,N_13232,N_13399);
or U13505 (N_13505,N_13384,N_13259);
and U13506 (N_13506,N_13330,N_13209);
or U13507 (N_13507,N_13360,N_13271);
nor U13508 (N_13508,N_13250,N_13349);
nor U13509 (N_13509,N_13334,N_13373);
nand U13510 (N_13510,N_13369,N_13212);
nand U13511 (N_13511,N_13341,N_13391);
or U13512 (N_13512,N_13357,N_13381);
or U13513 (N_13513,N_13386,N_13351);
or U13514 (N_13514,N_13375,N_13394);
nor U13515 (N_13515,N_13220,N_13293);
nor U13516 (N_13516,N_13381,N_13321);
and U13517 (N_13517,N_13397,N_13289);
or U13518 (N_13518,N_13238,N_13247);
nor U13519 (N_13519,N_13334,N_13350);
or U13520 (N_13520,N_13331,N_13340);
or U13521 (N_13521,N_13325,N_13376);
nor U13522 (N_13522,N_13224,N_13206);
and U13523 (N_13523,N_13252,N_13379);
nand U13524 (N_13524,N_13228,N_13389);
or U13525 (N_13525,N_13229,N_13322);
or U13526 (N_13526,N_13297,N_13386);
nand U13527 (N_13527,N_13240,N_13380);
nand U13528 (N_13528,N_13368,N_13261);
nand U13529 (N_13529,N_13355,N_13305);
nand U13530 (N_13530,N_13314,N_13324);
and U13531 (N_13531,N_13352,N_13286);
nor U13532 (N_13532,N_13201,N_13371);
or U13533 (N_13533,N_13230,N_13265);
and U13534 (N_13534,N_13389,N_13246);
and U13535 (N_13535,N_13241,N_13260);
nand U13536 (N_13536,N_13384,N_13271);
and U13537 (N_13537,N_13395,N_13322);
and U13538 (N_13538,N_13285,N_13308);
nor U13539 (N_13539,N_13324,N_13381);
or U13540 (N_13540,N_13307,N_13231);
or U13541 (N_13541,N_13225,N_13261);
or U13542 (N_13542,N_13221,N_13283);
or U13543 (N_13543,N_13271,N_13214);
and U13544 (N_13544,N_13276,N_13223);
nor U13545 (N_13545,N_13239,N_13308);
nor U13546 (N_13546,N_13226,N_13256);
and U13547 (N_13547,N_13228,N_13372);
nor U13548 (N_13548,N_13321,N_13266);
nor U13549 (N_13549,N_13281,N_13258);
and U13550 (N_13550,N_13261,N_13382);
nand U13551 (N_13551,N_13286,N_13322);
nor U13552 (N_13552,N_13312,N_13296);
nand U13553 (N_13553,N_13369,N_13337);
or U13554 (N_13554,N_13340,N_13319);
nor U13555 (N_13555,N_13309,N_13333);
xnor U13556 (N_13556,N_13300,N_13293);
and U13557 (N_13557,N_13295,N_13375);
nor U13558 (N_13558,N_13294,N_13239);
nand U13559 (N_13559,N_13262,N_13269);
or U13560 (N_13560,N_13338,N_13223);
and U13561 (N_13561,N_13319,N_13377);
or U13562 (N_13562,N_13232,N_13384);
or U13563 (N_13563,N_13208,N_13202);
nand U13564 (N_13564,N_13267,N_13299);
nor U13565 (N_13565,N_13302,N_13216);
nor U13566 (N_13566,N_13279,N_13262);
nor U13567 (N_13567,N_13214,N_13230);
nand U13568 (N_13568,N_13346,N_13373);
nand U13569 (N_13569,N_13264,N_13278);
nor U13570 (N_13570,N_13292,N_13299);
and U13571 (N_13571,N_13248,N_13399);
or U13572 (N_13572,N_13280,N_13287);
or U13573 (N_13573,N_13234,N_13214);
nand U13574 (N_13574,N_13358,N_13261);
and U13575 (N_13575,N_13378,N_13266);
or U13576 (N_13576,N_13333,N_13210);
nand U13577 (N_13577,N_13335,N_13366);
and U13578 (N_13578,N_13201,N_13267);
nor U13579 (N_13579,N_13240,N_13319);
and U13580 (N_13580,N_13286,N_13271);
nand U13581 (N_13581,N_13341,N_13274);
nand U13582 (N_13582,N_13311,N_13245);
nand U13583 (N_13583,N_13268,N_13265);
nor U13584 (N_13584,N_13209,N_13379);
and U13585 (N_13585,N_13266,N_13332);
nand U13586 (N_13586,N_13351,N_13238);
and U13587 (N_13587,N_13238,N_13350);
or U13588 (N_13588,N_13384,N_13333);
nor U13589 (N_13589,N_13266,N_13265);
and U13590 (N_13590,N_13256,N_13393);
nand U13591 (N_13591,N_13359,N_13221);
nor U13592 (N_13592,N_13221,N_13294);
nor U13593 (N_13593,N_13329,N_13220);
nor U13594 (N_13594,N_13209,N_13320);
or U13595 (N_13595,N_13328,N_13391);
nand U13596 (N_13596,N_13200,N_13221);
nand U13597 (N_13597,N_13338,N_13384);
and U13598 (N_13598,N_13275,N_13232);
or U13599 (N_13599,N_13282,N_13276);
nor U13600 (N_13600,N_13591,N_13414);
nand U13601 (N_13601,N_13447,N_13473);
nand U13602 (N_13602,N_13418,N_13485);
or U13603 (N_13603,N_13562,N_13403);
and U13604 (N_13604,N_13507,N_13512);
nand U13605 (N_13605,N_13555,N_13574);
and U13606 (N_13606,N_13504,N_13544);
or U13607 (N_13607,N_13419,N_13529);
and U13608 (N_13608,N_13505,N_13405);
xnor U13609 (N_13609,N_13582,N_13462);
nand U13610 (N_13610,N_13542,N_13596);
nor U13611 (N_13611,N_13571,N_13422);
and U13612 (N_13612,N_13444,N_13416);
nor U13613 (N_13613,N_13569,N_13423);
nor U13614 (N_13614,N_13537,N_13427);
or U13615 (N_13615,N_13404,N_13451);
and U13616 (N_13616,N_13411,N_13494);
and U13617 (N_13617,N_13522,N_13471);
nor U13618 (N_13618,N_13568,N_13420);
or U13619 (N_13619,N_13453,N_13580);
or U13620 (N_13620,N_13521,N_13465);
nor U13621 (N_13621,N_13502,N_13468);
and U13622 (N_13622,N_13531,N_13430);
nand U13623 (N_13623,N_13593,N_13527);
and U13624 (N_13624,N_13501,N_13449);
and U13625 (N_13625,N_13472,N_13470);
nand U13626 (N_13626,N_13532,N_13567);
or U13627 (N_13627,N_13459,N_13481);
and U13628 (N_13628,N_13415,N_13460);
and U13629 (N_13629,N_13429,N_13439);
nand U13630 (N_13630,N_13484,N_13587);
nand U13631 (N_13631,N_13466,N_13588);
or U13632 (N_13632,N_13592,N_13454);
and U13633 (N_13633,N_13495,N_13421);
and U13634 (N_13634,N_13450,N_13553);
nor U13635 (N_13635,N_13528,N_13402);
or U13636 (N_13636,N_13536,N_13488);
xnor U13637 (N_13637,N_13464,N_13575);
or U13638 (N_13638,N_13576,N_13540);
nand U13639 (N_13639,N_13518,N_13487);
or U13640 (N_13640,N_13517,N_13424);
nand U13641 (N_13641,N_13434,N_13483);
or U13642 (N_13642,N_13526,N_13486);
or U13643 (N_13643,N_13581,N_13566);
nor U13644 (N_13644,N_13557,N_13438);
and U13645 (N_13645,N_13598,N_13432);
or U13646 (N_13646,N_13476,N_13583);
nor U13647 (N_13647,N_13463,N_13428);
nand U13648 (N_13648,N_13508,N_13547);
and U13649 (N_13649,N_13577,N_13590);
or U13650 (N_13650,N_13477,N_13546);
nor U13651 (N_13651,N_13552,N_13509);
nand U13652 (N_13652,N_13426,N_13445);
nor U13653 (N_13653,N_13497,N_13589);
nor U13654 (N_13654,N_13493,N_13452);
and U13655 (N_13655,N_13417,N_13413);
and U13656 (N_13656,N_13530,N_13407);
or U13657 (N_13657,N_13584,N_13533);
or U13658 (N_13658,N_13482,N_13519);
or U13659 (N_13659,N_13457,N_13412);
and U13660 (N_13660,N_13561,N_13491);
nand U13661 (N_13661,N_13446,N_13543);
and U13662 (N_13662,N_13585,N_13539);
and U13663 (N_13663,N_13594,N_13578);
or U13664 (N_13664,N_13554,N_13523);
nand U13665 (N_13665,N_13513,N_13437);
or U13666 (N_13666,N_13538,N_13516);
or U13667 (N_13667,N_13560,N_13549);
and U13668 (N_13668,N_13525,N_13489);
nand U13669 (N_13669,N_13490,N_13406);
or U13670 (N_13670,N_13541,N_13436);
and U13671 (N_13671,N_13524,N_13558);
nand U13672 (N_13672,N_13448,N_13548);
or U13673 (N_13673,N_13579,N_13599);
and U13674 (N_13674,N_13559,N_13425);
xor U13675 (N_13675,N_13442,N_13455);
or U13676 (N_13676,N_13431,N_13469);
or U13677 (N_13677,N_13565,N_13534);
and U13678 (N_13678,N_13556,N_13492);
or U13679 (N_13679,N_13570,N_13433);
nor U13680 (N_13680,N_13503,N_13551);
or U13681 (N_13681,N_13456,N_13410);
or U13682 (N_13682,N_13564,N_13475);
nand U13683 (N_13683,N_13572,N_13458);
nand U13684 (N_13684,N_13496,N_13510);
xnor U13685 (N_13685,N_13573,N_13499);
nand U13686 (N_13686,N_13435,N_13443);
nand U13687 (N_13687,N_13595,N_13535);
xor U13688 (N_13688,N_13515,N_13511);
or U13689 (N_13689,N_13440,N_13586);
and U13690 (N_13690,N_13478,N_13409);
and U13691 (N_13691,N_13506,N_13498);
or U13692 (N_13692,N_13474,N_13480);
or U13693 (N_13693,N_13479,N_13461);
or U13694 (N_13694,N_13597,N_13401);
nand U13695 (N_13695,N_13500,N_13545);
nand U13696 (N_13696,N_13441,N_13408);
or U13697 (N_13697,N_13400,N_13467);
nand U13698 (N_13698,N_13520,N_13563);
or U13699 (N_13699,N_13514,N_13550);
or U13700 (N_13700,N_13508,N_13544);
nand U13701 (N_13701,N_13506,N_13404);
nor U13702 (N_13702,N_13560,N_13599);
and U13703 (N_13703,N_13430,N_13406);
and U13704 (N_13704,N_13571,N_13523);
and U13705 (N_13705,N_13584,N_13495);
and U13706 (N_13706,N_13529,N_13567);
and U13707 (N_13707,N_13439,N_13462);
and U13708 (N_13708,N_13406,N_13526);
xor U13709 (N_13709,N_13586,N_13405);
xnor U13710 (N_13710,N_13408,N_13492);
nand U13711 (N_13711,N_13432,N_13483);
and U13712 (N_13712,N_13466,N_13569);
nor U13713 (N_13713,N_13511,N_13505);
or U13714 (N_13714,N_13445,N_13554);
or U13715 (N_13715,N_13574,N_13538);
or U13716 (N_13716,N_13579,N_13487);
or U13717 (N_13717,N_13539,N_13514);
nand U13718 (N_13718,N_13538,N_13570);
nor U13719 (N_13719,N_13504,N_13414);
and U13720 (N_13720,N_13551,N_13533);
nand U13721 (N_13721,N_13582,N_13445);
nand U13722 (N_13722,N_13549,N_13491);
nor U13723 (N_13723,N_13411,N_13563);
and U13724 (N_13724,N_13519,N_13566);
and U13725 (N_13725,N_13467,N_13487);
nor U13726 (N_13726,N_13408,N_13514);
nand U13727 (N_13727,N_13494,N_13452);
and U13728 (N_13728,N_13456,N_13499);
or U13729 (N_13729,N_13429,N_13568);
nor U13730 (N_13730,N_13591,N_13401);
xnor U13731 (N_13731,N_13507,N_13537);
nand U13732 (N_13732,N_13533,N_13436);
nand U13733 (N_13733,N_13550,N_13582);
xor U13734 (N_13734,N_13525,N_13450);
nor U13735 (N_13735,N_13533,N_13401);
nand U13736 (N_13736,N_13599,N_13474);
and U13737 (N_13737,N_13497,N_13449);
and U13738 (N_13738,N_13513,N_13575);
nor U13739 (N_13739,N_13507,N_13495);
nor U13740 (N_13740,N_13418,N_13415);
or U13741 (N_13741,N_13485,N_13588);
nor U13742 (N_13742,N_13479,N_13431);
nor U13743 (N_13743,N_13466,N_13472);
nand U13744 (N_13744,N_13582,N_13477);
nand U13745 (N_13745,N_13595,N_13438);
nor U13746 (N_13746,N_13489,N_13424);
nand U13747 (N_13747,N_13400,N_13404);
nand U13748 (N_13748,N_13445,N_13541);
and U13749 (N_13749,N_13480,N_13509);
and U13750 (N_13750,N_13585,N_13513);
nor U13751 (N_13751,N_13440,N_13553);
and U13752 (N_13752,N_13491,N_13588);
nor U13753 (N_13753,N_13570,N_13459);
or U13754 (N_13754,N_13403,N_13459);
or U13755 (N_13755,N_13407,N_13410);
nor U13756 (N_13756,N_13563,N_13532);
and U13757 (N_13757,N_13491,N_13517);
nand U13758 (N_13758,N_13538,N_13511);
or U13759 (N_13759,N_13497,N_13405);
nand U13760 (N_13760,N_13519,N_13547);
and U13761 (N_13761,N_13512,N_13528);
nand U13762 (N_13762,N_13488,N_13508);
and U13763 (N_13763,N_13528,N_13400);
nor U13764 (N_13764,N_13414,N_13437);
or U13765 (N_13765,N_13456,N_13455);
xnor U13766 (N_13766,N_13574,N_13539);
nor U13767 (N_13767,N_13483,N_13597);
nor U13768 (N_13768,N_13593,N_13531);
or U13769 (N_13769,N_13545,N_13436);
or U13770 (N_13770,N_13509,N_13441);
and U13771 (N_13771,N_13496,N_13582);
and U13772 (N_13772,N_13519,N_13582);
and U13773 (N_13773,N_13539,N_13415);
or U13774 (N_13774,N_13423,N_13516);
nand U13775 (N_13775,N_13440,N_13530);
or U13776 (N_13776,N_13470,N_13582);
and U13777 (N_13777,N_13489,N_13517);
nand U13778 (N_13778,N_13586,N_13582);
and U13779 (N_13779,N_13446,N_13587);
nor U13780 (N_13780,N_13494,N_13406);
nor U13781 (N_13781,N_13434,N_13498);
and U13782 (N_13782,N_13508,N_13565);
nor U13783 (N_13783,N_13482,N_13536);
nor U13784 (N_13784,N_13588,N_13441);
nor U13785 (N_13785,N_13563,N_13419);
and U13786 (N_13786,N_13582,N_13480);
nand U13787 (N_13787,N_13428,N_13474);
and U13788 (N_13788,N_13401,N_13510);
or U13789 (N_13789,N_13471,N_13445);
or U13790 (N_13790,N_13468,N_13467);
and U13791 (N_13791,N_13534,N_13587);
xnor U13792 (N_13792,N_13591,N_13534);
nor U13793 (N_13793,N_13581,N_13598);
nand U13794 (N_13794,N_13587,N_13415);
and U13795 (N_13795,N_13557,N_13400);
or U13796 (N_13796,N_13595,N_13401);
and U13797 (N_13797,N_13557,N_13583);
nor U13798 (N_13798,N_13546,N_13570);
nor U13799 (N_13799,N_13459,N_13532);
nor U13800 (N_13800,N_13611,N_13672);
or U13801 (N_13801,N_13681,N_13741);
xnor U13802 (N_13802,N_13605,N_13738);
nor U13803 (N_13803,N_13615,N_13773);
nand U13804 (N_13804,N_13744,N_13732);
and U13805 (N_13805,N_13616,N_13790);
or U13806 (N_13806,N_13645,N_13683);
and U13807 (N_13807,N_13708,N_13657);
and U13808 (N_13808,N_13647,N_13627);
nor U13809 (N_13809,N_13677,N_13628);
nor U13810 (N_13810,N_13685,N_13792);
and U13811 (N_13811,N_13636,N_13658);
nand U13812 (N_13812,N_13676,N_13670);
nor U13813 (N_13813,N_13669,N_13652);
or U13814 (N_13814,N_13688,N_13609);
nand U13815 (N_13815,N_13602,N_13798);
or U13816 (N_13816,N_13715,N_13735);
or U13817 (N_13817,N_13679,N_13682);
nand U13818 (N_13818,N_13728,N_13778);
or U13819 (N_13819,N_13757,N_13797);
xor U13820 (N_13820,N_13664,N_13726);
nand U13821 (N_13821,N_13651,N_13606);
nor U13822 (N_13822,N_13720,N_13603);
nor U13823 (N_13823,N_13617,N_13665);
nand U13824 (N_13824,N_13642,N_13753);
and U13825 (N_13825,N_13774,N_13764);
nor U13826 (N_13826,N_13750,N_13644);
and U13827 (N_13827,N_13694,N_13788);
nor U13828 (N_13828,N_13746,N_13663);
nor U13829 (N_13829,N_13725,N_13748);
and U13830 (N_13830,N_13678,N_13646);
and U13831 (N_13831,N_13780,N_13695);
or U13832 (N_13832,N_13643,N_13731);
nor U13833 (N_13833,N_13723,N_13624);
nor U13834 (N_13834,N_13661,N_13660);
xor U13835 (N_13835,N_13648,N_13639);
and U13836 (N_13836,N_13618,N_13742);
nor U13837 (N_13837,N_13673,N_13693);
nor U13838 (N_13838,N_13640,N_13608);
or U13839 (N_13839,N_13722,N_13671);
nand U13840 (N_13840,N_13784,N_13667);
nor U13841 (N_13841,N_13745,N_13772);
nor U13842 (N_13842,N_13633,N_13601);
and U13843 (N_13843,N_13631,N_13758);
or U13844 (N_13844,N_13783,N_13704);
nor U13845 (N_13845,N_13786,N_13674);
and U13846 (N_13846,N_13655,N_13662);
and U13847 (N_13847,N_13696,N_13637);
and U13848 (N_13848,N_13789,N_13653);
and U13849 (N_13849,N_13727,N_13641);
and U13850 (N_13850,N_13769,N_13771);
nor U13851 (N_13851,N_13762,N_13703);
or U13852 (N_13852,N_13707,N_13796);
nor U13853 (N_13853,N_13760,N_13638);
and U13854 (N_13854,N_13759,N_13779);
or U13855 (N_13855,N_13659,N_13700);
nand U13856 (N_13856,N_13743,N_13709);
nor U13857 (N_13857,N_13716,N_13724);
nand U13858 (N_13858,N_13656,N_13620);
and U13859 (N_13859,N_13791,N_13730);
nor U13860 (N_13860,N_13747,N_13739);
nand U13861 (N_13861,N_13634,N_13755);
and U13862 (N_13862,N_13719,N_13699);
nand U13863 (N_13863,N_13734,N_13721);
or U13864 (N_13864,N_13714,N_13690);
and U13865 (N_13865,N_13689,N_13754);
nor U13866 (N_13866,N_13687,N_13770);
nor U13867 (N_13867,N_13701,N_13650);
and U13868 (N_13868,N_13702,N_13710);
or U13869 (N_13869,N_13787,N_13668);
nand U13870 (N_13870,N_13782,N_13765);
or U13871 (N_13871,N_13706,N_13626);
or U13872 (N_13872,N_13621,N_13619);
nand U13873 (N_13873,N_13733,N_13756);
nand U13874 (N_13874,N_13625,N_13632);
or U13875 (N_13875,N_13691,N_13705);
or U13876 (N_13876,N_13718,N_13623);
nor U13877 (N_13877,N_13795,N_13713);
and U13878 (N_13878,N_13600,N_13785);
or U13879 (N_13879,N_13761,N_13777);
nor U13880 (N_13880,N_13799,N_13794);
nor U13881 (N_13881,N_13675,N_13712);
and U13882 (N_13882,N_13629,N_13776);
and U13883 (N_13883,N_13680,N_13768);
or U13884 (N_13884,N_13751,N_13612);
nor U13885 (N_13885,N_13767,N_13740);
nand U13886 (N_13886,N_13749,N_13684);
or U13887 (N_13887,N_13610,N_13775);
or U13888 (N_13888,N_13793,N_13763);
nand U13889 (N_13889,N_13604,N_13613);
and U13890 (N_13890,N_13711,N_13766);
and U13891 (N_13891,N_13736,N_13752);
nand U13892 (N_13892,N_13654,N_13781);
and U13893 (N_13893,N_13692,N_13697);
nor U13894 (N_13894,N_13614,N_13607);
and U13895 (N_13895,N_13666,N_13737);
and U13896 (N_13896,N_13635,N_13698);
and U13897 (N_13897,N_13729,N_13630);
and U13898 (N_13898,N_13622,N_13649);
nor U13899 (N_13899,N_13686,N_13717);
nor U13900 (N_13900,N_13634,N_13797);
and U13901 (N_13901,N_13656,N_13632);
and U13902 (N_13902,N_13779,N_13600);
nor U13903 (N_13903,N_13621,N_13735);
or U13904 (N_13904,N_13749,N_13772);
and U13905 (N_13905,N_13783,N_13705);
and U13906 (N_13906,N_13672,N_13642);
or U13907 (N_13907,N_13757,N_13784);
or U13908 (N_13908,N_13702,N_13619);
and U13909 (N_13909,N_13776,N_13784);
nor U13910 (N_13910,N_13675,N_13671);
and U13911 (N_13911,N_13778,N_13604);
and U13912 (N_13912,N_13776,N_13701);
nor U13913 (N_13913,N_13710,N_13699);
nor U13914 (N_13914,N_13650,N_13767);
or U13915 (N_13915,N_13736,N_13678);
nand U13916 (N_13916,N_13616,N_13737);
nor U13917 (N_13917,N_13772,N_13785);
nand U13918 (N_13918,N_13784,N_13770);
nand U13919 (N_13919,N_13669,N_13675);
nand U13920 (N_13920,N_13777,N_13779);
nor U13921 (N_13921,N_13751,N_13623);
and U13922 (N_13922,N_13764,N_13667);
nand U13923 (N_13923,N_13786,N_13645);
or U13924 (N_13924,N_13740,N_13787);
nor U13925 (N_13925,N_13618,N_13684);
and U13926 (N_13926,N_13636,N_13627);
or U13927 (N_13927,N_13776,N_13766);
and U13928 (N_13928,N_13788,N_13718);
and U13929 (N_13929,N_13794,N_13785);
nand U13930 (N_13930,N_13740,N_13753);
nor U13931 (N_13931,N_13784,N_13680);
and U13932 (N_13932,N_13700,N_13628);
nor U13933 (N_13933,N_13697,N_13699);
nor U13934 (N_13934,N_13732,N_13722);
nor U13935 (N_13935,N_13747,N_13659);
and U13936 (N_13936,N_13621,N_13708);
and U13937 (N_13937,N_13778,N_13708);
or U13938 (N_13938,N_13752,N_13700);
or U13939 (N_13939,N_13735,N_13698);
nor U13940 (N_13940,N_13607,N_13727);
nand U13941 (N_13941,N_13783,N_13724);
and U13942 (N_13942,N_13617,N_13691);
nand U13943 (N_13943,N_13656,N_13741);
or U13944 (N_13944,N_13634,N_13654);
nand U13945 (N_13945,N_13645,N_13623);
nand U13946 (N_13946,N_13774,N_13778);
nor U13947 (N_13947,N_13767,N_13709);
or U13948 (N_13948,N_13606,N_13770);
and U13949 (N_13949,N_13654,N_13708);
nand U13950 (N_13950,N_13684,N_13686);
nand U13951 (N_13951,N_13601,N_13671);
nand U13952 (N_13952,N_13657,N_13693);
and U13953 (N_13953,N_13657,N_13645);
xnor U13954 (N_13954,N_13694,N_13770);
and U13955 (N_13955,N_13779,N_13739);
and U13956 (N_13956,N_13698,N_13710);
or U13957 (N_13957,N_13608,N_13647);
nor U13958 (N_13958,N_13706,N_13683);
and U13959 (N_13959,N_13715,N_13623);
or U13960 (N_13960,N_13744,N_13758);
or U13961 (N_13961,N_13705,N_13697);
nand U13962 (N_13962,N_13787,N_13691);
nand U13963 (N_13963,N_13664,N_13693);
nor U13964 (N_13964,N_13676,N_13797);
or U13965 (N_13965,N_13645,N_13792);
nor U13966 (N_13966,N_13688,N_13629);
or U13967 (N_13967,N_13613,N_13733);
and U13968 (N_13968,N_13641,N_13698);
nand U13969 (N_13969,N_13701,N_13794);
or U13970 (N_13970,N_13651,N_13698);
nand U13971 (N_13971,N_13657,N_13699);
or U13972 (N_13972,N_13726,N_13761);
nor U13973 (N_13973,N_13735,N_13714);
or U13974 (N_13974,N_13668,N_13649);
or U13975 (N_13975,N_13686,N_13784);
or U13976 (N_13976,N_13677,N_13772);
nor U13977 (N_13977,N_13755,N_13743);
nor U13978 (N_13978,N_13703,N_13669);
nor U13979 (N_13979,N_13603,N_13693);
or U13980 (N_13980,N_13791,N_13741);
and U13981 (N_13981,N_13739,N_13799);
or U13982 (N_13982,N_13772,N_13705);
nor U13983 (N_13983,N_13670,N_13745);
nand U13984 (N_13984,N_13758,N_13680);
nor U13985 (N_13985,N_13749,N_13621);
and U13986 (N_13986,N_13795,N_13617);
and U13987 (N_13987,N_13615,N_13619);
nand U13988 (N_13988,N_13751,N_13727);
nand U13989 (N_13989,N_13682,N_13666);
nand U13990 (N_13990,N_13690,N_13600);
nor U13991 (N_13991,N_13659,N_13709);
nor U13992 (N_13992,N_13667,N_13686);
nand U13993 (N_13993,N_13793,N_13673);
nor U13994 (N_13994,N_13668,N_13623);
nor U13995 (N_13995,N_13705,N_13678);
nor U13996 (N_13996,N_13750,N_13607);
nor U13997 (N_13997,N_13728,N_13693);
and U13998 (N_13998,N_13776,N_13799);
or U13999 (N_13999,N_13788,N_13607);
or U14000 (N_14000,N_13814,N_13903);
or U14001 (N_14001,N_13981,N_13897);
nand U14002 (N_14002,N_13902,N_13892);
nor U14003 (N_14003,N_13907,N_13895);
and U14004 (N_14004,N_13804,N_13839);
or U14005 (N_14005,N_13972,N_13984);
nor U14006 (N_14006,N_13935,N_13945);
nor U14007 (N_14007,N_13822,N_13968);
and U14008 (N_14008,N_13857,N_13863);
and U14009 (N_14009,N_13899,N_13974);
nor U14010 (N_14010,N_13921,N_13970);
nor U14011 (N_14011,N_13813,N_13978);
and U14012 (N_14012,N_13913,N_13983);
and U14013 (N_14013,N_13993,N_13842);
nor U14014 (N_14014,N_13948,N_13964);
and U14015 (N_14015,N_13809,N_13830);
or U14016 (N_14016,N_13947,N_13800);
or U14017 (N_14017,N_13930,N_13962);
or U14018 (N_14018,N_13889,N_13908);
nor U14019 (N_14019,N_13967,N_13919);
nor U14020 (N_14020,N_13990,N_13846);
nor U14021 (N_14021,N_13823,N_13805);
nand U14022 (N_14022,N_13819,N_13987);
and U14023 (N_14023,N_13950,N_13975);
and U14024 (N_14024,N_13906,N_13838);
or U14025 (N_14025,N_13837,N_13882);
or U14026 (N_14026,N_13946,N_13808);
and U14027 (N_14027,N_13931,N_13890);
and U14028 (N_14028,N_13900,N_13992);
and U14029 (N_14029,N_13843,N_13951);
or U14030 (N_14030,N_13850,N_13957);
nand U14031 (N_14031,N_13848,N_13818);
or U14032 (N_14032,N_13924,N_13883);
and U14033 (N_14033,N_13934,N_13852);
and U14034 (N_14034,N_13965,N_13834);
nand U14035 (N_14035,N_13801,N_13923);
nand U14036 (N_14036,N_13858,N_13835);
or U14037 (N_14037,N_13932,N_13865);
nand U14038 (N_14038,N_13994,N_13942);
nor U14039 (N_14039,N_13821,N_13916);
and U14040 (N_14040,N_13910,N_13862);
and U14041 (N_14041,N_13876,N_13803);
or U14042 (N_14042,N_13954,N_13977);
or U14043 (N_14043,N_13944,N_13941);
nor U14044 (N_14044,N_13917,N_13912);
nand U14045 (N_14045,N_13922,N_13870);
nand U14046 (N_14046,N_13898,N_13991);
nand U14047 (N_14047,N_13881,N_13926);
nor U14048 (N_14048,N_13864,N_13828);
or U14049 (N_14049,N_13938,N_13896);
and U14050 (N_14050,N_13980,N_13877);
nor U14051 (N_14051,N_13979,N_13847);
nand U14052 (N_14052,N_13929,N_13911);
nand U14053 (N_14053,N_13802,N_13996);
and U14054 (N_14054,N_13920,N_13925);
and U14055 (N_14055,N_13936,N_13999);
and U14056 (N_14056,N_13836,N_13976);
nor U14057 (N_14057,N_13820,N_13867);
or U14058 (N_14058,N_13869,N_13933);
nand U14059 (N_14059,N_13998,N_13995);
nand U14060 (N_14060,N_13958,N_13855);
and U14061 (N_14061,N_13806,N_13829);
and U14062 (N_14062,N_13918,N_13937);
or U14063 (N_14063,N_13915,N_13887);
or U14064 (N_14064,N_13914,N_13956);
nor U14065 (N_14065,N_13849,N_13841);
and U14066 (N_14066,N_13810,N_13815);
nand U14067 (N_14067,N_13856,N_13961);
nor U14068 (N_14068,N_13953,N_13879);
or U14069 (N_14069,N_13986,N_13872);
nand U14070 (N_14070,N_13853,N_13817);
nand U14071 (N_14071,N_13885,N_13989);
nor U14072 (N_14072,N_13826,N_13807);
nor U14073 (N_14073,N_13878,N_13901);
or U14074 (N_14074,N_13960,N_13845);
nand U14075 (N_14075,N_13971,N_13952);
and U14076 (N_14076,N_13825,N_13955);
and U14077 (N_14077,N_13868,N_13966);
and U14078 (N_14078,N_13812,N_13927);
nand U14079 (N_14079,N_13963,N_13851);
nand U14080 (N_14080,N_13988,N_13997);
or U14081 (N_14081,N_13844,N_13840);
and U14082 (N_14082,N_13866,N_13859);
or U14083 (N_14083,N_13949,N_13940);
or U14084 (N_14084,N_13982,N_13884);
or U14085 (N_14085,N_13831,N_13873);
nand U14086 (N_14086,N_13861,N_13905);
nand U14087 (N_14087,N_13969,N_13816);
or U14088 (N_14088,N_13893,N_13985);
nand U14089 (N_14089,N_13886,N_13894);
nor U14090 (N_14090,N_13832,N_13880);
nand U14091 (N_14091,N_13973,N_13904);
nand U14092 (N_14092,N_13854,N_13874);
nand U14093 (N_14093,N_13860,N_13824);
or U14094 (N_14094,N_13888,N_13827);
or U14095 (N_14095,N_13891,N_13928);
or U14096 (N_14096,N_13959,N_13909);
or U14097 (N_14097,N_13811,N_13833);
or U14098 (N_14098,N_13939,N_13875);
and U14099 (N_14099,N_13871,N_13943);
nor U14100 (N_14100,N_13807,N_13823);
nor U14101 (N_14101,N_13903,N_13828);
or U14102 (N_14102,N_13924,N_13801);
and U14103 (N_14103,N_13910,N_13858);
nor U14104 (N_14104,N_13904,N_13986);
nor U14105 (N_14105,N_13812,N_13834);
nor U14106 (N_14106,N_13817,N_13923);
nor U14107 (N_14107,N_13807,N_13815);
nand U14108 (N_14108,N_13973,N_13952);
nand U14109 (N_14109,N_13833,N_13925);
nand U14110 (N_14110,N_13935,N_13908);
nand U14111 (N_14111,N_13997,N_13863);
nand U14112 (N_14112,N_13975,N_13881);
and U14113 (N_14113,N_13931,N_13881);
and U14114 (N_14114,N_13864,N_13816);
and U14115 (N_14115,N_13948,N_13816);
nor U14116 (N_14116,N_13818,N_13867);
or U14117 (N_14117,N_13806,N_13973);
nand U14118 (N_14118,N_13931,N_13998);
or U14119 (N_14119,N_13979,N_13900);
nor U14120 (N_14120,N_13809,N_13845);
nor U14121 (N_14121,N_13983,N_13865);
nor U14122 (N_14122,N_13802,N_13899);
or U14123 (N_14123,N_13958,N_13999);
nand U14124 (N_14124,N_13839,N_13862);
nor U14125 (N_14125,N_13990,N_13871);
nand U14126 (N_14126,N_13946,N_13965);
nor U14127 (N_14127,N_13985,N_13934);
nor U14128 (N_14128,N_13947,N_13960);
nor U14129 (N_14129,N_13894,N_13834);
and U14130 (N_14130,N_13853,N_13871);
nor U14131 (N_14131,N_13846,N_13845);
and U14132 (N_14132,N_13890,N_13809);
nand U14133 (N_14133,N_13921,N_13896);
nor U14134 (N_14134,N_13998,N_13835);
nand U14135 (N_14135,N_13929,N_13869);
nand U14136 (N_14136,N_13906,N_13831);
or U14137 (N_14137,N_13898,N_13950);
and U14138 (N_14138,N_13878,N_13988);
nor U14139 (N_14139,N_13874,N_13916);
nand U14140 (N_14140,N_13948,N_13896);
nand U14141 (N_14141,N_13808,N_13911);
nor U14142 (N_14142,N_13837,N_13975);
and U14143 (N_14143,N_13931,N_13997);
or U14144 (N_14144,N_13882,N_13802);
and U14145 (N_14145,N_13860,N_13834);
nor U14146 (N_14146,N_13819,N_13897);
or U14147 (N_14147,N_13922,N_13917);
and U14148 (N_14148,N_13969,N_13939);
nor U14149 (N_14149,N_13897,N_13863);
nor U14150 (N_14150,N_13939,N_13819);
nand U14151 (N_14151,N_13920,N_13850);
nand U14152 (N_14152,N_13972,N_13977);
or U14153 (N_14153,N_13979,N_13886);
and U14154 (N_14154,N_13821,N_13946);
nor U14155 (N_14155,N_13864,N_13888);
or U14156 (N_14156,N_13892,N_13904);
or U14157 (N_14157,N_13855,N_13901);
nand U14158 (N_14158,N_13949,N_13934);
nor U14159 (N_14159,N_13971,N_13863);
nand U14160 (N_14160,N_13994,N_13895);
or U14161 (N_14161,N_13800,N_13883);
and U14162 (N_14162,N_13912,N_13809);
and U14163 (N_14163,N_13868,N_13851);
nor U14164 (N_14164,N_13950,N_13812);
and U14165 (N_14165,N_13851,N_13824);
nor U14166 (N_14166,N_13897,N_13870);
nand U14167 (N_14167,N_13850,N_13822);
nand U14168 (N_14168,N_13831,N_13922);
or U14169 (N_14169,N_13956,N_13938);
nor U14170 (N_14170,N_13882,N_13942);
and U14171 (N_14171,N_13890,N_13842);
and U14172 (N_14172,N_13958,N_13922);
nor U14173 (N_14173,N_13999,N_13969);
nor U14174 (N_14174,N_13847,N_13875);
nand U14175 (N_14175,N_13944,N_13982);
and U14176 (N_14176,N_13835,N_13845);
nor U14177 (N_14177,N_13968,N_13990);
nor U14178 (N_14178,N_13801,N_13838);
nor U14179 (N_14179,N_13837,N_13927);
nor U14180 (N_14180,N_13858,N_13825);
nand U14181 (N_14181,N_13826,N_13920);
nor U14182 (N_14182,N_13981,N_13863);
and U14183 (N_14183,N_13941,N_13803);
nor U14184 (N_14184,N_13925,N_13997);
or U14185 (N_14185,N_13893,N_13803);
nand U14186 (N_14186,N_13930,N_13831);
and U14187 (N_14187,N_13939,N_13903);
nand U14188 (N_14188,N_13888,N_13899);
nor U14189 (N_14189,N_13957,N_13849);
and U14190 (N_14190,N_13842,N_13840);
nand U14191 (N_14191,N_13954,N_13903);
or U14192 (N_14192,N_13981,N_13889);
or U14193 (N_14193,N_13974,N_13972);
and U14194 (N_14194,N_13999,N_13887);
or U14195 (N_14195,N_13859,N_13871);
or U14196 (N_14196,N_13861,N_13962);
and U14197 (N_14197,N_13998,N_13907);
nand U14198 (N_14198,N_13838,N_13805);
and U14199 (N_14199,N_13894,N_13857);
nor U14200 (N_14200,N_14016,N_14102);
and U14201 (N_14201,N_14034,N_14074);
nor U14202 (N_14202,N_14076,N_14081);
or U14203 (N_14203,N_14132,N_14199);
or U14204 (N_14204,N_14092,N_14111);
and U14205 (N_14205,N_14066,N_14113);
nand U14206 (N_14206,N_14163,N_14156);
nor U14207 (N_14207,N_14108,N_14017);
and U14208 (N_14208,N_14121,N_14170);
xnor U14209 (N_14209,N_14126,N_14174);
nor U14210 (N_14210,N_14166,N_14041);
nor U14211 (N_14211,N_14117,N_14114);
nor U14212 (N_14212,N_14173,N_14019);
or U14213 (N_14213,N_14013,N_14031);
and U14214 (N_14214,N_14022,N_14128);
or U14215 (N_14215,N_14079,N_14195);
nand U14216 (N_14216,N_14142,N_14043);
or U14217 (N_14217,N_14042,N_14062);
nand U14218 (N_14218,N_14065,N_14136);
nand U14219 (N_14219,N_14159,N_14137);
nor U14220 (N_14220,N_14165,N_14140);
or U14221 (N_14221,N_14009,N_14014);
nor U14222 (N_14222,N_14011,N_14098);
xor U14223 (N_14223,N_14033,N_14026);
or U14224 (N_14224,N_14146,N_14025);
nand U14225 (N_14225,N_14095,N_14130);
nand U14226 (N_14226,N_14143,N_14070);
nand U14227 (N_14227,N_14105,N_14197);
or U14228 (N_14228,N_14162,N_14188);
or U14229 (N_14229,N_14010,N_14157);
or U14230 (N_14230,N_14002,N_14180);
nand U14231 (N_14231,N_14153,N_14171);
nor U14232 (N_14232,N_14115,N_14110);
xor U14233 (N_14233,N_14052,N_14064);
nor U14234 (N_14234,N_14183,N_14134);
nand U14235 (N_14235,N_14067,N_14029);
xor U14236 (N_14236,N_14127,N_14186);
and U14237 (N_14237,N_14055,N_14191);
or U14238 (N_14238,N_14104,N_14051);
or U14239 (N_14239,N_14119,N_14151);
and U14240 (N_14240,N_14000,N_14047);
nand U14241 (N_14241,N_14129,N_14172);
nand U14242 (N_14242,N_14040,N_14145);
and U14243 (N_14243,N_14012,N_14150);
and U14244 (N_14244,N_14054,N_14085);
nor U14245 (N_14245,N_14155,N_14109);
nand U14246 (N_14246,N_14048,N_14141);
nand U14247 (N_14247,N_14160,N_14027);
xor U14248 (N_14248,N_14139,N_14090);
and U14249 (N_14249,N_14032,N_14149);
and U14250 (N_14250,N_14124,N_14101);
or U14251 (N_14251,N_14023,N_14072);
nor U14252 (N_14252,N_14168,N_14189);
nor U14253 (N_14253,N_14030,N_14063);
nand U14254 (N_14254,N_14148,N_14046);
and U14255 (N_14255,N_14039,N_14169);
nor U14256 (N_14256,N_14167,N_14177);
and U14257 (N_14257,N_14103,N_14122);
nand U14258 (N_14258,N_14193,N_14107);
nor U14259 (N_14259,N_14049,N_14087);
nor U14260 (N_14260,N_14158,N_14196);
and U14261 (N_14261,N_14198,N_14161);
nand U14262 (N_14262,N_14091,N_14094);
nor U14263 (N_14263,N_14083,N_14015);
or U14264 (N_14264,N_14018,N_14020);
nor U14265 (N_14265,N_14069,N_14123);
nand U14266 (N_14266,N_14006,N_14133);
or U14267 (N_14267,N_14024,N_14135);
nand U14268 (N_14268,N_14021,N_14037);
or U14269 (N_14269,N_14097,N_14008);
nor U14270 (N_14270,N_14053,N_14112);
nand U14271 (N_14271,N_14154,N_14088);
nor U14272 (N_14272,N_14185,N_14131);
nand U14273 (N_14273,N_14116,N_14082);
or U14274 (N_14274,N_14038,N_14073);
nand U14275 (N_14275,N_14084,N_14061);
nand U14276 (N_14276,N_14138,N_14007);
nand U14277 (N_14277,N_14176,N_14075);
and U14278 (N_14278,N_14175,N_14181);
nor U14279 (N_14279,N_14118,N_14096);
or U14280 (N_14280,N_14147,N_14144);
and U14281 (N_14281,N_14100,N_14093);
and U14282 (N_14282,N_14068,N_14152);
nand U14283 (N_14283,N_14099,N_14089);
nor U14284 (N_14284,N_14192,N_14071);
or U14285 (N_14285,N_14077,N_14001);
or U14286 (N_14286,N_14086,N_14182);
or U14287 (N_14287,N_14036,N_14028);
nor U14288 (N_14288,N_14003,N_14004);
nand U14289 (N_14289,N_14035,N_14190);
nand U14290 (N_14290,N_14005,N_14106);
and U14291 (N_14291,N_14060,N_14044);
nand U14292 (N_14292,N_14057,N_14058);
nor U14293 (N_14293,N_14059,N_14120);
nand U14294 (N_14294,N_14164,N_14080);
nor U14295 (N_14295,N_14179,N_14194);
and U14296 (N_14296,N_14184,N_14056);
nor U14297 (N_14297,N_14187,N_14178);
and U14298 (N_14298,N_14078,N_14125);
nand U14299 (N_14299,N_14045,N_14050);
or U14300 (N_14300,N_14007,N_14133);
nor U14301 (N_14301,N_14181,N_14008);
nor U14302 (N_14302,N_14166,N_14130);
or U14303 (N_14303,N_14120,N_14030);
or U14304 (N_14304,N_14109,N_14175);
or U14305 (N_14305,N_14035,N_14177);
and U14306 (N_14306,N_14128,N_14122);
nor U14307 (N_14307,N_14136,N_14018);
and U14308 (N_14308,N_14126,N_14014);
nor U14309 (N_14309,N_14166,N_14071);
nor U14310 (N_14310,N_14065,N_14029);
nor U14311 (N_14311,N_14098,N_14056);
or U14312 (N_14312,N_14150,N_14179);
nand U14313 (N_14313,N_14192,N_14157);
and U14314 (N_14314,N_14029,N_14084);
nor U14315 (N_14315,N_14117,N_14168);
or U14316 (N_14316,N_14091,N_14007);
nor U14317 (N_14317,N_14036,N_14173);
or U14318 (N_14318,N_14172,N_14184);
or U14319 (N_14319,N_14118,N_14038);
or U14320 (N_14320,N_14001,N_14110);
or U14321 (N_14321,N_14049,N_14156);
or U14322 (N_14322,N_14105,N_14177);
or U14323 (N_14323,N_14151,N_14004);
nand U14324 (N_14324,N_14181,N_14064);
and U14325 (N_14325,N_14066,N_14014);
nor U14326 (N_14326,N_14177,N_14042);
nor U14327 (N_14327,N_14024,N_14161);
nand U14328 (N_14328,N_14153,N_14199);
nand U14329 (N_14329,N_14174,N_14147);
and U14330 (N_14330,N_14170,N_14092);
or U14331 (N_14331,N_14177,N_14031);
and U14332 (N_14332,N_14187,N_14183);
and U14333 (N_14333,N_14076,N_14052);
and U14334 (N_14334,N_14167,N_14121);
nor U14335 (N_14335,N_14052,N_14041);
and U14336 (N_14336,N_14121,N_14020);
and U14337 (N_14337,N_14004,N_14021);
nand U14338 (N_14338,N_14026,N_14191);
or U14339 (N_14339,N_14139,N_14093);
or U14340 (N_14340,N_14181,N_14009);
and U14341 (N_14341,N_14150,N_14176);
nand U14342 (N_14342,N_14128,N_14000);
and U14343 (N_14343,N_14005,N_14063);
or U14344 (N_14344,N_14010,N_14084);
or U14345 (N_14345,N_14047,N_14009);
nand U14346 (N_14346,N_14180,N_14117);
nand U14347 (N_14347,N_14063,N_14100);
nand U14348 (N_14348,N_14132,N_14049);
and U14349 (N_14349,N_14126,N_14033);
and U14350 (N_14350,N_14129,N_14097);
or U14351 (N_14351,N_14114,N_14046);
or U14352 (N_14352,N_14119,N_14122);
nand U14353 (N_14353,N_14132,N_14009);
nand U14354 (N_14354,N_14139,N_14088);
nor U14355 (N_14355,N_14039,N_14185);
nor U14356 (N_14356,N_14022,N_14183);
nor U14357 (N_14357,N_14062,N_14073);
and U14358 (N_14358,N_14139,N_14014);
and U14359 (N_14359,N_14128,N_14117);
or U14360 (N_14360,N_14123,N_14028);
nand U14361 (N_14361,N_14118,N_14049);
or U14362 (N_14362,N_14126,N_14086);
nor U14363 (N_14363,N_14179,N_14070);
and U14364 (N_14364,N_14000,N_14174);
nand U14365 (N_14365,N_14161,N_14129);
nand U14366 (N_14366,N_14196,N_14199);
or U14367 (N_14367,N_14006,N_14176);
and U14368 (N_14368,N_14031,N_14128);
nor U14369 (N_14369,N_14194,N_14121);
nor U14370 (N_14370,N_14046,N_14065);
or U14371 (N_14371,N_14015,N_14134);
and U14372 (N_14372,N_14043,N_14049);
nand U14373 (N_14373,N_14085,N_14082);
or U14374 (N_14374,N_14114,N_14106);
or U14375 (N_14375,N_14021,N_14199);
and U14376 (N_14376,N_14100,N_14083);
nand U14377 (N_14377,N_14154,N_14135);
or U14378 (N_14378,N_14116,N_14020);
or U14379 (N_14379,N_14143,N_14174);
and U14380 (N_14380,N_14179,N_14011);
or U14381 (N_14381,N_14108,N_14198);
nor U14382 (N_14382,N_14067,N_14002);
nor U14383 (N_14383,N_14151,N_14023);
and U14384 (N_14384,N_14196,N_14069);
or U14385 (N_14385,N_14171,N_14024);
nand U14386 (N_14386,N_14001,N_14108);
or U14387 (N_14387,N_14068,N_14010);
and U14388 (N_14388,N_14135,N_14184);
xnor U14389 (N_14389,N_14021,N_14091);
and U14390 (N_14390,N_14030,N_14130);
nor U14391 (N_14391,N_14154,N_14024);
xor U14392 (N_14392,N_14060,N_14169);
and U14393 (N_14393,N_14101,N_14100);
nand U14394 (N_14394,N_14146,N_14199);
nor U14395 (N_14395,N_14003,N_14167);
nor U14396 (N_14396,N_14040,N_14068);
nor U14397 (N_14397,N_14143,N_14077);
nor U14398 (N_14398,N_14114,N_14018);
nor U14399 (N_14399,N_14156,N_14038);
and U14400 (N_14400,N_14287,N_14244);
nand U14401 (N_14401,N_14211,N_14210);
nand U14402 (N_14402,N_14222,N_14390);
nor U14403 (N_14403,N_14351,N_14288);
nor U14404 (N_14404,N_14346,N_14265);
nand U14405 (N_14405,N_14345,N_14201);
and U14406 (N_14406,N_14236,N_14282);
nor U14407 (N_14407,N_14347,N_14270);
or U14408 (N_14408,N_14259,N_14297);
and U14409 (N_14409,N_14387,N_14310);
or U14410 (N_14410,N_14314,N_14344);
and U14411 (N_14411,N_14227,N_14311);
and U14412 (N_14412,N_14257,N_14235);
and U14413 (N_14413,N_14367,N_14376);
nor U14414 (N_14414,N_14340,N_14226);
and U14415 (N_14415,N_14234,N_14299);
and U14416 (N_14416,N_14219,N_14321);
nor U14417 (N_14417,N_14341,N_14377);
nand U14418 (N_14418,N_14334,N_14372);
or U14419 (N_14419,N_14363,N_14212);
nor U14420 (N_14420,N_14239,N_14271);
nand U14421 (N_14421,N_14286,N_14399);
nand U14422 (N_14422,N_14240,N_14263);
nor U14423 (N_14423,N_14221,N_14216);
xor U14424 (N_14424,N_14229,N_14357);
nor U14425 (N_14425,N_14230,N_14324);
or U14426 (N_14426,N_14237,N_14252);
or U14427 (N_14427,N_14248,N_14253);
or U14428 (N_14428,N_14379,N_14382);
and U14429 (N_14429,N_14220,N_14395);
or U14430 (N_14430,N_14262,N_14392);
and U14431 (N_14431,N_14348,N_14213);
or U14432 (N_14432,N_14200,N_14255);
nand U14433 (N_14433,N_14251,N_14264);
nor U14434 (N_14434,N_14336,N_14293);
nand U14435 (N_14435,N_14319,N_14375);
nand U14436 (N_14436,N_14396,N_14300);
and U14437 (N_14437,N_14355,N_14394);
or U14438 (N_14438,N_14241,N_14281);
and U14439 (N_14439,N_14327,N_14374);
nor U14440 (N_14440,N_14381,N_14242);
and U14441 (N_14441,N_14247,N_14283);
nor U14442 (N_14442,N_14384,N_14391);
and U14443 (N_14443,N_14209,N_14385);
and U14444 (N_14444,N_14315,N_14316);
or U14445 (N_14445,N_14388,N_14302);
nand U14446 (N_14446,N_14368,N_14250);
nor U14447 (N_14447,N_14215,N_14232);
nand U14448 (N_14448,N_14223,N_14290);
nand U14449 (N_14449,N_14218,N_14266);
or U14450 (N_14450,N_14366,N_14380);
nor U14451 (N_14451,N_14398,N_14339);
nand U14452 (N_14452,N_14225,N_14360);
nand U14453 (N_14453,N_14298,N_14205);
and U14454 (N_14454,N_14304,N_14294);
or U14455 (N_14455,N_14356,N_14279);
and U14456 (N_14456,N_14397,N_14231);
nand U14457 (N_14457,N_14260,N_14343);
and U14458 (N_14458,N_14268,N_14358);
or U14459 (N_14459,N_14291,N_14272);
and U14460 (N_14460,N_14280,N_14354);
and U14461 (N_14461,N_14386,N_14254);
nand U14462 (N_14462,N_14329,N_14275);
nor U14463 (N_14463,N_14325,N_14238);
nor U14464 (N_14464,N_14365,N_14370);
nand U14465 (N_14465,N_14217,N_14258);
or U14466 (N_14466,N_14371,N_14362);
or U14467 (N_14467,N_14317,N_14331);
or U14468 (N_14468,N_14246,N_14301);
and U14469 (N_14469,N_14308,N_14233);
nor U14470 (N_14470,N_14249,N_14278);
and U14471 (N_14471,N_14276,N_14361);
nor U14472 (N_14472,N_14277,N_14228);
or U14473 (N_14473,N_14292,N_14338);
and U14474 (N_14474,N_14330,N_14323);
nand U14475 (N_14475,N_14332,N_14284);
or U14476 (N_14476,N_14349,N_14295);
nand U14477 (N_14477,N_14364,N_14359);
and U14478 (N_14478,N_14383,N_14378);
nor U14479 (N_14479,N_14369,N_14273);
or U14480 (N_14480,N_14322,N_14352);
nor U14481 (N_14481,N_14208,N_14305);
or U14482 (N_14482,N_14202,N_14224);
nor U14483 (N_14483,N_14389,N_14393);
nor U14484 (N_14484,N_14313,N_14207);
nor U14485 (N_14485,N_14289,N_14342);
nand U14486 (N_14486,N_14326,N_14269);
and U14487 (N_14487,N_14307,N_14296);
nand U14488 (N_14488,N_14214,N_14337);
nand U14489 (N_14489,N_14320,N_14206);
or U14490 (N_14490,N_14309,N_14267);
nor U14491 (N_14491,N_14303,N_14312);
nor U14492 (N_14492,N_14335,N_14245);
or U14493 (N_14493,N_14261,N_14350);
and U14494 (N_14494,N_14306,N_14274);
or U14495 (N_14495,N_14328,N_14203);
nor U14496 (N_14496,N_14333,N_14353);
or U14497 (N_14497,N_14256,N_14285);
or U14498 (N_14498,N_14318,N_14243);
or U14499 (N_14499,N_14373,N_14204);
or U14500 (N_14500,N_14366,N_14207);
or U14501 (N_14501,N_14272,N_14384);
nand U14502 (N_14502,N_14236,N_14201);
or U14503 (N_14503,N_14250,N_14284);
nand U14504 (N_14504,N_14284,N_14216);
and U14505 (N_14505,N_14364,N_14232);
nand U14506 (N_14506,N_14330,N_14297);
and U14507 (N_14507,N_14306,N_14335);
or U14508 (N_14508,N_14228,N_14211);
nor U14509 (N_14509,N_14245,N_14240);
and U14510 (N_14510,N_14209,N_14221);
or U14511 (N_14511,N_14203,N_14215);
nand U14512 (N_14512,N_14269,N_14386);
nand U14513 (N_14513,N_14259,N_14280);
nand U14514 (N_14514,N_14393,N_14388);
nor U14515 (N_14515,N_14361,N_14387);
and U14516 (N_14516,N_14292,N_14378);
nor U14517 (N_14517,N_14239,N_14282);
or U14518 (N_14518,N_14356,N_14399);
and U14519 (N_14519,N_14344,N_14368);
nor U14520 (N_14520,N_14345,N_14233);
nor U14521 (N_14521,N_14253,N_14226);
nand U14522 (N_14522,N_14244,N_14317);
and U14523 (N_14523,N_14372,N_14399);
nand U14524 (N_14524,N_14359,N_14330);
and U14525 (N_14525,N_14285,N_14200);
nand U14526 (N_14526,N_14242,N_14231);
xor U14527 (N_14527,N_14394,N_14379);
or U14528 (N_14528,N_14308,N_14392);
nand U14529 (N_14529,N_14251,N_14213);
and U14530 (N_14530,N_14253,N_14249);
and U14531 (N_14531,N_14382,N_14326);
and U14532 (N_14532,N_14264,N_14368);
nor U14533 (N_14533,N_14336,N_14255);
nor U14534 (N_14534,N_14357,N_14392);
and U14535 (N_14535,N_14389,N_14337);
nor U14536 (N_14536,N_14227,N_14329);
and U14537 (N_14537,N_14344,N_14384);
or U14538 (N_14538,N_14291,N_14280);
and U14539 (N_14539,N_14341,N_14309);
or U14540 (N_14540,N_14276,N_14295);
nand U14541 (N_14541,N_14388,N_14238);
and U14542 (N_14542,N_14262,N_14271);
nor U14543 (N_14543,N_14388,N_14283);
or U14544 (N_14544,N_14238,N_14314);
nand U14545 (N_14545,N_14375,N_14347);
or U14546 (N_14546,N_14348,N_14221);
xnor U14547 (N_14547,N_14220,N_14291);
and U14548 (N_14548,N_14202,N_14387);
nor U14549 (N_14549,N_14291,N_14253);
nor U14550 (N_14550,N_14380,N_14236);
and U14551 (N_14551,N_14275,N_14394);
and U14552 (N_14552,N_14365,N_14342);
nand U14553 (N_14553,N_14227,N_14392);
nor U14554 (N_14554,N_14273,N_14223);
nor U14555 (N_14555,N_14209,N_14273);
and U14556 (N_14556,N_14277,N_14301);
nor U14557 (N_14557,N_14274,N_14228);
nand U14558 (N_14558,N_14352,N_14317);
or U14559 (N_14559,N_14299,N_14235);
or U14560 (N_14560,N_14367,N_14342);
or U14561 (N_14561,N_14309,N_14371);
and U14562 (N_14562,N_14300,N_14216);
nor U14563 (N_14563,N_14270,N_14377);
and U14564 (N_14564,N_14366,N_14378);
xor U14565 (N_14565,N_14383,N_14259);
nand U14566 (N_14566,N_14396,N_14204);
and U14567 (N_14567,N_14236,N_14288);
nor U14568 (N_14568,N_14309,N_14378);
or U14569 (N_14569,N_14200,N_14353);
or U14570 (N_14570,N_14289,N_14317);
nor U14571 (N_14571,N_14296,N_14203);
nor U14572 (N_14572,N_14356,N_14331);
nand U14573 (N_14573,N_14269,N_14317);
or U14574 (N_14574,N_14248,N_14305);
nor U14575 (N_14575,N_14204,N_14256);
xor U14576 (N_14576,N_14285,N_14303);
nor U14577 (N_14577,N_14328,N_14387);
or U14578 (N_14578,N_14304,N_14334);
and U14579 (N_14579,N_14371,N_14245);
nand U14580 (N_14580,N_14308,N_14205);
and U14581 (N_14581,N_14355,N_14277);
or U14582 (N_14582,N_14266,N_14264);
or U14583 (N_14583,N_14329,N_14261);
nor U14584 (N_14584,N_14307,N_14278);
nor U14585 (N_14585,N_14359,N_14360);
nor U14586 (N_14586,N_14208,N_14397);
and U14587 (N_14587,N_14374,N_14358);
nand U14588 (N_14588,N_14397,N_14304);
and U14589 (N_14589,N_14326,N_14210);
or U14590 (N_14590,N_14338,N_14227);
and U14591 (N_14591,N_14247,N_14203);
nand U14592 (N_14592,N_14221,N_14358);
nor U14593 (N_14593,N_14279,N_14383);
or U14594 (N_14594,N_14298,N_14262);
or U14595 (N_14595,N_14391,N_14261);
nor U14596 (N_14596,N_14325,N_14358);
nor U14597 (N_14597,N_14368,N_14251);
nor U14598 (N_14598,N_14338,N_14334);
or U14599 (N_14599,N_14392,N_14367);
or U14600 (N_14600,N_14423,N_14457);
nand U14601 (N_14601,N_14436,N_14435);
nand U14602 (N_14602,N_14554,N_14520);
and U14603 (N_14603,N_14555,N_14408);
nand U14604 (N_14604,N_14533,N_14420);
and U14605 (N_14605,N_14479,N_14425);
or U14606 (N_14606,N_14483,N_14539);
or U14607 (N_14607,N_14490,N_14442);
nand U14608 (N_14608,N_14424,N_14407);
or U14609 (N_14609,N_14585,N_14411);
and U14610 (N_14610,N_14596,N_14454);
and U14611 (N_14611,N_14513,N_14584);
and U14612 (N_14612,N_14571,N_14519);
nor U14613 (N_14613,N_14589,N_14417);
nand U14614 (N_14614,N_14561,N_14484);
and U14615 (N_14615,N_14403,N_14450);
nand U14616 (N_14616,N_14598,N_14530);
or U14617 (N_14617,N_14400,N_14540);
nand U14618 (N_14618,N_14488,N_14577);
or U14619 (N_14619,N_14578,N_14437);
xnor U14620 (N_14620,N_14545,N_14592);
and U14621 (N_14621,N_14498,N_14458);
or U14622 (N_14622,N_14544,N_14568);
nor U14623 (N_14623,N_14579,N_14494);
nand U14624 (N_14624,N_14537,N_14444);
xnor U14625 (N_14625,N_14469,N_14470);
nor U14626 (N_14626,N_14431,N_14466);
nand U14627 (N_14627,N_14413,N_14524);
or U14628 (N_14628,N_14414,N_14416);
or U14629 (N_14629,N_14507,N_14471);
nand U14630 (N_14630,N_14587,N_14499);
and U14631 (N_14631,N_14401,N_14570);
and U14632 (N_14632,N_14556,N_14505);
or U14633 (N_14633,N_14586,N_14560);
nand U14634 (N_14634,N_14452,N_14481);
nor U14635 (N_14635,N_14482,N_14468);
nand U14636 (N_14636,N_14445,N_14492);
nand U14637 (N_14637,N_14493,N_14406);
and U14638 (N_14638,N_14478,N_14551);
and U14639 (N_14639,N_14575,N_14572);
nor U14640 (N_14640,N_14448,N_14449);
or U14641 (N_14641,N_14434,N_14566);
or U14642 (N_14642,N_14441,N_14569);
nand U14643 (N_14643,N_14538,N_14595);
or U14644 (N_14644,N_14504,N_14421);
or U14645 (N_14645,N_14463,N_14459);
and U14646 (N_14646,N_14467,N_14546);
xor U14647 (N_14647,N_14429,N_14487);
and U14648 (N_14648,N_14590,N_14548);
nand U14649 (N_14649,N_14502,N_14562);
xor U14650 (N_14650,N_14426,N_14485);
or U14651 (N_14651,N_14509,N_14486);
nor U14652 (N_14652,N_14491,N_14588);
or U14653 (N_14653,N_14440,N_14525);
nand U14654 (N_14654,N_14432,N_14541);
or U14655 (N_14655,N_14433,N_14419);
nor U14656 (N_14656,N_14547,N_14460);
nor U14657 (N_14657,N_14564,N_14543);
or U14658 (N_14658,N_14476,N_14402);
and U14659 (N_14659,N_14550,N_14517);
or U14660 (N_14660,N_14582,N_14472);
nand U14661 (N_14661,N_14514,N_14412);
nor U14662 (N_14662,N_14512,N_14522);
and U14663 (N_14663,N_14516,N_14573);
and U14664 (N_14664,N_14574,N_14558);
and U14665 (N_14665,N_14405,N_14511);
nor U14666 (N_14666,N_14475,N_14581);
nor U14667 (N_14667,N_14559,N_14456);
nor U14668 (N_14668,N_14536,N_14480);
or U14669 (N_14669,N_14534,N_14528);
nand U14670 (N_14670,N_14462,N_14474);
or U14671 (N_14671,N_14529,N_14497);
and U14672 (N_14672,N_14409,N_14477);
and U14673 (N_14673,N_14500,N_14489);
nor U14674 (N_14674,N_14535,N_14438);
nor U14675 (N_14675,N_14418,N_14567);
nand U14676 (N_14676,N_14597,N_14427);
nand U14677 (N_14677,N_14552,N_14549);
and U14678 (N_14678,N_14518,N_14542);
or U14679 (N_14679,N_14565,N_14508);
nor U14680 (N_14680,N_14446,N_14515);
nor U14681 (N_14681,N_14523,N_14422);
or U14682 (N_14682,N_14594,N_14591);
nand U14683 (N_14683,N_14593,N_14410);
and U14684 (N_14684,N_14451,N_14428);
or U14685 (N_14685,N_14461,N_14453);
or U14686 (N_14686,N_14430,N_14415);
nor U14687 (N_14687,N_14580,N_14439);
and U14688 (N_14688,N_14473,N_14443);
and U14689 (N_14689,N_14506,N_14501);
nand U14690 (N_14690,N_14521,N_14447);
nand U14691 (N_14691,N_14464,N_14599);
and U14692 (N_14692,N_14553,N_14503);
nor U14693 (N_14693,N_14557,N_14532);
nor U14694 (N_14694,N_14496,N_14531);
or U14695 (N_14695,N_14583,N_14404);
and U14696 (N_14696,N_14563,N_14527);
or U14697 (N_14697,N_14510,N_14526);
nor U14698 (N_14698,N_14455,N_14576);
and U14699 (N_14699,N_14465,N_14495);
nand U14700 (N_14700,N_14482,N_14484);
and U14701 (N_14701,N_14485,N_14526);
nor U14702 (N_14702,N_14485,N_14565);
nand U14703 (N_14703,N_14405,N_14554);
nor U14704 (N_14704,N_14469,N_14408);
nand U14705 (N_14705,N_14598,N_14550);
nand U14706 (N_14706,N_14466,N_14550);
nor U14707 (N_14707,N_14542,N_14496);
or U14708 (N_14708,N_14547,N_14563);
nor U14709 (N_14709,N_14526,N_14448);
nand U14710 (N_14710,N_14565,N_14577);
nand U14711 (N_14711,N_14437,N_14467);
nand U14712 (N_14712,N_14496,N_14420);
nor U14713 (N_14713,N_14412,N_14565);
nand U14714 (N_14714,N_14433,N_14540);
or U14715 (N_14715,N_14476,N_14576);
nand U14716 (N_14716,N_14538,N_14424);
and U14717 (N_14717,N_14494,N_14405);
nand U14718 (N_14718,N_14472,N_14527);
or U14719 (N_14719,N_14515,N_14507);
and U14720 (N_14720,N_14477,N_14499);
or U14721 (N_14721,N_14477,N_14445);
nand U14722 (N_14722,N_14503,N_14521);
and U14723 (N_14723,N_14505,N_14594);
nand U14724 (N_14724,N_14573,N_14451);
nor U14725 (N_14725,N_14404,N_14431);
nand U14726 (N_14726,N_14563,N_14562);
nand U14727 (N_14727,N_14469,N_14504);
and U14728 (N_14728,N_14569,N_14514);
or U14729 (N_14729,N_14487,N_14592);
nand U14730 (N_14730,N_14533,N_14538);
or U14731 (N_14731,N_14410,N_14512);
and U14732 (N_14732,N_14516,N_14591);
nand U14733 (N_14733,N_14485,N_14520);
nand U14734 (N_14734,N_14453,N_14571);
nor U14735 (N_14735,N_14502,N_14416);
or U14736 (N_14736,N_14524,N_14454);
or U14737 (N_14737,N_14513,N_14512);
and U14738 (N_14738,N_14431,N_14547);
nor U14739 (N_14739,N_14461,N_14472);
nor U14740 (N_14740,N_14585,N_14444);
and U14741 (N_14741,N_14477,N_14581);
nor U14742 (N_14742,N_14575,N_14442);
or U14743 (N_14743,N_14486,N_14597);
nor U14744 (N_14744,N_14553,N_14560);
and U14745 (N_14745,N_14577,N_14549);
or U14746 (N_14746,N_14547,N_14582);
and U14747 (N_14747,N_14591,N_14444);
nor U14748 (N_14748,N_14427,N_14524);
and U14749 (N_14749,N_14573,N_14517);
nor U14750 (N_14750,N_14498,N_14496);
or U14751 (N_14751,N_14420,N_14583);
nor U14752 (N_14752,N_14544,N_14466);
and U14753 (N_14753,N_14415,N_14411);
and U14754 (N_14754,N_14486,N_14446);
and U14755 (N_14755,N_14551,N_14499);
nand U14756 (N_14756,N_14498,N_14526);
xnor U14757 (N_14757,N_14551,N_14464);
nand U14758 (N_14758,N_14489,N_14433);
and U14759 (N_14759,N_14537,N_14522);
nand U14760 (N_14760,N_14455,N_14563);
nand U14761 (N_14761,N_14560,N_14411);
nand U14762 (N_14762,N_14461,N_14503);
nor U14763 (N_14763,N_14426,N_14572);
and U14764 (N_14764,N_14550,N_14472);
nor U14765 (N_14765,N_14534,N_14539);
nor U14766 (N_14766,N_14497,N_14484);
or U14767 (N_14767,N_14560,N_14508);
nand U14768 (N_14768,N_14457,N_14572);
nand U14769 (N_14769,N_14552,N_14401);
nor U14770 (N_14770,N_14428,N_14482);
nor U14771 (N_14771,N_14428,N_14518);
nor U14772 (N_14772,N_14529,N_14502);
or U14773 (N_14773,N_14449,N_14571);
or U14774 (N_14774,N_14406,N_14557);
or U14775 (N_14775,N_14401,N_14472);
nand U14776 (N_14776,N_14447,N_14551);
nand U14777 (N_14777,N_14592,N_14503);
nor U14778 (N_14778,N_14514,N_14457);
and U14779 (N_14779,N_14521,N_14569);
and U14780 (N_14780,N_14496,N_14560);
or U14781 (N_14781,N_14439,N_14523);
nand U14782 (N_14782,N_14583,N_14400);
and U14783 (N_14783,N_14590,N_14545);
nand U14784 (N_14784,N_14594,N_14468);
or U14785 (N_14785,N_14504,N_14546);
nor U14786 (N_14786,N_14444,N_14463);
nor U14787 (N_14787,N_14409,N_14436);
and U14788 (N_14788,N_14487,N_14427);
and U14789 (N_14789,N_14500,N_14460);
nand U14790 (N_14790,N_14460,N_14596);
and U14791 (N_14791,N_14419,N_14597);
and U14792 (N_14792,N_14452,N_14464);
nor U14793 (N_14793,N_14436,N_14524);
nand U14794 (N_14794,N_14557,N_14461);
and U14795 (N_14795,N_14493,N_14419);
nand U14796 (N_14796,N_14525,N_14528);
xnor U14797 (N_14797,N_14454,N_14459);
nand U14798 (N_14798,N_14532,N_14589);
nand U14799 (N_14799,N_14518,N_14440);
nor U14800 (N_14800,N_14750,N_14747);
and U14801 (N_14801,N_14693,N_14777);
or U14802 (N_14802,N_14645,N_14782);
nor U14803 (N_14803,N_14602,N_14752);
nor U14804 (N_14804,N_14657,N_14624);
nor U14805 (N_14805,N_14637,N_14716);
and U14806 (N_14806,N_14712,N_14700);
and U14807 (N_14807,N_14779,N_14688);
nor U14808 (N_14808,N_14607,N_14691);
or U14809 (N_14809,N_14652,N_14765);
and U14810 (N_14810,N_14695,N_14708);
or U14811 (N_14811,N_14687,N_14668);
nand U14812 (N_14812,N_14612,N_14773);
or U14813 (N_14813,N_14741,N_14678);
nor U14814 (N_14814,N_14726,N_14684);
nand U14815 (N_14815,N_14648,N_14659);
xnor U14816 (N_14816,N_14640,N_14646);
or U14817 (N_14817,N_14758,N_14605);
or U14818 (N_14818,N_14766,N_14699);
nor U14819 (N_14819,N_14757,N_14626);
nand U14820 (N_14820,N_14698,N_14743);
and U14821 (N_14821,N_14799,N_14650);
nor U14822 (N_14822,N_14636,N_14690);
nor U14823 (N_14823,N_14654,N_14729);
and U14824 (N_14824,N_14744,N_14632);
or U14825 (N_14825,N_14673,N_14732);
nor U14826 (N_14826,N_14711,N_14679);
nand U14827 (N_14827,N_14694,N_14721);
nand U14828 (N_14828,N_14745,N_14728);
nand U14829 (N_14829,N_14756,N_14629);
nand U14830 (N_14830,N_14770,N_14763);
nand U14831 (N_14831,N_14725,N_14760);
nor U14832 (N_14832,N_14786,N_14754);
or U14833 (N_14833,N_14735,N_14670);
and U14834 (N_14834,N_14739,N_14781);
and U14835 (N_14835,N_14671,N_14720);
and U14836 (N_14836,N_14748,N_14715);
nand U14837 (N_14837,N_14617,N_14669);
or U14838 (N_14838,N_14697,N_14610);
nor U14839 (N_14839,N_14631,N_14794);
nand U14840 (N_14840,N_14738,N_14666);
or U14841 (N_14841,N_14603,N_14775);
or U14842 (N_14842,N_14641,N_14730);
and U14843 (N_14843,N_14740,N_14622);
nor U14844 (N_14844,N_14649,N_14642);
and U14845 (N_14845,N_14625,N_14772);
nand U14846 (N_14846,N_14790,N_14664);
nand U14847 (N_14847,N_14681,N_14707);
nand U14848 (N_14848,N_14701,N_14719);
nor U14849 (N_14849,N_14616,N_14736);
and U14850 (N_14850,N_14660,N_14686);
or U14851 (N_14851,N_14768,N_14651);
nor U14852 (N_14852,N_14703,N_14611);
or U14853 (N_14853,N_14621,N_14710);
nor U14854 (N_14854,N_14665,N_14737);
or U14855 (N_14855,N_14791,N_14615);
or U14856 (N_14856,N_14689,N_14627);
nor U14857 (N_14857,N_14705,N_14600);
nand U14858 (N_14858,N_14682,N_14733);
nor U14859 (N_14859,N_14717,N_14742);
and U14860 (N_14860,N_14606,N_14731);
and U14861 (N_14861,N_14780,N_14696);
xor U14862 (N_14862,N_14683,N_14709);
nand U14863 (N_14863,N_14724,N_14619);
and U14864 (N_14864,N_14662,N_14685);
nor U14865 (N_14865,N_14706,N_14718);
nand U14866 (N_14866,N_14653,N_14787);
nand U14867 (N_14867,N_14788,N_14795);
nor U14868 (N_14868,N_14644,N_14778);
and U14869 (N_14869,N_14663,N_14702);
and U14870 (N_14870,N_14658,N_14769);
nor U14871 (N_14871,N_14789,N_14630);
and U14872 (N_14872,N_14628,N_14704);
nand U14873 (N_14873,N_14792,N_14643);
or U14874 (N_14874,N_14655,N_14618);
nor U14875 (N_14875,N_14713,N_14753);
nor U14876 (N_14876,N_14692,N_14634);
nand U14877 (N_14877,N_14722,N_14635);
nor U14878 (N_14878,N_14734,N_14759);
nand U14879 (N_14879,N_14751,N_14676);
nand U14880 (N_14880,N_14774,N_14656);
and U14881 (N_14881,N_14797,N_14755);
or U14882 (N_14882,N_14764,N_14783);
nand U14883 (N_14883,N_14647,N_14727);
or U14884 (N_14884,N_14601,N_14798);
nor U14885 (N_14885,N_14762,N_14620);
and U14886 (N_14886,N_14604,N_14661);
nor U14887 (N_14887,N_14675,N_14614);
nand U14888 (N_14888,N_14784,N_14667);
nor U14889 (N_14889,N_14746,N_14776);
nor U14890 (N_14890,N_14680,N_14723);
and U14891 (N_14891,N_14761,N_14672);
nor U14892 (N_14892,N_14639,N_14677);
or U14893 (N_14893,N_14638,N_14613);
or U14894 (N_14894,N_14623,N_14793);
and U14895 (N_14895,N_14767,N_14714);
and U14896 (N_14896,N_14674,N_14609);
nand U14897 (N_14897,N_14633,N_14749);
or U14898 (N_14898,N_14785,N_14796);
nand U14899 (N_14899,N_14771,N_14608);
nor U14900 (N_14900,N_14643,N_14687);
nor U14901 (N_14901,N_14714,N_14644);
nand U14902 (N_14902,N_14745,N_14640);
and U14903 (N_14903,N_14611,N_14731);
or U14904 (N_14904,N_14729,N_14749);
and U14905 (N_14905,N_14626,N_14752);
nor U14906 (N_14906,N_14677,N_14664);
and U14907 (N_14907,N_14796,N_14652);
nor U14908 (N_14908,N_14630,N_14723);
or U14909 (N_14909,N_14679,N_14623);
or U14910 (N_14910,N_14727,N_14612);
nand U14911 (N_14911,N_14615,N_14703);
nor U14912 (N_14912,N_14715,N_14669);
nor U14913 (N_14913,N_14697,N_14715);
nor U14914 (N_14914,N_14743,N_14683);
nor U14915 (N_14915,N_14733,N_14722);
xnor U14916 (N_14916,N_14795,N_14757);
nand U14917 (N_14917,N_14795,N_14717);
or U14918 (N_14918,N_14761,N_14781);
nor U14919 (N_14919,N_14615,N_14731);
or U14920 (N_14920,N_14632,N_14652);
nand U14921 (N_14921,N_14651,N_14783);
nand U14922 (N_14922,N_14754,N_14616);
nor U14923 (N_14923,N_14778,N_14767);
nand U14924 (N_14924,N_14711,N_14606);
or U14925 (N_14925,N_14630,N_14650);
nor U14926 (N_14926,N_14701,N_14665);
nor U14927 (N_14927,N_14667,N_14666);
and U14928 (N_14928,N_14705,N_14761);
nor U14929 (N_14929,N_14749,N_14745);
and U14930 (N_14930,N_14796,N_14792);
nand U14931 (N_14931,N_14608,N_14741);
and U14932 (N_14932,N_14679,N_14724);
or U14933 (N_14933,N_14798,N_14603);
and U14934 (N_14934,N_14748,N_14706);
or U14935 (N_14935,N_14634,N_14795);
and U14936 (N_14936,N_14608,N_14654);
nand U14937 (N_14937,N_14784,N_14756);
nor U14938 (N_14938,N_14603,N_14705);
nor U14939 (N_14939,N_14746,N_14773);
nor U14940 (N_14940,N_14794,N_14614);
or U14941 (N_14941,N_14756,N_14655);
and U14942 (N_14942,N_14640,N_14659);
and U14943 (N_14943,N_14626,N_14791);
and U14944 (N_14944,N_14687,N_14777);
nand U14945 (N_14945,N_14758,N_14757);
nand U14946 (N_14946,N_14738,N_14783);
or U14947 (N_14947,N_14718,N_14684);
nand U14948 (N_14948,N_14707,N_14634);
or U14949 (N_14949,N_14703,N_14769);
or U14950 (N_14950,N_14779,N_14757);
or U14951 (N_14951,N_14791,N_14794);
and U14952 (N_14952,N_14730,N_14630);
or U14953 (N_14953,N_14617,N_14666);
nor U14954 (N_14954,N_14710,N_14667);
and U14955 (N_14955,N_14717,N_14671);
nor U14956 (N_14956,N_14679,N_14755);
nand U14957 (N_14957,N_14614,N_14658);
nand U14958 (N_14958,N_14782,N_14731);
or U14959 (N_14959,N_14703,N_14777);
or U14960 (N_14960,N_14647,N_14629);
and U14961 (N_14961,N_14653,N_14732);
nand U14962 (N_14962,N_14671,N_14672);
and U14963 (N_14963,N_14630,N_14679);
nand U14964 (N_14964,N_14619,N_14650);
nor U14965 (N_14965,N_14770,N_14790);
and U14966 (N_14966,N_14678,N_14681);
nor U14967 (N_14967,N_14610,N_14705);
or U14968 (N_14968,N_14763,N_14776);
and U14969 (N_14969,N_14747,N_14782);
or U14970 (N_14970,N_14684,N_14722);
or U14971 (N_14971,N_14628,N_14681);
or U14972 (N_14972,N_14785,N_14688);
nor U14973 (N_14973,N_14638,N_14738);
nand U14974 (N_14974,N_14673,N_14683);
and U14975 (N_14975,N_14699,N_14678);
nand U14976 (N_14976,N_14747,N_14719);
nand U14977 (N_14977,N_14678,N_14644);
or U14978 (N_14978,N_14769,N_14750);
nand U14979 (N_14979,N_14740,N_14606);
nor U14980 (N_14980,N_14673,N_14710);
or U14981 (N_14981,N_14662,N_14630);
or U14982 (N_14982,N_14650,N_14693);
and U14983 (N_14983,N_14794,N_14700);
nor U14984 (N_14984,N_14692,N_14624);
nand U14985 (N_14985,N_14652,N_14711);
and U14986 (N_14986,N_14646,N_14742);
and U14987 (N_14987,N_14728,N_14691);
nor U14988 (N_14988,N_14702,N_14724);
or U14989 (N_14989,N_14664,N_14789);
nand U14990 (N_14990,N_14738,N_14604);
or U14991 (N_14991,N_14791,N_14705);
nand U14992 (N_14992,N_14606,N_14600);
nor U14993 (N_14993,N_14631,N_14770);
nor U14994 (N_14994,N_14644,N_14696);
and U14995 (N_14995,N_14789,N_14705);
or U14996 (N_14996,N_14600,N_14652);
or U14997 (N_14997,N_14733,N_14744);
or U14998 (N_14998,N_14756,N_14654);
nand U14999 (N_14999,N_14637,N_14659);
and U15000 (N_15000,N_14973,N_14848);
nor U15001 (N_15001,N_14831,N_14857);
nand U15002 (N_15002,N_14821,N_14808);
and U15003 (N_15003,N_14960,N_14981);
and U15004 (N_15004,N_14803,N_14852);
or U15005 (N_15005,N_14925,N_14820);
or U15006 (N_15006,N_14870,N_14955);
nor U15007 (N_15007,N_14875,N_14986);
nor U15008 (N_15008,N_14942,N_14900);
or U15009 (N_15009,N_14901,N_14853);
and U15010 (N_15010,N_14836,N_14982);
nor U15011 (N_15011,N_14984,N_14879);
or U15012 (N_15012,N_14936,N_14980);
or U15013 (N_15013,N_14866,N_14861);
or U15014 (N_15014,N_14834,N_14975);
nand U15015 (N_15015,N_14921,N_14881);
nand U15016 (N_15016,N_14903,N_14926);
or U15017 (N_15017,N_14871,N_14816);
and U15018 (N_15018,N_14924,N_14950);
and U15019 (N_15019,N_14892,N_14806);
nor U15020 (N_15020,N_14801,N_14948);
nor U15021 (N_15021,N_14867,N_14844);
and U15022 (N_15022,N_14911,N_14949);
nand U15023 (N_15023,N_14920,N_14931);
nor U15024 (N_15024,N_14883,N_14922);
nor U15025 (N_15025,N_14897,N_14945);
or U15026 (N_15026,N_14964,N_14958);
nand U15027 (N_15027,N_14993,N_14966);
nor U15028 (N_15028,N_14997,N_14858);
nand U15029 (N_15029,N_14890,N_14990);
nand U15030 (N_15030,N_14915,N_14873);
nand U15031 (N_15031,N_14855,N_14988);
or U15032 (N_15032,N_14951,N_14956);
nor U15033 (N_15033,N_14987,N_14826);
or U15034 (N_15034,N_14907,N_14946);
nor U15035 (N_15035,N_14817,N_14952);
or U15036 (N_15036,N_14869,N_14914);
nand U15037 (N_15037,N_14818,N_14823);
and U15038 (N_15038,N_14862,N_14916);
nor U15039 (N_15039,N_14887,N_14977);
nor U15040 (N_15040,N_14909,N_14846);
and U15041 (N_15041,N_14838,N_14830);
or U15042 (N_15042,N_14904,N_14800);
and U15043 (N_15043,N_14943,N_14910);
and U15044 (N_15044,N_14891,N_14804);
or U15045 (N_15045,N_14954,N_14983);
or U15046 (N_15046,N_14832,N_14840);
nor U15047 (N_15047,N_14835,N_14992);
nand U15048 (N_15048,N_14811,N_14906);
and U15049 (N_15049,N_14935,N_14849);
nand U15050 (N_15050,N_14930,N_14968);
and U15051 (N_15051,N_14919,N_14839);
nor U15052 (N_15052,N_14829,N_14885);
or U15053 (N_15053,N_14888,N_14863);
nor U15054 (N_15054,N_14991,N_14902);
xor U15055 (N_15055,N_14971,N_14933);
nor U15056 (N_15056,N_14841,N_14884);
nand U15057 (N_15057,N_14802,N_14938);
nand U15058 (N_15058,N_14939,N_14843);
nand U15059 (N_15059,N_14947,N_14989);
nand U15060 (N_15060,N_14918,N_14896);
nor U15061 (N_15061,N_14828,N_14882);
nor U15062 (N_15062,N_14995,N_14932);
nand U15063 (N_15063,N_14974,N_14959);
nand U15064 (N_15064,N_14827,N_14874);
and U15065 (N_15065,N_14994,N_14822);
nand U15066 (N_15066,N_14967,N_14850);
or U15067 (N_15067,N_14912,N_14998);
or U15068 (N_15068,N_14880,N_14917);
nor U15069 (N_15069,N_14859,N_14985);
and U15070 (N_15070,N_14941,N_14860);
and U15071 (N_15071,N_14889,N_14978);
and U15072 (N_15072,N_14813,N_14928);
and U15073 (N_15073,N_14805,N_14847);
nor U15074 (N_15074,N_14824,N_14953);
nor U15075 (N_15075,N_14877,N_14996);
and U15076 (N_15076,N_14999,N_14837);
nand U15077 (N_15077,N_14957,N_14940);
nor U15078 (N_15078,N_14970,N_14961);
nand U15079 (N_15079,N_14965,N_14865);
or U15080 (N_15080,N_14898,N_14845);
or U15081 (N_15081,N_14937,N_14908);
nor U15082 (N_15082,N_14929,N_14872);
nand U15083 (N_15083,N_14962,N_14923);
or U15084 (N_15084,N_14812,N_14876);
nor U15085 (N_15085,N_14833,N_14905);
nor U15086 (N_15086,N_14969,N_14894);
or U15087 (N_15087,N_14810,N_14934);
nor U15088 (N_15088,N_14878,N_14819);
and U15089 (N_15089,N_14864,N_14893);
nand U15090 (N_15090,N_14979,N_14814);
and U15091 (N_15091,N_14842,N_14886);
and U15092 (N_15092,N_14815,N_14809);
or U15093 (N_15093,N_14972,N_14976);
nor U15094 (N_15094,N_14856,N_14895);
and U15095 (N_15095,N_14807,N_14854);
or U15096 (N_15096,N_14825,N_14899);
and U15097 (N_15097,N_14868,N_14944);
or U15098 (N_15098,N_14927,N_14963);
and U15099 (N_15099,N_14851,N_14913);
or U15100 (N_15100,N_14971,N_14883);
nand U15101 (N_15101,N_14955,N_14810);
nand U15102 (N_15102,N_14815,N_14849);
nor U15103 (N_15103,N_14874,N_14800);
nand U15104 (N_15104,N_14823,N_14905);
nand U15105 (N_15105,N_14826,N_14833);
nand U15106 (N_15106,N_14830,N_14869);
nor U15107 (N_15107,N_14893,N_14967);
nand U15108 (N_15108,N_14970,N_14855);
nand U15109 (N_15109,N_14871,N_14827);
or U15110 (N_15110,N_14800,N_14959);
nand U15111 (N_15111,N_14924,N_14874);
and U15112 (N_15112,N_14860,N_14992);
or U15113 (N_15113,N_14875,N_14856);
nand U15114 (N_15114,N_14831,N_14980);
and U15115 (N_15115,N_14932,N_14852);
and U15116 (N_15116,N_14853,N_14861);
and U15117 (N_15117,N_14932,N_14845);
or U15118 (N_15118,N_14876,N_14863);
and U15119 (N_15119,N_14965,N_14871);
nor U15120 (N_15120,N_14941,N_14982);
nor U15121 (N_15121,N_14817,N_14953);
and U15122 (N_15122,N_14982,N_14915);
nor U15123 (N_15123,N_14912,N_14811);
xor U15124 (N_15124,N_14816,N_14951);
nor U15125 (N_15125,N_14993,N_14990);
nor U15126 (N_15126,N_14981,N_14836);
nand U15127 (N_15127,N_14888,N_14938);
or U15128 (N_15128,N_14897,N_14904);
nand U15129 (N_15129,N_14971,N_14921);
nand U15130 (N_15130,N_14832,N_14955);
nand U15131 (N_15131,N_14974,N_14988);
and U15132 (N_15132,N_14861,N_14850);
or U15133 (N_15133,N_14883,N_14830);
nor U15134 (N_15134,N_14879,N_14885);
nand U15135 (N_15135,N_14995,N_14842);
nor U15136 (N_15136,N_14940,N_14814);
or U15137 (N_15137,N_14951,N_14902);
or U15138 (N_15138,N_14886,N_14873);
nand U15139 (N_15139,N_14911,N_14980);
or U15140 (N_15140,N_14826,N_14953);
nor U15141 (N_15141,N_14867,N_14942);
or U15142 (N_15142,N_14852,N_14974);
or U15143 (N_15143,N_14927,N_14989);
nor U15144 (N_15144,N_14889,N_14917);
and U15145 (N_15145,N_14920,N_14918);
nor U15146 (N_15146,N_14970,N_14892);
and U15147 (N_15147,N_14873,N_14806);
and U15148 (N_15148,N_14951,N_14963);
and U15149 (N_15149,N_14915,N_14834);
or U15150 (N_15150,N_14860,N_14853);
nor U15151 (N_15151,N_14931,N_14877);
nor U15152 (N_15152,N_14831,N_14954);
or U15153 (N_15153,N_14935,N_14938);
or U15154 (N_15154,N_14813,N_14894);
nor U15155 (N_15155,N_14916,N_14897);
nor U15156 (N_15156,N_14926,N_14931);
nand U15157 (N_15157,N_14842,N_14824);
nand U15158 (N_15158,N_14859,N_14977);
and U15159 (N_15159,N_14965,N_14824);
and U15160 (N_15160,N_14837,N_14998);
and U15161 (N_15161,N_14804,N_14905);
nand U15162 (N_15162,N_14992,N_14945);
or U15163 (N_15163,N_14907,N_14880);
or U15164 (N_15164,N_14870,N_14962);
or U15165 (N_15165,N_14978,N_14964);
and U15166 (N_15166,N_14906,N_14836);
or U15167 (N_15167,N_14921,N_14948);
and U15168 (N_15168,N_14947,N_14843);
and U15169 (N_15169,N_14934,N_14851);
nand U15170 (N_15170,N_14853,N_14982);
or U15171 (N_15171,N_14861,N_14950);
nand U15172 (N_15172,N_14956,N_14944);
nor U15173 (N_15173,N_14969,N_14895);
nor U15174 (N_15174,N_14993,N_14984);
and U15175 (N_15175,N_14943,N_14855);
and U15176 (N_15176,N_14834,N_14803);
nor U15177 (N_15177,N_14812,N_14860);
or U15178 (N_15178,N_14855,N_14981);
nand U15179 (N_15179,N_14923,N_14994);
and U15180 (N_15180,N_14980,N_14945);
or U15181 (N_15181,N_14904,N_14866);
or U15182 (N_15182,N_14971,N_14817);
nor U15183 (N_15183,N_14971,N_14898);
and U15184 (N_15184,N_14989,N_14839);
nor U15185 (N_15185,N_14825,N_14929);
and U15186 (N_15186,N_14952,N_14821);
and U15187 (N_15187,N_14935,N_14810);
and U15188 (N_15188,N_14937,N_14898);
or U15189 (N_15189,N_14953,N_14950);
or U15190 (N_15190,N_14887,N_14961);
or U15191 (N_15191,N_14951,N_14849);
nand U15192 (N_15192,N_14986,N_14941);
or U15193 (N_15193,N_14845,N_14839);
nand U15194 (N_15194,N_14914,N_14945);
nand U15195 (N_15195,N_14984,N_14976);
or U15196 (N_15196,N_14937,N_14819);
and U15197 (N_15197,N_14822,N_14970);
nand U15198 (N_15198,N_14840,N_14800);
and U15199 (N_15199,N_14834,N_14839);
and U15200 (N_15200,N_15098,N_15001);
nand U15201 (N_15201,N_15168,N_15055);
or U15202 (N_15202,N_15139,N_15145);
nand U15203 (N_15203,N_15059,N_15113);
nand U15204 (N_15204,N_15179,N_15137);
and U15205 (N_15205,N_15181,N_15142);
and U15206 (N_15206,N_15032,N_15174);
nand U15207 (N_15207,N_15189,N_15000);
and U15208 (N_15208,N_15021,N_15080);
and U15209 (N_15209,N_15015,N_15195);
and U15210 (N_15210,N_15117,N_15044);
nor U15211 (N_15211,N_15081,N_15199);
nand U15212 (N_15212,N_15029,N_15194);
nand U15213 (N_15213,N_15188,N_15116);
and U15214 (N_15214,N_15156,N_15053);
and U15215 (N_15215,N_15014,N_15121);
nand U15216 (N_15216,N_15041,N_15045);
or U15217 (N_15217,N_15006,N_15025);
or U15218 (N_15218,N_15071,N_15038);
or U15219 (N_15219,N_15146,N_15026);
and U15220 (N_15220,N_15019,N_15018);
nor U15221 (N_15221,N_15182,N_15089);
or U15222 (N_15222,N_15196,N_15102);
nor U15223 (N_15223,N_15126,N_15099);
nand U15224 (N_15224,N_15064,N_15074);
or U15225 (N_15225,N_15009,N_15150);
or U15226 (N_15226,N_15086,N_15140);
nand U15227 (N_15227,N_15036,N_15193);
nand U15228 (N_15228,N_15110,N_15151);
nand U15229 (N_15229,N_15073,N_15136);
nor U15230 (N_15230,N_15020,N_15120);
nor U15231 (N_15231,N_15052,N_15085);
nor U15232 (N_15232,N_15147,N_15197);
nor U15233 (N_15233,N_15067,N_15063);
and U15234 (N_15234,N_15131,N_15092);
nand U15235 (N_15235,N_15163,N_15164);
nor U15236 (N_15236,N_15170,N_15106);
or U15237 (N_15237,N_15198,N_15167);
and U15238 (N_15238,N_15010,N_15042);
nor U15239 (N_15239,N_15191,N_15173);
and U15240 (N_15240,N_15076,N_15165);
nand U15241 (N_15241,N_15079,N_15039);
and U15242 (N_15242,N_15175,N_15097);
nand U15243 (N_15243,N_15155,N_15100);
or U15244 (N_15244,N_15144,N_15157);
nor U15245 (N_15245,N_15070,N_15128);
nand U15246 (N_15246,N_15088,N_15103);
and U15247 (N_15247,N_15125,N_15119);
or U15248 (N_15248,N_15122,N_15104);
and U15249 (N_15249,N_15037,N_15186);
and U15250 (N_15250,N_15031,N_15172);
or U15251 (N_15251,N_15033,N_15093);
and U15252 (N_15252,N_15095,N_15034);
or U15253 (N_15253,N_15008,N_15048);
or U15254 (N_15254,N_15187,N_15012);
or U15255 (N_15255,N_15030,N_15133);
xnor U15256 (N_15256,N_15083,N_15077);
nor U15257 (N_15257,N_15138,N_15016);
nor U15258 (N_15258,N_15148,N_15149);
nand U15259 (N_15259,N_15115,N_15158);
nor U15260 (N_15260,N_15192,N_15050);
and U15261 (N_15261,N_15024,N_15075);
nand U15262 (N_15262,N_15065,N_15028);
nand U15263 (N_15263,N_15169,N_15047);
or U15264 (N_15264,N_15162,N_15027);
or U15265 (N_15265,N_15087,N_15040);
or U15266 (N_15266,N_15013,N_15177);
nand U15267 (N_15267,N_15160,N_15022);
nand U15268 (N_15268,N_15096,N_15090);
or U15269 (N_15269,N_15124,N_15078);
nor U15270 (N_15270,N_15108,N_15058);
nor U15271 (N_15271,N_15084,N_15069);
nor U15272 (N_15272,N_15176,N_15062);
and U15273 (N_15273,N_15101,N_15123);
nand U15274 (N_15274,N_15094,N_15002);
nand U15275 (N_15275,N_15109,N_15035);
or U15276 (N_15276,N_15003,N_15134);
or U15277 (N_15277,N_15056,N_15161);
nand U15278 (N_15278,N_15135,N_15007);
nor U15279 (N_15279,N_15152,N_15054);
nor U15280 (N_15280,N_15143,N_15127);
nor U15281 (N_15281,N_15111,N_15049);
or U15282 (N_15282,N_15159,N_15072);
nor U15283 (N_15283,N_15107,N_15185);
nor U15284 (N_15284,N_15105,N_15184);
or U15285 (N_15285,N_15132,N_15060);
or U15286 (N_15286,N_15153,N_15118);
or U15287 (N_15287,N_15082,N_15004);
nand U15288 (N_15288,N_15171,N_15068);
and U15289 (N_15289,N_15114,N_15011);
nor U15290 (N_15290,N_15057,N_15166);
and U15291 (N_15291,N_15154,N_15005);
and U15292 (N_15292,N_15141,N_15046);
and U15293 (N_15293,N_15023,N_15043);
nor U15294 (N_15294,N_15183,N_15130);
and U15295 (N_15295,N_15051,N_15178);
nor U15296 (N_15296,N_15061,N_15112);
and U15297 (N_15297,N_15129,N_15017);
nor U15298 (N_15298,N_15066,N_15180);
nor U15299 (N_15299,N_15091,N_15190);
nor U15300 (N_15300,N_15139,N_15055);
and U15301 (N_15301,N_15157,N_15146);
or U15302 (N_15302,N_15143,N_15128);
or U15303 (N_15303,N_15031,N_15071);
and U15304 (N_15304,N_15112,N_15116);
or U15305 (N_15305,N_15002,N_15131);
and U15306 (N_15306,N_15070,N_15087);
nor U15307 (N_15307,N_15194,N_15060);
nand U15308 (N_15308,N_15135,N_15170);
or U15309 (N_15309,N_15179,N_15087);
and U15310 (N_15310,N_15165,N_15005);
or U15311 (N_15311,N_15054,N_15137);
nor U15312 (N_15312,N_15139,N_15137);
or U15313 (N_15313,N_15197,N_15024);
or U15314 (N_15314,N_15093,N_15022);
or U15315 (N_15315,N_15074,N_15163);
and U15316 (N_15316,N_15174,N_15018);
nand U15317 (N_15317,N_15025,N_15145);
nand U15318 (N_15318,N_15074,N_15125);
or U15319 (N_15319,N_15123,N_15078);
or U15320 (N_15320,N_15040,N_15016);
or U15321 (N_15321,N_15037,N_15081);
nor U15322 (N_15322,N_15094,N_15177);
or U15323 (N_15323,N_15136,N_15151);
nor U15324 (N_15324,N_15166,N_15175);
or U15325 (N_15325,N_15116,N_15091);
and U15326 (N_15326,N_15196,N_15016);
nor U15327 (N_15327,N_15187,N_15191);
or U15328 (N_15328,N_15052,N_15121);
or U15329 (N_15329,N_15131,N_15079);
and U15330 (N_15330,N_15133,N_15028);
and U15331 (N_15331,N_15113,N_15005);
and U15332 (N_15332,N_15162,N_15130);
nor U15333 (N_15333,N_15183,N_15043);
nor U15334 (N_15334,N_15048,N_15102);
or U15335 (N_15335,N_15044,N_15124);
or U15336 (N_15336,N_15188,N_15010);
or U15337 (N_15337,N_15145,N_15140);
or U15338 (N_15338,N_15074,N_15148);
nor U15339 (N_15339,N_15025,N_15036);
nand U15340 (N_15340,N_15114,N_15174);
or U15341 (N_15341,N_15059,N_15085);
nand U15342 (N_15342,N_15094,N_15019);
nand U15343 (N_15343,N_15177,N_15014);
and U15344 (N_15344,N_15097,N_15122);
nor U15345 (N_15345,N_15002,N_15165);
or U15346 (N_15346,N_15148,N_15095);
or U15347 (N_15347,N_15088,N_15187);
nand U15348 (N_15348,N_15178,N_15099);
nor U15349 (N_15349,N_15141,N_15198);
and U15350 (N_15350,N_15067,N_15030);
and U15351 (N_15351,N_15039,N_15018);
nor U15352 (N_15352,N_15047,N_15110);
and U15353 (N_15353,N_15063,N_15189);
and U15354 (N_15354,N_15138,N_15166);
and U15355 (N_15355,N_15008,N_15112);
and U15356 (N_15356,N_15036,N_15011);
or U15357 (N_15357,N_15076,N_15058);
and U15358 (N_15358,N_15133,N_15158);
and U15359 (N_15359,N_15007,N_15056);
and U15360 (N_15360,N_15117,N_15034);
or U15361 (N_15361,N_15015,N_15119);
and U15362 (N_15362,N_15174,N_15122);
nor U15363 (N_15363,N_15104,N_15169);
nand U15364 (N_15364,N_15012,N_15086);
nand U15365 (N_15365,N_15150,N_15061);
and U15366 (N_15366,N_15029,N_15172);
or U15367 (N_15367,N_15093,N_15046);
or U15368 (N_15368,N_15040,N_15033);
nand U15369 (N_15369,N_15166,N_15128);
nand U15370 (N_15370,N_15001,N_15125);
nand U15371 (N_15371,N_15064,N_15080);
or U15372 (N_15372,N_15049,N_15179);
nor U15373 (N_15373,N_15186,N_15148);
or U15374 (N_15374,N_15060,N_15171);
nand U15375 (N_15375,N_15122,N_15092);
nand U15376 (N_15376,N_15086,N_15082);
and U15377 (N_15377,N_15006,N_15012);
nor U15378 (N_15378,N_15010,N_15011);
nand U15379 (N_15379,N_15097,N_15094);
and U15380 (N_15380,N_15191,N_15067);
nand U15381 (N_15381,N_15107,N_15050);
or U15382 (N_15382,N_15174,N_15090);
nand U15383 (N_15383,N_15195,N_15185);
xnor U15384 (N_15384,N_15111,N_15082);
nand U15385 (N_15385,N_15063,N_15196);
nor U15386 (N_15386,N_15051,N_15176);
or U15387 (N_15387,N_15059,N_15005);
or U15388 (N_15388,N_15041,N_15093);
nor U15389 (N_15389,N_15192,N_15117);
nor U15390 (N_15390,N_15156,N_15049);
and U15391 (N_15391,N_15056,N_15165);
nand U15392 (N_15392,N_15154,N_15002);
or U15393 (N_15393,N_15174,N_15146);
nor U15394 (N_15394,N_15109,N_15132);
nor U15395 (N_15395,N_15039,N_15162);
and U15396 (N_15396,N_15155,N_15172);
nor U15397 (N_15397,N_15010,N_15121);
and U15398 (N_15398,N_15167,N_15085);
and U15399 (N_15399,N_15160,N_15151);
nor U15400 (N_15400,N_15257,N_15350);
nor U15401 (N_15401,N_15327,N_15214);
or U15402 (N_15402,N_15265,N_15365);
nand U15403 (N_15403,N_15288,N_15387);
nand U15404 (N_15404,N_15245,N_15330);
and U15405 (N_15405,N_15340,N_15316);
nor U15406 (N_15406,N_15283,N_15267);
and U15407 (N_15407,N_15374,N_15255);
nand U15408 (N_15408,N_15358,N_15342);
and U15409 (N_15409,N_15355,N_15321);
nor U15410 (N_15410,N_15392,N_15324);
or U15411 (N_15411,N_15377,N_15221);
or U15412 (N_15412,N_15210,N_15395);
and U15413 (N_15413,N_15236,N_15364);
nor U15414 (N_15414,N_15369,N_15273);
or U15415 (N_15415,N_15396,N_15278);
or U15416 (N_15416,N_15213,N_15252);
nand U15417 (N_15417,N_15372,N_15271);
nand U15418 (N_15418,N_15248,N_15289);
and U15419 (N_15419,N_15348,N_15353);
and U15420 (N_15420,N_15315,N_15212);
or U15421 (N_15421,N_15231,N_15336);
and U15422 (N_15422,N_15307,N_15200);
xnor U15423 (N_15423,N_15202,N_15375);
and U15424 (N_15424,N_15370,N_15258);
and U15425 (N_15425,N_15346,N_15379);
and U15426 (N_15426,N_15295,N_15241);
and U15427 (N_15427,N_15246,N_15222);
nor U15428 (N_15428,N_15243,N_15234);
and U15429 (N_15429,N_15360,N_15367);
and U15430 (N_15430,N_15207,N_15304);
or U15431 (N_15431,N_15384,N_15239);
nand U15432 (N_15432,N_15256,N_15293);
and U15433 (N_15433,N_15357,N_15263);
nand U15434 (N_15434,N_15359,N_15254);
and U15435 (N_15435,N_15389,N_15393);
and U15436 (N_15436,N_15276,N_15313);
or U15437 (N_15437,N_15284,N_15230);
and U15438 (N_15438,N_15294,N_15331);
nand U15439 (N_15439,N_15386,N_15272);
or U15440 (N_15440,N_15204,N_15223);
and U15441 (N_15441,N_15305,N_15363);
nor U15442 (N_15442,N_15242,N_15332);
nor U15443 (N_15443,N_15390,N_15268);
nand U15444 (N_15444,N_15322,N_15297);
nand U15445 (N_15445,N_15253,N_15317);
nand U15446 (N_15446,N_15391,N_15343);
nor U15447 (N_15447,N_15206,N_15306);
nand U15448 (N_15448,N_15249,N_15280);
nor U15449 (N_15449,N_15211,N_15262);
or U15450 (N_15450,N_15356,N_15266);
nor U15451 (N_15451,N_15261,N_15250);
or U15452 (N_15452,N_15328,N_15323);
nand U15453 (N_15453,N_15296,N_15291);
or U15454 (N_15454,N_15371,N_15217);
nand U15455 (N_15455,N_15325,N_15244);
or U15456 (N_15456,N_15208,N_15385);
and U15457 (N_15457,N_15347,N_15235);
nor U15458 (N_15458,N_15300,N_15344);
nand U15459 (N_15459,N_15398,N_15399);
or U15460 (N_15460,N_15352,N_15282);
and U15461 (N_15461,N_15251,N_15368);
or U15462 (N_15462,N_15281,N_15341);
nand U15463 (N_15463,N_15270,N_15274);
and U15464 (N_15464,N_15277,N_15335);
nand U15465 (N_15465,N_15318,N_15388);
or U15466 (N_15466,N_15203,N_15329);
nand U15467 (N_15467,N_15312,N_15381);
and U15468 (N_15468,N_15351,N_15205);
or U15469 (N_15469,N_15397,N_15290);
nor U15470 (N_15470,N_15238,N_15362);
nor U15471 (N_15471,N_15361,N_15233);
nand U15472 (N_15472,N_15378,N_15366);
nor U15473 (N_15473,N_15298,N_15259);
and U15474 (N_15474,N_15286,N_15319);
and U15475 (N_15475,N_15382,N_15209);
or U15476 (N_15476,N_15320,N_15247);
nand U15477 (N_15477,N_15201,N_15394);
nand U15478 (N_15478,N_15380,N_15287);
nand U15479 (N_15479,N_15334,N_15376);
or U15480 (N_15480,N_15269,N_15232);
or U15481 (N_15481,N_15326,N_15237);
or U15482 (N_15482,N_15338,N_15339);
or U15483 (N_15483,N_15333,N_15224);
and U15484 (N_15484,N_15228,N_15383);
and U15485 (N_15485,N_15308,N_15275);
and U15486 (N_15486,N_15279,N_15219);
and U15487 (N_15487,N_15299,N_15220);
and U15488 (N_15488,N_15226,N_15225);
nor U15489 (N_15489,N_15354,N_15240);
or U15490 (N_15490,N_15227,N_15216);
nor U15491 (N_15491,N_15373,N_15311);
and U15492 (N_15492,N_15314,N_15229);
or U15493 (N_15493,N_15264,N_15285);
nor U15494 (N_15494,N_15349,N_15309);
nor U15495 (N_15495,N_15302,N_15218);
or U15496 (N_15496,N_15310,N_15292);
or U15497 (N_15497,N_15337,N_15260);
nand U15498 (N_15498,N_15301,N_15303);
nor U15499 (N_15499,N_15215,N_15345);
nand U15500 (N_15500,N_15233,N_15283);
nor U15501 (N_15501,N_15281,N_15301);
nor U15502 (N_15502,N_15291,N_15381);
nand U15503 (N_15503,N_15381,N_15345);
nand U15504 (N_15504,N_15243,N_15324);
nor U15505 (N_15505,N_15254,N_15396);
and U15506 (N_15506,N_15243,N_15383);
and U15507 (N_15507,N_15359,N_15211);
or U15508 (N_15508,N_15222,N_15226);
and U15509 (N_15509,N_15370,N_15381);
and U15510 (N_15510,N_15324,N_15317);
nor U15511 (N_15511,N_15391,N_15296);
nand U15512 (N_15512,N_15381,N_15327);
and U15513 (N_15513,N_15223,N_15290);
or U15514 (N_15514,N_15364,N_15326);
nand U15515 (N_15515,N_15356,N_15384);
nand U15516 (N_15516,N_15264,N_15370);
nand U15517 (N_15517,N_15376,N_15295);
and U15518 (N_15518,N_15237,N_15271);
nor U15519 (N_15519,N_15211,N_15363);
nand U15520 (N_15520,N_15280,N_15399);
or U15521 (N_15521,N_15369,N_15328);
nand U15522 (N_15522,N_15273,N_15346);
nand U15523 (N_15523,N_15309,N_15271);
and U15524 (N_15524,N_15336,N_15232);
and U15525 (N_15525,N_15384,N_15323);
and U15526 (N_15526,N_15222,N_15383);
nor U15527 (N_15527,N_15216,N_15296);
nor U15528 (N_15528,N_15394,N_15223);
or U15529 (N_15529,N_15305,N_15309);
and U15530 (N_15530,N_15359,N_15247);
nor U15531 (N_15531,N_15390,N_15373);
nand U15532 (N_15532,N_15222,N_15272);
or U15533 (N_15533,N_15200,N_15238);
nor U15534 (N_15534,N_15286,N_15375);
and U15535 (N_15535,N_15217,N_15305);
nand U15536 (N_15536,N_15217,N_15386);
and U15537 (N_15537,N_15209,N_15331);
nor U15538 (N_15538,N_15392,N_15234);
and U15539 (N_15539,N_15393,N_15351);
nor U15540 (N_15540,N_15370,N_15305);
nand U15541 (N_15541,N_15287,N_15363);
and U15542 (N_15542,N_15299,N_15211);
or U15543 (N_15543,N_15236,N_15214);
or U15544 (N_15544,N_15201,N_15373);
nor U15545 (N_15545,N_15292,N_15373);
nand U15546 (N_15546,N_15312,N_15327);
nor U15547 (N_15547,N_15236,N_15295);
nor U15548 (N_15548,N_15377,N_15365);
and U15549 (N_15549,N_15360,N_15271);
and U15550 (N_15550,N_15357,N_15269);
nand U15551 (N_15551,N_15344,N_15369);
nor U15552 (N_15552,N_15264,N_15385);
and U15553 (N_15553,N_15219,N_15278);
or U15554 (N_15554,N_15220,N_15357);
and U15555 (N_15555,N_15226,N_15379);
nor U15556 (N_15556,N_15316,N_15374);
nand U15557 (N_15557,N_15373,N_15344);
nor U15558 (N_15558,N_15220,N_15358);
nor U15559 (N_15559,N_15303,N_15277);
nor U15560 (N_15560,N_15266,N_15287);
and U15561 (N_15561,N_15238,N_15369);
nand U15562 (N_15562,N_15307,N_15251);
or U15563 (N_15563,N_15316,N_15236);
nor U15564 (N_15564,N_15217,N_15241);
or U15565 (N_15565,N_15302,N_15279);
nand U15566 (N_15566,N_15244,N_15312);
and U15567 (N_15567,N_15208,N_15381);
and U15568 (N_15568,N_15253,N_15339);
and U15569 (N_15569,N_15357,N_15271);
and U15570 (N_15570,N_15305,N_15253);
nor U15571 (N_15571,N_15213,N_15354);
or U15572 (N_15572,N_15261,N_15219);
nor U15573 (N_15573,N_15305,N_15344);
or U15574 (N_15574,N_15299,N_15382);
nor U15575 (N_15575,N_15257,N_15388);
or U15576 (N_15576,N_15221,N_15241);
nand U15577 (N_15577,N_15361,N_15225);
nor U15578 (N_15578,N_15322,N_15254);
nand U15579 (N_15579,N_15257,N_15226);
nand U15580 (N_15580,N_15346,N_15329);
nor U15581 (N_15581,N_15327,N_15237);
nor U15582 (N_15582,N_15382,N_15387);
and U15583 (N_15583,N_15289,N_15268);
or U15584 (N_15584,N_15237,N_15290);
nand U15585 (N_15585,N_15285,N_15395);
or U15586 (N_15586,N_15350,N_15331);
nor U15587 (N_15587,N_15344,N_15257);
and U15588 (N_15588,N_15302,N_15239);
or U15589 (N_15589,N_15272,N_15311);
nor U15590 (N_15590,N_15251,N_15350);
nand U15591 (N_15591,N_15333,N_15200);
nor U15592 (N_15592,N_15361,N_15323);
and U15593 (N_15593,N_15362,N_15317);
nand U15594 (N_15594,N_15205,N_15302);
or U15595 (N_15595,N_15269,N_15385);
and U15596 (N_15596,N_15286,N_15377);
nor U15597 (N_15597,N_15311,N_15337);
nor U15598 (N_15598,N_15280,N_15243);
nand U15599 (N_15599,N_15279,N_15378);
nor U15600 (N_15600,N_15584,N_15429);
and U15601 (N_15601,N_15589,N_15598);
or U15602 (N_15602,N_15431,N_15573);
or U15603 (N_15603,N_15511,N_15553);
nor U15604 (N_15604,N_15585,N_15457);
or U15605 (N_15605,N_15599,N_15416);
and U15606 (N_15606,N_15540,N_15592);
and U15607 (N_15607,N_15593,N_15562);
nor U15608 (N_15608,N_15575,N_15543);
nand U15609 (N_15609,N_15474,N_15558);
and U15610 (N_15610,N_15446,N_15514);
and U15611 (N_15611,N_15521,N_15458);
nor U15612 (N_15612,N_15560,N_15591);
nor U15613 (N_15613,N_15570,N_15522);
nand U15614 (N_15614,N_15550,N_15491);
nor U15615 (N_15615,N_15421,N_15410);
and U15616 (N_15616,N_15500,N_15468);
or U15617 (N_15617,N_15564,N_15432);
nor U15618 (N_15618,N_15559,N_15417);
nand U15619 (N_15619,N_15469,N_15556);
nor U15620 (N_15620,N_15477,N_15502);
or U15621 (N_15621,N_15567,N_15404);
nand U15622 (N_15622,N_15463,N_15533);
nand U15623 (N_15623,N_15546,N_15479);
or U15624 (N_15624,N_15439,N_15569);
or U15625 (N_15625,N_15442,N_15541);
nor U15626 (N_15626,N_15434,N_15534);
nand U15627 (N_15627,N_15586,N_15552);
and U15628 (N_15628,N_15551,N_15563);
nand U15629 (N_15629,N_15437,N_15490);
nor U15630 (N_15630,N_15454,N_15496);
nor U15631 (N_15631,N_15588,N_15480);
nand U15632 (N_15632,N_15430,N_15509);
or U15633 (N_15633,N_15529,N_15595);
or U15634 (N_15634,N_15400,N_15535);
and U15635 (N_15635,N_15467,N_15579);
or U15636 (N_15636,N_15425,N_15508);
and U15637 (N_15637,N_15524,N_15472);
nor U15638 (N_15638,N_15532,N_15489);
or U15639 (N_15639,N_15494,N_15470);
nor U15640 (N_15640,N_15497,N_15428);
nand U15641 (N_15641,N_15418,N_15495);
nand U15642 (N_15642,N_15414,N_15413);
nor U15643 (N_15643,N_15440,N_15531);
nand U15644 (N_15644,N_15572,N_15459);
nand U15645 (N_15645,N_15561,N_15460);
nor U15646 (N_15646,N_15527,N_15433);
and U15647 (N_15647,N_15536,N_15487);
nor U15648 (N_15648,N_15453,N_15465);
nor U15649 (N_15649,N_15456,N_15568);
nor U15650 (N_15650,N_15517,N_15501);
nand U15651 (N_15651,N_15574,N_15498);
nand U15652 (N_15652,N_15451,N_15438);
or U15653 (N_15653,N_15525,N_15450);
nor U15654 (N_15654,N_15578,N_15499);
and U15655 (N_15655,N_15484,N_15476);
nor U15656 (N_15656,N_15462,N_15577);
nand U15657 (N_15657,N_15554,N_15581);
nor U15658 (N_15658,N_15455,N_15580);
nand U15659 (N_15659,N_15408,N_15587);
or U15660 (N_15660,N_15405,N_15449);
nand U15661 (N_15661,N_15447,N_15471);
or U15662 (N_15662,N_15519,N_15583);
or U15663 (N_15663,N_15526,N_15473);
or U15664 (N_15664,N_15566,N_15545);
or U15665 (N_15665,N_15466,N_15448);
nand U15666 (N_15666,N_15597,N_15503);
and U15667 (N_15667,N_15548,N_15401);
xnor U15668 (N_15668,N_15486,N_15590);
nor U15669 (N_15669,N_15409,N_15542);
nand U15670 (N_15670,N_15594,N_15424);
and U15671 (N_15671,N_15420,N_15537);
nand U15672 (N_15672,N_15407,N_15411);
nor U15673 (N_15673,N_15523,N_15403);
nor U15674 (N_15674,N_15571,N_15530);
or U15675 (N_15675,N_15427,N_15565);
or U15676 (N_15676,N_15544,N_15485);
nor U15677 (N_15677,N_15419,N_15436);
or U15678 (N_15678,N_15493,N_15475);
nand U15679 (N_15679,N_15481,N_15512);
nand U15680 (N_15680,N_15444,N_15505);
nand U15681 (N_15681,N_15528,N_15520);
nand U15682 (N_15682,N_15549,N_15426);
or U15683 (N_15683,N_15582,N_15596);
or U15684 (N_15684,N_15516,N_15507);
nand U15685 (N_15685,N_15482,N_15506);
nand U15686 (N_15686,N_15412,N_15515);
nor U15687 (N_15687,N_15461,N_15435);
nor U15688 (N_15688,N_15518,N_15538);
or U15689 (N_15689,N_15539,N_15478);
and U15690 (N_15690,N_15406,N_15422);
or U15691 (N_15691,N_15483,N_15423);
and U15692 (N_15692,N_15576,N_15488);
nor U15693 (N_15693,N_15510,N_15402);
and U15694 (N_15694,N_15513,N_15443);
or U15695 (N_15695,N_15415,N_15547);
or U15696 (N_15696,N_15555,N_15504);
nor U15697 (N_15697,N_15452,N_15492);
or U15698 (N_15698,N_15464,N_15445);
xor U15699 (N_15699,N_15557,N_15441);
or U15700 (N_15700,N_15521,N_15477);
or U15701 (N_15701,N_15422,N_15419);
nor U15702 (N_15702,N_15415,N_15516);
nand U15703 (N_15703,N_15437,N_15410);
or U15704 (N_15704,N_15447,N_15503);
nor U15705 (N_15705,N_15408,N_15584);
and U15706 (N_15706,N_15512,N_15501);
or U15707 (N_15707,N_15446,N_15402);
or U15708 (N_15708,N_15593,N_15523);
or U15709 (N_15709,N_15592,N_15496);
or U15710 (N_15710,N_15526,N_15490);
nor U15711 (N_15711,N_15484,N_15415);
or U15712 (N_15712,N_15520,N_15553);
and U15713 (N_15713,N_15443,N_15527);
and U15714 (N_15714,N_15515,N_15491);
and U15715 (N_15715,N_15422,N_15403);
nor U15716 (N_15716,N_15402,N_15454);
and U15717 (N_15717,N_15494,N_15563);
and U15718 (N_15718,N_15590,N_15464);
or U15719 (N_15719,N_15487,N_15432);
and U15720 (N_15720,N_15453,N_15427);
nand U15721 (N_15721,N_15404,N_15479);
and U15722 (N_15722,N_15449,N_15427);
and U15723 (N_15723,N_15511,N_15515);
and U15724 (N_15724,N_15493,N_15593);
nand U15725 (N_15725,N_15543,N_15547);
and U15726 (N_15726,N_15586,N_15428);
nand U15727 (N_15727,N_15541,N_15595);
and U15728 (N_15728,N_15508,N_15543);
nand U15729 (N_15729,N_15417,N_15534);
or U15730 (N_15730,N_15485,N_15597);
nor U15731 (N_15731,N_15455,N_15562);
nand U15732 (N_15732,N_15491,N_15414);
nor U15733 (N_15733,N_15557,N_15577);
nand U15734 (N_15734,N_15430,N_15429);
or U15735 (N_15735,N_15559,N_15526);
and U15736 (N_15736,N_15573,N_15503);
nand U15737 (N_15737,N_15424,N_15443);
or U15738 (N_15738,N_15557,N_15560);
nand U15739 (N_15739,N_15471,N_15460);
nor U15740 (N_15740,N_15486,N_15569);
and U15741 (N_15741,N_15597,N_15417);
and U15742 (N_15742,N_15429,N_15443);
nor U15743 (N_15743,N_15424,N_15567);
nand U15744 (N_15744,N_15567,N_15458);
nor U15745 (N_15745,N_15411,N_15527);
nand U15746 (N_15746,N_15571,N_15484);
nor U15747 (N_15747,N_15524,N_15437);
and U15748 (N_15748,N_15518,N_15521);
or U15749 (N_15749,N_15458,N_15529);
and U15750 (N_15750,N_15544,N_15433);
nand U15751 (N_15751,N_15571,N_15592);
or U15752 (N_15752,N_15433,N_15565);
nor U15753 (N_15753,N_15446,N_15470);
or U15754 (N_15754,N_15434,N_15504);
or U15755 (N_15755,N_15475,N_15497);
nor U15756 (N_15756,N_15476,N_15482);
nand U15757 (N_15757,N_15519,N_15595);
and U15758 (N_15758,N_15581,N_15536);
nand U15759 (N_15759,N_15455,N_15528);
and U15760 (N_15760,N_15565,N_15423);
nor U15761 (N_15761,N_15589,N_15414);
nand U15762 (N_15762,N_15469,N_15417);
nand U15763 (N_15763,N_15469,N_15431);
nand U15764 (N_15764,N_15474,N_15410);
nor U15765 (N_15765,N_15406,N_15466);
nand U15766 (N_15766,N_15561,N_15401);
nand U15767 (N_15767,N_15586,N_15529);
or U15768 (N_15768,N_15438,N_15498);
xnor U15769 (N_15769,N_15563,N_15584);
or U15770 (N_15770,N_15530,N_15506);
and U15771 (N_15771,N_15535,N_15466);
nor U15772 (N_15772,N_15534,N_15531);
and U15773 (N_15773,N_15462,N_15599);
nor U15774 (N_15774,N_15575,N_15591);
and U15775 (N_15775,N_15535,N_15458);
nand U15776 (N_15776,N_15426,N_15569);
nor U15777 (N_15777,N_15497,N_15531);
nand U15778 (N_15778,N_15507,N_15580);
or U15779 (N_15779,N_15426,N_15506);
or U15780 (N_15780,N_15481,N_15453);
and U15781 (N_15781,N_15508,N_15537);
nand U15782 (N_15782,N_15516,N_15552);
nor U15783 (N_15783,N_15557,N_15583);
and U15784 (N_15784,N_15580,N_15470);
xnor U15785 (N_15785,N_15596,N_15493);
nand U15786 (N_15786,N_15424,N_15421);
and U15787 (N_15787,N_15502,N_15484);
and U15788 (N_15788,N_15504,N_15418);
nor U15789 (N_15789,N_15426,N_15432);
and U15790 (N_15790,N_15590,N_15472);
nor U15791 (N_15791,N_15490,N_15436);
or U15792 (N_15792,N_15500,N_15537);
and U15793 (N_15793,N_15523,N_15487);
nor U15794 (N_15794,N_15517,N_15580);
or U15795 (N_15795,N_15524,N_15525);
nand U15796 (N_15796,N_15577,N_15555);
nor U15797 (N_15797,N_15589,N_15517);
and U15798 (N_15798,N_15444,N_15488);
and U15799 (N_15799,N_15519,N_15407);
and U15800 (N_15800,N_15614,N_15796);
nor U15801 (N_15801,N_15666,N_15779);
nand U15802 (N_15802,N_15706,N_15687);
nand U15803 (N_15803,N_15615,N_15729);
or U15804 (N_15804,N_15612,N_15608);
and U15805 (N_15805,N_15644,N_15625);
or U15806 (N_15806,N_15785,N_15777);
nor U15807 (N_15807,N_15726,N_15663);
and U15808 (N_15808,N_15699,N_15693);
nand U15809 (N_15809,N_15603,N_15708);
or U15810 (N_15810,N_15767,N_15634);
and U15811 (N_15811,N_15776,N_15607);
and U15812 (N_15812,N_15722,N_15732);
nor U15813 (N_15813,N_15733,N_15639);
and U15814 (N_15814,N_15703,N_15789);
or U15815 (N_15815,N_15642,N_15690);
or U15816 (N_15816,N_15788,N_15773);
nand U15817 (N_15817,N_15745,N_15684);
and U15818 (N_15818,N_15743,N_15637);
or U15819 (N_15819,N_15761,N_15650);
nor U15820 (N_15820,N_15681,N_15668);
nor U15821 (N_15821,N_15772,N_15600);
or U15822 (N_15822,N_15627,N_15655);
nor U15823 (N_15823,N_15756,N_15778);
nand U15824 (N_15824,N_15766,N_15604);
and U15825 (N_15825,N_15737,N_15638);
nor U15826 (N_15826,N_15654,N_15782);
or U15827 (N_15827,N_15674,N_15609);
or U15828 (N_15828,N_15771,N_15658);
or U15829 (N_15829,N_15629,N_15691);
or U15830 (N_15830,N_15799,N_15667);
and U15831 (N_15831,N_15657,N_15618);
and U15832 (N_15832,N_15739,N_15797);
nor U15833 (N_15833,N_15680,N_15685);
nand U15834 (N_15834,N_15721,N_15744);
xnor U15835 (N_15835,N_15723,N_15704);
and U15836 (N_15836,N_15780,N_15675);
nand U15837 (N_15837,N_15720,N_15613);
or U15838 (N_15838,N_15677,N_15665);
or U15839 (N_15839,N_15794,N_15734);
nand U15840 (N_15840,N_15716,N_15664);
nand U15841 (N_15841,N_15707,N_15755);
or U15842 (N_15842,N_15727,N_15646);
nor U15843 (N_15843,N_15701,N_15740);
nand U15844 (N_15844,N_15623,N_15730);
nand U15845 (N_15845,N_15750,N_15783);
or U15846 (N_15846,N_15651,N_15662);
nand U15847 (N_15847,N_15754,N_15728);
and U15848 (N_15848,N_15659,N_15624);
nor U15849 (N_15849,N_15645,N_15770);
xnor U15850 (N_15850,N_15610,N_15621);
nor U15851 (N_15851,N_15712,N_15619);
and U15852 (N_15852,N_15786,N_15736);
or U15853 (N_15853,N_15696,N_15747);
or U15854 (N_15854,N_15633,N_15764);
nor U15855 (N_15855,N_15602,N_15628);
nor U15856 (N_15856,N_15686,N_15688);
nor U15857 (N_15857,N_15702,N_15648);
nor U15858 (N_15858,N_15763,N_15749);
or U15859 (N_15859,N_15714,N_15606);
or U15860 (N_15860,N_15705,N_15724);
nand U15861 (N_15861,N_15735,N_15787);
or U15862 (N_15862,N_15718,N_15698);
nand U15863 (N_15863,N_15746,N_15713);
nor U15864 (N_15864,N_15611,N_15679);
nand U15865 (N_15865,N_15795,N_15669);
or U15866 (N_15866,N_15660,N_15768);
or U15867 (N_15867,N_15620,N_15601);
nor U15868 (N_15868,N_15700,N_15626);
and U15869 (N_15869,N_15678,N_15791);
and U15870 (N_15870,N_15682,N_15635);
nand U15871 (N_15871,N_15617,N_15774);
nor U15872 (N_15872,N_15653,N_15741);
nor U15873 (N_15873,N_15683,N_15762);
and U15874 (N_15874,N_15798,N_15643);
nand U15875 (N_15875,N_15652,N_15697);
nor U15876 (N_15876,N_15640,N_15759);
and U15877 (N_15877,N_15715,N_15753);
nor U15878 (N_15878,N_15631,N_15751);
nor U15879 (N_15879,N_15710,N_15632);
nor U15880 (N_15880,N_15622,N_15738);
nor U15881 (N_15881,N_15742,N_15673);
or U15882 (N_15882,N_15692,N_15752);
and U15883 (N_15883,N_15731,N_15641);
and U15884 (N_15884,N_15790,N_15636);
nor U15885 (N_15885,N_15616,N_15630);
and U15886 (N_15886,N_15765,N_15649);
xor U15887 (N_15887,N_15672,N_15792);
and U15888 (N_15888,N_15689,N_15748);
nor U15889 (N_15889,N_15670,N_15757);
nand U15890 (N_15890,N_15676,N_15719);
nor U15891 (N_15891,N_15725,N_15711);
nand U15892 (N_15892,N_15793,N_15656);
nor U15893 (N_15893,N_15717,N_15784);
nor U15894 (N_15894,N_15769,N_15695);
nand U15895 (N_15895,N_15671,N_15647);
nand U15896 (N_15896,N_15781,N_15661);
and U15897 (N_15897,N_15605,N_15758);
or U15898 (N_15898,N_15775,N_15709);
or U15899 (N_15899,N_15760,N_15694);
nand U15900 (N_15900,N_15690,N_15669);
or U15901 (N_15901,N_15633,N_15740);
or U15902 (N_15902,N_15700,N_15686);
and U15903 (N_15903,N_15672,N_15725);
nand U15904 (N_15904,N_15706,N_15704);
or U15905 (N_15905,N_15687,N_15686);
or U15906 (N_15906,N_15757,N_15777);
nand U15907 (N_15907,N_15672,N_15728);
nand U15908 (N_15908,N_15778,N_15799);
and U15909 (N_15909,N_15797,N_15635);
or U15910 (N_15910,N_15698,N_15627);
or U15911 (N_15911,N_15746,N_15654);
nand U15912 (N_15912,N_15643,N_15745);
nand U15913 (N_15913,N_15679,N_15764);
nand U15914 (N_15914,N_15760,N_15656);
nand U15915 (N_15915,N_15646,N_15783);
and U15916 (N_15916,N_15610,N_15728);
and U15917 (N_15917,N_15760,N_15777);
nor U15918 (N_15918,N_15637,N_15673);
and U15919 (N_15919,N_15779,N_15670);
nand U15920 (N_15920,N_15743,N_15667);
nand U15921 (N_15921,N_15749,N_15638);
or U15922 (N_15922,N_15635,N_15765);
nor U15923 (N_15923,N_15791,N_15715);
and U15924 (N_15924,N_15737,N_15654);
nand U15925 (N_15925,N_15662,N_15648);
nand U15926 (N_15926,N_15623,N_15678);
or U15927 (N_15927,N_15638,N_15732);
or U15928 (N_15928,N_15721,N_15727);
nand U15929 (N_15929,N_15651,N_15635);
nor U15930 (N_15930,N_15627,N_15753);
or U15931 (N_15931,N_15649,N_15674);
and U15932 (N_15932,N_15719,N_15648);
or U15933 (N_15933,N_15700,N_15673);
nand U15934 (N_15934,N_15768,N_15741);
nand U15935 (N_15935,N_15663,N_15799);
or U15936 (N_15936,N_15720,N_15624);
nor U15937 (N_15937,N_15770,N_15668);
nor U15938 (N_15938,N_15760,N_15766);
nand U15939 (N_15939,N_15673,N_15603);
nand U15940 (N_15940,N_15739,N_15748);
or U15941 (N_15941,N_15686,N_15783);
nor U15942 (N_15942,N_15689,N_15726);
nor U15943 (N_15943,N_15679,N_15724);
and U15944 (N_15944,N_15674,N_15762);
and U15945 (N_15945,N_15654,N_15697);
and U15946 (N_15946,N_15686,N_15610);
nor U15947 (N_15947,N_15779,N_15797);
nor U15948 (N_15948,N_15658,N_15681);
nand U15949 (N_15949,N_15732,N_15746);
nor U15950 (N_15950,N_15671,N_15793);
nor U15951 (N_15951,N_15798,N_15786);
and U15952 (N_15952,N_15684,N_15770);
nand U15953 (N_15953,N_15613,N_15646);
nand U15954 (N_15954,N_15625,N_15690);
nor U15955 (N_15955,N_15683,N_15795);
nand U15956 (N_15956,N_15779,N_15761);
nor U15957 (N_15957,N_15795,N_15655);
nand U15958 (N_15958,N_15743,N_15679);
or U15959 (N_15959,N_15726,N_15640);
and U15960 (N_15960,N_15631,N_15719);
and U15961 (N_15961,N_15694,N_15700);
or U15962 (N_15962,N_15749,N_15723);
nor U15963 (N_15963,N_15701,N_15731);
or U15964 (N_15964,N_15737,N_15760);
nor U15965 (N_15965,N_15705,N_15629);
and U15966 (N_15966,N_15671,N_15795);
and U15967 (N_15967,N_15772,N_15654);
or U15968 (N_15968,N_15751,N_15728);
and U15969 (N_15969,N_15623,N_15713);
and U15970 (N_15970,N_15713,N_15695);
nor U15971 (N_15971,N_15621,N_15633);
nor U15972 (N_15972,N_15745,N_15796);
nand U15973 (N_15973,N_15602,N_15773);
nor U15974 (N_15974,N_15699,N_15773);
nor U15975 (N_15975,N_15690,N_15659);
and U15976 (N_15976,N_15669,N_15793);
nand U15977 (N_15977,N_15618,N_15767);
or U15978 (N_15978,N_15684,N_15633);
nor U15979 (N_15979,N_15627,N_15634);
or U15980 (N_15980,N_15610,N_15795);
nand U15981 (N_15981,N_15699,N_15796);
and U15982 (N_15982,N_15726,N_15683);
and U15983 (N_15983,N_15661,N_15793);
and U15984 (N_15984,N_15725,N_15666);
and U15985 (N_15985,N_15775,N_15629);
nand U15986 (N_15986,N_15713,N_15748);
nor U15987 (N_15987,N_15710,N_15717);
nor U15988 (N_15988,N_15637,N_15741);
or U15989 (N_15989,N_15788,N_15738);
and U15990 (N_15990,N_15636,N_15679);
or U15991 (N_15991,N_15621,N_15734);
nand U15992 (N_15992,N_15718,N_15672);
and U15993 (N_15993,N_15623,N_15602);
or U15994 (N_15994,N_15771,N_15693);
or U15995 (N_15995,N_15775,N_15748);
and U15996 (N_15996,N_15658,N_15725);
or U15997 (N_15997,N_15798,N_15682);
and U15998 (N_15998,N_15694,N_15706);
or U15999 (N_15999,N_15776,N_15718);
nor U16000 (N_16000,N_15904,N_15878);
nor U16001 (N_16001,N_15921,N_15851);
or U16002 (N_16002,N_15979,N_15933);
nor U16003 (N_16003,N_15886,N_15838);
or U16004 (N_16004,N_15807,N_15910);
xor U16005 (N_16005,N_15951,N_15948);
and U16006 (N_16006,N_15902,N_15802);
or U16007 (N_16007,N_15827,N_15975);
and U16008 (N_16008,N_15994,N_15907);
nand U16009 (N_16009,N_15954,N_15881);
or U16010 (N_16010,N_15911,N_15997);
and U16011 (N_16011,N_15918,N_15847);
nor U16012 (N_16012,N_15831,N_15836);
or U16013 (N_16013,N_15858,N_15939);
or U16014 (N_16014,N_15984,N_15955);
or U16015 (N_16015,N_15859,N_15866);
or U16016 (N_16016,N_15823,N_15875);
or U16017 (N_16017,N_15914,N_15987);
nor U16018 (N_16018,N_15900,N_15894);
and U16019 (N_16019,N_15821,N_15814);
and U16020 (N_16020,N_15870,N_15924);
nand U16021 (N_16021,N_15868,N_15895);
nor U16022 (N_16022,N_15822,N_15839);
nor U16023 (N_16023,N_15801,N_15972);
and U16024 (N_16024,N_15936,N_15952);
or U16025 (N_16025,N_15983,N_15976);
and U16026 (N_16026,N_15857,N_15968);
nand U16027 (N_16027,N_15824,N_15891);
and U16028 (N_16028,N_15957,N_15956);
nor U16029 (N_16029,N_15930,N_15922);
or U16030 (N_16030,N_15962,N_15920);
nor U16031 (N_16031,N_15999,N_15888);
nand U16032 (N_16032,N_15863,N_15937);
and U16033 (N_16033,N_15817,N_15837);
nor U16034 (N_16034,N_15943,N_15800);
nor U16035 (N_16035,N_15880,N_15861);
nor U16036 (N_16036,N_15805,N_15826);
and U16037 (N_16037,N_15989,N_15816);
nor U16038 (N_16038,N_15990,N_15893);
nand U16039 (N_16039,N_15882,N_15873);
and U16040 (N_16040,N_15867,N_15843);
nand U16041 (N_16041,N_15828,N_15845);
nand U16042 (N_16042,N_15980,N_15929);
and U16043 (N_16043,N_15871,N_15852);
nor U16044 (N_16044,N_15927,N_15909);
nor U16045 (N_16045,N_15825,N_15982);
nand U16046 (N_16046,N_15967,N_15938);
nand U16047 (N_16047,N_15950,N_15865);
nand U16048 (N_16048,N_15813,N_15969);
or U16049 (N_16049,N_15815,N_15963);
nor U16050 (N_16050,N_15945,N_15974);
nor U16051 (N_16051,N_15947,N_15960);
or U16052 (N_16052,N_15915,N_15993);
nand U16053 (N_16053,N_15977,N_15812);
or U16054 (N_16054,N_15884,N_15995);
or U16055 (N_16055,N_15869,N_15832);
nor U16056 (N_16056,N_15917,N_15949);
nor U16057 (N_16057,N_15854,N_15964);
nand U16058 (N_16058,N_15897,N_15804);
nand U16059 (N_16059,N_15874,N_15986);
nand U16060 (N_16060,N_15885,N_15842);
and U16061 (N_16061,N_15953,N_15803);
and U16062 (N_16062,N_15853,N_15942);
nor U16063 (N_16063,N_15889,N_15926);
nor U16064 (N_16064,N_15965,N_15841);
nor U16065 (N_16065,N_15883,N_15806);
nand U16066 (N_16066,N_15988,N_15923);
and U16067 (N_16067,N_15834,N_15961);
nor U16068 (N_16068,N_15855,N_15932);
nand U16069 (N_16069,N_15970,N_15931);
or U16070 (N_16070,N_15919,N_15830);
or U16071 (N_16071,N_15856,N_15925);
and U16072 (N_16072,N_15908,N_15876);
and U16073 (N_16073,N_15809,N_15934);
and U16074 (N_16074,N_15946,N_15844);
nor U16075 (N_16075,N_15912,N_15887);
or U16076 (N_16076,N_15811,N_15860);
nand U16077 (N_16077,N_15890,N_15940);
or U16078 (N_16078,N_15810,N_15906);
nor U16079 (N_16079,N_15941,N_15849);
nor U16080 (N_16080,N_15862,N_15850);
nor U16081 (N_16081,N_15833,N_15835);
nand U16082 (N_16082,N_15991,N_15966);
or U16083 (N_16083,N_15928,N_15981);
nor U16084 (N_16084,N_15819,N_15840);
nand U16085 (N_16085,N_15896,N_15829);
nor U16086 (N_16086,N_15892,N_15905);
nor U16087 (N_16087,N_15944,N_15879);
and U16088 (N_16088,N_15971,N_15998);
or U16089 (N_16089,N_15820,N_15872);
or U16090 (N_16090,N_15808,N_15901);
nand U16091 (N_16091,N_15903,N_15958);
or U16092 (N_16092,N_15899,N_15959);
and U16093 (N_16093,N_15992,N_15877);
and U16094 (N_16094,N_15985,N_15973);
nor U16095 (N_16095,N_15996,N_15848);
or U16096 (N_16096,N_15935,N_15916);
and U16097 (N_16097,N_15846,N_15978);
or U16098 (N_16098,N_15864,N_15818);
or U16099 (N_16099,N_15913,N_15898);
or U16100 (N_16100,N_15959,N_15887);
or U16101 (N_16101,N_15824,N_15978);
nor U16102 (N_16102,N_15906,N_15942);
and U16103 (N_16103,N_15893,N_15885);
and U16104 (N_16104,N_15985,N_15820);
nand U16105 (N_16105,N_15818,N_15944);
or U16106 (N_16106,N_15909,N_15841);
nand U16107 (N_16107,N_15844,N_15951);
and U16108 (N_16108,N_15910,N_15857);
nor U16109 (N_16109,N_15916,N_15801);
or U16110 (N_16110,N_15904,N_15893);
and U16111 (N_16111,N_15912,N_15826);
and U16112 (N_16112,N_15957,N_15838);
and U16113 (N_16113,N_15919,N_15872);
nor U16114 (N_16114,N_15827,N_15891);
nand U16115 (N_16115,N_15822,N_15863);
and U16116 (N_16116,N_15881,N_15941);
nor U16117 (N_16117,N_15851,N_15858);
or U16118 (N_16118,N_15883,N_15808);
and U16119 (N_16119,N_15841,N_15889);
nor U16120 (N_16120,N_15840,N_15828);
nand U16121 (N_16121,N_15946,N_15950);
or U16122 (N_16122,N_15900,N_15807);
nor U16123 (N_16123,N_15947,N_15831);
or U16124 (N_16124,N_15851,N_15929);
or U16125 (N_16125,N_15978,N_15848);
nor U16126 (N_16126,N_15997,N_15865);
or U16127 (N_16127,N_15900,N_15988);
nor U16128 (N_16128,N_15918,N_15836);
nand U16129 (N_16129,N_15924,N_15883);
and U16130 (N_16130,N_15809,N_15961);
or U16131 (N_16131,N_15906,N_15973);
or U16132 (N_16132,N_15880,N_15936);
and U16133 (N_16133,N_15984,N_15810);
nor U16134 (N_16134,N_15966,N_15960);
nand U16135 (N_16135,N_15859,N_15993);
nand U16136 (N_16136,N_15866,N_15823);
or U16137 (N_16137,N_15951,N_15865);
nor U16138 (N_16138,N_15884,N_15895);
or U16139 (N_16139,N_15988,N_15912);
nand U16140 (N_16140,N_15808,N_15988);
nand U16141 (N_16141,N_15841,N_15933);
nor U16142 (N_16142,N_15974,N_15906);
nor U16143 (N_16143,N_15938,N_15997);
and U16144 (N_16144,N_15955,N_15808);
xor U16145 (N_16145,N_15944,N_15876);
nand U16146 (N_16146,N_15881,N_15955);
nand U16147 (N_16147,N_15961,N_15821);
nand U16148 (N_16148,N_15982,N_15817);
nand U16149 (N_16149,N_15824,N_15997);
or U16150 (N_16150,N_15822,N_15940);
and U16151 (N_16151,N_15970,N_15819);
and U16152 (N_16152,N_15898,N_15895);
or U16153 (N_16153,N_15911,N_15932);
nand U16154 (N_16154,N_15829,N_15984);
or U16155 (N_16155,N_15911,N_15953);
and U16156 (N_16156,N_15965,N_15810);
or U16157 (N_16157,N_15870,N_15968);
and U16158 (N_16158,N_15811,N_15897);
or U16159 (N_16159,N_15918,N_15925);
and U16160 (N_16160,N_15944,N_15889);
or U16161 (N_16161,N_15908,N_15808);
and U16162 (N_16162,N_15922,N_15876);
nand U16163 (N_16163,N_15927,N_15872);
and U16164 (N_16164,N_15968,N_15911);
nor U16165 (N_16165,N_15862,N_15889);
and U16166 (N_16166,N_15821,N_15823);
nand U16167 (N_16167,N_15801,N_15800);
and U16168 (N_16168,N_15805,N_15867);
and U16169 (N_16169,N_15876,N_15872);
or U16170 (N_16170,N_15912,N_15948);
nor U16171 (N_16171,N_15936,N_15860);
nor U16172 (N_16172,N_15867,N_15957);
nand U16173 (N_16173,N_15867,N_15952);
nand U16174 (N_16174,N_15953,N_15807);
nand U16175 (N_16175,N_15894,N_15825);
or U16176 (N_16176,N_15995,N_15803);
nand U16177 (N_16177,N_15873,N_15964);
nor U16178 (N_16178,N_15902,N_15846);
nand U16179 (N_16179,N_15933,N_15869);
nor U16180 (N_16180,N_15965,N_15882);
and U16181 (N_16181,N_15802,N_15995);
nand U16182 (N_16182,N_15810,N_15963);
xnor U16183 (N_16183,N_15854,N_15855);
and U16184 (N_16184,N_15946,N_15979);
nor U16185 (N_16185,N_15878,N_15925);
nor U16186 (N_16186,N_15843,N_15913);
and U16187 (N_16187,N_15915,N_15936);
and U16188 (N_16188,N_15891,N_15823);
nand U16189 (N_16189,N_15951,N_15811);
nand U16190 (N_16190,N_15968,N_15850);
nor U16191 (N_16191,N_15927,N_15896);
nor U16192 (N_16192,N_15914,N_15925);
nor U16193 (N_16193,N_15891,N_15923);
nor U16194 (N_16194,N_15860,N_15874);
and U16195 (N_16195,N_15919,N_15991);
nand U16196 (N_16196,N_15922,N_15940);
and U16197 (N_16197,N_15963,N_15927);
or U16198 (N_16198,N_15984,N_15936);
nand U16199 (N_16199,N_15819,N_15842);
and U16200 (N_16200,N_16113,N_16077);
nor U16201 (N_16201,N_16024,N_16175);
and U16202 (N_16202,N_16105,N_16144);
and U16203 (N_16203,N_16095,N_16172);
or U16204 (N_16204,N_16065,N_16187);
nor U16205 (N_16205,N_16013,N_16037);
nor U16206 (N_16206,N_16194,N_16064);
nor U16207 (N_16207,N_16153,N_16168);
or U16208 (N_16208,N_16179,N_16149);
nand U16209 (N_16209,N_16161,N_16189);
and U16210 (N_16210,N_16053,N_16009);
or U16211 (N_16211,N_16129,N_16177);
nor U16212 (N_16212,N_16085,N_16171);
or U16213 (N_16213,N_16030,N_16066);
nor U16214 (N_16214,N_16039,N_16002);
or U16215 (N_16215,N_16103,N_16049);
and U16216 (N_16216,N_16021,N_16032);
nand U16217 (N_16217,N_16136,N_16057);
or U16218 (N_16218,N_16010,N_16089);
nor U16219 (N_16219,N_16001,N_16146);
nand U16220 (N_16220,N_16139,N_16097);
or U16221 (N_16221,N_16166,N_16082);
and U16222 (N_16222,N_16059,N_16068);
and U16223 (N_16223,N_16070,N_16094);
and U16224 (N_16224,N_16034,N_16087);
or U16225 (N_16225,N_16080,N_16164);
nor U16226 (N_16226,N_16140,N_16199);
nor U16227 (N_16227,N_16167,N_16026);
nand U16228 (N_16228,N_16184,N_16124);
nor U16229 (N_16229,N_16008,N_16174);
nor U16230 (N_16230,N_16192,N_16137);
and U16231 (N_16231,N_16151,N_16190);
nor U16232 (N_16232,N_16117,N_16054);
or U16233 (N_16233,N_16035,N_16173);
and U16234 (N_16234,N_16178,N_16165);
nand U16235 (N_16235,N_16060,N_16134);
or U16236 (N_16236,N_16130,N_16047);
nor U16237 (N_16237,N_16118,N_16096);
and U16238 (N_16238,N_16023,N_16188);
and U16239 (N_16239,N_16029,N_16193);
nor U16240 (N_16240,N_16042,N_16091);
and U16241 (N_16241,N_16093,N_16160);
nor U16242 (N_16242,N_16079,N_16111);
and U16243 (N_16243,N_16148,N_16116);
nand U16244 (N_16244,N_16109,N_16098);
or U16245 (N_16245,N_16012,N_16055);
or U16246 (N_16246,N_16185,N_16015);
and U16247 (N_16247,N_16046,N_16033);
and U16248 (N_16248,N_16100,N_16019);
or U16249 (N_16249,N_16126,N_16076);
and U16250 (N_16250,N_16197,N_16004);
nor U16251 (N_16251,N_16000,N_16027);
and U16252 (N_16252,N_16031,N_16169);
nor U16253 (N_16253,N_16075,N_16016);
or U16254 (N_16254,N_16084,N_16186);
nand U16255 (N_16255,N_16198,N_16086);
or U16256 (N_16256,N_16063,N_16036);
and U16257 (N_16257,N_16128,N_16020);
nor U16258 (N_16258,N_16003,N_16011);
nand U16259 (N_16259,N_16088,N_16125);
or U16260 (N_16260,N_16078,N_16112);
nor U16261 (N_16261,N_16069,N_16156);
or U16262 (N_16262,N_16044,N_16041);
nand U16263 (N_16263,N_16145,N_16132);
nor U16264 (N_16264,N_16119,N_16017);
nor U16265 (N_16265,N_16007,N_16061);
nor U16266 (N_16266,N_16183,N_16050);
nor U16267 (N_16267,N_16018,N_16045);
or U16268 (N_16268,N_16141,N_16181);
or U16269 (N_16269,N_16022,N_16162);
and U16270 (N_16270,N_16147,N_16081);
nand U16271 (N_16271,N_16051,N_16028);
and U16272 (N_16272,N_16014,N_16180);
nor U16273 (N_16273,N_16101,N_16135);
and U16274 (N_16274,N_16196,N_16107);
xnor U16275 (N_16275,N_16052,N_16074);
nand U16276 (N_16276,N_16163,N_16072);
and U16277 (N_16277,N_16092,N_16108);
nand U16278 (N_16278,N_16090,N_16071);
nor U16279 (N_16279,N_16005,N_16158);
or U16280 (N_16280,N_16038,N_16157);
and U16281 (N_16281,N_16182,N_16131);
or U16282 (N_16282,N_16025,N_16056);
nor U16283 (N_16283,N_16143,N_16191);
or U16284 (N_16284,N_16121,N_16138);
nor U16285 (N_16285,N_16048,N_16102);
or U16286 (N_16286,N_16155,N_16142);
or U16287 (N_16287,N_16133,N_16127);
nand U16288 (N_16288,N_16120,N_16114);
nand U16289 (N_16289,N_16154,N_16115);
or U16290 (N_16290,N_16110,N_16006);
nand U16291 (N_16291,N_16104,N_16123);
nand U16292 (N_16292,N_16152,N_16083);
nor U16293 (N_16293,N_16176,N_16122);
or U16294 (N_16294,N_16195,N_16058);
or U16295 (N_16295,N_16170,N_16067);
or U16296 (N_16296,N_16043,N_16150);
nor U16297 (N_16297,N_16159,N_16062);
and U16298 (N_16298,N_16099,N_16040);
or U16299 (N_16299,N_16106,N_16073);
nor U16300 (N_16300,N_16158,N_16074);
nor U16301 (N_16301,N_16049,N_16136);
and U16302 (N_16302,N_16113,N_16061);
and U16303 (N_16303,N_16049,N_16146);
or U16304 (N_16304,N_16056,N_16082);
or U16305 (N_16305,N_16059,N_16062);
or U16306 (N_16306,N_16129,N_16009);
and U16307 (N_16307,N_16157,N_16185);
nand U16308 (N_16308,N_16026,N_16051);
and U16309 (N_16309,N_16037,N_16132);
or U16310 (N_16310,N_16079,N_16113);
nor U16311 (N_16311,N_16071,N_16002);
nand U16312 (N_16312,N_16060,N_16074);
nand U16313 (N_16313,N_16009,N_16101);
nand U16314 (N_16314,N_16147,N_16188);
and U16315 (N_16315,N_16129,N_16006);
and U16316 (N_16316,N_16021,N_16103);
and U16317 (N_16317,N_16166,N_16097);
xor U16318 (N_16318,N_16060,N_16120);
and U16319 (N_16319,N_16151,N_16003);
or U16320 (N_16320,N_16173,N_16001);
or U16321 (N_16321,N_16163,N_16025);
or U16322 (N_16322,N_16175,N_16044);
and U16323 (N_16323,N_16146,N_16142);
nor U16324 (N_16324,N_16030,N_16044);
nand U16325 (N_16325,N_16150,N_16033);
and U16326 (N_16326,N_16064,N_16199);
nand U16327 (N_16327,N_16047,N_16015);
nor U16328 (N_16328,N_16177,N_16061);
nand U16329 (N_16329,N_16014,N_16028);
and U16330 (N_16330,N_16120,N_16032);
xnor U16331 (N_16331,N_16108,N_16110);
xor U16332 (N_16332,N_16106,N_16091);
and U16333 (N_16333,N_16055,N_16073);
and U16334 (N_16334,N_16037,N_16186);
nor U16335 (N_16335,N_16090,N_16092);
or U16336 (N_16336,N_16050,N_16163);
nand U16337 (N_16337,N_16128,N_16070);
and U16338 (N_16338,N_16024,N_16137);
or U16339 (N_16339,N_16020,N_16070);
and U16340 (N_16340,N_16071,N_16109);
and U16341 (N_16341,N_16171,N_16139);
and U16342 (N_16342,N_16000,N_16155);
nand U16343 (N_16343,N_16146,N_16067);
and U16344 (N_16344,N_16048,N_16001);
and U16345 (N_16345,N_16030,N_16070);
nand U16346 (N_16346,N_16034,N_16133);
nor U16347 (N_16347,N_16086,N_16092);
nand U16348 (N_16348,N_16178,N_16058);
xor U16349 (N_16349,N_16025,N_16052);
nor U16350 (N_16350,N_16131,N_16082);
nand U16351 (N_16351,N_16074,N_16082);
nand U16352 (N_16352,N_16091,N_16072);
nor U16353 (N_16353,N_16189,N_16155);
nand U16354 (N_16354,N_16162,N_16164);
and U16355 (N_16355,N_16197,N_16175);
or U16356 (N_16356,N_16020,N_16122);
nor U16357 (N_16357,N_16060,N_16158);
nand U16358 (N_16358,N_16047,N_16021);
nand U16359 (N_16359,N_16180,N_16184);
or U16360 (N_16360,N_16081,N_16049);
and U16361 (N_16361,N_16054,N_16094);
and U16362 (N_16362,N_16178,N_16005);
nand U16363 (N_16363,N_16191,N_16084);
nor U16364 (N_16364,N_16012,N_16192);
nor U16365 (N_16365,N_16075,N_16063);
or U16366 (N_16366,N_16119,N_16149);
nand U16367 (N_16367,N_16047,N_16121);
nor U16368 (N_16368,N_16061,N_16014);
nor U16369 (N_16369,N_16167,N_16118);
and U16370 (N_16370,N_16058,N_16165);
nor U16371 (N_16371,N_16045,N_16037);
and U16372 (N_16372,N_16159,N_16138);
nor U16373 (N_16373,N_16195,N_16172);
nor U16374 (N_16374,N_16164,N_16157);
or U16375 (N_16375,N_16026,N_16044);
or U16376 (N_16376,N_16057,N_16160);
or U16377 (N_16377,N_16199,N_16024);
nor U16378 (N_16378,N_16178,N_16129);
nand U16379 (N_16379,N_16006,N_16096);
nand U16380 (N_16380,N_16105,N_16180);
nand U16381 (N_16381,N_16172,N_16037);
nand U16382 (N_16382,N_16180,N_16109);
and U16383 (N_16383,N_16126,N_16196);
or U16384 (N_16384,N_16100,N_16115);
and U16385 (N_16385,N_16127,N_16175);
nand U16386 (N_16386,N_16162,N_16001);
nor U16387 (N_16387,N_16188,N_16047);
nor U16388 (N_16388,N_16179,N_16023);
and U16389 (N_16389,N_16005,N_16128);
and U16390 (N_16390,N_16036,N_16090);
or U16391 (N_16391,N_16059,N_16185);
nand U16392 (N_16392,N_16071,N_16046);
nand U16393 (N_16393,N_16010,N_16123);
nor U16394 (N_16394,N_16096,N_16058);
nor U16395 (N_16395,N_16023,N_16029);
nor U16396 (N_16396,N_16119,N_16046);
or U16397 (N_16397,N_16142,N_16073);
or U16398 (N_16398,N_16039,N_16020);
or U16399 (N_16399,N_16016,N_16010);
and U16400 (N_16400,N_16372,N_16222);
or U16401 (N_16401,N_16244,N_16353);
or U16402 (N_16402,N_16348,N_16397);
nor U16403 (N_16403,N_16236,N_16294);
nand U16404 (N_16404,N_16333,N_16351);
nor U16405 (N_16405,N_16325,N_16335);
nor U16406 (N_16406,N_16210,N_16300);
or U16407 (N_16407,N_16259,N_16311);
and U16408 (N_16408,N_16323,N_16322);
nand U16409 (N_16409,N_16290,N_16398);
nor U16410 (N_16410,N_16279,N_16376);
nand U16411 (N_16411,N_16257,N_16378);
nor U16412 (N_16412,N_16373,N_16340);
and U16413 (N_16413,N_16223,N_16281);
nor U16414 (N_16414,N_16332,N_16326);
nor U16415 (N_16415,N_16374,N_16350);
and U16416 (N_16416,N_16271,N_16260);
nor U16417 (N_16417,N_16264,N_16215);
and U16418 (N_16418,N_16203,N_16273);
nor U16419 (N_16419,N_16337,N_16369);
nand U16420 (N_16420,N_16349,N_16368);
and U16421 (N_16421,N_16318,N_16390);
or U16422 (N_16422,N_16387,N_16352);
or U16423 (N_16423,N_16287,N_16275);
and U16424 (N_16424,N_16321,N_16317);
or U16425 (N_16425,N_16239,N_16367);
and U16426 (N_16426,N_16213,N_16250);
nor U16427 (N_16427,N_16370,N_16269);
nor U16428 (N_16428,N_16245,N_16396);
nand U16429 (N_16429,N_16230,N_16226);
and U16430 (N_16430,N_16330,N_16320);
and U16431 (N_16431,N_16209,N_16356);
and U16432 (N_16432,N_16355,N_16288);
and U16433 (N_16433,N_16202,N_16216);
or U16434 (N_16434,N_16383,N_16211);
nor U16435 (N_16435,N_16240,N_16346);
nor U16436 (N_16436,N_16261,N_16360);
nor U16437 (N_16437,N_16345,N_16225);
and U16438 (N_16438,N_16289,N_16357);
nand U16439 (N_16439,N_16293,N_16285);
nor U16440 (N_16440,N_16339,N_16319);
or U16441 (N_16441,N_16208,N_16393);
nand U16442 (N_16442,N_16305,N_16381);
or U16443 (N_16443,N_16299,N_16344);
nor U16444 (N_16444,N_16313,N_16280);
nand U16445 (N_16445,N_16206,N_16301);
and U16446 (N_16446,N_16231,N_16292);
or U16447 (N_16447,N_16302,N_16243);
and U16448 (N_16448,N_16291,N_16272);
nand U16449 (N_16449,N_16395,N_16307);
nor U16450 (N_16450,N_16265,N_16394);
nand U16451 (N_16451,N_16268,N_16392);
nand U16452 (N_16452,N_16227,N_16359);
nand U16453 (N_16453,N_16324,N_16286);
and U16454 (N_16454,N_16312,N_16229);
or U16455 (N_16455,N_16309,N_16364);
or U16456 (N_16456,N_16237,N_16331);
nand U16457 (N_16457,N_16253,N_16371);
and U16458 (N_16458,N_16219,N_16214);
nand U16459 (N_16459,N_16232,N_16385);
and U16460 (N_16460,N_16252,N_16251);
nor U16461 (N_16461,N_16218,N_16316);
and U16462 (N_16462,N_16388,N_16343);
nor U16463 (N_16463,N_16362,N_16212);
nand U16464 (N_16464,N_16283,N_16262);
nor U16465 (N_16465,N_16329,N_16217);
nor U16466 (N_16466,N_16327,N_16310);
nor U16467 (N_16467,N_16246,N_16205);
nand U16468 (N_16468,N_16270,N_16242);
nand U16469 (N_16469,N_16200,N_16278);
or U16470 (N_16470,N_16201,N_16220);
or U16471 (N_16471,N_16334,N_16267);
and U16472 (N_16472,N_16255,N_16336);
and U16473 (N_16473,N_16303,N_16306);
and U16474 (N_16474,N_16258,N_16233);
nand U16475 (N_16475,N_16391,N_16342);
nand U16476 (N_16476,N_16241,N_16314);
and U16477 (N_16477,N_16399,N_16254);
and U16478 (N_16478,N_16328,N_16224);
or U16479 (N_16479,N_16266,N_16238);
nand U16480 (N_16480,N_16384,N_16304);
nand U16481 (N_16481,N_16379,N_16375);
or U16482 (N_16482,N_16234,N_16365);
nand U16483 (N_16483,N_16377,N_16274);
and U16484 (N_16484,N_16380,N_16297);
nor U16485 (N_16485,N_16207,N_16296);
nand U16486 (N_16486,N_16363,N_16358);
nand U16487 (N_16487,N_16204,N_16247);
nand U16488 (N_16488,N_16249,N_16389);
nand U16489 (N_16489,N_16347,N_16277);
nor U16490 (N_16490,N_16256,N_16263);
and U16491 (N_16491,N_16284,N_16361);
and U16492 (N_16492,N_16341,N_16276);
nor U16493 (N_16493,N_16228,N_16382);
and U16494 (N_16494,N_16235,N_16298);
and U16495 (N_16495,N_16366,N_16282);
and U16496 (N_16496,N_16248,N_16221);
or U16497 (N_16497,N_16295,N_16386);
nand U16498 (N_16498,N_16354,N_16315);
nand U16499 (N_16499,N_16338,N_16308);
or U16500 (N_16500,N_16247,N_16206);
nand U16501 (N_16501,N_16212,N_16383);
nand U16502 (N_16502,N_16352,N_16249);
or U16503 (N_16503,N_16391,N_16325);
and U16504 (N_16504,N_16275,N_16331);
or U16505 (N_16505,N_16318,N_16331);
or U16506 (N_16506,N_16229,N_16300);
and U16507 (N_16507,N_16247,N_16288);
and U16508 (N_16508,N_16341,N_16201);
or U16509 (N_16509,N_16375,N_16359);
and U16510 (N_16510,N_16242,N_16347);
nor U16511 (N_16511,N_16267,N_16347);
nand U16512 (N_16512,N_16227,N_16229);
and U16513 (N_16513,N_16330,N_16321);
and U16514 (N_16514,N_16341,N_16292);
or U16515 (N_16515,N_16382,N_16220);
nor U16516 (N_16516,N_16228,N_16332);
xnor U16517 (N_16517,N_16217,N_16325);
or U16518 (N_16518,N_16397,N_16340);
and U16519 (N_16519,N_16318,N_16350);
or U16520 (N_16520,N_16320,N_16366);
or U16521 (N_16521,N_16283,N_16212);
and U16522 (N_16522,N_16229,N_16209);
nor U16523 (N_16523,N_16226,N_16391);
nand U16524 (N_16524,N_16308,N_16313);
nor U16525 (N_16525,N_16277,N_16349);
or U16526 (N_16526,N_16223,N_16218);
nor U16527 (N_16527,N_16207,N_16345);
and U16528 (N_16528,N_16275,N_16399);
nor U16529 (N_16529,N_16261,N_16318);
nor U16530 (N_16530,N_16291,N_16259);
and U16531 (N_16531,N_16297,N_16266);
or U16532 (N_16532,N_16314,N_16308);
nor U16533 (N_16533,N_16277,N_16247);
or U16534 (N_16534,N_16399,N_16223);
or U16535 (N_16535,N_16347,N_16327);
or U16536 (N_16536,N_16322,N_16390);
nor U16537 (N_16537,N_16264,N_16261);
or U16538 (N_16538,N_16292,N_16319);
or U16539 (N_16539,N_16316,N_16295);
nand U16540 (N_16540,N_16251,N_16243);
nand U16541 (N_16541,N_16243,N_16367);
or U16542 (N_16542,N_16232,N_16235);
nand U16543 (N_16543,N_16356,N_16233);
nand U16544 (N_16544,N_16246,N_16396);
nor U16545 (N_16545,N_16282,N_16347);
nor U16546 (N_16546,N_16381,N_16288);
nand U16547 (N_16547,N_16352,N_16365);
or U16548 (N_16548,N_16301,N_16263);
and U16549 (N_16549,N_16395,N_16269);
and U16550 (N_16550,N_16240,N_16293);
nor U16551 (N_16551,N_16232,N_16397);
nand U16552 (N_16552,N_16329,N_16398);
and U16553 (N_16553,N_16383,N_16368);
nor U16554 (N_16554,N_16248,N_16373);
nand U16555 (N_16555,N_16378,N_16313);
or U16556 (N_16556,N_16352,N_16348);
or U16557 (N_16557,N_16382,N_16237);
and U16558 (N_16558,N_16310,N_16201);
or U16559 (N_16559,N_16288,N_16380);
nand U16560 (N_16560,N_16298,N_16311);
nor U16561 (N_16561,N_16210,N_16388);
or U16562 (N_16562,N_16214,N_16302);
xnor U16563 (N_16563,N_16363,N_16398);
nand U16564 (N_16564,N_16200,N_16293);
nor U16565 (N_16565,N_16204,N_16330);
or U16566 (N_16566,N_16284,N_16342);
nor U16567 (N_16567,N_16391,N_16320);
and U16568 (N_16568,N_16361,N_16209);
xor U16569 (N_16569,N_16345,N_16244);
nor U16570 (N_16570,N_16352,N_16311);
nor U16571 (N_16571,N_16320,N_16220);
nand U16572 (N_16572,N_16349,N_16396);
nor U16573 (N_16573,N_16337,N_16373);
or U16574 (N_16574,N_16353,N_16233);
nor U16575 (N_16575,N_16317,N_16358);
and U16576 (N_16576,N_16377,N_16209);
nand U16577 (N_16577,N_16209,N_16367);
or U16578 (N_16578,N_16327,N_16295);
nor U16579 (N_16579,N_16242,N_16380);
or U16580 (N_16580,N_16368,N_16297);
or U16581 (N_16581,N_16370,N_16365);
and U16582 (N_16582,N_16383,N_16396);
nor U16583 (N_16583,N_16254,N_16333);
or U16584 (N_16584,N_16257,N_16307);
nor U16585 (N_16585,N_16245,N_16364);
nor U16586 (N_16586,N_16236,N_16332);
and U16587 (N_16587,N_16333,N_16288);
nor U16588 (N_16588,N_16399,N_16210);
or U16589 (N_16589,N_16201,N_16232);
and U16590 (N_16590,N_16218,N_16301);
nand U16591 (N_16591,N_16379,N_16244);
nand U16592 (N_16592,N_16337,N_16380);
or U16593 (N_16593,N_16379,N_16348);
and U16594 (N_16594,N_16372,N_16237);
and U16595 (N_16595,N_16343,N_16394);
and U16596 (N_16596,N_16274,N_16374);
and U16597 (N_16597,N_16360,N_16239);
nor U16598 (N_16598,N_16262,N_16343);
and U16599 (N_16599,N_16303,N_16268);
nand U16600 (N_16600,N_16427,N_16417);
nor U16601 (N_16601,N_16505,N_16448);
nor U16602 (N_16602,N_16476,N_16481);
nand U16603 (N_16603,N_16435,N_16533);
nand U16604 (N_16604,N_16509,N_16511);
and U16605 (N_16605,N_16591,N_16548);
and U16606 (N_16606,N_16491,N_16569);
and U16607 (N_16607,N_16459,N_16438);
nor U16608 (N_16608,N_16464,N_16447);
or U16609 (N_16609,N_16508,N_16560);
nand U16610 (N_16610,N_16406,N_16578);
and U16611 (N_16611,N_16573,N_16478);
and U16612 (N_16612,N_16428,N_16502);
nor U16613 (N_16613,N_16472,N_16504);
nand U16614 (N_16614,N_16544,N_16421);
or U16615 (N_16615,N_16506,N_16598);
or U16616 (N_16616,N_16554,N_16517);
nor U16617 (N_16617,N_16500,N_16561);
nand U16618 (N_16618,N_16543,N_16553);
or U16619 (N_16619,N_16531,N_16513);
and U16620 (N_16620,N_16430,N_16575);
or U16621 (N_16621,N_16455,N_16572);
or U16622 (N_16622,N_16526,N_16423);
nand U16623 (N_16623,N_16456,N_16532);
or U16624 (N_16624,N_16496,N_16462);
nand U16625 (N_16625,N_16530,N_16579);
and U16626 (N_16626,N_16468,N_16418);
or U16627 (N_16627,N_16477,N_16527);
nor U16628 (N_16628,N_16588,N_16539);
nor U16629 (N_16629,N_16587,N_16487);
xor U16630 (N_16630,N_16516,N_16484);
or U16631 (N_16631,N_16586,N_16465);
nor U16632 (N_16632,N_16528,N_16449);
and U16633 (N_16633,N_16415,N_16489);
nor U16634 (N_16634,N_16576,N_16471);
or U16635 (N_16635,N_16589,N_16545);
nand U16636 (N_16636,N_16454,N_16494);
nand U16637 (N_16637,N_16451,N_16542);
and U16638 (N_16638,N_16488,N_16410);
nor U16639 (N_16639,N_16444,N_16522);
nor U16640 (N_16640,N_16458,N_16479);
nor U16641 (N_16641,N_16424,N_16407);
nand U16642 (N_16642,N_16552,N_16434);
or U16643 (N_16643,N_16400,N_16453);
or U16644 (N_16644,N_16467,N_16597);
nand U16645 (N_16645,N_16524,N_16426);
nand U16646 (N_16646,N_16432,N_16409);
and U16647 (N_16647,N_16446,N_16596);
xor U16648 (N_16648,N_16535,N_16495);
or U16649 (N_16649,N_16412,N_16503);
nand U16650 (N_16650,N_16482,N_16583);
nor U16651 (N_16651,N_16450,N_16599);
nor U16652 (N_16652,N_16490,N_16515);
and U16653 (N_16653,N_16470,N_16556);
nand U16654 (N_16654,N_16562,N_16403);
nor U16655 (N_16655,N_16568,N_16540);
or U16656 (N_16656,N_16420,N_16534);
and U16657 (N_16657,N_16433,N_16520);
nand U16658 (N_16658,N_16431,N_16559);
and U16659 (N_16659,N_16518,N_16402);
nand U16660 (N_16660,N_16590,N_16404);
and U16661 (N_16661,N_16564,N_16510);
and U16662 (N_16662,N_16538,N_16567);
and U16663 (N_16663,N_16436,N_16512);
nand U16664 (N_16664,N_16577,N_16469);
nor U16665 (N_16665,N_16519,N_16550);
or U16666 (N_16666,N_16595,N_16525);
and U16667 (N_16667,N_16537,N_16440);
nand U16668 (N_16668,N_16486,N_16460);
or U16669 (N_16669,N_16461,N_16551);
and U16670 (N_16670,N_16582,N_16563);
or U16671 (N_16671,N_16584,N_16485);
and U16672 (N_16672,N_16442,N_16593);
and U16673 (N_16673,N_16555,N_16501);
nor U16674 (N_16674,N_16483,N_16523);
nand U16675 (N_16675,N_16429,N_16413);
and U16676 (N_16676,N_16514,N_16529);
nand U16677 (N_16677,N_16441,N_16457);
or U16678 (N_16678,N_16422,N_16414);
or U16679 (N_16679,N_16557,N_16594);
and U16680 (N_16680,N_16463,N_16498);
nand U16681 (N_16681,N_16425,N_16493);
or U16682 (N_16682,N_16492,N_16549);
nor U16683 (N_16683,N_16565,N_16497);
nor U16684 (N_16684,N_16580,N_16408);
nor U16685 (N_16685,N_16547,N_16452);
or U16686 (N_16686,N_16574,N_16480);
and U16687 (N_16687,N_16592,N_16566);
or U16688 (N_16688,N_16570,N_16581);
nor U16689 (N_16689,N_16536,N_16437);
nor U16690 (N_16690,N_16499,N_16439);
nor U16691 (N_16691,N_16541,N_16571);
and U16692 (N_16692,N_16416,N_16558);
nand U16693 (N_16693,N_16419,N_16401);
nor U16694 (N_16694,N_16474,N_16405);
and U16695 (N_16695,N_16443,N_16585);
or U16696 (N_16696,N_16473,N_16475);
nor U16697 (N_16697,N_16521,N_16466);
and U16698 (N_16698,N_16411,N_16546);
nand U16699 (N_16699,N_16445,N_16507);
or U16700 (N_16700,N_16499,N_16575);
nor U16701 (N_16701,N_16483,N_16513);
xnor U16702 (N_16702,N_16560,N_16422);
nor U16703 (N_16703,N_16541,N_16554);
or U16704 (N_16704,N_16560,N_16421);
nand U16705 (N_16705,N_16534,N_16470);
and U16706 (N_16706,N_16483,N_16552);
nand U16707 (N_16707,N_16554,N_16426);
or U16708 (N_16708,N_16499,N_16450);
nand U16709 (N_16709,N_16497,N_16572);
nor U16710 (N_16710,N_16449,N_16541);
xnor U16711 (N_16711,N_16578,N_16432);
and U16712 (N_16712,N_16549,N_16550);
nand U16713 (N_16713,N_16463,N_16595);
or U16714 (N_16714,N_16417,N_16403);
nand U16715 (N_16715,N_16550,N_16427);
or U16716 (N_16716,N_16420,N_16431);
and U16717 (N_16717,N_16544,N_16553);
nand U16718 (N_16718,N_16587,N_16550);
nor U16719 (N_16719,N_16547,N_16561);
and U16720 (N_16720,N_16477,N_16498);
and U16721 (N_16721,N_16557,N_16533);
nor U16722 (N_16722,N_16414,N_16467);
nor U16723 (N_16723,N_16520,N_16517);
and U16724 (N_16724,N_16423,N_16536);
nand U16725 (N_16725,N_16471,N_16422);
nor U16726 (N_16726,N_16572,N_16553);
and U16727 (N_16727,N_16463,N_16563);
nor U16728 (N_16728,N_16588,N_16431);
xor U16729 (N_16729,N_16411,N_16430);
and U16730 (N_16730,N_16465,N_16564);
and U16731 (N_16731,N_16575,N_16522);
nand U16732 (N_16732,N_16416,N_16449);
nor U16733 (N_16733,N_16531,N_16586);
and U16734 (N_16734,N_16578,N_16542);
or U16735 (N_16735,N_16529,N_16481);
and U16736 (N_16736,N_16408,N_16537);
xnor U16737 (N_16737,N_16426,N_16559);
nand U16738 (N_16738,N_16422,N_16533);
or U16739 (N_16739,N_16429,N_16524);
nand U16740 (N_16740,N_16538,N_16594);
and U16741 (N_16741,N_16531,N_16410);
nand U16742 (N_16742,N_16438,N_16479);
or U16743 (N_16743,N_16541,N_16584);
and U16744 (N_16744,N_16513,N_16451);
nor U16745 (N_16745,N_16444,N_16513);
and U16746 (N_16746,N_16530,N_16514);
nor U16747 (N_16747,N_16508,N_16515);
nor U16748 (N_16748,N_16487,N_16448);
nand U16749 (N_16749,N_16497,N_16590);
and U16750 (N_16750,N_16415,N_16501);
nand U16751 (N_16751,N_16469,N_16433);
nand U16752 (N_16752,N_16538,N_16412);
and U16753 (N_16753,N_16575,N_16469);
or U16754 (N_16754,N_16537,N_16552);
or U16755 (N_16755,N_16446,N_16569);
or U16756 (N_16756,N_16412,N_16444);
nand U16757 (N_16757,N_16526,N_16459);
nor U16758 (N_16758,N_16599,N_16425);
nand U16759 (N_16759,N_16501,N_16413);
or U16760 (N_16760,N_16485,N_16533);
or U16761 (N_16761,N_16540,N_16582);
or U16762 (N_16762,N_16563,N_16551);
and U16763 (N_16763,N_16553,N_16416);
or U16764 (N_16764,N_16419,N_16434);
nor U16765 (N_16765,N_16599,N_16587);
and U16766 (N_16766,N_16407,N_16509);
or U16767 (N_16767,N_16406,N_16562);
nor U16768 (N_16768,N_16533,N_16434);
nor U16769 (N_16769,N_16417,N_16580);
or U16770 (N_16770,N_16519,N_16524);
nand U16771 (N_16771,N_16505,N_16442);
nor U16772 (N_16772,N_16514,N_16598);
nor U16773 (N_16773,N_16553,N_16489);
nand U16774 (N_16774,N_16400,N_16495);
or U16775 (N_16775,N_16452,N_16417);
nor U16776 (N_16776,N_16570,N_16577);
or U16777 (N_16777,N_16435,N_16428);
and U16778 (N_16778,N_16454,N_16572);
nor U16779 (N_16779,N_16494,N_16576);
nand U16780 (N_16780,N_16461,N_16502);
or U16781 (N_16781,N_16573,N_16562);
and U16782 (N_16782,N_16561,N_16582);
nand U16783 (N_16783,N_16470,N_16537);
nand U16784 (N_16784,N_16466,N_16598);
or U16785 (N_16785,N_16490,N_16417);
or U16786 (N_16786,N_16496,N_16565);
nor U16787 (N_16787,N_16517,N_16443);
or U16788 (N_16788,N_16488,N_16549);
or U16789 (N_16789,N_16410,N_16460);
and U16790 (N_16790,N_16486,N_16515);
nand U16791 (N_16791,N_16536,N_16460);
and U16792 (N_16792,N_16515,N_16531);
nand U16793 (N_16793,N_16510,N_16433);
and U16794 (N_16794,N_16403,N_16587);
and U16795 (N_16795,N_16545,N_16449);
xnor U16796 (N_16796,N_16585,N_16507);
nand U16797 (N_16797,N_16475,N_16555);
nand U16798 (N_16798,N_16543,N_16585);
nand U16799 (N_16799,N_16501,N_16497);
and U16800 (N_16800,N_16735,N_16704);
xor U16801 (N_16801,N_16649,N_16729);
or U16802 (N_16802,N_16733,N_16744);
nor U16803 (N_16803,N_16765,N_16673);
and U16804 (N_16804,N_16776,N_16715);
nand U16805 (N_16805,N_16721,N_16774);
and U16806 (N_16806,N_16778,N_16630);
nand U16807 (N_16807,N_16753,N_16786);
nor U16808 (N_16808,N_16693,N_16757);
nor U16809 (N_16809,N_16615,N_16796);
or U16810 (N_16810,N_16766,N_16797);
and U16811 (N_16811,N_16707,N_16712);
and U16812 (N_16812,N_16708,N_16665);
and U16813 (N_16813,N_16762,N_16756);
or U16814 (N_16814,N_16706,N_16664);
nand U16815 (N_16815,N_16697,N_16679);
or U16816 (N_16816,N_16613,N_16621);
and U16817 (N_16817,N_16677,N_16675);
nor U16818 (N_16818,N_16787,N_16754);
or U16819 (N_16819,N_16763,N_16610);
or U16820 (N_16820,N_16768,N_16623);
or U16821 (N_16821,N_16724,N_16688);
nor U16822 (N_16822,N_16653,N_16777);
or U16823 (N_16823,N_16628,N_16607);
nor U16824 (N_16824,N_16798,N_16655);
nand U16825 (N_16825,N_16782,N_16726);
nand U16826 (N_16826,N_16760,N_16602);
nand U16827 (N_16827,N_16685,N_16625);
nor U16828 (N_16828,N_16711,N_16785);
nand U16829 (N_16829,N_16644,N_16738);
and U16830 (N_16830,N_16752,N_16694);
or U16831 (N_16831,N_16629,N_16784);
and U16832 (N_16832,N_16667,N_16713);
and U16833 (N_16833,N_16745,N_16661);
or U16834 (N_16834,N_16663,N_16641);
and U16835 (N_16835,N_16718,N_16692);
and U16836 (N_16836,N_16666,N_16648);
and U16837 (N_16837,N_16646,N_16794);
and U16838 (N_16838,N_16714,N_16651);
and U16839 (N_16839,N_16700,N_16790);
or U16840 (N_16840,N_16720,N_16639);
nand U16841 (N_16841,N_16702,N_16678);
nand U16842 (N_16842,N_16795,N_16771);
or U16843 (N_16843,N_16671,N_16716);
and U16844 (N_16844,N_16624,N_16789);
or U16845 (N_16845,N_16696,N_16660);
and U16846 (N_16846,N_16608,N_16681);
and U16847 (N_16847,N_16632,N_16638);
or U16848 (N_16848,N_16633,N_16634);
nor U16849 (N_16849,N_16670,N_16650);
and U16850 (N_16850,N_16751,N_16761);
or U16851 (N_16851,N_16618,N_16699);
and U16852 (N_16852,N_16643,N_16627);
nor U16853 (N_16853,N_16727,N_16701);
or U16854 (N_16854,N_16631,N_16769);
nand U16855 (N_16855,N_16799,N_16674);
nand U16856 (N_16856,N_16747,N_16705);
nor U16857 (N_16857,N_16779,N_16657);
nor U16858 (N_16858,N_16767,N_16686);
nor U16859 (N_16859,N_16749,N_16717);
nor U16860 (N_16860,N_16659,N_16750);
nor U16861 (N_16861,N_16676,N_16755);
nor U16862 (N_16862,N_16770,N_16680);
or U16863 (N_16863,N_16626,N_16672);
and U16864 (N_16864,N_16605,N_16722);
or U16865 (N_16865,N_16611,N_16736);
or U16866 (N_16866,N_16603,N_16617);
nor U16867 (N_16867,N_16645,N_16743);
nand U16868 (N_16868,N_16710,N_16616);
nand U16869 (N_16869,N_16601,N_16619);
and U16870 (N_16870,N_16773,N_16709);
and U16871 (N_16871,N_16662,N_16636);
and U16872 (N_16872,N_16654,N_16698);
nand U16873 (N_16873,N_16604,N_16691);
or U16874 (N_16874,N_16780,N_16637);
nor U16875 (N_16875,N_16606,N_16719);
and U16876 (N_16876,N_16759,N_16748);
nor U16877 (N_16877,N_16781,N_16791);
nor U16878 (N_16878,N_16622,N_16741);
or U16879 (N_16879,N_16620,N_16723);
and U16880 (N_16880,N_16668,N_16758);
and U16881 (N_16881,N_16793,N_16746);
or U16882 (N_16882,N_16734,N_16742);
and U16883 (N_16883,N_16656,N_16732);
and U16884 (N_16884,N_16725,N_16772);
nor U16885 (N_16885,N_16642,N_16737);
nor U16886 (N_16886,N_16775,N_16600);
or U16887 (N_16887,N_16703,N_16792);
and U16888 (N_16888,N_16684,N_16728);
nand U16889 (N_16889,N_16640,N_16682);
nand U16890 (N_16890,N_16683,N_16609);
nand U16891 (N_16891,N_16687,N_16612);
and U16892 (N_16892,N_16788,N_16614);
or U16893 (N_16893,N_16658,N_16647);
and U16894 (N_16894,N_16764,N_16695);
and U16895 (N_16895,N_16652,N_16669);
nor U16896 (N_16896,N_16731,N_16689);
and U16897 (N_16897,N_16783,N_16739);
nand U16898 (N_16898,N_16730,N_16635);
nor U16899 (N_16899,N_16740,N_16690);
or U16900 (N_16900,N_16616,N_16745);
or U16901 (N_16901,N_16603,N_16747);
or U16902 (N_16902,N_16772,N_16699);
or U16903 (N_16903,N_16616,N_16740);
nor U16904 (N_16904,N_16682,N_16734);
and U16905 (N_16905,N_16634,N_16698);
or U16906 (N_16906,N_16775,N_16678);
or U16907 (N_16907,N_16642,N_16603);
or U16908 (N_16908,N_16696,N_16665);
nor U16909 (N_16909,N_16742,N_16739);
or U16910 (N_16910,N_16625,N_16614);
or U16911 (N_16911,N_16636,N_16753);
nand U16912 (N_16912,N_16654,N_16766);
nor U16913 (N_16913,N_16788,N_16670);
and U16914 (N_16914,N_16632,N_16639);
nor U16915 (N_16915,N_16691,N_16768);
and U16916 (N_16916,N_16726,N_16781);
or U16917 (N_16917,N_16733,N_16750);
and U16918 (N_16918,N_16703,N_16769);
nor U16919 (N_16919,N_16647,N_16706);
or U16920 (N_16920,N_16712,N_16720);
nand U16921 (N_16921,N_16696,N_16738);
nand U16922 (N_16922,N_16682,N_16680);
nor U16923 (N_16923,N_16741,N_16725);
and U16924 (N_16924,N_16787,N_16633);
or U16925 (N_16925,N_16704,N_16614);
and U16926 (N_16926,N_16651,N_16798);
or U16927 (N_16927,N_16756,N_16793);
nand U16928 (N_16928,N_16777,N_16631);
or U16929 (N_16929,N_16647,N_16602);
nor U16930 (N_16930,N_16792,N_16795);
and U16931 (N_16931,N_16745,N_16670);
nor U16932 (N_16932,N_16785,N_16773);
nand U16933 (N_16933,N_16690,N_16620);
or U16934 (N_16934,N_16653,N_16799);
and U16935 (N_16935,N_16619,N_16748);
nor U16936 (N_16936,N_16716,N_16767);
nand U16937 (N_16937,N_16621,N_16654);
and U16938 (N_16938,N_16744,N_16621);
nor U16939 (N_16939,N_16732,N_16629);
and U16940 (N_16940,N_16736,N_16655);
nor U16941 (N_16941,N_16614,N_16738);
nor U16942 (N_16942,N_16640,N_16678);
or U16943 (N_16943,N_16763,N_16715);
and U16944 (N_16944,N_16701,N_16649);
nor U16945 (N_16945,N_16625,N_16644);
nor U16946 (N_16946,N_16668,N_16761);
nand U16947 (N_16947,N_16721,N_16616);
nor U16948 (N_16948,N_16799,N_16753);
nor U16949 (N_16949,N_16600,N_16682);
nand U16950 (N_16950,N_16779,N_16749);
nand U16951 (N_16951,N_16752,N_16732);
nand U16952 (N_16952,N_16637,N_16770);
nand U16953 (N_16953,N_16630,N_16764);
nand U16954 (N_16954,N_16629,N_16659);
or U16955 (N_16955,N_16636,N_16676);
nand U16956 (N_16956,N_16657,N_16642);
nand U16957 (N_16957,N_16791,N_16683);
nand U16958 (N_16958,N_16644,N_16714);
or U16959 (N_16959,N_16630,N_16788);
or U16960 (N_16960,N_16678,N_16661);
and U16961 (N_16961,N_16681,N_16794);
nor U16962 (N_16962,N_16678,N_16680);
nor U16963 (N_16963,N_16725,N_16693);
nor U16964 (N_16964,N_16780,N_16778);
nand U16965 (N_16965,N_16644,N_16662);
nand U16966 (N_16966,N_16637,N_16697);
or U16967 (N_16967,N_16697,N_16600);
or U16968 (N_16968,N_16633,N_16786);
nor U16969 (N_16969,N_16625,N_16705);
and U16970 (N_16970,N_16795,N_16615);
xnor U16971 (N_16971,N_16717,N_16676);
xnor U16972 (N_16972,N_16777,N_16750);
and U16973 (N_16973,N_16701,N_16683);
or U16974 (N_16974,N_16623,N_16746);
and U16975 (N_16975,N_16797,N_16733);
nand U16976 (N_16976,N_16783,N_16743);
nand U16977 (N_16977,N_16629,N_16735);
nor U16978 (N_16978,N_16692,N_16705);
or U16979 (N_16979,N_16679,N_16768);
and U16980 (N_16980,N_16613,N_16792);
nor U16981 (N_16981,N_16720,N_16660);
and U16982 (N_16982,N_16718,N_16654);
or U16983 (N_16983,N_16642,N_16785);
nand U16984 (N_16984,N_16659,N_16780);
and U16985 (N_16985,N_16798,N_16611);
or U16986 (N_16986,N_16751,N_16650);
nand U16987 (N_16987,N_16749,N_16714);
nor U16988 (N_16988,N_16677,N_16780);
or U16989 (N_16989,N_16638,N_16727);
nor U16990 (N_16990,N_16774,N_16664);
or U16991 (N_16991,N_16617,N_16731);
nor U16992 (N_16992,N_16647,N_16782);
nor U16993 (N_16993,N_16744,N_16742);
nand U16994 (N_16994,N_16602,N_16614);
nor U16995 (N_16995,N_16602,N_16744);
nand U16996 (N_16996,N_16647,N_16625);
or U16997 (N_16997,N_16772,N_16760);
or U16998 (N_16998,N_16700,N_16614);
nand U16999 (N_16999,N_16765,N_16720);
and U17000 (N_17000,N_16825,N_16979);
nand U17001 (N_17001,N_16859,N_16951);
and U17002 (N_17002,N_16891,N_16923);
nor U17003 (N_17003,N_16878,N_16896);
nor U17004 (N_17004,N_16901,N_16986);
and U17005 (N_17005,N_16948,N_16937);
and U17006 (N_17006,N_16930,N_16968);
or U17007 (N_17007,N_16829,N_16884);
or U17008 (N_17008,N_16964,N_16972);
or U17009 (N_17009,N_16864,N_16992);
and U17010 (N_17010,N_16830,N_16836);
and U17011 (N_17011,N_16820,N_16848);
nand U17012 (N_17012,N_16908,N_16926);
and U17013 (N_17013,N_16969,N_16854);
and U17014 (N_17014,N_16892,N_16952);
nand U17015 (N_17015,N_16936,N_16802);
or U17016 (N_17016,N_16987,N_16880);
and U17017 (N_17017,N_16837,N_16982);
and U17018 (N_17018,N_16897,N_16839);
nor U17019 (N_17019,N_16819,N_16996);
nor U17020 (N_17020,N_16920,N_16960);
or U17021 (N_17021,N_16882,N_16985);
nor U17022 (N_17022,N_16955,N_16902);
or U17023 (N_17023,N_16959,N_16803);
or U17024 (N_17024,N_16919,N_16885);
nand U17025 (N_17025,N_16856,N_16989);
nand U17026 (N_17026,N_16965,N_16924);
or U17027 (N_17027,N_16838,N_16917);
and U17028 (N_17028,N_16872,N_16971);
or U17029 (N_17029,N_16970,N_16912);
and U17030 (N_17030,N_16842,N_16811);
and U17031 (N_17031,N_16858,N_16801);
nand U17032 (N_17032,N_16906,N_16805);
and U17033 (N_17033,N_16871,N_16868);
and U17034 (N_17034,N_16949,N_16940);
nor U17035 (N_17035,N_16980,N_16904);
and U17036 (N_17036,N_16832,N_16874);
or U17037 (N_17037,N_16945,N_16883);
or U17038 (N_17038,N_16913,N_16855);
or U17039 (N_17039,N_16821,N_16953);
or U17040 (N_17040,N_16810,N_16943);
or U17041 (N_17041,N_16983,N_16835);
nor U17042 (N_17042,N_16990,N_16950);
and U17043 (N_17043,N_16978,N_16976);
nor U17044 (N_17044,N_16927,N_16847);
nor U17045 (N_17045,N_16881,N_16998);
nand U17046 (N_17046,N_16922,N_16935);
nor U17047 (N_17047,N_16999,N_16806);
nor U17048 (N_17048,N_16932,N_16958);
nand U17049 (N_17049,N_16929,N_16939);
nand U17050 (N_17050,N_16963,N_16911);
and U17051 (N_17051,N_16962,N_16840);
nor U17052 (N_17052,N_16894,N_16817);
or U17053 (N_17053,N_16934,N_16826);
nor U17054 (N_17054,N_16933,N_16841);
nand U17055 (N_17055,N_16869,N_16899);
nand U17056 (N_17056,N_16852,N_16898);
and U17057 (N_17057,N_16947,N_16991);
nand U17058 (N_17058,N_16857,N_16866);
and U17059 (N_17059,N_16824,N_16822);
nor U17060 (N_17060,N_16966,N_16977);
or U17061 (N_17061,N_16893,N_16946);
nand U17062 (N_17062,N_16827,N_16834);
and U17063 (N_17063,N_16918,N_16915);
nor U17064 (N_17064,N_16916,N_16823);
or U17065 (N_17065,N_16890,N_16907);
or U17066 (N_17066,N_16800,N_16921);
or U17067 (N_17067,N_16804,N_16875);
and U17068 (N_17068,N_16867,N_16815);
nor U17069 (N_17069,N_16863,N_16938);
nor U17070 (N_17070,N_16961,N_16931);
and U17071 (N_17071,N_16895,N_16993);
or U17072 (N_17072,N_16853,N_16809);
nand U17073 (N_17073,N_16944,N_16808);
and U17074 (N_17074,N_16900,N_16861);
nor U17075 (N_17075,N_16974,N_16957);
nand U17076 (N_17076,N_16879,N_16846);
nor U17077 (N_17077,N_16851,N_16975);
or U17078 (N_17078,N_16984,N_16967);
and U17079 (N_17079,N_16903,N_16850);
nand U17080 (N_17080,N_16865,N_16941);
and U17081 (N_17081,N_16860,N_16997);
or U17082 (N_17082,N_16887,N_16844);
or U17083 (N_17083,N_16845,N_16988);
nor U17084 (N_17084,N_16813,N_16910);
nor U17085 (N_17085,N_16814,N_16942);
or U17086 (N_17086,N_16973,N_16995);
nor U17087 (N_17087,N_16956,N_16849);
nor U17088 (N_17088,N_16981,N_16876);
nor U17089 (N_17089,N_16873,N_16828);
nor U17090 (N_17090,N_16870,N_16816);
and U17091 (N_17091,N_16807,N_16877);
and U17092 (N_17092,N_16889,N_16833);
nand U17093 (N_17093,N_16812,N_16928);
or U17094 (N_17094,N_16914,N_16909);
nor U17095 (N_17095,N_16886,N_16888);
nand U17096 (N_17096,N_16905,N_16862);
and U17097 (N_17097,N_16994,N_16954);
and U17098 (N_17098,N_16818,N_16831);
and U17099 (N_17099,N_16843,N_16925);
nand U17100 (N_17100,N_16933,N_16983);
and U17101 (N_17101,N_16985,N_16999);
nor U17102 (N_17102,N_16831,N_16976);
or U17103 (N_17103,N_16926,N_16956);
or U17104 (N_17104,N_16969,N_16861);
and U17105 (N_17105,N_16908,N_16852);
nor U17106 (N_17106,N_16887,N_16817);
and U17107 (N_17107,N_16863,N_16850);
and U17108 (N_17108,N_16829,N_16862);
or U17109 (N_17109,N_16967,N_16845);
or U17110 (N_17110,N_16977,N_16848);
nand U17111 (N_17111,N_16957,N_16893);
and U17112 (N_17112,N_16982,N_16933);
nor U17113 (N_17113,N_16923,N_16948);
or U17114 (N_17114,N_16983,N_16976);
nor U17115 (N_17115,N_16945,N_16906);
or U17116 (N_17116,N_16977,N_16897);
or U17117 (N_17117,N_16974,N_16832);
or U17118 (N_17118,N_16841,N_16953);
or U17119 (N_17119,N_16902,N_16982);
and U17120 (N_17120,N_16917,N_16921);
nor U17121 (N_17121,N_16975,N_16904);
nand U17122 (N_17122,N_16868,N_16982);
and U17123 (N_17123,N_16829,N_16899);
nor U17124 (N_17124,N_16992,N_16941);
and U17125 (N_17125,N_16986,N_16900);
and U17126 (N_17126,N_16968,N_16815);
and U17127 (N_17127,N_16999,N_16902);
nor U17128 (N_17128,N_16942,N_16972);
and U17129 (N_17129,N_16979,N_16888);
and U17130 (N_17130,N_16881,N_16859);
nand U17131 (N_17131,N_16868,N_16859);
nor U17132 (N_17132,N_16944,N_16914);
or U17133 (N_17133,N_16830,N_16813);
nand U17134 (N_17134,N_16938,N_16866);
nand U17135 (N_17135,N_16907,N_16811);
nor U17136 (N_17136,N_16981,N_16824);
or U17137 (N_17137,N_16945,N_16828);
or U17138 (N_17138,N_16914,N_16902);
xnor U17139 (N_17139,N_16834,N_16948);
nand U17140 (N_17140,N_16806,N_16915);
nand U17141 (N_17141,N_16894,N_16939);
and U17142 (N_17142,N_16807,N_16963);
nand U17143 (N_17143,N_16960,N_16825);
nand U17144 (N_17144,N_16811,N_16883);
nand U17145 (N_17145,N_16924,N_16858);
or U17146 (N_17146,N_16839,N_16833);
or U17147 (N_17147,N_16910,N_16950);
or U17148 (N_17148,N_16944,N_16953);
and U17149 (N_17149,N_16860,N_16993);
nor U17150 (N_17150,N_16959,N_16882);
nor U17151 (N_17151,N_16954,N_16909);
or U17152 (N_17152,N_16885,N_16894);
and U17153 (N_17153,N_16908,N_16992);
and U17154 (N_17154,N_16907,N_16985);
or U17155 (N_17155,N_16803,N_16899);
nand U17156 (N_17156,N_16886,N_16833);
and U17157 (N_17157,N_16996,N_16849);
or U17158 (N_17158,N_16844,N_16824);
nor U17159 (N_17159,N_16987,N_16925);
nand U17160 (N_17160,N_16992,N_16965);
nor U17161 (N_17161,N_16997,N_16835);
or U17162 (N_17162,N_16854,N_16966);
nand U17163 (N_17163,N_16934,N_16808);
nand U17164 (N_17164,N_16960,N_16837);
or U17165 (N_17165,N_16989,N_16840);
and U17166 (N_17166,N_16828,N_16940);
nand U17167 (N_17167,N_16836,N_16853);
or U17168 (N_17168,N_16812,N_16904);
and U17169 (N_17169,N_16831,N_16907);
nor U17170 (N_17170,N_16977,N_16819);
nand U17171 (N_17171,N_16874,N_16991);
nand U17172 (N_17172,N_16919,N_16832);
nor U17173 (N_17173,N_16989,N_16806);
and U17174 (N_17174,N_16841,N_16970);
nand U17175 (N_17175,N_16891,N_16996);
nor U17176 (N_17176,N_16924,N_16854);
nor U17177 (N_17177,N_16890,N_16934);
nand U17178 (N_17178,N_16963,N_16927);
nor U17179 (N_17179,N_16841,N_16891);
and U17180 (N_17180,N_16874,N_16906);
and U17181 (N_17181,N_16987,N_16899);
or U17182 (N_17182,N_16885,N_16828);
or U17183 (N_17183,N_16890,N_16872);
or U17184 (N_17184,N_16948,N_16947);
nand U17185 (N_17185,N_16831,N_16990);
nand U17186 (N_17186,N_16838,N_16898);
or U17187 (N_17187,N_16859,N_16821);
and U17188 (N_17188,N_16992,N_16820);
and U17189 (N_17189,N_16872,N_16981);
nand U17190 (N_17190,N_16924,N_16876);
nand U17191 (N_17191,N_16975,N_16861);
nand U17192 (N_17192,N_16894,N_16830);
nand U17193 (N_17193,N_16830,N_16837);
or U17194 (N_17194,N_16943,N_16959);
or U17195 (N_17195,N_16984,N_16994);
nor U17196 (N_17196,N_16800,N_16920);
and U17197 (N_17197,N_16809,N_16907);
or U17198 (N_17198,N_16867,N_16977);
nand U17199 (N_17199,N_16963,N_16817);
nand U17200 (N_17200,N_17137,N_17072);
nand U17201 (N_17201,N_17025,N_17195);
or U17202 (N_17202,N_17041,N_17058);
or U17203 (N_17203,N_17177,N_17009);
and U17204 (N_17204,N_17158,N_17198);
nand U17205 (N_17205,N_17044,N_17069);
nor U17206 (N_17206,N_17075,N_17095);
nand U17207 (N_17207,N_17164,N_17138);
nor U17208 (N_17208,N_17085,N_17123);
nand U17209 (N_17209,N_17030,N_17124);
or U17210 (N_17210,N_17129,N_17066);
nand U17211 (N_17211,N_17067,N_17178);
or U17212 (N_17212,N_17079,N_17115);
and U17213 (N_17213,N_17096,N_17100);
nor U17214 (N_17214,N_17188,N_17084);
and U17215 (N_17215,N_17043,N_17063);
nand U17216 (N_17216,N_17078,N_17003);
or U17217 (N_17217,N_17135,N_17150);
and U17218 (N_17218,N_17119,N_17033);
nand U17219 (N_17219,N_17017,N_17056);
nand U17220 (N_17220,N_17167,N_17073);
and U17221 (N_17221,N_17128,N_17105);
or U17222 (N_17222,N_17184,N_17130);
xor U17223 (N_17223,N_17170,N_17189);
or U17224 (N_17224,N_17097,N_17016);
nor U17225 (N_17225,N_17042,N_17051);
nand U17226 (N_17226,N_17156,N_17081);
nor U17227 (N_17227,N_17102,N_17133);
and U17228 (N_17228,N_17000,N_17020);
and U17229 (N_17229,N_17109,N_17174);
or U17230 (N_17230,N_17197,N_17054);
nor U17231 (N_17231,N_17172,N_17110);
nor U17232 (N_17232,N_17179,N_17099);
or U17233 (N_17233,N_17152,N_17071);
nand U17234 (N_17234,N_17168,N_17139);
nand U17235 (N_17235,N_17131,N_17015);
or U17236 (N_17236,N_17117,N_17059);
nor U17237 (N_17237,N_17161,N_17103);
nand U17238 (N_17238,N_17022,N_17087);
nand U17239 (N_17239,N_17140,N_17021);
and U17240 (N_17240,N_17194,N_17154);
nor U17241 (N_17241,N_17112,N_17053);
and U17242 (N_17242,N_17040,N_17171);
nor U17243 (N_17243,N_17036,N_17065);
and U17244 (N_17244,N_17091,N_17035);
or U17245 (N_17245,N_17104,N_17088);
nor U17246 (N_17246,N_17077,N_17142);
nand U17247 (N_17247,N_17143,N_17049);
or U17248 (N_17248,N_17196,N_17175);
or U17249 (N_17249,N_17173,N_17181);
nand U17250 (N_17250,N_17055,N_17192);
and U17251 (N_17251,N_17098,N_17176);
nand U17252 (N_17252,N_17070,N_17114);
nor U17253 (N_17253,N_17028,N_17111);
and U17254 (N_17254,N_17068,N_17180);
or U17255 (N_17255,N_17061,N_17151);
nand U17256 (N_17256,N_17132,N_17144);
nand U17257 (N_17257,N_17048,N_17157);
and U17258 (N_17258,N_17018,N_17107);
or U17259 (N_17259,N_17034,N_17193);
and U17260 (N_17260,N_17094,N_17012);
and U17261 (N_17261,N_17001,N_17046);
nand U17262 (N_17262,N_17011,N_17076);
nor U17263 (N_17263,N_17038,N_17106);
nand U17264 (N_17264,N_17019,N_17023);
and U17265 (N_17265,N_17125,N_17013);
or U17266 (N_17266,N_17005,N_17024);
nand U17267 (N_17267,N_17080,N_17136);
and U17268 (N_17268,N_17010,N_17008);
or U17269 (N_17269,N_17047,N_17146);
nand U17270 (N_17270,N_17182,N_17045);
and U17271 (N_17271,N_17050,N_17183);
and U17272 (N_17272,N_17090,N_17014);
and U17273 (N_17273,N_17166,N_17163);
nand U17274 (N_17274,N_17052,N_17169);
nand U17275 (N_17275,N_17064,N_17153);
nor U17276 (N_17276,N_17002,N_17083);
nand U17277 (N_17277,N_17149,N_17093);
and U17278 (N_17278,N_17108,N_17089);
and U17279 (N_17279,N_17147,N_17101);
nand U17280 (N_17280,N_17039,N_17155);
and U17281 (N_17281,N_17007,N_17145);
nand U17282 (N_17282,N_17118,N_17159);
nor U17283 (N_17283,N_17127,N_17092);
nor U17284 (N_17284,N_17057,N_17160);
nor U17285 (N_17285,N_17191,N_17031);
and U17286 (N_17286,N_17006,N_17148);
nand U17287 (N_17287,N_17165,N_17190);
or U17288 (N_17288,N_17037,N_17162);
nor U17289 (N_17289,N_17062,N_17027);
xnor U17290 (N_17290,N_17026,N_17186);
nor U17291 (N_17291,N_17126,N_17120);
and U17292 (N_17292,N_17199,N_17187);
nor U17293 (N_17293,N_17086,N_17060);
or U17294 (N_17294,N_17141,N_17074);
or U17295 (N_17295,N_17113,N_17134);
or U17296 (N_17296,N_17004,N_17082);
nor U17297 (N_17297,N_17121,N_17116);
nand U17298 (N_17298,N_17032,N_17122);
or U17299 (N_17299,N_17029,N_17185);
nand U17300 (N_17300,N_17174,N_17099);
nor U17301 (N_17301,N_17103,N_17092);
nor U17302 (N_17302,N_17153,N_17089);
nor U17303 (N_17303,N_17066,N_17162);
and U17304 (N_17304,N_17012,N_17161);
nand U17305 (N_17305,N_17181,N_17009);
xnor U17306 (N_17306,N_17178,N_17077);
or U17307 (N_17307,N_17004,N_17042);
or U17308 (N_17308,N_17141,N_17034);
and U17309 (N_17309,N_17064,N_17034);
nor U17310 (N_17310,N_17123,N_17178);
or U17311 (N_17311,N_17176,N_17050);
or U17312 (N_17312,N_17062,N_17176);
or U17313 (N_17313,N_17022,N_17084);
or U17314 (N_17314,N_17198,N_17103);
nor U17315 (N_17315,N_17001,N_17192);
or U17316 (N_17316,N_17152,N_17002);
or U17317 (N_17317,N_17123,N_17042);
xor U17318 (N_17318,N_17032,N_17031);
xnor U17319 (N_17319,N_17082,N_17021);
or U17320 (N_17320,N_17194,N_17119);
nor U17321 (N_17321,N_17145,N_17198);
and U17322 (N_17322,N_17072,N_17183);
and U17323 (N_17323,N_17170,N_17043);
nand U17324 (N_17324,N_17186,N_17192);
nor U17325 (N_17325,N_17056,N_17023);
nor U17326 (N_17326,N_17113,N_17174);
and U17327 (N_17327,N_17141,N_17189);
nand U17328 (N_17328,N_17059,N_17128);
nand U17329 (N_17329,N_17015,N_17136);
and U17330 (N_17330,N_17140,N_17180);
nor U17331 (N_17331,N_17033,N_17120);
nand U17332 (N_17332,N_17076,N_17110);
nor U17333 (N_17333,N_17026,N_17122);
and U17334 (N_17334,N_17163,N_17149);
nor U17335 (N_17335,N_17093,N_17160);
or U17336 (N_17336,N_17077,N_17088);
nand U17337 (N_17337,N_17096,N_17174);
nor U17338 (N_17338,N_17093,N_17186);
or U17339 (N_17339,N_17061,N_17114);
and U17340 (N_17340,N_17186,N_17131);
or U17341 (N_17341,N_17149,N_17058);
nor U17342 (N_17342,N_17017,N_17111);
and U17343 (N_17343,N_17198,N_17063);
and U17344 (N_17344,N_17189,N_17198);
and U17345 (N_17345,N_17154,N_17076);
nand U17346 (N_17346,N_17106,N_17137);
and U17347 (N_17347,N_17191,N_17121);
nor U17348 (N_17348,N_17004,N_17011);
nand U17349 (N_17349,N_17111,N_17112);
nand U17350 (N_17350,N_17138,N_17042);
nor U17351 (N_17351,N_17063,N_17010);
or U17352 (N_17352,N_17195,N_17173);
nand U17353 (N_17353,N_17033,N_17173);
nand U17354 (N_17354,N_17119,N_17036);
or U17355 (N_17355,N_17192,N_17167);
nor U17356 (N_17356,N_17082,N_17068);
or U17357 (N_17357,N_17173,N_17101);
or U17358 (N_17358,N_17113,N_17101);
or U17359 (N_17359,N_17182,N_17137);
and U17360 (N_17360,N_17020,N_17172);
nor U17361 (N_17361,N_17067,N_17014);
and U17362 (N_17362,N_17095,N_17190);
nand U17363 (N_17363,N_17048,N_17099);
and U17364 (N_17364,N_17082,N_17131);
nand U17365 (N_17365,N_17094,N_17088);
nand U17366 (N_17366,N_17195,N_17162);
and U17367 (N_17367,N_17170,N_17132);
nand U17368 (N_17368,N_17181,N_17000);
nor U17369 (N_17369,N_17099,N_17082);
or U17370 (N_17370,N_17189,N_17042);
and U17371 (N_17371,N_17056,N_17184);
or U17372 (N_17372,N_17184,N_17058);
and U17373 (N_17373,N_17180,N_17147);
nor U17374 (N_17374,N_17026,N_17015);
nand U17375 (N_17375,N_17013,N_17133);
nand U17376 (N_17376,N_17100,N_17090);
and U17377 (N_17377,N_17088,N_17175);
and U17378 (N_17378,N_17143,N_17009);
nand U17379 (N_17379,N_17061,N_17144);
or U17380 (N_17380,N_17029,N_17159);
or U17381 (N_17381,N_17175,N_17039);
or U17382 (N_17382,N_17155,N_17152);
nand U17383 (N_17383,N_17006,N_17152);
or U17384 (N_17384,N_17056,N_17198);
or U17385 (N_17385,N_17132,N_17031);
nand U17386 (N_17386,N_17191,N_17195);
xnor U17387 (N_17387,N_17017,N_17049);
nand U17388 (N_17388,N_17038,N_17064);
and U17389 (N_17389,N_17049,N_17046);
and U17390 (N_17390,N_17172,N_17124);
nand U17391 (N_17391,N_17036,N_17146);
or U17392 (N_17392,N_17089,N_17055);
nor U17393 (N_17393,N_17098,N_17140);
or U17394 (N_17394,N_17153,N_17018);
and U17395 (N_17395,N_17043,N_17078);
nand U17396 (N_17396,N_17108,N_17078);
or U17397 (N_17397,N_17000,N_17141);
and U17398 (N_17398,N_17137,N_17162);
nand U17399 (N_17399,N_17179,N_17023);
or U17400 (N_17400,N_17394,N_17273);
and U17401 (N_17401,N_17265,N_17278);
and U17402 (N_17402,N_17242,N_17294);
nor U17403 (N_17403,N_17210,N_17279);
and U17404 (N_17404,N_17285,N_17385);
and U17405 (N_17405,N_17244,N_17295);
and U17406 (N_17406,N_17274,N_17299);
or U17407 (N_17407,N_17374,N_17358);
nor U17408 (N_17408,N_17328,N_17325);
or U17409 (N_17409,N_17236,N_17340);
nand U17410 (N_17410,N_17221,N_17308);
or U17411 (N_17411,N_17332,N_17360);
nand U17412 (N_17412,N_17338,N_17241);
nor U17413 (N_17413,N_17219,N_17288);
nand U17414 (N_17414,N_17268,N_17378);
or U17415 (N_17415,N_17380,N_17264);
nor U17416 (N_17416,N_17346,N_17209);
and U17417 (N_17417,N_17387,N_17257);
or U17418 (N_17418,N_17375,N_17314);
or U17419 (N_17419,N_17362,N_17321);
and U17420 (N_17420,N_17329,N_17370);
nand U17421 (N_17421,N_17275,N_17245);
or U17422 (N_17422,N_17345,N_17309);
nor U17423 (N_17423,N_17343,N_17291);
or U17424 (N_17424,N_17276,N_17371);
and U17425 (N_17425,N_17263,N_17304);
nand U17426 (N_17426,N_17390,N_17366);
and U17427 (N_17427,N_17364,N_17280);
xor U17428 (N_17428,N_17222,N_17311);
or U17429 (N_17429,N_17317,N_17218);
nor U17430 (N_17430,N_17213,N_17373);
or U17431 (N_17431,N_17206,N_17339);
or U17432 (N_17432,N_17204,N_17305);
nand U17433 (N_17433,N_17212,N_17356);
or U17434 (N_17434,N_17246,N_17201);
or U17435 (N_17435,N_17324,N_17367);
or U17436 (N_17436,N_17251,N_17256);
and U17437 (N_17437,N_17389,N_17232);
and U17438 (N_17438,N_17271,N_17262);
nand U17439 (N_17439,N_17365,N_17319);
and U17440 (N_17440,N_17253,N_17301);
or U17441 (N_17441,N_17298,N_17216);
nor U17442 (N_17442,N_17229,N_17352);
nand U17443 (N_17443,N_17377,N_17284);
nand U17444 (N_17444,N_17272,N_17368);
nor U17445 (N_17445,N_17238,N_17335);
and U17446 (N_17446,N_17392,N_17283);
and U17447 (N_17447,N_17363,N_17330);
or U17448 (N_17448,N_17289,N_17313);
or U17449 (N_17449,N_17361,N_17228);
and U17450 (N_17450,N_17255,N_17217);
or U17451 (N_17451,N_17297,N_17260);
and U17452 (N_17452,N_17281,N_17296);
nor U17453 (N_17453,N_17359,N_17302);
or U17454 (N_17454,N_17220,N_17331);
nor U17455 (N_17455,N_17259,N_17351);
nor U17456 (N_17456,N_17282,N_17243);
and U17457 (N_17457,N_17290,N_17249);
and U17458 (N_17458,N_17261,N_17292);
or U17459 (N_17459,N_17396,N_17323);
nand U17460 (N_17460,N_17269,N_17258);
nand U17461 (N_17461,N_17334,N_17333);
nor U17462 (N_17462,N_17205,N_17235);
nor U17463 (N_17463,N_17266,N_17207);
nand U17464 (N_17464,N_17254,N_17208);
and U17465 (N_17465,N_17307,N_17315);
nor U17466 (N_17466,N_17395,N_17318);
or U17467 (N_17467,N_17383,N_17386);
nor U17468 (N_17468,N_17234,N_17239);
and U17469 (N_17469,N_17225,N_17200);
nand U17470 (N_17470,N_17341,N_17376);
and U17471 (N_17471,N_17286,N_17350);
nand U17472 (N_17472,N_17336,N_17349);
nand U17473 (N_17473,N_17300,N_17379);
or U17474 (N_17474,N_17337,N_17252);
or U17475 (N_17475,N_17287,N_17316);
or U17476 (N_17476,N_17381,N_17202);
and U17477 (N_17477,N_17270,N_17224);
and U17478 (N_17478,N_17354,N_17306);
nand U17479 (N_17479,N_17215,N_17326);
and U17480 (N_17480,N_17397,N_17230);
or U17481 (N_17481,N_17382,N_17247);
nand U17482 (N_17482,N_17322,N_17203);
and U17483 (N_17483,N_17293,N_17357);
nand U17484 (N_17484,N_17227,N_17353);
or U17485 (N_17485,N_17231,N_17384);
nand U17486 (N_17486,N_17369,N_17399);
nor U17487 (N_17487,N_17327,N_17372);
and U17488 (N_17488,N_17226,N_17355);
and U17489 (N_17489,N_17233,N_17248);
nor U17490 (N_17490,N_17237,N_17310);
and U17491 (N_17491,N_17342,N_17240);
or U17492 (N_17492,N_17344,N_17223);
nand U17493 (N_17493,N_17277,N_17214);
nand U17494 (N_17494,N_17303,N_17393);
nor U17495 (N_17495,N_17388,N_17398);
nor U17496 (N_17496,N_17267,N_17250);
or U17497 (N_17497,N_17211,N_17348);
nand U17498 (N_17498,N_17391,N_17347);
and U17499 (N_17499,N_17320,N_17312);
nor U17500 (N_17500,N_17283,N_17296);
and U17501 (N_17501,N_17209,N_17321);
and U17502 (N_17502,N_17292,N_17284);
nand U17503 (N_17503,N_17281,N_17223);
nand U17504 (N_17504,N_17371,N_17334);
nor U17505 (N_17505,N_17299,N_17204);
nand U17506 (N_17506,N_17374,N_17214);
nand U17507 (N_17507,N_17275,N_17398);
and U17508 (N_17508,N_17254,N_17288);
nor U17509 (N_17509,N_17281,N_17381);
nor U17510 (N_17510,N_17282,N_17238);
or U17511 (N_17511,N_17386,N_17225);
and U17512 (N_17512,N_17377,N_17311);
xor U17513 (N_17513,N_17296,N_17309);
and U17514 (N_17514,N_17257,N_17373);
or U17515 (N_17515,N_17368,N_17256);
nor U17516 (N_17516,N_17267,N_17218);
and U17517 (N_17517,N_17336,N_17297);
and U17518 (N_17518,N_17365,N_17377);
nand U17519 (N_17519,N_17394,N_17250);
or U17520 (N_17520,N_17353,N_17376);
and U17521 (N_17521,N_17279,N_17306);
nor U17522 (N_17522,N_17294,N_17286);
or U17523 (N_17523,N_17284,N_17205);
nor U17524 (N_17524,N_17293,N_17369);
nor U17525 (N_17525,N_17386,N_17259);
nor U17526 (N_17526,N_17398,N_17316);
nor U17527 (N_17527,N_17261,N_17273);
nand U17528 (N_17528,N_17349,N_17316);
nand U17529 (N_17529,N_17396,N_17293);
nor U17530 (N_17530,N_17344,N_17290);
nor U17531 (N_17531,N_17298,N_17274);
nor U17532 (N_17532,N_17249,N_17225);
and U17533 (N_17533,N_17213,N_17244);
nand U17534 (N_17534,N_17312,N_17245);
or U17535 (N_17535,N_17246,N_17290);
nor U17536 (N_17536,N_17392,N_17242);
nor U17537 (N_17537,N_17285,N_17223);
or U17538 (N_17538,N_17302,N_17239);
nor U17539 (N_17539,N_17280,N_17398);
and U17540 (N_17540,N_17372,N_17203);
or U17541 (N_17541,N_17271,N_17290);
nor U17542 (N_17542,N_17279,N_17264);
nor U17543 (N_17543,N_17386,N_17267);
nand U17544 (N_17544,N_17317,N_17248);
nor U17545 (N_17545,N_17318,N_17282);
or U17546 (N_17546,N_17355,N_17245);
nand U17547 (N_17547,N_17249,N_17315);
nor U17548 (N_17548,N_17351,N_17330);
nor U17549 (N_17549,N_17226,N_17396);
nor U17550 (N_17550,N_17273,N_17212);
nand U17551 (N_17551,N_17239,N_17350);
nand U17552 (N_17552,N_17272,N_17227);
nor U17553 (N_17553,N_17296,N_17354);
nor U17554 (N_17554,N_17318,N_17379);
nand U17555 (N_17555,N_17357,N_17200);
and U17556 (N_17556,N_17353,N_17270);
or U17557 (N_17557,N_17371,N_17222);
nand U17558 (N_17558,N_17289,N_17367);
nand U17559 (N_17559,N_17250,N_17290);
or U17560 (N_17560,N_17394,N_17229);
and U17561 (N_17561,N_17205,N_17273);
nor U17562 (N_17562,N_17306,N_17242);
and U17563 (N_17563,N_17256,N_17229);
nor U17564 (N_17564,N_17311,N_17247);
and U17565 (N_17565,N_17249,N_17324);
nand U17566 (N_17566,N_17249,N_17376);
nor U17567 (N_17567,N_17374,N_17347);
and U17568 (N_17568,N_17220,N_17338);
or U17569 (N_17569,N_17230,N_17299);
nand U17570 (N_17570,N_17333,N_17232);
nand U17571 (N_17571,N_17257,N_17380);
nor U17572 (N_17572,N_17335,N_17241);
nor U17573 (N_17573,N_17236,N_17358);
or U17574 (N_17574,N_17307,N_17254);
or U17575 (N_17575,N_17256,N_17283);
or U17576 (N_17576,N_17382,N_17376);
or U17577 (N_17577,N_17320,N_17330);
nand U17578 (N_17578,N_17208,N_17354);
nor U17579 (N_17579,N_17396,N_17299);
nor U17580 (N_17580,N_17229,N_17330);
and U17581 (N_17581,N_17374,N_17328);
nand U17582 (N_17582,N_17287,N_17293);
and U17583 (N_17583,N_17352,N_17204);
and U17584 (N_17584,N_17246,N_17226);
and U17585 (N_17585,N_17262,N_17393);
or U17586 (N_17586,N_17248,N_17360);
and U17587 (N_17587,N_17249,N_17346);
or U17588 (N_17588,N_17339,N_17306);
and U17589 (N_17589,N_17374,N_17327);
and U17590 (N_17590,N_17367,N_17341);
or U17591 (N_17591,N_17252,N_17242);
and U17592 (N_17592,N_17204,N_17302);
and U17593 (N_17593,N_17230,N_17343);
nand U17594 (N_17594,N_17310,N_17313);
or U17595 (N_17595,N_17397,N_17357);
or U17596 (N_17596,N_17369,N_17253);
and U17597 (N_17597,N_17273,N_17383);
nor U17598 (N_17598,N_17383,N_17323);
xnor U17599 (N_17599,N_17321,N_17258);
and U17600 (N_17600,N_17451,N_17490);
nor U17601 (N_17601,N_17592,N_17468);
or U17602 (N_17602,N_17542,N_17403);
nor U17603 (N_17603,N_17462,N_17552);
nand U17604 (N_17604,N_17424,N_17534);
nand U17605 (N_17605,N_17455,N_17537);
or U17606 (N_17606,N_17476,N_17503);
and U17607 (N_17607,N_17442,N_17544);
nor U17608 (N_17608,N_17591,N_17461);
or U17609 (N_17609,N_17555,N_17443);
and U17610 (N_17610,N_17524,N_17530);
and U17611 (N_17611,N_17449,N_17519);
and U17612 (N_17612,N_17472,N_17501);
and U17613 (N_17613,N_17431,N_17597);
and U17614 (N_17614,N_17415,N_17568);
nor U17615 (N_17615,N_17488,N_17412);
and U17616 (N_17616,N_17531,N_17535);
or U17617 (N_17617,N_17527,N_17520);
or U17618 (N_17618,N_17480,N_17594);
and U17619 (N_17619,N_17439,N_17562);
and U17620 (N_17620,N_17507,N_17511);
and U17621 (N_17621,N_17450,N_17598);
nor U17622 (N_17622,N_17437,N_17474);
or U17623 (N_17623,N_17436,N_17538);
and U17624 (N_17624,N_17465,N_17486);
nand U17625 (N_17625,N_17583,N_17593);
or U17626 (N_17626,N_17543,N_17540);
or U17627 (N_17627,N_17475,N_17549);
nand U17628 (N_17628,N_17518,N_17588);
nand U17629 (N_17629,N_17419,N_17584);
nor U17630 (N_17630,N_17509,N_17504);
and U17631 (N_17631,N_17513,N_17470);
nor U17632 (N_17632,N_17582,N_17407);
or U17633 (N_17633,N_17556,N_17590);
and U17634 (N_17634,N_17557,N_17495);
nand U17635 (N_17635,N_17473,N_17471);
nor U17636 (N_17636,N_17574,N_17550);
and U17637 (N_17637,N_17401,N_17454);
nor U17638 (N_17638,N_17510,N_17522);
nor U17639 (N_17639,N_17492,N_17571);
nor U17640 (N_17640,N_17573,N_17416);
nand U17641 (N_17641,N_17428,N_17400);
nor U17642 (N_17642,N_17498,N_17466);
or U17643 (N_17643,N_17438,N_17482);
nor U17644 (N_17644,N_17484,N_17560);
and U17645 (N_17645,N_17413,N_17599);
and U17646 (N_17646,N_17423,N_17499);
and U17647 (N_17647,N_17529,N_17577);
and U17648 (N_17648,N_17508,N_17460);
and U17649 (N_17649,N_17506,N_17464);
and U17650 (N_17650,N_17414,N_17576);
and U17651 (N_17651,N_17585,N_17570);
and U17652 (N_17652,N_17487,N_17422);
and U17653 (N_17653,N_17533,N_17447);
nor U17654 (N_17654,N_17569,N_17528);
nor U17655 (N_17655,N_17558,N_17425);
nand U17656 (N_17656,N_17417,N_17467);
nand U17657 (N_17657,N_17581,N_17463);
or U17658 (N_17658,N_17502,N_17514);
nor U17659 (N_17659,N_17559,N_17516);
or U17660 (N_17660,N_17469,N_17493);
or U17661 (N_17661,N_17515,N_17408);
nor U17662 (N_17662,N_17435,N_17579);
nand U17663 (N_17663,N_17551,N_17446);
nor U17664 (N_17664,N_17572,N_17481);
nor U17665 (N_17665,N_17445,N_17405);
nand U17666 (N_17666,N_17477,N_17409);
or U17667 (N_17667,N_17526,N_17497);
nor U17668 (N_17668,N_17548,N_17406);
nand U17669 (N_17669,N_17404,N_17567);
xnor U17670 (N_17670,N_17561,N_17532);
and U17671 (N_17671,N_17433,N_17578);
or U17672 (N_17672,N_17411,N_17596);
and U17673 (N_17673,N_17586,N_17483);
and U17674 (N_17674,N_17410,N_17563);
xor U17675 (N_17675,N_17575,N_17491);
or U17676 (N_17676,N_17500,N_17517);
and U17677 (N_17677,N_17494,N_17547);
nand U17678 (N_17678,N_17536,N_17485);
nand U17679 (N_17679,N_17444,N_17565);
nor U17680 (N_17680,N_17521,N_17523);
or U17681 (N_17681,N_17505,N_17453);
nor U17682 (N_17682,N_17564,N_17420);
or U17683 (N_17683,N_17512,N_17459);
and U17684 (N_17684,N_17434,N_17427);
and U17685 (N_17685,N_17496,N_17589);
or U17686 (N_17686,N_17545,N_17489);
xnor U17687 (N_17687,N_17426,N_17458);
or U17688 (N_17688,N_17402,N_17566);
and U17689 (N_17689,N_17452,N_17580);
or U17690 (N_17690,N_17595,N_17441);
nand U17691 (N_17691,N_17418,N_17457);
and U17692 (N_17692,N_17456,N_17448);
and U17693 (N_17693,N_17430,N_17440);
or U17694 (N_17694,N_17553,N_17539);
or U17695 (N_17695,N_17429,N_17479);
or U17696 (N_17696,N_17587,N_17421);
or U17697 (N_17697,N_17546,N_17432);
nand U17698 (N_17698,N_17525,N_17541);
or U17699 (N_17699,N_17478,N_17554);
and U17700 (N_17700,N_17597,N_17429);
nand U17701 (N_17701,N_17485,N_17487);
nor U17702 (N_17702,N_17488,N_17439);
or U17703 (N_17703,N_17555,N_17532);
or U17704 (N_17704,N_17508,N_17472);
nor U17705 (N_17705,N_17416,N_17424);
nor U17706 (N_17706,N_17546,N_17482);
nand U17707 (N_17707,N_17548,N_17505);
nor U17708 (N_17708,N_17550,N_17583);
and U17709 (N_17709,N_17585,N_17466);
nor U17710 (N_17710,N_17469,N_17492);
nand U17711 (N_17711,N_17556,N_17526);
nand U17712 (N_17712,N_17497,N_17562);
nand U17713 (N_17713,N_17582,N_17589);
and U17714 (N_17714,N_17586,N_17421);
nand U17715 (N_17715,N_17515,N_17485);
or U17716 (N_17716,N_17401,N_17480);
and U17717 (N_17717,N_17552,N_17496);
nand U17718 (N_17718,N_17499,N_17539);
nor U17719 (N_17719,N_17544,N_17440);
and U17720 (N_17720,N_17502,N_17530);
xnor U17721 (N_17721,N_17499,N_17573);
or U17722 (N_17722,N_17473,N_17508);
and U17723 (N_17723,N_17407,N_17467);
or U17724 (N_17724,N_17489,N_17481);
nor U17725 (N_17725,N_17468,N_17521);
nor U17726 (N_17726,N_17409,N_17480);
nand U17727 (N_17727,N_17583,N_17406);
nand U17728 (N_17728,N_17585,N_17472);
or U17729 (N_17729,N_17404,N_17593);
or U17730 (N_17730,N_17508,N_17405);
nand U17731 (N_17731,N_17411,N_17563);
or U17732 (N_17732,N_17598,N_17481);
or U17733 (N_17733,N_17509,N_17478);
and U17734 (N_17734,N_17491,N_17542);
and U17735 (N_17735,N_17470,N_17558);
nor U17736 (N_17736,N_17510,N_17596);
nand U17737 (N_17737,N_17511,N_17530);
nor U17738 (N_17738,N_17485,N_17458);
or U17739 (N_17739,N_17568,N_17414);
and U17740 (N_17740,N_17516,N_17475);
and U17741 (N_17741,N_17525,N_17455);
or U17742 (N_17742,N_17594,N_17467);
or U17743 (N_17743,N_17488,N_17549);
nor U17744 (N_17744,N_17468,N_17429);
nand U17745 (N_17745,N_17583,N_17426);
nand U17746 (N_17746,N_17497,N_17423);
nand U17747 (N_17747,N_17571,N_17457);
nand U17748 (N_17748,N_17421,N_17519);
nand U17749 (N_17749,N_17451,N_17598);
nor U17750 (N_17750,N_17544,N_17430);
or U17751 (N_17751,N_17526,N_17440);
and U17752 (N_17752,N_17438,N_17409);
and U17753 (N_17753,N_17404,N_17497);
nand U17754 (N_17754,N_17410,N_17448);
and U17755 (N_17755,N_17549,N_17414);
nand U17756 (N_17756,N_17465,N_17434);
nor U17757 (N_17757,N_17535,N_17593);
nor U17758 (N_17758,N_17404,N_17599);
nand U17759 (N_17759,N_17453,N_17596);
and U17760 (N_17760,N_17410,N_17413);
or U17761 (N_17761,N_17537,N_17571);
and U17762 (N_17762,N_17491,N_17597);
nor U17763 (N_17763,N_17535,N_17465);
nand U17764 (N_17764,N_17471,N_17440);
and U17765 (N_17765,N_17494,N_17539);
nand U17766 (N_17766,N_17569,N_17426);
and U17767 (N_17767,N_17416,N_17510);
and U17768 (N_17768,N_17405,N_17433);
nand U17769 (N_17769,N_17509,N_17473);
or U17770 (N_17770,N_17516,N_17445);
nor U17771 (N_17771,N_17584,N_17430);
nand U17772 (N_17772,N_17498,N_17571);
and U17773 (N_17773,N_17598,N_17571);
or U17774 (N_17774,N_17587,N_17462);
xor U17775 (N_17775,N_17414,N_17459);
or U17776 (N_17776,N_17532,N_17504);
and U17777 (N_17777,N_17445,N_17442);
nand U17778 (N_17778,N_17471,N_17534);
nor U17779 (N_17779,N_17561,N_17413);
xnor U17780 (N_17780,N_17501,N_17552);
nand U17781 (N_17781,N_17556,N_17546);
nand U17782 (N_17782,N_17550,N_17467);
nand U17783 (N_17783,N_17419,N_17503);
nand U17784 (N_17784,N_17451,N_17478);
nand U17785 (N_17785,N_17495,N_17595);
nor U17786 (N_17786,N_17590,N_17559);
and U17787 (N_17787,N_17457,N_17480);
nor U17788 (N_17788,N_17512,N_17417);
nand U17789 (N_17789,N_17418,N_17508);
and U17790 (N_17790,N_17418,N_17522);
xnor U17791 (N_17791,N_17475,N_17436);
or U17792 (N_17792,N_17550,N_17507);
nand U17793 (N_17793,N_17404,N_17569);
and U17794 (N_17794,N_17513,N_17569);
nor U17795 (N_17795,N_17502,N_17406);
or U17796 (N_17796,N_17590,N_17417);
xor U17797 (N_17797,N_17496,N_17588);
and U17798 (N_17798,N_17412,N_17406);
nor U17799 (N_17799,N_17416,N_17519);
nand U17800 (N_17800,N_17797,N_17695);
nand U17801 (N_17801,N_17650,N_17606);
or U17802 (N_17802,N_17779,N_17787);
and U17803 (N_17803,N_17723,N_17624);
and U17804 (N_17804,N_17740,N_17700);
nor U17805 (N_17805,N_17639,N_17601);
nand U17806 (N_17806,N_17649,N_17789);
or U17807 (N_17807,N_17655,N_17702);
nand U17808 (N_17808,N_17753,N_17630);
nor U17809 (N_17809,N_17666,N_17759);
nor U17810 (N_17810,N_17646,N_17696);
nand U17811 (N_17811,N_17664,N_17620);
nand U17812 (N_17812,N_17713,N_17707);
nand U17813 (N_17813,N_17640,N_17660);
and U17814 (N_17814,N_17767,N_17791);
or U17815 (N_17815,N_17608,N_17651);
nor U17816 (N_17816,N_17637,N_17626);
nor U17817 (N_17817,N_17619,N_17751);
or U17818 (N_17818,N_17761,N_17647);
nand U17819 (N_17819,N_17720,N_17652);
and U17820 (N_17820,N_17677,N_17692);
and U17821 (N_17821,N_17605,N_17636);
or U17822 (N_17822,N_17673,N_17795);
nor U17823 (N_17823,N_17641,N_17718);
or U17824 (N_17824,N_17788,N_17726);
nand U17825 (N_17825,N_17722,N_17676);
and U17826 (N_17826,N_17776,N_17772);
xnor U17827 (N_17827,N_17682,N_17623);
and U17828 (N_17828,N_17735,N_17771);
and U17829 (N_17829,N_17627,N_17631);
or U17830 (N_17830,N_17749,N_17711);
or U17831 (N_17831,N_17780,N_17687);
nand U17832 (N_17832,N_17680,N_17763);
or U17833 (N_17833,N_17685,N_17739);
nand U17834 (N_17834,N_17633,N_17796);
nor U17835 (N_17835,N_17773,N_17667);
or U17836 (N_17836,N_17790,N_17609);
or U17837 (N_17837,N_17690,N_17777);
nand U17838 (N_17838,N_17629,N_17669);
and U17839 (N_17839,N_17625,N_17738);
or U17840 (N_17840,N_17600,N_17703);
nand U17841 (N_17841,N_17643,N_17716);
and U17842 (N_17842,N_17748,N_17634);
or U17843 (N_17843,N_17757,N_17607);
nor U17844 (N_17844,N_17662,N_17781);
nor U17845 (N_17845,N_17701,N_17622);
nor U17846 (N_17846,N_17628,N_17674);
nor U17847 (N_17847,N_17648,N_17783);
or U17848 (N_17848,N_17733,N_17708);
or U17849 (N_17849,N_17745,N_17766);
or U17850 (N_17850,N_17792,N_17719);
or U17851 (N_17851,N_17750,N_17712);
and U17852 (N_17852,N_17671,N_17727);
and U17853 (N_17853,N_17769,N_17747);
nand U17854 (N_17854,N_17621,N_17746);
nor U17855 (N_17855,N_17699,N_17778);
and U17856 (N_17856,N_17758,N_17752);
nand U17857 (N_17857,N_17618,N_17678);
nand U17858 (N_17858,N_17765,N_17775);
nor U17859 (N_17859,N_17675,N_17786);
and U17860 (N_17860,N_17668,N_17697);
and U17861 (N_17861,N_17706,N_17689);
and U17862 (N_17862,N_17617,N_17684);
nand U17863 (N_17863,N_17764,N_17782);
nand U17864 (N_17864,N_17612,N_17635);
and U17865 (N_17865,N_17611,N_17709);
and U17866 (N_17866,N_17683,N_17760);
or U17867 (N_17867,N_17604,N_17741);
nor U17868 (N_17868,N_17693,N_17691);
or U17869 (N_17869,N_17725,N_17661);
nor U17870 (N_17870,N_17762,N_17616);
nor U17871 (N_17871,N_17614,N_17659);
nor U17872 (N_17872,N_17704,N_17721);
nand U17873 (N_17873,N_17742,N_17686);
xnor U17874 (N_17874,N_17715,N_17732);
or U17875 (N_17875,N_17705,N_17657);
or U17876 (N_17876,N_17658,N_17724);
and U17877 (N_17877,N_17714,N_17602);
nor U17878 (N_17878,N_17799,N_17793);
or U17879 (N_17879,N_17615,N_17656);
or U17880 (N_17880,N_17785,N_17654);
nor U17881 (N_17881,N_17717,N_17698);
nand U17882 (N_17882,N_17645,N_17756);
and U17883 (N_17883,N_17784,N_17734);
and U17884 (N_17884,N_17665,N_17754);
nand U17885 (N_17885,N_17679,N_17736);
nand U17886 (N_17886,N_17798,N_17688);
or U17887 (N_17887,N_17603,N_17770);
or U17888 (N_17888,N_17644,N_17730);
and U17889 (N_17889,N_17613,N_17638);
nor U17890 (N_17890,N_17728,N_17610);
or U17891 (N_17891,N_17744,N_17681);
and U17892 (N_17892,N_17755,N_17653);
nand U17893 (N_17893,N_17774,N_17663);
nor U17894 (N_17894,N_17737,N_17670);
and U17895 (N_17895,N_17694,N_17632);
nor U17896 (N_17896,N_17768,N_17642);
nand U17897 (N_17897,N_17710,N_17672);
nand U17898 (N_17898,N_17743,N_17731);
and U17899 (N_17899,N_17729,N_17794);
and U17900 (N_17900,N_17644,N_17722);
and U17901 (N_17901,N_17695,N_17754);
nor U17902 (N_17902,N_17669,N_17721);
or U17903 (N_17903,N_17678,N_17627);
nor U17904 (N_17904,N_17613,N_17601);
nand U17905 (N_17905,N_17741,N_17683);
nand U17906 (N_17906,N_17727,N_17756);
nor U17907 (N_17907,N_17793,N_17779);
and U17908 (N_17908,N_17640,N_17700);
or U17909 (N_17909,N_17770,N_17754);
nor U17910 (N_17910,N_17694,N_17657);
or U17911 (N_17911,N_17748,N_17667);
and U17912 (N_17912,N_17751,N_17720);
nor U17913 (N_17913,N_17747,N_17660);
and U17914 (N_17914,N_17707,N_17632);
and U17915 (N_17915,N_17738,N_17759);
nand U17916 (N_17916,N_17619,N_17653);
and U17917 (N_17917,N_17764,N_17766);
and U17918 (N_17918,N_17667,N_17659);
nor U17919 (N_17919,N_17764,N_17613);
nor U17920 (N_17920,N_17689,N_17637);
nand U17921 (N_17921,N_17683,N_17744);
nand U17922 (N_17922,N_17735,N_17687);
and U17923 (N_17923,N_17796,N_17600);
nand U17924 (N_17924,N_17768,N_17624);
and U17925 (N_17925,N_17660,N_17654);
nand U17926 (N_17926,N_17743,N_17641);
and U17927 (N_17927,N_17639,N_17775);
and U17928 (N_17928,N_17688,N_17766);
nor U17929 (N_17929,N_17733,N_17779);
and U17930 (N_17930,N_17695,N_17648);
or U17931 (N_17931,N_17726,N_17791);
nor U17932 (N_17932,N_17665,N_17619);
and U17933 (N_17933,N_17740,N_17760);
nor U17934 (N_17934,N_17708,N_17698);
nand U17935 (N_17935,N_17625,N_17645);
and U17936 (N_17936,N_17794,N_17780);
and U17937 (N_17937,N_17695,N_17758);
and U17938 (N_17938,N_17743,N_17610);
xor U17939 (N_17939,N_17706,N_17605);
or U17940 (N_17940,N_17724,N_17678);
nand U17941 (N_17941,N_17693,N_17767);
nand U17942 (N_17942,N_17771,N_17683);
nand U17943 (N_17943,N_17778,N_17758);
nor U17944 (N_17944,N_17744,N_17780);
or U17945 (N_17945,N_17603,N_17631);
or U17946 (N_17946,N_17799,N_17687);
nand U17947 (N_17947,N_17658,N_17756);
nor U17948 (N_17948,N_17715,N_17616);
or U17949 (N_17949,N_17773,N_17640);
nor U17950 (N_17950,N_17699,N_17604);
and U17951 (N_17951,N_17745,N_17678);
nor U17952 (N_17952,N_17735,N_17621);
and U17953 (N_17953,N_17706,N_17770);
nand U17954 (N_17954,N_17665,N_17780);
or U17955 (N_17955,N_17606,N_17716);
and U17956 (N_17956,N_17656,N_17786);
nand U17957 (N_17957,N_17779,N_17659);
nor U17958 (N_17958,N_17650,N_17674);
nand U17959 (N_17959,N_17783,N_17743);
and U17960 (N_17960,N_17712,N_17609);
nand U17961 (N_17961,N_17793,N_17669);
nand U17962 (N_17962,N_17694,N_17623);
nand U17963 (N_17963,N_17722,N_17692);
or U17964 (N_17964,N_17663,N_17731);
nor U17965 (N_17965,N_17732,N_17798);
nor U17966 (N_17966,N_17771,N_17637);
and U17967 (N_17967,N_17680,N_17773);
or U17968 (N_17968,N_17668,N_17751);
nand U17969 (N_17969,N_17712,N_17739);
and U17970 (N_17970,N_17741,N_17761);
nor U17971 (N_17971,N_17772,N_17792);
nor U17972 (N_17972,N_17719,N_17669);
and U17973 (N_17973,N_17714,N_17636);
nand U17974 (N_17974,N_17644,N_17735);
or U17975 (N_17975,N_17695,N_17682);
nor U17976 (N_17976,N_17732,N_17741);
nor U17977 (N_17977,N_17726,N_17637);
nand U17978 (N_17978,N_17662,N_17600);
nand U17979 (N_17979,N_17760,N_17651);
or U17980 (N_17980,N_17652,N_17675);
and U17981 (N_17981,N_17795,N_17638);
and U17982 (N_17982,N_17663,N_17672);
and U17983 (N_17983,N_17666,N_17660);
nor U17984 (N_17984,N_17758,N_17772);
nand U17985 (N_17985,N_17600,N_17629);
nand U17986 (N_17986,N_17687,N_17769);
nand U17987 (N_17987,N_17652,N_17604);
nand U17988 (N_17988,N_17639,N_17739);
or U17989 (N_17989,N_17753,N_17670);
and U17990 (N_17990,N_17782,N_17736);
or U17991 (N_17991,N_17767,N_17715);
nand U17992 (N_17992,N_17777,N_17614);
and U17993 (N_17993,N_17604,N_17607);
nor U17994 (N_17994,N_17715,N_17756);
and U17995 (N_17995,N_17677,N_17704);
or U17996 (N_17996,N_17793,N_17603);
and U17997 (N_17997,N_17794,N_17749);
and U17998 (N_17998,N_17716,N_17658);
nand U17999 (N_17999,N_17723,N_17769);
and U18000 (N_18000,N_17999,N_17895);
nor U18001 (N_18001,N_17950,N_17929);
nor U18002 (N_18002,N_17813,N_17932);
nand U18003 (N_18003,N_17982,N_17877);
or U18004 (N_18004,N_17904,N_17892);
and U18005 (N_18005,N_17921,N_17947);
nor U18006 (N_18006,N_17946,N_17860);
and U18007 (N_18007,N_17882,N_17839);
nand U18008 (N_18008,N_17807,N_17937);
and U18009 (N_18009,N_17925,N_17900);
nor U18010 (N_18010,N_17881,N_17893);
nor U18011 (N_18011,N_17919,N_17806);
or U18012 (N_18012,N_17983,N_17909);
nand U18013 (N_18013,N_17965,N_17942);
or U18014 (N_18014,N_17811,N_17966);
nor U18015 (N_18015,N_17988,N_17916);
and U18016 (N_18016,N_17803,N_17976);
xnor U18017 (N_18017,N_17908,N_17869);
nand U18018 (N_18018,N_17961,N_17912);
nor U18019 (N_18019,N_17867,N_17948);
nor U18020 (N_18020,N_17801,N_17923);
nand U18021 (N_18021,N_17933,N_17943);
nand U18022 (N_18022,N_17858,N_17967);
or U18023 (N_18023,N_17821,N_17805);
or U18024 (N_18024,N_17838,N_17851);
and U18025 (N_18025,N_17915,N_17934);
and U18026 (N_18026,N_17956,N_17986);
nand U18027 (N_18027,N_17927,N_17833);
nor U18028 (N_18028,N_17917,N_17889);
and U18029 (N_18029,N_17940,N_17853);
or U18030 (N_18030,N_17864,N_17953);
nor U18031 (N_18031,N_17969,N_17876);
or U18032 (N_18032,N_17826,N_17959);
nor U18033 (N_18033,N_17854,N_17879);
and U18034 (N_18034,N_17842,N_17989);
or U18035 (N_18035,N_17981,N_17987);
nand U18036 (N_18036,N_17861,N_17824);
nor U18037 (N_18037,N_17905,N_17939);
nand U18038 (N_18038,N_17998,N_17993);
nand U18039 (N_18039,N_17804,N_17852);
or U18040 (N_18040,N_17836,N_17949);
nand U18041 (N_18041,N_17840,N_17902);
nor U18042 (N_18042,N_17935,N_17883);
nor U18043 (N_18043,N_17859,N_17870);
nand U18044 (N_18044,N_17931,N_17812);
nor U18045 (N_18045,N_17868,N_17907);
and U18046 (N_18046,N_17825,N_17897);
and U18047 (N_18047,N_17835,N_17984);
nand U18048 (N_18048,N_17880,N_17847);
nand U18049 (N_18049,N_17928,N_17894);
and U18050 (N_18050,N_17862,N_17960);
or U18051 (N_18051,N_17941,N_17848);
nand U18052 (N_18052,N_17898,N_17954);
nand U18053 (N_18053,N_17816,N_17944);
or U18054 (N_18054,N_17834,N_17913);
or U18055 (N_18055,N_17885,N_17957);
nand U18056 (N_18056,N_17841,N_17963);
nand U18057 (N_18057,N_17971,N_17996);
nand U18058 (N_18058,N_17992,N_17964);
nor U18059 (N_18059,N_17846,N_17962);
nand U18060 (N_18060,N_17810,N_17903);
nand U18061 (N_18061,N_17936,N_17832);
and U18062 (N_18062,N_17977,N_17856);
xor U18063 (N_18063,N_17844,N_17910);
and U18064 (N_18064,N_17850,N_17849);
or U18065 (N_18065,N_17970,N_17828);
and U18066 (N_18066,N_17878,N_17820);
and U18067 (N_18067,N_17918,N_17823);
or U18068 (N_18068,N_17814,N_17817);
or U18069 (N_18069,N_17926,N_17899);
nand U18070 (N_18070,N_17955,N_17920);
nor U18071 (N_18071,N_17974,N_17887);
or U18072 (N_18072,N_17831,N_17975);
or U18073 (N_18073,N_17924,N_17827);
nor U18074 (N_18074,N_17865,N_17991);
and U18075 (N_18075,N_17980,N_17930);
xnor U18076 (N_18076,N_17994,N_17997);
and U18077 (N_18077,N_17843,N_17873);
and U18078 (N_18078,N_17990,N_17973);
or U18079 (N_18079,N_17815,N_17800);
nor U18080 (N_18080,N_17857,N_17978);
or U18081 (N_18081,N_17891,N_17872);
nor U18082 (N_18082,N_17985,N_17875);
nand U18083 (N_18083,N_17938,N_17888);
nand U18084 (N_18084,N_17886,N_17979);
nand U18085 (N_18085,N_17802,N_17819);
or U18086 (N_18086,N_17922,N_17837);
nand U18087 (N_18087,N_17866,N_17808);
or U18088 (N_18088,N_17995,N_17822);
or U18089 (N_18089,N_17951,N_17945);
nand U18090 (N_18090,N_17890,N_17818);
and U18091 (N_18091,N_17829,N_17901);
nor U18092 (N_18092,N_17914,N_17958);
and U18093 (N_18093,N_17863,N_17874);
nor U18094 (N_18094,N_17845,N_17911);
nand U18095 (N_18095,N_17968,N_17884);
nor U18096 (N_18096,N_17830,N_17906);
or U18097 (N_18097,N_17809,N_17855);
or U18098 (N_18098,N_17952,N_17972);
nor U18099 (N_18099,N_17896,N_17871);
and U18100 (N_18100,N_17877,N_17989);
nor U18101 (N_18101,N_17855,N_17859);
nor U18102 (N_18102,N_17937,N_17854);
nand U18103 (N_18103,N_17827,N_17807);
and U18104 (N_18104,N_17971,N_17804);
and U18105 (N_18105,N_17990,N_17957);
nand U18106 (N_18106,N_17907,N_17855);
and U18107 (N_18107,N_17951,N_17830);
and U18108 (N_18108,N_17992,N_17910);
and U18109 (N_18109,N_17918,N_17837);
or U18110 (N_18110,N_17809,N_17837);
or U18111 (N_18111,N_17940,N_17802);
nor U18112 (N_18112,N_17965,N_17875);
and U18113 (N_18113,N_17959,N_17983);
and U18114 (N_18114,N_17980,N_17905);
and U18115 (N_18115,N_17801,N_17996);
and U18116 (N_18116,N_17847,N_17877);
nor U18117 (N_18117,N_17821,N_17986);
nand U18118 (N_18118,N_17951,N_17917);
nor U18119 (N_18119,N_17927,N_17897);
and U18120 (N_18120,N_17835,N_17931);
nor U18121 (N_18121,N_17936,N_17845);
and U18122 (N_18122,N_17942,N_17918);
or U18123 (N_18123,N_17857,N_17836);
nand U18124 (N_18124,N_17939,N_17841);
nand U18125 (N_18125,N_17895,N_17867);
nor U18126 (N_18126,N_17862,N_17889);
and U18127 (N_18127,N_17846,N_17971);
nand U18128 (N_18128,N_17817,N_17879);
or U18129 (N_18129,N_17890,N_17856);
and U18130 (N_18130,N_17972,N_17884);
xnor U18131 (N_18131,N_17937,N_17923);
and U18132 (N_18132,N_17910,N_17946);
or U18133 (N_18133,N_17838,N_17969);
or U18134 (N_18134,N_17849,N_17930);
nor U18135 (N_18135,N_17926,N_17915);
or U18136 (N_18136,N_17944,N_17875);
nand U18137 (N_18137,N_17944,N_17857);
nand U18138 (N_18138,N_17988,N_17929);
or U18139 (N_18139,N_17846,N_17809);
and U18140 (N_18140,N_17918,N_17970);
or U18141 (N_18141,N_17885,N_17830);
or U18142 (N_18142,N_17992,N_17919);
nor U18143 (N_18143,N_17805,N_17935);
nor U18144 (N_18144,N_17950,N_17964);
nand U18145 (N_18145,N_17959,N_17850);
and U18146 (N_18146,N_17959,N_17973);
nand U18147 (N_18147,N_17838,N_17942);
or U18148 (N_18148,N_17926,N_17881);
nand U18149 (N_18149,N_17950,N_17970);
and U18150 (N_18150,N_17860,N_17967);
and U18151 (N_18151,N_17979,N_17969);
xor U18152 (N_18152,N_17890,N_17837);
or U18153 (N_18153,N_17828,N_17897);
nand U18154 (N_18154,N_17806,N_17884);
nand U18155 (N_18155,N_17975,N_17849);
nor U18156 (N_18156,N_17883,N_17965);
or U18157 (N_18157,N_17875,N_17876);
nor U18158 (N_18158,N_17919,N_17947);
nand U18159 (N_18159,N_17867,N_17808);
nor U18160 (N_18160,N_17869,N_17949);
or U18161 (N_18161,N_17946,N_17819);
nand U18162 (N_18162,N_17994,N_17887);
and U18163 (N_18163,N_17881,N_17940);
or U18164 (N_18164,N_17831,N_17989);
and U18165 (N_18165,N_17997,N_17866);
nor U18166 (N_18166,N_17934,N_17865);
nand U18167 (N_18167,N_17969,N_17843);
and U18168 (N_18168,N_17847,N_17923);
nor U18169 (N_18169,N_17826,N_17874);
nor U18170 (N_18170,N_17893,N_17824);
nand U18171 (N_18171,N_17942,N_17852);
nand U18172 (N_18172,N_17873,N_17831);
nand U18173 (N_18173,N_17936,N_17950);
nor U18174 (N_18174,N_17841,N_17980);
nor U18175 (N_18175,N_17959,N_17876);
or U18176 (N_18176,N_17924,N_17843);
or U18177 (N_18177,N_17995,N_17846);
xnor U18178 (N_18178,N_17971,N_17878);
and U18179 (N_18179,N_17814,N_17829);
nor U18180 (N_18180,N_17844,N_17963);
and U18181 (N_18181,N_17865,N_17860);
nor U18182 (N_18182,N_17934,N_17834);
nor U18183 (N_18183,N_17876,N_17830);
nand U18184 (N_18184,N_17968,N_17991);
and U18185 (N_18185,N_17998,N_17865);
or U18186 (N_18186,N_17896,N_17898);
or U18187 (N_18187,N_17929,N_17965);
nand U18188 (N_18188,N_17811,N_17902);
and U18189 (N_18189,N_17954,N_17976);
nand U18190 (N_18190,N_17959,N_17868);
nand U18191 (N_18191,N_17995,N_17851);
nor U18192 (N_18192,N_17848,N_17929);
or U18193 (N_18193,N_17834,N_17922);
or U18194 (N_18194,N_17901,N_17917);
nor U18195 (N_18195,N_17975,N_17930);
or U18196 (N_18196,N_17846,N_17975);
nand U18197 (N_18197,N_17817,N_17875);
nand U18198 (N_18198,N_17939,N_17952);
nand U18199 (N_18199,N_17943,N_17838);
nor U18200 (N_18200,N_18109,N_18122);
and U18201 (N_18201,N_18187,N_18143);
nand U18202 (N_18202,N_18192,N_18150);
nand U18203 (N_18203,N_18072,N_18000);
nand U18204 (N_18204,N_18060,N_18044);
and U18205 (N_18205,N_18160,N_18119);
nor U18206 (N_18206,N_18046,N_18134);
nand U18207 (N_18207,N_18085,N_18196);
and U18208 (N_18208,N_18091,N_18080);
nor U18209 (N_18209,N_18132,N_18041);
and U18210 (N_18210,N_18069,N_18076);
nand U18211 (N_18211,N_18012,N_18089);
nor U18212 (N_18212,N_18023,N_18179);
or U18213 (N_18213,N_18026,N_18099);
and U18214 (N_18214,N_18038,N_18024);
or U18215 (N_18215,N_18074,N_18015);
nor U18216 (N_18216,N_18031,N_18198);
nor U18217 (N_18217,N_18040,N_18156);
and U18218 (N_18218,N_18093,N_18059);
or U18219 (N_18219,N_18182,N_18083);
nor U18220 (N_18220,N_18006,N_18184);
nand U18221 (N_18221,N_18186,N_18007);
nand U18222 (N_18222,N_18016,N_18079);
nand U18223 (N_18223,N_18062,N_18126);
nor U18224 (N_18224,N_18029,N_18128);
nor U18225 (N_18225,N_18125,N_18051);
nand U18226 (N_18226,N_18195,N_18153);
and U18227 (N_18227,N_18148,N_18088);
nor U18228 (N_18228,N_18170,N_18141);
nand U18229 (N_18229,N_18139,N_18121);
nor U18230 (N_18230,N_18193,N_18004);
and U18231 (N_18231,N_18147,N_18131);
nor U18232 (N_18232,N_18105,N_18114);
or U18233 (N_18233,N_18057,N_18096);
and U18234 (N_18234,N_18108,N_18100);
and U18235 (N_18235,N_18138,N_18166);
or U18236 (N_18236,N_18036,N_18117);
and U18237 (N_18237,N_18053,N_18102);
nor U18238 (N_18238,N_18142,N_18037);
nand U18239 (N_18239,N_18173,N_18033);
nor U18240 (N_18240,N_18052,N_18106);
and U18241 (N_18241,N_18162,N_18055);
nor U18242 (N_18242,N_18043,N_18118);
and U18243 (N_18243,N_18068,N_18094);
and U18244 (N_18244,N_18071,N_18161);
and U18245 (N_18245,N_18073,N_18191);
and U18246 (N_18246,N_18017,N_18020);
nor U18247 (N_18247,N_18078,N_18097);
or U18248 (N_18248,N_18155,N_18154);
nand U18249 (N_18249,N_18169,N_18075);
nand U18250 (N_18250,N_18087,N_18077);
nand U18251 (N_18251,N_18005,N_18149);
and U18252 (N_18252,N_18144,N_18098);
or U18253 (N_18253,N_18110,N_18181);
and U18254 (N_18254,N_18066,N_18022);
or U18255 (N_18255,N_18045,N_18164);
nand U18256 (N_18256,N_18009,N_18030);
nor U18257 (N_18257,N_18190,N_18027);
and U18258 (N_18258,N_18034,N_18129);
or U18259 (N_18259,N_18130,N_18002);
or U18260 (N_18260,N_18157,N_18058);
or U18261 (N_18261,N_18003,N_18177);
or U18262 (N_18262,N_18035,N_18103);
nand U18263 (N_18263,N_18112,N_18146);
nor U18264 (N_18264,N_18048,N_18197);
nand U18265 (N_18265,N_18188,N_18104);
xor U18266 (N_18266,N_18070,N_18019);
nand U18267 (N_18267,N_18171,N_18199);
and U18268 (N_18268,N_18064,N_18140);
or U18269 (N_18269,N_18127,N_18152);
or U18270 (N_18270,N_18111,N_18175);
and U18271 (N_18271,N_18174,N_18047);
and U18272 (N_18272,N_18158,N_18065);
nand U18273 (N_18273,N_18189,N_18159);
nor U18274 (N_18274,N_18137,N_18063);
and U18275 (N_18275,N_18050,N_18135);
or U18276 (N_18276,N_18101,N_18123);
nand U18277 (N_18277,N_18194,N_18136);
xnor U18278 (N_18278,N_18185,N_18082);
and U18279 (N_18279,N_18011,N_18049);
nor U18280 (N_18280,N_18013,N_18151);
or U18281 (N_18281,N_18001,N_18061);
nand U18282 (N_18282,N_18124,N_18120);
and U18283 (N_18283,N_18084,N_18113);
and U18284 (N_18284,N_18090,N_18042);
nor U18285 (N_18285,N_18163,N_18167);
nor U18286 (N_18286,N_18032,N_18176);
nor U18287 (N_18287,N_18168,N_18025);
nor U18288 (N_18288,N_18178,N_18067);
and U18289 (N_18289,N_18021,N_18180);
nor U18290 (N_18290,N_18086,N_18145);
nor U18291 (N_18291,N_18018,N_18010);
nand U18292 (N_18292,N_18081,N_18172);
and U18293 (N_18293,N_18183,N_18039);
or U18294 (N_18294,N_18008,N_18165);
nor U18295 (N_18295,N_18028,N_18092);
nor U18296 (N_18296,N_18056,N_18133);
nand U18297 (N_18297,N_18095,N_18014);
and U18298 (N_18298,N_18054,N_18107);
and U18299 (N_18299,N_18115,N_18116);
or U18300 (N_18300,N_18103,N_18047);
nor U18301 (N_18301,N_18010,N_18198);
nor U18302 (N_18302,N_18158,N_18071);
and U18303 (N_18303,N_18045,N_18167);
or U18304 (N_18304,N_18071,N_18061);
and U18305 (N_18305,N_18067,N_18027);
nor U18306 (N_18306,N_18160,N_18108);
nand U18307 (N_18307,N_18116,N_18085);
and U18308 (N_18308,N_18012,N_18092);
and U18309 (N_18309,N_18067,N_18167);
or U18310 (N_18310,N_18017,N_18032);
nor U18311 (N_18311,N_18135,N_18031);
nor U18312 (N_18312,N_18064,N_18143);
nor U18313 (N_18313,N_18008,N_18085);
nor U18314 (N_18314,N_18141,N_18089);
nand U18315 (N_18315,N_18116,N_18070);
nand U18316 (N_18316,N_18153,N_18042);
nand U18317 (N_18317,N_18148,N_18188);
nand U18318 (N_18318,N_18142,N_18139);
nand U18319 (N_18319,N_18142,N_18075);
nand U18320 (N_18320,N_18049,N_18069);
nor U18321 (N_18321,N_18077,N_18189);
nand U18322 (N_18322,N_18000,N_18101);
nor U18323 (N_18323,N_18100,N_18020);
nand U18324 (N_18324,N_18136,N_18016);
nand U18325 (N_18325,N_18183,N_18093);
or U18326 (N_18326,N_18121,N_18046);
or U18327 (N_18327,N_18015,N_18081);
nor U18328 (N_18328,N_18075,N_18153);
nor U18329 (N_18329,N_18056,N_18093);
and U18330 (N_18330,N_18143,N_18158);
nand U18331 (N_18331,N_18169,N_18065);
or U18332 (N_18332,N_18194,N_18077);
and U18333 (N_18333,N_18194,N_18020);
nand U18334 (N_18334,N_18186,N_18054);
or U18335 (N_18335,N_18171,N_18151);
and U18336 (N_18336,N_18019,N_18118);
nand U18337 (N_18337,N_18189,N_18132);
nand U18338 (N_18338,N_18153,N_18099);
nor U18339 (N_18339,N_18122,N_18098);
or U18340 (N_18340,N_18183,N_18136);
nand U18341 (N_18341,N_18021,N_18158);
xnor U18342 (N_18342,N_18175,N_18189);
nor U18343 (N_18343,N_18191,N_18059);
or U18344 (N_18344,N_18143,N_18154);
or U18345 (N_18345,N_18128,N_18166);
xor U18346 (N_18346,N_18129,N_18076);
and U18347 (N_18347,N_18114,N_18014);
nor U18348 (N_18348,N_18044,N_18003);
nor U18349 (N_18349,N_18004,N_18102);
or U18350 (N_18350,N_18095,N_18046);
or U18351 (N_18351,N_18010,N_18074);
and U18352 (N_18352,N_18120,N_18194);
nor U18353 (N_18353,N_18180,N_18050);
nor U18354 (N_18354,N_18089,N_18007);
nor U18355 (N_18355,N_18098,N_18165);
nand U18356 (N_18356,N_18126,N_18025);
and U18357 (N_18357,N_18113,N_18129);
nor U18358 (N_18358,N_18199,N_18000);
nor U18359 (N_18359,N_18034,N_18130);
nand U18360 (N_18360,N_18056,N_18066);
nor U18361 (N_18361,N_18180,N_18184);
or U18362 (N_18362,N_18128,N_18025);
and U18363 (N_18363,N_18085,N_18061);
or U18364 (N_18364,N_18181,N_18070);
nand U18365 (N_18365,N_18022,N_18085);
and U18366 (N_18366,N_18087,N_18176);
nor U18367 (N_18367,N_18115,N_18102);
nand U18368 (N_18368,N_18090,N_18046);
and U18369 (N_18369,N_18023,N_18031);
or U18370 (N_18370,N_18135,N_18130);
nor U18371 (N_18371,N_18048,N_18177);
nand U18372 (N_18372,N_18152,N_18137);
or U18373 (N_18373,N_18012,N_18143);
nor U18374 (N_18374,N_18008,N_18088);
and U18375 (N_18375,N_18179,N_18102);
nor U18376 (N_18376,N_18013,N_18145);
and U18377 (N_18377,N_18124,N_18117);
nor U18378 (N_18378,N_18012,N_18083);
nand U18379 (N_18379,N_18092,N_18165);
nand U18380 (N_18380,N_18045,N_18141);
nor U18381 (N_18381,N_18017,N_18061);
nand U18382 (N_18382,N_18102,N_18137);
nand U18383 (N_18383,N_18043,N_18199);
nand U18384 (N_18384,N_18029,N_18086);
and U18385 (N_18385,N_18036,N_18152);
or U18386 (N_18386,N_18115,N_18114);
nor U18387 (N_18387,N_18003,N_18172);
or U18388 (N_18388,N_18046,N_18037);
nand U18389 (N_18389,N_18035,N_18192);
or U18390 (N_18390,N_18093,N_18009);
nor U18391 (N_18391,N_18104,N_18087);
or U18392 (N_18392,N_18103,N_18033);
and U18393 (N_18393,N_18022,N_18182);
or U18394 (N_18394,N_18025,N_18033);
nor U18395 (N_18395,N_18003,N_18017);
nand U18396 (N_18396,N_18063,N_18197);
nand U18397 (N_18397,N_18006,N_18050);
nor U18398 (N_18398,N_18019,N_18137);
nor U18399 (N_18399,N_18088,N_18173);
and U18400 (N_18400,N_18276,N_18334);
nand U18401 (N_18401,N_18370,N_18267);
nand U18402 (N_18402,N_18294,N_18331);
and U18403 (N_18403,N_18371,N_18242);
nor U18404 (N_18404,N_18323,N_18224);
nand U18405 (N_18405,N_18306,N_18304);
nand U18406 (N_18406,N_18289,N_18253);
nor U18407 (N_18407,N_18303,N_18333);
and U18408 (N_18408,N_18216,N_18375);
nor U18409 (N_18409,N_18384,N_18219);
and U18410 (N_18410,N_18277,N_18229);
nor U18411 (N_18411,N_18374,N_18260);
nand U18412 (N_18412,N_18344,N_18360);
or U18413 (N_18413,N_18317,N_18214);
xor U18414 (N_18414,N_18350,N_18366);
and U18415 (N_18415,N_18330,N_18337);
or U18416 (N_18416,N_18359,N_18209);
nor U18417 (N_18417,N_18223,N_18314);
nor U18418 (N_18418,N_18272,N_18358);
nand U18419 (N_18419,N_18288,N_18285);
nand U18420 (N_18420,N_18259,N_18365);
and U18421 (N_18421,N_18220,N_18227);
nand U18422 (N_18422,N_18269,N_18257);
xnor U18423 (N_18423,N_18393,N_18212);
nor U18424 (N_18424,N_18222,N_18316);
or U18425 (N_18425,N_18273,N_18327);
or U18426 (N_18426,N_18200,N_18263);
nand U18427 (N_18427,N_18286,N_18310);
nand U18428 (N_18428,N_18213,N_18324);
nand U18429 (N_18429,N_18287,N_18387);
and U18430 (N_18430,N_18210,N_18398);
or U18431 (N_18431,N_18347,N_18228);
and U18432 (N_18432,N_18352,N_18315);
nand U18433 (N_18433,N_18329,N_18308);
nand U18434 (N_18434,N_18397,N_18231);
and U18435 (N_18435,N_18215,N_18250);
nor U18436 (N_18436,N_18355,N_18258);
nand U18437 (N_18437,N_18338,N_18299);
or U18438 (N_18438,N_18206,N_18379);
nand U18439 (N_18439,N_18280,N_18394);
and U18440 (N_18440,N_18364,N_18270);
nor U18441 (N_18441,N_18348,N_18311);
and U18442 (N_18442,N_18262,N_18318);
and U18443 (N_18443,N_18268,N_18255);
nand U18444 (N_18444,N_18254,N_18335);
and U18445 (N_18445,N_18266,N_18246);
or U18446 (N_18446,N_18353,N_18251);
and U18447 (N_18447,N_18332,N_18373);
and U18448 (N_18448,N_18325,N_18377);
or U18449 (N_18449,N_18271,N_18217);
nand U18450 (N_18450,N_18345,N_18381);
or U18451 (N_18451,N_18321,N_18305);
nand U18452 (N_18452,N_18367,N_18320);
nand U18453 (N_18453,N_18221,N_18351);
and U18454 (N_18454,N_18386,N_18357);
and U18455 (N_18455,N_18207,N_18342);
nand U18456 (N_18456,N_18233,N_18201);
or U18457 (N_18457,N_18298,N_18237);
and U18458 (N_18458,N_18248,N_18346);
and U18459 (N_18459,N_18247,N_18378);
nand U18460 (N_18460,N_18389,N_18380);
or U18461 (N_18461,N_18278,N_18283);
and U18462 (N_18462,N_18309,N_18261);
nand U18463 (N_18463,N_18225,N_18362);
nand U18464 (N_18464,N_18336,N_18243);
nand U18465 (N_18465,N_18249,N_18244);
or U18466 (N_18466,N_18234,N_18290);
and U18467 (N_18467,N_18382,N_18363);
nor U18468 (N_18468,N_18313,N_18300);
or U18469 (N_18469,N_18343,N_18238);
xnor U18470 (N_18470,N_18291,N_18226);
nor U18471 (N_18471,N_18395,N_18203);
nand U18472 (N_18472,N_18349,N_18296);
or U18473 (N_18473,N_18274,N_18385);
nand U18474 (N_18474,N_18293,N_18328);
or U18475 (N_18475,N_18340,N_18307);
or U18476 (N_18476,N_18383,N_18295);
and U18477 (N_18477,N_18275,N_18376);
nor U18478 (N_18478,N_18399,N_18235);
and U18479 (N_18479,N_18211,N_18281);
nand U18480 (N_18480,N_18372,N_18319);
nand U18481 (N_18481,N_18391,N_18284);
nand U18482 (N_18482,N_18265,N_18369);
or U18483 (N_18483,N_18252,N_18301);
xnor U18484 (N_18484,N_18264,N_18356);
or U18485 (N_18485,N_18322,N_18240);
and U18486 (N_18486,N_18230,N_18392);
nor U18487 (N_18487,N_18302,N_18354);
nand U18488 (N_18488,N_18236,N_18292);
or U18489 (N_18489,N_18339,N_18361);
nand U18490 (N_18490,N_18204,N_18256);
and U18491 (N_18491,N_18205,N_18239);
and U18492 (N_18492,N_18208,N_18218);
nand U18493 (N_18493,N_18326,N_18245);
or U18494 (N_18494,N_18297,N_18241);
nor U18495 (N_18495,N_18368,N_18388);
or U18496 (N_18496,N_18202,N_18390);
nor U18497 (N_18497,N_18232,N_18312);
or U18498 (N_18498,N_18282,N_18396);
nor U18499 (N_18499,N_18279,N_18341);
and U18500 (N_18500,N_18335,N_18363);
or U18501 (N_18501,N_18230,N_18283);
and U18502 (N_18502,N_18370,N_18318);
nor U18503 (N_18503,N_18210,N_18209);
and U18504 (N_18504,N_18229,N_18299);
and U18505 (N_18505,N_18259,N_18286);
or U18506 (N_18506,N_18207,N_18300);
nand U18507 (N_18507,N_18385,N_18380);
or U18508 (N_18508,N_18299,N_18269);
and U18509 (N_18509,N_18320,N_18200);
nor U18510 (N_18510,N_18292,N_18270);
nand U18511 (N_18511,N_18265,N_18361);
nor U18512 (N_18512,N_18218,N_18309);
and U18513 (N_18513,N_18223,N_18342);
nor U18514 (N_18514,N_18287,N_18359);
or U18515 (N_18515,N_18347,N_18354);
or U18516 (N_18516,N_18330,N_18232);
and U18517 (N_18517,N_18229,N_18372);
or U18518 (N_18518,N_18288,N_18303);
or U18519 (N_18519,N_18345,N_18301);
and U18520 (N_18520,N_18244,N_18376);
or U18521 (N_18521,N_18330,N_18283);
or U18522 (N_18522,N_18374,N_18369);
and U18523 (N_18523,N_18224,N_18244);
nor U18524 (N_18524,N_18233,N_18363);
and U18525 (N_18525,N_18319,N_18235);
or U18526 (N_18526,N_18250,N_18286);
and U18527 (N_18527,N_18359,N_18366);
nand U18528 (N_18528,N_18239,N_18329);
nand U18529 (N_18529,N_18287,N_18297);
or U18530 (N_18530,N_18223,N_18369);
nand U18531 (N_18531,N_18238,N_18297);
or U18532 (N_18532,N_18211,N_18300);
and U18533 (N_18533,N_18240,N_18201);
or U18534 (N_18534,N_18298,N_18254);
or U18535 (N_18535,N_18274,N_18383);
nand U18536 (N_18536,N_18313,N_18378);
nand U18537 (N_18537,N_18258,N_18368);
nand U18538 (N_18538,N_18232,N_18381);
nand U18539 (N_18539,N_18280,N_18345);
nor U18540 (N_18540,N_18361,N_18203);
nand U18541 (N_18541,N_18296,N_18224);
nand U18542 (N_18542,N_18332,N_18376);
nor U18543 (N_18543,N_18358,N_18203);
or U18544 (N_18544,N_18390,N_18303);
nor U18545 (N_18545,N_18394,N_18258);
nor U18546 (N_18546,N_18370,N_18214);
nor U18547 (N_18547,N_18226,N_18259);
and U18548 (N_18548,N_18331,N_18255);
nor U18549 (N_18549,N_18350,N_18299);
nand U18550 (N_18550,N_18224,N_18267);
nor U18551 (N_18551,N_18384,N_18357);
or U18552 (N_18552,N_18308,N_18330);
nand U18553 (N_18553,N_18267,N_18203);
nor U18554 (N_18554,N_18227,N_18216);
and U18555 (N_18555,N_18217,N_18294);
and U18556 (N_18556,N_18316,N_18355);
or U18557 (N_18557,N_18234,N_18353);
nand U18558 (N_18558,N_18279,N_18333);
and U18559 (N_18559,N_18358,N_18387);
and U18560 (N_18560,N_18310,N_18285);
nor U18561 (N_18561,N_18317,N_18348);
nor U18562 (N_18562,N_18252,N_18333);
and U18563 (N_18563,N_18303,N_18354);
nor U18564 (N_18564,N_18228,N_18363);
nand U18565 (N_18565,N_18259,N_18275);
or U18566 (N_18566,N_18240,N_18306);
nor U18567 (N_18567,N_18219,N_18289);
nor U18568 (N_18568,N_18331,N_18306);
nor U18569 (N_18569,N_18273,N_18321);
and U18570 (N_18570,N_18388,N_18274);
nand U18571 (N_18571,N_18391,N_18249);
nand U18572 (N_18572,N_18258,N_18339);
or U18573 (N_18573,N_18229,N_18232);
or U18574 (N_18574,N_18317,N_18356);
or U18575 (N_18575,N_18245,N_18274);
and U18576 (N_18576,N_18202,N_18276);
or U18577 (N_18577,N_18257,N_18313);
nand U18578 (N_18578,N_18284,N_18280);
nand U18579 (N_18579,N_18225,N_18207);
nand U18580 (N_18580,N_18261,N_18327);
nor U18581 (N_18581,N_18301,N_18362);
nor U18582 (N_18582,N_18248,N_18383);
nand U18583 (N_18583,N_18391,N_18293);
and U18584 (N_18584,N_18216,N_18316);
nand U18585 (N_18585,N_18260,N_18316);
nor U18586 (N_18586,N_18225,N_18258);
or U18587 (N_18587,N_18280,N_18229);
and U18588 (N_18588,N_18386,N_18389);
and U18589 (N_18589,N_18369,N_18389);
and U18590 (N_18590,N_18378,N_18328);
nand U18591 (N_18591,N_18357,N_18295);
and U18592 (N_18592,N_18380,N_18208);
nor U18593 (N_18593,N_18368,N_18386);
and U18594 (N_18594,N_18334,N_18369);
xnor U18595 (N_18595,N_18276,N_18312);
or U18596 (N_18596,N_18338,N_18262);
nand U18597 (N_18597,N_18373,N_18342);
nand U18598 (N_18598,N_18337,N_18216);
nand U18599 (N_18599,N_18227,N_18366);
nand U18600 (N_18600,N_18412,N_18551);
and U18601 (N_18601,N_18504,N_18482);
nand U18602 (N_18602,N_18544,N_18578);
nor U18603 (N_18603,N_18450,N_18521);
nand U18604 (N_18604,N_18507,N_18524);
nor U18605 (N_18605,N_18403,N_18523);
or U18606 (N_18606,N_18468,N_18500);
or U18607 (N_18607,N_18470,N_18447);
nand U18608 (N_18608,N_18552,N_18406);
or U18609 (N_18609,N_18461,N_18596);
or U18610 (N_18610,N_18430,N_18416);
nand U18611 (N_18611,N_18593,N_18543);
or U18612 (N_18612,N_18590,N_18548);
nor U18613 (N_18613,N_18539,N_18565);
or U18614 (N_18614,N_18553,N_18518);
or U18615 (N_18615,N_18560,N_18437);
or U18616 (N_18616,N_18558,N_18452);
and U18617 (N_18617,N_18555,N_18574);
nand U18618 (N_18618,N_18449,N_18567);
or U18619 (N_18619,N_18425,N_18443);
or U18620 (N_18620,N_18448,N_18409);
and U18621 (N_18621,N_18480,N_18444);
nand U18622 (N_18622,N_18534,N_18421);
or U18623 (N_18623,N_18428,N_18554);
nor U18624 (N_18624,N_18549,N_18458);
nand U18625 (N_18625,N_18445,N_18464);
or U18626 (N_18626,N_18556,N_18575);
or U18627 (N_18627,N_18513,N_18426);
nand U18628 (N_18628,N_18431,N_18442);
nor U18629 (N_18629,N_18400,N_18429);
or U18630 (N_18630,N_18503,N_18572);
nor U18631 (N_18631,N_18533,N_18446);
nand U18632 (N_18632,N_18517,N_18414);
nand U18633 (N_18633,N_18547,N_18440);
xor U18634 (N_18634,N_18516,N_18487);
nand U18635 (N_18635,N_18459,N_18413);
or U18636 (N_18636,N_18581,N_18420);
or U18637 (N_18637,N_18514,N_18410);
or U18638 (N_18638,N_18502,N_18474);
nor U18639 (N_18639,N_18599,N_18479);
nor U18640 (N_18640,N_18454,N_18419);
or U18641 (N_18641,N_18436,N_18490);
and U18642 (N_18642,N_18569,N_18540);
or U18643 (N_18643,N_18485,N_18417);
and U18644 (N_18644,N_18492,N_18453);
and U18645 (N_18645,N_18491,N_18463);
nand U18646 (N_18646,N_18597,N_18531);
or U18647 (N_18647,N_18477,N_18481);
or U18648 (N_18648,N_18471,N_18594);
and U18649 (N_18649,N_18573,N_18465);
nor U18650 (N_18650,N_18562,N_18592);
or U18651 (N_18651,N_18501,N_18579);
or U18652 (N_18652,N_18422,N_18435);
nor U18653 (N_18653,N_18561,N_18402);
nor U18654 (N_18654,N_18499,N_18401);
nand U18655 (N_18655,N_18484,N_18589);
nor U18656 (N_18656,N_18432,N_18576);
and U18657 (N_18657,N_18472,N_18585);
or U18658 (N_18658,N_18509,N_18530);
nor U18659 (N_18659,N_18498,N_18489);
or U18660 (N_18660,N_18525,N_18456);
nand U18661 (N_18661,N_18423,N_18510);
and U18662 (N_18662,N_18418,N_18529);
nand U18663 (N_18663,N_18404,N_18469);
nand U18664 (N_18664,N_18522,N_18494);
xnor U18665 (N_18665,N_18515,N_18538);
or U18666 (N_18666,N_18546,N_18493);
or U18667 (N_18667,N_18462,N_18495);
and U18668 (N_18668,N_18587,N_18563);
or U18669 (N_18669,N_18520,N_18455);
nand U18670 (N_18670,N_18536,N_18588);
nor U18671 (N_18671,N_18571,N_18473);
nor U18672 (N_18672,N_18506,N_18566);
xnor U18673 (N_18673,N_18564,N_18405);
nand U18674 (N_18674,N_18586,N_18535);
and U18675 (N_18675,N_18584,N_18570);
and U18676 (N_18676,N_18568,N_18527);
nand U18677 (N_18677,N_18550,N_18407);
or U18678 (N_18678,N_18537,N_18411);
or U18679 (N_18679,N_18583,N_18486);
nor U18680 (N_18680,N_18438,N_18591);
or U18681 (N_18681,N_18434,N_18457);
and U18682 (N_18682,N_18559,N_18476);
nor U18683 (N_18683,N_18460,N_18512);
nor U18684 (N_18684,N_18439,N_18408);
and U18685 (N_18685,N_18542,N_18508);
or U18686 (N_18686,N_18427,N_18577);
nand U18687 (N_18687,N_18532,N_18466);
nand U18688 (N_18688,N_18505,N_18541);
nand U18689 (N_18689,N_18433,N_18526);
or U18690 (N_18690,N_18595,N_18478);
nand U18691 (N_18691,N_18545,N_18528);
xnor U18692 (N_18692,N_18475,N_18483);
or U18693 (N_18693,N_18415,N_18451);
and U18694 (N_18694,N_18496,N_18467);
nor U18695 (N_18695,N_18580,N_18582);
nand U18696 (N_18696,N_18598,N_18497);
nor U18697 (N_18697,N_18557,N_18488);
and U18698 (N_18698,N_18441,N_18424);
and U18699 (N_18699,N_18519,N_18511);
nand U18700 (N_18700,N_18462,N_18569);
nor U18701 (N_18701,N_18485,N_18525);
nor U18702 (N_18702,N_18557,N_18594);
and U18703 (N_18703,N_18420,N_18443);
nor U18704 (N_18704,N_18592,N_18500);
nand U18705 (N_18705,N_18491,N_18592);
nor U18706 (N_18706,N_18543,N_18549);
xor U18707 (N_18707,N_18450,N_18479);
nor U18708 (N_18708,N_18490,N_18565);
nor U18709 (N_18709,N_18537,N_18568);
or U18710 (N_18710,N_18465,N_18507);
nand U18711 (N_18711,N_18514,N_18582);
or U18712 (N_18712,N_18459,N_18503);
or U18713 (N_18713,N_18528,N_18432);
nor U18714 (N_18714,N_18526,N_18478);
nor U18715 (N_18715,N_18478,N_18529);
or U18716 (N_18716,N_18514,N_18591);
nand U18717 (N_18717,N_18401,N_18462);
nand U18718 (N_18718,N_18415,N_18544);
and U18719 (N_18719,N_18489,N_18403);
or U18720 (N_18720,N_18556,N_18550);
nor U18721 (N_18721,N_18595,N_18522);
or U18722 (N_18722,N_18572,N_18494);
and U18723 (N_18723,N_18551,N_18404);
and U18724 (N_18724,N_18581,N_18478);
nand U18725 (N_18725,N_18489,N_18537);
nor U18726 (N_18726,N_18553,N_18494);
nand U18727 (N_18727,N_18417,N_18459);
nand U18728 (N_18728,N_18411,N_18498);
nor U18729 (N_18729,N_18519,N_18407);
and U18730 (N_18730,N_18598,N_18555);
nand U18731 (N_18731,N_18555,N_18483);
nand U18732 (N_18732,N_18446,N_18465);
nor U18733 (N_18733,N_18460,N_18449);
or U18734 (N_18734,N_18552,N_18468);
xor U18735 (N_18735,N_18576,N_18508);
nor U18736 (N_18736,N_18432,N_18411);
nand U18737 (N_18737,N_18497,N_18471);
nor U18738 (N_18738,N_18595,N_18581);
nor U18739 (N_18739,N_18501,N_18463);
and U18740 (N_18740,N_18503,N_18589);
nor U18741 (N_18741,N_18478,N_18448);
nand U18742 (N_18742,N_18558,N_18548);
and U18743 (N_18743,N_18425,N_18576);
or U18744 (N_18744,N_18513,N_18461);
and U18745 (N_18745,N_18588,N_18464);
and U18746 (N_18746,N_18525,N_18470);
or U18747 (N_18747,N_18529,N_18536);
and U18748 (N_18748,N_18571,N_18458);
or U18749 (N_18749,N_18433,N_18557);
and U18750 (N_18750,N_18596,N_18559);
and U18751 (N_18751,N_18414,N_18582);
nand U18752 (N_18752,N_18446,N_18478);
or U18753 (N_18753,N_18468,N_18402);
and U18754 (N_18754,N_18565,N_18463);
nor U18755 (N_18755,N_18426,N_18412);
and U18756 (N_18756,N_18414,N_18522);
and U18757 (N_18757,N_18578,N_18486);
nor U18758 (N_18758,N_18583,N_18484);
nor U18759 (N_18759,N_18502,N_18401);
nand U18760 (N_18760,N_18400,N_18553);
nand U18761 (N_18761,N_18539,N_18516);
nor U18762 (N_18762,N_18411,N_18592);
nor U18763 (N_18763,N_18559,N_18439);
nor U18764 (N_18764,N_18424,N_18504);
and U18765 (N_18765,N_18549,N_18401);
nor U18766 (N_18766,N_18589,N_18461);
nand U18767 (N_18767,N_18511,N_18504);
or U18768 (N_18768,N_18431,N_18429);
or U18769 (N_18769,N_18450,N_18549);
and U18770 (N_18770,N_18548,N_18471);
or U18771 (N_18771,N_18573,N_18506);
and U18772 (N_18772,N_18474,N_18599);
and U18773 (N_18773,N_18436,N_18485);
or U18774 (N_18774,N_18431,N_18515);
nor U18775 (N_18775,N_18515,N_18497);
nand U18776 (N_18776,N_18576,N_18448);
and U18777 (N_18777,N_18492,N_18509);
or U18778 (N_18778,N_18510,N_18483);
and U18779 (N_18779,N_18506,N_18479);
nand U18780 (N_18780,N_18494,N_18423);
or U18781 (N_18781,N_18517,N_18440);
or U18782 (N_18782,N_18419,N_18406);
and U18783 (N_18783,N_18588,N_18546);
nor U18784 (N_18784,N_18487,N_18542);
nand U18785 (N_18785,N_18520,N_18522);
or U18786 (N_18786,N_18436,N_18506);
and U18787 (N_18787,N_18528,N_18429);
and U18788 (N_18788,N_18577,N_18451);
nand U18789 (N_18789,N_18438,N_18580);
nor U18790 (N_18790,N_18543,N_18490);
or U18791 (N_18791,N_18418,N_18550);
and U18792 (N_18792,N_18502,N_18508);
or U18793 (N_18793,N_18572,N_18569);
nor U18794 (N_18794,N_18415,N_18418);
nor U18795 (N_18795,N_18511,N_18466);
or U18796 (N_18796,N_18547,N_18428);
nand U18797 (N_18797,N_18483,N_18459);
or U18798 (N_18798,N_18545,N_18558);
or U18799 (N_18799,N_18596,N_18419);
and U18800 (N_18800,N_18685,N_18631);
nand U18801 (N_18801,N_18665,N_18797);
and U18802 (N_18802,N_18681,N_18611);
nand U18803 (N_18803,N_18799,N_18738);
nand U18804 (N_18804,N_18645,N_18750);
nand U18805 (N_18805,N_18709,N_18766);
and U18806 (N_18806,N_18615,N_18668);
or U18807 (N_18807,N_18635,N_18722);
nand U18808 (N_18808,N_18667,N_18654);
or U18809 (N_18809,N_18632,N_18680);
nand U18810 (N_18810,N_18623,N_18693);
and U18811 (N_18811,N_18794,N_18741);
nand U18812 (N_18812,N_18637,N_18703);
and U18813 (N_18813,N_18776,N_18661);
or U18814 (N_18814,N_18716,N_18610);
nor U18815 (N_18815,N_18713,N_18727);
nand U18816 (N_18816,N_18639,N_18760);
nand U18817 (N_18817,N_18790,N_18763);
or U18818 (N_18818,N_18717,N_18644);
nand U18819 (N_18819,N_18748,N_18715);
nor U18820 (N_18820,N_18793,N_18612);
nor U18821 (N_18821,N_18744,N_18636);
nand U18822 (N_18822,N_18792,N_18652);
nand U18823 (N_18823,N_18777,N_18755);
and U18824 (N_18824,N_18603,N_18704);
nand U18825 (N_18825,N_18616,N_18607);
nand U18826 (N_18826,N_18735,N_18779);
or U18827 (N_18827,N_18706,N_18682);
and U18828 (N_18828,N_18745,N_18698);
nor U18829 (N_18829,N_18786,N_18729);
nand U18830 (N_18830,N_18768,N_18638);
nor U18831 (N_18831,N_18605,N_18740);
nand U18832 (N_18832,N_18702,N_18630);
or U18833 (N_18833,N_18769,N_18624);
xor U18834 (N_18834,N_18718,N_18604);
nor U18835 (N_18835,N_18778,N_18707);
nand U18836 (N_18836,N_18601,N_18684);
nand U18837 (N_18837,N_18772,N_18697);
or U18838 (N_18838,N_18765,N_18640);
nor U18839 (N_18839,N_18730,N_18747);
nor U18840 (N_18840,N_18619,N_18686);
nand U18841 (N_18841,N_18659,N_18660);
and U18842 (N_18842,N_18737,N_18771);
or U18843 (N_18843,N_18666,N_18758);
and U18844 (N_18844,N_18609,N_18731);
nor U18845 (N_18845,N_18663,N_18699);
or U18846 (N_18846,N_18627,N_18618);
or U18847 (N_18847,N_18648,N_18711);
or U18848 (N_18848,N_18764,N_18724);
or U18849 (N_18849,N_18798,N_18783);
nand U18850 (N_18850,N_18762,N_18708);
and U18851 (N_18851,N_18678,N_18608);
and U18852 (N_18852,N_18787,N_18677);
or U18853 (N_18853,N_18626,N_18761);
nand U18854 (N_18854,N_18683,N_18710);
nor U18855 (N_18855,N_18617,N_18705);
or U18856 (N_18856,N_18655,N_18628);
and U18857 (N_18857,N_18767,N_18620);
and U18858 (N_18858,N_18700,N_18679);
nand U18859 (N_18859,N_18657,N_18753);
nand U18860 (N_18860,N_18791,N_18796);
nand U18861 (N_18861,N_18746,N_18734);
and U18862 (N_18862,N_18651,N_18725);
and U18863 (N_18863,N_18642,N_18614);
and U18864 (N_18864,N_18742,N_18712);
nor U18865 (N_18865,N_18784,N_18774);
nor U18866 (N_18866,N_18795,N_18739);
xnor U18867 (N_18867,N_18775,N_18752);
nor U18868 (N_18868,N_18650,N_18600);
and U18869 (N_18869,N_18692,N_18656);
and U18870 (N_18870,N_18641,N_18749);
nor U18871 (N_18871,N_18613,N_18723);
and U18872 (N_18872,N_18728,N_18714);
or U18873 (N_18873,N_18751,N_18633);
or U18874 (N_18874,N_18754,N_18647);
or U18875 (N_18875,N_18743,N_18653);
xnor U18876 (N_18876,N_18675,N_18643);
or U18877 (N_18877,N_18646,N_18780);
nand U18878 (N_18878,N_18672,N_18756);
nand U18879 (N_18879,N_18658,N_18759);
and U18880 (N_18880,N_18669,N_18721);
and U18881 (N_18881,N_18625,N_18689);
nor U18882 (N_18882,N_18662,N_18736);
or U18883 (N_18883,N_18732,N_18785);
nor U18884 (N_18884,N_18757,N_18719);
nand U18885 (N_18885,N_18634,N_18694);
nand U18886 (N_18886,N_18781,N_18688);
and U18887 (N_18887,N_18701,N_18674);
or U18888 (N_18888,N_18782,N_18691);
or U18889 (N_18889,N_18602,N_18788);
or U18890 (N_18890,N_18670,N_18621);
and U18891 (N_18891,N_18726,N_18733);
and U18892 (N_18892,N_18770,N_18696);
nand U18893 (N_18893,N_18687,N_18664);
or U18894 (N_18894,N_18606,N_18676);
or U18895 (N_18895,N_18773,N_18622);
nand U18896 (N_18896,N_18649,N_18789);
nand U18897 (N_18897,N_18695,N_18629);
nand U18898 (N_18898,N_18671,N_18690);
nor U18899 (N_18899,N_18720,N_18673);
nand U18900 (N_18900,N_18705,N_18664);
or U18901 (N_18901,N_18776,N_18705);
nor U18902 (N_18902,N_18618,N_18698);
nand U18903 (N_18903,N_18609,N_18651);
nor U18904 (N_18904,N_18600,N_18612);
or U18905 (N_18905,N_18745,N_18692);
nand U18906 (N_18906,N_18787,N_18721);
or U18907 (N_18907,N_18745,N_18718);
nand U18908 (N_18908,N_18638,N_18663);
nor U18909 (N_18909,N_18679,N_18770);
nor U18910 (N_18910,N_18611,N_18661);
and U18911 (N_18911,N_18744,N_18637);
nand U18912 (N_18912,N_18723,N_18728);
nor U18913 (N_18913,N_18710,N_18612);
nor U18914 (N_18914,N_18715,N_18754);
nand U18915 (N_18915,N_18630,N_18668);
and U18916 (N_18916,N_18618,N_18759);
or U18917 (N_18917,N_18753,N_18666);
and U18918 (N_18918,N_18614,N_18629);
nor U18919 (N_18919,N_18691,N_18675);
or U18920 (N_18920,N_18780,N_18656);
nor U18921 (N_18921,N_18744,N_18770);
and U18922 (N_18922,N_18694,N_18606);
or U18923 (N_18923,N_18617,N_18753);
nand U18924 (N_18924,N_18631,N_18617);
or U18925 (N_18925,N_18612,N_18604);
or U18926 (N_18926,N_18754,N_18747);
and U18927 (N_18927,N_18702,N_18716);
or U18928 (N_18928,N_18668,N_18758);
and U18929 (N_18929,N_18643,N_18683);
nand U18930 (N_18930,N_18758,N_18664);
nor U18931 (N_18931,N_18626,N_18647);
or U18932 (N_18932,N_18741,N_18764);
nor U18933 (N_18933,N_18673,N_18625);
nand U18934 (N_18934,N_18736,N_18699);
and U18935 (N_18935,N_18648,N_18608);
nor U18936 (N_18936,N_18792,N_18722);
and U18937 (N_18937,N_18761,N_18766);
nand U18938 (N_18938,N_18649,N_18776);
nor U18939 (N_18939,N_18770,N_18721);
or U18940 (N_18940,N_18646,N_18796);
and U18941 (N_18941,N_18620,N_18784);
or U18942 (N_18942,N_18668,N_18656);
nor U18943 (N_18943,N_18728,N_18761);
or U18944 (N_18944,N_18606,N_18716);
and U18945 (N_18945,N_18769,N_18774);
or U18946 (N_18946,N_18783,N_18699);
nor U18947 (N_18947,N_18623,N_18648);
or U18948 (N_18948,N_18750,N_18753);
and U18949 (N_18949,N_18747,N_18779);
nand U18950 (N_18950,N_18690,N_18760);
nand U18951 (N_18951,N_18729,N_18617);
nor U18952 (N_18952,N_18645,N_18772);
nor U18953 (N_18953,N_18607,N_18710);
nor U18954 (N_18954,N_18608,N_18643);
or U18955 (N_18955,N_18631,N_18751);
and U18956 (N_18956,N_18684,N_18765);
or U18957 (N_18957,N_18608,N_18744);
and U18958 (N_18958,N_18770,N_18789);
or U18959 (N_18959,N_18725,N_18716);
nand U18960 (N_18960,N_18625,N_18721);
nand U18961 (N_18961,N_18715,N_18707);
and U18962 (N_18962,N_18601,N_18673);
or U18963 (N_18963,N_18776,N_18700);
and U18964 (N_18964,N_18645,N_18605);
nand U18965 (N_18965,N_18626,N_18693);
nand U18966 (N_18966,N_18680,N_18685);
and U18967 (N_18967,N_18688,N_18763);
and U18968 (N_18968,N_18695,N_18785);
or U18969 (N_18969,N_18732,N_18625);
nand U18970 (N_18970,N_18717,N_18686);
or U18971 (N_18971,N_18799,N_18724);
nor U18972 (N_18972,N_18670,N_18738);
nand U18973 (N_18973,N_18715,N_18724);
or U18974 (N_18974,N_18600,N_18736);
and U18975 (N_18975,N_18643,N_18621);
or U18976 (N_18976,N_18788,N_18687);
nor U18977 (N_18977,N_18788,N_18745);
nor U18978 (N_18978,N_18781,N_18720);
nand U18979 (N_18979,N_18612,N_18734);
and U18980 (N_18980,N_18781,N_18641);
nor U18981 (N_18981,N_18740,N_18623);
or U18982 (N_18982,N_18738,N_18792);
nor U18983 (N_18983,N_18799,N_18731);
and U18984 (N_18984,N_18644,N_18674);
and U18985 (N_18985,N_18706,N_18614);
or U18986 (N_18986,N_18736,N_18664);
nand U18987 (N_18987,N_18766,N_18613);
nand U18988 (N_18988,N_18771,N_18724);
nand U18989 (N_18989,N_18726,N_18761);
nand U18990 (N_18990,N_18704,N_18717);
or U18991 (N_18991,N_18713,N_18791);
nand U18992 (N_18992,N_18795,N_18695);
nand U18993 (N_18993,N_18745,N_18626);
xor U18994 (N_18994,N_18799,N_18640);
or U18995 (N_18995,N_18707,N_18687);
nand U18996 (N_18996,N_18620,N_18668);
or U18997 (N_18997,N_18728,N_18633);
nor U18998 (N_18998,N_18675,N_18757);
or U18999 (N_18999,N_18709,N_18677);
xor U19000 (N_19000,N_18951,N_18993);
nand U19001 (N_19001,N_18939,N_18895);
and U19002 (N_19002,N_18904,N_18845);
nand U19003 (N_19003,N_18958,N_18956);
nor U19004 (N_19004,N_18924,N_18852);
nand U19005 (N_19005,N_18869,N_18960);
nor U19006 (N_19006,N_18982,N_18827);
or U19007 (N_19007,N_18806,N_18955);
nor U19008 (N_19008,N_18944,N_18810);
or U19009 (N_19009,N_18882,N_18858);
or U19010 (N_19010,N_18971,N_18844);
nand U19011 (N_19011,N_18866,N_18973);
and U19012 (N_19012,N_18945,N_18848);
or U19013 (N_19013,N_18921,N_18991);
and U19014 (N_19014,N_18879,N_18830);
nand U19015 (N_19015,N_18872,N_18861);
or U19016 (N_19016,N_18963,N_18829);
and U19017 (N_19017,N_18930,N_18822);
xor U19018 (N_19018,N_18820,N_18984);
or U19019 (N_19019,N_18851,N_18906);
and U19020 (N_19020,N_18868,N_18957);
nand U19021 (N_19021,N_18886,N_18997);
nand U19022 (N_19022,N_18938,N_18880);
nand U19023 (N_19023,N_18913,N_18846);
and U19024 (N_19024,N_18950,N_18855);
or U19025 (N_19025,N_18853,N_18987);
or U19026 (N_19026,N_18926,N_18874);
nor U19027 (N_19027,N_18899,N_18915);
and U19028 (N_19028,N_18969,N_18877);
nor U19029 (N_19029,N_18940,N_18870);
nor U19030 (N_19030,N_18812,N_18917);
nand U19031 (N_19031,N_18922,N_18834);
or U19032 (N_19032,N_18936,N_18994);
nand U19033 (N_19033,N_18892,N_18875);
nand U19034 (N_19034,N_18989,N_18811);
nand U19035 (N_19035,N_18948,N_18954);
nand U19036 (N_19036,N_18802,N_18966);
nor U19037 (N_19037,N_18985,N_18801);
nor U19038 (N_19038,N_18932,N_18931);
or U19039 (N_19039,N_18967,N_18817);
and U19040 (N_19040,N_18813,N_18929);
and U19041 (N_19041,N_18975,N_18864);
or U19042 (N_19042,N_18857,N_18839);
and U19043 (N_19043,N_18981,N_18900);
nor U19044 (N_19044,N_18964,N_18953);
nand U19045 (N_19045,N_18952,N_18998);
and U19046 (N_19046,N_18933,N_18891);
nor U19047 (N_19047,N_18901,N_18808);
or U19048 (N_19048,N_18972,N_18934);
or U19049 (N_19049,N_18821,N_18884);
and U19050 (N_19050,N_18837,N_18843);
nor U19051 (N_19051,N_18878,N_18867);
nor U19052 (N_19052,N_18842,N_18840);
nand U19053 (N_19053,N_18847,N_18961);
nor U19054 (N_19054,N_18909,N_18873);
or U19055 (N_19055,N_18863,N_18977);
nor U19056 (N_19056,N_18941,N_18907);
and U19057 (N_19057,N_18831,N_18974);
nand U19058 (N_19058,N_18928,N_18800);
and U19059 (N_19059,N_18947,N_18916);
and U19060 (N_19060,N_18894,N_18980);
nand U19061 (N_19061,N_18949,N_18914);
nand U19062 (N_19062,N_18912,N_18856);
or U19063 (N_19063,N_18807,N_18908);
nand U19064 (N_19064,N_18920,N_18942);
or U19065 (N_19065,N_18819,N_18816);
nor U19066 (N_19066,N_18897,N_18978);
nand U19067 (N_19067,N_18903,N_18890);
nand U19068 (N_19068,N_18832,N_18988);
nor U19069 (N_19069,N_18825,N_18970);
and U19070 (N_19070,N_18996,N_18905);
nand U19071 (N_19071,N_18881,N_18809);
and U19072 (N_19072,N_18946,N_18818);
nand U19073 (N_19073,N_18871,N_18992);
nand U19074 (N_19074,N_18910,N_18876);
nand U19075 (N_19075,N_18889,N_18862);
nand U19076 (N_19076,N_18911,N_18865);
nor U19077 (N_19077,N_18918,N_18824);
and U19078 (N_19078,N_18990,N_18887);
nand U19079 (N_19079,N_18896,N_18841);
nor U19080 (N_19080,N_18925,N_18962);
and U19081 (N_19081,N_18823,N_18836);
nor U19082 (N_19082,N_18923,N_18883);
and U19083 (N_19083,N_18898,N_18999);
and U19084 (N_19084,N_18919,N_18927);
nor U19085 (N_19085,N_18943,N_18833);
nand U19086 (N_19086,N_18976,N_18835);
or U19087 (N_19087,N_18854,N_18959);
nand U19088 (N_19088,N_18965,N_18986);
or U19089 (N_19089,N_18968,N_18902);
or U19090 (N_19090,N_18893,N_18935);
nand U19091 (N_19091,N_18859,N_18814);
nor U19092 (N_19092,N_18860,N_18850);
or U19093 (N_19093,N_18995,N_18838);
xnor U19094 (N_19094,N_18826,N_18888);
nor U19095 (N_19095,N_18828,N_18983);
and U19096 (N_19096,N_18979,N_18885);
or U19097 (N_19097,N_18815,N_18849);
and U19098 (N_19098,N_18805,N_18937);
nand U19099 (N_19099,N_18803,N_18804);
or U19100 (N_19100,N_18840,N_18977);
or U19101 (N_19101,N_18975,N_18843);
nand U19102 (N_19102,N_18933,N_18928);
nand U19103 (N_19103,N_18874,N_18958);
and U19104 (N_19104,N_18908,N_18920);
nor U19105 (N_19105,N_18922,N_18990);
or U19106 (N_19106,N_18836,N_18969);
nand U19107 (N_19107,N_18897,N_18963);
or U19108 (N_19108,N_18966,N_18964);
nor U19109 (N_19109,N_18804,N_18871);
nor U19110 (N_19110,N_18988,N_18956);
nand U19111 (N_19111,N_18912,N_18921);
nor U19112 (N_19112,N_18824,N_18809);
or U19113 (N_19113,N_18890,N_18918);
nand U19114 (N_19114,N_18971,N_18822);
or U19115 (N_19115,N_18963,N_18984);
or U19116 (N_19116,N_18950,N_18914);
nor U19117 (N_19117,N_18903,N_18929);
or U19118 (N_19118,N_18985,N_18963);
nor U19119 (N_19119,N_18973,N_18901);
nand U19120 (N_19120,N_18995,N_18946);
and U19121 (N_19121,N_18938,N_18877);
and U19122 (N_19122,N_18909,N_18949);
and U19123 (N_19123,N_18821,N_18829);
or U19124 (N_19124,N_18985,N_18845);
or U19125 (N_19125,N_18940,N_18819);
or U19126 (N_19126,N_18910,N_18810);
nand U19127 (N_19127,N_18895,N_18965);
and U19128 (N_19128,N_18984,N_18979);
and U19129 (N_19129,N_18809,N_18914);
or U19130 (N_19130,N_18909,N_18856);
and U19131 (N_19131,N_18886,N_18992);
nor U19132 (N_19132,N_18838,N_18993);
and U19133 (N_19133,N_18884,N_18816);
and U19134 (N_19134,N_18952,N_18903);
and U19135 (N_19135,N_18895,N_18887);
nand U19136 (N_19136,N_18993,N_18810);
or U19137 (N_19137,N_18962,N_18996);
nand U19138 (N_19138,N_18914,N_18909);
and U19139 (N_19139,N_18942,N_18946);
or U19140 (N_19140,N_18845,N_18851);
or U19141 (N_19141,N_18960,N_18827);
nor U19142 (N_19142,N_18800,N_18878);
or U19143 (N_19143,N_18816,N_18851);
or U19144 (N_19144,N_18882,N_18994);
or U19145 (N_19145,N_18830,N_18935);
nand U19146 (N_19146,N_18843,N_18821);
or U19147 (N_19147,N_18873,N_18828);
and U19148 (N_19148,N_18904,N_18918);
nand U19149 (N_19149,N_18894,N_18872);
or U19150 (N_19150,N_18830,N_18894);
nor U19151 (N_19151,N_18915,N_18886);
nor U19152 (N_19152,N_18819,N_18840);
or U19153 (N_19153,N_18913,N_18986);
nor U19154 (N_19154,N_18990,N_18949);
and U19155 (N_19155,N_18875,N_18866);
or U19156 (N_19156,N_18963,N_18880);
nand U19157 (N_19157,N_18998,N_18938);
and U19158 (N_19158,N_18842,N_18854);
or U19159 (N_19159,N_18886,N_18971);
or U19160 (N_19160,N_18933,N_18938);
nor U19161 (N_19161,N_18810,N_18815);
or U19162 (N_19162,N_18841,N_18907);
and U19163 (N_19163,N_18863,N_18906);
nor U19164 (N_19164,N_18971,N_18995);
and U19165 (N_19165,N_18832,N_18990);
and U19166 (N_19166,N_18891,N_18851);
or U19167 (N_19167,N_18987,N_18983);
nor U19168 (N_19168,N_18976,N_18807);
nor U19169 (N_19169,N_18855,N_18897);
and U19170 (N_19170,N_18970,N_18899);
and U19171 (N_19171,N_18916,N_18969);
nor U19172 (N_19172,N_18938,N_18847);
nor U19173 (N_19173,N_18891,N_18909);
nor U19174 (N_19174,N_18964,N_18967);
nand U19175 (N_19175,N_18831,N_18991);
nor U19176 (N_19176,N_18827,N_18923);
nor U19177 (N_19177,N_18847,N_18914);
nor U19178 (N_19178,N_18928,N_18984);
nor U19179 (N_19179,N_18892,N_18891);
or U19180 (N_19180,N_18878,N_18805);
and U19181 (N_19181,N_18984,N_18903);
nor U19182 (N_19182,N_18846,N_18911);
and U19183 (N_19183,N_18926,N_18875);
nor U19184 (N_19184,N_18992,N_18826);
or U19185 (N_19185,N_18955,N_18887);
and U19186 (N_19186,N_18994,N_18974);
nor U19187 (N_19187,N_18824,N_18901);
and U19188 (N_19188,N_18832,N_18899);
nor U19189 (N_19189,N_18813,N_18938);
or U19190 (N_19190,N_18929,N_18994);
nand U19191 (N_19191,N_18933,N_18973);
nand U19192 (N_19192,N_18928,N_18829);
nor U19193 (N_19193,N_18966,N_18876);
nand U19194 (N_19194,N_18818,N_18859);
and U19195 (N_19195,N_18955,N_18967);
and U19196 (N_19196,N_18970,N_18871);
or U19197 (N_19197,N_18917,N_18823);
nor U19198 (N_19198,N_18802,N_18804);
and U19199 (N_19199,N_18925,N_18856);
nor U19200 (N_19200,N_19197,N_19155);
nand U19201 (N_19201,N_19023,N_19083);
nand U19202 (N_19202,N_19071,N_19124);
and U19203 (N_19203,N_19118,N_19182);
or U19204 (N_19204,N_19077,N_19054);
and U19205 (N_19205,N_19151,N_19040);
nor U19206 (N_19206,N_19060,N_19089);
nor U19207 (N_19207,N_19165,N_19007);
or U19208 (N_19208,N_19114,N_19195);
and U19209 (N_19209,N_19048,N_19059);
nand U19210 (N_19210,N_19135,N_19075);
nor U19211 (N_19211,N_19061,N_19019);
nor U19212 (N_19212,N_19103,N_19171);
nor U19213 (N_19213,N_19084,N_19021);
or U19214 (N_19214,N_19009,N_19175);
nand U19215 (N_19215,N_19018,N_19126);
nor U19216 (N_19216,N_19157,N_19123);
nor U19217 (N_19217,N_19108,N_19092);
nand U19218 (N_19218,N_19022,N_19037);
or U19219 (N_19219,N_19193,N_19051);
nand U19220 (N_19220,N_19039,N_19082);
nand U19221 (N_19221,N_19131,N_19091);
nor U19222 (N_19222,N_19121,N_19035);
nor U19223 (N_19223,N_19189,N_19156);
or U19224 (N_19224,N_19130,N_19000);
or U19225 (N_19225,N_19183,N_19029);
nand U19226 (N_19226,N_19113,N_19145);
or U19227 (N_19227,N_19096,N_19172);
or U19228 (N_19228,N_19147,N_19167);
nand U19229 (N_19229,N_19105,N_19137);
or U19230 (N_19230,N_19134,N_19187);
and U19231 (N_19231,N_19170,N_19042);
and U19232 (N_19232,N_19120,N_19176);
or U19233 (N_19233,N_19033,N_19116);
nor U19234 (N_19234,N_19094,N_19179);
nor U19235 (N_19235,N_19140,N_19027);
nor U19236 (N_19236,N_19136,N_19138);
and U19237 (N_19237,N_19057,N_19196);
nand U19238 (N_19238,N_19072,N_19093);
or U19239 (N_19239,N_19199,N_19133);
nand U19240 (N_19240,N_19166,N_19177);
nand U19241 (N_19241,N_19034,N_19032);
or U19242 (N_19242,N_19122,N_19159);
or U19243 (N_19243,N_19086,N_19049);
nand U19244 (N_19244,N_19005,N_19050);
and U19245 (N_19245,N_19112,N_19044);
and U19246 (N_19246,N_19031,N_19064);
nand U19247 (N_19247,N_19181,N_19062);
nor U19248 (N_19248,N_19191,N_19160);
or U19249 (N_19249,N_19173,N_19192);
and U19250 (N_19250,N_19163,N_19041);
nor U19251 (N_19251,N_19106,N_19111);
or U19252 (N_19252,N_19168,N_19047);
nand U19253 (N_19253,N_19107,N_19017);
nand U19254 (N_19254,N_19098,N_19080);
or U19255 (N_19255,N_19067,N_19025);
nor U19256 (N_19256,N_19012,N_19078);
or U19257 (N_19257,N_19125,N_19014);
nor U19258 (N_19258,N_19081,N_19065);
nand U19259 (N_19259,N_19006,N_19198);
or U19260 (N_19260,N_19026,N_19178);
and U19261 (N_19261,N_19070,N_19119);
nand U19262 (N_19262,N_19164,N_19085);
or U19263 (N_19263,N_19194,N_19148);
or U19264 (N_19264,N_19004,N_19110);
and U19265 (N_19265,N_19028,N_19150);
or U19266 (N_19266,N_19190,N_19180);
and U19267 (N_19267,N_19141,N_19066);
nand U19268 (N_19268,N_19079,N_19127);
or U19269 (N_19269,N_19188,N_19045);
or U19270 (N_19270,N_19146,N_19153);
or U19271 (N_19271,N_19104,N_19088);
nor U19272 (N_19272,N_19008,N_19169);
or U19273 (N_19273,N_19011,N_19144);
nor U19274 (N_19274,N_19090,N_19016);
nor U19275 (N_19275,N_19158,N_19043);
and U19276 (N_19276,N_19149,N_19139);
or U19277 (N_19277,N_19046,N_19102);
or U19278 (N_19278,N_19087,N_19053);
nor U19279 (N_19279,N_19100,N_19015);
nand U19280 (N_19280,N_19013,N_19030);
and U19281 (N_19281,N_19010,N_19128);
or U19282 (N_19282,N_19052,N_19101);
nor U19283 (N_19283,N_19099,N_19117);
and U19284 (N_19284,N_19038,N_19132);
and U19285 (N_19285,N_19063,N_19056);
nand U19286 (N_19286,N_19058,N_19186);
nand U19287 (N_19287,N_19184,N_19069);
or U19288 (N_19288,N_19068,N_19115);
and U19289 (N_19289,N_19002,N_19152);
or U19290 (N_19290,N_19143,N_19097);
nor U19291 (N_19291,N_19129,N_19024);
nand U19292 (N_19292,N_19020,N_19161);
and U19293 (N_19293,N_19095,N_19073);
xnor U19294 (N_19294,N_19036,N_19074);
or U19295 (N_19295,N_19109,N_19003);
nor U19296 (N_19296,N_19076,N_19142);
nand U19297 (N_19297,N_19055,N_19174);
or U19298 (N_19298,N_19001,N_19154);
and U19299 (N_19299,N_19162,N_19185);
and U19300 (N_19300,N_19080,N_19181);
nand U19301 (N_19301,N_19016,N_19097);
nand U19302 (N_19302,N_19162,N_19081);
or U19303 (N_19303,N_19053,N_19146);
nand U19304 (N_19304,N_19109,N_19114);
or U19305 (N_19305,N_19179,N_19013);
nor U19306 (N_19306,N_19119,N_19127);
nand U19307 (N_19307,N_19145,N_19040);
and U19308 (N_19308,N_19031,N_19075);
and U19309 (N_19309,N_19143,N_19157);
or U19310 (N_19310,N_19144,N_19028);
nand U19311 (N_19311,N_19086,N_19092);
nand U19312 (N_19312,N_19138,N_19144);
nand U19313 (N_19313,N_19184,N_19172);
and U19314 (N_19314,N_19060,N_19006);
nor U19315 (N_19315,N_19082,N_19007);
nand U19316 (N_19316,N_19105,N_19194);
and U19317 (N_19317,N_19184,N_19133);
nor U19318 (N_19318,N_19057,N_19049);
or U19319 (N_19319,N_19067,N_19031);
nor U19320 (N_19320,N_19070,N_19141);
or U19321 (N_19321,N_19183,N_19053);
nand U19322 (N_19322,N_19075,N_19094);
nand U19323 (N_19323,N_19121,N_19167);
nor U19324 (N_19324,N_19059,N_19080);
nor U19325 (N_19325,N_19083,N_19166);
nand U19326 (N_19326,N_19019,N_19087);
nor U19327 (N_19327,N_19011,N_19044);
nand U19328 (N_19328,N_19122,N_19043);
nand U19329 (N_19329,N_19169,N_19096);
nor U19330 (N_19330,N_19033,N_19163);
xnor U19331 (N_19331,N_19009,N_19011);
and U19332 (N_19332,N_19030,N_19115);
nor U19333 (N_19333,N_19028,N_19185);
and U19334 (N_19334,N_19185,N_19108);
nor U19335 (N_19335,N_19130,N_19081);
nor U19336 (N_19336,N_19181,N_19063);
nand U19337 (N_19337,N_19016,N_19105);
or U19338 (N_19338,N_19081,N_19164);
nand U19339 (N_19339,N_19055,N_19092);
or U19340 (N_19340,N_19031,N_19011);
and U19341 (N_19341,N_19084,N_19185);
nand U19342 (N_19342,N_19055,N_19062);
nor U19343 (N_19343,N_19161,N_19056);
or U19344 (N_19344,N_19046,N_19166);
and U19345 (N_19345,N_19098,N_19154);
or U19346 (N_19346,N_19030,N_19191);
nand U19347 (N_19347,N_19048,N_19068);
nor U19348 (N_19348,N_19063,N_19060);
nor U19349 (N_19349,N_19056,N_19098);
nand U19350 (N_19350,N_19122,N_19044);
and U19351 (N_19351,N_19066,N_19007);
nand U19352 (N_19352,N_19095,N_19161);
nor U19353 (N_19353,N_19107,N_19166);
nor U19354 (N_19354,N_19096,N_19106);
nor U19355 (N_19355,N_19084,N_19049);
and U19356 (N_19356,N_19151,N_19012);
nand U19357 (N_19357,N_19011,N_19137);
nor U19358 (N_19358,N_19166,N_19172);
nand U19359 (N_19359,N_19099,N_19156);
and U19360 (N_19360,N_19128,N_19003);
or U19361 (N_19361,N_19127,N_19198);
and U19362 (N_19362,N_19026,N_19073);
nor U19363 (N_19363,N_19178,N_19115);
nand U19364 (N_19364,N_19025,N_19147);
nand U19365 (N_19365,N_19150,N_19049);
or U19366 (N_19366,N_19182,N_19149);
and U19367 (N_19367,N_19011,N_19118);
nor U19368 (N_19368,N_19143,N_19020);
and U19369 (N_19369,N_19174,N_19056);
nand U19370 (N_19370,N_19114,N_19074);
and U19371 (N_19371,N_19071,N_19175);
and U19372 (N_19372,N_19108,N_19022);
or U19373 (N_19373,N_19197,N_19008);
or U19374 (N_19374,N_19018,N_19127);
and U19375 (N_19375,N_19171,N_19059);
or U19376 (N_19376,N_19043,N_19114);
or U19377 (N_19377,N_19157,N_19009);
nor U19378 (N_19378,N_19109,N_19186);
and U19379 (N_19379,N_19168,N_19073);
nand U19380 (N_19380,N_19064,N_19184);
nor U19381 (N_19381,N_19159,N_19140);
and U19382 (N_19382,N_19114,N_19182);
nor U19383 (N_19383,N_19127,N_19066);
nand U19384 (N_19384,N_19153,N_19013);
nor U19385 (N_19385,N_19002,N_19177);
or U19386 (N_19386,N_19039,N_19067);
and U19387 (N_19387,N_19072,N_19105);
and U19388 (N_19388,N_19106,N_19167);
or U19389 (N_19389,N_19051,N_19151);
and U19390 (N_19390,N_19059,N_19023);
xnor U19391 (N_19391,N_19163,N_19192);
nand U19392 (N_19392,N_19112,N_19037);
nor U19393 (N_19393,N_19134,N_19188);
or U19394 (N_19394,N_19164,N_19151);
nand U19395 (N_19395,N_19056,N_19048);
nor U19396 (N_19396,N_19091,N_19024);
nand U19397 (N_19397,N_19059,N_19081);
nor U19398 (N_19398,N_19100,N_19189);
or U19399 (N_19399,N_19136,N_19026);
or U19400 (N_19400,N_19357,N_19323);
or U19401 (N_19401,N_19309,N_19388);
and U19402 (N_19402,N_19272,N_19392);
or U19403 (N_19403,N_19360,N_19335);
nand U19404 (N_19404,N_19206,N_19374);
nand U19405 (N_19405,N_19365,N_19297);
or U19406 (N_19406,N_19282,N_19203);
nor U19407 (N_19407,N_19338,N_19217);
or U19408 (N_19408,N_19271,N_19398);
nor U19409 (N_19409,N_19292,N_19351);
nand U19410 (N_19410,N_19300,N_19243);
xnor U19411 (N_19411,N_19332,N_19370);
nor U19412 (N_19412,N_19240,N_19210);
nand U19413 (N_19413,N_19298,N_19304);
nand U19414 (N_19414,N_19204,N_19220);
nor U19415 (N_19415,N_19399,N_19391);
nand U19416 (N_19416,N_19395,N_19228);
or U19417 (N_19417,N_19205,N_19285);
xnor U19418 (N_19418,N_19366,N_19222);
nor U19419 (N_19419,N_19382,N_19242);
nor U19420 (N_19420,N_19373,N_19287);
nor U19421 (N_19421,N_19266,N_19369);
and U19422 (N_19422,N_19384,N_19393);
or U19423 (N_19423,N_19302,N_19311);
nor U19424 (N_19424,N_19362,N_19371);
nand U19425 (N_19425,N_19284,N_19320);
or U19426 (N_19426,N_19264,N_19263);
nor U19427 (N_19427,N_19308,N_19315);
or U19428 (N_19428,N_19299,N_19232);
and U19429 (N_19429,N_19278,N_19231);
or U19430 (N_19430,N_19314,N_19303);
nor U19431 (N_19431,N_19295,N_19214);
nor U19432 (N_19432,N_19250,N_19313);
nor U19433 (N_19433,N_19239,N_19219);
nor U19434 (N_19434,N_19305,N_19229);
nor U19435 (N_19435,N_19353,N_19349);
nand U19436 (N_19436,N_19213,N_19248);
nor U19437 (N_19437,N_19241,N_19211);
and U19438 (N_19438,N_19318,N_19301);
nor U19439 (N_19439,N_19319,N_19346);
or U19440 (N_19440,N_19208,N_19316);
and U19441 (N_19441,N_19288,N_19277);
nand U19442 (N_19442,N_19380,N_19212);
and U19443 (N_19443,N_19201,N_19317);
and U19444 (N_19444,N_19330,N_19367);
nand U19445 (N_19445,N_19223,N_19363);
nor U19446 (N_19446,N_19251,N_19227);
nor U19447 (N_19447,N_19368,N_19356);
or U19448 (N_19448,N_19347,N_19236);
and U19449 (N_19449,N_19389,N_19269);
and U19450 (N_19450,N_19387,N_19336);
and U19451 (N_19451,N_19390,N_19234);
nand U19452 (N_19452,N_19247,N_19310);
nor U19453 (N_19453,N_19230,N_19255);
nor U19454 (N_19454,N_19257,N_19262);
or U19455 (N_19455,N_19396,N_19345);
nand U19456 (N_19456,N_19221,N_19326);
nand U19457 (N_19457,N_19215,N_19286);
or U19458 (N_19458,N_19274,N_19378);
or U19459 (N_19459,N_19273,N_19216);
nor U19460 (N_19460,N_19359,N_19394);
nand U19461 (N_19461,N_19361,N_19294);
and U19462 (N_19462,N_19265,N_19244);
or U19463 (N_19463,N_19275,N_19268);
or U19464 (N_19464,N_19253,N_19328);
nor U19465 (N_19465,N_19372,N_19276);
or U19466 (N_19466,N_19226,N_19267);
nor U19467 (N_19467,N_19377,N_19340);
nor U19468 (N_19468,N_19381,N_19337);
or U19469 (N_19469,N_19290,N_19348);
nand U19470 (N_19470,N_19209,N_19283);
or U19471 (N_19471,N_19296,N_19200);
and U19472 (N_19472,N_19280,N_19379);
nor U19473 (N_19473,N_19339,N_19306);
or U19474 (N_19474,N_19341,N_19261);
and U19475 (N_19475,N_19385,N_19343);
nor U19476 (N_19476,N_19342,N_19307);
nand U19477 (N_19477,N_19333,N_19355);
and U19478 (N_19478,N_19354,N_19324);
nor U19479 (N_19479,N_19270,N_19375);
or U19480 (N_19480,N_19224,N_19321);
or U19481 (N_19481,N_19238,N_19235);
nand U19482 (N_19482,N_19376,N_19252);
nand U19483 (N_19483,N_19256,N_19289);
and U19484 (N_19484,N_19325,N_19386);
and U19485 (N_19485,N_19344,N_19334);
nand U19486 (N_19486,N_19352,N_19329);
or U19487 (N_19487,N_19281,N_19383);
and U19488 (N_19488,N_19260,N_19245);
and U19489 (N_19489,N_19312,N_19233);
or U19490 (N_19490,N_19207,N_19291);
or U19491 (N_19491,N_19279,N_19322);
nand U19492 (N_19492,N_19254,N_19202);
nand U19493 (N_19493,N_19358,N_19327);
and U19494 (N_19494,N_19258,N_19293);
nand U19495 (N_19495,N_19331,N_19364);
or U19496 (N_19496,N_19246,N_19350);
nor U19497 (N_19497,N_19397,N_19259);
or U19498 (N_19498,N_19237,N_19249);
or U19499 (N_19499,N_19225,N_19218);
or U19500 (N_19500,N_19355,N_19397);
nor U19501 (N_19501,N_19363,N_19303);
nor U19502 (N_19502,N_19275,N_19233);
nor U19503 (N_19503,N_19280,N_19226);
or U19504 (N_19504,N_19370,N_19371);
nand U19505 (N_19505,N_19370,N_19310);
or U19506 (N_19506,N_19274,N_19299);
or U19507 (N_19507,N_19306,N_19303);
nand U19508 (N_19508,N_19262,N_19375);
or U19509 (N_19509,N_19324,N_19207);
and U19510 (N_19510,N_19216,N_19221);
nand U19511 (N_19511,N_19364,N_19356);
and U19512 (N_19512,N_19282,N_19345);
nand U19513 (N_19513,N_19211,N_19340);
or U19514 (N_19514,N_19331,N_19358);
nand U19515 (N_19515,N_19382,N_19282);
and U19516 (N_19516,N_19369,N_19247);
nor U19517 (N_19517,N_19327,N_19237);
or U19518 (N_19518,N_19373,N_19323);
or U19519 (N_19519,N_19264,N_19289);
or U19520 (N_19520,N_19381,N_19214);
and U19521 (N_19521,N_19200,N_19343);
and U19522 (N_19522,N_19235,N_19276);
nand U19523 (N_19523,N_19295,N_19300);
and U19524 (N_19524,N_19395,N_19301);
or U19525 (N_19525,N_19371,N_19276);
and U19526 (N_19526,N_19332,N_19298);
nor U19527 (N_19527,N_19306,N_19209);
nor U19528 (N_19528,N_19325,N_19327);
nand U19529 (N_19529,N_19360,N_19210);
nand U19530 (N_19530,N_19381,N_19278);
nor U19531 (N_19531,N_19320,N_19323);
nor U19532 (N_19532,N_19209,N_19290);
and U19533 (N_19533,N_19230,N_19398);
nor U19534 (N_19534,N_19380,N_19303);
nor U19535 (N_19535,N_19296,N_19290);
nor U19536 (N_19536,N_19363,N_19240);
or U19537 (N_19537,N_19308,N_19383);
or U19538 (N_19538,N_19262,N_19267);
nor U19539 (N_19539,N_19210,N_19364);
nand U19540 (N_19540,N_19336,N_19327);
nor U19541 (N_19541,N_19309,N_19354);
or U19542 (N_19542,N_19252,N_19222);
nor U19543 (N_19543,N_19287,N_19350);
or U19544 (N_19544,N_19253,N_19250);
and U19545 (N_19545,N_19288,N_19270);
or U19546 (N_19546,N_19291,N_19273);
nand U19547 (N_19547,N_19211,N_19206);
and U19548 (N_19548,N_19397,N_19292);
nor U19549 (N_19549,N_19220,N_19237);
and U19550 (N_19550,N_19370,N_19246);
nor U19551 (N_19551,N_19347,N_19232);
nor U19552 (N_19552,N_19388,N_19334);
nor U19553 (N_19553,N_19308,N_19268);
or U19554 (N_19554,N_19250,N_19342);
and U19555 (N_19555,N_19379,N_19278);
nand U19556 (N_19556,N_19326,N_19361);
and U19557 (N_19557,N_19368,N_19325);
or U19558 (N_19558,N_19357,N_19216);
nand U19559 (N_19559,N_19307,N_19363);
nand U19560 (N_19560,N_19210,N_19343);
nor U19561 (N_19561,N_19368,N_19308);
or U19562 (N_19562,N_19279,N_19395);
and U19563 (N_19563,N_19255,N_19239);
nand U19564 (N_19564,N_19260,N_19311);
nand U19565 (N_19565,N_19210,N_19267);
and U19566 (N_19566,N_19379,N_19315);
nor U19567 (N_19567,N_19386,N_19277);
nor U19568 (N_19568,N_19376,N_19216);
and U19569 (N_19569,N_19223,N_19347);
nor U19570 (N_19570,N_19354,N_19207);
and U19571 (N_19571,N_19217,N_19285);
or U19572 (N_19572,N_19263,N_19220);
or U19573 (N_19573,N_19331,N_19347);
nand U19574 (N_19574,N_19301,N_19327);
nor U19575 (N_19575,N_19286,N_19267);
or U19576 (N_19576,N_19314,N_19323);
and U19577 (N_19577,N_19204,N_19251);
nor U19578 (N_19578,N_19349,N_19221);
and U19579 (N_19579,N_19236,N_19289);
nor U19580 (N_19580,N_19361,N_19234);
or U19581 (N_19581,N_19376,N_19355);
nor U19582 (N_19582,N_19369,N_19326);
nor U19583 (N_19583,N_19227,N_19299);
nand U19584 (N_19584,N_19363,N_19388);
and U19585 (N_19585,N_19331,N_19301);
or U19586 (N_19586,N_19213,N_19276);
nand U19587 (N_19587,N_19224,N_19387);
or U19588 (N_19588,N_19210,N_19237);
or U19589 (N_19589,N_19295,N_19306);
and U19590 (N_19590,N_19277,N_19251);
nor U19591 (N_19591,N_19291,N_19235);
nand U19592 (N_19592,N_19276,N_19203);
or U19593 (N_19593,N_19236,N_19206);
nor U19594 (N_19594,N_19270,N_19234);
or U19595 (N_19595,N_19395,N_19319);
nand U19596 (N_19596,N_19232,N_19384);
nor U19597 (N_19597,N_19252,N_19272);
and U19598 (N_19598,N_19394,N_19237);
or U19599 (N_19599,N_19213,N_19204);
nand U19600 (N_19600,N_19476,N_19427);
nor U19601 (N_19601,N_19419,N_19429);
or U19602 (N_19602,N_19405,N_19411);
nor U19603 (N_19603,N_19408,N_19466);
or U19604 (N_19604,N_19410,N_19467);
nor U19605 (N_19605,N_19432,N_19531);
or U19606 (N_19606,N_19569,N_19453);
or U19607 (N_19607,N_19500,N_19479);
or U19608 (N_19608,N_19440,N_19480);
and U19609 (N_19609,N_19435,N_19527);
nor U19610 (N_19610,N_19556,N_19524);
nor U19611 (N_19611,N_19592,N_19469);
and U19612 (N_19612,N_19528,N_19497);
nand U19613 (N_19613,N_19523,N_19428);
nand U19614 (N_19614,N_19442,N_19406);
or U19615 (N_19615,N_19549,N_19543);
nor U19616 (N_19616,N_19544,N_19578);
or U19617 (N_19617,N_19594,N_19464);
and U19618 (N_19618,N_19548,N_19484);
and U19619 (N_19619,N_19417,N_19489);
nor U19620 (N_19620,N_19590,N_19572);
nor U19621 (N_19621,N_19584,N_19552);
or U19622 (N_19622,N_19533,N_19538);
nand U19623 (N_19623,N_19449,N_19424);
nand U19624 (N_19624,N_19537,N_19474);
nor U19625 (N_19625,N_19542,N_19456);
or U19626 (N_19626,N_19502,N_19468);
and U19627 (N_19627,N_19444,N_19501);
nor U19628 (N_19628,N_19526,N_19595);
and U19629 (N_19629,N_19460,N_19520);
xor U19630 (N_19630,N_19496,N_19522);
and U19631 (N_19631,N_19525,N_19512);
nand U19632 (N_19632,N_19492,N_19498);
nor U19633 (N_19633,N_19562,N_19452);
or U19634 (N_19634,N_19530,N_19482);
xnor U19635 (N_19635,N_19493,N_19439);
and U19636 (N_19636,N_19574,N_19521);
or U19637 (N_19637,N_19515,N_19506);
and U19638 (N_19638,N_19553,N_19458);
or U19639 (N_19639,N_19471,N_19588);
and U19640 (N_19640,N_19573,N_19407);
or U19641 (N_19641,N_19483,N_19475);
nor U19642 (N_19642,N_19566,N_19580);
and U19643 (N_19643,N_19599,N_19504);
and U19644 (N_19644,N_19462,N_19490);
and U19645 (N_19645,N_19536,N_19532);
nand U19646 (N_19646,N_19447,N_19455);
and U19647 (N_19647,N_19583,N_19400);
nand U19648 (N_19648,N_19454,N_19461);
and U19649 (N_19649,N_19423,N_19582);
or U19650 (N_19650,N_19593,N_19567);
and U19651 (N_19651,N_19403,N_19494);
and U19652 (N_19652,N_19575,N_19422);
or U19653 (N_19653,N_19414,N_19441);
nor U19654 (N_19654,N_19518,N_19491);
and U19655 (N_19655,N_19517,N_19557);
nor U19656 (N_19656,N_19431,N_19465);
or U19657 (N_19657,N_19534,N_19418);
xor U19658 (N_19658,N_19587,N_19508);
and U19659 (N_19659,N_19499,N_19409);
nor U19660 (N_19660,N_19473,N_19412);
and U19661 (N_19661,N_19510,N_19563);
and U19662 (N_19662,N_19540,N_19433);
nor U19663 (N_19663,N_19436,N_19558);
and U19664 (N_19664,N_19535,N_19519);
and U19665 (N_19665,N_19568,N_19564);
nand U19666 (N_19666,N_19488,N_19416);
nand U19667 (N_19667,N_19434,N_19457);
and U19668 (N_19668,N_19486,N_19514);
nand U19669 (N_19669,N_19560,N_19463);
nand U19670 (N_19670,N_19547,N_19529);
and U19671 (N_19671,N_19551,N_19413);
or U19672 (N_19672,N_19404,N_19445);
or U19673 (N_19673,N_19443,N_19545);
or U19674 (N_19674,N_19425,N_19585);
nor U19675 (N_19675,N_19546,N_19507);
and U19676 (N_19676,N_19470,N_19511);
nor U19677 (N_19677,N_19550,N_19415);
nor U19678 (N_19678,N_19487,N_19451);
or U19679 (N_19679,N_19450,N_19561);
or U19680 (N_19680,N_19426,N_19586);
and U19681 (N_19681,N_19555,N_19420);
nor U19682 (N_19682,N_19513,N_19598);
nor U19683 (N_19683,N_19589,N_19430);
nor U19684 (N_19684,N_19577,N_19571);
nor U19685 (N_19685,N_19472,N_19597);
nand U19686 (N_19686,N_19541,N_19448);
xnor U19687 (N_19687,N_19576,N_19438);
or U19688 (N_19688,N_19579,N_19516);
or U19689 (N_19689,N_19477,N_19481);
nor U19690 (N_19690,N_19591,N_19459);
or U19691 (N_19691,N_19401,N_19437);
nor U19692 (N_19692,N_19509,N_19581);
nor U19693 (N_19693,N_19446,N_19596);
nand U19694 (N_19694,N_19505,N_19559);
or U19695 (N_19695,N_19554,N_19503);
nor U19696 (N_19696,N_19478,N_19539);
xor U19697 (N_19697,N_19421,N_19485);
and U19698 (N_19698,N_19570,N_19495);
nor U19699 (N_19699,N_19402,N_19565);
and U19700 (N_19700,N_19517,N_19504);
and U19701 (N_19701,N_19409,N_19476);
nand U19702 (N_19702,N_19584,N_19419);
and U19703 (N_19703,N_19590,N_19538);
and U19704 (N_19704,N_19466,N_19511);
nand U19705 (N_19705,N_19467,N_19501);
and U19706 (N_19706,N_19406,N_19508);
nand U19707 (N_19707,N_19581,N_19493);
nor U19708 (N_19708,N_19491,N_19481);
or U19709 (N_19709,N_19445,N_19454);
nand U19710 (N_19710,N_19558,N_19598);
nand U19711 (N_19711,N_19506,N_19594);
and U19712 (N_19712,N_19502,N_19432);
or U19713 (N_19713,N_19482,N_19443);
and U19714 (N_19714,N_19594,N_19567);
nor U19715 (N_19715,N_19417,N_19595);
nand U19716 (N_19716,N_19421,N_19491);
or U19717 (N_19717,N_19549,N_19402);
or U19718 (N_19718,N_19556,N_19566);
nor U19719 (N_19719,N_19464,N_19487);
or U19720 (N_19720,N_19598,N_19448);
or U19721 (N_19721,N_19487,N_19482);
nand U19722 (N_19722,N_19413,N_19488);
and U19723 (N_19723,N_19577,N_19459);
nor U19724 (N_19724,N_19459,N_19448);
nor U19725 (N_19725,N_19424,N_19412);
or U19726 (N_19726,N_19452,N_19404);
nand U19727 (N_19727,N_19518,N_19556);
and U19728 (N_19728,N_19558,N_19491);
or U19729 (N_19729,N_19555,N_19416);
and U19730 (N_19730,N_19530,N_19568);
and U19731 (N_19731,N_19573,N_19547);
nor U19732 (N_19732,N_19483,N_19521);
nand U19733 (N_19733,N_19490,N_19558);
and U19734 (N_19734,N_19524,N_19515);
nand U19735 (N_19735,N_19514,N_19584);
nor U19736 (N_19736,N_19510,N_19531);
or U19737 (N_19737,N_19464,N_19460);
nand U19738 (N_19738,N_19442,N_19541);
or U19739 (N_19739,N_19580,N_19456);
nand U19740 (N_19740,N_19422,N_19563);
or U19741 (N_19741,N_19446,N_19576);
or U19742 (N_19742,N_19534,N_19481);
nor U19743 (N_19743,N_19537,N_19541);
and U19744 (N_19744,N_19420,N_19594);
nor U19745 (N_19745,N_19434,N_19465);
nor U19746 (N_19746,N_19527,N_19543);
and U19747 (N_19747,N_19493,N_19520);
or U19748 (N_19748,N_19514,N_19511);
nand U19749 (N_19749,N_19424,N_19467);
nor U19750 (N_19750,N_19477,N_19580);
nor U19751 (N_19751,N_19532,N_19427);
nor U19752 (N_19752,N_19559,N_19595);
nor U19753 (N_19753,N_19525,N_19514);
xor U19754 (N_19754,N_19532,N_19505);
or U19755 (N_19755,N_19510,N_19404);
or U19756 (N_19756,N_19437,N_19452);
or U19757 (N_19757,N_19456,N_19596);
nor U19758 (N_19758,N_19559,N_19453);
nor U19759 (N_19759,N_19482,N_19423);
nand U19760 (N_19760,N_19477,N_19597);
and U19761 (N_19761,N_19585,N_19409);
and U19762 (N_19762,N_19597,N_19585);
or U19763 (N_19763,N_19444,N_19528);
nor U19764 (N_19764,N_19508,N_19471);
and U19765 (N_19765,N_19487,N_19495);
or U19766 (N_19766,N_19473,N_19559);
nor U19767 (N_19767,N_19401,N_19456);
nor U19768 (N_19768,N_19576,N_19479);
or U19769 (N_19769,N_19583,N_19409);
or U19770 (N_19770,N_19464,N_19453);
and U19771 (N_19771,N_19536,N_19422);
and U19772 (N_19772,N_19482,N_19493);
or U19773 (N_19773,N_19510,N_19529);
and U19774 (N_19774,N_19536,N_19486);
and U19775 (N_19775,N_19578,N_19434);
and U19776 (N_19776,N_19560,N_19431);
and U19777 (N_19777,N_19565,N_19536);
or U19778 (N_19778,N_19562,N_19419);
or U19779 (N_19779,N_19498,N_19548);
nor U19780 (N_19780,N_19507,N_19561);
or U19781 (N_19781,N_19491,N_19428);
and U19782 (N_19782,N_19528,N_19435);
nor U19783 (N_19783,N_19450,N_19440);
and U19784 (N_19784,N_19491,N_19454);
nand U19785 (N_19785,N_19430,N_19431);
and U19786 (N_19786,N_19510,N_19478);
nor U19787 (N_19787,N_19542,N_19472);
nand U19788 (N_19788,N_19574,N_19409);
nor U19789 (N_19789,N_19589,N_19493);
or U19790 (N_19790,N_19528,N_19483);
nand U19791 (N_19791,N_19570,N_19538);
or U19792 (N_19792,N_19428,N_19404);
nand U19793 (N_19793,N_19459,N_19473);
nand U19794 (N_19794,N_19515,N_19556);
or U19795 (N_19795,N_19561,N_19437);
nor U19796 (N_19796,N_19465,N_19568);
nor U19797 (N_19797,N_19467,N_19592);
nand U19798 (N_19798,N_19477,N_19400);
nand U19799 (N_19799,N_19438,N_19437);
nand U19800 (N_19800,N_19606,N_19769);
or U19801 (N_19801,N_19641,N_19630);
nand U19802 (N_19802,N_19620,N_19723);
and U19803 (N_19803,N_19777,N_19709);
nand U19804 (N_19804,N_19730,N_19706);
or U19805 (N_19805,N_19719,N_19711);
or U19806 (N_19806,N_19757,N_19629);
nor U19807 (N_19807,N_19790,N_19664);
or U19808 (N_19808,N_19604,N_19728);
nand U19809 (N_19809,N_19765,N_19619);
and U19810 (N_19810,N_19603,N_19639);
nor U19811 (N_19811,N_19694,N_19775);
nand U19812 (N_19812,N_19633,N_19774);
nand U19813 (N_19813,N_19667,N_19761);
and U19814 (N_19814,N_19725,N_19679);
nand U19815 (N_19815,N_19680,N_19672);
nor U19816 (N_19816,N_19759,N_19710);
or U19817 (N_19817,N_19707,N_19685);
nand U19818 (N_19818,N_19654,N_19754);
nand U19819 (N_19819,N_19767,N_19718);
or U19820 (N_19820,N_19651,N_19635);
or U19821 (N_19821,N_19677,N_19744);
and U19822 (N_19822,N_19722,N_19770);
and U19823 (N_19823,N_19780,N_19650);
nand U19824 (N_19824,N_19737,N_19632);
nand U19825 (N_19825,N_19657,N_19652);
and U19826 (N_19826,N_19787,N_19748);
nand U19827 (N_19827,N_19771,N_19640);
nor U19828 (N_19828,N_19613,N_19760);
or U19829 (N_19829,N_19683,N_19697);
nand U19830 (N_19830,N_19668,N_19624);
nor U19831 (N_19831,N_19681,N_19621);
or U19832 (N_19832,N_19691,N_19705);
or U19833 (N_19833,N_19782,N_19779);
and U19834 (N_19834,N_19669,N_19671);
and U19835 (N_19835,N_19716,N_19720);
or U19836 (N_19836,N_19623,N_19655);
and U19837 (N_19837,N_19773,N_19762);
nand U19838 (N_19838,N_19763,N_19628);
nor U19839 (N_19839,N_19721,N_19778);
or U19840 (N_19840,N_19605,N_19627);
nand U19841 (N_19841,N_19612,N_19643);
or U19842 (N_19842,N_19699,N_19766);
or U19843 (N_19843,N_19786,N_19638);
nand U19844 (N_19844,N_19740,N_19794);
nand U19845 (N_19845,N_19758,N_19739);
and U19846 (N_19846,N_19684,N_19653);
nand U19847 (N_19847,N_19648,N_19752);
nor U19848 (N_19848,N_19611,N_19665);
and U19849 (N_19849,N_19625,N_19663);
and U19850 (N_19850,N_19675,N_19749);
nor U19851 (N_19851,N_19676,N_19670);
and U19852 (N_19852,N_19726,N_19714);
nand U19853 (N_19853,N_19791,N_19674);
or U19854 (N_19854,N_19678,N_19713);
and U19855 (N_19855,N_19636,N_19702);
and U19856 (N_19856,N_19661,N_19626);
and U19857 (N_19857,N_19717,N_19736);
nor U19858 (N_19858,N_19634,N_19658);
nand U19859 (N_19859,N_19799,N_19729);
or U19860 (N_19860,N_19743,N_19733);
and U19861 (N_19861,N_19781,N_19637);
nand U19862 (N_19862,N_19755,N_19610);
nand U19863 (N_19863,N_19689,N_19768);
or U19864 (N_19864,N_19792,N_19789);
or U19865 (N_19865,N_19704,N_19693);
and U19866 (N_19866,N_19695,N_19798);
nand U19867 (N_19867,N_19647,N_19682);
nand U19868 (N_19868,N_19690,N_19631);
nor U19869 (N_19869,N_19642,N_19738);
nor U19870 (N_19870,N_19602,N_19724);
and U19871 (N_19871,N_19731,N_19646);
and U19872 (N_19872,N_19747,N_19700);
nand U19873 (N_19873,N_19764,N_19795);
or U19874 (N_19874,N_19735,N_19659);
nand U19875 (N_19875,N_19784,N_19715);
and U19876 (N_19876,N_19756,N_19607);
or U19877 (N_19877,N_19617,N_19796);
and U19878 (N_19878,N_19616,N_19696);
nand U19879 (N_19879,N_19666,N_19698);
or U19880 (N_19880,N_19753,N_19692);
nand U19881 (N_19881,N_19734,N_19797);
nand U19882 (N_19882,N_19673,N_19688);
and U19883 (N_19883,N_19622,N_19609);
nor U19884 (N_19884,N_19741,N_19732);
nand U19885 (N_19885,N_19742,N_19712);
and U19886 (N_19886,N_19708,N_19783);
nand U19887 (N_19887,N_19660,N_19776);
nor U19888 (N_19888,N_19656,N_19614);
or U19889 (N_19889,N_19751,N_19746);
or U19890 (N_19890,N_19750,N_19615);
and U19891 (N_19891,N_19745,N_19645);
nand U19892 (N_19892,N_19600,N_19703);
nand U19893 (N_19893,N_19727,N_19772);
or U19894 (N_19894,N_19793,N_19785);
nand U19895 (N_19895,N_19701,N_19649);
and U19896 (N_19896,N_19788,N_19618);
nor U19897 (N_19897,N_19662,N_19601);
or U19898 (N_19898,N_19687,N_19644);
or U19899 (N_19899,N_19608,N_19686);
nand U19900 (N_19900,N_19729,N_19614);
nand U19901 (N_19901,N_19683,N_19738);
nor U19902 (N_19902,N_19670,N_19671);
nor U19903 (N_19903,N_19601,N_19790);
nor U19904 (N_19904,N_19659,N_19654);
nor U19905 (N_19905,N_19700,N_19764);
nand U19906 (N_19906,N_19794,N_19788);
nand U19907 (N_19907,N_19691,N_19708);
nand U19908 (N_19908,N_19753,N_19799);
xor U19909 (N_19909,N_19698,N_19628);
nor U19910 (N_19910,N_19636,N_19788);
nor U19911 (N_19911,N_19751,N_19621);
nor U19912 (N_19912,N_19680,N_19734);
or U19913 (N_19913,N_19721,N_19792);
and U19914 (N_19914,N_19725,N_19658);
or U19915 (N_19915,N_19691,N_19672);
and U19916 (N_19916,N_19759,N_19617);
nand U19917 (N_19917,N_19795,N_19725);
nand U19918 (N_19918,N_19717,N_19700);
or U19919 (N_19919,N_19789,N_19791);
nor U19920 (N_19920,N_19716,N_19703);
and U19921 (N_19921,N_19631,N_19693);
or U19922 (N_19922,N_19661,N_19653);
nand U19923 (N_19923,N_19607,N_19692);
or U19924 (N_19924,N_19719,N_19635);
and U19925 (N_19925,N_19785,N_19733);
xnor U19926 (N_19926,N_19750,N_19644);
nor U19927 (N_19927,N_19641,N_19721);
nand U19928 (N_19928,N_19798,N_19643);
and U19929 (N_19929,N_19631,N_19731);
nor U19930 (N_19930,N_19705,N_19735);
and U19931 (N_19931,N_19745,N_19734);
and U19932 (N_19932,N_19740,N_19635);
nand U19933 (N_19933,N_19781,N_19679);
nor U19934 (N_19934,N_19787,N_19750);
nor U19935 (N_19935,N_19667,N_19699);
nor U19936 (N_19936,N_19681,N_19635);
and U19937 (N_19937,N_19690,N_19686);
and U19938 (N_19938,N_19799,N_19765);
nand U19939 (N_19939,N_19661,N_19632);
or U19940 (N_19940,N_19607,N_19616);
nand U19941 (N_19941,N_19728,N_19700);
nand U19942 (N_19942,N_19652,N_19638);
or U19943 (N_19943,N_19645,N_19770);
nand U19944 (N_19944,N_19666,N_19683);
nand U19945 (N_19945,N_19709,N_19685);
or U19946 (N_19946,N_19632,N_19735);
nor U19947 (N_19947,N_19675,N_19764);
or U19948 (N_19948,N_19651,N_19626);
and U19949 (N_19949,N_19670,N_19612);
nand U19950 (N_19950,N_19614,N_19674);
nor U19951 (N_19951,N_19704,N_19663);
nand U19952 (N_19952,N_19719,N_19657);
or U19953 (N_19953,N_19650,N_19686);
and U19954 (N_19954,N_19663,N_19679);
or U19955 (N_19955,N_19619,N_19616);
nand U19956 (N_19956,N_19647,N_19661);
and U19957 (N_19957,N_19708,N_19634);
or U19958 (N_19958,N_19610,N_19756);
nand U19959 (N_19959,N_19610,N_19795);
nor U19960 (N_19960,N_19703,N_19663);
nor U19961 (N_19961,N_19625,N_19614);
or U19962 (N_19962,N_19651,N_19663);
and U19963 (N_19963,N_19735,N_19620);
and U19964 (N_19964,N_19706,N_19645);
nor U19965 (N_19965,N_19775,N_19721);
and U19966 (N_19966,N_19681,N_19795);
xor U19967 (N_19967,N_19616,N_19769);
or U19968 (N_19968,N_19702,N_19648);
nand U19969 (N_19969,N_19734,N_19799);
nand U19970 (N_19970,N_19646,N_19783);
nand U19971 (N_19971,N_19753,N_19665);
and U19972 (N_19972,N_19747,N_19623);
nand U19973 (N_19973,N_19627,N_19680);
nand U19974 (N_19974,N_19725,N_19717);
and U19975 (N_19975,N_19713,N_19715);
nand U19976 (N_19976,N_19614,N_19697);
and U19977 (N_19977,N_19753,N_19663);
nor U19978 (N_19978,N_19719,N_19676);
nand U19979 (N_19979,N_19705,N_19716);
and U19980 (N_19980,N_19606,N_19641);
or U19981 (N_19981,N_19752,N_19716);
or U19982 (N_19982,N_19616,N_19645);
and U19983 (N_19983,N_19749,N_19690);
or U19984 (N_19984,N_19713,N_19704);
and U19985 (N_19985,N_19688,N_19659);
or U19986 (N_19986,N_19678,N_19645);
or U19987 (N_19987,N_19725,N_19633);
nor U19988 (N_19988,N_19711,N_19746);
and U19989 (N_19989,N_19649,N_19638);
nor U19990 (N_19990,N_19773,N_19781);
nor U19991 (N_19991,N_19737,N_19744);
and U19992 (N_19992,N_19654,N_19697);
nand U19993 (N_19993,N_19772,N_19746);
or U19994 (N_19994,N_19787,N_19620);
or U19995 (N_19995,N_19723,N_19770);
nor U19996 (N_19996,N_19760,N_19658);
nand U19997 (N_19997,N_19616,N_19743);
nand U19998 (N_19998,N_19704,N_19779);
nor U19999 (N_19999,N_19758,N_19644);
or U20000 (N_20000,N_19958,N_19965);
and U20001 (N_20001,N_19833,N_19894);
nor U20002 (N_20002,N_19966,N_19838);
or U20003 (N_20003,N_19898,N_19967);
and U20004 (N_20004,N_19982,N_19826);
nor U20005 (N_20005,N_19812,N_19872);
and U20006 (N_20006,N_19849,N_19910);
nor U20007 (N_20007,N_19928,N_19880);
or U20008 (N_20008,N_19996,N_19904);
or U20009 (N_20009,N_19953,N_19816);
and U20010 (N_20010,N_19808,N_19871);
nor U20011 (N_20011,N_19890,N_19860);
nor U20012 (N_20012,N_19825,N_19823);
and U20013 (N_20013,N_19807,N_19803);
nand U20014 (N_20014,N_19869,N_19886);
and U20015 (N_20015,N_19931,N_19964);
or U20016 (N_20016,N_19853,N_19915);
or U20017 (N_20017,N_19862,N_19804);
nor U20018 (N_20018,N_19989,N_19911);
or U20019 (N_20019,N_19882,N_19809);
and U20020 (N_20020,N_19839,N_19938);
nor U20021 (N_20021,N_19888,N_19828);
or U20022 (N_20022,N_19933,N_19935);
and U20023 (N_20023,N_19820,N_19829);
and U20024 (N_20024,N_19802,N_19857);
nand U20025 (N_20025,N_19929,N_19875);
nand U20026 (N_20026,N_19831,N_19902);
nand U20027 (N_20027,N_19856,N_19817);
or U20028 (N_20028,N_19845,N_19813);
nor U20029 (N_20029,N_19811,N_19979);
or U20030 (N_20030,N_19987,N_19976);
and U20031 (N_20031,N_19939,N_19969);
or U20032 (N_20032,N_19920,N_19879);
and U20033 (N_20033,N_19986,N_19995);
nor U20034 (N_20034,N_19892,N_19961);
or U20035 (N_20035,N_19924,N_19948);
or U20036 (N_20036,N_19973,N_19836);
or U20037 (N_20037,N_19889,N_19927);
and U20038 (N_20038,N_19909,N_19873);
nor U20039 (N_20039,N_19819,N_19992);
and U20040 (N_20040,N_19844,N_19918);
and U20041 (N_20041,N_19901,N_19952);
and U20042 (N_20042,N_19859,N_19868);
nor U20043 (N_20043,N_19994,N_19903);
or U20044 (N_20044,N_19821,N_19981);
nand U20045 (N_20045,N_19908,N_19876);
and U20046 (N_20046,N_19993,N_19887);
nor U20047 (N_20047,N_19858,N_19932);
nor U20048 (N_20048,N_19841,N_19930);
nand U20049 (N_20049,N_19801,N_19834);
nor U20050 (N_20050,N_19970,N_19891);
and U20051 (N_20051,N_19847,N_19960);
nand U20052 (N_20052,N_19865,N_19916);
or U20053 (N_20053,N_19878,N_19835);
or U20054 (N_20054,N_19944,N_19934);
nor U20055 (N_20055,N_19840,N_19925);
and U20056 (N_20056,N_19842,N_19963);
nand U20057 (N_20057,N_19863,N_19913);
nand U20058 (N_20058,N_19852,N_19955);
or U20059 (N_20059,N_19936,N_19814);
nand U20060 (N_20060,N_19824,N_19900);
or U20061 (N_20061,N_19980,N_19827);
or U20062 (N_20062,N_19943,N_19899);
nand U20063 (N_20063,N_19861,N_19956);
and U20064 (N_20064,N_19937,N_19850);
nor U20065 (N_20065,N_19884,N_19949);
and U20066 (N_20066,N_19972,N_19962);
or U20067 (N_20067,N_19805,N_19977);
or U20068 (N_20068,N_19957,N_19830);
nand U20069 (N_20069,N_19810,N_19974);
and U20070 (N_20070,N_19983,N_19907);
nor U20071 (N_20071,N_19855,N_19837);
and U20072 (N_20072,N_19941,N_19922);
and U20073 (N_20073,N_19870,N_19906);
nand U20074 (N_20074,N_19946,N_19999);
nor U20075 (N_20075,N_19893,N_19897);
nor U20076 (N_20076,N_19984,N_19971);
nor U20077 (N_20077,N_19951,N_19954);
nor U20078 (N_20078,N_19881,N_19945);
and U20079 (N_20079,N_19968,N_19998);
and U20080 (N_20080,N_19990,N_19806);
nand U20081 (N_20081,N_19926,N_19818);
and U20082 (N_20082,N_19896,N_19874);
and U20083 (N_20083,N_19988,N_19997);
nor U20084 (N_20084,N_19912,N_19877);
nor U20085 (N_20085,N_19917,N_19800);
nor U20086 (N_20086,N_19885,N_19867);
or U20087 (N_20087,N_19975,N_19959);
nand U20088 (N_20088,N_19851,N_19864);
or U20089 (N_20089,N_19947,N_19848);
nor U20090 (N_20090,N_19905,N_19815);
nor U20091 (N_20091,N_19854,N_19921);
and U20092 (N_20092,N_19883,N_19991);
nor U20093 (N_20093,N_19919,N_19832);
nand U20094 (N_20094,N_19822,N_19940);
nand U20095 (N_20095,N_19895,N_19846);
nor U20096 (N_20096,N_19843,N_19866);
nand U20097 (N_20097,N_19942,N_19923);
or U20098 (N_20098,N_19978,N_19950);
nand U20099 (N_20099,N_19914,N_19985);
nand U20100 (N_20100,N_19910,N_19895);
nor U20101 (N_20101,N_19882,N_19913);
nor U20102 (N_20102,N_19912,N_19986);
and U20103 (N_20103,N_19947,N_19833);
xnor U20104 (N_20104,N_19951,N_19825);
nor U20105 (N_20105,N_19918,N_19854);
and U20106 (N_20106,N_19925,N_19980);
or U20107 (N_20107,N_19960,N_19952);
nor U20108 (N_20108,N_19813,N_19805);
nor U20109 (N_20109,N_19993,N_19907);
nand U20110 (N_20110,N_19855,N_19948);
and U20111 (N_20111,N_19887,N_19972);
and U20112 (N_20112,N_19914,N_19958);
and U20113 (N_20113,N_19996,N_19989);
or U20114 (N_20114,N_19835,N_19907);
nor U20115 (N_20115,N_19808,N_19826);
or U20116 (N_20116,N_19939,N_19847);
or U20117 (N_20117,N_19821,N_19835);
and U20118 (N_20118,N_19932,N_19922);
nor U20119 (N_20119,N_19859,N_19822);
nor U20120 (N_20120,N_19971,N_19872);
and U20121 (N_20121,N_19834,N_19963);
and U20122 (N_20122,N_19832,N_19937);
and U20123 (N_20123,N_19817,N_19883);
or U20124 (N_20124,N_19825,N_19855);
nand U20125 (N_20125,N_19884,N_19900);
or U20126 (N_20126,N_19934,N_19933);
nor U20127 (N_20127,N_19928,N_19841);
or U20128 (N_20128,N_19916,N_19808);
nand U20129 (N_20129,N_19951,N_19926);
or U20130 (N_20130,N_19867,N_19903);
and U20131 (N_20131,N_19812,N_19911);
nor U20132 (N_20132,N_19899,N_19874);
nor U20133 (N_20133,N_19839,N_19899);
nand U20134 (N_20134,N_19986,N_19981);
nand U20135 (N_20135,N_19869,N_19918);
nand U20136 (N_20136,N_19934,N_19972);
and U20137 (N_20137,N_19821,N_19881);
nand U20138 (N_20138,N_19844,N_19897);
or U20139 (N_20139,N_19937,N_19902);
and U20140 (N_20140,N_19871,N_19986);
or U20141 (N_20141,N_19928,N_19945);
or U20142 (N_20142,N_19820,N_19862);
or U20143 (N_20143,N_19960,N_19813);
and U20144 (N_20144,N_19915,N_19842);
nor U20145 (N_20145,N_19945,N_19825);
nor U20146 (N_20146,N_19870,N_19928);
nor U20147 (N_20147,N_19936,N_19975);
or U20148 (N_20148,N_19902,N_19820);
nor U20149 (N_20149,N_19876,N_19869);
nand U20150 (N_20150,N_19874,N_19857);
nand U20151 (N_20151,N_19863,N_19926);
nor U20152 (N_20152,N_19901,N_19819);
nor U20153 (N_20153,N_19964,N_19847);
or U20154 (N_20154,N_19881,N_19981);
or U20155 (N_20155,N_19950,N_19998);
or U20156 (N_20156,N_19978,N_19999);
nor U20157 (N_20157,N_19817,N_19802);
nor U20158 (N_20158,N_19874,N_19839);
or U20159 (N_20159,N_19861,N_19824);
and U20160 (N_20160,N_19861,N_19943);
nand U20161 (N_20161,N_19816,N_19971);
or U20162 (N_20162,N_19934,N_19882);
xnor U20163 (N_20163,N_19927,N_19906);
nand U20164 (N_20164,N_19959,N_19910);
nand U20165 (N_20165,N_19965,N_19823);
or U20166 (N_20166,N_19940,N_19826);
and U20167 (N_20167,N_19843,N_19974);
nor U20168 (N_20168,N_19958,N_19830);
or U20169 (N_20169,N_19889,N_19954);
nand U20170 (N_20170,N_19880,N_19878);
or U20171 (N_20171,N_19966,N_19977);
or U20172 (N_20172,N_19947,N_19959);
nand U20173 (N_20173,N_19920,N_19853);
nand U20174 (N_20174,N_19869,N_19809);
or U20175 (N_20175,N_19998,N_19803);
and U20176 (N_20176,N_19848,N_19996);
and U20177 (N_20177,N_19819,N_19945);
nor U20178 (N_20178,N_19899,N_19824);
and U20179 (N_20179,N_19835,N_19809);
nand U20180 (N_20180,N_19874,N_19941);
nand U20181 (N_20181,N_19831,N_19915);
and U20182 (N_20182,N_19897,N_19972);
and U20183 (N_20183,N_19884,N_19964);
nand U20184 (N_20184,N_19896,N_19955);
nor U20185 (N_20185,N_19900,N_19874);
and U20186 (N_20186,N_19942,N_19917);
nand U20187 (N_20187,N_19933,N_19812);
and U20188 (N_20188,N_19806,N_19976);
nor U20189 (N_20189,N_19971,N_19890);
or U20190 (N_20190,N_19853,N_19913);
or U20191 (N_20191,N_19876,N_19858);
nor U20192 (N_20192,N_19808,N_19869);
or U20193 (N_20193,N_19847,N_19965);
nor U20194 (N_20194,N_19980,N_19918);
nor U20195 (N_20195,N_19822,N_19813);
nand U20196 (N_20196,N_19870,N_19822);
and U20197 (N_20197,N_19888,N_19895);
nand U20198 (N_20198,N_19991,N_19885);
and U20199 (N_20199,N_19806,N_19950);
and U20200 (N_20200,N_20174,N_20122);
nand U20201 (N_20201,N_20152,N_20193);
and U20202 (N_20202,N_20087,N_20145);
nand U20203 (N_20203,N_20118,N_20175);
or U20204 (N_20204,N_20127,N_20028);
and U20205 (N_20205,N_20165,N_20082);
nor U20206 (N_20206,N_20015,N_20000);
nand U20207 (N_20207,N_20185,N_20141);
xnor U20208 (N_20208,N_20159,N_20044);
nor U20209 (N_20209,N_20113,N_20137);
or U20210 (N_20210,N_20142,N_20121);
nor U20211 (N_20211,N_20149,N_20077);
or U20212 (N_20212,N_20022,N_20032);
nand U20213 (N_20213,N_20001,N_20154);
nand U20214 (N_20214,N_20008,N_20095);
nand U20215 (N_20215,N_20194,N_20055);
or U20216 (N_20216,N_20023,N_20172);
nor U20217 (N_20217,N_20140,N_20130);
xnor U20218 (N_20218,N_20078,N_20094);
and U20219 (N_20219,N_20106,N_20100);
nor U20220 (N_20220,N_20104,N_20050);
or U20221 (N_20221,N_20182,N_20116);
nor U20222 (N_20222,N_20092,N_20009);
nand U20223 (N_20223,N_20052,N_20156);
or U20224 (N_20224,N_20160,N_20021);
and U20225 (N_20225,N_20072,N_20187);
nor U20226 (N_20226,N_20128,N_20170);
nand U20227 (N_20227,N_20199,N_20099);
or U20228 (N_20228,N_20024,N_20198);
nand U20229 (N_20229,N_20006,N_20117);
nand U20230 (N_20230,N_20083,N_20071);
and U20231 (N_20231,N_20003,N_20062);
and U20232 (N_20232,N_20186,N_20042);
or U20233 (N_20233,N_20011,N_20060);
nor U20234 (N_20234,N_20169,N_20017);
and U20235 (N_20235,N_20153,N_20014);
nand U20236 (N_20236,N_20178,N_20059);
nor U20237 (N_20237,N_20041,N_20181);
nor U20238 (N_20238,N_20089,N_20047);
and U20239 (N_20239,N_20111,N_20012);
and U20240 (N_20240,N_20135,N_20007);
or U20241 (N_20241,N_20136,N_20162);
or U20242 (N_20242,N_20037,N_20048);
and U20243 (N_20243,N_20068,N_20123);
and U20244 (N_20244,N_20076,N_20105);
or U20245 (N_20245,N_20036,N_20080);
or U20246 (N_20246,N_20109,N_20053);
nor U20247 (N_20247,N_20013,N_20163);
and U20248 (N_20248,N_20084,N_20039);
nand U20249 (N_20249,N_20025,N_20016);
or U20250 (N_20250,N_20091,N_20073);
and U20251 (N_20251,N_20129,N_20144);
and U20252 (N_20252,N_20031,N_20030);
or U20253 (N_20253,N_20086,N_20067);
nor U20254 (N_20254,N_20146,N_20019);
nor U20255 (N_20255,N_20098,N_20102);
nand U20256 (N_20256,N_20132,N_20115);
nor U20257 (N_20257,N_20110,N_20108);
nand U20258 (N_20258,N_20191,N_20061);
nor U20259 (N_20259,N_20069,N_20033);
or U20260 (N_20260,N_20004,N_20190);
nor U20261 (N_20261,N_20029,N_20079);
nor U20262 (N_20262,N_20075,N_20049);
or U20263 (N_20263,N_20179,N_20088);
nand U20264 (N_20264,N_20035,N_20070);
nor U20265 (N_20265,N_20066,N_20161);
nor U20266 (N_20266,N_20064,N_20096);
and U20267 (N_20267,N_20051,N_20151);
or U20268 (N_20268,N_20119,N_20167);
nand U20269 (N_20269,N_20155,N_20056);
nand U20270 (N_20270,N_20057,N_20195);
nand U20271 (N_20271,N_20157,N_20101);
or U20272 (N_20272,N_20045,N_20107);
nor U20273 (N_20273,N_20114,N_20085);
and U20274 (N_20274,N_20046,N_20150);
nand U20275 (N_20275,N_20131,N_20093);
or U20276 (N_20276,N_20005,N_20112);
nand U20277 (N_20277,N_20143,N_20180);
nand U20278 (N_20278,N_20063,N_20177);
nand U20279 (N_20279,N_20124,N_20034);
or U20280 (N_20280,N_20147,N_20018);
nand U20281 (N_20281,N_20125,N_20065);
and U20282 (N_20282,N_20196,N_20126);
nand U20283 (N_20283,N_20134,N_20103);
and U20284 (N_20284,N_20090,N_20197);
or U20285 (N_20285,N_20002,N_20139);
nand U20286 (N_20286,N_20164,N_20040);
nand U20287 (N_20287,N_20168,N_20097);
and U20288 (N_20288,N_20043,N_20171);
nor U20289 (N_20289,N_20148,N_20133);
or U20290 (N_20290,N_20188,N_20038);
and U20291 (N_20291,N_20189,N_20166);
nand U20292 (N_20292,N_20183,N_20081);
and U20293 (N_20293,N_20184,N_20120);
or U20294 (N_20294,N_20026,N_20010);
xor U20295 (N_20295,N_20020,N_20074);
nand U20296 (N_20296,N_20176,N_20158);
nand U20297 (N_20297,N_20027,N_20058);
nand U20298 (N_20298,N_20054,N_20192);
nand U20299 (N_20299,N_20173,N_20138);
and U20300 (N_20300,N_20171,N_20068);
and U20301 (N_20301,N_20021,N_20062);
or U20302 (N_20302,N_20019,N_20059);
and U20303 (N_20303,N_20000,N_20174);
and U20304 (N_20304,N_20183,N_20083);
xnor U20305 (N_20305,N_20186,N_20076);
or U20306 (N_20306,N_20072,N_20032);
and U20307 (N_20307,N_20035,N_20160);
nor U20308 (N_20308,N_20096,N_20035);
and U20309 (N_20309,N_20028,N_20124);
nor U20310 (N_20310,N_20085,N_20058);
nor U20311 (N_20311,N_20062,N_20103);
and U20312 (N_20312,N_20119,N_20057);
nand U20313 (N_20313,N_20171,N_20163);
nand U20314 (N_20314,N_20092,N_20087);
nand U20315 (N_20315,N_20163,N_20107);
and U20316 (N_20316,N_20099,N_20151);
nor U20317 (N_20317,N_20157,N_20142);
and U20318 (N_20318,N_20008,N_20072);
and U20319 (N_20319,N_20123,N_20104);
and U20320 (N_20320,N_20116,N_20122);
or U20321 (N_20321,N_20099,N_20044);
nor U20322 (N_20322,N_20192,N_20161);
or U20323 (N_20323,N_20179,N_20147);
nand U20324 (N_20324,N_20152,N_20016);
nor U20325 (N_20325,N_20125,N_20075);
or U20326 (N_20326,N_20048,N_20019);
nor U20327 (N_20327,N_20169,N_20037);
and U20328 (N_20328,N_20128,N_20052);
nor U20329 (N_20329,N_20036,N_20018);
and U20330 (N_20330,N_20144,N_20058);
or U20331 (N_20331,N_20160,N_20079);
and U20332 (N_20332,N_20177,N_20011);
nand U20333 (N_20333,N_20066,N_20135);
or U20334 (N_20334,N_20031,N_20017);
and U20335 (N_20335,N_20187,N_20175);
nand U20336 (N_20336,N_20157,N_20016);
and U20337 (N_20337,N_20173,N_20103);
and U20338 (N_20338,N_20124,N_20011);
nand U20339 (N_20339,N_20130,N_20003);
or U20340 (N_20340,N_20075,N_20162);
or U20341 (N_20341,N_20133,N_20040);
nand U20342 (N_20342,N_20157,N_20172);
xor U20343 (N_20343,N_20119,N_20136);
nor U20344 (N_20344,N_20155,N_20196);
and U20345 (N_20345,N_20108,N_20021);
xor U20346 (N_20346,N_20030,N_20198);
or U20347 (N_20347,N_20154,N_20139);
or U20348 (N_20348,N_20159,N_20036);
nor U20349 (N_20349,N_20156,N_20124);
nand U20350 (N_20350,N_20068,N_20095);
nand U20351 (N_20351,N_20057,N_20060);
and U20352 (N_20352,N_20067,N_20127);
or U20353 (N_20353,N_20113,N_20132);
nand U20354 (N_20354,N_20088,N_20138);
nor U20355 (N_20355,N_20104,N_20040);
and U20356 (N_20356,N_20120,N_20021);
or U20357 (N_20357,N_20069,N_20013);
and U20358 (N_20358,N_20166,N_20097);
nor U20359 (N_20359,N_20058,N_20188);
nand U20360 (N_20360,N_20145,N_20090);
or U20361 (N_20361,N_20172,N_20169);
and U20362 (N_20362,N_20059,N_20030);
or U20363 (N_20363,N_20152,N_20138);
nor U20364 (N_20364,N_20026,N_20168);
nand U20365 (N_20365,N_20013,N_20047);
and U20366 (N_20366,N_20059,N_20120);
or U20367 (N_20367,N_20172,N_20158);
nor U20368 (N_20368,N_20078,N_20104);
or U20369 (N_20369,N_20000,N_20161);
nor U20370 (N_20370,N_20163,N_20111);
nor U20371 (N_20371,N_20102,N_20113);
nand U20372 (N_20372,N_20130,N_20105);
or U20373 (N_20373,N_20199,N_20092);
and U20374 (N_20374,N_20034,N_20199);
nand U20375 (N_20375,N_20187,N_20111);
xor U20376 (N_20376,N_20198,N_20167);
and U20377 (N_20377,N_20187,N_20058);
nor U20378 (N_20378,N_20099,N_20047);
nor U20379 (N_20379,N_20073,N_20113);
nor U20380 (N_20380,N_20111,N_20027);
nand U20381 (N_20381,N_20099,N_20131);
nand U20382 (N_20382,N_20012,N_20040);
and U20383 (N_20383,N_20073,N_20076);
nand U20384 (N_20384,N_20151,N_20140);
nor U20385 (N_20385,N_20137,N_20184);
or U20386 (N_20386,N_20084,N_20096);
nand U20387 (N_20387,N_20179,N_20124);
or U20388 (N_20388,N_20081,N_20001);
and U20389 (N_20389,N_20193,N_20010);
nand U20390 (N_20390,N_20078,N_20097);
nand U20391 (N_20391,N_20007,N_20021);
or U20392 (N_20392,N_20024,N_20151);
and U20393 (N_20393,N_20186,N_20070);
nand U20394 (N_20394,N_20107,N_20094);
nor U20395 (N_20395,N_20198,N_20095);
nor U20396 (N_20396,N_20014,N_20009);
xor U20397 (N_20397,N_20019,N_20155);
nand U20398 (N_20398,N_20132,N_20006);
nand U20399 (N_20399,N_20076,N_20106);
nor U20400 (N_20400,N_20373,N_20399);
or U20401 (N_20401,N_20244,N_20284);
or U20402 (N_20402,N_20338,N_20218);
nor U20403 (N_20403,N_20209,N_20362);
xnor U20404 (N_20404,N_20271,N_20272);
nand U20405 (N_20405,N_20319,N_20278);
or U20406 (N_20406,N_20255,N_20350);
or U20407 (N_20407,N_20379,N_20391);
nor U20408 (N_20408,N_20355,N_20242);
nor U20409 (N_20409,N_20266,N_20384);
or U20410 (N_20410,N_20365,N_20201);
or U20411 (N_20411,N_20285,N_20220);
xor U20412 (N_20412,N_20260,N_20394);
nor U20413 (N_20413,N_20308,N_20232);
nand U20414 (N_20414,N_20389,N_20213);
nand U20415 (N_20415,N_20323,N_20382);
or U20416 (N_20416,N_20225,N_20240);
nand U20417 (N_20417,N_20301,N_20320);
and U20418 (N_20418,N_20352,N_20318);
or U20419 (N_20419,N_20307,N_20316);
or U20420 (N_20420,N_20297,N_20235);
nor U20421 (N_20421,N_20296,N_20273);
and U20422 (N_20422,N_20359,N_20254);
or U20423 (N_20423,N_20287,N_20292);
and U20424 (N_20424,N_20356,N_20205);
nor U20425 (N_20425,N_20290,N_20357);
nand U20426 (N_20426,N_20239,N_20396);
or U20427 (N_20427,N_20336,N_20380);
nor U20428 (N_20428,N_20354,N_20325);
nor U20429 (N_20429,N_20317,N_20293);
nand U20430 (N_20430,N_20219,N_20358);
nand U20431 (N_20431,N_20253,N_20224);
nand U20432 (N_20432,N_20264,N_20376);
nand U20433 (N_20433,N_20223,N_20361);
or U20434 (N_20434,N_20314,N_20304);
nand U20435 (N_20435,N_20206,N_20249);
nand U20436 (N_20436,N_20247,N_20252);
or U20437 (N_20437,N_20360,N_20309);
or U20438 (N_20438,N_20286,N_20305);
and U20439 (N_20439,N_20246,N_20299);
or U20440 (N_20440,N_20234,N_20364);
nor U20441 (N_20441,N_20333,N_20230);
nor U20442 (N_20442,N_20215,N_20310);
or U20443 (N_20443,N_20383,N_20274);
and U20444 (N_20444,N_20270,N_20367);
and U20445 (N_20445,N_20261,N_20294);
or U20446 (N_20446,N_20257,N_20298);
nor U20447 (N_20447,N_20222,N_20275);
or U20448 (N_20448,N_20289,N_20236);
nor U20449 (N_20449,N_20324,N_20353);
or U20450 (N_20450,N_20334,N_20217);
or U20451 (N_20451,N_20214,N_20243);
nor U20452 (N_20452,N_20200,N_20245);
nand U20453 (N_20453,N_20368,N_20229);
or U20454 (N_20454,N_20340,N_20381);
or U20455 (N_20455,N_20395,N_20241);
or U20456 (N_20456,N_20306,N_20372);
or U20457 (N_20457,N_20371,N_20250);
xor U20458 (N_20458,N_20363,N_20313);
and U20459 (N_20459,N_20231,N_20335);
and U20460 (N_20460,N_20375,N_20328);
nor U20461 (N_20461,N_20393,N_20398);
nor U20462 (N_20462,N_20221,N_20349);
nor U20463 (N_20463,N_20295,N_20210);
and U20464 (N_20464,N_20212,N_20202);
nor U20465 (N_20465,N_20347,N_20263);
nor U20466 (N_20466,N_20262,N_20300);
and U20467 (N_20467,N_20326,N_20339);
nand U20468 (N_20468,N_20233,N_20311);
nand U20469 (N_20469,N_20321,N_20277);
nor U20470 (N_20470,N_20303,N_20228);
nand U20471 (N_20471,N_20211,N_20388);
and U20472 (N_20472,N_20283,N_20267);
nand U20473 (N_20473,N_20342,N_20280);
or U20474 (N_20474,N_20344,N_20227);
and U20475 (N_20475,N_20345,N_20248);
or U20476 (N_20476,N_20276,N_20377);
nor U20477 (N_20477,N_20302,N_20397);
or U20478 (N_20478,N_20332,N_20259);
or U20479 (N_20479,N_20386,N_20237);
and U20480 (N_20480,N_20258,N_20279);
nor U20481 (N_20481,N_20322,N_20251);
and U20482 (N_20482,N_20208,N_20369);
nand U20483 (N_20483,N_20256,N_20341);
nand U20484 (N_20484,N_20337,N_20351);
and U20485 (N_20485,N_20312,N_20374);
nor U20486 (N_20486,N_20387,N_20330);
nand U20487 (N_20487,N_20226,N_20385);
and U20488 (N_20488,N_20390,N_20378);
or U20489 (N_20489,N_20216,N_20238);
and U20490 (N_20490,N_20370,N_20203);
xor U20491 (N_20491,N_20315,N_20366);
nand U20492 (N_20492,N_20282,N_20291);
nand U20493 (N_20493,N_20268,N_20204);
and U20494 (N_20494,N_20207,N_20392);
nor U20495 (N_20495,N_20288,N_20269);
and U20496 (N_20496,N_20348,N_20281);
and U20497 (N_20497,N_20343,N_20329);
or U20498 (N_20498,N_20265,N_20331);
or U20499 (N_20499,N_20327,N_20346);
or U20500 (N_20500,N_20392,N_20224);
or U20501 (N_20501,N_20382,N_20256);
nand U20502 (N_20502,N_20333,N_20236);
and U20503 (N_20503,N_20396,N_20377);
nor U20504 (N_20504,N_20249,N_20235);
nand U20505 (N_20505,N_20279,N_20334);
nand U20506 (N_20506,N_20266,N_20395);
nand U20507 (N_20507,N_20298,N_20324);
or U20508 (N_20508,N_20360,N_20206);
or U20509 (N_20509,N_20294,N_20272);
and U20510 (N_20510,N_20257,N_20262);
nor U20511 (N_20511,N_20286,N_20395);
or U20512 (N_20512,N_20320,N_20246);
nor U20513 (N_20513,N_20263,N_20327);
nor U20514 (N_20514,N_20282,N_20218);
nor U20515 (N_20515,N_20271,N_20346);
or U20516 (N_20516,N_20381,N_20356);
nand U20517 (N_20517,N_20200,N_20272);
and U20518 (N_20518,N_20352,N_20399);
nor U20519 (N_20519,N_20370,N_20285);
nand U20520 (N_20520,N_20298,N_20348);
nand U20521 (N_20521,N_20262,N_20366);
or U20522 (N_20522,N_20303,N_20233);
or U20523 (N_20523,N_20277,N_20307);
nand U20524 (N_20524,N_20374,N_20244);
nor U20525 (N_20525,N_20307,N_20295);
nand U20526 (N_20526,N_20212,N_20372);
or U20527 (N_20527,N_20288,N_20266);
nand U20528 (N_20528,N_20206,N_20248);
nand U20529 (N_20529,N_20244,N_20220);
nand U20530 (N_20530,N_20243,N_20373);
nand U20531 (N_20531,N_20392,N_20214);
and U20532 (N_20532,N_20343,N_20259);
nor U20533 (N_20533,N_20308,N_20215);
or U20534 (N_20534,N_20367,N_20200);
nand U20535 (N_20535,N_20362,N_20320);
nor U20536 (N_20536,N_20363,N_20371);
or U20537 (N_20537,N_20326,N_20387);
or U20538 (N_20538,N_20267,N_20395);
or U20539 (N_20539,N_20331,N_20289);
nor U20540 (N_20540,N_20279,N_20283);
xnor U20541 (N_20541,N_20231,N_20259);
and U20542 (N_20542,N_20216,N_20210);
nor U20543 (N_20543,N_20306,N_20397);
nand U20544 (N_20544,N_20265,N_20276);
and U20545 (N_20545,N_20383,N_20253);
and U20546 (N_20546,N_20329,N_20256);
and U20547 (N_20547,N_20209,N_20373);
or U20548 (N_20548,N_20250,N_20290);
and U20549 (N_20549,N_20398,N_20330);
nor U20550 (N_20550,N_20260,N_20265);
or U20551 (N_20551,N_20221,N_20299);
or U20552 (N_20552,N_20220,N_20342);
nor U20553 (N_20553,N_20269,N_20358);
nand U20554 (N_20554,N_20397,N_20247);
or U20555 (N_20555,N_20205,N_20332);
or U20556 (N_20556,N_20345,N_20326);
nand U20557 (N_20557,N_20336,N_20343);
or U20558 (N_20558,N_20313,N_20371);
or U20559 (N_20559,N_20330,N_20272);
nand U20560 (N_20560,N_20233,N_20324);
nand U20561 (N_20561,N_20387,N_20323);
nor U20562 (N_20562,N_20389,N_20220);
and U20563 (N_20563,N_20201,N_20240);
or U20564 (N_20564,N_20279,N_20224);
nor U20565 (N_20565,N_20338,N_20272);
nor U20566 (N_20566,N_20337,N_20220);
nand U20567 (N_20567,N_20395,N_20301);
nand U20568 (N_20568,N_20364,N_20356);
nor U20569 (N_20569,N_20259,N_20357);
or U20570 (N_20570,N_20232,N_20277);
nor U20571 (N_20571,N_20357,N_20261);
and U20572 (N_20572,N_20234,N_20286);
or U20573 (N_20573,N_20347,N_20207);
or U20574 (N_20574,N_20389,N_20302);
nor U20575 (N_20575,N_20359,N_20378);
nand U20576 (N_20576,N_20280,N_20374);
nand U20577 (N_20577,N_20350,N_20262);
or U20578 (N_20578,N_20361,N_20333);
nor U20579 (N_20579,N_20225,N_20378);
nand U20580 (N_20580,N_20279,N_20259);
nand U20581 (N_20581,N_20294,N_20382);
nor U20582 (N_20582,N_20307,N_20368);
or U20583 (N_20583,N_20205,N_20301);
or U20584 (N_20584,N_20355,N_20253);
and U20585 (N_20585,N_20357,N_20214);
nand U20586 (N_20586,N_20344,N_20294);
or U20587 (N_20587,N_20217,N_20366);
xnor U20588 (N_20588,N_20372,N_20248);
nor U20589 (N_20589,N_20258,N_20275);
or U20590 (N_20590,N_20229,N_20219);
and U20591 (N_20591,N_20356,N_20383);
nand U20592 (N_20592,N_20296,N_20244);
and U20593 (N_20593,N_20310,N_20304);
nor U20594 (N_20594,N_20252,N_20283);
or U20595 (N_20595,N_20396,N_20322);
nor U20596 (N_20596,N_20328,N_20225);
and U20597 (N_20597,N_20218,N_20243);
nor U20598 (N_20598,N_20302,N_20399);
and U20599 (N_20599,N_20327,N_20294);
and U20600 (N_20600,N_20464,N_20477);
nand U20601 (N_20601,N_20554,N_20453);
or U20602 (N_20602,N_20434,N_20489);
nor U20603 (N_20603,N_20508,N_20580);
nand U20604 (N_20604,N_20476,N_20466);
and U20605 (N_20605,N_20407,N_20403);
and U20606 (N_20606,N_20447,N_20475);
and U20607 (N_20607,N_20412,N_20436);
nand U20608 (N_20608,N_20585,N_20571);
nor U20609 (N_20609,N_20472,N_20425);
nand U20610 (N_20610,N_20449,N_20423);
nor U20611 (N_20611,N_20536,N_20558);
nand U20612 (N_20612,N_20594,N_20576);
or U20613 (N_20613,N_20530,N_20456);
nand U20614 (N_20614,N_20599,N_20433);
nand U20615 (N_20615,N_20481,N_20550);
nand U20616 (N_20616,N_20442,N_20471);
and U20617 (N_20617,N_20406,N_20465);
nor U20618 (N_20618,N_20593,N_20428);
or U20619 (N_20619,N_20549,N_20467);
or U20620 (N_20620,N_20498,N_20409);
nor U20621 (N_20621,N_20596,N_20445);
nor U20622 (N_20622,N_20437,N_20517);
nor U20623 (N_20623,N_20555,N_20458);
nor U20624 (N_20624,N_20420,N_20452);
nand U20625 (N_20625,N_20521,N_20419);
or U20626 (N_20626,N_20418,N_20551);
or U20627 (N_20627,N_20504,N_20413);
and U20628 (N_20628,N_20483,N_20572);
nor U20629 (N_20629,N_20509,N_20541);
or U20630 (N_20630,N_20589,N_20562);
and U20631 (N_20631,N_20538,N_20523);
or U20632 (N_20632,N_20525,N_20546);
and U20633 (N_20633,N_20402,N_20564);
nand U20634 (N_20634,N_20410,N_20513);
or U20635 (N_20635,N_20516,N_20505);
nand U20636 (N_20636,N_20539,N_20527);
nor U20637 (N_20637,N_20454,N_20443);
nand U20638 (N_20638,N_20469,N_20426);
nand U20639 (N_20639,N_20537,N_20584);
or U20640 (N_20640,N_20520,N_20540);
nor U20641 (N_20641,N_20518,N_20470);
nand U20642 (N_20642,N_20491,N_20422);
or U20643 (N_20643,N_20569,N_20446);
nand U20644 (N_20644,N_20573,N_20457);
nor U20645 (N_20645,N_20512,N_20500);
nor U20646 (N_20646,N_20432,N_20482);
nor U20647 (N_20647,N_20577,N_20514);
nand U20648 (N_20648,N_20548,N_20408);
nor U20649 (N_20649,N_20460,N_20528);
or U20650 (N_20650,N_20496,N_20568);
and U20651 (N_20651,N_20424,N_20502);
and U20652 (N_20652,N_20455,N_20598);
and U20653 (N_20653,N_20444,N_20430);
or U20654 (N_20654,N_20533,N_20439);
or U20655 (N_20655,N_20590,N_20544);
and U20656 (N_20656,N_20438,N_20493);
nor U20657 (N_20657,N_20526,N_20582);
nor U20658 (N_20658,N_20566,N_20515);
nor U20659 (N_20659,N_20480,N_20435);
nor U20660 (N_20660,N_20559,N_20440);
or U20661 (N_20661,N_20567,N_20583);
nor U20662 (N_20662,N_20417,N_20415);
nor U20663 (N_20663,N_20400,N_20459);
and U20664 (N_20664,N_20542,N_20570);
nor U20665 (N_20665,N_20473,N_20556);
and U20666 (N_20666,N_20597,N_20522);
nand U20667 (N_20667,N_20488,N_20474);
or U20668 (N_20668,N_20545,N_20427);
and U20669 (N_20669,N_20578,N_20416);
nand U20670 (N_20670,N_20479,N_20451);
or U20671 (N_20671,N_20450,N_20462);
and U20672 (N_20672,N_20501,N_20586);
nand U20673 (N_20673,N_20507,N_20574);
or U20674 (N_20674,N_20486,N_20543);
xnor U20675 (N_20675,N_20441,N_20552);
nor U20676 (N_20676,N_20581,N_20511);
nor U20677 (N_20677,N_20563,N_20487);
nand U20678 (N_20678,N_20404,N_20519);
or U20679 (N_20679,N_20510,N_20414);
nor U20680 (N_20680,N_20506,N_20531);
or U20681 (N_20681,N_20495,N_20503);
or U20682 (N_20682,N_20592,N_20499);
or U20683 (N_20683,N_20494,N_20421);
nand U20684 (N_20684,N_20565,N_20497);
nand U20685 (N_20685,N_20448,N_20547);
and U20686 (N_20686,N_20561,N_20490);
or U20687 (N_20687,N_20591,N_20478);
nand U20688 (N_20688,N_20588,N_20405);
nand U20689 (N_20689,N_20587,N_20401);
nor U20690 (N_20690,N_20411,N_20535);
and U20691 (N_20691,N_20484,N_20534);
or U20692 (N_20692,N_20485,N_20468);
and U20693 (N_20693,N_20463,N_20492);
or U20694 (N_20694,N_20553,N_20429);
nand U20695 (N_20695,N_20431,N_20575);
and U20696 (N_20696,N_20529,N_20557);
nor U20697 (N_20697,N_20461,N_20595);
nand U20698 (N_20698,N_20532,N_20524);
nand U20699 (N_20699,N_20560,N_20579);
and U20700 (N_20700,N_20493,N_20435);
or U20701 (N_20701,N_20479,N_20573);
or U20702 (N_20702,N_20509,N_20415);
or U20703 (N_20703,N_20486,N_20525);
nor U20704 (N_20704,N_20590,N_20545);
or U20705 (N_20705,N_20493,N_20474);
nand U20706 (N_20706,N_20552,N_20488);
nor U20707 (N_20707,N_20426,N_20535);
or U20708 (N_20708,N_20590,N_20468);
nand U20709 (N_20709,N_20573,N_20452);
nor U20710 (N_20710,N_20567,N_20570);
xor U20711 (N_20711,N_20453,N_20463);
or U20712 (N_20712,N_20441,N_20483);
and U20713 (N_20713,N_20528,N_20459);
nand U20714 (N_20714,N_20595,N_20407);
nor U20715 (N_20715,N_20522,N_20458);
or U20716 (N_20716,N_20552,N_20578);
nand U20717 (N_20717,N_20567,N_20462);
nor U20718 (N_20718,N_20584,N_20581);
nand U20719 (N_20719,N_20460,N_20549);
and U20720 (N_20720,N_20540,N_20505);
and U20721 (N_20721,N_20414,N_20595);
nand U20722 (N_20722,N_20538,N_20504);
or U20723 (N_20723,N_20453,N_20502);
and U20724 (N_20724,N_20423,N_20461);
or U20725 (N_20725,N_20588,N_20510);
nand U20726 (N_20726,N_20579,N_20577);
or U20727 (N_20727,N_20424,N_20401);
nand U20728 (N_20728,N_20570,N_20496);
nand U20729 (N_20729,N_20587,N_20499);
nor U20730 (N_20730,N_20424,N_20556);
or U20731 (N_20731,N_20566,N_20593);
nor U20732 (N_20732,N_20547,N_20549);
nand U20733 (N_20733,N_20581,N_20407);
and U20734 (N_20734,N_20593,N_20451);
nor U20735 (N_20735,N_20401,N_20594);
and U20736 (N_20736,N_20563,N_20462);
xnor U20737 (N_20737,N_20539,N_20411);
and U20738 (N_20738,N_20596,N_20558);
and U20739 (N_20739,N_20560,N_20510);
nand U20740 (N_20740,N_20469,N_20443);
or U20741 (N_20741,N_20564,N_20554);
and U20742 (N_20742,N_20418,N_20548);
or U20743 (N_20743,N_20538,N_20426);
nor U20744 (N_20744,N_20547,N_20555);
nor U20745 (N_20745,N_20401,N_20407);
nor U20746 (N_20746,N_20459,N_20539);
and U20747 (N_20747,N_20507,N_20532);
or U20748 (N_20748,N_20469,N_20460);
and U20749 (N_20749,N_20558,N_20443);
or U20750 (N_20750,N_20462,N_20524);
or U20751 (N_20751,N_20561,N_20460);
or U20752 (N_20752,N_20404,N_20494);
nor U20753 (N_20753,N_20427,N_20567);
nand U20754 (N_20754,N_20577,N_20588);
or U20755 (N_20755,N_20454,N_20521);
or U20756 (N_20756,N_20405,N_20517);
and U20757 (N_20757,N_20535,N_20437);
nor U20758 (N_20758,N_20559,N_20421);
nand U20759 (N_20759,N_20466,N_20463);
nor U20760 (N_20760,N_20550,N_20591);
and U20761 (N_20761,N_20475,N_20571);
nor U20762 (N_20762,N_20478,N_20408);
or U20763 (N_20763,N_20561,N_20416);
nor U20764 (N_20764,N_20467,N_20526);
nand U20765 (N_20765,N_20450,N_20416);
nor U20766 (N_20766,N_20568,N_20444);
nor U20767 (N_20767,N_20533,N_20487);
nand U20768 (N_20768,N_20513,N_20415);
or U20769 (N_20769,N_20569,N_20405);
and U20770 (N_20770,N_20542,N_20423);
or U20771 (N_20771,N_20519,N_20557);
or U20772 (N_20772,N_20504,N_20491);
nand U20773 (N_20773,N_20515,N_20582);
or U20774 (N_20774,N_20557,N_20445);
nor U20775 (N_20775,N_20463,N_20550);
or U20776 (N_20776,N_20537,N_20499);
nand U20777 (N_20777,N_20479,N_20432);
or U20778 (N_20778,N_20567,N_20494);
or U20779 (N_20779,N_20574,N_20493);
or U20780 (N_20780,N_20414,N_20577);
nor U20781 (N_20781,N_20560,N_20415);
nand U20782 (N_20782,N_20474,N_20489);
nor U20783 (N_20783,N_20471,N_20548);
nor U20784 (N_20784,N_20505,N_20450);
nand U20785 (N_20785,N_20484,N_20585);
nor U20786 (N_20786,N_20542,N_20520);
nor U20787 (N_20787,N_20573,N_20423);
and U20788 (N_20788,N_20562,N_20437);
or U20789 (N_20789,N_20527,N_20422);
nand U20790 (N_20790,N_20491,N_20552);
nand U20791 (N_20791,N_20483,N_20490);
nand U20792 (N_20792,N_20535,N_20499);
nand U20793 (N_20793,N_20569,N_20532);
nor U20794 (N_20794,N_20420,N_20574);
nor U20795 (N_20795,N_20426,N_20400);
nor U20796 (N_20796,N_20530,N_20522);
nor U20797 (N_20797,N_20401,N_20586);
nand U20798 (N_20798,N_20439,N_20498);
and U20799 (N_20799,N_20402,N_20478);
or U20800 (N_20800,N_20657,N_20662);
nand U20801 (N_20801,N_20649,N_20761);
nor U20802 (N_20802,N_20631,N_20742);
nand U20803 (N_20803,N_20672,N_20633);
nand U20804 (N_20804,N_20629,N_20799);
or U20805 (N_20805,N_20783,N_20676);
or U20806 (N_20806,N_20729,N_20609);
nor U20807 (N_20807,N_20777,N_20767);
and U20808 (N_20808,N_20647,N_20764);
nand U20809 (N_20809,N_20719,N_20720);
nor U20810 (N_20810,N_20710,N_20787);
nor U20811 (N_20811,N_20715,N_20610);
or U20812 (N_20812,N_20660,N_20788);
and U20813 (N_20813,N_20686,N_20754);
nor U20814 (N_20814,N_20775,N_20648);
or U20815 (N_20815,N_20727,N_20785);
or U20816 (N_20816,N_20658,N_20630);
or U20817 (N_20817,N_20701,N_20721);
and U20818 (N_20818,N_20759,N_20704);
nor U20819 (N_20819,N_20697,N_20691);
nor U20820 (N_20820,N_20753,N_20746);
nand U20821 (N_20821,N_20650,N_20778);
and U20822 (N_20822,N_20750,N_20693);
nor U20823 (N_20823,N_20705,N_20646);
nor U20824 (N_20824,N_20690,N_20780);
nand U20825 (N_20825,N_20644,N_20632);
nand U20826 (N_20826,N_20794,N_20659);
nor U20827 (N_20827,N_20613,N_20669);
and U20828 (N_20828,N_20699,N_20665);
or U20829 (N_20829,N_20616,N_20674);
nand U20830 (N_20830,N_20656,N_20752);
or U20831 (N_20831,N_20714,N_20680);
nor U20832 (N_20832,N_20703,N_20792);
nand U20833 (N_20833,N_20735,N_20702);
nand U20834 (N_20834,N_20639,N_20700);
nor U20835 (N_20835,N_20677,N_20653);
nand U20836 (N_20836,N_20620,N_20698);
or U20837 (N_20837,N_20755,N_20689);
and U20838 (N_20838,N_20741,N_20793);
and U20839 (N_20839,N_20790,N_20762);
nor U20840 (N_20840,N_20604,N_20760);
nor U20841 (N_20841,N_20751,N_20772);
nand U20842 (N_20842,N_20743,N_20723);
nor U20843 (N_20843,N_20694,N_20687);
and U20844 (N_20844,N_20776,N_20756);
or U20845 (N_20845,N_20725,N_20744);
nor U20846 (N_20846,N_20685,N_20605);
nor U20847 (N_20847,N_20706,N_20625);
and U20848 (N_20848,N_20724,N_20722);
nor U20849 (N_20849,N_20765,N_20600);
nand U20850 (N_20850,N_20758,N_20675);
nand U20851 (N_20851,N_20607,N_20798);
nand U20852 (N_20852,N_20717,N_20654);
nor U20853 (N_20853,N_20622,N_20748);
and U20854 (N_20854,N_20627,N_20683);
and U20855 (N_20855,N_20711,N_20664);
or U20856 (N_20856,N_20695,N_20641);
nand U20857 (N_20857,N_20626,N_20713);
nand U20858 (N_20858,N_20636,N_20730);
or U20859 (N_20859,N_20796,N_20770);
and U20860 (N_20860,N_20668,N_20749);
nor U20861 (N_20861,N_20786,N_20635);
nor U20862 (N_20862,N_20673,N_20769);
nand U20863 (N_20863,N_20709,N_20617);
and U20864 (N_20864,N_20745,N_20682);
nor U20865 (N_20865,N_20681,N_20651);
or U20866 (N_20866,N_20679,N_20784);
nor U20867 (N_20867,N_20612,N_20789);
and U20868 (N_20868,N_20779,N_20726);
and U20869 (N_20869,N_20708,N_20640);
or U20870 (N_20870,N_20712,N_20740);
or U20871 (N_20871,N_20628,N_20603);
or U20872 (N_20872,N_20738,N_20663);
and U20873 (N_20873,N_20614,N_20757);
or U20874 (N_20874,N_20606,N_20688);
nor U20875 (N_20875,N_20716,N_20623);
and U20876 (N_20876,N_20739,N_20791);
or U20877 (N_20877,N_20692,N_20661);
nor U20878 (N_20878,N_20782,N_20747);
and U20879 (N_20879,N_20670,N_20642);
nor U20880 (N_20880,N_20718,N_20601);
nand U20881 (N_20881,N_20734,N_20652);
and U20882 (N_20882,N_20763,N_20781);
nor U20883 (N_20883,N_20643,N_20696);
and U20884 (N_20884,N_20773,N_20634);
or U20885 (N_20885,N_20637,N_20602);
nand U20886 (N_20886,N_20678,N_20671);
or U20887 (N_20887,N_20608,N_20731);
or U20888 (N_20888,N_20707,N_20766);
nor U20889 (N_20889,N_20666,N_20733);
and U20890 (N_20890,N_20618,N_20736);
and U20891 (N_20891,N_20615,N_20684);
and U20892 (N_20892,N_20611,N_20797);
xor U20893 (N_20893,N_20737,N_20768);
nand U20894 (N_20894,N_20655,N_20667);
nor U20895 (N_20895,N_20621,N_20645);
and U20896 (N_20896,N_20728,N_20732);
and U20897 (N_20897,N_20771,N_20624);
nand U20898 (N_20898,N_20774,N_20795);
and U20899 (N_20899,N_20619,N_20638);
nor U20900 (N_20900,N_20638,N_20714);
nand U20901 (N_20901,N_20766,N_20747);
and U20902 (N_20902,N_20734,N_20763);
nand U20903 (N_20903,N_20660,N_20727);
or U20904 (N_20904,N_20687,N_20793);
nor U20905 (N_20905,N_20755,N_20617);
and U20906 (N_20906,N_20610,N_20708);
and U20907 (N_20907,N_20636,N_20669);
or U20908 (N_20908,N_20728,N_20629);
or U20909 (N_20909,N_20734,N_20783);
or U20910 (N_20910,N_20732,N_20651);
nand U20911 (N_20911,N_20702,N_20700);
and U20912 (N_20912,N_20623,N_20634);
nor U20913 (N_20913,N_20668,N_20612);
nand U20914 (N_20914,N_20759,N_20709);
or U20915 (N_20915,N_20634,N_20611);
and U20916 (N_20916,N_20680,N_20612);
or U20917 (N_20917,N_20686,N_20622);
and U20918 (N_20918,N_20733,N_20792);
or U20919 (N_20919,N_20770,N_20627);
and U20920 (N_20920,N_20690,N_20605);
or U20921 (N_20921,N_20625,N_20651);
or U20922 (N_20922,N_20627,N_20624);
nor U20923 (N_20923,N_20604,N_20795);
nand U20924 (N_20924,N_20657,N_20665);
nand U20925 (N_20925,N_20783,N_20669);
and U20926 (N_20926,N_20729,N_20624);
or U20927 (N_20927,N_20791,N_20748);
nand U20928 (N_20928,N_20709,N_20623);
nor U20929 (N_20929,N_20703,N_20724);
or U20930 (N_20930,N_20763,N_20736);
nor U20931 (N_20931,N_20776,N_20657);
nand U20932 (N_20932,N_20785,N_20620);
or U20933 (N_20933,N_20654,N_20734);
nor U20934 (N_20934,N_20785,N_20792);
nor U20935 (N_20935,N_20798,N_20784);
nor U20936 (N_20936,N_20739,N_20606);
and U20937 (N_20937,N_20645,N_20727);
or U20938 (N_20938,N_20623,N_20790);
and U20939 (N_20939,N_20777,N_20610);
nor U20940 (N_20940,N_20679,N_20642);
nor U20941 (N_20941,N_20677,N_20645);
and U20942 (N_20942,N_20719,N_20744);
or U20943 (N_20943,N_20710,N_20672);
and U20944 (N_20944,N_20677,N_20721);
nand U20945 (N_20945,N_20721,N_20766);
nand U20946 (N_20946,N_20605,N_20781);
nand U20947 (N_20947,N_20680,N_20791);
or U20948 (N_20948,N_20765,N_20678);
nand U20949 (N_20949,N_20633,N_20735);
nand U20950 (N_20950,N_20749,N_20602);
nor U20951 (N_20951,N_20688,N_20600);
nor U20952 (N_20952,N_20781,N_20734);
nor U20953 (N_20953,N_20774,N_20711);
nor U20954 (N_20954,N_20652,N_20787);
or U20955 (N_20955,N_20696,N_20745);
and U20956 (N_20956,N_20704,N_20676);
or U20957 (N_20957,N_20706,N_20724);
and U20958 (N_20958,N_20699,N_20740);
nor U20959 (N_20959,N_20728,N_20673);
nand U20960 (N_20960,N_20659,N_20684);
and U20961 (N_20961,N_20724,N_20622);
nand U20962 (N_20962,N_20710,N_20629);
or U20963 (N_20963,N_20680,N_20780);
or U20964 (N_20964,N_20712,N_20631);
nor U20965 (N_20965,N_20795,N_20712);
nand U20966 (N_20966,N_20798,N_20641);
nand U20967 (N_20967,N_20639,N_20785);
and U20968 (N_20968,N_20741,N_20671);
and U20969 (N_20969,N_20685,N_20760);
or U20970 (N_20970,N_20731,N_20663);
nor U20971 (N_20971,N_20715,N_20709);
nand U20972 (N_20972,N_20724,N_20749);
and U20973 (N_20973,N_20690,N_20698);
or U20974 (N_20974,N_20795,N_20689);
nor U20975 (N_20975,N_20771,N_20690);
nand U20976 (N_20976,N_20795,N_20624);
xor U20977 (N_20977,N_20602,N_20748);
nand U20978 (N_20978,N_20766,N_20622);
nor U20979 (N_20979,N_20688,N_20658);
nor U20980 (N_20980,N_20701,N_20730);
nor U20981 (N_20981,N_20778,N_20677);
or U20982 (N_20982,N_20729,N_20728);
nand U20983 (N_20983,N_20660,N_20624);
or U20984 (N_20984,N_20796,N_20756);
nor U20985 (N_20985,N_20736,N_20718);
and U20986 (N_20986,N_20767,N_20704);
and U20987 (N_20987,N_20669,N_20750);
and U20988 (N_20988,N_20709,N_20691);
nor U20989 (N_20989,N_20690,N_20715);
or U20990 (N_20990,N_20656,N_20684);
or U20991 (N_20991,N_20741,N_20768);
nand U20992 (N_20992,N_20607,N_20736);
and U20993 (N_20993,N_20630,N_20710);
nand U20994 (N_20994,N_20783,N_20612);
or U20995 (N_20995,N_20768,N_20615);
and U20996 (N_20996,N_20751,N_20728);
or U20997 (N_20997,N_20658,N_20757);
and U20998 (N_20998,N_20640,N_20634);
nand U20999 (N_20999,N_20658,N_20676);
and U21000 (N_21000,N_20930,N_20871);
or U21001 (N_21001,N_20963,N_20847);
and U21002 (N_21002,N_20857,N_20834);
nor U21003 (N_21003,N_20993,N_20926);
nor U21004 (N_21004,N_20814,N_20985);
nand U21005 (N_21005,N_20815,N_20896);
nand U21006 (N_21006,N_20906,N_20932);
and U21007 (N_21007,N_20875,N_20910);
nand U21008 (N_21008,N_20803,N_20839);
or U21009 (N_21009,N_20971,N_20947);
or U21010 (N_21010,N_20841,N_20830);
or U21011 (N_21011,N_20995,N_20821);
nor U21012 (N_21012,N_20991,N_20935);
nor U21013 (N_21013,N_20914,N_20923);
or U21014 (N_21014,N_20917,N_20825);
or U21015 (N_21015,N_20913,N_20800);
or U21016 (N_21016,N_20946,N_20883);
nor U21017 (N_21017,N_20809,N_20873);
or U21018 (N_21018,N_20812,N_20874);
and U21019 (N_21019,N_20826,N_20822);
nor U21020 (N_21020,N_20843,N_20885);
and U21021 (N_21021,N_20832,N_20924);
and U21022 (N_21022,N_20992,N_20855);
or U21023 (N_21023,N_20864,N_20999);
nor U21024 (N_21024,N_20901,N_20900);
and U21025 (N_21025,N_20919,N_20860);
nor U21026 (N_21026,N_20844,N_20911);
or U21027 (N_21027,N_20816,N_20967);
nand U21028 (N_21028,N_20813,N_20863);
nor U21029 (N_21029,N_20819,N_20884);
or U21030 (N_21030,N_20944,N_20850);
nand U21031 (N_21031,N_20876,N_20804);
and U21032 (N_21032,N_20977,N_20962);
nand U21033 (N_21033,N_20805,N_20820);
and U21034 (N_21034,N_20909,N_20888);
and U21035 (N_21035,N_20808,N_20966);
and U21036 (N_21036,N_20867,N_20802);
or U21037 (N_21037,N_20929,N_20972);
or U21038 (N_21038,N_20856,N_20903);
nor U21039 (N_21039,N_20976,N_20892);
xnor U21040 (N_21040,N_20954,N_20978);
and U21041 (N_21041,N_20949,N_20945);
and U21042 (N_21042,N_20958,N_20968);
nor U21043 (N_21043,N_20965,N_20810);
or U21044 (N_21044,N_20907,N_20891);
nand U21045 (N_21045,N_20941,N_20899);
or U21046 (N_21046,N_20940,N_20865);
nand U21047 (N_21047,N_20838,N_20937);
nand U21048 (N_21048,N_20886,N_20955);
nand U21049 (N_21049,N_20952,N_20854);
nand U21050 (N_21050,N_20837,N_20928);
nor U21051 (N_21051,N_20973,N_20893);
and U21052 (N_21052,N_20931,N_20922);
nand U21053 (N_21053,N_20898,N_20806);
nor U21054 (N_21054,N_20936,N_20984);
nand U21055 (N_21055,N_20964,N_20957);
nand U21056 (N_21056,N_20878,N_20969);
nor U21057 (N_21057,N_20953,N_20934);
or U21058 (N_21058,N_20861,N_20938);
nand U21059 (N_21059,N_20882,N_20987);
nor U21060 (N_21060,N_20840,N_20996);
nor U21061 (N_21061,N_20948,N_20982);
nand U21062 (N_21062,N_20890,N_20927);
nor U21063 (N_21063,N_20869,N_20879);
or U21064 (N_21064,N_20974,N_20951);
nand U21065 (N_21065,N_20902,N_20859);
nor U21066 (N_21066,N_20872,N_20866);
nand U21067 (N_21067,N_20918,N_20994);
nand U21068 (N_21068,N_20894,N_20858);
and U21069 (N_21069,N_20933,N_20998);
nor U21070 (N_21070,N_20912,N_20960);
or U21071 (N_21071,N_20836,N_20811);
nor U21072 (N_21072,N_20942,N_20823);
or U21073 (N_21073,N_20904,N_20915);
and U21074 (N_21074,N_20835,N_20950);
and U21075 (N_21075,N_20921,N_20897);
nand U21076 (N_21076,N_20925,N_20989);
nor U21077 (N_21077,N_20920,N_20997);
and U21078 (N_21078,N_20979,N_20905);
nand U21079 (N_21079,N_20981,N_20970);
or U21080 (N_21080,N_20990,N_20956);
nand U21081 (N_21081,N_20846,N_20880);
xnor U21082 (N_21082,N_20862,N_20939);
nor U21083 (N_21083,N_20853,N_20961);
and U21084 (N_21084,N_20983,N_20988);
nor U21085 (N_21085,N_20959,N_20852);
nor U21086 (N_21086,N_20975,N_20881);
nand U21087 (N_21087,N_20980,N_20848);
nand U21088 (N_21088,N_20807,N_20943);
nor U21089 (N_21089,N_20851,N_20845);
nor U21090 (N_21090,N_20824,N_20817);
nand U21091 (N_21091,N_20833,N_20829);
nand U21092 (N_21092,N_20842,N_20916);
nand U21093 (N_21093,N_20908,N_20889);
and U21094 (N_21094,N_20868,N_20801);
and U21095 (N_21095,N_20827,N_20986);
or U21096 (N_21096,N_20895,N_20828);
and U21097 (N_21097,N_20831,N_20887);
or U21098 (N_21098,N_20849,N_20877);
nor U21099 (N_21099,N_20870,N_20818);
or U21100 (N_21100,N_20862,N_20899);
or U21101 (N_21101,N_20946,N_20954);
nor U21102 (N_21102,N_20816,N_20930);
and U21103 (N_21103,N_20932,N_20886);
and U21104 (N_21104,N_20944,N_20805);
nor U21105 (N_21105,N_20898,N_20868);
nand U21106 (N_21106,N_20861,N_20918);
nand U21107 (N_21107,N_20816,N_20865);
or U21108 (N_21108,N_20857,N_20946);
or U21109 (N_21109,N_20870,N_20859);
nor U21110 (N_21110,N_20873,N_20981);
nand U21111 (N_21111,N_20937,N_20853);
and U21112 (N_21112,N_20925,N_20914);
nand U21113 (N_21113,N_20822,N_20879);
nand U21114 (N_21114,N_20912,N_20888);
nor U21115 (N_21115,N_20915,N_20945);
or U21116 (N_21116,N_20869,N_20898);
or U21117 (N_21117,N_20875,N_20924);
or U21118 (N_21118,N_20921,N_20974);
and U21119 (N_21119,N_20899,N_20840);
nand U21120 (N_21120,N_20892,N_20939);
nor U21121 (N_21121,N_20825,N_20854);
nand U21122 (N_21122,N_20975,N_20827);
or U21123 (N_21123,N_20886,N_20937);
nor U21124 (N_21124,N_20980,N_20956);
and U21125 (N_21125,N_20806,N_20860);
nand U21126 (N_21126,N_20961,N_20861);
nor U21127 (N_21127,N_20973,N_20803);
nor U21128 (N_21128,N_20808,N_20999);
or U21129 (N_21129,N_20924,N_20939);
nor U21130 (N_21130,N_20999,N_20945);
nor U21131 (N_21131,N_20985,N_20837);
nor U21132 (N_21132,N_20984,N_20990);
and U21133 (N_21133,N_20970,N_20869);
and U21134 (N_21134,N_20921,N_20935);
or U21135 (N_21135,N_20908,N_20971);
nor U21136 (N_21136,N_20976,N_20935);
and U21137 (N_21137,N_20923,N_20824);
or U21138 (N_21138,N_20946,N_20992);
and U21139 (N_21139,N_20943,N_20887);
nor U21140 (N_21140,N_20846,N_20885);
nand U21141 (N_21141,N_20814,N_20857);
or U21142 (N_21142,N_20954,N_20867);
nand U21143 (N_21143,N_20920,N_20951);
nor U21144 (N_21144,N_20939,N_20852);
nand U21145 (N_21145,N_20887,N_20928);
nor U21146 (N_21146,N_20997,N_20991);
or U21147 (N_21147,N_20898,N_20852);
nand U21148 (N_21148,N_20805,N_20824);
nor U21149 (N_21149,N_20842,N_20829);
or U21150 (N_21150,N_20833,N_20822);
nand U21151 (N_21151,N_20818,N_20869);
nor U21152 (N_21152,N_20823,N_20957);
nand U21153 (N_21153,N_20903,N_20981);
or U21154 (N_21154,N_20898,N_20835);
nor U21155 (N_21155,N_20855,N_20967);
nor U21156 (N_21156,N_20866,N_20827);
and U21157 (N_21157,N_20831,N_20812);
nor U21158 (N_21158,N_20887,N_20839);
or U21159 (N_21159,N_20853,N_20908);
nor U21160 (N_21160,N_20957,N_20837);
nor U21161 (N_21161,N_20868,N_20864);
or U21162 (N_21162,N_20979,N_20973);
and U21163 (N_21163,N_20814,N_20809);
or U21164 (N_21164,N_20926,N_20818);
and U21165 (N_21165,N_20900,N_20903);
nor U21166 (N_21166,N_20912,N_20878);
nor U21167 (N_21167,N_20903,N_20972);
nor U21168 (N_21168,N_20847,N_20939);
and U21169 (N_21169,N_20902,N_20858);
and U21170 (N_21170,N_20963,N_20916);
nand U21171 (N_21171,N_20948,N_20845);
and U21172 (N_21172,N_20849,N_20901);
and U21173 (N_21173,N_20934,N_20930);
or U21174 (N_21174,N_20822,N_20915);
and U21175 (N_21175,N_20867,N_20890);
xnor U21176 (N_21176,N_20909,N_20887);
and U21177 (N_21177,N_20999,N_20876);
or U21178 (N_21178,N_20913,N_20810);
nor U21179 (N_21179,N_20808,N_20924);
or U21180 (N_21180,N_20831,N_20924);
or U21181 (N_21181,N_20855,N_20851);
or U21182 (N_21182,N_20809,N_20824);
or U21183 (N_21183,N_20976,N_20884);
nand U21184 (N_21184,N_20880,N_20831);
or U21185 (N_21185,N_20817,N_20950);
nor U21186 (N_21186,N_20886,N_20849);
nor U21187 (N_21187,N_20919,N_20909);
or U21188 (N_21188,N_20916,N_20892);
and U21189 (N_21189,N_20924,N_20805);
nor U21190 (N_21190,N_20964,N_20927);
or U21191 (N_21191,N_20987,N_20909);
nand U21192 (N_21192,N_20869,N_20800);
and U21193 (N_21193,N_20956,N_20925);
and U21194 (N_21194,N_20806,N_20810);
nor U21195 (N_21195,N_20909,N_20975);
and U21196 (N_21196,N_20879,N_20996);
or U21197 (N_21197,N_20960,N_20972);
and U21198 (N_21198,N_20802,N_20977);
or U21199 (N_21199,N_20881,N_20837);
and U21200 (N_21200,N_21112,N_21041);
nand U21201 (N_21201,N_21035,N_21192);
nand U21202 (N_21202,N_21072,N_21169);
and U21203 (N_21203,N_21151,N_21125);
and U21204 (N_21204,N_21045,N_21084);
or U21205 (N_21205,N_21066,N_21160);
nand U21206 (N_21206,N_21166,N_21038);
and U21207 (N_21207,N_21080,N_21088);
or U21208 (N_21208,N_21176,N_21056);
and U21209 (N_21209,N_21193,N_21065);
nand U21210 (N_21210,N_21092,N_21191);
or U21211 (N_21211,N_21006,N_21033);
nor U21212 (N_21212,N_21113,N_21040);
nor U21213 (N_21213,N_21198,N_21139);
and U21214 (N_21214,N_21094,N_21182);
nor U21215 (N_21215,N_21147,N_21070);
nor U21216 (N_21216,N_21052,N_21172);
nand U21217 (N_21217,N_21102,N_21087);
nand U21218 (N_21218,N_21150,N_21091);
and U21219 (N_21219,N_21077,N_21188);
and U21220 (N_21220,N_21116,N_21068);
or U21221 (N_21221,N_21111,N_21099);
and U21222 (N_21222,N_21141,N_21007);
or U21223 (N_21223,N_21046,N_21109);
nand U21224 (N_21224,N_21011,N_21089);
or U21225 (N_21225,N_21181,N_21009);
or U21226 (N_21226,N_21135,N_21002);
nor U21227 (N_21227,N_21034,N_21130);
nand U21228 (N_21228,N_21042,N_21095);
and U21229 (N_21229,N_21026,N_21104);
nor U21230 (N_21230,N_21067,N_21164);
or U21231 (N_21231,N_21143,N_21144);
nand U21232 (N_21232,N_21179,N_21013);
nor U21233 (N_21233,N_21133,N_21050);
nand U21234 (N_21234,N_21024,N_21060);
and U21235 (N_21235,N_21146,N_21027);
nor U21236 (N_21236,N_21163,N_21054);
nand U21237 (N_21237,N_21051,N_21162);
nor U21238 (N_21238,N_21184,N_21189);
nand U21239 (N_21239,N_21173,N_21145);
nand U21240 (N_21240,N_21103,N_21069);
nor U21241 (N_21241,N_21093,N_21016);
or U21242 (N_21242,N_21017,N_21129);
nor U21243 (N_21243,N_21121,N_21155);
nor U21244 (N_21244,N_21124,N_21115);
nor U21245 (N_21245,N_21174,N_21106);
and U21246 (N_21246,N_21048,N_21148);
nor U21247 (N_21247,N_21128,N_21197);
or U21248 (N_21248,N_21071,N_21161);
or U21249 (N_21249,N_21190,N_21074);
or U21250 (N_21250,N_21186,N_21175);
nor U21251 (N_21251,N_21196,N_21015);
and U21252 (N_21252,N_21098,N_21142);
or U21253 (N_21253,N_21108,N_21123);
and U21254 (N_21254,N_21136,N_21047);
nand U21255 (N_21255,N_21180,N_21185);
nand U21256 (N_21256,N_21014,N_21000);
or U21257 (N_21257,N_21018,N_21120);
and U21258 (N_21258,N_21167,N_21001);
or U21259 (N_21259,N_21158,N_21075);
nand U21260 (N_21260,N_21153,N_21171);
or U21261 (N_21261,N_21012,N_21025);
nor U21262 (N_21262,N_21183,N_21081);
and U21263 (N_21263,N_21083,N_21096);
or U21264 (N_21264,N_21101,N_21177);
or U21265 (N_21265,N_21061,N_21079);
nand U21266 (N_21266,N_21010,N_21097);
and U21267 (N_21267,N_21063,N_21059);
or U21268 (N_21268,N_21031,N_21187);
nand U21269 (N_21269,N_21126,N_21049);
and U21270 (N_21270,N_21064,N_21029);
nand U21271 (N_21271,N_21127,N_21023);
or U21272 (N_21272,N_21076,N_21152);
nand U21273 (N_21273,N_21085,N_21131);
nor U21274 (N_21274,N_21039,N_21119);
or U21275 (N_21275,N_21058,N_21003);
nor U21276 (N_21276,N_21043,N_21082);
or U21277 (N_21277,N_21055,N_21030);
nor U21278 (N_21278,N_21086,N_21100);
nand U21279 (N_21279,N_21020,N_21154);
or U21280 (N_21280,N_21149,N_21078);
nor U21281 (N_21281,N_21019,N_21137);
nor U21282 (N_21282,N_21105,N_21165);
nor U21283 (N_21283,N_21110,N_21022);
or U21284 (N_21284,N_21118,N_21156);
or U21285 (N_21285,N_21159,N_21008);
and U21286 (N_21286,N_21157,N_21028);
or U21287 (N_21287,N_21138,N_21021);
or U21288 (N_21288,N_21036,N_21132);
nand U21289 (N_21289,N_21004,N_21195);
and U21290 (N_21290,N_21199,N_21037);
and U21291 (N_21291,N_21073,N_21005);
nor U21292 (N_21292,N_21032,N_21053);
and U21293 (N_21293,N_21117,N_21194);
and U21294 (N_21294,N_21057,N_21062);
or U21295 (N_21295,N_21170,N_21044);
nor U21296 (N_21296,N_21178,N_21122);
nor U21297 (N_21297,N_21107,N_21140);
or U21298 (N_21298,N_21114,N_21134);
or U21299 (N_21299,N_21090,N_21168);
and U21300 (N_21300,N_21011,N_21051);
and U21301 (N_21301,N_21164,N_21172);
nor U21302 (N_21302,N_21066,N_21140);
or U21303 (N_21303,N_21101,N_21180);
and U21304 (N_21304,N_21142,N_21198);
or U21305 (N_21305,N_21138,N_21183);
nand U21306 (N_21306,N_21171,N_21088);
nand U21307 (N_21307,N_21102,N_21092);
and U21308 (N_21308,N_21129,N_21174);
nand U21309 (N_21309,N_21136,N_21143);
nor U21310 (N_21310,N_21009,N_21187);
nand U21311 (N_21311,N_21135,N_21100);
nand U21312 (N_21312,N_21190,N_21118);
xnor U21313 (N_21313,N_21046,N_21113);
nand U21314 (N_21314,N_21128,N_21071);
or U21315 (N_21315,N_21118,N_21079);
or U21316 (N_21316,N_21005,N_21168);
nor U21317 (N_21317,N_21056,N_21195);
or U21318 (N_21318,N_21183,N_21048);
and U21319 (N_21319,N_21102,N_21081);
nor U21320 (N_21320,N_21085,N_21056);
and U21321 (N_21321,N_21132,N_21055);
nand U21322 (N_21322,N_21170,N_21050);
or U21323 (N_21323,N_21007,N_21154);
and U21324 (N_21324,N_21050,N_21185);
and U21325 (N_21325,N_21068,N_21198);
or U21326 (N_21326,N_21073,N_21061);
nand U21327 (N_21327,N_21112,N_21048);
nand U21328 (N_21328,N_21179,N_21046);
xnor U21329 (N_21329,N_21129,N_21044);
nor U21330 (N_21330,N_21028,N_21009);
nor U21331 (N_21331,N_21005,N_21152);
nor U21332 (N_21332,N_21095,N_21011);
or U21333 (N_21333,N_21178,N_21104);
nand U21334 (N_21334,N_21016,N_21153);
nor U21335 (N_21335,N_21196,N_21060);
nor U21336 (N_21336,N_21165,N_21004);
nand U21337 (N_21337,N_21058,N_21067);
or U21338 (N_21338,N_21171,N_21137);
nand U21339 (N_21339,N_21186,N_21139);
and U21340 (N_21340,N_21078,N_21162);
or U21341 (N_21341,N_21038,N_21169);
nand U21342 (N_21342,N_21060,N_21031);
and U21343 (N_21343,N_21083,N_21023);
nand U21344 (N_21344,N_21109,N_21156);
and U21345 (N_21345,N_21119,N_21095);
or U21346 (N_21346,N_21118,N_21068);
nand U21347 (N_21347,N_21190,N_21177);
and U21348 (N_21348,N_21099,N_21053);
or U21349 (N_21349,N_21139,N_21074);
and U21350 (N_21350,N_21114,N_21012);
and U21351 (N_21351,N_21121,N_21199);
nor U21352 (N_21352,N_21080,N_21115);
or U21353 (N_21353,N_21163,N_21111);
nand U21354 (N_21354,N_21144,N_21020);
nor U21355 (N_21355,N_21039,N_21058);
nand U21356 (N_21356,N_21084,N_21005);
or U21357 (N_21357,N_21101,N_21164);
or U21358 (N_21358,N_21112,N_21089);
nor U21359 (N_21359,N_21145,N_21098);
nor U21360 (N_21360,N_21109,N_21139);
and U21361 (N_21361,N_21102,N_21026);
or U21362 (N_21362,N_21180,N_21154);
nor U21363 (N_21363,N_21054,N_21100);
nand U21364 (N_21364,N_21180,N_21059);
or U21365 (N_21365,N_21018,N_21189);
and U21366 (N_21366,N_21089,N_21123);
nand U21367 (N_21367,N_21131,N_21048);
xor U21368 (N_21368,N_21067,N_21138);
nor U21369 (N_21369,N_21190,N_21003);
nand U21370 (N_21370,N_21033,N_21131);
or U21371 (N_21371,N_21108,N_21013);
nand U21372 (N_21372,N_21169,N_21163);
and U21373 (N_21373,N_21153,N_21013);
or U21374 (N_21374,N_21065,N_21045);
and U21375 (N_21375,N_21096,N_21112);
or U21376 (N_21376,N_21166,N_21049);
and U21377 (N_21377,N_21001,N_21004);
or U21378 (N_21378,N_21192,N_21151);
nor U21379 (N_21379,N_21182,N_21009);
or U21380 (N_21380,N_21084,N_21138);
or U21381 (N_21381,N_21140,N_21087);
or U21382 (N_21382,N_21083,N_21057);
or U21383 (N_21383,N_21126,N_21175);
and U21384 (N_21384,N_21061,N_21147);
nand U21385 (N_21385,N_21183,N_21142);
nand U21386 (N_21386,N_21097,N_21029);
and U21387 (N_21387,N_21155,N_21015);
or U21388 (N_21388,N_21003,N_21031);
nand U21389 (N_21389,N_21101,N_21149);
and U21390 (N_21390,N_21012,N_21076);
and U21391 (N_21391,N_21161,N_21158);
and U21392 (N_21392,N_21169,N_21131);
nor U21393 (N_21393,N_21174,N_21042);
nor U21394 (N_21394,N_21062,N_21050);
and U21395 (N_21395,N_21078,N_21093);
nand U21396 (N_21396,N_21102,N_21118);
nor U21397 (N_21397,N_21133,N_21197);
xor U21398 (N_21398,N_21044,N_21161);
or U21399 (N_21399,N_21052,N_21061);
nand U21400 (N_21400,N_21289,N_21278);
nand U21401 (N_21401,N_21388,N_21251);
and U21402 (N_21402,N_21305,N_21373);
or U21403 (N_21403,N_21262,N_21308);
nand U21404 (N_21404,N_21304,N_21383);
or U21405 (N_21405,N_21212,N_21232);
and U21406 (N_21406,N_21258,N_21244);
nand U21407 (N_21407,N_21378,N_21322);
or U21408 (N_21408,N_21276,N_21353);
nand U21409 (N_21409,N_21303,N_21345);
nor U21410 (N_21410,N_21346,N_21341);
nand U21411 (N_21411,N_21310,N_21386);
or U21412 (N_21412,N_21285,N_21270);
nor U21413 (N_21413,N_21209,N_21249);
nand U21414 (N_21414,N_21274,N_21288);
or U21415 (N_21415,N_21349,N_21313);
nand U21416 (N_21416,N_21290,N_21306);
nor U21417 (N_21417,N_21340,N_21237);
or U21418 (N_21418,N_21375,N_21355);
or U21419 (N_21419,N_21217,N_21216);
and U21420 (N_21420,N_21269,N_21362);
or U21421 (N_21421,N_21339,N_21256);
nand U21422 (N_21422,N_21384,N_21297);
and U21423 (N_21423,N_21202,N_21321);
or U21424 (N_21424,N_21371,N_21385);
and U21425 (N_21425,N_21343,N_21268);
and U21426 (N_21426,N_21380,N_21215);
nor U21427 (N_21427,N_21358,N_21391);
or U21428 (N_21428,N_21365,N_21210);
or U21429 (N_21429,N_21281,N_21377);
and U21430 (N_21430,N_21267,N_21379);
and U21431 (N_21431,N_21337,N_21243);
or U21432 (N_21432,N_21300,N_21245);
or U21433 (N_21433,N_21361,N_21374);
and U21434 (N_21434,N_21253,N_21309);
nor U21435 (N_21435,N_21342,N_21208);
or U21436 (N_21436,N_21221,N_21330);
nor U21437 (N_21437,N_21204,N_21318);
nor U21438 (N_21438,N_21236,N_21273);
nand U21439 (N_21439,N_21316,N_21201);
or U21440 (N_21440,N_21338,N_21241);
and U21441 (N_21441,N_21364,N_21296);
and U21442 (N_21442,N_21298,N_21291);
and U21443 (N_21443,N_21336,N_21360);
nand U21444 (N_21444,N_21226,N_21248);
or U21445 (N_21445,N_21246,N_21206);
nor U21446 (N_21446,N_21302,N_21282);
nor U21447 (N_21447,N_21266,N_21240);
nor U21448 (N_21448,N_21219,N_21222);
nor U21449 (N_21449,N_21272,N_21214);
and U21450 (N_21450,N_21294,N_21223);
and U21451 (N_21451,N_21315,N_21354);
nand U21452 (N_21452,N_21363,N_21367);
and U21453 (N_21453,N_21234,N_21277);
and U21454 (N_21454,N_21356,N_21242);
and U21455 (N_21455,N_21327,N_21397);
and U21456 (N_21456,N_21334,N_21359);
and U21457 (N_21457,N_21366,N_21254);
nor U21458 (N_21458,N_21200,N_21252);
and U21459 (N_21459,N_21311,N_21392);
and U21460 (N_21460,N_21283,N_21275);
and U21461 (N_21461,N_21207,N_21324);
or U21462 (N_21462,N_21229,N_21329);
and U21463 (N_21463,N_21319,N_21260);
nand U21464 (N_21464,N_21203,N_21331);
or U21465 (N_21465,N_21328,N_21286);
nor U21466 (N_21466,N_21265,N_21227);
and U21467 (N_21467,N_21398,N_21352);
nor U21468 (N_21468,N_21280,N_21394);
nand U21469 (N_21469,N_21351,N_21213);
or U21470 (N_21470,N_21368,N_21399);
or U21471 (N_21471,N_21225,N_21261);
and U21472 (N_21472,N_21325,N_21332);
or U21473 (N_21473,N_21220,N_21357);
or U21474 (N_21474,N_21271,N_21382);
and U21475 (N_21475,N_21228,N_21333);
and U21476 (N_21476,N_21259,N_21369);
or U21477 (N_21477,N_21307,N_21299);
nor U21478 (N_21478,N_21370,N_21247);
or U21479 (N_21479,N_21372,N_21292);
and U21480 (N_21480,N_21317,N_21395);
nor U21481 (N_21481,N_21393,N_21344);
and U21482 (N_21482,N_21314,N_21287);
nor U21483 (N_21483,N_21224,N_21205);
and U21484 (N_21484,N_21293,N_21211);
nand U21485 (N_21485,N_21250,N_21257);
and U21486 (N_21486,N_21239,N_21312);
or U21487 (N_21487,N_21279,N_21233);
nand U21488 (N_21488,N_21348,N_21381);
nor U21489 (N_21489,N_21235,N_21347);
nor U21490 (N_21490,N_21389,N_21396);
and U21491 (N_21491,N_21231,N_21387);
nor U21492 (N_21492,N_21284,N_21301);
and U21493 (N_21493,N_21264,N_21390);
nor U21494 (N_21494,N_21255,N_21326);
nor U21495 (N_21495,N_21238,N_21323);
nand U21496 (N_21496,N_21295,N_21320);
nand U21497 (N_21497,N_21335,N_21350);
and U21498 (N_21498,N_21230,N_21376);
nand U21499 (N_21499,N_21263,N_21218);
or U21500 (N_21500,N_21337,N_21332);
and U21501 (N_21501,N_21310,N_21352);
nor U21502 (N_21502,N_21255,N_21390);
and U21503 (N_21503,N_21374,N_21279);
nor U21504 (N_21504,N_21321,N_21372);
or U21505 (N_21505,N_21224,N_21362);
and U21506 (N_21506,N_21305,N_21376);
nor U21507 (N_21507,N_21341,N_21308);
or U21508 (N_21508,N_21298,N_21350);
or U21509 (N_21509,N_21386,N_21290);
and U21510 (N_21510,N_21328,N_21232);
nand U21511 (N_21511,N_21204,N_21216);
nor U21512 (N_21512,N_21384,N_21361);
or U21513 (N_21513,N_21389,N_21363);
or U21514 (N_21514,N_21326,N_21206);
nand U21515 (N_21515,N_21230,N_21327);
and U21516 (N_21516,N_21364,N_21299);
or U21517 (N_21517,N_21384,N_21244);
and U21518 (N_21518,N_21358,N_21366);
xor U21519 (N_21519,N_21394,N_21242);
or U21520 (N_21520,N_21270,N_21393);
nand U21521 (N_21521,N_21345,N_21290);
nand U21522 (N_21522,N_21288,N_21233);
and U21523 (N_21523,N_21354,N_21341);
nand U21524 (N_21524,N_21313,N_21385);
or U21525 (N_21525,N_21366,N_21302);
and U21526 (N_21526,N_21358,N_21228);
nor U21527 (N_21527,N_21218,N_21277);
and U21528 (N_21528,N_21301,N_21374);
nor U21529 (N_21529,N_21210,N_21213);
or U21530 (N_21530,N_21392,N_21339);
and U21531 (N_21531,N_21346,N_21205);
nand U21532 (N_21532,N_21314,N_21305);
nand U21533 (N_21533,N_21282,N_21297);
nor U21534 (N_21534,N_21210,N_21230);
nand U21535 (N_21535,N_21367,N_21329);
and U21536 (N_21536,N_21229,N_21360);
nor U21537 (N_21537,N_21380,N_21289);
and U21538 (N_21538,N_21229,N_21251);
or U21539 (N_21539,N_21237,N_21256);
or U21540 (N_21540,N_21254,N_21231);
nor U21541 (N_21541,N_21228,N_21206);
nor U21542 (N_21542,N_21331,N_21384);
nor U21543 (N_21543,N_21266,N_21358);
or U21544 (N_21544,N_21382,N_21207);
and U21545 (N_21545,N_21303,N_21359);
and U21546 (N_21546,N_21357,N_21372);
nand U21547 (N_21547,N_21340,N_21382);
or U21548 (N_21548,N_21256,N_21312);
and U21549 (N_21549,N_21308,N_21230);
nand U21550 (N_21550,N_21305,N_21285);
and U21551 (N_21551,N_21352,N_21388);
and U21552 (N_21552,N_21230,N_21381);
or U21553 (N_21553,N_21364,N_21274);
or U21554 (N_21554,N_21351,N_21222);
and U21555 (N_21555,N_21364,N_21271);
or U21556 (N_21556,N_21363,N_21271);
nand U21557 (N_21557,N_21399,N_21299);
nand U21558 (N_21558,N_21279,N_21394);
or U21559 (N_21559,N_21290,N_21324);
or U21560 (N_21560,N_21394,N_21284);
and U21561 (N_21561,N_21358,N_21265);
nor U21562 (N_21562,N_21393,N_21331);
nor U21563 (N_21563,N_21259,N_21301);
or U21564 (N_21564,N_21319,N_21373);
nor U21565 (N_21565,N_21239,N_21270);
or U21566 (N_21566,N_21380,N_21268);
nor U21567 (N_21567,N_21245,N_21264);
nand U21568 (N_21568,N_21222,N_21262);
and U21569 (N_21569,N_21232,N_21312);
nand U21570 (N_21570,N_21231,N_21204);
or U21571 (N_21571,N_21266,N_21208);
nand U21572 (N_21572,N_21262,N_21390);
nand U21573 (N_21573,N_21222,N_21325);
nand U21574 (N_21574,N_21213,N_21329);
and U21575 (N_21575,N_21391,N_21394);
and U21576 (N_21576,N_21341,N_21350);
or U21577 (N_21577,N_21239,N_21282);
and U21578 (N_21578,N_21246,N_21335);
or U21579 (N_21579,N_21316,N_21202);
or U21580 (N_21580,N_21369,N_21258);
nand U21581 (N_21581,N_21368,N_21245);
and U21582 (N_21582,N_21362,N_21226);
or U21583 (N_21583,N_21301,N_21364);
nand U21584 (N_21584,N_21313,N_21334);
nand U21585 (N_21585,N_21268,N_21261);
or U21586 (N_21586,N_21356,N_21341);
xnor U21587 (N_21587,N_21275,N_21248);
nor U21588 (N_21588,N_21368,N_21361);
and U21589 (N_21589,N_21328,N_21397);
and U21590 (N_21590,N_21318,N_21220);
and U21591 (N_21591,N_21304,N_21371);
nor U21592 (N_21592,N_21273,N_21281);
nor U21593 (N_21593,N_21265,N_21341);
and U21594 (N_21594,N_21392,N_21233);
nand U21595 (N_21595,N_21291,N_21249);
or U21596 (N_21596,N_21288,N_21258);
or U21597 (N_21597,N_21229,N_21258);
or U21598 (N_21598,N_21313,N_21368);
or U21599 (N_21599,N_21257,N_21379);
or U21600 (N_21600,N_21434,N_21472);
nand U21601 (N_21601,N_21569,N_21429);
nor U21602 (N_21602,N_21437,N_21425);
nand U21603 (N_21603,N_21498,N_21465);
or U21604 (N_21604,N_21448,N_21418);
or U21605 (N_21605,N_21409,N_21497);
and U21606 (N_21606,N_21536,N_21502);
or U21607 (N_21607,N_21424,N_21401);
or U21608 (N_21608,N_21572,N_21592);
and U21609 (N_21609,N_21556,N_21526);
and U21610 (N_21610,N_21438,N_21552);
or U21611 (N_21611,N_21520,N_21451);
and U21612 (N_21612,N_21554,N_21488);
or U21613 (N_21613,N_21586,N_21478);
nand U21614 (N_21614,N_21486,N_21559);
nor U21615 (N_21615,N_21583,N_21585);
or U21616 (N_21616,N_21582,N_21435);
and U21617 (N_21617,N_21541,N_21504);
nor U21618 (N_21618,N_21514,N_21473);
or U21619 (N_21619,N_21519,N_21527);
and U21620 (N_21620,N_21494,N_21469);
nor U21621 (N_21621,N_21579,N_21479);
nor U21622 (N_21622,N_21551,N_21561);
and U21623 (N_21623,N_21443,N_21470);
or U21624 (N_21624,N_21593,N_21450);
and U21625 (N_21625,N_21464,N_21462);
nand U21626 (N_21626,N_21542,N_21534);
or U21627 (N_21627,N_21512,N_21532);
nor U21628 (N_21628,N_21510,N_21524);
or U21629 (N_21629,N_21525,N_21528);
and U21630 (N_21630,N_21531,N_21405);
or U21631 (N_21631,N_21463,N_21505);
nor U21632 (N_21632,N_21508,N_21454);
and U21633 (N_21633,N_21589,N_21545);
and U21634 (N_21634,N_21546,N_21402);
and U21635 (N_21635,N_21557,N_21482);
nand U21636 (N_21636,N_21491,N_21408);
nor U21637 (N_21637,N_21460,N_21596);
and U21638 (N_21638,N_21456,N_21550);
nor U21639 (N_21639,N_21446,N_21417);
and U21640 (N_21640,N_21507,N_21477);
nor U21641 (N_21641,N_21598,N_21544);
nor U21642 (N_21642,N_21495,N_21447);
or U21643 (N_21643,N_21407,N_21576);
and U21644 (N_21644,N_21501,N_21474);
nor U21645 (N_21645,N_21577,N_21578);
nor U21646 (N_21646,N_21433,N_21499);
and U21647 (N_21647,N_21471,N_21436);
nor U21648 (N_21648,N_21580,N_21500);
nor U21649 (N_21649,N_21573,N_21503);
or U21650 (N_21650,N_21420,N_21419);
nor U21651 (N_21651,N_21530,N_21410);
and U21652 (N_21652,N_21571,N_21567);
nand U21653 (N_21653,N_21404,N_21412);
or U21654 (N_21654,N_21568,N_21475);
nand U21655 (N_21655,N_21584,N_21476);
or U21656 (N_21656,N_21575,N_21485);
nor U21657 (N_21657,N_21518,N_21467);
nand U21658 (N_21658,N_21558,N_21509);
nor U21659 (N_21659,N_21427,N_21513);
nor U21660 (N_21660,N_21432,N_21423);
or U21661 (N_21661,N_21445,N_21588);
or U21662 (N_21662,N_21547,N_21483);
nor U21663 (N_21663,N_21440,N_21400);
nor U21664 (N_21664,N_21529,N_21493);
nand U21665 (N_21665,N_21422,N_21539);
or U21666 (N_21666,N_21516,N_21564);
nand U21667 (N_21667,N_21570,N_21587);
and U21668 (N_21668,N_21549,N_21565);
nand U21669 (N_21669,N_21406,N_21459);
or U21670 (N_21670,N_21449,N_21597);
nand U21671 (N_21671,N_21574,N_21444);
or U21672 (N_21672,N_21431,N_21413);
or U21673 (N_21673,N_21492,N_21535);
and U21674 (N_21674,N_21453,N_21411);
or U21675 (N_21675,N_21555,N_21458);
and U21676 (N_21676,N_21562,N_21428);
and U21677 (N_21677,N_21511,N_21538);
nand U21678 (N_21678,N_21415,N_21457);
nor U21679 (N_21679,N_21533,N_21506);
or U21680 (N_21680,N_21416,N_21487);
nor U21681 (N_21681,N_21439,N_21548);
and U21682 (N_21682,N_21403,N_21414);
and U21683 (N_21683,N_21523,N_21481);
or U21684 (N_21684,N_21461,N_21484);
nor U21685 (N_21685,N_21591,N_21468);
nand U21686 (N_21686,N_21563,N_21590);
nor U21687 (N_21687,N_21452,N_21515);
and U21688 (N_21688,N_21599,N_21553);
nor U21689 (N_21689,N_21466,N_21489);
nand U21690 (N_21690,N_21490,N_21430);
nor U21691 (N_21691,N_21517,N_21496);
or U21692 (N_21692,N_21543,N_21566);
nand U21693 (N_21693,N_21540,N_21581);
and U21694 (N_21694,N_21480,N_21442);
and U21695 (N_21695,N_21421,N_21441);
nor U21696 (N_21696,N_21560,N_21521);
and U21697 (N_21697,N_21455,N_21595);
or U21698 (N_21698,N_21426,N_21537);
and U21699 (N_21699,N_21522,N_21594);
or U21700 (N_21700,N_21476,N_21519);
or U21701 (N_21701,N_21479,N_21443);
nand U21702 (N_21702,N_21557,N_21425);
and U21703 (N_21703,N_21509,N_21536);
nand U21704 (N_21704,N_21421,N_21482);
or U21705 (N_21705,N_21527,N_21402);
xnor U21706 (N_21706,N_21423,N_21404);
nor U21707 (N_21707,N_21539,N_21573);
or U21708 (N_21708,N_21447,N_21439);
and U21709 (N_21709,N_21552,N_21496);
and U21710 (N_21710,N_21544,N_21595);
xor U21711 (N_21711,N_21584,N_21599);
or U21712 (N_21712,N_21573,N_21576);
nor U21713 (N_21713,N_21517,N_21526);
nand U21714 (N_21714,N_21520,N_21584);
or U21715 (N_21715,N_21462,N_21448);
and U21716 (N_21716,N_21563,N_21507);
and U21717 (N_21717,N_21577,N_21413);
or U21718 (N_21718,N_21417,N_21509);
or U21719 (N_21719,N_21587,N_21425);
nor U21720 (N_21720,N_21492,N_21408);
or U21721 (N_21721,N_21530,N_21409);
or U21722 (N_21722,N_21527,N_21566);
or U21723 (N_21723,N_21503,N_21534);
nor U21724 (N_21724,N_21489,N_21505);
nand U21725 (N_21725,N_21416,N_21562);
and U21726 (N_21726,N_21504,N_21501);
nor U21727 (N_21727,N_21544,N_21537);
nor U21728 (N_21728,N_21489,N_21593);
nor U21729 (N_21729,N_21468,N_21440);
or U21730 (N_21730,N_21417,N_21410);
nor U21731 (N_21731,N_21580,N_21450);
nand U21732 (N_21732,N_21506,N_21507);
or U21733 (N_21733,N_21432,N_21516);
nor U21734 (N_21734,N_21483,N_21429);
and U21735 (N_21735,N_21479,N_21591);
nor U21736 (N_21736,N_21452,N_21421);
or U21737 (N_21737,N_21462,N_21482);
or U21738 (N_21738,N_21485,N_21544);
and U21739 (N_21739,N_21474,N_21530);
and U21740 (N_21740,N_21581,N_21404);
nand U21741 (N_21741,N_21556,N_21409);
nor U21742 (N_21742,N_21559,N_21498);
and U21743 (N_21743,N_21502,N_21549);
nand U21744 (N_21744,N_21529,N_21497);
or U21745 (N_21745,N_21521,N_21495);
or U21746 (N_21746,N_21443,N_21453);
and U21747 (N_21747,N_21519,N_21571);
nand U21748 (N_21748,N_21567,N_21422);
and U21749 (N_21749,N_21447,N_21416);
or U21750 (N_21750,N_21495,N_21524);
or U21751 (N_21751,N_21487,N_21465);
or U21752 (N_21752,N_21496,N_21599);
or U21753 (N_21753,N_21481,N_21435);
or U21754 (N_21754,N_21532,N_21554);
and U21755 (N_21755,N_21526,N_21427);
nor U21756 (N_21756,N_21502,N_21591);
nor U21757 (N_21757,N_21455,N_21490);
and U21758 (N_21758,N_21568,N_21485);
or U21759 (N_21759,N_21556,N_21536);
nor U21760 (N_21760,N_21453,N_21540);
or U21761 (N_21761,N_21518,N_21582);
xor U21762 (N_21762,N_21438,N_21406);
or U21763 (N_21763,N_21580,N_21484);
or U21764 (N_21764,N_21460,N_21568);
nand U21765 (N_21765,N_21558,N_21518);
or U21766 (N_21766,N_21581,N_21437);
and U21767 (N_21767,N_21411,N_21485);
nor U21768 (N_21768,N_21450,N_21516);
nand U21769 (N_21769,N_21450,N_21590);
and U21770 (N_21770,N_21506,N_21534);
or U21771 (N_21771,N_21494,N_21457);
or U21772 (N_21772,N_21583,N_21558);
or U21773 (N_21773,N_21570,N_21493);
and U21774 (N_21774,N_21450,N_21549);
nor U21775 (N_21775,N_21463,N_21460);
nand U21776 (N_21776,N_21429,N_21460);
nand U21777 (N_21777,N_21461,N_21506);
nand U21778 (N_21778,N_21414,N_21519);
or U21779 (N_21779,N_21509,N_21412);
and U21780 (N_21780,N_21452,N_21598);
nand U21781 (N_21781,N_21436,N_21408);
or U21782 (N_21782,N_21415,N_21564);
or U21783 (N_21783,N_21422,N_21472);
nand U21784 (N_21784,N_21477,N_21525);
nand U21785 (N_21785,N_21497,N_21511);
nand U21786 (N_21786,N_21405,N_21402);
and U21787 (N_21787,N_21525,N_21506);
and U21788 (N_21788,N_21501,N_21423);
or U21789 (N_21789,N_21417,N_21440);
nor U21790 (N_21790,N_21428,N_21571);
or U21791 (N_21791,N_21449,N_21599);
nand U21792 (N_21792,N_21503,N_21561);
nand U21793 (N_21793,N_21418,N_21583);
and U21794 (N_21794,N_21583,N_21450);
or U21795 (N_21795,N_21463,N_21536);
or U21796 (N_21796,N_21556,N_21545);
and U21797 (N_21797,N_21534,N_21567);
and U21798 (N_21798,N_21562,N_21493);
nor U21799 (N_21799,N_21555,N_21587);
or U21800 (N_21800,N_21794,N_21755);
nor U21801 (N_21801,N_21674,N_21733);
nor U21802 (N_21802,N_21691,N_21738);
nand U21803 (N_21803,N_21688,N_21641);
and U21804 (N_21804,N_21721,N_21769);
nor U21805 (N_21805,N_21763,N_21671);
nor U21806 (N_21806,N_21609,N_21726);
or U21807 (N_21807,N_21635,N_21602);
nand U21808 (N_21808,N_21631,N_21613);
or U21809 (N_21809,N_21686,N_21772);
nor U21810 (N_21810,N_21665,N_21657);
nor U21811 (N_21811,N_21681,N_21714);
or U21812 (N_21812,N_21630,N_21709);
or U21813 (N_21813,N_21797,N_21679);
xor U21814 (N_21814,N_21642,N_21699);
nor U21815 (N_21815,N_21713,N_21718);
or U21816 (N_21816,N_21644,N_21742);
nand U21817 (N_21817,N_21623,N_21637);
or U21818 (N_21818,N_21778,N_21664);
or U21819 (N_21819,N_21711,N_21694);
or U21820 (N_21820,N_21650,N_21689);
nand U21821 (N_21821,N_21608,N_21678);
or U21822 (N_21822,N_21632,N_21607);
or U21823 (N_21823,N_21649,N_21652);
nor U21824 (N_21824,N_21698,N_21676);
or U21825 (N_21825,N_21616,N_21728);
or U21826 (N_21826,N_21750,N_21793);
nor U21827 (N_21827,N_21754,N_21775);
and U21828 (N_21828,N_21760,N_21693);
or U21829 (N_21829,N_21682,N_21612);
nor U21830 (N_21830,N_21625,N_21670);
nand U21831 (N_21831,N_21675,N_21727);
and U21832 (N_21832,N_21606,N_21618);
nand U21833 (N_21833,N_21791,N_21747);
or U21834 (N_21834,N_21774,N_21777);
or U21835 (N_21835,N_21725,N_21740);
or U21836 (N_21836,N_21767,N_21729);
or U21837 (N_21837,N_21762,N_21704);
nor U21838 (N_21838,N_21759,N_21716);
nand U21839 (N_21839,N_21666,N_21601);
nand U21840 (N_21840,N_21799,N_21603);
nor U21841 (N_21841,N_21661,N_21781);
nor U21842 (N_21842,N_21614,N_21706);
and U21843 (N_21843,N_21771,N_21605);
nor U21844 (N_21844,N_21654,N_21796);
and U21845 (N_21845,N_21707,N_21786);
and U21846 (N_21846,N_21627,N_21667);
nor U21847 (N_21847,N_21732,N_21708);
nand U21848 (N_21848,N_21756,N_21792);
and U21849 (N_21849,N_21722,N_21701);
or U21850 (N_21850,N_21735,N_21761);
or U21851 (N_21851,N_21651,N_21672);
and U21852 (N_21852,N_21749,N_21684);
and U21853 (N_21853,N_21783,N_21653);
nor U21854 (N_21854,N_21787,N_21734);
nor U21855 (N_21855,N_21628,N_21660);
and U21856 (N_21856,N_21638,N_21739);
nor U21857 (N_21857,N_21798,N_21604);
or U21858 (N_21858,N_21695,N_21622);
nor U21859 (N_21859,N_21719,N_21626);
nor U21860 (N_21860,N_21776,N_21692);
and U21861 (N_21861,N_21745,N_21668);
nor U21862 (N_21862,N_21615,N_21677);
nor U21863 (N_21863,N_21766,N_21753);
nor U21864 (N_21864,N_21751,N_21789);
or U21865 (N_21865,N_21737,N_21683);
nand U21866 (N_21866,N_21770,N_21785);
and U21867 (N_21867,N_21700,N_21712);
nor U21868 (N_21868,N_21647,N_21768);
nand U21869 (N_21869,N_21629,N_21784);
nand U21870 (N_21870,N_21648,N_21658);
nor U21871 (N_21871,N_21743,N_21780);
nand U21872 (N_21872,N_21752,N_21639);
or U21873 (N_21873,N_21710,N_21673);
nor U21874 (N_21874,N_21720,N_21619);
and U21875 (N_21875,N_21782,N_21773);
and U21876 (N_21876,N_21788,N_21633);
or U21877 (N_21877,N_21731,N_21663);
or U21878 (N_21878,N_21705,N_21600);
nor U21879 (N_21879,N_21640,N_21757);
nor U21880 (N_21880,N_21645,N_21715);
and U21881 (N_21881,N_21643,N_21723);
nand U21882 (N_21882,N_21636,N_21779);
and U21883 (N_21883,N_21659,N_21611);
nor U21884 (N_21884,N_21610,N_21617);
and U21885 (N_21885,N_21736,N_21655);
nor U21886 (N_21886,N_21741,N_21680);
nand U21887 (N_21887,N_21687,N_21634);
and U21888 (N_21888,N_21746,N_21764);
or U21889 (N_21889,N_21748,N_21765);
nand U21890 (N_21890,N_21621,N_21685);
and U21891 (N_21891,N_21744,N_21724);
or U21892 (N_21892,N_21620,N_21758);
nor U21893 (N_21893,N_21646,N_21795);
or U21894 (N_21894,N_21717,N_21790);
or U21895 (N_21895,N_21662,N_21697);
and U21896 (N_21896,N_21703,N_21702);
nand U21897 (N_21897,N_21669,N_21624);
nand U21898 (N_21898,N_21730,N_21656);
nand U21899 (N_21899,N_21690,N_21696);
and U21900 (N_21900,N_21750,N_21728);
or U21901 (N_21901,N_21607,N_21750);
nand U21902 (N_21902,N_21770,N_21692);
nand U21903 (N_21903,N_21644,N_21665);
and U21904 (N_21904,N_21763,N_21704);
nand U21905 (N_21905,N_21720,N_21663);
nor U21906 (N_21906,N_21782,N_21776);
nor U21907 (N_21907,N_21686,N_21756);
nor U21908 (N_21908,N_21778,N_21680);
nor U21909 (N_21909,N_21628,N_21614);
or U21910 (N_21910,N_21761,N_21675);
and U21911 (N_21911,N_21743,N_21685);
nand U21912 (N_21912,N_21607,N_21693);
or U21913 (N_21913,N_21798,N_21626);
or U21914 (N_21914,N_21678,N_21697);
nor U21915 (N_21915,N_21628,N_21698);
nand U21916 (N_21916,N_21748,N_21678);
or U21917 (N_21917,N_21657,N_21654);
and U21918 (N_21918,N_21718,N_21772);
or U21919 (N_21919,N_21700,N_21710);
or U21920 (N_21920,N_21619,N_21711);
and U21921 (N_21921,N_21601,N_21776);
xnor U21922 (N_21922,N_21648,N_21675);
nor U21923 (N_21923,N_21652,N_21682);
or U21924 (N_21924,N_21613,N_21726);
or U21925 (N_21925,N_21611,N_21679);
nor U21926 (N_21926,N_21741,N_21744);
or U21927 (N_21927,N_21777,N_21658);
nand U21928 (N_21928,N_21627,N_21630);
nor U21929 (N_21929,N_21694,N_21735);
and U21930 (N_21930,N_21642,N_21785);
nand U21931 (N_21931,N_21600,N_21685);
xor U21932 (N_21932,N_21636,N_21743);
and U21933 (N_21933,N_21652,N_21621);
nor U21934 (N_21934,N_21770,N_21635);
or U21935 (N_21935,N_21689,N_21626);
nor U21936 (N_21936,N_21649,N_21725);
nand U21937 (N_21937,N_21693,N_21704);
nor U21938 (N_21938,N_21724,N_21772);
nand U21939 (N_21939,N_21720,N_21729);
and U21940 (N_21940,N_21787,N_21791);
or U21941 (N_21941,N_21678,N_21620);
nand U21942 (N_21942,N_21657,N_21672);
nand U21943 (N_21943,N_21690,N_21725);
nor U21944 (N_21944,N_21716,N_21795);
nor U21945 (N_21945,N_21697,N_21772);
and U21946 (N_21946,N_21762,N_21680);
nor U21947 (N_21947,N_21788,N_21694);
nand U21948 (N_21948,N_21695,N_21771);
and U21949 (N_21949,N_21759,N_21672);
or U21950 (N_21950,N_21683,N_21642);
and U21951 (N_21951,N_21623,N_21667);
or U21952 (N_21952,N_21758,N_21702);
nor U21953 (N_21953,N_21659,N_21658);
or U21954 (N_21954,N_21692,N_21683);
nand U21955 (N_21955,N_21630,N_21675);
and U21956 (N_21956,N_21774,N_21797);
nor U21957 (N_21957,N_21794,N_21607);
or U21958 (N_21958,N_21670,N_21647);
or U21959 (N_21959,N_21703,N_21665);
nor U21960 (N_21960,N_21731,N_21660);
and U21961 (N_21961,N_21601,N_21627);
and U21962 (N_21962,N_21602,N_21622);
or U21963 (N_21963,N_21784,N_21777);
nand U21964 (N_21964,N_21706,N_21770);
and U21965 (N_21965,N_21691,N_21730);
or U21966 (N_21966,N_21765,N_21636);
and U21967 (N_21967,N_21735,N_21616);
and U21968 (N_21968,N_21711,N_21768);
nand U21969 (N_21969,N_21676,N_21729);
or U21970 (N_21970,N_21710,N_21621);
nor U21971 (N_21971,N_21655,N_21700);
and U21972 (N_21972,N_21640,N_21630);
nor U21973 (N_21973,N_21788,N_21796);
nor U21974 (N_21974,N_21760,N_21710);
nor U21975 (N_21975,N_21686,N_21603);
or U21976 (N_21976,N_21639,N_21660);
nand U21977 (N_21977,N_21746,N_21783);
nor U21978 (N_21978,N_21688,N_21707);
nand U21979 (N_21979,N_21740,N_21698);
or U21980 (N_21980,N_21707,N_21797);
nand U21981 (N_21981,N_21748,N_21743);
or U21982 (N_21982,N_21779,N_21673);
nor U21983 (N_21983,N_21760,N_21713);
nor U21984 (N_21984,N_21779,N_21642);
nand U21985 (N_21985,N_21690,N_21665);
and U21986 (N_21986,N_21788,N_21639);
nand U21987 (N_21987,N_21693,N_21663);
nand U21988 (N_21988,N_21790,N_21772);
and U21989 (N_21989,N_21607,N_21630);
nor U21990 (N_21990,N_21773,N_21699);
nor U21991 (N_21991,N_21663,N_21616);
nor U21992 (N_21992,N_21697,N_21698);
and U21993 (N_21993,N_21745,N_21722);
nor U21994 (N_21994,N_21694,N_21636);
nor U21995 (N_21995,N_21659,N_21650);
nor U21996 (N_21996,N_21667,N_21679);
nand U21997 (N_21997,N_21725,N_21673);
or U21998 (N_21998,N_21602,N_21614);
or U21999 (N_21999,N_21736,N_21616);
and U22000 (N_22000,N_21826,N_21839);
or U22001 (N_22001,N_21999,N_21842);
and U22002 (N_22002,N_21963,N_21947);
or U22003 (N_22003,N_21880,N_21968);
or U22004 (N_22004,N_21894,N_21971);
and U22005 (N_22005,N_21828,N_21917);
nor U22006 (N_22006,N_21812,N_21970);
and U22007 (N_22007,N_21984,N_21909);
or U22008 (N_22008,N_21813,N_21902);
nor U22009 (N_22009,N_21822,N_21884);
nor U22010 (N_22010,N_21879,N_21997);
nor U22011 (N_22011,N_21849,N_21921);
nand U22012 (N_22012,N_21843,N_21919);
or U22013 (N_22013,N_21885,N_21900);
nor U22014 (N_22014,N_21960,N_21941);
nand U22015 (N_22015,N_21804,N_21993);
nand U22016 (N_22016,N_21867,N_21852);
and U22017 (N_22017,N_21801,N_21950);
nand U22018 (N_22018,N_21987,N_21864);
or U22019 (N_22019,N_21914,N_21929);
nor U22020 (N_22020,N_21996,N_21943);
and U22021 (N_22021,N_21868,N_21861);
xor U22022 (N_22022,N_21860,N_21969);
or U22023 (N_22023,N_21892,N_21815);
or U22024 (N_22024,N_21944,N_21857);
or U22025 (N_22025,N_21869,N_21962);
nand U22026 (N_22026,N_21800,N_21928);
nor U22027 (N_22027,N_21827,N_21859);
nand U22028 (N_22028,N_21851,N_21817);
nand U22029 (N_22029,N_21846,N_21854);
nand U22030 (N_22030,N_21973,N_21953);
or U22031 (N_22031,N_21856,N_21980);
and U22032 (N_22032,N_21871,N_21954);
and U22033 (N_22033,N_21844,N_21904);
and U22034 (N_22034,N_21898,N_21937);
or U22035 (N_22035,N_21916,N_21865);
nand U22036 (N_22036,N_21903,N_21994);
nor U22037 (N_22037,N_21926,N_21887);
nor U22038 (N_22038,N_21870,N_21949);
or U22039 (N_22039,N_21818,N_21920);
nand U22040 (N_22040,N_21823,N_21991);
nand U22041 (N_22041,N_21875,N_21932);
or U22042 (N_22042,N_21803,N_21862);
and U22043 (N_22043,N_21811,N_21893);
or U22044 (N_22044,N_21866,N_21863);
or U22045 (N_22045,N_21907,N_21913);
nand U22046 (N_22046,N_21830,N_21981);
nand U22047 (N_22047,N_21837,N_21967);
or U22048 (N_22048,N_21848,N_21992);
and U22049 (N_22049,N_21995,N_21912);
and U22050 (N_22050,N_21957,N_21936);
nor U22051 (N_22051,N_21964,N_21986);
nor U22052 (N_22052,N_21922,N_21972);
or U22053 (N_22053,N_21891,N_21850);
nor U22054 (N_22054,N_21908,N_21935);
nor U22055 (N_22055,N_21877,N_21951);
nor U22056 (N_22056,N_21940,N_21858);
and U22057 (N_22057,N_21910,N_21924);
and U22058 (N_22058,N_21878,N_21965);
and U22059 (N_22059,N_21821,N_21853);
nor U22060 (N_22060,N_21927,N_21840);
nor U22061 (N_22061,N_21874,N_21808);
nor U22062 (N_22062,N_21883,N_21923);
nand U22063 (N_22063,N_21959,N_21855);
nor U22064 (N_22064,N_21974,N_21825);
and U22065 (N_22065,N_21824,N_21841);
nand U22066 (N_22066,N_21989,N_21966);
nor U22067 (N_22067,N_21925,N_21977);
or U22068 (N_22068,N_21905,N_21948);
or U22069 (N_22069,N_21814,N_21901);
and U22070 (N_22070,N_21835,N_21881);
nor U22071 (N_22071,N_21895,N_21831);
nand U22072 (N_22072,N_21847,N_21930);
nand U22073 (N_22073,N_21888,N_21956);
or U22074 (N_22074,N_21942,N_21873);
or U22075 (N_22075,N_21938,N_21988);
nor U22076 (N_22076,N_21899,N_21805);
xor U22077 (N_22077,N_21998,N_21889);
and U22078 (N_22078,N_21985,N_21890);
nand U22079 (N_22079,N_21975,N_21906);
nand U22080 (N_22080,N_21809,N_21836);
nand U22081 (N_22081,N_21918,N_21806);
and U22082 (N_22082,N_21829,N_21946);
and U22083 (N_22083,N_21976,N_21915);
nand U22084 (N_22084,N_21931,N_21896);
nor U22085 (N_22085,N_21882,N_21945);
nor U22086 (N_22086,N_21990,N_21819);
or U22087 (N_22087,N_21886,N_21939);
nor U22088 (N_22088,N_21832,N_21876);
and U22089 (N_22089,N_21807,N_21872);
and U22090 (N_22090,N_21961,N_21952);
and U22091 (N_22091,N_21820,N_21911);
and U22092 (N_22092,N_21845,N_21838);
nor U22093 (N_22093,N_21834,N_21955);
nor U22094 (N_22094,N_21958,N_21897);
nor U22095 (N_22095,N_21983,N_21978);
or U22096 (N_22096,N_21982,N_21933);
nor U22097 (N_22097,N_21934,N_21833);
nand U22098 (N_22098,N_21810,N_21802);
and U22099 (N_22099,N_21979,N_21816);
or U22100 (N_22100,N_21849,N_21848);
nor U22101 (N_22101,N_21879,N_21822);
or U22102 (N_22102,N_21984,N_21940);
and U22103 (N_22103,N_21946,N_21882);
nor U22104 (N_22104,N_21831,N_21883);
nor U22105 (N_22105,N_21959,N_21823);
nor U22106 (N_22106,N_21863,N_21824);
or U22107 (N_22107,N_21946,N_21924);
and U22108 (N_22108,N_21913,N_21888);
or U22109 (N_22109,N_21964,N_21806);
nand U22110 (N_22110,N_21987,N_21910);
and U22111 (N_22111,N_21831,N_21995);
or U22112 (N_22112,N_21959,N_21859);
or U22113 (N_22113,N_21846,N_21912);
or U22114 (N_22114,N_21809,N_21997);
and U22115 (N_22115,N_21869,N_21997);
nor U22116 (N_22116,N_21821,N_21969);
nand U22117 (N_22117,N_21870,N_21827);
nor U22118 (N_22118,N_21893,N_21923);
nor U22119 (N_22119,N_21885,N_21809);
or U22120 (N_22120,N_21973,N_21866);
and U22121 (N_22121,N_21857,N_21981);
nor U22122 (N_22122,N_21826,N_21963);
and U22123 (N_22123,N_21838,N_21875);
or U22124 (N_22124,N_21991,N_21843);
nand U22125 (N_22125,N_21903,N_21964);
and U22126 (N_22126,N_21902,N_21895);
nand U22127 (N_22127,N_21866,N_21952);
and U22128 (N_22128,N_21819,N_21984);
or U22129 (N_22129,N_21807,N_21926);
and U22130 (N_22130,N_21941,N_21913);
and U22131 (N_22131,N_21845,N_21982);
nand U22132 (N_22132,N_21950,N_21905);
or U22133 (N_22133,N_21878,N_21830);
or U22134 (N_22134,N_21863,N_21839);
nand U22135 (N_22135,N_21962,N_21904);
nor U22136 (N_22136,N_21823,N_21885);
and U22137 (N_22137,N_21948,N_21911);
xor U22138 (N_22138,N_21979,N_21872);
nand U22139 (N_22139,N_21885,N_21901);
and U22140 (N_22140,N_21818,N_21953);
nand U22141 (N_22141,N_21846,N_21896);
and U22142 (N_22142,N_21850,N_21867);
nand U22143 (N_22143,N_21849,N_21904);
nor U22144 (N_22144,N_21807,N_21980);
nand U22145 (N_22145,N_21842,N_21884);
nand U22146 (N_22146,N_21916,N_21995);
nand U22147 (N_22147,N_21871,N_21868);
nor U22148 (N_22148,N_21929,N_21813);
xor U22149 (N_22149,N_21874,N_21931);
nor U22150 (N_22150,N_21846,N_21801);
nor U22151 (N_22151,N_21847,N_21895);
nand U22152 (N_22152,N_21835,N_21981);
or U22153 (N_22153,N_21808,N_21888);
nand U22154 (N_22154,N_21939,N_21840);
and U22155 (N_22155,N_21816,N_21855);
nor U22156 (N_22156,N_21915,N_21925);
or U22157 (N_22157,N_21933,N_21818);
nor U22158 (N_22158,N_21886,N_21806);
or U22159 (N_22159,N_21923,N_21865);
and U22160 (N_22160,N_21990,N_21939);
nor U22161 (N_22161,N_21983,N_21837);
nor U22162 (N_22162,N_21935,N_21962);
or U22163 (N_22163,N_21993,N_21932);
and U22164 (N_22164,N_21980,N_21804);
nand U22165 (N_22165,N_21981,N_21896);
nand U22166 (N_22166,N_21867,N_21917);
or U22167 (N_22167,N_21862,N_21885);
nor U22168 (N_22168,N_21864,N_21901);
nor U22169 (N_22169,N_21968,N_21970);
or U22170 (N_22170,N_21869,N_21956);
nand U22171 (N_22171,N_21883,N_21978);
or U22172 (N_22172,N_21897,N_21807);
and U22173 (N_22173,N_21907,N_21802);
nand U22174 (N_22174,N_21894,N_21827);
nor U22175 (N_22175,N_21891,N_21923);
and U22176 (N_22176,N_21917,N_21984);
and U22177 (N_22177,N_21994,N_21990);
nor U22178 (N_22178,N_21872,N_21985);
nand U22179 (N_22179,N_21932,N_21980);
nand U22180 (N_22180,N_21963,N_21919);
and U22181 (N_22181,N_21978,N_21873);
nand U22182 (N_22182,N_21853,N_21874);
nor U22183 (N_22183,N_21859,N_21847);
and U22184 (N_22184,N_21949,N_21914);
or U22185 (N_22185,N_21938,N_21863);
nor U22186 (N_22186,N_21865,N_21985);
or U22187 (N_22187,N_21937,N_21893);
or U22188 (N_22188,N_21920,N_21866);
and U22189 (N_22189,N_21929,N_21933);
nor U22190 (N_22190,N_21988,N_21911);
and U22191 (N_22191,N_21951,N_21820);
nand U22192 (N_22192,N_21870,N_21805);
nor U22193 (N_22193,N_21897,N_21869);
nand U22194 (N_22194,N_21822,N_21901);
or U22195 (N_22195,N_21831,N_21834);
and U22196 (N_22196,N_21983,N_21825);
nand U22197 (N_22197,N_21831,N_21989);
nor U22198 (N_22198,N_21841,N_21982);
and U22199 (N_22199,N_21837,N_21843);
or U22200 (N_22200,N_22007,N_22074);
nor U22201 (N_22201,N_22178,N_22153);
and U22202 (N_22202,N_22079,N_22140);
nand U22203 (N_22203,N_22134,N_22086);
and U22204 (N_22204,N_22040,N_22002);
nor U22205 (N_22205,N_22022,N_22013);
and U22206 (N_22206,N_22023,N_22073);
nor U22207 (N_22207,N_22129,N_22076);
or U22208 (N_22208,N_22052,N_22124);
and U22209 (N_22209,N_22060,N_22045);
or U22210 (N_22210,N_22097,N_22191);
nand U22211 (N_22211,N_22198,N_22151);
and U22212 (N_22212,N_22121,N_22021);
and U22213 (N_22213,N_22003,N_22020);
or U22214 (N_22214,N_22176,N_22039);
nor U22215 (N_22215,N_22179,N_22172);
nor U22216 (N_22216,N_22102,N_22113);
nand U22217 (N_22217,N_22085,N_22148);
and U22218 (N_22218,N_22037,N_22028);
and U22219 (N_22219,N_22080,N_22057);
and U22220 (N_22220,N_22087,N_22107);
nor U22221 (N_22221,N_22033,N_22042);
nor U22222 (N_22222,N_22159,N_22062);
nand U22223 (N_22223,N_22110,N_22070);
and U22224 (N_22224,N_22145,N_22162);
and U22225 (N_22225,N_22167,N_22075);
nor U22226 (N_22226,N_22049,N_22182);
or U22227 (N_22227,N_22029,N_22166);
or U22228 (N_22228,N_22160,N_22193);
and U22229 (N_22229,N_22053,N_22025);
nand U22230 (N_22230,N_22063,N_22018);
nand U22231 (N_22231,N_22184,N_22005);
or U22232 (N_22232,N_22109,N_22058);
or U22233 (N_22233,N_22032,N_22051);
nand U22234 (N_22234,N_22137,N_22048);
and U22235 (N_22235,N_22047,N_22177);
nand U22236 (N_22236,N_22089,N_22041);
nor U22237 (N_22237,N_22146,N_22072);
or U22238 (N_22238,N_22117,N_22108);
nor U22239 (N_22239,N_22006,N_22138);
or U22240 (N_22240,N_22059,N_22044);
nor U22241 (N_22241,N_22016,N_22128);
and U22242 (N_22242,N_22118,N_22010);
or U22243 (N_22243,N_22157,N_22067);
or U22244 (N_22244,N_22185,N_22046);
nand U22245 (N_22245,N_22194,N_22071);
nand U22246 (N_22246,N_22169,N_22119);
and U22247 (N_22247,N_22190,N_22019);
nand U22248 (N_22248,N_22161,N_22174);
and U22249 (N_22249,N_22014,N_22186);
or U22250 (N_22250,N_22171,N_22066);
and U22251 (N_22251,N_22154,N_22143);
nand U22252 (N_22252,N_22175,N_22165);
and U22253 (N_22253,N_22027,N_22034);
nor U22254 (N_22254,N_22054,N_22188);
and U22255 (N_22255,N_22030,N_22164);
or U22256 (N_22256,N_22088,N_22015);
and U22257 (N_22257,N_22081,N_22149);
nand U22258 (N_22258,N_22096,N_22064);
or U22259 (N_22259,N_22084,N_22111);
or U22260 (N_22260,N_22105,N_22150);
nand U22261 (N_22261,N_22077,N_22126);
nor U22262 (N_22262,N_22093,N_22197);
and U22263 (N_22263,N_22133,N_22173);
nand U22264 (N_22264,N_22196,N_22061);
and U22265 (N_22265,N_22180,N_22031);
nor U22266 (N_22266,N_22115,N_22170);
or U22267 (N_22267,N_22116,N_22004);
and U22268 (N_22268,N_22158,N_22132);
and U22269 (N_22269,N_22035,N_22192);
xor U22270 (N_22270,N_22024,N_22112);
or U22271 (N_22271,N_22101,N_22009);
nor U22272 (N_22272,N_22092,N_22136);
nor U22273 (N_22273,N_22130,N_22125);
nand U22274 (N_22274,N_22091,N_22106);
and U22275 (N_22275,N_22095,N_22012);
nor U22276 (N_22276,N_22104,N_22103);
and U22277 (N_22277,N_22189,N_22120);
or U22278 (N_22278,N_22139,N_22187);
nand U22279 (N_22279,N_22055,N_22098);
and U22280 (N_22280,N_22123,N_22122);
and U22281 (N_22281,N_22099,N_22008);
nor U22282 (N_22282,N_22141,N_22001);
and U22283 (N_22283,N_22017,N_22168);
nor U22284 (N_22284,N_22114,N_22038);
nor U22285 (N_22285,N_22131,N_22163);
or U22286 (N_22286,N_22056,N_22183);
nor U22287 (N_22287,N_22147,N_22078);
and U22288 (N_22288,N_22036,N_22144);
nand U22289 (N_22289,N_22090,N_22156);
or U22290 (N_22290,N_22100,N_22050);
nor U22291 (N_22291,N_22094,N_22181);
or U22292 (N_22292,N_22152,N_22026);
nand U22293 (N_22293,N_22069,N_22155);
nor U22294 (N_22294,N_22135,N_22195);
nor U22295 (N_22295,N_22082,N_22011);
and U22296 (N_22296,N_22199,N_22068);
nand U22297 (N_22297,N_22000,N_22127);
and U22298 (N_22298,N_22083,N_22043);
nor U22299 (N_22299,N_22065,N_22142);
or U22300 (N_22300,N_22009,N_22099);
nand U22301 (N_22301,N_22056,N_22076);
nor U22302 (N_22302,N_22074,N_22055);
nor U22303 (N_22303,N_22125,N_22082);
or U22304 (N_22304,N_22185,N_22159);
or U22305 (N_22305,N_22096,N_22068);
or U22306 (N_22306,N_22174,N_22181);
nand U22307 (N_22307,N_22065,N_22108);
nor U22308 (N_22308,N_22117,N_22054);
nand U22309 (N_22309,N_22103,N_22116);
and U22310 (N_22310,N_22177,N_22115);
and U22311 (N_22311,N_22018,N_22163);
nor U22312 (N_22312,N_22071,N_22047);
nor U22313 (N_22313,N_22115,N_22076);
nor U22314 (N_22314,N_22176,N_22198);
or U22315 (N_22315,N_22145,N_22157);
or U22316 (N_22316,N_22161,N_22178);
nand U22317 (N_22317,N_22087,N_22055);
and U22318 (N_22318,N_22015,N_22026);
and U22319 (N_22319,N_22135,N_22044);
or U22320 (N_22320,N_22076,N_22160);
or U22321 (N_22321,N_22057,N_22042);
nor U22322 (N_22322,N_22016,N_22020);
nor U22323 (N_22323,N_22052,N_22115);
nor U22324 (N_22324,N_22157,N_22158);
or U22325 (N_22325,N_22037,N_22136);
and U22326 (N_22326,N_22100,N_22150);
nor U22327 (N_22327,N_22172,N_22067);
nor U22328 (N_22328,N_22026,N_22002);
or U22329 (N_22329,N_22164,N_22119);
and U22330 (N_22330,N_22162,N_22036);
nor U22331 (N_22331,N_22159,N_22130);
or U22332 (N_22332,N_22058,N_22011);
and U22333 (N_22333,N_22065,N_22031);
and U22334 (N_22334,N_22198,N_22130);
nor U22335 (N_22335,N_22122,N_22003);
or U22336 (N_22336,N_22104,N_22021);
and U22337 (N_22337,N_22104,N_22058);
nand U22338 (N_22338,N_22031,N_22014);
nand U22339 (N_22339,N_22006,N_22036);
or U22340 (N_22340,N_22080,N_22064);
or U22341 (N_22341,N_22107,N_22114);
or U22342 (N_22342,N_22071,N_22088);
nand U22343 (N_22343,N_22080,N_22144);
nand U22344 (N_22344,N_22024,N_22162);
nand U22345 (N_22345,N_22179,N_22154);
and U22346 (N_22346,N_22183,N_22165);
or U22347 (N_22347,N_22061,N_22008);
nand U22348 (N_22348,N_22183,N_22198);
nand U22349 (N_22349,N_22077,N_22139);
nand U22350 (N_22350,N_22003,N_22129);
nand U22351 (N_22351,N_22046,N_22118);
xor U22352 (N_22352,N_22078,N_22131);
nor U22353 (N_22353,N_22117,N_22066);
and U22354 (N_22354,N_22151,N_22134);
or U22355 (N_22355,N_22079,N_22100);
nand U22356 (N_22356,N_22083,N_22004);
or U22357 (N_22357,N_22141,N_22126);
nand U22358 (N_22358,N_22104,N_22191);
or U22359 (N_22359,N_22162,N_22159);
nor U22360 (N_22360,N_22096,N_22114);
nand U22361 (N_22361,N_22104,N_22038);
nand U22362 (N_22362,N_22149,N_22063);
nand U22363 (N_22363,N_22023,N_22186);
nor U22364 (N_22364,N_22103,N_22188);
and U22365 (N_22365,N_22068,N_22088);
nand U22366 (N_22366,N_22034,N_22135);
nor U22367 (N_22367,N_22137,N_22113);
or U22368 (N_22368,N_22076,N_22182);
or U22369 (N_22369,N_22138,N_22196);
or U22370 (N_22370,N_22061,N_22128);
and U22371 (N_22371,N_22191,N_22045);
or U22372 (N_22372,N_22160,N_22143);
nor U22373 (N_22373,N_22178,N_22080);
and U22374 (N_22374,N_22113,N_22126);
and U22375 (N_22375,N_22129,N_22049);
and U22376 (N_22376,N_22013,N_22102);
and U22377 (N_22377,N_22144,N_22153);
and U22378 (N_22378,N_22190,N_22125);
and U22379 (N_22379,N_22132,N_22179);
or U22380 (N_22380,N_22086,N_22184);
nand U22381 (N_22381,N_22051,N_22160);
and U22382 (N_22382,N_22078,N_22000);
or U22383 (N_22383,N_22070,N_22105);
and U22384 (N_22384,N_22100,N_22055);
and U22385 (N_22385,N_22116,N_22122);
or U22386 (N_22386,N_22151,N_22176);
and U22387 (N_22387,N_22113,N_22090);
or U22388 (N_22388,N_22024,N_22121);
nand U22389 (N_22389,N_22165,N_22114);
or U22390 (N_22390,N_22006,N_22132);
or U22391 (N_22391,N_22105,N_22031);
or U22392 (N_22392,N_22100,N_22070);
and U22393 (N_22393,N_22100,N_22144);
and U22394 (N_22394,N_22021,N_22135);
nand U22395 (N_22395,N_22114,N_22134);
nor U22396 (N_22396,N_22073,N_22083);
nor U22397 (N_22397,N_22169,N_22064);
nor U22398 (N_22398,N_22181,N_22121);
and U22399 (N_22399,N_22183,N_22078);
or U22400 (N_22400,N_22240,N_22396);
nor U22401 (N_22401,N_22370,N_22316);
and U22402 (N_22402,N_22306,N_22215);
nor U22403 (N_22403,N_22318,N_22393);
nor U22404 (N_22404,N_22303,N_22224);
and U22405 (N_22405,N_22247,N_22276);
and U22406 (N_22406,N_22234,N_22295);
nand U22407 (N_22407,N_22255,N_22283);
nor U22408 (N_22408,N_22333,N_22357);
nor U22409 (N_22409,N_22207,N_22201);
and U22410 (N_22410,N_22289,N_22266);
or U22411 (N_22411,N_22375,N_22397);
nor U22412 (N_22412,N_22273,N_22244);
and U22413 (N_22413,N_22205,N_22389);
nand U22414 (N_22414,N_22299,N_22391);
and U22415 (N_22415,N_22204,N_22225);
or U22416 (N_22416,N_22336,N_22359);
and U22417 (N_22417,N_22304,N_22291);
and U22418 (N_22418,N_22223,N_22288);
and U22419 (N_22419,N_22249,N_22216);
and U22420 (N_22420,N_22380,N_22355);
and U22421 (N_22421,N_22233,N_22279);
nand U22422 (N_22422,N_22226,N_22275);
or U22423 (N_22423,N_22331,N_22392);
or U22424 (N_22424,N_22250,N_22314);
or U22425 (N_22425,N_22285,N_22214);
and U22426 (N_22426,N_22372,N_22200);
nand U22427 (N_22427,N_22310,N_22259);
nor U22428 (N_22428,N_22344,N_22352);
nor U22429 (N_22429,N_22366,N_22222);
or U22430 (N_22430,N_22229,N_22277);
or U22431 (N_22431,N_22383,N_22252);
or U22432 (N_22432,N_22230,N_22329);
nor U22433 (N_22433,N_22217,N_22354);
and U22434 (N_22434,N_22361,N_22311);
or U22435 (N_22435,N_22236,N_22203);
nand U22436 (N_22436,N_22210,N_22343);
or U22437 (N_22437,N_22272,N_22341);
nor U22438 (N_22438,N_22385,N_22309);
nor U22439 (N_22439,N_22258,N_22360);
nor U22440 (N_22440,N_22245,N_22256);
and U22441 (N_22441,N_22339,N_22209);
and U22442 (N_22442,N_22251,N_22376);
or U22443 (N_22443,N_22330,N_22335);
or U22444 (N_22444,N_22294,N_22293);
and U22445 (N_22445,N_22313,N_22325);
nand U22446 (N_22446,N_22282,N_22248);
nand U22447 (N_22447,N_22300,N_22395);
and U22448 (N_22448,N_22351,N_22269);
nand U22449 (N_22449,N_22262,N_22296);
or U22450 (N_22450,N_22362,N_22267);
and U22451 (N_22451,N_22246,N_22323);
nor U22452 (N_22452,N_22378,N_22235);
and U22453 (N_22453,N_22253,N_22328);
nand U22454 (N_22454,N_22238,N_22371);
or U22455 (N_22455,N_22321,N_22346);
or U22456 (N_22456,N_22349,N_22394);
and U22457 (N_22457,N_22347,N_22202);
nor U22458 (N_22458,N_22369,N_22211);
and U22459 (N_22459,N_22334,N_22308);
or U22460 (N_22460,N_22367,N_22358);
nand U22461 (N_22461,N_22337,N_22254);
or U22462 (N_22462,N_22208,N_22356);
nor U22463 (N_22463,N_22232,N_22284);
nor U22464 (N_22464,N_22218,N_22302);
nor U22465 (N_22465,N_22265,N_22219);
nor U22466 (N_22466,N_22292,N_22281);
or U22467 (N_22467,N_22312,N_22220);
or U22468 (N_22468,N_22237,N_22384);
or U22469 (N_22469,N_22264,N_22301);
or U22470 (N_22470,N_22206,N_22363);
and U22471 (N_22471,N_22348,N_22365);
and U22472 (N_22472,N_22298,N_22278);
nor U22473 (N_22473,N_22243,N_22242);
and U22474 (N_22474,N_22315,N_22379);
and U22475 (N_22475,N_22274,N_22374);
nand U22476 (N_22476,N_22350,N_22268);
or U22477 (N_22477,N_22212,N_22317);
or U22478 (N_22478,N_22239,N_22327);
and U22479 (N_22479,N_22307,N_22382);
nand U22480 (N_22480,N_22338,N_22332);
and U22481 (N_22481,N_22320,N_22270);
and U22482 (N_22482,N_22388,N_22373);
or U22483 (N_22483,N_22287,N_22377);
nor U22484 (N_22484,N_22241,N_22290);
and U22485 (N_22485,N_22228,N_22398);
nor U22486 (N_22486,N_22257,N_22368);
nand U22487 (N_22487,N_22286,N_22390);
and U22488 (N_22488,N_22326,N_22324);
or U22489 (N_22489,N_22340,N_22213);
or U22490 (N_22490,N_22271,N_22221);
or U22491 (N_22491,N_22381,N_22319);
nor U22492 (N_22492,N_22297,N_22345);
nor U22493 (N_22493,N_22227,N_22260);
or U22494 (N_22494,N_22280,N_22364);
or U22495 (N_22495,N_22305,N_22263);
nand U22496 (N_22496,N_22386,N_22387);
nor U22497 (N_22497,N_22261,N_22342);
or U22498 (N_22498,N_22231,N_22353);
or U22499 (N_22499,N_22322,N_22399);
nand U22500 (N_22500,N_22301,N_22335);
xnor U22501 (N_22501,N_22295,N_22324);
and U22502 (N_22502,N_22310,N_22360);
nor U22503 (N_22503,N_22226,N_22272);
nand U22504 (N_22504,N_22321,N_22370);
nand U22505 (N_22505,N_22367,N_22256);
or U22506 (N_22506,N_22329,N_22275);
and U22507 (N_22507,N_22269,N_22251);
or U22508 (N_22508,N_22372,N_22252);
or U22509 (N_22509,N_22315,N_22227);
and U22510 (N_22510,N_22245,N_22282);
nor U22511 (N_22511,N_22269,N_22324);
or U22512 (N_22512,N_22334,N_22281);
and U22513 (N_22513,N_22335,N_22298);
nand U22514 (N_22514,N_22297,N_22307);
or U22515 (N_22515,N_22371,N_22367);
or U22516 (N_22516,N_22281,N_22243);
nand U22517 (N_22517,N_22226,N_22289);
nand U22518 (N_22518,N_22231,N_22314);
nor U22519 (N_22519,N_22200,N_22388);
nor U22520 (N_22520,N_22238,N_22200);
xnor U22521 (N_22521,N_22259,N_22334);
and U22522 (N_22522,N_22388,N_22286);
nor U22523 (N_22523,N_22232,N_22396);
or U22524 (N_22524,N_22352,N_22307);
and U22525 (N_22525,N_22222,N_22341);
or U22526 (N_22526,N_22366,N_22392);
nor U22527 (N_22527,N_22296,N_22361);
or U22528 (N_22528,N_22264,N_22237);
or U22529 (N_22529,N_22282,N_22213);
and U22530 (N_22530,N_22273,N_22384);
or U22531 (N_22531,N_22236,N_22246);
nor U22532 (N_22532,N_22294,N_22246);
or U22533 (N_22533,N_22301,N_22362);
or U22534 (N_22534,N_22300,N_22393);
or U22535 (N_22535,N_22281,N_22203);
nand U22536 (N_22536,N_22267,N_22374);
and U22537 (N_22537,N_22311,N_22336);
nand U22538 (N_22538,N_22378,N_22375);
nor U22539 (N_22539,N_22201,N_22253);
nand U22540 (N_22540,N_22227,N_22258);
and U22541 (N_22541,N_22375,N_22368);
or U22542 (N_22542,N_22206,N_22392);
nand U22543 (N_22543,N_22250,N_22332);
or U22544 (N_22544,N_22262,N_22355);
and U22545 (N_22545,N_22283,N_22218);
and U22546 (N_22546,N_22351,N_22391);
and U22547 (N_22547,N_22236,N_22279);
and U22548 (N_22548,N_22211,N_22399);
nor U22549 (N_22549,N_22267,N_22383);
xor U22550 (N_22550,N_22249,N_22220);
and U22551 (N_22551,N_22330,N_22305);
or U22552 (N_22552,N_22313,N_22252);
and U22553 (N_22553,N_22378,N_22239);
and U22554 (N_22554,N_22278,N_22284);
and U22555 (N_22555,N_22274,N_22266);
and U22556 (N_22556,N_22299,N_22280);
nand U22557 (N_22557,N_22296,N_22293);
nor U22558 (N_22558,N_22289,N_22202);
or U22559 (N_22559,N_22281,N_22207);
or U22560 (N_22560,N_22214,N_22243);
or U22561 (N_22561,N_22279,N_22353);
or U22562 (N_22562,N_22354,N_22253);
nor U22563 (N_22563,N_22271,N_22274);
nand U22564 (N_22564,N_22364,N_22346);
or U22565 (N_22565,N_22224,N_22252);
and U22566 (N_22566,N_22216,N_22269);
nor U22567 (N_22567,N_22275,N_22251);
xor U22568 (N_22568,N_22284,N_22215);
nand U22569 (N_22569,N_22286,N_22227);
nor U22570 (N_22570,N_22299,N_22348);
nand U22571 (N_22571,N_22322,N_22353);
nand U22572 (N_22572,N_22387,N_22203);
or U22573 (N_22573,N_22208,N_22207);
and U22574 (N_22574,N_22357,N_22346);
and U22575 (N_22575,N_22281,N_22348);
nand U22576 (N_22576,N_22285,N_22312);
nor U22577 (N_22577,N_22372,N_22338);
and U22578 (N_22578,N_22291,N_22335);
and U22579 (N_22579,N_22349,N_22304);
and U22580 (N_22580,N_22334,N_22263);
and U22581 (N_22581,N_22398,N_22256);
nor U22582 (N_22582,N_22274,N_22330);
and U22583 (N_22583,N_22301,N_22323);
nor U22584 (N_22584,N_22367,N_22303);
and U22585 (N_22585,N_22274,N_22246);
and U22586 (N_22586,N_22276,N_22209);
nand U22587 (N_22587,N_22293,N_22203);
and U22588 (N_22588,N_22200,N_22256);
and U22589 (N_22589,N_22396,N_22351);
nand U22590 (N_22590,N_22325,N_22243);
and U22591 (N_22591,N_22239,N_22330);
and U22592 (N_22592,N_22340,N_22204);
nand U22593 (N_22593,N_22231,N_22207);
and U22594 (N_22594,N_22285,N_22291);
or U22595 (N_22595,N_22337,N_22370);
or U22596 (N_22596,N_22274,N_22270);
nand U22597 (N_22597,N_22217,N_22246);
or U22598 (N_22598,N_22396,N_22200);
xnor U22599 (N_22599,N_22204,N_22384);
nor U22600 (N_22600,N_22470,N_22536);
and U22601 (N_22601,N_22518,N_22462);
nor U22602 (N_22602,N_22446,N_22433);
or U22603 (N_22603,N_22497,N_22574);
nand U22604 (N_22604,N_22508,N_22480);
and U22605 (N_22605,N_22461,N_22570);
and U22606 (N_22606,N_22488,N_22465);
nand U22607 (N_22607,N_22595,N_22554);
nor U22608 (N_22608,N_22439,N_22427);
nand U22609 (N_22609,N_22469,N_22597);
nand U22610 (N_22610,N_22434,N_22413);
nand U22611 (N_22611,N_22441,N_22416);
nand U22612 (N_22612,N_22510,N_22576);
nor U22613 (N_22613,N_22475,N_22507);
or U22614 (N_22614,N_22501,N_22517);
and U22615 (N_22615,N_22449,N_22535);
or U22616 (N_22616,N_22460,N_22579);
and U22617 (N_22617,N_22424,N_22590);
nor U22618 (N_22618,N_22455,N_22513);
nand U22619 (N_22619,N_22509,N_22494);
or U22620 (N_22620,N_22514,N_22437);
nor U22621 (N_22621,N_22563,N_22489);
nand U22622 (N_22622,N_22580,N_22559);
nand U22623 (N_22623,N_22546,N_22528);
nor U22624 (N_22624,N_22426,N_22459);
nand U22625 (N_22625,N_22400,N_22532);
nand U22626 (N_22626,N_22537,N_22567);
or U22627 (N_22627,N_22582,N_22538);
nor U22628 (N_22628,N_22587,N_22432);
and U22629 (N_22629,N_22534,N_22406);
nor U22630 (N_22630,N_22421,N_22473);
or U22631 (N_22631,N_22599,N_22474);
nor U22632 (N_22632,N_22542,N_22479);
nor U22633 (N_22633,N_22577,N_22436);
nand U22634 (N_22634,N_22447,N_22578);
and U22635 (N_22635,N_22451,N_22458);
or U22636 (N_22636,N_22594,N_22504);
nor U22637 (N_22637,N_22521,N_22409);
nand U22638 (N_22638,N_22463,N_22467);
nor U22639 (N_22639,N_22551,N_22429);
nor U22640 (N_22640,N_22540,N_22499);
nand U22641 (N_22641,N_22516,N_22456);
nand U22642 (N_22642,N_22407,N_22565);
or U22643 (N_22643,N_22571,N_22547);
nor U22644 (N_22644,N_22589,N_22404);
nand U22645 (N_22645,N_22530,N_22544);
and U22646 (N_22646,N_22558,N_22556);
and U22647 (N_22647,N_22503,N_22525);
nand U22648 (N_22648,N_22482,N_22506);
nor U22649 (N_22649,N_22529,N_22471);
nand U22650 (N_22650,N_22592,N_22572);
or U22651 (N_22651,N_22428,N_22512);
or U22652 (N_22652,N_22598,N_22402);
nand U22653 (N_22653,N_22453,N_22533);
nor U22654 (N_22654,N_22522,N_22573);
nand U22655 (N_22655,N_22477,N_22410);
nor U22656 (N_22656,N_22562,N_22586);
nand U22657 (N_22657,N_22430,N_22549);
nor U22658 (N_22658,N_22412,N_22591);
and U22659 (N_22659,N_22583,N_22519);
nor U22660 (N_22660,N_22575,N_22481);
or U22661 (N_22661,N_22440,N_22492);
nor U22662 (N_22662,N_22478,N_22444);
or U22663 (N_22663,N_22431,N_22566);
nor U22664 (N_22664,N_22545,N_22466);
nor U22665 (N_22665,N_22448,N_22496);
nand U22666 (N_22666,N_22584,N_22560);
or U22667 (N_22667,N_22472,N_22422);
and U22668 (N_22668,N_22505,N_22568);
nand U22669 (N_22669,N_22581,N_22450);
nor U22670 (N_22670,N_22411,N_22435);
or U22671 (N_22671,N_22561,N_22443);
xnor U22672 (N_22672,N_22550,N_22423);
and U22673 (N_22673,N_22495,N_22442);
and U22674 (N_22674,N_22539,N_22564);
nand U22675 (N_22675,N_22527,N_22419);
or U22676 (N_22676,N_22493,N_22548);
and U22677 (N_22677,N_22523,N_22593);
or U22678 (N_22678,N_22531,N_22543);
and U22679 (N_22679,N_22526,N_22585);
nand U22680 (N_22680,N_22405,N_22438);
or U22681 (N_22681,N_22596,N_22515);
nand U22682 (N_22682,N_22415,N_22511);
nor U22683 (N_22683,N_22425,N_22486);
nand U22684 (N_22684,N_22418,N_22498);
or U22685 (N_22685,N_22420,N_22464);
nor U22686 (N_22686,N_22417,N_22401);
nor U22687 (N_22687,N_22487,N_22457);
nor U22688 (N_22688,N_22468,N_22569);
and U22689 (N_22689,N_22484,N_22476);
nand U22690 (N_22690,N_22541,N_22408);
nor U22691 (N_22691,N_22524,N_22452);
or U22692 (N_22692,N_22520,N_22491);
nor U22693 (N_22693,N_22502,N_22588);
nor U22694 (N_22694,N_22490,N_22557);
nand U22695 (N_22695,N_22414,N_22403);
and U22696 (N_22696,N_22485,N_22483);
and U22697 (N_22697,N_22552,N_22445);
nor U22698 (N_22698,N_22555,N_22553);
nor U22699 (N_22699,N_22454,N_22500);
and U22700 (N_22700,N_22544,N_22426);
and U22701 (N_22701,N_22534,N_22456);
and U22702 (N_22702,N_22544,N_22425);
and U22703 (N_22703,N_22462,N_22546);
and U22704 (N_22704,N_22428,N_22475);
nand U22705 (N_22705,N_22524,N_22446);
nor U22706 (N_22706,N_22593,N_22526);
nor U22707 (N_22707,N_22413,N_22557);
nor U22708 (N_22708,N_22467,N_22519);
nand U22709 (N_22709,N_22423,N_22569);
and U22710 (N_22710,N_22503,N_22476);
nor U22711 (N_22711,N_22537,N_22431);
nor U22712 (N_22712,N_22539,N_22547);
and U22713 (N_22713,N_22509,N_22421);
nand U22714 (N_22714,N_22559,N_22416);
and U22715 (N_22715,N_22556,N_22440);
nand U22716 (N_22716,N_22514,N_22418);
nor U22717 (N_22717,N_22530,N_22421);
nand U22718 (N_22718,N_22432,N_22482);
and U22719 (N_22719,N_22535,N_22481);
or U22720 (N_22720,N_22548,N_22419);
nor U22721 (N_22721,N_22496,N_22579);
or U22722 (N_22722,N_22437,N_22495);
nor U22723 (N_22723,N_22441,N_22508);
or U22724 (N_22724,N_22589,N_22424);
nor U22725 (N_22725,N_22506,N_22559);
and U22726 (N_22726,N_22514,N_22519);
nor U22727 (N_22727,N_22556,N_22500);
or U22728 (N_22728,N_22558,N_22435);
nor U22729 (N_22729,N_22421,N_22454);
nand U22730 (N_22730,N_22414,N_22440);
or U22731 (N_22731,N_22428,N_22511);
nor U22732 (N_22732,N_22412,N_22529);
nor U22733 (N_22733,N_22443,N_22453);
nor U22734 (N_22734,N_22470,N_22524);
and U22735 (N_22735,N_22437,N_22581);
nand U22736 (N_22736,N_22495,N_22447);
nand U22737 (N_22737,N_22493,N_22535);
or U22738 (N_22738,N_22421,N_22450);
nor U22739 (N_22739,N_22557,N_22507);
and U22740 (N_22740,N_22462,N_22585);
nor U22741 (N_22741,N_22560,N_22586);
and U22742 (N_22742,N_22445,N_22567);
or U22743 (N_22743,N_22574,N_22576);
and U22744 (N_22744,N_22477,N_22429);
and U22745 (N_22745,N_22565,N_22572);
and U22746 (N_22746,N_22573,N_22450);
or U22747 (N_22747,N_22437,N_22593);
nand U22748 (N_22748,N_22584,N_22468);
nand U22749 (N_22749,N_22520,N_22404);
and U22750 (N_22750,N_22412,N_22488);
or U22751 (N_22751,N_22416,N_22529);
or U22752 (N_22752,N_22430,N_22503);
or U22753 (N_22753,N_22489,N_22557);
or U22754 (N_22754,N_22491,N_22531);
nor U22755 (N_22755,N_22413,N_22438);
and U22756 (N_22756,N_22567,N_22469);
or U22757 (N_22757,N_22549,N_22525);
nor U22758 (N_22758,N_22545,N_22417);
nand U22759 (N_22759,N_22479,N_22544);
xor U22760 (N_22760,N_22478,N_22429);
or U22761 (N_22761,N_22541,N_22453);
nand U22762 (N_22762,N_22563,N_22456);
and U22763 (N_22763,N_22430,N_22518);
nor U22764 (N_22764,N_22532,N_22519);
nor U22765 (N_22765,N_22595,N_22559);
and U22766 (N_22766,N_22573,N_22402);
or U22767 (N_22767,N_22579,N_22400);
nor U22768 (N_22768,N_22466,N_22467);
and U22769 (N_22769,N_22413,N_22539);
nor U22770 (N_22770,N_22478,N_22449);
and U22771 (N_22771,N_22512,N_22523);
nor U22772 (N_22772,N_22570,N_22548);
and U22773 (N_22773,N_22442,N_22427);
nand U22774 (N_22774,N_22580,N_22410);
nor U22775 (N_22775,N_22458,N_22587);
or U22776 (N_22776,N_22547,N_22412);
nor U22777 (N_22777,N_22488,N_22558);
and U22778 (N_22778,N_22469,N_22481);
nand U22779 (N_22779,N_22437,N_22407);
nand U22780 (N_22780,N_22481,N_22493);
and U22781 (N_22781,N_22497,N_22501);
or U22782 (N_22782,N_22596,N_22508);
nand U22783 (N_22783,N_22421,N_22400);
or U22784 (N_22784,N_22597,N_22491);
nand U22785 (N_22785,N_22560,N_22549);
nand U22786 (N_22786,N_22474,N_22593);
or U22787 (N_22787,N_22529,N_22488);
or U22788 (N_22788,N_22571,N_22467);
nor U22789 (N_22789,N_22440,N_22523);
nand U22790 (N_22790,N_22512,N_22524);
nor U22791 (N_22791,N_22550,N_22463);
nand U22792 (N_22792,N_22542,N_22556);
or U22793 (N_22793,N_22530,N_22401);
nand U22794 (N_22794,N_22475,N_22433);
nand U22795 (N_22795,N_22518,N_22412);
or U22796 (N_22796,N_22460,N_22587);
nand U22797 (N_22797,N_22482,N_22406);
nor U22798 (N_22798,N_22435,N_22512);
or U22799 (N_22799,N_22460,N_22575);
nor U22800 (N_22800,N_22659,N_22768);
nand U22801 (N_22801,N_22775,N_22777);
or U22802 (N_22802,N_22641,N_22694);
and U22803 (N_22803,N_22649,N_22741);
nor U22804 (N_22804,N_22677,N_22791);
nand U22805 (N_22805,N_22733,N_22731);
or U22806 (N_22806,N_22755,N_22767);
or U22807 (N_22807,N_22667,N_22758);
and U22808 (N_22808,N_22732,N_22662);
and U22809 (N_22809,N_22725,N_22717);
nand U22810 (N_22810,N_22653,N_22640);
and U22811 (N_22811,N_22693,N_22799);
nor U22812 (N_22812,N_22751,N_22718);
or U22813 (N_22813,N_22771,N_22645);
nand U22814 (N_22814,N_22619,N_22686);
and U22815 (N_22815,N_22715,N_22626);
or U22816 (N_22816,N_22704,N_22685);
nand U22817 (N_22817,N_22719,N_22726);
and U22818 (N_22818,N_22683,N_22784);
or U22819 (N_22819,N_22708,N_22690);
nor U22820 (N_22820,N_22663,N_22600);
and U22821 (N_22821,N_22696,N_22754);
or U22822 (N_22822,N_22773,N_22648);
or U22823 (N_22823,N_22643,N_22700);
or U22824 (N_22824,N_22607,N_22692);
nor U22825 (N_22825,N_22756,N_22671);
or U22826 (N_22826,N_22706,N_22613);
nor U22827 (N_22827,N_22609,N_22669);
nor U22828 (N_22828,N_22749,N_22769);
nor U22829 (N_22829,N_22727,N_22794);
nand U22830 (N_22830,N_22605,N_22670);
nor U22831 (N_22831,N_22697,N_22778);
nand U22832 (N_22832,N_22631,N_22743);
nor U22833 (N_22833,N_22765,N_22637);
nand U22834 (N_22834,N_22632,N_22709);
xor U22835 (N_22835,N_22698,N_22621);
nor U22836 (N_22836,N_22703,N_22699);
nor U22837 (N_22837,N_22622,N_22646);
nand U22838 (N_22838,N_22797,N_22748);
and U22839 (N_22839,N_22624,N_22740);
and U22840 (N_22840,N_22614,N_22790);
or U22841 (N_22841,N_22716,N_22608);
nor U22842 (N_22842,N_22687,N_22720);
and U22843 (N_22843,N_22774,N_22764);
nand U22844 (N_22844,N_22654,N_22753);
and U22845 (N_22845,N_22695,N_22782);
and U22846 (N_22846,N_22652,N_22616);
nor U22847 (N_22847,N_22636,N_22747);
nand U22848 (N_22848,N_22745,N_22750);
nor U22849 (N_22849,N_22757,N_22639);
and U22850 (N_22850,N_22779,N_22776);
or U22851 (N_22851,N_22658,N_22635);
nand U22852 (N_22852,N_22701,N_22739);
xnor U22853 (N_22853,N_22655,N_22735);
nand U22854 (N_22854,N_22752,N_22647);
nand U22855 (N_22855,N_22656,N_22642);
and U22856 (N_22856,N_22788,N_22644);
nand U22857 (N_22857,N_22787,N_22734);
or U22858 (N_22858,N_22672,N_22761);
nor U22859 (N_22859,N_22618,N_22763);
nand U22860 (N_22860,N_22630,N_22786);
or U22861 (N_22861,N_22759,N_22678);
or U22862 (N_22862,N_22665,N_22660);
nand U22863 (N_22863,N_22675,N_22606);
nand U22864 (N_22864,N_22628,N_22783);
nand U22865 (N_22865,N_22680,N_22657);
and U22866 (N_22866,N_22766,N_22603);
and U22867 (N_22867,N_22664,N_22676);
nor U22868 (N_22868,N_22666,N_22684);
or U22869 (N_22869,N_22798,N_22689);
nor U22870 (N_22870,N_22623,N_22723);
or U22871 (N_22871,N_22729,N_22702);
or U22872 (N_22872,N_22707,N_22673);
and U22873 (N_22873,N_22651,N_22770);
nor U22874 (N_22874,N_22772,N_22789);
nand U22875 (N_22875,N_22712,N_22610);
xnor U22876 (N_22876,N_22730,N_22721);
nand U22877 (N_22877,N_22620,N_22793);
nor U22878 (N_22878,N_22746,N_22611);
nor U22879 (N_22879,N_22681,N_22710);
and U22880 (N_22880,N_22674,N_22629);
nor U22881 (N_22881,N_22682,N_22602);
and U22882 (N_22882,N_22780,N_22615);
nand U22883 (N_22883,N_22744,N_22762);
nor U22884 (N_22884,N_22650,N_22724);
nor U22885 (N_22885,N_22617,N_22691);
and U22886 (N_22886,N_22796,N_22627);
nand U22887 (N_22887,N_22785,N_22737);
and U22888 (N_22888,N_22711,N_22795);
nand U22889 (N_22889,N_22688,N_22661);
and U22890 (N_22890,N_22713,N_22792);
nor U22891 (N_22891,N_22634,N_22604);
and U22892 (N_22892,N_22601,N_22781);
nor U22893 (N_22893,N_22633,N_22722);
nand U22894 (N_22894,N_22612,N_22679);
and U22895 (N_22895,N_22738,N_22736);
nand U22896 (N_22896,N_22668,N_22705);
and U22897 (N_22897,N_22742,N_22714);
nand U22898 (N_22898,N_22760,N_22638);
or U22899 (N_22899,N_22625,N_22728);
and U22900 (N_22900,N_22741,N_22781);
nand U22901 (N_22901,N_22674,N_22692);
xnor U22902 (N_22902,N_22774,N_22665);
or U22903 (N_22903,N_22685,N_22713);
and U22904 (N_22904,N_22667,N_22666);
or U22905 (N_22905,N_22627,N_22711);
and U22906 (N_22906,N_22601,N_22797);
nor U22907 (N_22907,N_22670,N_22743);
or U22908 (N_22908,N_22687,N_22667);
nand U22909 (N_22909,N_22781,N_22792);
and U22910 (N_22910,N_22777,N_22678);
nor U22911 (N_22911,N_22611,N_22640);
nor U22912 (N_22912,N_22716,N_22613);
and U22913 (N_22913,N_22789,N_22667);
nand U22914 (N_22914,N_22622,N_22707);
or U22915 (N_22915,N_22603,N_22701);
or U22916 (N_22916,N_22709,N_22641);
and U22917 (N_22917,N_22735,N_22727);
nor U22918 (N_22918,N_22630,N_22713);
nand U22919 (N_22919,N_22694,N_22773);
nor U22920 (N_22920,N_22712,N_22713);
or U22921 (N_22921,N_22620,N_22689);
nand U22922 (N_22922,N_22692,N_22787);
nand U22923 (N_22923,N_22667,N_22717);
and U22924 (N_22924,N_22786,N_22640);
and U22925 (N_22925,N_22766,N_22604);
or U22926 (N_22926,N_22788,N_22638);
nand U22927 (N_22927,N_22712,N_22622);
nand U22928 (N_22928,N_22680,N_22722);
nand U22929 (N_22929,N_22751,N_22628);
or U22930 (N_22930,N_22728,N_22635);
nor U22931 (N_22931,N_22732,N_22600);
nor U22932 (N_22932,N_22710,N_22650);
nor U22933 (N_22933,N_22664,N_22723);
nor U22934 (N_22934,N_22730,N_22631);
and U22935 (N_22935,N_22680,N_22703);
nor U22936 (N_22936,N_22767,N_22665);
or U22937 (N_22937,N_22748,N_22624);
nor U22938 (N_22938,N_22787,N_22702);
nor U22939 (N_22939,N_22687,N_22615);
or U22940 (N_22940,N_22780,N_22755);
nor U22941 (N_22941,N_22693,N_22707);
nor U22942 (N_22942,N_22739,N_22755);
or U22943 (N_22943,N_22657,N_22764);
or U22944 (N_22944,N_22705,N_22618);
and U22945 (N_22945,N_22711,N_22645);
nor U22946 (N_22946,N_22725,N_22738);
and U22947 (N_22947,N_22713,N_22638);
nor U22948 (N_22948,N_22728,N_22641);
and U22949 (N_22949,N_22673,N_22655);
or U22950 (N_22950,N_22750,N_22709);
or U22951 (N_22951,N_22657,N_22634);
nand U22952 (N_22952,N_22617,N_22785);
or U22953 (N_22953,N_22638,N_22671);
nor U22954 (N_22954,N_22710,N_22638);
nand U22955 (N_22955,N_22717,N_22722);
or U22956 (N_22956,N_22696,N_22688);
and U22957 (N_22957,N_22784,N_22637);
or U22958 (N_22958,N_22674,N_22630);
and U22959 (N_22959,N_22748,N_22689);
nand U22960 (N_22960,N_22759,N_22795);
nand U22961 (N_22961,N_22715,N_22677);
nor U22962 (N_22962,N_22676,N_22743);
and U22963 (N_22963,N_22790,N_22688);
nor U22964 (N_22964,N_22756,N_22796);
nor U22965 (N_22965,N_22607,N_22725);
and U22966 (N_22966,N_22703,N_22650);
or U22967 (N_22967,N_22687,N_22766);
nand U22968 (N_22968,N_22755,N_22783);
nor U22969 (N_22969,N_22672,N_22633);
nand U22970 (N_22970,N_22660,N_22792);
nand U22971 (N_22971,N_22772,N_22616);
and U22972 (N_22972,N_22623,N_22667);
or U22973 (N_22973,N_22732,N_22697);
nor U22974 (N_22974,N_22744,N_22761);
nand U22975 (N_22975,N_22657,N_22602);
nand U22976 (N_22976,N_22783,N_22753);
nor U22977 (N_22977,N_22699,N_22655);
nor U22978 (N_22978,N_22671,N_22747);
nand U22979 (N_22979,N_22667,N_22781);
and U22980 (N_22980,N_22714,N_22704);
or U22981 (N_22981,N_22640,N_22776);
and U22982 (N_22982,N_22786,N_22765);
or U22983 (N_22983,N_22778,N_22744);
or U22984 (N_22984,N_22658,N_22682);
and U22985 (N_22985,N_22668,N_22774);
and U22986 (N_22986,N_22637,N_22698);
nand U22987 (N_22987,N_22662,N_22648);
and U22988 (N_22988,N_22602,N_22695);
nand U22989 (N_22989,N_22798,N_22618);
or U22990 (N_22990,N_22658,N_22637);
nand U22991 (N_22991,N_22713,N_22795);
and U22992 (N_22992,N_22664,N_22604);
or U22993 (N_22993,N_22722,N_22603);
nand U22994 (N_22994,N_22755,N_22605);
nor U22995 (N_22995,N_22695,N_22631);
nand U22996 (N_22996,N_22678,N_22714);
nand U22997 (N_22997,N_22663,N_22704);
or U22998 (N_22998,N_22756,N_22769);
nor U22999 (N_22999,N_22635,N_22752);
and U23000 (N_23000,N_22996,N_22842);
or U23001 (N_23001,N_22954,N_22866);
and U23002 (N_23002,N_22906,N_22821);
nand U23003 (N_23003,N_22802,N_22991);
and U23004 (N_23004,N_22835,N_22897);
nor U23005 (N_23005,N_22965,N_22914);
nand U23006 (N_23006,N_22930,N_22800);
nand U23007 (N_23007,N_22831,N_22856);
or U23008 (N_23008,N_22823,N_22890);
or U23009 (N_23009,N_22977,N_22907);
nor U23010 (N_23010,N_22913,N_22833);
nor U23011 (N_23011,N_22865,N_22942);
or U23012 (N_23012,N_22959,N_22994);
nor U23013 (N_23013,N_22916,N_22868);
or U23014 (N_23014,N_22889,N_22829);
and U23015 (N_23015,N_22982,N_22815);
nor U23016 (N_23016,N_22891,N_22872);
or U23017 (N_23017,N_22813,N_22984);
and U23018 (N_23018,N_22816,N_22944);
and U23019 (N_23019,N_22808,N_22989);
or U23020 (N_23020,N_22883,N_22923);
and U23021 (N_23021,N_22938,N_22966);
nor U23022 (N_23022,N_22971,N_22998);
nor U23023 (N_23023,N_22893,N_22843);
nand U23024 (N_23024,N_22812,N_22926);
nor U23025 (N_23025,N_22892,N_22929);
or U23026 (N_23026,N_22811,N_22937);
and U23027 (N_23027,N_22894,N_22976);
nand U23028 (N_23028,N_22839,N_22841);
or U23029 (N_23029,N_22853,N_22973);
and U23030 (N_23030,N_22832,N_22881);
nand U23031 (N_23031,N_22805,N_22900);
and U23032 (N_23032,N_22836,N_22895);
or U23033 (N_23033,N_22884,N_22845);
or U23034 (N_23034,N_22828,N_22952);
nand U23035 (N_23035,N_22864,N_22902);
nor U23036 (N_23036,N_22887,N_22896);
and U23037 (N_23037,N_22936,N_22904);
nor U23038 (N_23038,N_22974,N_22869);
nor U23039 (N_23039,N_22978,N_22983);
nand U23040 (N_23040,N_22874,N_22879);
nor U23041 (N_23041,N_22909,N_22880);
or U23042 (N_23042,N_22803,N_22859);
and U23043 (N_23043,N_22981,N_22995);
or U23044 (N_23044,N_22817,N_22899);
nor U23045 (N_23045,N_22992,N_22920);
nor U23046 (N_23046,N_22871,N_22844);
xor U23047 (N_23047,N_22878,N_22943);
and U23048 (N_23048,N_22986,N_22955);
nor U23049 (N_23049,N_22935,N_22933);
nand U23050 (N_23050,N_22888,N_22898);
nand U23051 (N_23051,N_22905,N_22963);
or U23052 (N_23052,N_22969,N_22931);
xor U23053 (N_23053,N_22840,N_22928);
or U23054 (N_23054,N_22858,N_22985);
or U23055 (N_23055,N_22950,N_22988);
nand U23056 (N_23056,N_22870,N_22960);
nor U23057 (N_23057,N_22990,N_22948);
nand U23058 (N_23058,N_22818,N_22951);
or U23059 (N_23059,N_22956,N_22970);
or U23060 (N_23060,N_22968,N_22910);
or U23061 (N_23061,N_22860,N_22857);
and U23062 (N_23062,N_22847,N_22886);
or U23063 (N_23063,N_22806,N_22908);
and U23064 (N_23064,N_22827,N_22953);
nor U23065 (N_23065,N_22993,N_22851);
nand U23066 (N_23066,N_22958,N_22918);
nor U23067 (N_23067,N_22838,N_22924);
or U23068 (N_23068,N_22901,N_22975);
nor U23069 (N_23069,N_22807,N_22987);
or U23070 (N_23070,N_22939,N_22822);
and U23071 (N_23071,N_22876,N_22825);
and U23072 (N_23072,N_22873,N_22932);
nand U23073 (N_23073,N_22862,N_22867);
nand U23074 (N_23074,N_22945,N_22979);
nor U23075 (N_23075,N_22852,N_22967);
nand U23076 (N_23076,N_22941,N_22972);
or U23077 (N_23077,N_22940,N_22980);
or U23078 (N_23078,N_22849,N_22885);
nand U23079 (N_23079,N_22921,N_22826);
nor U23080 (N_23080,N_22911,N_22877);
nand U23081 (N_23081,N_22882,N_22934);
or U23082 (N_23082,N_22925,N_22947);
nor U23083 (N_23083,N_22855,N_22915);
nor U23084 (N_23084,N_22949,N_22919);
nand U23085 (N_23085,N_22854,N_22861);
and U23086 (N_23086,N_22810,N_22804);
xor U23087 (N_23087,N_22903,N_22964);
and U23088 (N_23088,N_22830,N_22824);
and U23089 (N_23089,N_22809,N_22837);
or U23090 (N_23090,N_22819,N_22946);
or U23091 (N_23091,N_22846,N_22997);
nand U23092 (N_23092,N_22850,N_22875);
nor U23093 (N_23093,N_22927,N_22957);
or U23094 (N_23094,N_22917,N_22999);
nand U23095 (N_23095,N_22820,N_22814);
and U23096 (N_23096,N_22922,N_22848);
nor U23097 (N_23097,N_22834,N_22962);
and U23098 (N_23098,N_22912,N_22961);
and U23099 (N_23099,N_22863,N_22801);
and U23100 (N_23100,N_22966,N_22973);
nor U23101 (N_23101,N_22863,N_22885);
nand U23102 (N_23102,N_22882,N_22812);
and U23103 (N_23103,N_22982,N_22883);
nor U23104 (N_23104,N_22809,N_22980);
nor U23105 (N_23105,N_22934,N_22975);
nor U23106 (N_23106,N_22863,N_22838);
and U23107 (N_23107,N_22949,N_22851);
nor U23108 (N_23108,N_22846,N_22813);
or U23109 (N_23109,N_22938,N_22826);
and U23110 (N_23110,N_22965,N_22821);
and U23111 (N_23111,N_22940,N_22917);
xor U23112 (N_23112,N_22888,N_22802);
and U23113 (N_23113,N_22947,N_22932);
or U23114 (N_23114,N_22871,N_22966);
nand U23115 (N_23115,N_22904,N_22856);
and U23116 (N_23116,N_22963,N_22949);
nand U23117 (N_23117,N_22940,N_22962);
nor U23118 (N_23118,N_22946,N_22889);
nand U23119 (N_23119,N_22830,N_22892);
nor U23120 (N_23120,N_22856,N_22923);
and U23121 (N_23121,N_22832,N_22943);
and U23122 (N_23122,N_22915,N_22952);
and U23123 (N_23123,N_22867,N_22988);
nand U23124 (N_23124,N_22816,N_22930);
or U23125 (N_23125,N_22851,N_22905);
or U23126 (N_23126,N_22952,N_22872);
nor U23127 (N_23127,N_22921,N_22814);
and U23128 (N_23128,N_22914,N_22970);
nand U23129 (N_23129,N_22977,N_22953);
nor U23130 (N_23130,N_22936,N_22906);
and U23131 (N_23131,N_22958,N_22942);
nor U23132 (N_23132,N_22852,N_22823);
nand U23133 (N_23133,N_22824,N_22986);
nor U23134 (N_23134,N_22891,N_22953);
nand U23135 (N_23135,N_22984,N_22906);
and U23136 (N_23136,N_22978,N_22902);
nand U23137 (N_23137,N_22969,N_22983);
or U23138 (N_23138,N_22969,N_22978);
and U23139 (N_23139,N_22840,N_22895);
nand U23140 (N_23140,N_22968,N_22983);
or U23141 (N_23141,N_22800,N_22990);
and U23142 (N_23142,N_22810,N_22986);
nor U23143 (N_23143,N_22806,N_22967);
and U23144 (N_23144,N_22985,N_22805);
and U23145 (N_23145,N_22962,N_22983);
or U23146 (N_23146,N_22866,N_22850);
and U23147 (N_23147,N_22874,N_22803);
nand U23148 (N_23148,N_22953,N_22982);
or U23149 (N_23149,N_22843,N_22847);
and U23150 (N_23150,N_22908,N_22877);
nor U23151 (N_23151,N_22881,N_22835);
nand U23152 (N_23152,N_22862,N_22958);
nand U23153 (N_23153,N_22804,N_22915);
nand U23154 (N_23154,N_22879,N_22870);
nand U23155 (N_23155,N_22911,N_22904);
or U23156 (N_23156,N_22858,N_22884);
and U23157 (N_23157,N_22954,N_22935);
or U23158 (N_23158,N_22964,N_22959);
nor U23159 (N_23159,N_22981,N_22930);
or U23160 (N_23160,N_22837,N_22993);
nor U23161 (N_23161,N_22828,N_22852);
and U23162 (N_23162,N_22909,N_22992);
or U23163 (N_23163,N_22996,N_22872);
nand U23164 (N_23164,N_22990,N_22844);
and U23165 (N_23165,N_22838,N_22902);
nor U23166 (N_23166,N_22964,N_22869);
or U23167 (N_23167,N_22922,N_22940);
or U23168 (N_23168,N_22810,N_22985);
or U23169 (N_23169,N_22840,N_22957);
or U23170 (N_23170,N_22983,N_22887);
nor U23171 (N_23171,N_22841,N_22978);
nand U23172 (N_23172,N_22812,N_22841);
and U23173 (N_23173,N_22968,N_22838);
nand U23174 (N_23174,N_22928,N_22944);
or U23175 (N_23175,N_22830,N_22872);
nand U23176 (N_23176,N_22953,N_22951);
nor U23177 (N_23177,N_22866,N_22821);
and U23178 (N_23178,N_22974,N_22922);
and U23179 (N_23179,N_22841,N_22930);
nand U23180 (N_23180,N_22892,N_22822);
and U23181 (N_23181,N_22823,N_22966);
nand U23182 (N_23182,N_22843,N_22896);
nor U23183 (N_23183,N_22811,N_22903);
nand U23184 (N_23184,N_22875,N_22989);
or U23185 (N_23185,N_22884,N_22829);
and U23186 (N_23186,N_22828,N_22862);
or U23187 (N_23187,N_22854,N_22837);
or U23188 (N_23188,N_22800,N_22915);
nor U23189 (N_23189,N_22938,N_22941);
nor U23190 (N_23190,N_22808,N_22974);
and U23191 (N_23191,N_22830,N_22874);
nand U23192 (N_23192,N_22993,N_22843);
and U23193 (N_23193,N_22867,N_22856);
nand U23194 (N_23194,N_22934,N_22814);
or U23195 (N_23195,N_22868,N_22815);
and U23196 (N_23196,N_22905,N_22832);
nor U23197 (N_23197,N_22876,N_22944);
nand U23198 (N_23198,N_22847,N_22863);
nand U23199 (N_23199,N_22984,N_22874);
or U23200 (N_23200,N_23183,N_23142);
or U23201 (N_23201,N_23044,N_23076);
and U23202 (N_23202,N_23192,N_23109);
nor U23203 (N_23203,N_23057,N_23111);
nand U23204 (N_23204,N_23022,N_23098);
or U23205 (N_23205,N_23036,N_23184);
nand U23206 (N_23206,N_23029,N_23107);
nand U23207 (N_23207,N_23150,N_23053);
nand U23208 (N_23208,N_23063,N_23071);
nand U23209 (N_23209,N_23108,N_23198);
nor U23210 (N_23210,N_23123,N_23035);
nand U23211 (N_23211,N_23138,N_23081);
and U23212 (N_23212,N_23084,N_23015);
nor U23213 (N_23213,N_23086,N_23020);
nor U23214 (N_23214,N_23180,N_23065);
nor U23215 (N_23215,N_23026,N_23025);
nor U23216 (N_23216,N_23147,N_23012);
and U23217 (N_23217,N_23125,N_23181);
nand U23218 (N_23218,N_23083,N_23165);
or U23219 (N_23219,N_23007,N_23050);
nor U23220 (N_23220,N_23006,N_23103);
nand U23221 (N_23221,N_23173,N_23024);
or U23222 (N_23222,N_23092,N_23042);
nand U23223 (N_23223,N_23095,N_23068);
and U23224 (N_23224,N_23161,N_23117);
nand U23225 (N_23225,N_23159,N_23049);
nand U23226 (N_23226,N_23119,N_23152);
nand U23227 (N_23227,N_23001,N_23014);
or U23228 (N_23228,N_23003,N_23045);
nor U23229 (N_23229,N_23191,N_23043);
nor U23230 (N_23230,N_23114,N_23187);
nand U23231 (N_23231,N_23130,N_23164);
nor U23232 (N_23232,N_23115,N_23112);
nand U23233 (N_23233,N_23113,N_23101);
and U23234 (N_23234,N_23193,N_23118);
and U23235 (N_23235,N_23028,N_23177);
or U23236 (N_23236,N_23163,N_23188);
and U23237 (N_23237,N_23079,N_23032);
or U23238 (N_23238,N_23122,N_23061);
or U23239 (N_23239,N_23008,N_23174);
and U23240 (N_23240,N_23039,N_23033);
or U23241 (N_23241,N_23156,N_23054);
or U23242 (N_23242,N_23088,N_23145);
nor U23243 (N_23243,N_23167,N_23153);
or U23244 (N_23244,N_23186,N_23091);
or U23245 (N_23245,N_23023,N_23128);
or U23246 (N_23246,N_23131,N_23062);
or U23247 (N_23247,N_23148,N_23066);
and U23248 (N_23248,N_23051,N_23157);
nor U23249 (N_23249,N_23176,N_23059);
and U23250 (N_23250,N_23077,N_23089);
nand U23251 (N_23251,N_23064,N_23124);
nor U23252 (N_23252,N_23005,N_23196);
and U23253 (N_23253,N_23046,N_23052);
nor U23254 (N_23254,N_23170,N_23047);
and U23255 (N_23255,N_23137,N_23013);
or U23256 (N_23256,N_23027,N_23171);
and U23257 (N_23257,N_23011,N_23040);
or U23258 (N_23258,N_23141,N_23190);
or U23259 (N_23259,N_23060,N_23197);
nor U23260 (N_23260,N_23078,N_23155);
and U23261 (N_23261,N_23075,N_23034);
and U23262 (N_23262,N_23019,N_23082);
and U23263 (N_23263,N_23185,N_23126);
and U23264 (N_23264,N_23085,N_23055);
and U23265 (N_23265,N_23151,N_23182);
and U23266 (N_23266,N_23168,N_23143);
nor U23267 (N_23267,N_23132,N_23017);
or U23268 (N_23268,N_23194,N_23090);
nor U23269 (N_23269,N_23121,N_23016);
or U23270 (N_23270,N_23144,N_23067);
or U23271 (N_23271,N_23110,N_23136);
or U23272 (N_23272,N_23056,N_23133);
or U23273 (N_23273,N_23175,N_23139);
nor U23274 (N_23274,N_23093,N_23178);
nand U23275 (N_23275,N_23002,N_23069);
and U23276 (N_23276,N_23097,N_23189);
or U23277 (N_23277,N_23102,N_23074);
and U23278 (N_23278,N_23096,N_23094);
or U23279 (N_23279,N_23169,N_23104);
and U23280 (N_23280,N_23135,N_23146);
xnor U23281 (N_23281,N_23058,N_23162);
or U23282 (N_23282,N_23195,N_23166);
and U23283 (N_23283,N_23172,N_23041);
and U23284 (N_23284,N_23149,N_23099);
and U23285 (N_23285,N_23105,N_23199);
nand U23286 (N_23286,N_23127,N_23037);
and U23287 (N_23287,N_23038,N_23158);
nor U23288 (N_23288,N_23048,N_23000);
nor U23289 (N_23289,N_23120,N_23134);
nand U23290 (N_23290,N_23087,N_23004);
and U23291 (N_23291,N_23129,N_23140);
and U23292 (N_23292,N_23010,N_23031);
and U23293 (N_23293,N_23073,N_23018);
nor U23294 (N_23294,N_23030,N_23154);
and U23295 (N_23295,N_23100,N_23179);
and U23296 (N_23296,N_23116,N_23021);
or U23297 (N_23297,N_23080,N_23070);
nor U23298 (N_23298,N_23106,N_23009);
or U23299 (N_23299,N_23160,N_23072);
nor U23300 (N_23300,N_23121,N_23029);
nor U23301 (N_23301,N_23152,N_23040);
and U23302 (N_23302,N_23143,N_23015);
nand U23303 (N_23303,N_23199,N_23092);
or U23304 (N_23304,N_23017,N_23000);
nand U23305 (N_23305,N_23184,N_23067);
nor U23306 (N_23306,N_23019,N_23142);
or U23307 (N_23307,N_23070,N_23104);
and U23308 (N_23308,N_23089,N_23040);
or U23309 (N_23309,N_23076,N_23176);
and U23310 (N_23310,N_23188,N_23020);
nor U23311 (N_23311,N_23187,N_23098);
nand U23312 (N_23312,N_23168,N_23185);
nand U23313 (N_23313,N_23022,N_23175);
nand U23314 (N_23314,N_23057,N_23070);
nand U23315 (N_23315,N_23180,N_23077);
and U23316 (N_23316,N_23153,N_23125);
and U23317 (N_23317,N_23092,N_23063);
or U23318 (N_23318,N_23090,N_23165);
nand U23319 (N_23319,N_23072,N_23186);
nand U23320 (N_23320,N_23026,N_23022);
or U23321 (N_23321,N_23172,N_23064);
nor U23322 (N_23322,N_23123,N_23073);
or U23323 (N_23323,N_23169,N_23067);
nor U23324 (N_23324,N_23116,N_23083);
and U23325 (N_23325,N_23070,N_23197);
and U23326 (N_23326,N_23070,N_23189);
nor U23327 (N_23327,N_23050,N_23145);
nor U23328 (N_23328,N_23116,N_23058);
or U23329 (N_23329,N_23001,N_23133);
nor U23330 (N_23330,N_23161,N_23135);
nand U23331 (N_23331,N_23136,N_23162);
nor U23332 (N_23332,N_23189,N_23065);
nand U23333 (N_23333,N_23119,N_23125);
nor U23334 (N_23334,N_23080,N_23045);
nor U23335 (N_23335,N_23020,N_23168);
nand U23336 (N_23336,N_23154,N_23082);
nand U23337 (N_23337,N_23156,N_23191);
and U23338 (N_23338,N_23183,N_23001);
or U23339 (N_23339,N_23039,N_23144);
nor U23340 (N_23340,N_23152,N_23091);
xnor U23341 (N_23341,N_23156,N_23133);
and U23342 (N_23342,N_23187,N_23105);
nor U23343 (N_23343,N_23007,N_23169);
nor U23344 (N_23344,N_23003,N_23012);
and U23345 (N_23345,N_23109,N_23047);
or U23346 (N_23346,N_23071,N_23033);
and U23347 (N_23347,N_23134,N_23021);
nand U23348 (N_23348,N_23085,N_23168);
or U23349 (N_23349,N_23127,N_23187);
or U23350 (N_23350,N_23018,N_23022);
or U23351 (N_23351,N_23162,N_23099);
or U23352 (N_23352,N_23024,N_23181);
or U23353 (N_23353,N_23174,N_23048);
and U23354 (N_23354,N_23164,N_23192);
nor U23355 (N_23355,N_23139,N_23034);
and U23356 (N_23356,N_23147,N_23190);
nor U23357 (N_23357,N_23129,N_23040);
or U23358 (N_23358,N_23122,N_23187);
or U23359 (N_23359,N_23120,N_23059);
or U23360 (N_23360,N_23154,N_23051);
or U23361 (N_23361,N_23117,N_23088);
nor U23362 (N_23362,N_23107,N_23156);
and U23363 (N_23363,N_23096,N_23115);
or U23364 (N_23364,N_23003,N_23178);
or U23365 (N_23365,N_23172,N_23076);
nand U23366 (N_23366,N_23172,N_23059);
nand U23367 (N_23367,N_23169,N_23192);
nor U23368 (N_23368,N_23071,N_23126);
nor U23369 (N_23369,N_23180,N_23053);
nor U23370 (N_23370,N_23190,N_23041);
nor U23371 (N_23371,N_23181,N_23166);
nand U23372 (N_23372,N_23132,N_23182);
nor U23373 (N_23373,N_23163,N_23152);
or U23374 (N_23374,N_23081,N_23102);
nor U23375 (N_23375,N_23013,N_23021);
nand U23376 (N_23376,N_23112,N_23135);
or U23377 (N_23377,N_23038,N_23106);
or U23378 (N_23378,N_23119,N_23098);
or U23379 (N_23379,N_23190,N_23165);
or U23380 (N_23380,N_23147,N_23131);
or U23381 (N_23381,N_23113,N_23109);
nor U23382 (N_23382,N_23107,N_23198);
nand U23383 (N_23383,N_23018,N_23087);
nand U23384 (N_23384,N_23173,N_23101);
or U23385 (N_23385,N_23061,N_23072);
nand U23386 (N_23386,N_23087,N_23073);
or U23387 (N_23387,N_23163,N_23012);
xnor U23388 (N_23388,N_23107,N_23149);
nor U23389 (N_23389,N_23033,N_23024);
nand U23390 (N_23390,N_23016,N_23124);
nor U23391 (N_23391,N_23103,N_23099);
or U23392 (N_23392,N_23003,N_23066);
or U23393 (N_23393,N_23092,N_23077);
nor U23394 (N_23394,N_23141,N_23033);
xor U23395 (N_23395,N_23011,N_23069);
or U23396 (N_23396,N_23139,N_23149);
or U23397 (N_23397,N_23192,N_23075);
nand U23398 (N_23398,N_23185,N_23009);
nor U23399 (N_23399,N_23179,N_23170);
and U23400 (N_23400,N_23256,N_23388);
nor U23401 (N_23401,N_23208,N_23313);
nor U23402 (N_23402,N_23340,N_23297);
or U23403 (N_23403,N_23322,N_23241);
and U23404 (N_23404,N_23350,N_23369);
or U23405 (N_23405,N_23367,N_23220);
or U23406 (N_23406,N_23396,N_23378);
nand U23407 (N_23407,N_23376,N_23343);
nor U23408 (N_23408,N_23300,N_23301);
nand U23409 (N_23409,N_23392,N_23289);
nor U23410 (N_23410,N_23279,N_23280);
or U23411 (N_23411,N_23287,N_23206);
nor U23412 (N_23412,N_23371,N_23203);
and U23413 (N_23413,N_23382,N_23219);
nor U23414 (N_23414,N_23293,N_23318);
and U23415 (N_23415,N_23271,N_23336);
nand U23416 (N_23416,N_23387,N_23227);
and U23417 (N_23417,N_23363,N_23215);
and U23418 (N_23418,N_23218,N_23224);
xnor U23419 (N_23419,N_23207,N_23211);
nor U23420 (N_23420,N_23267,N_23238);
nand U23421 (N_23421,N_23335,N_23290);
nor U23422 (N_23422,N_23282,N_23303);
and U23423 (N_23423,N_23223,N_23352);
nor U23424 (N_23424,N_23307,N_23283);
or U23425 (N_23425,N_23345,N_23353);
or U23426 (N_23426,N_23366,N_23295);
or U23427 (N_23427,N_23284,N_23298);
or U23428 (N_23428,N_23358,N_23397);
or U23429 (N_23429,N_23234,N_23212);
nor U23430 (N_23430,N_23320,N_23391);
or U23431 (N_23431,N_23221,N_23253);
or U23432 (N_23432,N_23329,N_23385);
nand U23433 (N_23433,N_23276,N_23317);
nand U23434 (N_23434,N_23373,N_23246);
or U23435 (N_23435,N_23309,N_23304);
or U23436 (N_23436,N_23327,N_23200);
and U23437 (N_23437,N_23326,N_23359);
nor U23438 (N_23438,N_23312,N_23395);
nand U23439 (N_23439,N_23277,N_23296);
or U23440 (N_23440,N_23244,N_23245);
xor U23441 (N_23441,N_23201,N_23252);
nor U23442 (N_23442,N_23229,N_23249);
or U23443 (N_23443,N_23226,N_23377);
and U23444 (N_23444,N_23344,N_23266);
or U23445 (N_23445,N_23254,N_23275);
nor U23446 (N_23446,N_23324,N_23250);
and U23447 (N_23447,N_23214,N_23262);
nand U23448 (N_23448,N_23231,N_23374);
nor U23449 (N_23449,N_23240,N_23398);
xnor U23450 (N_23450,N_23386,N_23264);
and U23451 (N_23451,N_23325,N_23232);
or U23452 (N_23452,N_23269,N_23235);
and U23453 (N_23453,N_23354,N_23311);
and U23454 (N_23454,N_23286,N_23360);
nor U23455 (N_23455,N_23233,N_23355);
and U23456 (N_23456,N_23251,N_23339);
nand U23457 (N_23457,N_23202,N_23236);
or U23458 (N_23458,N_23308,N_23299);
or U23459 (N_23459,N_23257,N_23292);
nor U23460 (N_23460,N_23230,N_23323);
or U23461 (N_23461,N_23394,N_23368);
nand U23462 (N_23462,N_23259,N_23332);
nand U23463 (N_23463,N_23383,N_23362);
nand U23464 (N_23464,N_23268,N_23380);
and U23465 (N_23465,N_23260,N_23361);
nand U23466 (N_23466,N_23204,N_23316);
nand U23467 (N_23467,N_23210,N_23381);
and U23468 (N_23468,N_23228,N_23349);
nor U23469 (N_23469,N_23393,N_23225);
nor U23470 (N_23470,N_23278,N_23364);
or U23471 (N_23471,N_23205,N_23239);
nand U23472 (N_23472,N_23285,N_23222);
or U23473 (N_23473,N_23237,N_23384);
nor U23474 (N_23474,N_23263,N_23370);
or U23475 (N_23475,N_23247,N_23291);
nand U23476 (N_23476,N_23288,N_23294);
and U23477 (N_23477,N_23372,N_23310);
nor U23478 (N_23478,N_23351,N_23338);
nand U23479 (N_23479,N_23399,N_23217);
and U23480 (N_23480,N_23389,N_23333);
nand U23481 (N_23481,N_23213,N_23346);
nand U23482 (N_23482,N_23216,N_23342);
or U23483 (N_23483,N_23328,N_23341);
and U23484 (N_23484,N_23261,N_23305);
nand U23485 (N_23485,N_23270,N_23302);
nor U23486 (N_23486,N_23356,N_23321);
or U23487 (N_23487,N_23242,N_23390);
nor U23488 (N_23488,N_23265,N_23274);
or U23489 (N_23489,N_23375,N_23379);
and U23490 (N_23490,N_23306,N_23258);
or U23491 (N_23491,N_23337,N_23248);
nor U23492 (N_23492,N_23348,N_23272);
or U23493 (N_23493,N_23334,N_23243);
and U23494 (N_23494,N_23331,N_23357);
and U23495 (N_23495,N_23281,N_23255);
nand U23496 (N_23496,N_23330,N_23273);
and U23497 (N_23497,N_23209,N_23319);
and U23498 (N_23498,N_23365,N_23347);
nor U23499 (N_23499,N_23315,N_23314);
and U23500 (N_23500,N_23253,N_23328);
nor U23501 (N_23501,N_23342,N_23237);
nand U23502 (N_23502,N_23285,N_23267);
or U23503 (N_23503,N_23284,N_23257);
and U23504 (N_23504,N_23354,N_23292);
nand U23505 (N_23505,N_23244,N_23282);
nor U23506 (N_23506,N_23252,N_23356);
or U23507 (N_23507,N_23225,N_23375);
and U23508 (N_23508,N_23316,N_23315);
xor U23509 (N_23509,N_23309,N_23276);
or U23510 (N_23510,N_23240,N_23226);
or U23511 (N_23511,N_23311,N_23388);
and U23512 (N_23512,N_23264,N_23367);
or U23513 (N_23513,N_23398,N_23209);
or U23514 (N_23514,N_23212,N_23201);
nand U23515 (N_23515,N_23230,N_23370);
nand U23516 (N_23516,N_23237,N_23216);
nor U23517 (N_23517,N_23388,N_23355);
nand U23518 (N_23518,N_23295,N_23253);
or U23519 (N_23519,N_23388,N_23354);
nor U23520 (N_23520,N_23215,N_23213);
nand U23521 (N_23521,N_23231,N_23279);
nand U23522 (N_23522,N_23247,N_23374);
or U23523 (N_23523,N_23215,N_23248);
nor U23524 (N_23524,N_23237,N_23393);
or U23525 (N_23525,N_23299,N_23309);
and U23526 (N_23526,N_23353,N_23323);
or U23527 (N_23527,N_23224,N_23215);
or U23528 (N_23528,N_23369,N_23381);
and U23529 (N_23529,N_23242,N_23285);
nand U23530 (N_23530,N_23272,N_23318);
nand U23531 (N_23531,N_23203,N_23335);
or U23532 (N_23532,N_23355,N_23223);
nand U23533 (N_23533,N_23302,N_23208);
and U23534 (N_23534,N_23329,N_23282);
nand U23535 (N_23535,N_23361,N_23269);
or U23536 (N_23536,N_23398,N_23315);
nor U23537 (N_23537,N_23290,N_23348);
nand U23538 (N_23538,N_23222,N_23294);
nand U23539 (N_23539,N_23251,N_23221);
nor U23540 (N_23540,N_23375,N_23274);
nor U23541 (N_23541,N_23295,N_23373);
nor U23542 (N_23542,N_23319,N_23353);
and U23543 (N_23543,N_23300,N_23383);
nand U23544 (N_23544,N_23372,N_23281);
or U23545 (N_23545,N_23202,N_23294);
or U23546 (N_23546,N_23387,N_23281);
nand U23547 (N_23547,N_23372,N_23386);
nand U23548 (N_23548,N_23324,N_23352);
and U23549 (N_23549,N_23208,N_23233);
nand U23550 (N_23550,N_23225,N_23251);
and U23551 (N_23551,N_23349,N_23360);
nor U23552 (N_23552,N_23266,N_23225);
nand U23553 (N_23553,N_23286,N_23236);
or U23554 (N_23554,N_23395,N_23363);
nor U23555 (N_23555,N_23320,N_23221);
and U23556 (N_23556,N_23382,N_23392);
nor U23557 (N_23557,N_23322,N_23399);
nor U23558 (N_23558,N_23398,N_23363);
or U23559 (N_23559,N_23263,N_23284);
or U23560 (N_23560,N_23260,N_23303);
nor U23561 (N_23561,N_23309,N_23283);
and U23562 (N_23562,N_23281,N_23225);
and U23563 (N_23563,N_23251,N_23354);
nor U23564 (N_23564,N_23338,N_23221);
and U23565 (N_23565,N_23265,N_23208);
and U23566 (N_23566,N_23250,N_23243);
or U23567 (N_23567,N_23294,N_23218);
or U23568 (N_23568,N_23286,N_23340);
nor U23569 (N_23569,N_23267,N_23208);
and U23570 (N_23570,N_23326,N_23342);
and U23571 (N_23571,N_23309,N_23203);
nor U23572 (N_23572,N_23384,N_23284);
and U23573 (N_23573,N_23356,N_23357);
and U23574 (N_23574,N_23341,N_23279);
and U23575 (N_23575,N_23341,N_23390);
or U23576 (N_23576,N_23204,N_23255);
or U23577 (N_23577,N_23296,N_23332);
or U23578 (N_23578,N_23210,N_23296);
or U23579 (N_23579,N_23385,N_23227);
or U23580 (N_23580,N_23276,N_23233);
nand U23581 (N_23581,N_23353,N_23264);
nand U23582 (N_23582,N_23361,N_23247);
or U23583 (N_23583,N_23354,N_23355);
or U23584 (N_23584,N_23338,N_23385);
nand U23585 (N_23585,N_23229,N_23223);
or U23586 (N_23586,N_23288,N_23362);
or U23587 (N_23587,N_23292,N_23255);
nor U23588 (N_23588,N_23265,N_23383);
nand U23589 (N_23589,N_23314,N_23271);
or U23590 (N_23590,N_23253,N_23358);
nor U23591 (N_23591,N_23202,N_23246);
nand U23592 (N_23592,N_23398,N_23222);
and U23593 (N_23593,N_23201,N_23234);
and U23594 (N_23594,N_23244,N_23222);
and U23595 (N_23595,N_23289,N_23368);
and U23596 (N_23596,N_23303,N_23388);
nand U23597 (N_23597,N_23266,N_23393);
and U23598 (N_23598,N_23303,N_23200);
and U23599 (N_23599,N_23398,N_23296);
nand U23600 (N_23600,N_23589,N_23535);
nand U23601 (N_23601,N_23410,N_23594);
or U23602 (N_23602,N_23404,N_23415);
and U23603 (N_23603,N_23474,N_23492);
nand U23604 (N_23604,N_23424,N_23524);
or U23605 (N_23605,N_23591,N_23443);
and U23606 (N_23606,N_23427,N_23523);
nand U23607 (N_23607,N_23599,N_23555);
and U23608 (N_23608,N_23511,N_23406);
nor U23609 (N_23609,N_23408,N_23539);
or U23610 (N_23610,N_23537,N_23432);
and U23611 (N_23611,N_23436,N_23417);
or U23612 (N_23612,N_23510,N_23453);
or U23613 (N_23613,N_23440,N_23407);
nand U23614 (N_23614,N_23439,N_23503);
and U23615 (N_23615,N_23585,N_23531);
nor U23616 (N_23616,N_23463,N_23558);
or U23617 (N_23617,N_23400,N_23456);
or U23618 (N_23618,N_23540,N_23501);
or U23619 (N_23619,N_23551,N_23566);
and U23620 (N_23620,N_23491,N_23556);
and U23621 (N_23621,N_23465,N_23461);
nor U23622 (N_23622,N_23457,N_23513);
nor U23623 (N_23623,N_23434,N_23418);
or U23624 (N_23624,N_23420,N_23536);
nand U23625 (N_23625,N_23419,N_23578);
nand U23626 (N_23626,N_23553,N_23442);
nor U23627 (N_23627,N_23516,N_23543);
nand U23628 (N_23628,N_23401,N_23502);
nor U23629 (N_23629,N_23528,N_23507);
nor U23630 (N_23630,N_23582,N_23476);
or U23631 (N_23631,N_23431,N_23549);
nor U23632 (N_23632,N_23544,N_23506);
and U23633 (N_23633,N_23557,N_23519);
or U23634 (N_23634,N_23478,N_23455);
nand U23635 (N_23635,N_23490,N_23562);
nor U23636 (N_23636,N_23547,N_23517);
nand U23637 (N_23637,N_23448,N_23527);
nand U23638 (N_23638,N_23571,N_23560);
and U23639 (N_23639,N_23485,N_23489);
nand U23640 (N_23640,N_23581,N_23534);
nor U23641 (N_23641,N_23405,N_23550);
or U23642 (N_23642,N_23561,N_23409);
or U23643 (N_23643,N_23593,N_23435);
and U23644 (N_23644,N_23422,N_23493);
and U23645 (N_23645,N_23569,N_23446);
or U23646 (N_23646,N_23450,N_23580);
and U23647 (N_23647,N_23542,N_23473);
and U23648 (N_23648,N_23468,N_23497);
nor U23649 (N_23649,N_23423,N_23466);
nor U23650 (N_23650,N_23426,N_23402);
nand U23651 (N_23651,N_23509,N_23499);
nand U23652 (N_23652,N_23574,N_23521);
nand U23653 (N_23653,N_23564,N_23575);
nand U23654 (N_23654,N_23508,N_23546);
nand U23655 (N_23655,N_23486,N_23532);
or U23656 (N_23656,N_23487,N_23538);
nand U23657 (N_23657,N_23471,N_23579);
and U23658 (N_23658,N_23458,N_23412);
or U23659 (N_23659,N_23573,N_23597);
nor U23660 (N_23660,N_23460,N_23462);
and U23661 (N_23661,N_23498,N_23559);
and U23662 (N_23662,N_23421,N_23568);
and U23663 (N_23663,N_23477,N_23587);
or U23664 (N_23664,N_23577,N_23411);
or U23665 (N_23665,N_23595,N_23592);
or U23666 (N_23666,N_23541,N_23576);
or U23667 (N_23667,N_23526,N_23570);
and U23668 (N_23668,N_23530,N_23469);
or U23669 (N_23669,N_23583,N_23533);
or U23670 (N_23670,N_23480,N_23449);
nand U23671 (N_23671,N_23433,N_23467);
nor U23672 (N_23672,N_23552,N_23414);
and U23673 (N_23673,N_23572,N_23554);
nor U23674 (N_23674,N_23565,N_23494);
and U23675 (N_23675,N_23430,N_23548);
and U23676 (N_23676,N_23413,N_23437);
nand U23677 (N_23677,N_23584,N_23481);
nand U23678 (N_23678,N_23596,N_23403);
or U23679 (N_23679,N_23483,N_23484);
nand U23680 (N_23680,N_23444,N_23464);
xor U23681 (N_23681,N_23598,N_23512);
or U23682 (N_23682,N_23590,N_23500);
or U23683 (N_23683,N_23452,N_23515);
nor U23684 (N_23684,N_23514,N_23525);
nor U23685 (N_23685,N_23586,N_23496);
nor U23686 (N_23686,N_23488,N_23447);
nor U23687 (N_23687,N_23505,N_23425);
and U23688 (N_23688,N_23495,N_23567);
nor U23689 (N_23689,N_23482,N_23451);
nand U23690 (N_23690,N_23520,N_23459);
nand U23691 (N_23691,N_23454,N_23588);
and U23692 (N_23692,N_23429,N_23479);
nand U23693 (N_23693,N_23518,N_23545);
nor U23694 (N_23694,N_23438,N_23470);
nor U23695 (N_23695,N_23529,N_23428);
or U23696 (N_23696,N_23445,N_23472);
nand U23697 (N_23697,N_23563,N_23504);
nor U23698 (N_23698,N_23441,N_23522);
nand U23699 (N_23699,N_23475,N_23416);
or U23700 (N_23700,N_23437,N_23520);
nand U23701 (N_23701,N_23583,N_23536);
or U23702 (N_23702,N_23409,N_23417);
nand U23703 (N_23703,N_23492,N_23412);
or U23704 (N_23704,N_23559,N_23588);
nor U23705 (N_23705,N_23449,N_23494);
nor U23706 (N_23706,N_23406,N_23437);
and U23707 (N_23707,N_23529,N_23584);
nand U23708 (N_23708,N_23436,N_23481);
nor U23709 (N_23709,N_23596,N_23518);
or U23710 (N_23710,N_23436,N_23534);
and U23711 (N_23711,N_23446,N_23421);
nor U23712 (N_23712,N_23452,N_23499);
nand U23713 (N_23713,N_23577,N_23465);
or U23714 (N_23714,N_23535,N_23507);
and U23715 (N_23715,N_23467,N_23471);
nand U23716 (N_23716,N_23426,N_23498);
or U23717 (N_23717,N_23442,N_23422);
and U23718 (N_23718,N_23521,N_23582);
nor U23719 (N_23719,N_23540,N_23469);
and U23720 (N_23720,N_23558,N_23573);
and U23721 (N_23721,N_23438,N_23499);
and U23722 (N_23722,N_23532,N_23467);
nand U23723 (N_23723,N_23443,N_23518);
and U23724 (N_23724,N_23543,N_23425);
or U23725 (N_23725,N_23484,N_23486);
nor U23726 (N_23726,N_23478,N_23444);
nor U23727 (N_23727,N_23535,N_23555);
nor U23728 (N_23728,N_23485,N_23434);
nor U23729 (N_23729,N_23424,N_23471);
and U23730 (N_23730,N_23545,N_23596);
nor U23731 (N_23731,N_23474,N_23515);
nor U23732 (N_23732,N_23596,N_23552);
or U23733 (N_23733,N_23443,N_23428);
or U23734 (N_23734,N_23493,N_23469);
nand U23735 (N_23735,N_23454,N_23580);
or U23736 (N_23736,N_23413,N_23509);
nor U23737 (N_23737,N_23549,N_23436);
nand U23738 (N_23738,N_23526,N_23595);
nand U23739 (N_23739,N_23527,N_23468);
and U23740 (N_23740,N_23543,N_23592);
nor U23741 (N_23741,N_23542,N_23539);
or U23742 (N_23742,N_23489,N_23498);
nand U23743 (N_23743,N_23451,N_23526);
and U23744 (N_23744,N_23546,N_23597);
nand U23745 (N_23745,N_23542,N_23471);
nand U23746 (N_23746,N_23543,N_23579);
nor U23747 (N_23747,N_23597,N_23515);
nand U23748 (N_23748,N_23475,N_23512);
or U23749 (N_23749,N_23415,N_23523);
nand U23750 (N_23750,N_23474,N_23409);
nand U23751 (N_23751,N_23526,N_23475);
nand U23752 (N_23752,N_23562,N_23405);
and U23753 (N_23753,N_23402,N_23528);
or U23754 (N_23754,N_23595,N_23425);
nor U23755 (N_23755,N_23419,N_23415);
nor U23756 (N_23756,N_23528,N_23494);
nor U23757 (N_23757,N_23446,N_23517);
or U23758 (N_23758,N_23492,N_23490);
nand U23759 (N_23759,N_23428,N_23513);
nor U23760 (N_23760,N_23467,N_23595);
nor U23761 (N_23761,N_23520,N_23549);
nand U23762 (N_23762,N_23466,N_23400);
nand U23763 (N_23763,N_23549,N_23519);
nand U23764 (N_23764,N_23508,N_23521);
nand U23765 (N_23765,N_23404,N_23464);
nand U23766 (N_23766,N_23497,N_23425);
nand U23767 (N_23767,N_23585,N_23525);
or U23768 (N_23768,N_23552,N_23570);
nor U23769 (N_23769,N_23489,N_23481);
nand U23770 (N_23770,N_23523,N_23593);
nor U23771 (N_23771,N_23555,N_23433);
and U23772 (N_23772,N_23553,N_23481);
and U23773 (N_23773,N_23502,N_23497);
or U23774 (N_23774,N_23571,N_23440);
nand U23775 (N_23775,N_23406,N_23513);
nand U23776 (N_23776,N_23450,N_23551);
or U23777 (N_23777,N_23511,N_23499);
nand U23778 (N_23778,N_23411,N_23441);
nand U23779 (N_23779,N_23428,N_23456);
or U23780 (N_23780,N_23598,N_23451);
nor U23781 (N_23781,N_23498,N_23537);
or U23782 (N_23782,N_23524,N_23453);
nand U23783 (N_23783,N_23596,N_23444);
nand U23784 (N_23784,N_23453,N_23418);
nor U23785 (N_23785,N_23420,N_23435);
or U23786 (N_23786,N_23497,N_23543);
nor U23787 (N_23787,N_23431,N_23453);
nand U23788 (N_23788,N_23447,N_23451);
and U23789 (N_23789,N_23403,N_23489);
and U23790 (N_23790,N_23499,N_23536);
nand U23791 (N_23791,N_23544,N_23444);
nor U23792 (N_23792,N_23588,N_23537);
and U23793 (N_23793,N_23566,N_23424);
and U23794 (N_23794,N_23500,N_23457);
nand U23795 (N_23795,N_23599,N_23525);
nand U23796 (N_23796,N_23450,N_23531);
and U23797 (N_23797,N_23510,N_23534);
and U23798 (N_23798,N_23539,N_23562);
and U23799 (N_23799,N_23413,N_23434);
and U23800 (N_23800,N_23746,N_23775);
nor U23801 (N_23801,N_23632,N_23780);
nor U23802 (N_23802,N_23677,N_23769);
or U23803 (N_23803,N_23636,N_23797);
and U23804 (N_23804,N_23793,N_23633);
and U23805 (N_23805,N_23680,N_23760);
or U23806 (N_23806,N_23694,N_23754);
xnor U23807 (N_23807,N_23741,N_23728);
or U23808 (N_23808,N_23716,N_23798);
xor U23809 (N_23809,N_23799,N_23655);
or U23810 (N_23810,N_23722,N_23704);
nand U23811 (N_23811,N_23649,N_23740);
and U23812 (N_23812,N_23618,N_23707);
or U23813 (N_23813,N_23782,N_23752);
nand U23814 (N_23814,N_23624,N_23773);
or U23815 (N_23815,N_23674,N_23725);
or U23816 (N_23816,N_23604,N_23622);
nand U23817 (N_23817,N_23646,N_23685);
or U23818 (N_23818,N_23724,N_23714);
or U23819 (N_23819,N_23616,N_23692);
nor U23820 (N_23820,N_23702,N_23788);
nand U23821 (N_23821,N_23734,N_23687);
and U23822 (N_23822,N_23600,N_23672);
and U23823 (N_23823,N_23638,N_23750);
nor U23824 (N_23824,N_23609,N_23777);
and U23825 (N_23825,N_23665,N_23663);
nand U23826 (N_23826,N_23779,N_23682);
nor U23827 (N_23827,N_23642,N_23676);
and U23828 (N_23828,N_23664,N_23648);
nand U23829 (N_23829,N_23711,N_23698);
or U23830 (N_23830,N_23673,N_23643);
nor U23831 (N_23831,N_23607,N_23768);
and U23832 (N_23832,N_23617,N_23789);
or U23833 (N_23833,N_23668,N_23690);
xnor U23834 (N_23834,N_23771,N_23742);
or U23835 (N_23835,N_23686,N_23675);
and U23836 (N_23836,N_23611,N_23612);
nand U23837 (N_23837,N_23651,N_23657);
nand U23838 (N_23838,N_23745,N_23653);
nand U23839 (N_23839,N_23732,N_23733);
nor U23840 (N_23840,N_23739,N_23645);
nand U23841 (N_23841,N_23628,N_23776);
nand U23842 (N_23842,N_23757,N_23613);
nand U23843 (N_23843,N_23783,N_23689);
nand U23844 (N_23844,N_23606,N_23747);
xor U23845 (N_23845,N_23667,N_23627);
and U23846 (N_23846,N_23659,N_23608);
and U23847 (N_23847,N_23736,N_23637);
nor U23848 (N_23848,N_23790,N_23630);
nand U23849 (N_23849,N_23635,N_23602);
or U23850 (N_23850,N_23703,N_23666);
and U23851 (N_23851,N_23691,N_23761);
or U23852 (N_23852,N_23652,N_23601);
or U23853 (N_23853,N_23727,N_23656);
and U23854 (N_23854,N_23759,N_23772);
or U23855 (N_23855,N_23658,N_23774);
or U23856 (N_23856,N_23765,N_23700);
nand U23857 (N_23857,N_23709,N_23626);
nand U23858 (N_23858,N_23660,N_23786);
nor U23859 (N_23859,N_23753,N_23620);
nor U23860 (N_23860,N_23719,N_23758);
and U23861 (N_23861,N_23726,N_23644);
nand U23862 (N_23862,N_23708,N_23621);
nand U23863 (N_23863,N_23785,N_23794);
nor U23864 (N_23864,N_23603,N_23705);
nor U23865 (N_23865,N_23737,N_23623);
nor U23866 (N_23866,N_23693,N_23715);
and U23867 (N_23867,N_23684,N_23770);
nand U23868 (N_23868,N_23751,N_23729);
nand U23869 (N_23869,N_23696,N_23763);
nor U23870 (N_23870,N_23756,N_23661);
and U23871 (N_23871,N_23695,N_23662);
nand U23872 (N_23872,N_23641,N_23681);
and U23873 (N_23873,N_23767,N_23766);
nor U23874 (N_23874,N_23697,N_23744);
and U23875 (N_23875,N_23631,N_23762);
and U23876 (N_23876,N_23683,N_23670);
or U23877 (N_23877,N_23795,N_23679);
nor U23878 (N_23878,N_23625,N_23678);
or U23879 (N_23879,N_23605,N_23723);
nor U23880 (N_23880,N_23688,N_23743);
nand U23881 (N_23881,N_23735,N_23634);
nor U23882 (N_23882,N_23720,N_23701);
and U23883 (N_23883,N_23614,N_23640);
nand U23884 (N_23884,N_23610,N_23749);
nor U23885 (N_23885,N_23738,N_23731);
nand U23886 (N_23886,N_23717,N_23781);
and U23887 (N_23887,N_23650,N_23706);
nor U23888 (N_23888,N_23784,N_23712);
nor U23889 (N_23889,N_23778,N_23721);
or U23890 (N_23890,N_23654,N_23619);
and U23891 (N_23891,N_23615,N_23671);
and U23892 (N_23892,N_23764,N_23718);
nand U23893 (N_23893,N_23792,N_23796);
or U23894 (N_23894,N_23791,N_23669);
xor U23895 (N_23895,N_23629,N_23748);
nor U23896 (N_23896,N_23730,N_23699);
and U23897 (N_23897,N_23710,N_23755);
nor U23898 (N_23898,N_23787,N_23713);
nor U23899 (N_23899,N_23647,N_23639);
or U23900 (N_23900,N_23733,N_23690);
or U23901 (N_23901,N_23784,N_23798);
nand U23902 (N_23902,N_23752,N_23762);
and U23903 (N_23903,N_23648,N_23754);
or U23904 (N_23904,N_23767,N_23707);
xnor U23905 (N_23905,N_23706,N_23620);
or U23906 (N_23906,N_23789,N_23633);
and U23907 (N_23907,N_23695,N_23716);
nand U23908 (N_23908,N_23750,N_23683);
or U23909 (N_23909,N_23734,N_23728);
nand U23910 (N_23910,N_23688,N_23726);
nor U23911 (N_23911,N_23737,N_23621);
nand U23912 (N_23912,N_23785,N_23774);
nand U23913 (N_23913,N_23751,N_23702);
nor U23914 (N_23914,N_23731,N_23715);
and U23915 (N_23915,N_23671,N_23626);
nor U23916 (N_23916,N_23647,N_23645);
or U23917 (N_23917,N_23638,N_23676);
nor U23918 (N_23918,N_23646,N_23738);
nor U23919 (N_23919,N_23764,N_23724);
nand U23920 (N_23920,N_23643,N_23654);
or U23921 (N_23921,N_23798,N_23767);
nand U23922 (N_23922,N_23785,N_23722);
nand U23923 (N_23923,N_23693,N_23647);
or U23924 (N_23924,N_23706,N_23641);
nand U23925 (N_23925,N_23713,N_23759);
nor U23926 (N_23926,N_23672,N_23713);
and U23927 (N_23927,N_23725,N_23750);
nand U23928 (N_23928,N_23624,N_23696);
or U23929 (N_23929,N_23797,N_23618);
and U23930 (N_23930,N_23702,N_23667);
and U23931 (N_23931,N_23768,N_23761);
and U23932 (N_23932,N_23680,N_23740);
nand U23933 (N_23933,N_23778,N_23645);
or U23934 (N_23934,N_23705,N_23723);
and U23935 (N_23935,N_23750,N_23652);
nor U23936 (N_23936,N_23791,N_23774);
or U23937 (N_23937,N_23634,N_23778);
nor U23938 (N_23938,N_23655,N_23745);
nand U23939 (N_23939,N_23657,N_23664);
nand U23940 (N_23940,N_23680,N_23739);
or U23941 (N_23941,N_23632,N_23734);
nand U23942 (N_23942,N_23608,N_23791);
and U23943 (N_23943,N_23654,N_23739);
and U23944 (N_23944,N_23652,N_23628);
or U23945 (N_23945,N_23602,N_23771);
nand U23946 (N_23946,N_23625,N_23735);
and U23947 (N_23947,N_23727,N_23744);
or U23948 (N_23948,N_23612,N_23798);
or U23949 (N_23949,N_23637,N_23605);
nand U23950 (N_23950,N_23604,N_23745);
nor U23951 (N_23951,N_23641,N_23704);
or U23952 (N_23952,N_23730,N_23781);
and U23953 (N_23953,N_23616,N_23712);
or U23954 (N_23954,N_23610,N_23746);
and U23955 (N_23955,N_23679,N_23602);
and U23956 (N_23956,N_23649,N_23791);
or U23957 (N_23957,N_23645,N_23766);
or U23958 (N_23958,N_23705,N_23792);
nor U23959 (N_23959,N_23685,N_23618);
nand U23960 (N_23960,N_23651,N_23718);
nand U23961 (N_23961,N_23737,N_23606);
nor U23962 (N_23962,N_23733,N_23652);
and U23963 (N_23963,N_23719,N_23672);
nand U23964 (N_23964,N_23693,N_23611);
nand U23965 (N_23965,N_23785,N_23702);
or U23966 (N_23966,N_23710,N_23791);
nand U23967 (N_23967,N_23682,N_23665);
nor U23968 (N_23968,N_23777,N_23798);
or U23969 (N_23969,N_23698,N_23789);
nor U23970 (N_23970,N_23619,N_23766);
nand U23971 (N_23971,N_23640,N_23703);
and U23972 (N_23972,N_23711,N_23619);
or U23973 (N_23973,N_23677,N_23770);
or U23974 (N_23974,N_23720,N_23628);
xor U23975 (N_23975,N_23689,N_23705);
nor U23976 (N_23976,N_23740,N_23644);
nand U23977 (N_23977,N_23728,N_23649);
nor U23978 (N_23978,N_23679,N_23785);
nand U23979 (N_23979,N_23603,N_23622);
and U23980 (N_23980,N_23646,N_23681);
nor U23981 (N_23981,N_23765,N_23708);
nor U23982 (N_23982,N_23741,N_23637);
nor U23983 (N_23983,N_23768,N_23602);
nand U23984 (N_23984,N_23764,N_23765);
and U23985 (N_23985,N_23760,N_23745);
nand U23986 (N_23986,N_23653,N_23704);
nand U23987 (N_23987,N_23663,N_23650);
nand U23988 (N_23988,N_23705,N_23730);
and U23989 (N_23989,N_23757,N_23748);
or U23990 (N_23990,N_23777,N_23675);
or U23991 (N_23991,N_23739,N_23702);
nor U23992 (N_23992,N_23604,N_23705);
and U23993 (N_23993,N_23717,N_23797);
nand U23994 (N_23994,N_23604,N_23737);
or U23995 (N_23995,N_23751,N_23626);
or U23996 (N_23996,N_23704,N_23657);
or U23997 (N_23997,N_23676,N_23778);
nor U23998 (N_23998,N_23712,N_23706);
nor U23999 (N_23999,N_23698,N_23680);
and U24000 (N_24000,N_23901,N_23981);
nor U24001 (N_24001,N_23977,N_23812);
and U24002 (N_24002,N_23867,N_23876);
or U24003 (N_24003,N_23990,N_23813);
or U24004 (N_24004,N_23970,N_23999);
nand U24005 (N_24005,N_23856,N_23834);
nor U24006 (N_24006,N_23826,N_23900);
nor U24007 (N_24007,N_23829,N_23963);
and U24008 (N_24008,N_23845,N_23904);
or U24009 (N_24009,N_23943,N_23953);
or U24010 (N_24010,N_23914,N_23831);
nor U24011 (N_24011,N_23884,N_23907);
nor U24012 (N_24012,N_23950,N_23869);
nor U24013 (N_24013,N_23806,N_23930);
nor U24014 (N_24014,N_23874,N_23957);
and U24015 (N_24015,N_23807,N_23891);
or U24016 (N_24016,N_23971,N_23935);
and U24017 (N_24017,N_23846,N_23879);
nand U24018 (N_24018,N_23903,N_23882);
or U24019 (N_24019,N_23853,N_23897);
nand U24020 (N_24020,N_23938,N_23960);
and U24021 (N_24021,N_23912,N_23989);
and U24022 (N_24022,N_23955,N_23862);
and U24023 (N_24023,N_23850,N_23858);
or U24024 (N_24024,N_23898,N_23985);
and U24025 (N_24025,N_23899,N_23896);
or U24026 (N_24026,N_23998,N_23937);
and U24027 (N_24027,N_23860,N_23934);
and U24028 (N_24028,N_23958,N_23841);
xor U24029 (N_24029,N_23811,N_23959);
nor U24030 (N_24030,N_23929,N_23933);
nor U24031 (N_24031,N_23984,N_23865);
and U24032 (N_24032,N_23997,N_23996);
and U24033 (N_24033,N_23817,N_23964);
and U24034 (N_24034,N_23942,N_23951);
and U24035 (N_24035,N_23828,N_23819);
or U24036 (N_24036,N_23859,N_23800);
and U24037 (N_24037,N_23824,N_23823);
nor U24038 (N_24038,N_23895,N_23928);
and U24039 (N_24039,N_23894,N_23804);
nor U24040 (N_24040,N_23983,N_23843);
nand U24041 (N_24041,N_23972,N_23848);
and U24042 (N_24042,N_23923,N_23818);
nand U24043 (N_24043,N_23851,N_23905);
or U24044 (N_24044,N_23978,N_23821);
nor U24045 (N_24045,N_23952,N_23889);
nor U24046 (N_24046,N_23885,N_23988);
and U24047 (N_24047,N_23892,N_23936);
and U24048 (N_24048,N_23808,N_23920);
nand U24049 (N_24049,N_23939,N_23864);
or U24050 (N_24050,N_23995,N_23968);
nor U24051 (N_24051,N_23815,N_23852);
and U24052 (N_24052,N_23872,N_23967);
nor U24053 (N_24053,N_23847,N_23866);
nor U24054 (N_24054,N_23922,N_23875);
nor U24055 (N_24055,N_23814,N_23809);
nand U24056 (N_24056,N_23954,N_23941);
nor U24057 (N_24057,N_23947,N_23991);
nand U24058 (N_24058,N_23890,N_23857);
and U24059 (N_24059,N_23916,N_23986);
nor U24060 (N_24060,N_23915,N_23810);
and U24061 (N_24061,N_23993,N_23982);
and U24062 (N_24062,N_23835,N_23927);
or U24063 (N_24063,N_23822,N_23913);
nor U24064 (N_24064,N_23802,N_23946);
or U24065 (N_24065,N_23909,N_23868);
nand U24066 (N_24066,N_23837,N_23918);
nand U24067 (N_24067,N_23979,N_23994);
nand U24068 (N_24068,N_23966,N_23883);
or U24069 (N_24069,N_23962,N_23805);
or U24070 (N_24070,N_23801,N_23840);
and U24071 (N_24071,N_23973,N_23842);
or U24072 (N_24072,N_23925,N_23871);
or U24073 (N_24073,N_23906,N_23877);
and U24074 (N_24074,N_23980,N_23880);
or U24075 (N_24075,N_23803,N_23917);
or U24076 (N_24076,N_23854,N_23976);
nor U24077 (N_24077,N_23832,N_23839);
nand U24078 (N_24078,N_23836,N_23908);
or U24079 (N_24079,N_23873,N_23969);
and U24080 (N_24080,N_23945,N_23992);
or U24081 (N_24081,N_23919,N_23887);
nor U24082 (N_24082,N_23924,N_23940);
and U24083 (N_24083,N_23974,N_23987);
or U24084 (N_24084,N_23861,N_23910);
and U24085 (N_24085,N_23878,N_23833);
or U24086 (N_24086,N_23886,N_23849);
and U24087 (N_24087,N_23911,N_23965);
or U24088 (N_24088,N_23944,N_23863);
or U24089 (N_24089,N_23902,N_23948);
or U24090 (N_24090,N_23855,N_23844);
or U24091 (N_24091,N_23820,N_23888);
nor U24092 (N_24092,N_23921,N_23975);
nand U24093 (N_24093,N_23825,N_23881);
nor U24094 (N_24094,N_23949,N_23830);
or U24095 (N_24095,N_23931,N_23932);
nand U24096 (N_24096,N_23926,N_23838);
or U24097 (N_24097,N_23816,N_23956);
nand U24098 (N_24098,N_23870,N_23827);
nor U24099 (N_24099,N_23961,N_23893);
and U24100 (N_24100,N_23836,N_23923);
nor U24101 (N_24101,N_23800,N_23985);
and U24102 (N_24102,N_23817,N_23960);
or U24103 (N_24103,N_23948,N_23996);
or U24104 (N_24104,N_23973,N_23963);
nor U24105 (N_24105,N_23974,N_23996);
nor U24106 (N_24106,N_23955,N_23967);
and U24107 (N_24107,N_23965,N_23825);
nor U24108 (N_24108,N_23808,N_23933);
nor U24109 (N_24109,N_23813,N_23914);
nor U24110 (N_24110,N_23960,N_23830);
and U24111 (N_24111,N_23849,N_23918);
nor U24112 (N_24112,N_23937,N_23943);
or U24113 (N_24113,N_23943,N_23997);
nand U24114 (N_24114,N_23962,N_23806);
nand U24115 (N_24115,N_23995,N_23864);
nand U24116 (N_24116,N_23801,N_23961);
and U24117 (N_24117,N_23953,N_23997);
and U24118 (N_24118,N_23950,N_23926);
nor U24119 (N_24119,N_23808,N_23834);
and U24120 (N_24120,N_23910,N_23915);
or U24121 (N_24121,N_23939,N_23854);
or U24122 (N_24122,N_23947,N_23855);
and U24123 (N_24123,N_23811,N_23905);
nor U24124 (N_24124,N_23883,N_23853);
or U24125 (N_24125,N_23943,N_23917);
or U24126 (N_24126,N_23904,N_23860);
nand U24127 (N_24127,N_23830,N_23868);
or U24128 (N_24128,N_23986,N_23843);
and U24129 (N_24129,N_23864,N_23863);
nand U24130 (N_24130,N_23957,N_23953);
or U24131 (N_24131,N_23926,N_23947);
and U24132 (N_24132,N_23920,N_23821);
nor U24133 (N_24133,N_23897,N_23869);
or U24134 (N_24134,N_23990,N_23857);
and U24135 (N_24135,N_23966,N_23933);
nand U24136 (N_24136,N_23904,N_23928);
or U24137 (N_24137,N_23959,N_23921);
nor U24138 (N_24138,N_23861,N_23925);
or U24139 (N_24139,N_23991,N_23896);
nand U24140 (N_24140,N_23950,N_23966);
and U24141 (N_24141,N_23941,N_23913);
nand U24142 (N_24142,N_23861,N_23931);
nor U24143 (N_24143,N_23814,N_23972);
and U24144 (N_24144,N_23984,N_23945);
or U24145 (N_24145,N_23810,N_23914);
nand U24146 (N_24146,N_23880,N_23988);
and U24147 (N_24147,N_23807,N_23914);
nor U24148 (N_24148,N_23829,N_23917);
or U24149 (N_24149,N_23980,N_23909);
nand U24150 (N_24150,N_23834,N_23998);
nor U24151 (N_24151,N_23887,N_23912);
and U24152 (N_24152,N_23953,N_23899);
or U24153 (N_24153,N_23940,N_23860);
or U24154 (N_24154,N_23852,N_23849);
and U24155 (N_24155,N_23958,N_23868);
and U24156 (N_24156,N_23985,N_23956);
and U24157 (N_24157,N_23916,N_23859);
nand U24158 (N_24158,N_23955,N_23913);
or U24159 (N_24159,N_23848,N_23834);
or U24160 (N_24160,N_23978,N_23931);
nor U24161 (N_24161,N_23909,N_23835);
and U24162 (N_24162,N_23815,N_23945);
nand U24163 (N_24163,N_23901,N_23989);
nand U24164 (N_24164,N_23880,N_23930);
nand U24165 (N_24165,N_23892,N_23842);
nor U24166 (N_24166,N_23997,N_23976);
nand U24167 (N_24167,N_23833,N_23814);
or U24168 (N_24168,N_23964,N_23860);
nor U24169 (N_24169,N_23826,N_23975);
or U24170 (N_24170,N_23951,N_23923);
nand U24171 (N_24171,N_23925,N_23858);
or U24172 (N_24172,N_23901,N_23916);
or U24173 (N_24173,N_23963,N_23859);
nor U24174 (N_24174,N_23914,N_23985);
nor U24175 (N_24175,N_23805,N_23842);
and U24176 (N_24176,N_23878,N_23897);
or U24177 (N_24177,N_23827,N_23987);
or U24178 (N_24178,N_23830,N_23849);
nor U24179 (N_24179,N_23995,N_23842);
or U24180 (N_24180,N_23869,N_23894);
nor U24181 (N_24181,N_23854,N_23881);
and U24182 (N_24182,N_23995,N_23881);
and U24183 (N_24183,N_23953,N_23993);
nand U24184 (N_24184,N_23817,N_23834);
nor U24185 (N_24185,N_23978,N_23876);
and U24186 (N_24186,N_23925,N_23909);
or U24187 (N_24187,N_23932,N_23915);
nor U24188 (N_24188,N_23819,N_23833);
nand U24189 (N_24189,N_23939,N_23825);
nand U24190 (N_24190,N_23808,N_23943);
nand U24191 (N_24191,N_23843,N_23837);
nor U24192 (N_24192,N_23959,N_23865);
nor U24193 (N_24193,N_23890,N_23858);
or U24194 (N_24194,N_23900,N_23802);
nor U24195 (N_24195,N_23990,N_23947);
nor U24196 (N_24196,N_23861,N_23897);
nand U24197 (N_24197,N_23905,N_23996);
nand U24198 (N_24198,N_23932,N_23984);
nand U24199 (N_24199,N_23935,N_23800);
and U24200 (N_24200,N_24159,N_24165);
nand U24201 (N_24201,N_24116,N_24038);
nand U24202 (N_24202,N_24077,N_24083);
or U24203 (N_24203,N_24158,N_24109);
or U24204 (N_24204,N_24113,N_24167);
nand U24205 (N_24205,N_24126,N_24039);
and U24206 (N_24206,N_24028,N_24164);
and U24207 (N_24207,N_24068,N_24074);
nor U24208 (N_24208,N_24062,N_24081);
nand U24209 (N_24209,N_24193,N_24034);
nor U24210 (N_24210,N_24124,N_24067);
and U24211 (N_24211,N_24198,N_24080);
nor U24212 (N_24212,N_24170,N_24131);
and U24213 (N_24213,N_24138,N_24139);
nand U24214 (N_24214,N_24020,N_24182);
nor U24215 (N_24215,N_24179,N_24105);
and U24216 (N_24216,N_24063,N_24168);
xor U24217 (N_24217,N_24075,N_24045);
or U24218 (N_24218,N_24030,N_24108);
and U24219 (N_24219,N_24180,N_24102);
nand U24220 (N_24220,N_24043,N_24119);
or U24221 (N_24221,N_24190,N_24042);
nor U24222 (N_24222,N_24064,N_24162);
and U24223 (N_24223,N_24163,N_24145);
and U24224 (N_24224,N_24153,N_24014);
and U24225 (N_24225,N_24098,N_24169);
nor U24226 (N_24226,N_24194,N_24007);
nor U24227 (N_24227,N_24029,N_24050);
or U24228 (N_24228,N_24053,N_24186);
and U24229 (N_24229,N_24023,N_24104);
or U24230 (N_24230,N_24025,N_24171);
nor U24231 (N_24231,N_24079,N_24175);
xor U24232 (N_24232,N_24066,N_24183);
nor U24233 (N_24233,N_24122,N_24059);
nand U24234 (N_24234,N_24152,N_24094);
nand U24235 (N_24235,N_24147,N_24088);
and U24236 (N_24236,N_24149,N_24093);
or U24237 (N_24237,N_24128,N_24140);
nand U24238 (N_24238,N_24044,N_24151);
nand U24239 (N_24239,N_24117,N_24001);
and U24240 (N_24240,N_24087,N_24176);
and U24241 (N_24241,N_24107,N_24054);
and U24242 (N_24242,N_24056,N_24095);
nor U24243 (N_24243,N_24103,N_24082);
xor U24244 (N_24244,N_24099,N_24195);
nor U24245 (N_24245,N_24010,N_24049);
or U24246 (N_24246,N_24037,N_24052);
or U24247 (N_24247,N_24137,N_24005);
nand U24248 (N_24248,N_24060,N_24129);
nand U24249 (N_24249,N_24016,N_24185);
nand U24250 (N_24250,N_24013,N_24199);
nor U24251 (N_24251,N_24046,N_24154);
or U24252 (N_24252,N_24166,N_24112);
or U24253 (N_24253,N_24156,N_24026);
and U24254 (N_24254,N_24033,N_24084);
nand U24255 (N_24255,N_24173,N_24000);
and U24256 (N_24256,N_24127,N_24178);
or U24257 (N_24257,N_24032,N_24090);
or U24258 (N_24258,N_24143,N_24161);
nand U24259 (N_24259,N_24027,N_24189);
nor U24260 (N_24260,N_24071,N_24115);
xor U24261 (N_24261,N_24004,N_24196);
and U24262 (N_24262,N_24073,N_24036);
or U24263 (N_24263,N_24142,N_24132);
nand U24264 (N_24264,N_24015,N_24006);
and U24265 (N_24265,N_24047,N_24091);
or U24266 (N_24266,N_24121,N_24002);
nand U24267 (N_24267,N_24110,N_24191);
or U24268 (N_24268,N_24061,N_24076);
or U24269 (N_24269,N_24141,N_24011);
nand U24270 (N_24270,N_24085,N_24078);
xor U24271 (N_24271,N_24065,N_24181);
and U24272 (N_24272,N_24031,N_24012);
nor U24273 (N_24273,N_24174,N_24144);
nor U24274 (N_24274,N_24177,N_24184);
or U24275 (N_24275,N_24187,N_24072);
nor U24276 (N_24276,N_24192,N_24022);
and U24277 (N_24277,N_24021,N_24041);
or U24278 (N_24278,N_24086,N_24009);
nand U24279 (N_24279,N_24130,N_24155);
nor U24280 (N_24280,N_24070,N_24035);
nor U24281 (N_24281,N_24057,N_24106);
or U24282 (N_24282,N_24048,N_24096);
and U24283 (N_24283,N_24133,N_24069);
nor U24284 (N_24284,N_24114,N_24188);
nand U24285 (N_24285,N_24017,N_24146);
or U24286 (N_24286,N_24089,N_24136);
nand U24287 (N_24287,N_24003,N_24040);
nor U24288 (N_24288,N_24058,N_24097);
nand U24289 (N_24289,N_24150,N_24019);
nor U24290 (N_24290,N_24125,N_24101);
nand U24291 (N_24291,N_24160,N_24118);
nor U24292 (N_24292,N_24024,N_24135);
or U24293 (N_24293,N_24148,N_24172);
and U24294 (N_24294,N_24111,N_24008);
and U24295 (N_24295,N_24120,N_24018);
nand U24296 (N_24296,N_24123,N_24092);
nand U24297 (N_24297,N_24055,N_24197);
and U24298 (N_24298,N_24051,N_24134);
and U24299 (N_24299,N_24157,N_24100);
nor U24300 (N_24300,N_24019,N_24087);
or U24301 (N_24301,N_24028,N_24197);
nor U24302 (N_24302,N_24121,N_24150);
or U24303 (N_24303,N_24081,N_24094);
and U24304 (N_24304,N_24041,N_24011);
nand U24305 (N_24305,N_24152,N_24026);
and U24306 (N_24306,N_24096,N_24144);
and U24307 (N_24307,N_24036,N_24179);
or U24308 (N_24308,N_24176,N_24024);
nor U24309 (N_24309,N_24127,N_24112);
nand U24310 (N_24310,N_24199,N_24113);
nor U24311 (N_24311,N_24016,N_24120);
or U24312 (N_24312,N_24014,N_24154);
and U24313 (N_24313,N_24166,N_24007);
nand U24314 (N_24314,N_24016,N_24114);
nand U24315 (N_24315,N_24127,N_24175);
and U24316 (N_24316,N_24186,N_24182);
nor U24317 (N_24317,N_24169,N_24139);
and U24318 (N_24318,N_24151,N_24124);
and U24319 (N_24319,N_24187,N_24103);
nand U24320 (N_24320,N_24086,N_24066);
and U24321 (N_24321,N_24028,N_24042);
and U24322 (N_24322,N_24077,N_24188);
or U24323 (N_24323,N_24078,N_24027);
or U24324 (N_24324,N_24015,N_24041);
nand U24325 (N_24325,N_24027,N_24143);
or U24326 (N_24326,N_24153,N_24004);
nand U24327 (N_24327,N_24133,N_24091);
or U24328 (N_24328,N_24157,N_24092);
or U24329 (N_24329,N_24034,N_24081);
and U24330 (N_24330,N_24192,N_24178);
and U24331 (N_24331,N_24167,N_24073);
nor U24332 (N_24332,N_24115,N_24163);
nand U24333 (N_24333,N_24075,N_24123);
or U24334 (N_24334,N_24171,N_24001);
nor U24335 (N_24335,N_24071,N_24193);
and U24336 (N_24336,N_24115,N_24171);
nand U24337 (N_24337,N_24070,N_24189);
nor U24338 (N_24338,N_24145,N_24131);
or U24339 (N_24339,N_24032,N_24195);
nor U24340 (N_24340,N_24165,N_24137);
and U24341 (N_24341,N_24007,N_24072);
nor U24342 (N_24342,N_24167,N_24181);
or U24343 (N_24343,N_24143,N_24087);
nand U24344 (N_24344,N_24164,N_24189);
and U24345 (N_24345,N_24113,N_24069);
nand U24346 (N_24346,N_24125,N_24086);
nor U24347 (N_24347,N_24079,N_24108);
and U24348 (N_24348,N_24075,N_24072);
nor U24349 (N_24349,N_24163,N_24002);
and U24350 (N_24350,N_24041,N_24162);
nor U24351 (N_24351,N_24120,N_24197);
nand U24352 (N_24352,N_24196,N_24138);
nor U24353 (N_24353,N_24136,N_24043);
or U24354 (N_24354,N_24042,N_24093);
nand U24355 (N_24355,N_24019,N_24024);
nor U24356 (N_24356,N_24078,N_24007);
and U24357 (N_24357,N_24015,N_24176);
nor U24358 (N_24358,N_24036,N_24011);
or U24359 (N_24359,N_24188,N_24090);
nor U24360 (N_24360,N_24147,N_24003);
or U24361 (N_24361,N_24045,N_24120);
or U24362 (N_24362,N_24172,N_24005);
nand U24363 (N_24363,N_24040,N_24061);
nor U24364 (N_24364,N_24168,N_24049);
or U24365 (N_24365,N_24117,N_24158);
nand U24366 (N_24366,N_24190,N_24089);
or U24367 (N_24367,N_24029,N_24129);
nor U24368 (N_24368,N_24183,N_24194);
nor U24369 (N_24369,N_24193,N_24165);
and U24370 (N_24370,N_24021,N_24147);
and U24371 (N_24371,N_24140,N_24078);
nand U24372 (N_24372,N_24082,N_24193);
and U24373 (N_24373,N_24085,N_24002);
or U24374 (N_24374,N_24128,N_24070);
nand U24375 (N_24375,N_24154,N_24020);
and U24376 (N_24376,N_24148,N_24065);
or U24377 (N_24377,N_24035,N_24139);
nor U24378 (N_24378,N_24160,N_24133);
nand U24379 (N_24379,N_24104,N_24009);
or U24380 (N_24380,N_24006,N_24158);
nand U24381 (N_24381,N_24089,N_24199);
and U24382 (N_24382,N_24080,N_24135);
or U24383 (N_24383,N_24191,N_24102);
nand U24384 (N_24384,N_24034,N_24004);
nor U24385 (N_24385,N_24199,N_24188);
and U24386 (N_24386,N_24154,N_24179);
nand U24387 (N_24387,N_24073,N_24162);
or U24388 (N_24388,N_24127,N_24117);
or U24389 (N_24389,N_24125,N_24022);
or U24390 (N_24390,N_24093,N_24111);
or U24391 (N_24391,N_24043,N_24118);
or U24392 (N_24392,N_24109,N_24183);
nand U24393 (N_24393,N_24197,N_24161);
nand U24394 (N_24394,N_24194,N_24100);
nor U24395 (N_24395,N_24094,N_24071);
or U24396 (N_24396,N_24097,N_24102);
or U24397 (N_24397,N_24106,N_24138);
and U24398 (N_24398,N_24117,N_24181);
or U24399 (N_24399,N_24002,N_24034);
nor U24400 (N_24400,N_24381,N_24243);
xor U24401 (N_24401,N_24344,N_24386);
nand U24402 (N_24402,N_24220,N_24390);
nand U24403 (N_24403,N_24217,N_24302);
xnor U24404 (N_24404,N_24277,N_24256);
or U24405 (N_24405,N_24311,N_24367);
nand U24406 (N_24406,N_24341,N_24272);
or U24407 (N_24407,N_24225,N_24259);
nand U24408 (N_24408,N_24203,N_24373);
nand U24409 (N_24409,N_24249,N_24216);
and U24410 (N_24410,N_24202,N_24205);
nand U24411 (N_24411,N_24287,N_24339);
and U24412 (N_24412,N_24263,N_24240);
nor U24413 (N_24413,N_24210,N_24332);
nand U24414 (N_24414,N_24251,N_24239);
nand U24415 (N_24415,N_24276,N_24310);
nor U24416 (N_24416,N_24275,N_24234);
nor U24417 (N_24417,N_24340,N_24201);
nand U24418 (N_24418,N_24365,N_24290);
or U24419 (N_24419,N_24289,N_24244);
and U24420 (N_24420,N_24229,N_24308);
nor U24421 (N_24421,N_24253,N_24250);
or U24422 (N_24422,N_24285,N_24392);
nor U24423 (N_24423,N_24296,N_24343);
nand U24424 (N_24424,N_24221,N_24380);
nor U24425 (N_24425,N_24375,N_24314);
nor U24426 (N_24426,N_24294,N_24334);
nand U24427 (N_24427,N_24328,N_24355);
nand U24428 (N_24428,N_24204,N_24260);
nand U24429 (N_24429,N_24208,N_24255);
nand U24430 (N_24430,N_24316,N_24342);
and U24431 (N_24431,N_24298,N_24223);
and U24432 (N_24432,N_24378,N_24286);
or U24433 (N_24433,N_24379,N_24218);
or U24434 (N_24434,N_24293,N_24211);
nor U24435 (N_24435,N_24371,N_24319);
and U24436 (N_24436,N_24318,N_24213);
nor U24437 (N_24437,N_24335,N_24370);
and U24438 (N_24438,N_24393,N_24333);
nor U24439 (N_24439,N_24299,N_24215);
and U24440 (N_24440,N_24317,N_24200);
nand U24441 (N_24441,N_24304,N_24329);
or U24442 (N_24442,N_24309,N_24228);
and U24443 (N_24443,N_24362,N_24238);
nor U24444 (N_24444,N_24323,N_24245);
or U24445 (N_24445,N_24288,N_24389);
nand U24446 (N_24446,N_24206,N_24391);
and U24447 (N_24447,N_24231,N_24399);
and U24448 (N_24448,N_24372,N_24274);
nor U24449 (N_24449,N_24324,N_24377);
and U24450 (N_24450,N_24254,N_24320);
or U24451 (N_24451,N_24325,N_24257);
nand U24452 (N_24452,N_24265,N_24395);
nor U24453 (N_24453,N_24350,N_24360);
or U24454 (N_24454,N_24322,N_24338);
or U24455 (N_24455,N_24292,N_24353);
or U24456 (N_24456,N_24214,N_24305);
or U24457 (N_24457,N_24351,N_24226);
or U24458 (N_24458,N_24383,N_24356);
nand U24459 (N_24459,N_24326,N_24232);
and U24460 (N_24460,N_24266,N_24282);
and U24461 (N_24461,N_24284,N_24261);
nand U24462 (N_24462,N_24387,N_24306);
nor U24463 (N_24463,N_24264,N_24283);
or U24464 (N_24464,N_24397,N_24291);
and U24465 (N_24465,N_24273,N_24331);
or U24466 (N_24466,N_24352,N_24242);
nand U24467 (N_24467,N_24315,N_24348);
nand U24468 (N_24468,N_24269,N_24366);
nand U24469 (N_24469,N_24252,N_24224);
and U24470 (N_24470,N_24303,N_24233);
nor U24471 (N_24471,N_24230,N_24345);
and U24472 (N_24472,N_24297,N_24258);
nor U24473 (N_24473,N_24336,N_24347);
or U24474 (N_24474,N_24394,N_24374);
or U24475 (N_24475,N_24270,N_24337);
nand U24476 (N_24476,N_24237,N_24384);
and U24477 (N_24477,N_24271,N_24268);
nor U24478 (N_24478,N_24219,N_24398);
nor U24479 (N_24479,N_24222,N_24300);
nand U24480 (N_24480,N_24364,N_24236);
nor U24481 (N_24481,N_24262,N_24376);
nor U24482 (N_24482,N_24246,N_24212);
nor U24483 (N_24483,N_24369,N_24388);
or U24484 (N_24484,N_24267,N_24278);
nor U24485 (N_24485,N_24321,N_24209);
nand U24486 (N_24486,N_24385,N_24357);
and U24487 (N_24487,N_24279,N_24382);
and U24488 (N_24488,N_24307,N_24301);
nand U24489 (N_24489,N_24247,N_24295);
and U24490 (N_24490,N_24349,N_24363);
nor U24491 (N_24491,N_24396,N_24241);
nand U24492 (N_24492,N_24248,N_24281);
nand U24493 (N_24493,N_24235,N_24354);
or U24494 (N_24494,N_24361,N_24227);
nor U24495 (N_24495,N_24368,N_24313);
nor U24496 (N_24496,N_24330,N_24312);
nand U24497 (N_24497,N_24280,N_24346);
and U24498 (N_24498,N_24327,N_24207);
or U24499 (N_24499,N_24359,N_24358);
nand U24500 (N_24500,N_24212,N_24386);
nor U24501 (N_24501,N_24247,N_24254);
nand U24502 (N_24502,N_24236,N_24315);
or U24503 (N_24503,N_24353,N_24338);
nor U24504 (N_24504,N_24221,N_24389);
nor U24505 (N_24505,N_24293,N_24311);
or U24506 (N_24506,N_24333,N_24298);
nor U24507 (N_24507,N_24267,N_24230);
and U24508 (N_24508,N_24276,N_24242);
nor U24509 (N_24509,N_24296,N_24371);
and U24510 (N_24510,N_24202,N_24309);
or U24511 (N_24511,N_24283,N_24353);
or U24512 (N_24512,N_24219,N_24232);
nor U24513 (N_24513,N_24391,N_24334);
and U24514 (N_24514,N_24241,N_24238);
nor U24515 (N_24515,N_24357,N_24330);
nand U24516 (N_24516,N_24201,N_24230);
nand U24517 (N_24517,N_24386,N_24293);
or U24518 (N_24518,N_24269,N_24287);
nand U24519 (N_24519,N_24341,N_24298);
nor U24520 (N_24520,N_24209,N_24386);
or U24521 (N_24521,N_24395,N_24262);
or U24522 (N_24522,N_24236,N_24382);
nand U24523 (N_24523,N_24395,N_24225);
or U24524 (N_24524,N_24393,N_24261);
nor U24525 (N_24525,N_24385,N_24254);
nor U24526 (N_24526,N_24299,N_24309);
nor U24527 (N_24527,N_24348,N_24286);
nand U24528 (N_24528,N_24362,N_24319);
nand U24529 (N_24529,N_24318,N_24337);
nand U24530 (N_24530,N_24237,N_24356);
nand U24531 (N_24531,N_24231,N_24218);
nand U24532 (N_24532,N_24388,N_24337);
and U24533 (N_24533,N_24357,N_24302);
nand U24534 (N_24534,N_24274,N_24237);
or U24535 (N_24535,N_24286,N_24258);
or U24536 (N_24536,N_24343,N_24269);
or U24537 (N_24537,N_24282,N_24355);
and U24538 (N_24538,N_24399,N_24350);
and U24539 (N_24539,N_24267,N_24307);
nor U24540 (N_24540,N_24215,N_24383);
nand U24541 (N_24541,N_24238,N_24244);
nand U24542 (N_24542,N_24396,N_24208);
nor U24543 (N_24543,N_24325,N_24215);
and U24544 (N_24544,N_24308,N_24267);
or U24545 (N_24545,N_24318,N_24277);
and U24546 (N_24546,N_24275,N_24212);
or U24547 (N_24547,N_24288,N_24229);
nand U24548 (N_24548,N_24302,N_24256);
and U24549 (N_24549,N_24241,N_24217);
and U24550 (N_24550,N_24308,N_24300);
nor U24551 (N_24551,N_24364,N_24308);
nand U24552 (N_24552,N_24399,N_24342);
and U24553 (N_24553,N_24381,N_24274);
nand U24554 (N_24554,N_24215,N_24358);
nand U24555 (N_24555,N_24290,N_24293);
and U24556 (N_24556,N_24267,N_24333);
and U24557 (N_24557,N_24342,N_24387);
nand U24558 (N_24558,N_24374,N_24259);
nand U24559 (N_24559,N_24399,N_24395);
nand U24560 (N_24560,N_24257,N_24326);
and U24561 (N_24561,N_24387,N_24212);
and U24562 (N_24562,N_24241,N_24224);
nor U24563 (N_24563,N_24352,N_24291);
nand U24564 (N_24564,N_24271,N_24316);
and U24565 (N_24565,N_24375,N_24354);
or U24566 (N_24566,N_24399,N_24228);
and U24567 (N_24567,N_24201,N_24363);
or U24568 (N_24568,N_24289,N_24383);
or U24569 (N_24569,N_24268,N_24260);
nor U24570 (N_24570,N_24366,N_24261);
nor U24571 (N_24571,N_24205,N_24269);
nand U24572 (N_24572,N_24289,N_24283);
or U24573 (N_24573,N_24208,N_24304);
or U24574 (N_24574,N_24327,N_24345);
nor U24575 (N_24575,N_24397,N_24370);
nor U24576 (N_24576,N_24393,N_24315);
or U24577 (N_24577,N_24320,N_24267);
and U24578 (N_24578,N_24384,N_24238);
nand U24579 (N_24579,N_24247,N_24332);
nor U24580 (N_24580,N_24366,N_24265);
nand U24581 (N_24581,N_24342,N_24271);
or U24582 (N_24582,N_24294,N_24320);
nor U24583 (N_24583,N_24364,N_24366);
and U24584 (N_24584,N_24344,N_24235);
or U24585 (N_24585,N_24316,N_24317);
and U24586 (N_24586,N_24257,N_24385);
and U24587 (N_24587,N_24285,N_24349);
nand U24588 (N_24588,N_24349,N_24262);
or U24589 (N_24589,N_24226,N_24258);
nor U24590 (N_24590,N_24322,N_24285);
and U24591 (N_24591,N_24263,N_24274);
nor U24592 (N_24592,N_24278,N_24271);
and U24593 (N_24593,N_24317,N_24362);
and U24594 (N_24594,N_24371,N_24274);
or U24595 (N_24595,N_24350,N_24354);
or U24596 (N_24596,N_24236,N_24262);
nand U24597 (N_24597,N_24214,N_24375);
nand U24598 (N_24598,N_24222,N_24288);
nor U24599 (N_24599,N_24398,N_24254);
and U24600 (N_24600,N_24470,N_24456);
nand U24601 (N_24601,N_24497,N_24504);
or U24602 (N_24602,N_24467,N_24458);
nand U24603 (N_24603,N_24483,N_24465);
or U24604 (N_24604,N_24546,N_24455);
and U24605 (N_24605,N_24518,N_24473);
or U24606 (N_24606,N_24535,N_24431);
nand U24607 (N_24607,N_24434,N_24451);
and U24608 (N_24608,N_24475,N_24493);
and U24609 (N_24609,N_24511,N_24583);
nand U24610 (N_24610,N_24510,N_24489);
and U24611 (N_24611,N_24527,N_24472);
and U24612 (N_24612,N_24592,N_24477);
and U24613 (N_24613,N_24449,N_24594);
nand U24614 (N_24614,N_24521,N_24550);
nand U24615 (N_24615,N_24507,N_24519);
nor U24616 (N_24616,N_24464,N_24516);
and U24617 (N_24617,N_24542,N_24404);
and U24618 (N_24618,N_24578,N_24453);
and U24619 (N_24619,N_24570,N_24462);
nor U24620 (N_24620,N_24500,N_24424);
and U24621 (N_24621,N_24530,N_24534);
or U24622 (N_24622,N_24556,N_24436);
nor U24623 (N_24623,N_24414,N_24421);
nand U24624 (N_24624,N_24433,N_24501);
nand U24625 (N_24625,N_24597,N_24599);
nor U24626 (N_24626,N_24405,N_24509);
nor U24627 (N_24627,N_24533,N_24491);
or U24628 (N_24628,N_24558,N_24595);
and U24629 (N_24629,N_24478,N_24568);
or U24630 (N_24630,N_24413,N_24480);
nor U24631 (N_24631,N_24569,N_24498);
nor U24632 (N_24632,N_24551,N_24564);
nand U24633 (N_24633,N_24440,N_24416);
or U24634 (N_24634,N_24466,N_24549);
nor U24635 (N_24635,N_24459,N_24446);
and U24636 (N_24636,N_24415,N_24585);
nand U24637 (N_24637,N_24574,N_24523);
or U24638 (N_24638,N_24441,N_24494);
or U24639 (N_24639,N_24409,N_24591);
and U24640 (N_24640,N_24596,N_24430);
nor U24641 (N_24641,N_24513,N_24577);
and U24642 (N_24642,N_24548,N_24575);
nand U24643 (N_24643,N_24418,N_24437);
nand U24644 (N_24644,N_24492,N_24487);
nor U24645 (N_24645,N_24508,N_24422);
nand U24646 (N_24646,N_24426,N_24539);
nand U24647 (N_24647,N_24536,N_24484);
nand U24648 (N_24648,N_24584,N_24543);
nor U24649 (N_24649,N_24520,N_24555);
nand U24650 (N_24650,N_24435,N_24410);
and U24651 (N_24651,N_24566,N_24529);
or U24652 (N_24652,N_24496,N_24559);
nand U24653 (N_24653,N_24402,N_24531);
nor U24654 (N_24654,N_24485,N_24463);
or U24655 (N_24655,N_24454,N_24432);
and U24656 (N_24656,N_24579,N_24517);
nor U24657 (N_24657,N_24447,N_24452);
nor U24658 (N_24658,N_24544,N_24428);
or U24659 (N_24659,N_24460,N_24528);
nand U24660 (N_24660,N_24427,N_24571);
and U24661 (N_24661,N_24554,N_24442);
nor U24662 (N_24662,N_24407,N_24417);
or U24663 (N_24663,N_24503,N_24547);
or U24664 (N_24664,N_24502,N_24469);
nand U24665 (N_24665,N_24406,N_24412);
nor U24666 (N_24666,N_24524,N_24450);
nor U24667 (N_24667,N_24429,N_24481);
or U24668 (N_24668,N_24580,N_24438);
or U24669 (N_24669,N_24423,N_24490);
and U24670 (N_24670,N_24589,N_24495);
nor U24671 (N_24671,N_24461,N_24486);
nor U24672 (N_24672,N_24532,N_24588);
nor U24673 (N_24673,N_24562,N_24479);
nor U24674 (N_24674,N_24514,N_24587);
and U24675 (N_24675,N_24563,N_24537);
or U24676 (N_24676,N_24411,N_24590);
or U24677 (N_24677,N_24443,N_24474);
or U24678 (N_24678,N_24541,N_24561);
or U24679 (N_24679,N_24586,N_24482);
and U24680 (N_24680,N_24476,N_24565);
or U24681 (N_24681,N_24515,N_24552);
and U24682 (N_24682,N_24420,N_24598);
or U24683 (N_24683,N_24419,N_24499);
and U24684 (N_24684,N_24444,N_24576);
and U24685 (N_24685,N_24522,N_24567);
or U24686 (N_24686,N_24538,N_24526);
or U24687 (N_24687,N_24525,N_24582);
nor U24688 (N_24688,N_24439,N_24488);
nand U24689 (N_24689,N_24545,N_24408);
and U24690 (N_24690,N_24593,N_24401);
or U24691 (N_24691,N_24506,N_24581);
and U24692 (N_24692,N_24471,N_24448);
and U24693 (N_24693,N_24400,N_24403);
xor U24694 (N_24694,N_24468,N_24560);
and U24695 (N_24695,N_24512,N_24445);
nand U24696 (N_24696,N_24425,N_24557);
and U24697 (N_24697,N_24553,N_24540);
or U24698 (N_24698,N_24505,N_24573);
and U24699 (N_24699,N_24457,N_24572);
nor U24700 (N_24700,N_24486,N_24587);
nor U24701 (N_24701,N_24500,N_24547);
or U24702 (N_24702,N_24487,N_24551);
nand U24703 (N_24703,N_24553,N_24521);
nor U24704 (N_24704,N_24436,N_24451);
nor U24705 (N_24705,N_24549,N_24488);
nand U24706 (N_24706,N_24463,N_24455);
and U24707 (N_24707,N_24492,N_24462);
nand U24708 (N_24708,N_24427,N_24513);
nand U24709 (N_24709,N_24542,N_24534);
nand U24710 (N_24710,N_24426,N_24546);
or U24711 (N_24711,N_24485,N_24411);
and U24712 (N_24712,N_24433,N_24525);
or U24713 (N_24713,N_24520,N_24515);
nand U24714 (N_24714,N_24443,N_24492);
nand U24715 (N_24715,N_24538,N_24501);
and U24716 (N_24716,N_24573,N_24422);
nand U24717 (N_24717,N_24501,N_24458);
or U24718 (N_24718,N_24493,N_24447);
and U24719 (N_24719,N_24476,N_24522);
and U24720 (N_24720,N_24461,N_24566);
nand U24721 (N_24721,N_24463,N_24554);
nand U24722 (N_24722,N_24475,N_24530);
or U24723 (N_24723,N_24439,N_24531);
nor U24724 (N_24724,N_24419,N_24503);
or U24725 (N_24725,N_24576,N_24415);
or U24726 (N_24726,N_24507,N_24460);
or U24727 (N_24727,N_24413,N_24559);
and U24728 (N_24728,N_24477,N_24567);
nand U24729 (N_24729,N_24470,N_24575);
and U24730 (N_24730,N_24452,N_24577);
xor U24731 (N_24731,N_24412,N_24444);
or U24732 (N_24732,N_24441,N_24495);
or U24733 (N_24733,N_24533,N_24463);
or U24734 (N_24734,N_24563,N_24408);
nor U24735 (N_24735,N_24454,N_24429);
or U24736 (N_24736,N_24452,N_24545);
and U24737 (N_24737,N_24569,N_24578);
nor U24738 (N_24738,N_24555,N_24415);
or U24739 (N_24739,N_24458,N_24477);
nor U24740 (N_24740,N_24523,N_24509);
and U24741 (N_24741,N_24590,N_24490);
or U24742 (N_24742,N_24594,N_24586);
nand U24743 (N_24743,N_24442,N_24543);
and U24744 (N_24744,N_24422,N_24482);
or U24745 (N_24745,N_24468,N_24555);
nor U24746 (N_24746,N_24445,N_24596);
nor U24747 (N_24747,N_24489,N_24497);
nor U24748 (N_24748,N_24424,N_24454);
or U24749 (N_24749,N_24483,N_24470);
or U24750 (N_24750,N_24447,N_24539);
and U24751 (N_24751,N_24568,N_24441);
or U24752 (N_24752,N_24424,N_24564);
nor U24753 (N_24753,N_24474,N_24524);
xor U24754 (N_24754,N_24484,N_24512);
nor U24755 (N_24755,N_24531,N_24403);
or U24756 (N_24756,N_24493,N_24405);
nand U24757 (N_24757,N_24482,N_24541);
and U24758 (N_24758,N_24473,N_24446);
nand U24759 (N_24759,N_24474,N_24484);
or U24760 (N_24760,N_24485,N_24427);
nor U24761 (N_24761,N_24536,N_24541);
and U24762 (N_24762,N_24401,N_24427);
nand U24763 (N_24763,N_24585,N_24464);
and U24764 (N_24764,N_24595,N_24420);
nor U24765 (N_24765,N_24448,N_24544);
and U24766 (N_24766,N_24475,N_24574);
or U24767 (N_24767,N_24456,N_24563);
or U24768 (N_24768,N_24421,N_24551);
nand U24769 (N_24769,N_24464,N_24450);
nand U24770 (N_24770,N_24480,N_24419);
nor U24771 (N_24771,N_24402,N_24453);
nand U24772 (N_24772,N_24575,N_24547);
nand U24773 (N_24773,N_24522,N_24591);
nand U24774 (N_24774,N_24582,N_24581);
or U24775 (N_24775,N_24458,N_24599);
and U24776 (N_24776,N_24574,N_24427);
nor U24777 (N_24777,N_24448,N_24443);
and U24778 (N_24778,N_24517,N_24499);
and U24779 (N_24779,N_24520,N_24401);
and U24780 (N_24780,N_24438,N_24568);
and U24781 (N_24781,N_24541,N_24469);
nand U24782 (N_24782,N_24595,N_24541);
or U24783 (N_24783,N_24528,N_24511);
or U24784 (N_24784,N_24444,N_24512);
nor U24785 (N_24785,N_24465,N_24408);
nand U24786 (N_24786,N_24461,N_24407);
nor U24787 (N_24787,N_24575,N_24577);
or U24788 (N_24788,N_24469,N_24417);
nand U24789 (N_24789,N_24586,N_24564);
and U24790 (N_24790,N_24422,N_24552);
and U24791 (N_24791,N_24408,N_24431);
nor U24792 (N_24792,N_24595,N_24574);
or U24793 (N_24793,N_24497,N_24483);
nor U24794 (N_24794,N_24552,N_24554);
nor U24795 (N_24795,N_24529,N_24543);
and U24796 (N_24796,N_24493,N_24441);
nand U24797 (N_24797,N_24529,N_24415);
and U24798 (N_24798,N_24595,N_24578);
nor U24799 (N_24799,N_24422,N_24468);
nor U24800 (N_24800,N_24677,N_24625);
and U24801 (N_24801,N_24714,N_24771);
and U24802 (N_24802,N_24605,N_24708);
and U24803 (N_24803,N_24770,N_24729);
nand U24804 (N_24804,N_24673,N_24669);
or U24805 (N_24805,N_24765,N_24734);
and U24806 (N_24806,N_24624,N_24755);
or U24807 (N_24807,N_24618,N_24644);
and U24808 (N_24808,N_24776,N_24617);
or U24809 (N_24809,N_24719,N_24649);
and U24810 (N_24810,N_24757,N_24693);
nor U24811 (N_24811,N_24799,N_24684);
or U24812 (N_24812,N_24657,N_24759);
nor U24813 (N_24813,N_24750,N_24730);
nor U24814 (N_24814,N_24790,N_24738);
nand U24815 (N_24815,N_24655,N_24678);
and U24816 (N_24816,N_24740,N_24762);
nor U24817 (N_24817,N_24721,N_24751);
and U24818 (N_24818,N_24722,N_24769);
nand U24819 (N_24819,N_24793,N_24603);
nand U24820 (N_24820,N_24746,N_24748);
nor U24821 (N_24821,N_24761,N_24646);
and U24822 (N_24822,N_24731,N_24703);
or U24823 (N_24823,N_24629,N_24783);
nor U24824 (N_24824,N_24781,N_24668);
nand U24825 (N_24825,N_24660,N_24743);
and U24826 (N_24826,N_24697,N_24700);
nand U24827 (N_24827,N_24623,N_24726);
and U24828 (N_24828,N_24752,N_24779);
and U24829 (N_24829,N_24616,N_24753);
nand U24830 (N_24830,N_24733,N_24737);
and U24831 (N_24831,N_24780,N_24732);
nor U24832 (N_24832,N_24688,N_24787);
or U24833 (N_24833,N_24745,N_24635);
and U24834 (N_24834,N_24621,N_24648);
or U24835 (N_24835,N_24797,N_24675);
or U24836 (N_24836,N_24736,N_24701);
nand U24837 (N_24837,N_24710,N_24613);
nand U24838 (N_24838,N_24667,N_24695);
nor U24839 (N_24839,N_24606,N_24768);
nand U24840 (N_24840,N_24760,N_24723);
nand U24841 (N_24841,N_24676,N_24614);
nor U24842 (N_24842,N_24601,N_24767);
or U24843 (N_24843,N_24786,N_24682);
or U24844 (N_24844,N_24662,N_24609);
nand U24845 (N_24845,N_24691,N_24720);
nor U24846 (N_24846,N_24631,N_24670);
or U24847 (N_24847,N_24756,N_24619);
nand U24848 (N_24848,N_24633,N_24634);
or U24849 (N_24849,N_24653,N_24689);
nor U24850 (N_24850,N_24764,N_24711);
and U24851 (N_24851,N_24702,N_24792);
nor U24852 (N_24852,N_24774,N_24641);
and U24853 (N_24853,N_24604,N_24742);
and U24854 (N_24854,N_24663,N_24686);
nor U24855 (N_24855,N_24699,N_24666);
nand U24856 (N_24856,N_24639,N_24717);
nand U24857 (N_24857,N_24766,N_24758);
nand U24858 (N_24858,N_24656,N_24671);
and U24859 (N_24859,N_24795,N_24725);
or U24860 (N_24860,N_24704,N_24687);
nand U24861 (N_24861,N_24778,N_24643);
and U24862 (N_24862,N_24685,N_24782);
and U24863 (N_24863,N_24652,N_24785);
nor U24864 (N_24864,N_24715,N_24681);
or U24865 (N_24865,N_24716,N_24791);
or U24866 (N_24866,N_24680,N_24674);
nor U24867 (N_24867,N_24788,N_24658);
or U24868 (N_24868,N_24718,N_24630);
nor U24869 (N_24869,N_24741,N_24705);
nor U24870 (N_24870,N_24650,N_24698);
xor U24871 (N_24871,N_24727,N_24744);
and U24872 (N_24872,N_24707,N_24610);
nand U24873 (N_24873,N_24647,N_24713);
and U24874 (N_24874,N_24735,N_24638);
nor U24875 (N_24875,N_24608,N_24724);
nor U24876 (N_24876,N_24645,N_24709);
nand U24877 (N_24877,N_24620,N_24784);
or U24878 (N_24878,N_24754,N_24665);
nor U24879 (N_24879,N_24636,N_24749);
and U24880 (N_24880,N_24612,N_24773);
or U24881 (N_24881,N_24626,N_24600);
nor U24882 (N_24882,N_24706,N_24777);
or U24883 (N_24883,N_24664,N_24712);
and U24884 (N_24884,N_24651,N_24794);
nor U24885 (N_24885,N_24615,N_24637);
and U24886 (N_24886,N_24659,N_24728);
or U24887 (N_24887,N_24772,N_24796);
and U24888 (N_24888,N_24690,N_24694);
or U24889 (N_24889,N_24692,N_24763);
or U24890 (N_24890,N_24640,N_24661);
and U24891 (N_24891,N_24798,N_24627);
nor U24892 (N_24892,N_24789,N_24642);
nor U24893 (N_24893,N_24622,N_24628);
nor U24894 (N_24894,N_24683,N_24775);
or U24895 (N_24895,N_24632,N_24654);
and U24896 (N_24896,N_24607,N_24739);
or U24897 (N_24897,N_24602,N_24696);
nand U24898 (N_24898,N_24679,N_24747);
and U24899 (N_24899,N_24611,N_24672);
nor U24900 (N_24900,N_24716,N_24661);
or U24901 (N_24901,N_24722,N_24667);
nand U24902 (N_24902,N_24626,N_24704);
xnor U24903 (N_24903,N_24615,N_24712);
nand U24904 (N_24904,N_24606,N_24689);
or U24905 (N_24905,N_24717,N_24631);
nand U24906 (N_24906,N_24699,N_24799);
and U24907 (N_24907,N_24685,N_24759);
nor U24908 (N_24908,N_24746,N_24656);
nand U24909 (N_24909,N_24649,N_24789);
and U24910 (N_24910,N_24719,N_24624);
nand U24911 (N_24911,N_24701,N_24723);
nor U24912 (N_24912,N_24724,N_24755);
nand U24913 (N_24913,N_24697,N_24658);
and U24914 (N_24914,N_24793,N_24644);
nor U24915 (N_24915,N_24710,N_24794);
and U24916 (N_24916,N_24727,N_24664);
nor U24917 (N_24917,N_24790,N_24670);
nor U24918 (N_24918,N_24601,N_24757);
nand U24919 (N_24919,N_24605,N_24673);
or U24920 (N_24920,N_24630,N_24641);
or U24921 (N_24921,N_24721,N_24625);
and U24922 (N_24922,N_24704,N_24612);
nor U24923 (N_24923,N_24650,N_24710);
or U24924 (N_24924,N_24669,N_24765);
or U24925 (N_24925,N_24655,N_24752);
nand U24926 (N_24926,N_24608,N_24616);
or U24927 (N_24927,N_24727,N_24678);
and U24928 (N_24928,N_24619,N_24711);
or U24929 (N_24929,N_24755,N_24732);
and U24930 (N_24930,N_24671,N_24751);
and U24931 (N_24931,N_24623,N_24621);
nand U24932 (N_24932,N_24691,N_24630);
nand U24933 (N_24933,N_24609,N_24718);
and U24934 (N_24934,N_24656,N_24633);
nand U24935 (N_24935,N_24622,N_24726);
and U24936 (N_24936,N_24796,N_24779);
nand U24937 (N_24937,N_24602,N_24729);
nor U24938 (N_24938,N_24647,N_24694);
or U24939 (N_24939,N_24720,N_24708);
nor U24940 (N_24940,N_24659,N_24615);
or U24941 (N_24941,N_24694,N_24631);
and U24942 (N_24942,N_24687,N_24609);
nor U24943 (N_24943,N_24670,N_24775);
nand U24944 (N_24944,N_24794,N_24758);
and U24945 (N_24945,N_24754,N_24655);
or U24946 (N_24946,N_24637,N_24707);
nor U24947 (N_24947,N_24797,N_24620);
or U24948 (N_24948,N_24767,N_24632);
and U24949 (N_24949,N_24642,N_24625);
and U24950 (N_24950,N_24762,N_24650);
nor U24951 (N_24951,N_24756,N_24683);
nor U24952 (N_24952,N_24786,N_24674);
nor U24953 (N_24953,N_24707,N_24677);
and U24954 (N_24954,N_24684,N_24607);
and U24955 (N_24955,N_24719,N_24638);
or U24956 (N_24956,N_24601,N_24632);
nand U24957 (N_24957,N_24703,N_24667);
or U24958 (N_24958,N_24783,N_24668);
nand U24959 (N_24959,N_24716,N_24665);
or U24960 (N_24960,N_24691,N_24745);
or U24961 (N_24961,N_24776,N_24693);
nand U24962 (N_24962,N_24770,N_24708);
nand U24963 (N_24963,N_24726,N_24678);
nand U24964 (N_24964,N_24646,N_24779);
nand U24965 (N_24965,N_24768,N_24604);
and U24966 (N_24966,N_24733,N_24605);
nor U24967 (N_24967,N_24770,N_24655);
and U24968 (N_24968,N_24617,N_24626);
and U24969 (N_24969,N_24713,N_24634);
and U24970 (N_24970,N_24764,N_24739);
or U24971 (N_24971,N_24733,N_24703);
nor U24972 (N_24972,N_24746,N_24719);
nor U24973 (N_24973,N_24705,N_24679);
and U24974 (N_24974,N_24746,N_24600);
nor U24975 (N_24975,N_24677,N_24739);
nand U24976 (N_24976,N_24717,N_24762);
nor U24977 (N_24977,N_24762,N_24694);
xnor U24978 (N_24978,N_24656,N_24688);
nor U24979 (N_24979,N_24787,N_24677);
nand U24980 (N_24980,N_24663,N_24681);
and U24981 (N_24981,N_24779,N_24791);
nand U24982 (N_24982,N_24730,N_24752);
and U24983 (N_24983,N_24659,N_24706);
nand U24984 (N_24984,N_24606,N_24785);
or U24985 (N_24985,N_24736,N_24788);
nand U24986 (N_24986,N_24632,N_24631);
nor U24987 (N_24987,N_24714,N_24757);
or U24988 (N_24988,N_24612,N_24756);
nor U24989 (N_24989,N_24752,N_24621);
nor U24990 (N_24990,N_24778,N_24709);
or U24991 (N_24991,N_24600,N_24619);
nand U24992 (N_24992,N_24677,N_24672);
or U24993 (N_24993,N_24765,N_24680);
and U24994 (N_24994,N_24616,N_24659);
nor U24995 (N_24995,N_24718,N_24772);
and U24996 (N_24996,N_24704,N_24667);
and U24997 (N_24997,N_24661,N_24605);
nand U24998 (N_24998,N_24703,N_24628);
nand U24999 (N_24999,N_24699,N_24711);
nand UO_0 (O_0,N_24974,N_24882);
and UO_1 (O_1,N_24907,N_24804);
and UO_2 (O_2,N_24959,N_24931);
and UO_3 (O_3,N_24998,N_24828);
and UO_4 (O_4,N_24890,N_24855);
nand UO_5 (O_5,N_24909,N_24952);
nand UO_6 (O_6,N_24991,N_24878);
nand UO_7 (O_7,N_24930,N_24995);
or UO_8 (O_8,N_24865,N_24918);
and UO_9 (O_9,N_24928,N_24910);
and UO_10 (O_10,N_24946,N_24999);
nor UO_11 (O_11,N_24836,N_24872);
nand UO_12 (O_12,N_24874,N_24885);
or UO_13 (O_13,N_24832,N_24927);
or UO_14 (O_14,N_24802,N_24870);
and UO_15 (O_15,N_24863,N_24876);
nor UO_16 (O_16,N_24869,N_24902);
nand UO_17 (O_17,N_24895,N_24925);
or UO_18 (O_18,N_24912,N_24950);
or UO_19 (O_19,N_24958,N_24987);
nand UO_20 (O_20,N_24824,N_24818);
nand UO_21 (O_21,N_24911,N_24941);
and UO_22 (O_22,N_24973,N_24823);
or UO_23 (O_23,N_24924,N_24962);
and UO_24 (O_24,N_24810,N_24913);
and UO_25 (O_25,N_24985,N_24813);
and UO_26 (O_26,N_24881,N_24990);
nand UO_27 (O_27,N_24826,N_24969);
nand UO_28 (O_28,N_24850,N_24948);
nor UO_29 (O_29,N_24843,N_24866);
nand UO_30 (O_30,N_24822,N_24967);
nand UO_31 (O_31,N_24805,N_24961);
or UO_32 (O_32,N_24965,N_24968);
and UO_33 (O_33,N_24875,N_24966);
nand UO_34 (O_34,N_24880,N_24945);
or UO_35 (O_35,N_24846,N_24923);
or UO_36 (O_36,N_24915,N_24879);
nor UO_37 (O_37,N_24980,N_24817);
or UO_38 (O_38,N_24994,N_24920);
nor UO_39 (O_39,N_24979,N_24898);
and UO_40 (O_40,N_24949,N_24864);
nor UO_41 (O_41,N_24988,N_24889);
or UO_42 (O_42,N_24975,N_24856);
nand UO_43 (O_43,N_24908,N_24976);
nor UO_44 (O_44,N_24947,N_24996);
or UO_45 (O_45,N_24926,N_24960);
and UO_46 (O_46,N_24933,N_24989);
nand UO_47 (O_47,N_24992,N_24862);
or UO_48 (O_48,N_24821,N_24834);
nor UO_49 (O_49,N_24997,N_24883);
or UO_50 (O_50,N_24904,N_24859);
nor UO_51 (O_51,N_24993,N_24944);
nand UO_52 (O_52,N_24851,N_24951);
or UO_53 (O_53,N_24837,N_24953);
nand UO_54 (O_54,N_24914,N_24841);
nand UO_55 (O_55,N_24936,N_24825);
or UO_56 (O_56,N_24984,N_24839);
and UO_57 (O_57,N_24886,N_24943);
and UO_58 (O_58,N_24887,N_24820);
or UO_59 (O_59,N_24964,N_24814);
and UO_60 (O_60,N_24844,N_24840);
nor UO_61 (O_61,N_24972,N_24929);
and UO_62 (O_62,N_24807,N_24983);
nand UO_63 (O_63,N_24819,N_24917);
or UO_64 (O_64,N_24981,N_24891);
and UO_65 (O_65,N_24970,N_24831);
nand UO_66 (O_66,N_24899,N_24977);
nor UO_67 (O_67,N_24986,N_24860);
nor UO_68 (O_68,N_24861,N_24811);
or UO_69 (O_69,N_24892,N_24901);
nand UO_70 (O_70,N_24815,N_24934);
and UO_71 (O_71,N_24808,N_24982);
nor UO_72 (O_72,N_24900,N_24978);
nand UO_73 (O_73,N_24838,N_24942);
nor UO_74 (O_74,N_24919,N_24827);
xor UO_75 (O_75,N_24963,N_24854);
or UO_76 (O_76,N_24957,N_24801);
and UO_77 (O_77,N_24829,N_24896);
nor UO_78 (O_78,N_24857,N_24845);
nand UO_79 (O_79,N_24847,N_24858);
and UO_80 (O_80,N_24939,N_24868);
nor UO_81 (O_81,N_24888,N_24906);
nand UO_82 (O_82,N_24921,N_24905);
and UO_83 (O_83,N_24833,N_24937);
nor UO_84 (O_84,N_24867,N_24852);
and UO_85 (O_85,N_24897,N_24842);
nand UO_86 (O_86,N_24806,N_24971);
nand UO_87 (O_87,N_24894,N_24938);
nor UO_88 (O_88,N_24956,N_24954);
and UO_89 (O_89,N_24884,N_24955);
and UO_90 (O_90,N_24935,N_24809);
and UO_91 (O_91,N_24853,N_24816);
or UO_92 (O_92,N_24800,N_24893);
nand UO_93 (O_93,N_24877,N_24849);
or UO_94 (O_94,N_24932,N_24803);
and UO_95 (O_95,N_24812,N_24940);
or UO_96 (O_96,N_24922,N_24916);
or UO_97 (O_97,N_24871,N_24873);
nand UO_98 (O_98,N_24830,N_24848);
nand UO_99 (O_99,N_24835,N_24903);
or UO_100 (O_100,N_24927,N_24835);
and UO_101 (O_101,N_24970,N_24931);
nor UO_102 (O_102,N_24837,N_24822);
and UO_103 (O_103,N_24850,N_24822);
and UO_104 (O_104,N_24826,N_24953);
and UO_105 (O_105,N_24926,N_24867);
and UO_106 (O_106,N_24888,N_24850);
and UO_107 (O_107,N_24841,N_24846);
nor UO_108 (O_108,N_24963,N_24838);
nand UO_109 (O_109,N_24900,N_24808);
and UO_110 (O_110,N_24888,N_24932);
and UO_111 (O_111,N_24858,N_24836);
and UO_112 (O_112,N_24832,N_24837);
nor UO_113 (O_113,N_24817,N_24921);
nor UO_114 (O_114,N_24860,N_24980);
and UO_115 (O_115,N_24959,N_24812);
and UO_116 (O_116,N_24968,N_24932);
nor UO_117 (O_117,N_24955,N_24834);
nor UO_118 (O_118,N_24888,N_24986);
nor UO_119 (O_119,N_24918,N_24983);
and UO_120 (O_120,N_24970,N_24802);
nor UO_121 (O_121,N_24932,N_24805);
nand UO_122 (O_122,N_24904,N_24867);
or UO_123 (O_123,N_24994,N_24842);
nor UO_124 (O_124,N_24888,N_24882);
or UO_125 (O_125,N_24904,N_24820);
and UO_126 (O_126,N_24957,N_24839);
or UO_127 (O_127,N_24965,N_24820);
and UO_128 (O_128,N_24858,N_24912);
nor UO_129 (O_129,N_24836,N_24849);
nand UO_130 (O_130,N_24989,N_24883);
and UO_131 (O_131,N_24900,N_24996);
nor UO_132 (O_132,N_24804,N_24947);
nand UO_133 (O_133,N_24907,N_24845);
nor UO_134 (O_134,N_24970,N_24958);
or UO_135 (O_135,N_24875,N_24898);
nand UO_136 (O_136,N_24825,N_24839);
or UO_137 (O_137,N_24988,N_24981);
nor UO_138 (O_138,N_24931,N_24880);
nand UO_139 (O_139,N_24959,N_24913);
nor UO_140 (O_140,N_24991,N_24913);
or UO_141 (O_141,N_24949,N_24963);
nand UO_142 (O_142,N_24919,N_24917);
or UO_143 (O_143,N_24833,N_24987);
nand UO_144 (O_144,N_24962,N_24893);
nor UO_145 (O_145,N_24893,N_24841);
and UO_146 (O_146,N_24811,N_24911);
nand UO_147 (O_147,N_24864,N_24943);
and UO_148 (O_148,N_24846,N_24873);
or UO_149 (O_149,N_24963,N_24910);
and UO_150 (O_150,N_24961,N_24837);
and UO_151 (O_151,N_24963,N_24973);
nor UO_152 (O_152,N_24948,N_24970);
nand UO_153 (O_153,N_24979,N_24986);
or UO_154 (O_154,N_24884,N_24810);
nor UO_155 (O_155,N_24853,N_24963);
nand UO_156 (O_156,N_24849,N_24869);
nand UO_157 (O_157,N_24975,N_24938);
nor UO_158 (O_158,N_24847,N_24904);
nand UO_159 (O_159,N_24950,N_24991);
and UO_160 (O_160,N_24840,N_24945);
nand UO_161 (O_161,N_24996,N_24834);
nand UO_162 (O_162,N_24861,N_24844);
or UO_163 (O_163,N_24919,N_24889);
nand UO_164 (O_164,N_24918,N_24903);
and UO_165 (O_165,N_24949,N_24957);
or UO_166 (O_166,N_24902,N_24885);
or UO_167 (O_167,N_24862,N_24939);
and UO_168 (O_168,N_24908,N_24834);
or UO_169 (O_169,N_24988,N_24958);
nand UO_170 (O_170,N_24982,N_24968);
nand UO_171 (O_171,N_24850,N_24885);
or UO_172 (O_172,N_24801,N_24964);
and UO_173 (O_173,N_24991,N_24867);
and UO_174 (O_174,N_24972,N_24809);
nand UO_175 (O_175,N_24969,N_24867);
nor UO_176 (O_176,N_24874,N_24806);
nor UO_177 (O_177,N_24824,N_24958);
and UO_178 (O_178,N_24908,N_24860);
nand UO_179 (O_179,N_24993,N_24979);
nand UO_180 (O_180,N_24863,N_24915);
nor UO_181 (O_181,N_24815,N_24877);
or UO_182 (O_182,N_24858,N_24937);
nor UO_183 (O_183,N_24806,N_24929);
nand UO_184 (O_184,N_24945,N_24886);
and UO_185 (O_185,N_24993,N_24965);
and UO_186 (O_186,N_24984,N_24948);
or UO_187 (O_187,N_24871,N_24991);
and UO_188 (O_188,N_24800,N_24881);
nand UO_189 (O_189,N_24864,N_24979);
nand UO_190 (O_190,N_24926,N_24929);
nand UO_191 (O_191,N_24822,N_24915);
nor UO_192 (O_192,N_24946,N_24866);
or UO_193 (O_193,N_24886,N_24835);
and UO_194 (O_194,N_24949,N_24867);
and UO_195 (O_195,N_24938,N_24820);
and UO_196 (O_196,N_24986,N_24848);
nor UO_197 (O_197,N_24989,N_24861);
or UO_198 (O_198,N_24972,N_24941);
and UO_199 (O_199,N_24806,N_24816);
nand UO_200 (O_200,N_24853,N_24980);
or UO_201 (O_201,N_24893,N_24969);
nor UO_202 (O_202,N_24947,N_24944);
nor UO_203 (O_203,N_24949,N_24891);
nand UO_204 (O_204,N_24845,N_24849);
or UO_205 (O_205,N_24868,N_24852);
and UO_206 (O_206,N_24800,N_24806);
xnor UO_207 (O_207,N_24981,N_24873);
and UO_208 (O_208,N_24885,N_24813);
nand UO_209 (O_209,N_24976,N_24819);
nand UO_210 (O_210,N_24892,N_24884);
nand UO_211 (O_211,N_24883,N_24988);
nand UO_212 (O_212,N_24864,N_24813);
nor UO_213 (O_213,N_24826,N_24866);
nor UO_214 (O_214,N_24958,N_24915);
nand UO_215 (O_215,N_24869,N_24909);
nor UO_216 (O_216,N_24838,N_24904);
and UO_217 (O_217,N_24983,N_24846);
or UO_218 (O_218,N_24956,N_24911);
nor UO_219 (O_219,N_24812,N_24983);
nand UO_220 (O_220,N_24860,N_24820);
nand UO_221 (O_221,N_24884,N_24984);
nand UO_222 (O_222,N_24955,N_24963);
or UO_223 (O_223,N_24881,N_24828);
nand UO_224 (O_224,N_24945,N_24838);
nor UO_225 (O_225,N_24810,N_24877);
or UO_226 (O_226,N_24942,N_24862);
or UO_227 (O_227,N_24805,N_24878);
nor UO_228 (O_228,N_24861,N_24968);
nor UO_229 (O_229,N_24935,N_24892);
nand UO_230 (O_230,N_24800,N_24897);
or UO_231 (O_231,N_24827,N_24880);
nor UO_232 (O_232,N_24933,N_24823);
or UO_233 (O_233,N_24928,N_24869);
or UO_234 (O_234,N_24865,N_24973);
nand UO_235 (O_235,N_24838,N_24969);
nor UO_236 (O_236,N_24954,N_24857);
or UO_237 (O_237,N_24876,N_24891);
or UO_238 (O_238,N_24998,N_24888);
nor UO_239 (O_239,N_24970,N_24930);
nor UO_240 (O_240,N_24880,N_24972);
nor UO_241 (O_241,N_24816,N_24964);
nand UO_242 (O_242,N_24821,N_24867);
nor UO_243 (O_243,N_24920,N_24897);
or UO_244 (O_244,N_24902,N_24849);
nand UO_245 (O_245,N_24966,N_24917);
nand UO_246 (O_246,N_24849,N_24933);
nand UO_247 (O_247,N_24964,N_24914);
nand UO_248 (O_248,N_24921,N_24944);
nand UO_249 (O_249,N_24949,N_24865);
nor UO_250 (O_250,N_24881,N_24803);
nor UO_251 (O_251,N_24878,N_24948);
nand UO_252 (O_252,N_24817,N_24944);
xor UO_253 (O_253,N_24823,N_24853);
nand UO_254 (O_254,N_24952,N_24973);
or UO_255 (O_255,N_24905,N_24924);
or UO_256 (O_256,N_24929,N_24990);
and UO_257 (O_257,N_24808,N_24902);
nand UO_258 (O_258,N_24890,N_24818);
nand UO_259 (O_259,N_24953,N_24948);
or UO_260 (O_260,N_24864,N_24988);
nand UO_261 (O_261,N_24978,N_24808);
nand UO_262 (O_262,N_24801,N_24911);
nand UO_263 (O_263,N_24888,N_24810);
nor UO_264 (O_264,N_24800,N_24926);
or UO_265 (O_265,N_24978,N_24888);
nor UO_266 (O_266,N_24940,N_24996);
nand UO_267 (O_267,N_24813,N_24922);
or UO_268 (O_268,N_24932,N_24905);
nor UO_269 (O_269,N_24840,N_24964);
nor UO_270 (O_270,N_24977,N_24970);
nand UO_271 (O_271,N_24989,N_24970);
or UO_272 (O_272,N_24850,N_24837);
nor UO_273 (O_273,N_24894,N_24968);
nand UO_274 (O_274,N_24964,N_24948);
and UO_275 (O_275,N_24901,N_24826);
and UO_276 (O_276,N_24942,N_24940);
nand UO_277 (O_277,N_24894,N_24839);
and UO_278 (O_278,N_24860,N_24926);
or UO_279 (O_279,N_24827,N_24866);
or UO_280 (O_280,N_24908,N_24897);
nand UO_281 (O_281,N_24950,N_24845);
nor UO_282 (O_282,N_24948,N_24820);
or UO_283 (O_283,N_24925,N_24932);
or UO_284 (O_284,N_24884,N_24812);
or UO_285 (O_285,N_24878,N_24801);
nand UO_286 (O_286,N_24881,N_24812);
nor UO_287 (O_287,N_24985,N_24863);
nand UO_288 (O_288,N_24970,N_24848);
nor UO_289 (O_289,N_24982,N_24992);
and UO_290 (O_290,N_24958,N_24880);
or UO_291 (O_291,N_24900,N_24990);
or UO_292 (O_292,N_24912,N_24965);
or UO_293 (O_293,N_24903,N_24815);
and UO_294 (O_294,N_24881,N_24908);
or UO_295 (O_295,N_24861,N_24906);
and UO_296 (O_296,N_24820,N_24987);
and UO_297 (O_297,N_24900,N_24849);
nand UO_298 (O_298,N_24851,N_24901);
nor UO_299 (O_299,N_24989,N_24900);
nor UO_300 (O_300,N_24949,N_24805);
xor UO_301 (O_301,N_24852,N_24847);
nand UO_302 (O_302,N_24895,N_24872);
or UO_303 (O_303,N_24944,N_24914);
or UO_304 (O_304,N_24917,N_24884);
and UO_305 (O_305,N_24913,N_24857);
nand UO_306 (O_306,N_24865,N_24915);
or UO_307 (O_307,N_24842,N_24974);
or UO_308 (O_308,N_24843,N_24858);
or UO_309 (O_309,N_24930,N_24865);
nor UO_310 (O_310,N_24827,N_24868);
and UO_311 (O_311,N_24963,N_24830);
and UO_312 (O_312,N_24927,N_24930);
nor UO_313 (O_313,N_24810,N_24954);
or UO_314 (O_314,N_24903,N_24826);
xnor UO_315 (O_315,N_24962,N_24832);
nor UO_316 (O_316,N_24962,N_24895);
or UO_317 (O_317,N_24885,N_24869);
nor UO_318 (O_318,N_24917,N_24867);
or UO_319 (O_319,N_24907,N_24864);
or UO_320 (O_320,N_24822,N_24813);
and UO_321 (O_321,N_24973,N_24811);
nor UO_322 (O_322,N_24958,N_24900);
or UO_323 (O_323,N_24970,N_24950);
nand UO_324 (O_324,N_24958,N_24837);
nor UO_325 (O_325,N_24943,N_24999);
nand UO_326 (O_326,N_24868,N_24913);
and UO_327 (O_327,N_24972,N_24903);
nor UO_328 (O_328,N_24806,N_24928);
or UO_329 (O_329,N_24801,N_24982);
nand UO_330 (O_330,N_24819,N_24860);
nor UO_331 (O_331,N_24901,N_24978);
or UO_332 (O_332,N_24842,N_24891);
nand UO_333 (O_333,N_24856,N_24903);
or UO_334 (O_334,N_24807,N_24893);
nand UO_335 (O_335,N_24999,N_24908);
nor UO_336 (O_336,N_24988,N_24994);
and UO_337 (O_337,N_24970,N_24809);
and UO_338 (O_338,N_24960,N_24832);
and UO_339 (O_339,N_24947,N_24964);
nand UO_340 (O_340,N_24850,N_24874);
and UO_341 (O_341,N_24929,N_24988);
nor UO_342 (O_342,N_24957,N_24987);
or UO_343 (O_343,N_24842,N_24860);
nor UO_344 (O_344,N_24963,N_24831);
and UO_345 (O_345,N_24933,N_24886);
or UO_346 (O_346,N_24820,N_24934);
and UO_347 (O_347,N_24802,N_24994);
nor UO_348 (O_348,N_24966,N_24859);
nand UO_349 (O_349,N_24808,N_24864);
and UO_350 (O_350,N_24845,N_24901);
or UO_351 (O_351,N_24850,N_24938);
nor UO_352 (O_352,N_24916,N_24933);
nand UO_353 (O_353,N_24969,N_24810);
nor UO_354 (O_354,N_24900,N_24829);
or UO_355 (O_355,N_24860,N_24987);
or UO_356 (O_356,N_24864,N_24931);
nor UO_357 (O_357,N_24929,N_24823);
or UO_358 (O_358,N_24974,N_24935);
and UO_359 (O_359,N_24936,N_24873);
nand UO_360 (O_360,N_24945,N_24990);
or UO_361 (O_361,N_24879,N_24859);
or UO_362 (O_362,N_24958,N_24916);
and UO_363 (O_363,N_24905,N_24941);
or UO_364 (O_364,N_24930,N_24802);
or UO_365 (O_365,N_24973,N_24966);
nand UO_366 (O_366,N_24921,N_24883);
and UO_367 (O_367,N_24974,N_24955);
nor UO_368 (O_368,N_24972,N_24890);
or UO_369 (O_369,N_24853,N_24804);
and UO_370 (O_370,N_24904,N_24879);
or UO_371 (O_371,N_24847,N_24834);
or UO_372 (O_372,N_24902,N_24856);
or UO_373 (O_373,N_24851,N_24931);
nor UO_374 (O_374,N_24888,N_24875);
nand UO_375 (O_375,N_24835,N_24937);
or UO_376 (O_376,N_24970,N_24916);
and UO_377 (O_377,N_24800,N_24994);
or UO_378 (O_378,N_24871,N_24865);
and UO_379 (O_379,N_24873,N_24985);
and UO_380 (O_380,N_24945,N_24943);
or UO_381 (O_381,N_24928,N_24879);
and UO_382 (O_382,N_24816,N_24962);
or UO_383 (O_383,N_24867,N_24921);
nor UO_384 (O_384,N_24885,N_24922);
nand UO_385 (O_385,N_24933,N_24936);
and UO_386 (O_386,N_24935,N_24877);
and UO_387 (O_387,N_24849,N_24807);
and UO_388 (O_388,N_24982,N_24990);
or UO_389 (O_389,N_24970,N_24917);
or UO_390 (O_390,N_24887,N_24953);
and UO_391 (O_391,N_24904,N_24921);
or UO_392 (O_392,N_24914,N_24809);
and UO_393 (O_393,N_24888,N_24969);
nor UO_394 (O_394,N_24860,N_24834);
or UO_395 (O_395,N_24817,N_24975);
nor UO_396 (O_396,N_24993,N_24960);
nor UO_397 (O_397,N_24818,N_24877);
or UO_398 (O_398,N_24919,N_24911);
and UO_399 (O_399,N_24837,N_24903);
or UO_400 (O_400,N_24901,N_24848);
and UO_401 (O_401,N_24800,N_24896);
nor UO_402 (O_402,N_24952,N_24868);
nor UO_403 (O_403,N_24809,N_24801);
nand UO_404 (O_404,N_24910,N_24923);
nor UO_405 (O_405,N_24938,N_24841);
nor UO_406 (O_406,N_24979,N_24931);
nand UO_407 (O_407,N_24995,N_24907);
and UO_408 (O_408,N_24968,N_24846);
and UO_409 (O_409,N_24954,N_24888);
nor UO_410 (O_410,N_24929,N_24899);
or UO_411 (O_411,N_24949,N_24855);
or UO_412 (O_412,N_24999,N_24975);
nand UO_413 (O_413,N_24878,N_24821);
and UO_414 (O_414,N_24845,N_24938);
or UO_415 (O_415,N_24807,N_24984);
and UO_416 (O_416,N_24999,N_24890);
and UO_417 (O_417,N_24887,N_24891);
or UO_418 (O_418,N_24938,N_24960);
or UO_419 (O_419,N_24866,N_24847);
or UO_420 (O_420,N_24862,N_24967);
nor UO_421 (O_421,N_24804,N_24883);
nor UO_422 (O_422,N_24891,N_24810);
and UO_423 (O_423,N_24884,N_24887);
xnor UO_424 (O_424,N_24987,N_24924);
xnor UO_425 (O_425,N_24852,N_24828);
and UO_426 (O_426,N_24906,N_24820);
nor UO_427 (O_427,N_24818,N_24883);
and UO_428 (O_428,N_24823,N_24872);
and UO_429 (O_429,N_24918,N_24945);
or UO_430 (O_430,N_24805,N_24942);
nor UO_431 (O_431,N_24995,N_24988);
or UO_432 (O_432,N_24954,N_24968);
and UO_433 (O_433,N_24811,N_24951);
and UO_434 (O_434,N_24985,N_24996);
and UO_435 (O_435,N_24993,N_24840);
or UO_436 (O_436,N_24853,N_24835);
nand UO_437 (O_437,N_24962,N_24966);
nor UO_438 (O_438,N_24948,N_24882);
nand UO_439 (O_439,N_24833,N_24827);
nand UO_440 (O_440,N_24969,N_24971);
and UO_441 (O_441,N_24924,N_24849);
or UO_442 (O_442,N_24930,N_24859);
nor UO_443 (O_443,N_24814,N_24935);
or UO_444 (O_444,N_24845,N_24931);
nand UO_445 (O_445,N_24968,N_24803);
nand UO_446 (O_446,N_24812,N_24831);
nand UO_447 (O_447,N_24812,N_24920);
xnor UO_448 (O_448,N_24915,N_24808);
nor UO_449 (O_449,N_24896,N_24835);
nand UO_450 (O_450,N_24976,N_24893);
nand UO_451 (O_451,N_24825,N_24935);
nand UO_452 (O_452,N_24996,N_24895);
nand UO_453 (O_453,N_24993,N_24948);
and UO_454 (O_454,N_24819,N_24808);
nor UO_455 (O_455,N_24950,N_24978);
nor UO_456 (O_456,N_24814,N_24832);
and UO_457 (O_457,N_24845,N_24804);
xor UO_458 (O_458,N_24851,N_24954);
and UO_459 (O_459,N_24907,N_24905);
nand UO_460 (O_460,N_24859,N_24938);
nor UO_461 (O_461,N_24820,N_24841);
or UO_462 (O_462,N_24944,N_24813);
nor UO_463 (O_463,N_24890,N_24974);
or UO_464 (O_464,N_24868,N_24930);
nand UO_465 (O_465,N_24889,N_24968);
or UO_466 (O_466,N_24943,N_24879);
or UO_467 (O_467,N_24810,N_24881);
nor UO_468 (O_468,N_24805,N_24811);
nand UO_469 (O_469,N_24846,N_24827);
nor UO_470 (O_470,N_24942,N_24809);
or UO_471 (O_471,N_24934,N_24955);
and UO_472 (O_472,N_24926,N_24966);
and UO_473 (O_473,N_24925,N_24997);
and UO_474 (O_474,N_24976,N_24925);
nand UO_475 (O_475,N_24836,N_24965);
nor UO_476 (O_476,N_24969,N_24837);
and UO_477 (O_477,N_24838,N_24916);
or UO_478 (O_478,N_24835,N_24998);
and UO_479 (O_479,N_24943,N_24894);
nand UO_480 (O_480,N_24837,N_24876);
and UO_481 (O_481,N_24827,N_24858);
nand UO_482 (O_482,N_24991,N_24806);
and UO_483 (O_483,N_24951,N_24943);
nor UO_484 (O_484,N_24991,N_24949);
nand UO_485 (O_485,N_24945,N_24893);
nand UO_486 (O_486,N_24917,N_24920);
nand UO_487 (O_487,N_24909,N_24955);
nor UO_488 (O_488,N_24819,N_24940);
nand UO_489 (O_489,N_24942,N_24826);
or UO_490 (O_490,N_24878,N_24852);
and UO_491 (O_491,N_24914,N_24830);
or UO_492 (O_492,N_24952,N_24859);
nor UO_493 (O_493,N_24897,N_24953);
xnor UO_494 (O_494,N_24909,N_24980);
nand UO_495 (O_495,N_24850,N_24952);
nand UO_496 (O_496,N_24826,N_24874);
nor UO_497 (O_497,N_24863,N_24924);
nor UO_498 (O_498,N_24862,N_24830);
and UO_499 (O_499,N_24887,N_24922);
or UO_500 (O_500,N_24997,N_24944);
nor UO_501 (O_501,N_24887,N_24920);
nor UO_502 (O_502,N_24977,N_24939);
and UO_503 (O_503,N_24987,N_24965);
nand UO_504 (O_504,N_24918,N_24897);
or UO_505 (O_505,N_24826,N_24949);
or UO_506 (O_506,N_24885,N_24990);
or UO_507 (O_507,N_24854,N_24898);
nand UO_508 (O_508,N_24831,N_24968);
nand UO_509 (O_509,N_24861,N_24953);
and UO_510 (O_510,N_24939,N_24981);
xor UO_511 (O_511,N_24990,N_24912);
nand UO_512 (O_512,N_24938,N_24979);
nand UO_513 (O_513,N_24888,N_24941);
nand UO_514 (O_514,N_24893,N_24809);
nand UO_515 (O_515,N_24988,N_24916);
or UO_516 (O_516,N_24874,N_24899);
and UO_517 (O_517,N_24957,N_24808);
or UO_518 (O_518,N_24830,N_24973);
nand UO_519 (O_519,N_24896,N_24885);
or UO_520 (O_520,N_24993,N_24848);
and UO_521 (O_521,N_24864,N_24903);
nor UO_522 (O_522,N_24808,N_24913);
or UO_523 (O_523,N_24966,N_24980);
nor UO_524 (O_524,N_24836,N_24961);
nor UO_525 (O_525,N_24871,N_24898);
and UO_526 (O_526,N_24907,N_24964);
nand UO_527 (O_527,N_24885,N_24951);
nor UO_528 (O_528,N_24822,N_24873);
and UO_529 (O_529,N_24967,N_24876);
nand UO_530 (O_530,N_24874,N_24872);
and UO_531 (O_531,N_24907,N_24847);
nor UO_532 (O_532,N_24804,N_24914);
or UO_533 (O_533,N_24840,N_24904);
and UO_534 (O_534,N_24991,N_24832);
nand UO_535 (O_535,N_24834,N_24867);
and UO_536 (O_536,N_24953,N_24986);
nor UO_537 (O_537,N_24801,N_24855);
nor UO_538 (O_538,N_24931,N_24923);
and UO_539 (O_539,N_24855,N_24894);
nand UO_540 (O_540,N_24813,N_24963);
nand UO_541 (O_541,N_24953,N_24995);
nand UO_542 (O_542,N_24818,N_24852);
and UO_543 (O_543,N_24871,N_24880);
nor UO_544 (O_544,N_24891,N_24967);
nand UO_545 (O_545,N_24852,N_24805);
nand UO_546 (O_546,N_24820,N_24856);
nand UO_547 (O_547,N_24832,N_24876);
nand UO_548 (O_548,N_24897,N_24843);
or UO_549 (O_549,N_24993,N_24845);
nand UO_550 (O_550,N_24996,N_24968);
or UO_551 (O_551,N_24870,N_24978);
or UO_552 (O_552,N_24877,N_24873);
nand UO_553 (O_553,N_24867,N_24888);
or UO_554 (O_554,N_24881,N_24900);
and UO_555 (O_555,N_24914,N_24816);
and UO_556 (O_556,N_24997,N_24950);
nor UO_557 (O_557,N_24821,N_24963);
and UO_558 (O_558,N_24949,N_24827);
and UO_559 (O_559,N_24999,N_24892);
and UO_560 (O_560,N_24874,N_24904);
nand UO_561 (O_561,N_24957,N_24803);
nand UO_562 (O_562,N_24966,N_24982);
or UO_563 (O_563,N_24860,N_24972);
nor UO_564 (O_564,N_24991,N_24822);
nor UO_565 (O_565,N_24999,N_24995);
or UO_566 (O_566,N_24995,N_24857);
and UO_567 (O_567,N_24882,N_24945);
nand UO_568 (O_568,N_24995,N_24830);
or UO_569 (O_569,N_24834,N_24972);
nand UO_570 (O_570,N_24978,N_24885);
xor UO_571 (O_571,N_24904,N_24932);
nand UO_572 (O_572,N_24809,N_24834);
or UO_573 (O_573,N_24857,N_24963);
nand UO_574 (O_574,N_24911,N_24853);
xnor UO_575 (O_575,N_24958,N_24845);
nor UO_576 (O_576,N_24878,N_24884);
and UO_577 (O_577,N_24811,N_24945);
nand UO_578 (O_578,N_24985,N_24834);
and UO_579 (O_579,N_24840,N_24924);
and UO_580 (O_580,N_24844,N_24822);
nand UO_581 (O_581,N_24808,N_24868);
nand UO_582 (O_582,N_24886,N_24801);
nand UO_583 (O_583,N_24962,N_24849);
and UO_584 (O_584,N_24889,N_24853);
and UO_585 (O_585,N_24884,N_24965);
nand UO_586 (O_586,N_24944,N_24806);
or UO_587 (O_587,N_24833,N_24907);
nor UO_588 (O_588,N_24931,N_24862);
nand UO_589 (O_589,N_24923,N_24987);
nor UO_590 (O_590,N_24922,N_24886);
and UO_591 (O_591,N_24982,N_24850);
or UO_592 (O_592,N_24817,N_24961);
or UO_593 (O_593,N_24826,N_24876);
nor UO_594 (O_594,N_24940,N_24900);
nand UO_595 (O_595,N_24846,N_24812);
or UO_596 (O_596,N_24986,N_24938);
nand UO_597 (O_597,N_24920,N_24904);
nor UO_598 (O_598,N_24846,N_24918);
nand UO_599 (O_599,N_24928,N_24993);
nor UO_600 (O_600,N_24907,N_24953);
or UO_601 (O_601,N_24842,N_24800);
nand UO_602 (O_602,N_24853,N_24998);
or UO_603 (O_603,N_24900,N_24896);
or UO_604 (O_604,N_24936,N_24885);
nand UO_605 (O_605,N_24876,N_24845);
and UO_606 (O_606,N_24955,N_24855);
nor UO_607 (O_607,N_24824,N_24905);
and UO_608 (O_608,N_24808,N_24994);
or UO_609 (O_609,N_24996,N_24804);
nand UO_610 (O_610,N_24846,N_24952);
or UO_611 (O_611,N_24847,N_24863);
nor UO_612 (O_612,N_24876,N_24860);
or UO_613 (O_613,N_24907,N_24858);
nor UO_614 (O_614,N_24804,N_24961);
nand UO_615 (O_615,N_24931,N_24890);
and UO_616 (O_616,N_24956,N_24915);
nor UO_617 (O_617,N_24979,N_24921);
nor UO_618 (O_618,N_24978,N_24993);
xor UO_619 (O_619,N_24930,N_24964);
and UO_620 (O_620,N_24843,N_24903);
xnor UO_621 (O_621,N_24883,N_24839);
nor UO_622 (O_622,N_24994,N_24831);
nand UO_623 (O_623,N_24840,N_24994);
nand UO_624 (O_624,N_24827,N_24905);
and UO_625 (O_625,N_24921,N_24841);
nand UO_626 (O_626,N_24881,N_24964);
and UO_627 (O_627,N_24836,N_24890);
and UO_628 (O_628,N_24822,N_24807);
or UO_629 (O_629,N_24928,N_24830);
and UO_630 (O_630,N_24856,N_24994);
and UO_631 (O_631,N_24815,N_24823);
or UO_632 (O_632,N_24955,N_24835);
nor UO_633 (O_633,N_24985,N_24822);
nor UO_634 (O_634,N_24927,N_24879);
or UO_635 (O_635,N_24924,N_24992);
nand UO_636 (O_636,N_24895,N_24854);
and UO_637 (O_637,N_24961,N_24907);
nor UO_638 (O_638,N_24958,N_24812);
or UO_639 (O_639,N_24807,N_24958);
nand UO_640 (O_640,N_24917,N_24902);
nand UO_641 (O_641,N_24982,N_24999);
and UO_642 (O_642,N_24856,N_24924);
and UO_643 (O_643,N_24877,N_24943);
and UO_644 (O_644,N_24851,N_24948);
nand UO_645 (O_645,N_24912,N_24896);
nor UO_646 (O_646,N_24947,N_24974);
and UO_647 (O_647,N_24959,N_24988);
nand UO_648 (O_648,N_24957,N_24841);
nand UO_649 (O_649,N_24940,N_24896);
nor UO_650 (O_650,N_24991,N_24842);
and UO_651 (O_651,N_24875,N_24927);
or UO_652 (O_652,N_24815,N_24884);
nand UO_653 (O_653,N_24812,N_24945);
nor UO_654 (O_654,N_24914,N_24833);
nor UO_655 (O_655,N_24972,N_24915);
or UO_656 (O_656,N_24811,N_24967);
and UO_657 (O_657,N_24872,N_24984);
or UO_658 (O_658,N_24818,N_24859);
and UO_659 (O_659,N_24998,N_24893);
nand UO_660 (O_660,N_24992,N_24881);
nor UO_661 (O_661,N_24970,N_24915);
and UO_662 (O_662,N_24813,N_24995);
nor UO_663 (O_663,N_24922,N_24935);
nor UO_664 (O_664,N_24868,N_24985);
nand UO_665 (O_665,N_24826,N_24803);
nand UO_666 (O_666,N_24969,N_24805);
or UO_667 (O_667,N_24991,N_24804);
or UO_668 (O_668,N_24911,N_24957);
and UO_669 (O_669,N_24914,N_24815);
and UO_670 (O_670,N_24880,N_24967);
and UO_671 (O_671,N_24807,N_24808);
or UO_672 (O_672,N_24904,N_24842);
and UO_673 (O_673,N_24989,N_24878);
nor UO_674 (O_674,N_24889,N_24993);
or UO_675 (O_675,N_24847,N_24897);
nor UO_676 (O_676,N_24934,N_24960);
nor UO_677 (O_677,N_24858,N_24909);
nand UO_678 (O_678,N_24955,N_24806);
nand UO_679 (O_679,N_24891,N_24862);
or UO_680 (O_680,N_24962,N_24980);
nand UO_681 (O_681,N_24955,N_24973);
nor UO_682 (O_682,N_24831,N_24961);
or UO_683 (O_683,N_24976,N_24851);
and UO_684 (O_684,N_24969,N_24902);
or UO_685 (O_685,N_24952,N_24986);
and UO_686 (O_686,N_24984,N_24906);
nor UO_687 (O_687,N_24824,N_24836);
nor UO_688 (O_688,N_24956,N_24818);
or UO_689 (O_689,N_24830,N_24950);
nand UO_690 (O_690,N_24852,N_24840);
nand UO_691 (O_691,N_24927,N_24968);
and UO_692 (O_692,N_24827,N_24860);
nor UO_693 (O_693,N_24801,N_24814);
and UO_694 (O_694,N_24880,N_24830);
or UO_695 (O_695,N_24972,N_24969);
and UO_696 (O_696,N_24844,N_24809);
nand UO_697 (O_697,N_24871,N_24842);
and UO_698 (O_698,N_24938,N_24970);
and UO_699 (O_699,N_24877,N_24866);
or UO_700 (O_700,N_24935,N_24815);
or UO_701 (O_701,N_24821,N_24889);
nand UO_702 (O_702,N_24821,N_24829);
or UO_703 (O_703,N_24863,N_24842);
and UO_704 (O_704,N_24942,N_24917);
and UO_705 (O_705,N_24991,N_24966);
and UO_706 (O_706,N_24908,N_24867);
or UO_707 (O_707,N_24837,N_24918);
nor UO_708 (O_708,N_24822,N_24949);
and UO_709 (O_709,N_24877,N_24970);
nor UO_710 (O_710,N_24895,N_24848);
nand UO_711 (O_711,N_24913,N_24978);
nand UO_712 (O_712,N_24933,N_24911);
and UO_713 (O_713,N_24846,N_24924);
nand UO_714 (O_714,N_24988,N_24848);
nor UO_715 (O_715,N_24894,N_24901);
or UO_716 (O_716,N_24942,N_24976);
nand UO_717 (O_717,N_24804,N_24827);
or UO_718 (O_718,N_24919,N_24985);
or UO_719 (O_719,N_24864,N_24953);
nand UO_720 (O_720,N_24955,N_24862);
and UO_721 (O_721,N_24944,N_24842);
nor UO_722 (O_722,N_24837,N_24952);
nand UO_723 (O_723,N_24938,N_24917);
and UO_724 (O_724,N_24902,N_24819);
nand UO_725 (O_725,N_24975,N_24979);
nand UO_726 (O_726,N_24854,N_24850);
nor UO_727 (O_727,N_24957,N_24929);
nor UO_728 (O_728,N_24872,N_24936);
and UO_729 (O_729,N_24920,N_24870);
and UO_730 (O_730,N_24858,N_24957);
or UO_731 (O_731,N_24887,N_24810);
xor UO_732 (O_732,N_24840,N_24957);
and UO_733 (O_733,N_24928,N_24917);
and UO_734 (O_734,N_24816,N_24866);
nand UO_735 (O_735,N_24822,N_24954);
nor UO_736 (O_736,N_24884,N_24959);
nand UO_737 (O_737,N_24943,N_24870);
nand UO_738 (O_738,N_24921,N_24909);
nor UO_739 (O_739,N_24933,N_24964);
nand UO_740 (O_740,N_24879,N_24954);
nor UO_741 (O_741,N_24948,N_24822);
nand UO_742 (O_742,N_24976,N_24927);
or UO_743 (O_743,N_24973,N_24924);
nor UO_744 (O_744,N_24805,N_24999);
and UO_745 (O_745,N_24935,N_24882);
nand UO_746 (O_746,N_24870,N_24955);
or UO_747 (O_747,N_24891,N_24955);
and UO_748 (O_748,N_24885,N_24912);
or UO_749 (O_749,N_24888,N_24975);
and UO_750 (O_750,N_24982,N_24917);
nand UO_751 (O_751,N_24959,N_24957);
nand UO_752 (O_752,N_24806,N_24895);
nor UO_753 (O_753,N_24954,N_24824);
and UO_754 (O_754,N_24872,N_24920);
nor UO_755 (O_755,N_24977,N_24826);
nor UO_756 (O_756,N_24931,N_24980);
and UO_757 (O_757,N_24978,N_24840);
and UO_758 (O_758,N_24835,N_24985);
and UO_759 (O_759,N_24809,N_24800);
and UO_760 (O_760,N_24983,N_24811);
nand UO_761 (O_761,N_24894,N_24922);
or UO_762 (O_762,N_24977,N_24851);
or UO_763 (O_763,N_24805,N_24849);
nand UO_764 (O_764,N_24806,N_24986);
and UO_765 (O_765,N_24841,N_24951);
or UO_766 (O_766,N_24974,N_24994);
and UO_767 (O_767,N_24971,N_24861);
nor UO_768 (O_768,N_24874,N_24883);
or UO_769 (O_769,N_24804,N_24806);
and UO_770 (O_770,N_24928,N_24805);
nand UO_771 (O_771,N_24903,N_24887);
nand UO_772 (O_772,N_24924,N_24891);
and UO_773 (O_773,N_24853,N_24933);
nor UO_774 (O_774,N_24907,N_24826);
nand UO_775 (O_775,N_24940,N_24851);
nand UO_776 (O_776,N_24911,N_24880);
nor UO_777 (O_777,N_24815,N_24889);
or UO_778 (O_778,N_24851,N_24939);
nor UO_779 (O_779,N_24908,N_24951);
nor UO_780 (O_780,N_24806,N_24919);
nor UO_781 (O_781,N_24908,N_24984);
and UO_782 (O_782,N_24912,N_24817);
nor UO_783 (O_783,N_24914,N_24915);
nand UO_784 (O_784,N_24831,N_24949);
nor UO_785 (O_785,N_24917,N_24990);
nor UO_786 (O_786,N_24880,N_24981);
or UO_787 (O_787,N_24877,N_24853);
and UO_788 (O_788,N_24946,N_24964);
and UO_789 (O_789,N_24971,N_24908);
and UO_790 (O_790,N_24953,N_24919);
nand UO_791 (O_791,N_24927,N_24895);
nor UO_792 (O_792,N_24964,N_24896);
and UO_793 (O_793,N_24974,N_24920);
nor UO_794 (O_794,N_24928,N_24839);
and UO_795 (O_795,N_24876,N_24994);
or UO_796 (O_796,N_24980,N_24811);
or UO_797 (O_797,N_24943,N_24818);
nor UO_798 (O_798,N_24998,N_24899);
nor UO_799 (O_799,N_24976,N_24932);
and UO_800 (O_800,N_24858,N_24825);
nand UO_801 (O_801,N_24880,N_24842);
nor UO_802 (O_802,N_24974,N_24834);
and UO_803 (O_803,N_24966,N_24943);
and UO_804 (O_804,N_24892,N_24827);
nor UO_805 (O_805,N_24942,N_24908);
and UO_806 (O_806,N_24885,N_24825);
nor UO_807 (O_807,N_24813,N_24909);
nand UO_808 (O_808,N_24802,N_24881);
or UO_809 (O_809,N_24973,N_24841);
nor UO_810 (O_810,N_24948,N_24922);
nor UO_811 (O_811,N_24959,N_24830);
or UO_812 (O_812,N_24834,N_24827);
nor UO_813 (O_813,N_24981,N_24911);
nand UO_814 (O_814,N_24915,N_24929);
nor UO_815 (O_815,N_24952,N_24845);
nor UO_816 (O_816,N_24918,N_24896);
and UO_817 (O_817,N_24959,N_24869);
and UO_818 (O_818,N_24951,N_24984);
or UO_819 (O_819,N_24974,N_24900);
nor UO_820 (O_820,N_24857,N_24818);
nor UO_821 (O_821,N_24846,N_24836);
nand UO_822 (O_822,N_24915,N_24885);
nor UO_823 (O_823,N_24952,N_24831);
or UO_824 (O_824,N_24838,N_24892);
and UO_825 (O_825,N_24967,N_24808);
nor UO_826 (O_826,N_24994,N_24852);
and UO_827 (O_827,N_24963,N_24880);
and UO_828 (O_828,N_24969,N_24956);
and UO_829 (O_829,N_24940,N_24915);
nor UO_830 (O_830,N_24998,N_24966);
and UO_831 (O_831,N_24811,N_24814);
nor UO_832 (O_832,N_24869,N_24815);
and UO_833 (O_833,N_24849,N_24811);
and UO_834 (O_834,N_24934,N_24881);
or UO_835 (O_835,N_24965,N_24953);
nand UO_836 (O_836,N_24953,N_24970);
nor UO_837 (O_837,N_24831,N_24900);
or UO_838 (O_838,N_24840,N_24874);
and UO_839 (O_839,N_24908,N_24843);
nand UO_840 (O_840,N_24846,N_24855);
nand UO_841 (O_841,N_24982,N_24891);
and UO_842 (O_842,N_24862,N_24994);
nor UO_843 (O_843,N_24994,N_24836);
nor UO_844 (O_844,N_24888,N_24995);
and UO_845 (O_845,N_24880,N_24927);
nand UO_846 (O_846,N_24959,N_24936);
nor UO_847 (O_847,N_24884,N_24951);
or UO_848 (O_848,N_24934,N_24813);
or UO_849 (O_849,N_24934,N_24944);
nor UO_850 (O_850,N_24932,N_24846);
and UO_851 (O_851,N_24889,N_24851);
nor UO_852 (O_852,N_24996,N_24837);
or UO_853 (O_853,N_24838,N_24951);
nor UO_854 (O_854,N_24803,N_24812);
nand UO_855 (O_855,N_24819,N_24833);
nand UO_856 (O_856,N_24992,N_24946);
and UO_857 (O_857,N_24947,N_24990);
nor UO_858 (O_858,N_24874,N_24845);
nor UO_859 (O_859,N_24934,N_24918);
or UO_860 (O_860,N_24892,N_24847);
nor UO_861 (O_861,N_24896,N_24999);
and UO_862 (O_862,N_24820,N_24916);
nor UO_863 (O_863,N_24914,N_24912);
or UO_864 (O_864,N_24971,N_24943);
nand UO_865 (O_865,N_24952,N_24953);
and UO_866 (O_866,N_24961,N_24993);
nand UO_867 (O_867,N_24860,N_24945);
nand UO_868 (O_868,N_24975,N_24863);
or UO_869 (O_869,N_24869,N_24829);
or UO_870 (O_870,N_24839,N_24838);
and UO_871 (O_871,N_24806,N_24851);
nor UO_872 (O_872,N_24859,N_24939);
or UO_873 (O_873,N_24948,N_24857);
and UO_874 (O_874,N_24877,N_24920);
nand UO_875 (O_875,N_24994,N_24991);
nand UO_876 (O_876,N_24893,N_24981);
nand UO_877 (O_877,N_24968,N_24903);
or UO_878 (O_878,N_24904,N_24805);
or UO_879 (O_879,N_24908,N_24821);
nand UO_880 (O_880,N_24806,N_24890);
and UO_881 (O_881,N_24913,N_24903);
nand UO_882 (O_882,N_24978,N_24819);
nand UO_883 (O_883,N_24810,N_24880);
and UO_884 (O_884,N_24852,N_24845);
nor UO_885 (O_885,N_24938,N_24889);
nor UO_886 (O_886,N_24905,N_24937);
or UO_887 (O_887,N_24999,N_24984);
xnor UO_888 (O_888,N_24912,N_24898);
or UO_889 (O_889,N_24860,N_24920);
and UO_890 (O_890,N_24911,N_24951);
xnor UO_891 (O_891,N_24977,N_24934);
and UO_892 (O_892,N_24875,N_24999);
nor UO_893 (O_893,N_24805,N_24831);
or UO_894 (O_894,N_24871,N_24995);
xor UO_895 (O_895,N_24958,N_24802);
or UO_896 (O_896,N_24800,N_24959);
nand UO_897 (O_897,N_24907,N_24872);
nor UO_898 (O_898,N_24998,N_24959);
or UO_899 (O_899,N_24938,N_24945);
nand UO_900 (O_900,N_24977,N_24838);
nor UO_901 (O_901,N_24891,N_24855);
and UO_902 (O_902,N_24866,N_24860);
and UO_903 (O_903,N_24991,N_24868);
and UO_904 (O_904,N_24835,N_24861);
nor UO_905 (O_905,N_24914,N_24858);
and UO_906 (O_906,N_24979,N_24852);
and UO_907 (O_907,N_24948,N_24977);
and UO_908 (O_908,N_24976,N_24831);
nand UO_909 (O_909,N_24823,N_24895);
or UO_910 (O_910,N_24801,N_24894);
or UO_911 (O_911,N_24890,N_24832);
nand UO_912 (O_912,N_24841,N_24868);
or UO_913 (O_913,N_24903,N_24999);
nand UO_914 (O_914,N_24964,N_24928);
nor UO_915 (O_915,N_24902,N_24810);
nor UO_916 (O_916,N_24956,N_24873);
nor UO_917 (O_917,N_24951,N_24878);
nor UO_918 (O_918,N_24896,N_24956);
or UO_919 (O_919,N_24967,N_24907);
or UO_920 (O_920,N_24978,N_24903);
and UO_921 (O_921,N_24815,N_24956);
or UO_922 (O_922,N_24992,N_24974);
and UO_923 (O_923,N_24910,N_24874);
nand UO_924 (O_924,N_24909,N_24974);
or UO_925 (O_925,N_24811,N_24933);
or UO_926 (O_926,N_24907,N_24935);
nor UO_927 (O_927,N_24961,N_24930);
and UO_928 (O_928,N_24932,N_24828);
xnor UO_929 (O_929,N_24816,N_24957);
and UO_930 (O_930,N_24839,N_24820);
or UO_931 (O_931,N_24941,N_24979);
or UO_932 (O_932,N_24869,N_24817);
and UO_933 (O_933,N_24858,N_24835);
and UO_934 (O_934,N_24979,N_24880);
nand UO_935 (O_935,N_24921,N_24866);
nand UO_936 (O_936,N_24813,N_24828);
or UO_937 (O_937,N_24836,N_24852);
nand UO_938 (O_938,N_24840,N_24919);
and UO_939 (O_939,N_24815,N_24954);
or UO_940 (O_940,N_24859,N_24850);
nand UO_941 (O_941,N_24996,N_24803);
and UO_942 (O_942,N_24956,N_24882);
nand UO_943 (O_943,N_24852,N_24984);
nor UO_944 (O_944,N_24882,N_24814);
or UO_945 (O_945,N_24911,N_24964);
or UO_946 (O_946,N_24996,N_24881);
or UO_947 (O_947,N_24957,N_24965);
nand UO_948 (O_948,N_24837,N_24931);
or UO_949 (O_949,N_24941,N_24938);
or UO_950 (O_950,N_24819,N_24838);
or UO_951 (O_951,N_24981,N_24829);
nor UO_952 (O_952,N_24925,N_24942);
nor UO_953 (O_953,N_24822,N_24958);
nor UO_954 (O_954,N_24814,N_24886);
or UO_955 (O_955,N_24927,N_24936);
nor UO_956 (O_956,N_24858,N_24991);
nor UO_957 (O_957,N_24997,N_24908);
and UO_958 (O_958,N_24883,N_24992);
and UO_959 (O_959,N_24950,N_24849);
or UO_960 (O_960,N_24950,N_24840);
or UO_961 (O_961,N_24994,N_24815);
and UO_962 (O_962,N_24825,N_24938);
or UO_963 (O_963,N_24895,N_24849);
nand UO_964 (O_964,N_24831,N_24959);
or UO_965 (O_965,N_24879,N_24856);
and UO_966 (O_966,N_24873,N_24802);
nand UO_967 (O_967,N_24842,N_24992);
or UO_968 (O_968,N_24912,N_24829);
nand UO_969 (O_969,N_24892,N_24963);
or UO_970 (O_970,N_24963,N_24847);
nand UO_971 (O_971,N_24963,N_24881);
and UO_972 (O_972,N_24998,N_24815);
nand UO_973 (O_973,N_24965,N_24964);
nand UO_974 (O_974,N_24924,N_24819);
and UO_975 (O_975,N_24930,N_24960);
and UO_976 (O_976,N_24941,N_24991);
nor UO_977 (O_977,N_24917,N_24912);
nand UO_978 (O_978,N_24920,N_24875);
or UO_979 (O_979,N_24857,N_24988);
nand UO_980 (O_980,N_24976,N_24842);
nand UO_981 (O_981,N_24820,N_24903);
and UO_982 (O_982,N_24852,N_24949);
nor UO_983 (O_983,N_24984,N_24853);
and UO_984 (O_984,N_24811,N_24996);
nand UO_985 (O_985,N_24868,N_24918);
nand UO_986 (O_986,N_24896,N_24979);
or UO_987 (O_987,N_24924,N_24860);
and UO_988 (O_988,N_24976,N_24989);
nor UO_989 (O_989,N_24974,N_24984);
nand UO_990 (O_990,N_24845,N_24803);
or UO_991 (O_991,N_24925,N_24999);
nor UO_992 (O_992,N_24972,N_24904);
nor UO_993 (O_993,N_24977,N_24981);
nand UO_994 (O_994,N_24976,N_24850);
nor UO_995 (O_995,N_24848,N_24935);
or UO_996 (O_996,N_24981,N_24933);
or UO_997 (O_997,N_24867,N_24801);
nor UO_998 (O_998,N_24898,N_24903);
or UO_999 (O_999,N_24864,N_24833);
and UO_1000 (O_1000,N_24916,N_24892);
nand UO_1001 (O_1001,N_24947,N_24849);
nand UO_1002 (O_1002,N_24843,N_24930);
nand UO_1003 (O_1003,N_24984,N_24979);
or UO_1004 (O_1004,N_24944,N_24839);
and UO_1005 (O_1005,N_24877,N_24972);
nand UO_1006 (O_1006,N_24820,N_24800);
or UO_1007 (O_1007,N_24978,N_24943);
or UO_1008 (O_1008,N_24889,N_24979);
nor UO_1009 (O_1009,N_24852,N_24917);
and UO_1010 (O_1010,N_24897,N_24980);
and UO_1011 (O_1011,N_24919,N_24943);
nand UO_1012 (O_1012,N_24814,N_24911);
or UO_1013 (O_1013,N_24950,N_24945);
and UO_1014 (O_1014,N_24806,N_24956);
or UO_1015 (O_1015,N_24902,N_24995);
nand UO_1016 (O_1016,N_24818,N_24826);
and UO_1017 (O_1017,N_24955,N_24838);
nand UO_1018 (O_1018,N_24857,N_24984);
nor UO_1019 (O_1019,N_24962,N_24968);
nand UO_1020 (O_1020,N_24836,N_24962);
or UO_1021 (O_1021,N_24896,N_24984);
nand UO_1022 (O_1022,N_24923,N_24825);
nand UO_1023 (O_1023,N_24993,N_24931);
and UO_1024 (O_1024,N_24835,N_24977);
nand UO_1025 (O_1025,N_24988,N_24971);
or UO_1026 (O_1026,N_24900,N_24957);
nand UO_1027 (O_1027,N_24890,N_24810);
nor UO_1028 (O_1028,N_24807,N_24989);
or UO_1029 (O_1029,N_24913,N_24990);
or UO_1030 (O_1030,N_24893,N_24889);
and UO_1031 (O_1031,N_24879,N_24989);
or UO_1032 (O_1032,N_24909,N_24820);
nand UO_1033 (O_1033,N_24800,N_24859);
or UO_1034 (O_1034,N_24802,N_24985);
nand UO_1035 (O_1035,N_24990,N_24970);
and UO_1036 (O_1036,N_24981,N_24899);
nand UO_1037 (O_1037,N_24850,N_24995);
or UO_1038 (O_1038,N_24917,N_24801);
or UO_1039 (O_1039,N_24934,N_24988);
nand UO_1040 (O_1040,N_24887,N_24989);
nor UO_1041 (O_1041,N_24883,N_24854);
nor UO_1042 (O_1042,N_24988,N_24869);
nor UO_1043 (O_1043,N_24814,N_24995);
or UO_1044 (O_1044,N_24909,N_24802);
or UO_1045 (O_1045,N_24814,N_24977);
and UO_1046 (O_1046,N_24835,N_24986);
and UO_1047 (O_1047,N_24964,N_24989);
nor UO_1048 (O_1048,N_24922,N_24954);
nor UO_1049 (O_1049,N_24886,N_24806);
nor UO_1050 (O_1050,N_24958,N_24932);
nor UO_1051 (O_1051,N_24847,N_24896);
nor UO_1052 (O_1052,N_24837,N_24902);
nor UO_1053 (O_1053,N_24950,N_24919);
and UO_1054 (O_1054,N_24915,N_24892);
nor UO_1055 (O_1055,N_24912,N_24899);
nor UO_1056 (O_1056,N_24981,N_24934);
nand UO_1057 (O_1057,N_24896,N_24888);
or UO_1058 (O_1058,N_24913,N_24906);
or UO_1059 (O_1059,N_24881,N_24893);
nor UO_1060 (O_1060,N_24806,N_24941);
nor UO_1061 (O_1061,N_24981,N_24813);
nand UO_1062 (O_1062,N_24834,N_24903);
or UO_1063 (O_1063,N_24967,N_24988);
nor UO_1064 (O_1064,N_24972,N_24957);
nand UO_1065 (O_1065,N_24938,N_24924);
and UO_1066 (O_1066,N_24902,N_24915);
nand UO_1067 (O_1067,N_24899,N_24872);
nor UO_1068 (O_1068,N_24828,N_24912);
nor UO_1069 (O_1069,N_24953,N_24902);
and UO_1070 (O_1070,N_24991,N_24942);
or UO_1071 (O_1071,N_24854,N_24814);
nand UO_1072 (O_1072,N_24878,N_24843);
nand UO_1073 (O_1073,N_24874,N_24954);
and UO_1074 (O_1074,N_24976,N_24905);
nor UO_1075 (O_1075,N_24970,N_24822);
and UO_1076 (O_1076,N_24965,N_24905);
nor UO_1077 (O_1077,N_24945,N_24979);
nor UO_1078 (O_1078,N_24851,N_24829);
or UO_1079 (O_1079,N_24829,N_24801);
and UO_1080 (O_1080,N_24869,N_24870);
or UO_1081 (O_1081,N_24829,N_24998);
and UO_1082 (O_1082,N_24952,N_24810);
or UO_1083 (O_1083,N_24986,N_24969);
nor UO_1084 (O_1084,N_24955,N_24987);
nor UO_1085 (O_1085,N_24871,N_24946);
and UO_1086 (O_1086,N_24996,N_24868);
xor UO_1087 (O_1087,N_24833,N_24806);
nor UO_1088 (O_1088,N_24825,N_24851);
or UO_1089 (O_1089,N_24831,N_24954);
nor UO_1090 (O_1090,N_24948,N_24982);
nor UO_1091 (O_1091,N_24946,N_24816);
and UO_1092 (O_1092,N_24939,N_24809);
and UO_1093 (O_1093,N_24980,N_24863);
nand UO_1094 (O_1094,N_24895,N_24885);
or UO_1095 (O_1095,N_24934,N_24939);
or UO_1096 (O_1096,N_24867,N_24897);
or UO_1097 (O_1097,N_24827,N_24876);
nor UO_1098 (O_1098,N_24865,N_24919);
and UO_1099 (O_1099,N_24969,N_24872);
and UO_1100 (O_1100,N_24975,N_24922);
or UO_1101 (O_1101,N_24827,N_24960);
nand UO_1102 (O_1102,N_24819,N_24849);
or UO_1103 (O_1103,N_24835,N_24940);
or UO_1104 (O_1104,N_24868,N_24957);
nor UO_1105 (O_1105,N_24810,N_24948);
and UO_1106 (O_1106,N_24908,N_24995);
nand UO_1107 (O_1107,N_24846,N_24935);
and UO_1108 (O_1108,N_24851,N_24950);
nand UO_1109 (O_1109,N_24906,N_24917);
nor UO_1110 (O_1110,N_24997,N_24941);
or UO_1111 (O_1111,N_24944,N_24815);
nand UO_1112 (O_1112,N_24943,N_24890);
and UO_1113 (O_1113,N_24820,N_24999);
nor UO_1114 (O_1114,N_24983,N_24966);
or UO_1115 (O_1115,N_24920,N_24851);
nor UO_1116 (O_1116,N_24849,N_24868);
or UO_1117 (O_1117,N_24841,N_24834);
and UO_1118 (O_1118,N_24820,N_24899);
nand UO_1119 (O_1119,N_24857,N_24848);
or UO_1120 (O_1120,N_24864,N_24834);
nand UO_1121 (O_1121,N_24894,N_24887);
nor UO_1122 (O_1122,N_24941,N_24934);
nor UO_1123 (O_1123,N_24926,N_24836);
nand UO_1124 (O_1124,N_24969,N_24943);
and UO_1125 (O_1125,N_24892,N_24899);
and UO_1126 (O_1126,N_24844,N_24814);
nand UO_1127 (O_1127,N_24823,N_24931);
nor UO_1128 (O_1128,N_24811,N_24930);
and UO_1129 (O_1129,N_24923,N_24970);
and UO_1130 (O_1130,N_24872,N_24876);
or UO_1131 (O_1131,N_24854,N_24861);
nand UO_1132 (O_1132,N_24861,N_24875);
nor UO_1133 (O_1133,N_24869,N_24888);
nor UO_1134 (O_1134,N_24875,N_24918);
nand UO_1135 (O_1135,N_24871,N_24945);
or UO_1136 (O_1136,N_24890,N_24906);
nor UO_1137 (O_1137,N_24964,N_24910);
or UO_1138 (O_1138,N_24967,N_24875);
nor UO_1139 (O_1139,N_24914,N_24890);
nand UO_1140 (O_1140,N_24953,N_24957);
and UO_1141 (O_1141,N_24858,N_24815);
nor UO_1142 (O_1142,N_24903,N_24909);
or UO_1143 (O_1143,N_24922,N_24822);
and UO_1144 (O_1144,N_24852,N_24883);
nand UO_1145 (O_1145,N_24874,N_24879);
and UO_1146 (O_1146,N_24896,N_24987);
or UO_1147 (O_1147,N_24992,N_24903);
nand UO_1148 (O_1148,N_24944,N_24919);
or UO_1149 (O_1149,N_24932,N_24877);
or UO_1150 (O_1150,N_24960,N_24811);
nor UO_1151 (O_1151,N_24844,N_24898);
or UO_1152 (O_1152,N_24820,N_24967);
nand UO_1153 (O_1153,N_24977,N_24905);
nand UO_1154 (O_1154,N_24912,N_24842);
and UO_1155 (O_1155,N_24942,N_24845);
and UO_1156 (O_1156,N_24869,N_24912);
nor UO_1157 (O_1157,N_24998,N_24951);
nand UO_1158 (O_1158,N_24859,N_24851);
and UO_1159 (O_1159,N_24826,N_24865);
nor UO_1160 (O_1160,N_24933,N_24860);
nand UO_1161 (O_1161,N_24948,N_24885);
or UO_1162 (O_1162,N_24942,N_24965);
nor UO_1163 (O_1163,N_24888,N_24821);
nand UO_1164 (O_1164,N_24964,N_24867);
or UO_1165 (O_1165,N_24844,N_24965);
nand UO_1166 (O_1166,N_24885,N_24975);
nand UO_1167 (O_1167,N_24980,N_24847);
and UO_1168 (O_1168,N_24865,N_24837);
nor UO_1169 (O_1169,N_24979,N_24856);
nor UO_1170 (O_1170,N_24945,N_24913);
nor UO_1171 (O_1171,N_24939,N_24990);
or UO_1172 (O_1172,N_24983,N_24897);
nor UO_1173 (O_1173,N_24856,N_24985);
nor UO_1174 (O_1174,N_24976,N_24904);
or UO_1175 (O_1175,N_24918,N_24834);
or UO_1176 (O_1176,N_24835,N_24969);
or UO_1177 (O_1177,N_24989,N_24830);
and UO_1178 (O_1178,N_24895,N_24859);
and UO_1179 (O_1179,N_24936,N_24853);
nand UO_1180 (O_1180,N_24898,N_24996);
and UO_1181 (O_1181,N_24982,N_24818);
nor UO_1182 (O_1182,N_24976,N_24848);
nand UO_1183 (O_1183,N_24914,N_24917);
nor UO_1184 (O_1184,N_24982,N_24823);
nand UO_1185 (O_1185,N_24937,N_24868);
and UO_1186 (O_1186,N_24964,N_24849);
nor UO_1187 (O_1187,N_24825,N_24918);
or UO_1188 (O_1188,N_24837,N_24809);
nand UO_1189 (O_1189,N_24862,N_24991);
nand UO_1190 (O_1190,N_24934,N_24808);
nor UO_1191 (O_1191,N_24964,N_24870);
nor UO_1192 (O_1192,N_24873,N_24832);
or UO_1193 (O_1193,N_24829,N_24864);
nand UO_1194 (O_1194,N_24886,N_24810);
and UO_1195 (O_1195,N_24847,N_24999);
nand UO_1196 (O_1196,N_24818,N_24957);
and UO_1197 (O_1197,N_24944,N_24986);
nor UO_1198 (O_1198,N_24865,N_24996);
nor UO_1199 (O_1199,N_24867,N_24856);
nand UO_1200 (O_1200,N_24985,N_24894);
nor UO_1201 (O_1201,N_24847,N_24868);
or UO_1202 (O_1202,N_24983,N_24976);
nor UO_1203 (O_1203,N_24847,N_24829);
nor UO_1204 (O_1204,N_24808,N_24878);
nand UO_1205 (O_1205,N_24991,N_24929);
nand UO_1206 (O_1206,N_24891,N_24957);
nor UO_1207 (O_1207,N_24806,N_24893);
and UO_1208 (O_1208,N_24874,N_24809);
or UO_1209 (O_1209,N_24905,N_24823);
and UO_1210 (O_1210,N_24999,N_24804);
and UO_1211 (O_1211,N_24972,N_24988);
or UO_1212 (O_1212,N_24867,N_24911);
nand UO_1213 (O_1213,N_24944,N_24970);
or UO_1214 (O_1214,N_24856,N_24822);
nor UO_1215 (O_1215,N_24989,N_24809);
nand UO_1216 (O_1216,N_24968,N_24802);
or UO_1217 (O_1217,N_24958,N_24947);
and UO_1218 (O_1218,N_24935,N_24872);
and UO_1219 (O_1219,N_24859,N_24969);
and UO_1220 (O_1220,N_24906,N_24967);
and UO_1221 (O_1221,N_24826,N_24973);
nand UO_1222 (O_1222,N_24938,N_24883);
and UO_1223 (O_1223,N_24937,N_24994);
nor UO_1224 (O_1224,N_24868,N_24954);
or UO_1225 (O_1225,N_24847,N_24838);
nor UO_1226 (O_1226,N_24956,N_24997);
and UO_1227 (O_1227,N_24922,N_24930);
xor UO_1228 (O_1228,N_24934,N_24906);
nand UO_1229 (O_1229,N_24830,N_24900);
and UO_1230 (O_1230,N_24813,N_24916);
nor UO_1231 (O_1231,N_24948,N_24821);
and UO_1232 (O_1232,N_24829,N_24815);
nor UO_1233 (O_1233,N_24899,N_24863);
nand UO_1234 (O_1234,N_24906,N_24879);
nor UO_1235 (O_1235,N_24906,N_24811);
or UO_1236 (O_1236,N_24990,N_24847);
nand UO_1237 (O_1237,N_24942,N_24998);
nand UO_1238 (O_1238,N_24823,N_24829);
or UO_1239 (O_1239,N_24912,N_24934);
nand UO_1240 (O_1240,N_24904,N_24899);
or UO_1241 (O_1241,N_24818,N_24817);
and UO_1242 (O_1242,N_24858,N_24823);
nand UO_1243 (O_1243,N_24982,N_24863);
nor UO_1244 (O_1244,N_24874,N_24959);
nand UO_1245 (O_1245,N_24850,N_24968);
or UO_1246 (O_1246,N_24960,N_24871);
or UO_1247 (O_1247,N_24892,N_24886);
nand UO_1248 (O_1248,N_24968,N_24909);
nand UO_1249 (O_1249,N_24874,N_24923);
nand UO_1250 (O_1250,N_24900,N_24817);
and UO_1251 (O_1251,N_24884,N_24926);
or UO_1252 (O_1252,N_24812,N_24950);
and UO_1253 (O_1253,N_24835,N_24843);
and UO_1254 (O_1254,N_24909,N_24857);
or UO_1255 (O_1255,N_24808,N_24872);
and UO_1256 (O_1256,N_24929,N_24822);
nand UO_1257 (O_1257,N_24892,N_24833);
and UO_1258 (O_1258,N_24893,N_24888);
and UO_1259 (O_1259,N_24953,N_24836);
or UO_1260 (O_1260,N_24851,N_24865);
or UO_1261 (O_1261,N_24964,N_24842);
or UO_1262 (O_1262,N_24910,N_24986);
nand UO_1263 (O_1263,N_24889,N_24937);
nor UO_1264 (O_1264,N_24943,N_24867);
nor UO_1265 (O_1265,N_24850,N_24895);
or UO_1266 (O_1266,N_24948,N_24973);
and UO_1267 (O_1267,N_24850,N_24956);
or UO_1268 (O_1268,N_24869,N_24895);
or UO_1269 (O_1269,N_24878,N_24800);
and UO_1270 (O_1270,N_24970,N_24903);
or UO_1271 (O_1271,N_24901,N_24949);
or UO_1272 (O_1272,N_24965,N_24924);
and UO_1273 (O_1273,N_24933,N_24999);
nand UO_1274 (O_1274,N_24837,N_24971);
or UO_1275 (O_1275,N_24986,N_24834);
nand UO_1276 (O_1276,N_24910,N_24979);
nand UO_1277 (O_1277,N_24815,N_24904);
nand UO_1278 (O_1278,N_24828,N_24948);
nor UO_1279 (O_1279,N_24905,N_24807);
nor UO_1280 (O_1280,N_24969,N_24858);
nor UO_1281 (O_1281,N_24901,N_24985);
nor UO_1282 (O_1282,N_24874,N_24985);
nor UO_1283 (O_1283,N_24890,N_24929);
nor UO_1284 (O_1284,N_24985,N_24806);
or UO_1285 (O_1285,N_24989,N_24875);
nor UO_1286 (O_1286,N_24896,N_24858);
nand UO_1287 (O_1287,N_24974,N_24805);
nand UO_1288 (O_1288,N_24838,N_24938);
nand UO_1289 (O_1289,N_24965,N_24909);
nor UO_1290 (O_1290,N_24969,N_24855);
nand UO_1291 (O_1291,N_24856,N_24875);
and UO_1292 (O_1292,N_24858,N_24919);
nor UO_1293 (O_1293,N_24922,N_24856);
nand UO_1294 (O_1294,N_24859,N_24816);
nand UO_1295 (O_1295,N_24996,N_24872);
xnor UO_1296 (O_1296,N_24974,N_24999);
and UO_1297 (O_1297,N_24961,N_24976);
or UO_1298 (O_1298,N_24962,N_24828);
and UO_1299 (O_1299,N_24867,N_24861);
or UO_1300 (O_1300,N_24890,N_24973);
or UO_1301 (O_1301,N_24951,N_24867);
nand UO_1302 (O_1302,N_24961,N_24832);
or UO_1303 (O_1303,N_24891,N_24802);
nor UO_1304 (O_1304,N_24971,N_24924);
nand UO_1305 (O_1305,N_24805,N_24989);
nand UO_1306 (O_1306,N_24838,N_24933);
nor UO_1307 (O_1307,N_24891,N_24974);
nor UO_1308 (O_1308,N_24979,N_24920);
and UO_1309 (O_1309,N_24821,N_24988);
nand UO_1310 (O_1310,N_24991,N_24830);
or UO_1311 (O_1311,N_24832,N_24826);
and UO_1312 (O_1312,N_24900,N_24925);
and UO_1313 (O_1313,N_24956,N_24889);
nor UO_1314 (O_1314,N_24985,N_24876);
xnor UO_1315 (O_1315,N_24905,N_24813);
or UO_1316 (O_1316,N_24975,N_24858);
nand UO_1317 (O_1317,N_24800,N_24889);
nand UO_1318 (O_1318,N_24800,N_24840);
nor UO_1319 (O_1319,N_24831,N_24936);
nor UO_1320 (O_1320,N_24925,N_24960);
nand UO_1321 (O_1321,N_24880,N_24847);
nor UO_1322 (O_1322,N_24832,N_24883);
nor UO_1323 (O_1323,N_24801,N_24963);
nand UO_1324 (O_1324,N_24966,N_24806);
nand UO_1325 (O_1325,N_24886,N_24831);
nand UO_1326 (O_1326,N_24909,N_24918);
and UO_1327 (O_1327,N_24942,N_24886);
nand UO_1328 (O_1328,N_24874,N_24855);
or UO_1329 (O_1329,N_24974,N_24990);
or UO_1330 (O_1330,N_24907,N_24942);
nor UO_1331 (O_1331,N_24988,N_24875);
and UO_1332 (O_1332,N_24860,N_24939);
nand UO_1333 (O_1333,N_24891,N_24825);
nor UO_1334 (O_1334,N_24989,N_24920);
or UO_1335 (O_1335,N_24999,N_24810);
and UO_1336 (O_1336,N_24846,N_24943);
nand UO_1337 (O_1337,N_24846,N_24974);
nor UO_1338 (O_1338,N_24984,N_24814);
or UO_1339 (O_1339,N_24836,N_24839);
or UO_1340 (O_1340,N_24905,N_24913);
nor UO_1341 (O_1341,N_24848,N_24947);
and UO_1342 (O_1342,N_24907,N_24914);
and UO_1343 (O_1343,N_24998,N_24881);
xnor UO_1344 (O_1344,N_24946,N_24879);
and UO_1345 (O_1345,N_24903,N_24916);
or UO_1346 (O_1346,N_24806,N_24925);
nor UO_1347 (O_1347,N_24981,N_24821);
nor UO_1348 (O_1348,N_24962,N_24905);
or UO_1349 (O_1349,N_24924,N_24932);
or UO_1350 (O_1350,N_24999,N_24826);
or UO_1351 (O_1351,N_24850,N_24811);
or UO_1352 (O_1352,N_24959,N_24808);
nor UO_1353 (O_1353,N_24888,N_24928);
or UO_1354 (O_1354,N_24888,N_24830);
nand UO_1355 (O_1355,N_24930,N_24957);
or UO_1356 (O_1356,N_24970,N_24918);
nor UO_1357 (O_1357,N_24816,N_24996);
or UO_1358 (O_1358,N_24915,N_24840);
or UO_1359 (O_1359,N_24817,N_24808);
nand UO_1360 (O_1360,N_24899,N_24876);
or UO_1361 (O_1361,N_24978,N_24948);
or UO_1362 (O_1362,N_24920,N_24898);
and UO_1363 (O_1363,N_24856,N_24827);
or UO_1364 (O_1364,N_24866,N_24919);
nand UO_1365 (O_1365,N_24953,N_24892);
or UO_1366 (O_1366,N_24896,N_24848);
nor UO_1367 (O_1367,N_24810,N_24907);
and UO_1368 (O_1368,N_24871,N_24936);
nor UO_1369 (O_1369,N_24961,N_24950);
nand UO_1370 (O_1370,N_24943,N_24828);
nor UO_1371 (O_1371,N_24864,N_24817);
or UO_1372 (O_1372,N_24804,N_24979);
nor UO_1373 (O_1373,N_24887,N_24990);
or UO_1374 (O_1374,N_24833,N_24985);
and UO_1375 (O_1375,N_24924,N_24915);
or UO_1376 (O_1376,N_24917,N_24944);
nand UO_1377 (O_1377,N_24978,N_24886);
nor UO_1378 (O_1378,N_24937,N_24946);
nor UO_1379 (O_1379,N_24831,N_24876);
nand UO_1380 (O_1380,N_24878,N_24955);
nand UO_1381 (O_1381,N_24833,N_24885);
and UO_1382 (O_1382,N_24856,N_24802);
nor UO_1383 (O_1383,N_24823,N_24855);
nor UO_1384 (O_1384,N_24860,N_24916);
nand UO_1385 (O_1385,N_24857,N_24867);
or UO_1386 (O_1386,N_24868,N_24975);
nor UO_1387 (O_1387,N_24806,N_24904);
or UO_1388 (O_1388,N_24951,N_24834);
or UO_1389 (O_1389,N_24835,N_24864);
nand UO_1390 (O_1390,N_24839,N_24827);
or UO_1391 (O_1391,N_24819,N_24948);
or UO_1392 (O_1392,N_24884,N_24879);
and UO_1393 (O_1393,N_24842,N_24803);
and UO_1394 (O_1394,N_24930,N_24939);
nand UO_1395 (O_1395,N_24933,N_24890);
nand UO_1396 (O_1396,N_24830,N_24829);
or UO_1397 (O_1397,N_24974,N_24938);
or UO_1398 (O_1398,N_24978,N_24892);
and UO_1399 (O_1399,N_24951,N_24993);
and UO_1400 (O_1400,N_24842,N_24889);
and UO_1401 (O_1401,N_24952,N_24854);
or UO_1402 (O_1402,N_24929,N_24896);
nor UO_1403 (O_1403,N_24838,N_24911);
nor UO_1404 (O_1404,N_24812,N_24826);
nand UO_1405 (O_1405,N_24948,N_24928);
and UO_1406 (O_1406,N_24931,N_24992);
and UO_1407 (O_1407,N_24818,N_24967);
nor UO_1408 (O_1408,N_24877,N_24921);
or UO_1409 (O_1409,N_24993,N_24839);
nor UO_1410 (O_1410,N_24842,N_24921);
nor UO_1411 (O_1411,N_24899,N_24871);
nor UO_1412 (O_1412,N_24896,N_24855);
nor UO_1413 (O_1413,N_24950,N_24988);
nand UO_1414 (O_1414,N_24902,N_24983);
or UO_1415 (O_1415,N_24875,N_24951);
and UO_1416 (O_1416,N_24914,N_24935);
and UO_1417 (O_1417,N_24841,N_24949);
nor UO_1418 (O_1418,N_24981,N_24943);
nor UO_1419 (O_1419,N_24852,N_24964);
or UO_1420 (O_1420,N_24903,N_24908);
and UO_1421 (O_1421,N_24932,N_24839);
or UO_1422 (O_1422,N_24932,N_24808);
or UO_1423 (O_1423,N_24818,N_24925);
nor UO_1424 (O_1424,N_24928,N_24831);
and UO_1425 (O_1425,N_24876,N_24883);
nor UO_1426 (O_1426,N_24877,N_24813);
xnor UO_1427 (O_1427,N_24952,N_24979);
or UO_1428 (O_1428,N_24988,N_24850);
and UO_1429 (O_1429,N_24818,N_24808);
nand UO_1430 (O_1430,N_24801,N_24955);
or UO_1431 (O_1431,N_24816,N_24861);
or UO_1432 (O_1432,N_24958,N_24943);
nor UO_1433 (O_1433,N_24880,N_24922);
nor UO_1434 (O_1434,N_24879,N_24896);
nand UO_1435 (O_1435,N_24874,N_24847);
nor UO_1436 (O_1436,N_24995,N_24943);
and UO_1437 (O_1437,N_24924,N_24867);
nor UO_1438 (O_1438,N_24908,N_24921);
nand UO_1439 (O_1439,N_24882,N_24917);
nor UO_1440 (O_1440,N_24868,N_24972);
nand UO_1441 (O_1441,N_24912,N_24976);
nor UO_1442 (O_1442,N_24988,N_24873);
or UO_1443 (O_1443,N_24802,N_24995);
and UO_1444 (O_1444,N_24949,N_24970);
nand UO_1445 (O_1445,N_24866,N_24907);
xnor UO_1446 (O_1446,N_24977,N_24964);
or UO_1447 (O_1447,N_24927,N_24854);
nor UO_1448 (O_1448,N_24833,N_24871);
and UO_1449 (O_1449,N_24831,N_24853);
and UO_1450 (O_1450,N_24963,N_24934);
nand UO_1451 (O_1451,N_24925,N_24805);
nor UO_1452 (O_1452,N_24810,N_24945);
or UO_1453 (O_1453,N_24974,N_24985);
or UO_1454 (O_1454,N_24990,N_24866);
nor UO_1455 (O_1455,N_24832,N_24929);
nor UO_1456 (O_1456,N_24870,N_24844);
nand UO_1457 (O_1457,N_24910,N_24834);
nor UO_1458 (O_1458,N_24837,N_24977);
and UO_1459 (O_1459,N_24813,N_24895);
nor UO_1460 (O_1460,N_24826,N_24921);
nor UO_1461 (O_1461,N_24858,N_24800);
and UO_1462 (O_1462,N_24849,N_24885);
nor UO_1463 (O_1463,N_24920,N_24952);
or UO_1464 (O_1464,N_24872,N_24844);
nand UO_1465 (O_1465,N_24852,N_24923);
or UO_1466 (O_1466,N_24912,N_24931);
and UO_1467 (O_1467,N_24805,N_24975);
or UO_1468 (O_1468,N_24938,N_24983);
or UO_1469 (O_1469,N_24955,N_24840);
nor UO_1470 (O_1470,N_24884,N_24974);
nor UO_1471 (O_1471,N_24804,N_24930);
nand UO_1472 (O_1472,N_24952,N_24862);
and UO_1473 (O_1473,N_24877,N_24958);
and UO_1474 (O_1474,N_24957,N_24960);
or UO_1475 (O_1475,N_24990,N_24940);
nor UO_1476 (O_1476,N_24891,N_24922);
or UO_1477 (O_1477,N_24884,N_24800);
and UO_1478 (O_1478,N_24884,N_24890);
xnor UO_1479 (O_1479,N_24875,N_24806);
nor UO_1480 (O_1480,N_24822,N_24826);
and UO_1481 (O_1481,N_24847,N_24953);
and UO_1482 (O_1482,N_24986,N_24846);
nor UO_1483 (O_1483,N_24992,N_24890);
and UO_1484 (O_1484,N_24911,N_24915);
and UO_1485 (O_1485,N_24902,N_24999);
nand UO_1486 (O_1486,N_24827,N_24835);
nor UO_1487 (O_1487,N_24804,N_24906);
and UO_1488 (O_1488,N_24811,N_24869);
nor UO_1489 (O_1489,N_24951,N_24974);
nor UO_1490 (O_1490,N_24837,N_24905);
nand UO_1491 (O_1491,N_24939,N_24873);
nor UO_1492 (O_1492,N_24915,N_24810);
nor UO_1493 (O_1493,N_24942,N_24901);
or UO_1494 (O_1494,N_24845,N_24911);
and UO_1495 (O_1495,N_24856,N_24858);
or UO_1496 (O_1496,N_24802,N_24821);
or UO_1497 (O_1497,N_24856,N_24951);
nand UO_1498 (O_1498,N_24896,N_24933);
nand UO_1499 (O_1499,N_24988,N_24853);
nand UO_1500 (O_1500,N_24954,N_24870);
or UO_1501 (O_1501,N_24863,N_24859);
or UO_1502 (O_1502,N_24859,N_24871);
or UO_1503 (O_1503,N_24856,N_24925);
or UO_1504 (O_1504,N_24852,N_24970);
nor UO_1505 (O_1505,N_24963,N_24977);
nor UO_1506 (O_1506,N_24927,N_24850);
nand UO_1507 (O_1507,N_24877,N_24807);
or UO_1508 (O_1508,N_24858,N_24974);
and UO_1509 (O_1509,N_24915,N_24949);
nand UO_1510 (O_1510,N_24952,N_24840);
nand UO_1511 (O_1511,N_24974,N_24914);
and UO_1512 (O_1512,N_24868,N_24870);
or UO_1513 (O_1513,N_24903,N_24907);
nor UO_1514 (O_1514,N_24988,N_24804);
nor UO_1515 (O_1515,N_24801,N_24960);
or UO_1516 (O_1516,N_24841,N_24859);
nor UO_1517 (O_1517,N_24944,N_24848);
nand UO_1518 (O_1518,N_24859,N_24978);
nand UO_1519 (O_1519,N_24935,N_24921);
nand UO_1520 (O_1520,N_24808,N_24874);
nand UO_1521 (O_1521,N_24998,N_24867);
and UO_1522 (O_1522,N_24990,N_24888);
and UO_1523 (O_1523,N_24959,N_24836);
or UO_1524 (O_1524,N_24961,N_24847);
nor UO_1525 (O_1525,N_24935,N_24875);
and UO_1526 (O_1526,N_24929,N_24952);
nor UO_1527 (O_1527,N_24859,N_24906);
or UO_1528 (O_1528,N_24890,N_24830);
and UO_1529 (O_1529,N_24935,N_24828);
and UO_1530 (O_1530,N_24912,N_24810);
nand UO_1531 (O_1531,N_24925,N_24974);
or UO_1532 (O_1532,N_24896,N_24817);
nand UO_1533 (O_1533,N_24961,N_24815);
nor UO_1534 (O_1534,N_24961,N_24866);
or UO_1535 (O_1535,N_24889,N_24810);
and UO_1536 (O_1536,N_24812,N_24937);
or UO_1537 (O_1537,N_24984,N_24882);
or UO_1538 (O_1538,N_24812,N_24900);
nor UO_1539 (O_1539,N_24802,N_24848);
or UO_1540 (O_1540,N_24953,N_24839);
and UO_1541 (O_1541,N_24840,N_24866);
or UO_1542 (O_1542,N_24925,N_24865);
nor UO_1543 (O_1543,N_24836,N_24810);
nand UO_1544 (O_1544,N_24959,N_24933);
nand UO_1545 (O_1545,N_24956,N_24992);
and UO_1546 (O_1546,N_24831,N_24826);
or UO_1547 (O_1547,N_24819,N_24830);
nand UO_1548 (O_1548,N_24847,N_24936);
or UO_1549 (O_1549,N_24863,N_24812);
nor UO_1550 (O_1550,N_24997,N_24955);
nand UO_1551 (O_1551,N_24813,N_24820);
nor UO_1552 (O_1552,N_24932,N_24870);
or UO_1553 (O_1553,N_24895,N_24999);
or UO_1554 (O_1554,N_24840,N_24908);
nor UO_1555 (O_1555,N_24985,N_24890);
and UO_1556 (O_1556,N_24825,N_24943);
and UO_1557 (O_1557,N_24905,N_24930);
or UO_1558 (O_1558,N_24949,N_24834);
nor UO_1559 (O_1559,N_24977,N_24800);
nand UO_1560 (O_1560,N_24920,N_24808);
and UO_1561 (O_1561,N_24851,N_24904);
or UO_1562 (O_1562,N_24996,N_24929);
nand UO_1563 (O_1563,N_24977,N_24957);
and UO_1564 (O_1564,N_24902,N_24890);
nor UO_1565 (O_1565,N_24974,N_24803);
nand UO_1566 (O_1566,N_24909,N_24855);
or UO_1567 (O_1567,N_24890,N_24860);
or UO_1568 (O_1568,N_24976,N_24926);
nor UO_1569 (O_1569,N_24847,N_24881);
or UO_1570 (O_1570,N_24884,N_24839);
or UO_1571 (O_1571,N_24970,N_24853);
or UO_1572 (O_1572,N_24975,N_24940);
or UO_1573 (O_1573,N_24991,N_24928);
nor UO_1574 (O_1574,N_24854,N_24977);
nand UO_1575 (O_1575,N_24948,N_24954);
nand UO_1576 (O_1576,N_24986,N_24977);
nor UO_1577 (O_1577,N_24962,N_24822);
nand UO_1578 (O_1578,N_24875,N_24860);
or UO_1579 (O_1579,N_24997,N_24824);
or UO_1580 (O_1580,N_24842,N_24847);
or UO_1581 (O_1581,N_24994,N_24910);
or UO_1582 (O_1582,N_24902,N_24813);
nor UO_1583 (O_1583,N_24961,N_24998);
or UO_1584 (O_1584,N_24868,N_24910);
xor UO_1585 (O_1585,N_24990,N_24820);
or UO_1586 (O_1586,N_24923,N_24855);
nor UO_1587 (O_1587,N_24955,N_24901);
nor UO_1588 (O_1588,N_24998,N_24925);
nor UO_1589 (O_1589,N_24901,N_24804);
and UO_1590 (O_1590,N_24977,N_24822);
and UO_1591 (O_1591,N_24970,N_24947);
nor UO_1592 (O_1592,N_24925,N_24862);
nand UO_1593 (O_1593,N_24988,N_24892);
nor UO_1594 (O_1594,N_24978,N_24957);
or UO_1595 (O_1595,N_24860,N_24802);
nand UO_1596 (O_1596,N_24810,N_24927);
and UO_1597 (O_1597,N_24993,N_24922);
nor UO_1598 (O_1598,N_24910,N_24961);
nand UO_1599 (O_1599,N_24989,N_24996);
and UO_1600 (O_1600,N_24837,N_24867);
nor UO_1601 (O_1601,N_24995,N_24898);
or UO_1602 (O_1602,N_24813,N_24805);
or UO_1603 (O_1603,N_24862,N_24860);
and UO_1604 (O_1604,N_24868,N_24817);
and UO_1605 (O_1605,N_24966,N_24801);
or UO_1606 (O_1606,N_24995,N_24852);
nand UO_1607 (O_1607,N_24845,N_24972);
nor UO_1608 (O_1608,N_24907,N_24918);
and UO_1609 (O_1609,N_24809,N_24946);
or UO_1610 (O_1610,N_24810,N_24807);
nand UO_1611 (O_1611,N_24997,N_24926);
xor UO_1612 (O_1612,N_24916,N_24992);
nor UO_1613 (O_1613,N_24899,N_24829);
nor UO_1614 (O_1614,N_24994,N_24981);
and UO_1615 (O_1615,N_24854,N_24809);
and UO_1616 (O_1616,N_24960,N_24916);
nand UO_1617 (O_1617,N_24912,N_24929);
and UO_1618 (O_1618,N_24868,N_24891);
or UO_1619 (O_1619,N_24935,N_24890);
nand UO_1620 (O_1620,N_24953,N_24830);
and UO_1621 (O_1621,N_24807,N_24813);
or UO_1622 (O_1622,N_24953,N_24821);
nand UO_1623 (O_1623,N_24921,N_24976);
and UO_1624 (O_1624,N_24904,N_24893);
and UO_1625 (O_1625,N_24936,N_24863);
and UO_1626 (O_1626,N_24860,N_24832);
and UO_1627 (O_1627,N_24826,N_24988);
or UO_1628 (O_1628,N_24993,N_24849);
nor UO_1629 (O_1629,N_24800,N_24835);
or UO_1630 (O_1630,N_24876,N_24813);
and UO_1631 (O_1631,N_24967,N_24993);
and UO_1632 (O_1632,N_24859,N_24896);
nor UO_1633 (O_1633,N_24866,N_24979);
nand UO_1634 (O_1634,N_24944,N_24804);
or UO_1635 (O_1635,N_24940,N_24939);
nor UO_1636 (O_1636,N_24814,N_24808);
or UO_1637 (O_1637,N_24988,N_24841);
or UO_1638 (O_1638,N_24930,N_24937);
xor UO_1639 (O_1639,N_24899,N_24964);
nand UO_1640 (O_1640,N_24945,N_24814);
and UO_1641 (O_1641,N_24814,N_24940);
or UO_1642 (O_1642,N_24949,N_24908);
nor UO_1643 (O_1643,N_24904,N_24977);
nand UO_1644 (O_1644,N_24914,N_24954);
or UO_1645 (O_1645,N_24830,N_24908);
or UO_1646 (O_1646,N_24907,N_24922);
and UO_1647 (O_1647,N_24966,N_24972);
or UO_1648 (O_1648,N_24959,N_24969);
nor UO_1649 (O_1649,N_24860,N_24976);
or UO_1650 (O_1650,N_24852,N_24846);
and UO_1651 (O_1651,N_24951,N_24979);
nor UO_1652 (O_1652,N_24962,N_24978);
or UO_1653 (O_1653,N_24889,N_24994);
or UO_1654 (O_1654,N_24902,N_24801);
nand UO_1655 (O_1655,N_24884,N_24976);
nand UO_1656 (O_1656,N_24843,N_24931);
nor UO_1657 (O_1657,N_24850,N_24981);
nand UO_1658 (O_1658,N_24992,N_24922);
nand UO_1659 (O_1659,N_24998,N_24920);
and UO_1660 (O_1660,N_24877,N_24956);
nand UO_1661 (O_1661,N_24875,N_24889);
nand UO_1662 (O_1662,N_24922,N_24921);
and UO_1663 (O_1663,N_24926,N_24898);
and UO_1664 (O_1664,N_24921,N_24939);
or UO_1665 (O_1665,N_24980,N_24831);
nor UO_1666 (O_1666,N_24926,N_24851);
and UO_1667 (O_1667,N_24932,N_24923);
and UO_1668 (O_1668,N_24806,N_24988);
nor UO_1669 (O_1669,N_24994,N_24968);
nand UO_1670 (O_1670,N_24858,N_24861);
nand UO_1671 (O_1671,N_24975,N_24964);
and UO_1672 (O_1672,N_24924,N_24957);
or UO_1673 (O_1673,N_24959,N_24978);
nor UO_1674 (O_1674,N_24878,N_24942);
and UO_1675 (O_1675,N_24993,N_24923);
nor UO_1676 (O_1676,N_24955,N_24990);
or UO_1677 (O_1677,N_24806,N_24959);
and UO_1678 (O_1678,N_24977,N_24930);
nor UO_1679 (O_1679,N_24859,N_24842);
xnor UO_1680 (O_1680,N_24811,N_24918);
and UO_1681 (O_1681,N_24964,N_24815);
or UO_1682 (O_1682,N_24947,N_24886);
nor UO_1683 (O_1683,N_24856,N_24958);
nor UO_1684 (O_1684,N_24933,N_24899);
and UO_1685 (O_1685,N_24972,N_24909);
and UO_1686 (O_1686,N_24965,N_24885);
nor UO_1687 (O_1687,N_24877,N_24822);
nand UO_1688 (O_1688,N_24830,N_24828);
nand UO_1689 (O_1689,N_24887,N_24859);
nand UO_1690 (O_1690,N_24995,N_24979);
or UO_1691 (O_1691,N_24967,N_24816);
nand UO_1692 (O_1692,N_24831,N_24923);
or UO_1693 (O_1693,N_24807,N_24987);
or UO_1694 (O_1694,N_24806,N_24982);
xnor UO_1695 (O_1695,N_24999,N_24914);
or UO_1696 (O_1696,N_24923,N_24849);
or UO_1697 (O_1697,N_24891,N_24950);
or UO_1698 (O_1698,N_24940,N_24929);
nand UO_1699 (O_1699,N_24811,N_24979);
nor UO_1700 (O_1700,N_24857,N_24953);
nand UO_1701 (O_1701,N_24924,N_24900);
nand UO_1702 (O_1702,N_24868,N_24904);
and UO_1703 (O_1703,N_24998,N_24854);
or UO_1704 (O_1704,N_24823,N_24809);
xor UO_1705 (O_1705,N_24955,N_24847);
or UO_1706 (O_1706,N_24870,N_24979);
nor UO_1707 (O_1707,N_24823,N_24956);
nand UO_1708 (O_1708,N_24991,N_24936);
nor UO_1709 (O_1709,N_24832,N_24866);
and UO_1710 (O_1710,N_24902,N_24815);
nand UO_1711 (O_1711,N_24888,N_24894);
nor UO_1712 (O_1712,N_24840,N_24938);
nand UO_1713 (O_1713,N_24949,N_24999);
or UO_1714 (O_1714,N_24938,N_24948);
nor UO_1715 (O_1715,N_24992,N_24914);
nand UO_1716 (O_1716,N_24981,N_24818);
nor UO_1717 (O_1717,N_24945,N_24931);
or UO_1718 (O_1718,N_24878,N_24869);
and UO_1719 (O_1719,N_24855,N_24982);
and UO_1720 (O_1720,N_24866,N_24962);
or UO_1721 (O_1721,N_24905,N_24844);
nand UO_1722 (O_1722,N_24985,N_24841);
nor UO_1723 (O_1723,N_24881,N_24898);
and UO_1724 (O_1724,N_24926,N_24991);
nand UO_1725 (O_1725,N_24991,N_24983);
or UO_1726 (O_1726,N_24976,N_24873);
and UO_1727 (O_1727,N_24920,N_24817);
nor UO_1728 (O_1728,N_24967,N_24881);
and UO_1729 (O_1729,N_24963,N_24802);
or UO_1730 (O_1730,N_24890,N_24930);
nand UO_1731 (O_1731,N_24819,N_24881);
nand UO_1732 (O_1732,N_24802,N_24834);
nor UO_1733 (O_1733,N_24996,N_24820);
or UO_1734 (O_1734,N_24961,N_24856);
nor UO_1735 (O_1735,N_24922,N_24970);
nor UO_1736 (O_1736,N_24877,N_24947);
or UO_1737 (O_1737,N_24954,N_24994);
nor UO_1738 (O_1738,N_24804,N_24902);
and UO_1739 (O_1739,N_24848,N_24916);
and UO_1740 (O_1740,N_24815,N_24906);
or UO_1741 (O_1741,N_24828,N_24990);
or UO_1742 (O_1742,N_24896,N_24907);
nand UO_1743 (O_1743,N_24915,N_24948);
nor UO_1744 (O_1744,N_24967,N_24814);
or UO_1745 (O_1745,N_24808,N_24903);
nor UO_1746 (O_1746,N_24893,N_24949);
or UO_1747 (O_1747,N_24873,N_24801);
nand UO_1748 (O_1748,N_24802,N_24997);
or UO_1749 (O_1749,N_24850,N_24998);
or UO_1750 (O_1750,N_24860,N_24966);
nor UO_1751 (O_1751,N_24883,N_24952);
xnor UO_1752 (O_1752,N_24974,N_24877);
and UO_1753 (O_1753,N_24916,N_24863);
and UO_1754 (O_1754,N_24991,N_24916);
nor UO_1755 (O_1755,N_24880,N_24866);
or UO_1756 (O_1756,N_24896,N_24815);
nand UO_1757 (O_1757,N_24861,N_24815);
or UO_1758 (O_1758,N_24992,N_24950);
or UO_1759 (O_1759,N_24962,N_24818);
nand UO_1760 (O_1760,N_24812,N_24964);
or UO_1761 (O_1761,N_24954,N_24809);
nand UO_1762 (O_1762,N_24806,N_24992);
or UO_1763 (O_1763,N_24870,N_24985);
nor UO_1764 (O_1764,N_24812,N_24936);
and UO_1765 (O_1765,N_24953,N_24906);
nor UO_1766 (O_1766,N_24896,N_24966);
or UO_1767 (O_1767,N_24946,N_24972);
nand UO_1768 (O_1768,N_24975,N_24828);
nand UO_1769 (O_1769,N_24919,N_24930);
or UO_1770 (O_1770,N_24837,N_24880);
or UO_1771 (O_1771,N_24930,N_24870);
and UO_1772 (O_1772,N_24815,N_24939);
nand UO_1773 (O_1773,N_24949,N_24836);
and UO_1774 (O_1774,N_24996,N_24897);
or UO_1775 (O_1775,N_24909,N_24906);
nor UO_1776 (O_1776,N_24855,N_24926);
or UO_1777 (O_1777,N_24904,N_24934);
nand UO_1778 (O_1778,N_24992,N_24994);
or UO_1779 (O_1779,N_24866,N_24904);
or UO_1780 (O_1780,N_24929,N_24967);
or UO_1781 (O_1781,N_24929,N_24999);
nand UO_1782 (O_1782,N_24812,N_24834);
nor UO_1783 (O_1783,N_24812,N_24979);
nor UO_1784 (O_1784,N_24953,N_24950);
and UO_1785 (O_1785,N_24942,N_24994);
nand UO_1786 (O_1786,N_24958,N_24926);
or UO_1787 (O_1787,N_24830,N_24938);
nor UO_1788 (O_1788,N_24964,N_24939);
and UO_1789 (O_1789,N_24885,N_24929);
nor UO_1790 (O_1790,N_24804,N_24833);
nor UO_1791 (O_1791,N_24953,N_24998);
and UO_1792 (O_1792,N_24844,N_24918);
nor UO_1793 (O_1793,N_24976,N_24817);
and UO_1794 (O_1794,N_24926,N_24979);
and UO_1795 (O_1795,N_24828,N_24857);
nor UO_1796 (O_1796,N_24850,N_24857);
nand UO_1797 (O_1797,N_24921,N_24910);
and UO_1798 (O_1798,N_24900,N_24866);
or UO_1799 (O_1799,N_24914,N_24901);
nand UO_1800 (O_1800,N_24912,N_24839);
nand UO_1801 (O_1801,N_24859,N_24826);
nor UO_1802 (O_1802,N_24909,N_24924);
nand UO_1803 (O_1803,N_24848,N_24943);
nor UO_1804 (O_1804,N_24918,N_24878);
or UO_1805 (O_1805,N_24910,N_24990);
or UO_1806 (O_1806,N_24932,N_24855);
nor UO_1807 (O_1807,N_24827,N_24927);
or UO_1808 (O_1808,N_24986,N_24845);
and UO_1809 (O_1809,N_24808,N_24854);
nor UO_1810 (O_1810,N_24807,N_24992);
nor UO_1811 (O_1811,N_24862,N_24883);
nor UO_1812 (O_1812,N_24812,N_24868);
and UO_1813 (O_1813,N_24864,N_24932);
and UO_1814 (O_1814,N_24800,N_24829);
or UO_1815 (O_1815,N_24950,N_24842);
or UO_1816 (O_1816,N_24961,N_24893);
nand UO_1817 (O_1817,N_24838,N_24971);
or UO_1818 (O_1818,N_24931,N_24882);
nand UO_1819 (O_1819,N_24816,N_24911);
nor UO_1820 (O_1820,N_24970,N_24801);
or UO_1821 (O_1821,N_24885,N_24828);
or UO_1822 (O_1822,N_24971,N_24996);
and UO_1823 (O_1823,N_24977,N_24993);
or UO_1824 (O_1824,N_24867,N_24831);
and UO_1825 (O_1825,N_24868,N_24885);
and UO_1826 (O_1826,N_24865,N_24951);
nor UO_1827 (O_1827,N_24895,N_24974);
nand UO_1828 (O_1828,N_24934,N_24825);
nand UO_1829 (O_1829,N_24940,N_24984);
nand UO_1830 (O_1830,N_24927,N_24825);
and UO_1831 (O_1831,N_24835,N_24828);
and UO_1832 (O_1832,N_24971,N_24951);
nor UO_1833 (O_1833,N_24897,N_24878);
nor UO_1834 (O_1834,N_24919,N_24862);
or UO_1835 (O_1835,N_24919,N_24967);
nor UO_1836 (O_1836,N_24802,N_24943);
nor UO_1837 (O_1837,N_24834,N_24800);
nand UO_1838 (O_1838,N_24984,N_24989);
nand UO_1839 (O_1839,N_24845,N_24835);
and UO_1840 (O_1840,N_24909,N_24862);
and UO_1841 (O_1841,N_24960,N_24817);
nand UO_1842 (O_1842,N_24871,N_24928);
and UO_1843 (O_1843,N_24944,N_24865);
nand UO_1844 (O_1844,N_24956,N_24955);
and UO_1845 (O_1845,N_24965,N_24823);
and UO_1846 (O_1846,N_24898,N_24867);
and UO_1847 (O_1847,N_24981,N_24996);
or UO_1848 (O_1848,N_24965,N_24814);
nor UO_1849 (O_1849,N_24938,N_24903);
or UO_1850 (O_1850,N_24902,N_24918);
nor UO_1851 (O_1851,N_24922,N_24967);
and UO_1852 (O_1852,N_24881,N_24932);
nand UO_1853 (O_1853,N_24992,N_24871);
nand UO_1854 (O_1854,N_24853,N_24810);
and UO_1855 (O_1855,N_24925,N_24831);
and UO_1856 (O_1856,N_24838,N_24982);
and UO_1857 (O_1857,N_24907,N_24908);
or UO_1858 (O_1858,N_24899,N_24906);
nand UO_1859 (O_1859,N_24954,N_24985);
nor UO_1860 (O_1860,N_24946,N_24890);
nand UO_1861 (O_1861,N_24984,N_24841);
xnor UO_1862 (O_1862,N_24892,N_24849);
and UO_1863 (O_1863,N_24884,N_24987);
or UO_1864 (O_1864,N_24992,N_24980);
or UO_1865 (O_1865,N_24844,N_24991);
and UO_1866 (O_1866,N_24892,N_24807);
and UO_1867 (O_1867,N_24907,N_24817);
nand UO_1868 (O_1868,N_24883,N_24869);
and UO_1869 (O_1869,N_24924,N_24848);
nor UO_1870 (O_1870,N_24860,N_24968);
nand UO_1871 (O_1871,N_24972,N_24872);
nand UO_1872 (O_1872,N_24964,N_24906);
or UO_1873 (O_1873,N_24811,N_24916);
or UO_1874 (O_1874,N_24877,N_24992);
or UO_1875 (O_1875,N_24826,N_24904);
and UO_1876 (O_1876,N_24946,N_24912);
nand UO_1877 (O_1877,N_24872,N_24894);
nor UO_1878 (O_1878,N_24931,N_24816);
or UO_1879 (O_1879,N_24805,N_24860);
nor UO_1880 (O_1880,N_24928,N_24974);
nand UO_1881 (O_1881,N_24966,N_24833);
or UO_1882 (O_1882,N_24992,N_24896);
nand UO_1883 (O_1883,N_24991,N_24864);
and UO_1884 (O_1884,N_24856,N_24990);
nand UO_1885 (O_1885,N_24944,N_24807);
nand UO_1886 (O_1886,N_24833,N_24924);
nor UO_1887 (O_1887,N_24917,N_24907);
nand UO_1888 (O_1888,N_24998,N_24818);
and UO_1889 (O_1889,N_24896,N_24983);
and UO_1890 (O_1890,N_24997,N_24823);
and UO_1891 (O_1891,N_24969,N_24975);
nand UO_1892 (O_1892,N_24923,N_24994);
and UO_1893 (O_1893,N_24824,N_24856);
and UO_1894 (O_1894,N_24833,N_24825);
or UO_1895 (O_1895,N_24838,N_24967);
nand UO_1896 (O_1896,N_24974,N_24833);
or UO_1897 (O_1897,N_24968,N_24830);
nand UO_1898 (O_1898,N_24892,N_24860);
nand UO_1899 (O_1899,N_24959,N_24926);
nand UO_1900 (O_1900,N_24853,N_24920);
and UO_1901 (O_1901,N_24844,N_24974);
nor UO_1902 (O_1902,N_24926,N_24995);
and UO_1903 (O_1903,N_24893,N_24989);
nor UO_1904 (O_1904,N_24887,N_24925);
nand UO_1905 (O_1905,N_24853,N_24964);
nand UO_1906 (O_1906,N_24819,N_24980);
nor UO_1907 (O_1907,N_24946,N_24852);
nand UO_1908 (O_1908,N_24932,N_24916);
and UO_1909 (O_1909,N_24892,N_24834);
nand UO_1910 (O_1910,N_24993,N_24812);
or UO_1911 (O_1911,N_24947,N_24885);
nand UO_1912 (O_1912,N_24892,N_24924);
and UO_1913 (O_1913,N_24877,N_24894);
nor UO_1914 (O_1914,N_24858,N_24801);
and UO_1915 (O_1915,N_24839,N_24940);
xor UO_1916 (O_1916,N_24897,N_24927);
nand UO_1917 (O_1917,N_24946,N_24901);
and UO_1918 (O_1918,N_24989,N_24873);
nand UO_1919 (O_1919,N_24954,N_24808);
and UO_1920 (O_1920,N_24947,N_24884);
or UO_1921 (O_1921,N_24862,N_24877);
nor UO_1922 (O_1922,N_24839,N_24914);
or UO_1923 (O_1923,N_24959,N_24947);
nand UO_1924 (O_1924,N_24803,N_24884);
and UO_1925 (O_1925,N_24971,N_24961);
nor UO_1926 (O_1926,N_24902,N_24800);
nor UO_1927 (O_1927,N_24882,N_24856);
or UO_1928 (O_1928,N_24922,N_24968);
nand UO_1929 (O_1929,N_24858,N_24819);
nand UO_1930 (O_1930,N_24878,N_24850);
nand UO_1931 (O_1931,N_24887,N_24909);
or UO_1932 (O_1932,N_24849,N_24818);
nand UO_1933 (O_1933,N_24806,N_24894);
nor UO_1934 (O_1934,N_24891,N_24892);
or UO_1935 (O_1935,N_24969,N_24871);
nand UO_1936 (O_1936,N_24918,N_24986);
and UO_1937 (O_1937,N_24964,N_24829);
nor UO_1938 (O_1938,N_24866,N_24980);
nor UO_1939 (O_1939,N_24992,N_24884);
and UO_1940 (O_1940,N_24960,N_24861);
or UO_1941 (O_1941,N_24808,N_24845);
nor UO_1942 (O_1942,N_24881,N_24969);
or UO_1943 (O_1943,N_24803,N_24858);
nor UO_1944 (O_1944,N_24874,N_24944);
nand UO_1945 (O_1945,N_24834,N_24913);
or UO_1946 (O_1946,N_24974,N_24868);
nor UO_1947 (O_1947,N_24972,N_24853);
or UO_1948 (O_1948,N_24883,N_24831);
and UO_1949 (O_1949,N_24992,N_24848);
nand UO_1950 (O_1950,N_24860,N_24870);
xnor UO_1951 (O_1951,N_24912,N_24845);
nand UO_1952 (O_1952,N_24961,N_24806);
and UO_1953 (O_1953,N_24954,N_24855);
or UO_1954 (O_1954,N_24852,N_24912);
nor UO_1955 (O_1955,N_24958,N_24950);
nand UO_1956 (O_1956,N_24881,N_24868);
or UO_1957 (O_1957,N_24874,N_24937);
nand UO_1958 (O_1958,N_24956,N_24831);
and UO_1959 (O_1959,N_24926,N_24887);
and UO_1960 (O_1960,N_24990,N_24854);
nor UO_1961 (O_1961,N_24934,N_24802);
nand UO_1962 (O_1962,N_24998,N_24886);
nor UO_1963 (O_1963,N_24902,N_24850);
or UO_1964 (O_1964,N_24943,N_24847);
nand UO_1965 (O_1965,N_24811,N_24885);
or UO_1966 (O_1966,N_24915,N_24828);
nand UO_1967 (O_1967,N_24966,N_24898);
and UO_1968 (O_1968,N_24946,N_24903);
nor UO_1969 (O_1969,N_24896,N_24892);
and UO_1970 (O_1970,N_24831,N_24851);
nor UO_1971 (O_1971,N_24985,N_24899);
nor UO_1972 (O_1972,N_24860,N_24871);
nand UO_1973 (O_1973,N_24867,N_24864);
or UO_1974 (O_1974,N_24988,N_24866);
xnor UO_1975 (O_1975,N_24900,N_24932);
and UO_1976 (O_1976,N_24830,N_24857);
nand UO_1977 (O_1977,N_24843,N_24848);
nand UO_1978 (O_1978,N_24876,N_24830);
and UO_1979 (O_1979,N_24843,N_24988);
or UO_1980 (O_1980,N_24928,N_24883);
nand UO_1981 (O_1981,N_24810,N_24849);
nor UO_1982 (O_1982,N_24817,N_24822);
nor UO_1983 (O_1983,N_24977,N_24848);
or UO_1984 (O_1984,N_24876,N_24878);
and UO_1985 (O_1985,N_24888,N_24809);
nand UO_1986 (O_1986,N_24853,N_24847);
or UO_1987 (O_1987,N_24837,N_24886);
or UO_1988 (O_1988,N_24855,N_24975);
and UO_1989 (O_1989,N_24819,N_24817);
and UO_1990 (O_1990,N_24807,N_24887);
nor UO_1991 (O_1991,N_24930,N_24947);
nand UO_1992 (O_1992,N_24800,N_24856);
nand UO_1993 (O_1993,N_24903,N_24949);
and UO_1994 (O_1994,N_24861,N_24856);
or UO_1995 (O_1995,N_24960,N_24915);
and UO_1996 (O_1996,N_24861,N_24965);
and UO_1997 (O_1997,N_24941,N_24976);
nor UO_1998 (O_1998,N_24983,N_24986);
or UO_1999 (O_1999,N_24952,N_24878);
or UO_2000 (O_2000,N_24834,N_24804);
nand UO_2001 (O_2001,N_24922,N_24848);
nand UO_2002 (O_2002,N_24981,N_24881);
or UO_2003 (O_2003,N_24830,N_24863);
or UO_2004 (O_2004,N_24912,N_24974);
and UO_2005 (O_2005,N_24934,N_24935);
and UO_2006 (O_2006,N_24889,N_24913);
or UO_2007 (O_2007,N_24895,N_24810);
nor UO_2008 (O_2008,N_24880,N_24907);
nor UO_2009 (O_2009,N_24825,N_24975);
and UO_2010 (O_2010,N_24853,N_24956);
nor UO_2011 (O_2011,N_24994,N_24863);
or UO_2012 (O_2012,N_24965,N_24976);
nand UO_2013 (O_2013,N_24934,N_24816);
nand UO_2014 (O_2014,N_24933,N_24848);
or UO_2015 (O_2015,N_24811,N_24887);
nand UO_2016 (O_2016,N_24908,N_24864);
nand UO_2017 (O_2017,N_24914,N_24846);
or UO_2018 (O_2018,N_24996,N_24903);
nand UO_2019 (O_2019,N_24849,N_24838);
or UO_2020 (O_2020,N_24887,N_24997);
nand UO_2021 (O_2021,N_24921,N_24924);
or UO_2022 (O_2022,N_24935,N_24883);
or UO_2023 (O_2023,N_24827,N_24974);
nand UO_2024 (O_2024,N_24869,N_24843);
and UO_2025 (O_2025,N_24880,N_24914);
xnor UO_2026 (O_2026,N_24801,N_24984);
nand UO_2027 (O_2027,N_24974,N_24829);
or UO_2028 (O_2028,N_24823,N_24826);
and UO_2029 (O_2029,N_24857,N_24977);
nor UO_2030 (O_2030,N_24990,N_24927);
nand UO_2031 (O_2031,N_24818,N_24876);
or UO_2032 (O_2032,N_24907,N_24992);
or UO_2033 (O_2033,N_24802,N_24955);
and UO_2034 (O_2034,N_24990,N_24874);
or UO_2035 (O_2035,N_24934,N_24966);
and UO_2036 (O_2036,N_24858,N_24972);
nor UO_2037 (O_2037,N_24983,N_24845);
nand UO_2038 (O_2038,N_24990,N_24916);
or UO_2039 (O_2039,N_24999,N_24811);
nand UO_2040 (O_2040,N_24934,N_24805);
nand UO_2041 (O_2041,N_24849,N_24974);
and UO_2042 (O_2042,N_24863,N_24939);
and UO_2043 (O_2043,N_24907,N_24956);
or UO_2044 (O_2044,N_24848,N_24932);
or UO_2045 (O_2045,N_24845,N_24824);
or UO_2046 (O_2046,N_24842,N_24827);
and UO_2047 (O_2047,N_24837,N_24899);
and UO_2048 (O_2048,N_24974,N_24944);
or UO_2049 (O_2049,N_24802,N_24937);
and UO_2050 (O_2050,N_24988,N_24939);
nor UO_2051 (O_2051,N_24879,N_24832);
or UO_2052 (O_2052,N_24910,N_24905);
nor UO_2053 (O_2053,N_24873,N_24903);
nand UO_2054 (O_2054,N_24921,N_24812);
nand UO_2055 (O_2055,N_24934,N_24832);
or UO_2056 (O_2056,N_24907,N_24848);
nand UO_2057 (O_2057,N_24923,N_24860);
or UO_2058 (O_2058,N_24942,N_24818);
and UO_2059 (O_2059,N_24951,N_24899);
or UO_2060 (O_2060,N_24957,N_24920);
or UO_2061 (O_2061,N_24990,N_24833);
nor UO_2062 (O_2062,N_24955,N_24800);
nor UO_2063 (O_2063,N_24838,N_24978);
nand UO_2064 (O_2064,N_24971,N_24953);
or UO_2065 (O_2065,N_24825,N_24817);
nor UO_2066 (O_2066,N_24934,N_24978);
nor UO_2067 (O_2067,N_24977,N_24989);
or UO_2068 (O_2068,N_24905,N_24894);
nor UO_2069 (O_2069,N_24919,N_24945);
nor UO_2070 (O_2070,N_24957,N_24964);
nor UO_2071 (O_2071,N_24924,N_24926);
nor UO_2072 (O_2072,N_24939,N_24965);
or UO_2073 (O_2073,N_24872,N_24814);
or UO_2074 (O_2074,N_24915,N_24877);
nor UO_2075 (O_2075,N_24814,N_24923);
or UO_2076 (O_2076,N_24927,N_24945);
nor UO_2077 (O_2077,N_24860,N_24811);
nand UO_2078 (O_2078,N_24968,N_24865);
and UO_2079 (O_2079,N_24867,N_24846);
nand UO_2080 (O_2080,N_24913,N_24829);
and UO_2081 (O_2081,N_24832,N_24976);
nand UO_2082 (O_2082,N_24838,N_24979);
and UO_2083 (O_2083,N_24927,N_24873);
nor UO_2084 (O_2084,N_24978,N_24815);
and UO_2085 (O_2085,N_24982,N_24869);
or UO_2086 (O_2086,N_24917,N_24863);
and UO_2087 (O_2087,N_24924,N_24991);
or UO_2088 (O_2088,N_24907,N_24962);
nor UO_2089 (O_2089,N_24943,N_24916);
or UO_2090 (O_2090,N_24848,N_24928);
xnor UO_2091 (O_2091,N_24964,N_24872);
and UO_2092 (O_2092,N_24899,N_24806);
and UO_2093 (O_2093,N_24995,N_24806);
or UO_2094 (O_2094,N_24833,N_24829);
nand UO_2095 (O_2095,N_24866,N_24825);
and UO_2096 (O_2096,N_24896,N_24823);
nor UO_2097 (O_2097,N_24930,N_24925);
nand UO_2098 (O_2098,N_24851,N_24824);
nor UO_2099 (O_2099,N_24958,N_24889);
nor UO_2100 (O_2100,N_24864,N_24913);
nor UO_2101 (O_2101,N_24943,N_24836);
nand UO_2102 (O_2102,N_24956,N_24867);
and UO_2103 (O_2103,N_24907,N_24969);
or UO_2104 (O_2104,N_24865,N_24934);
and UO_2105 (O_2105,N_24935,N_24842);
nor UO_2106 (O_2106,N_24898,N_24944);
nand UO_2107 (O_2107,N_24888,N_24873);
nor UO_2108 (O_2108,N_24929,N_24882);
or UO_2109 (O_2109,N_24941,N_24996);
nor UO_2110 (O_2110,N_24808,N_24835);
nand UO_2111 (O_2111,N_24881,N_24838);
or UO_2112 (O_2112,N_24999,N_24917);
and UO_2113 (O_2113,N_24967,N_24932);
and UO_2114 (O_2114,N_24871,N_24944);
nand UO_2115 (O_2115,N_24844,N_24955);
nor UO_2116 (O_2116,N_24888,N_24960);
or UO_2117 (O_2117,N_24951,N_24941);
and UO_2118 (O_2118,N_24876,N_24812);
and UO_2119 (O_2119,N_24959,N_24893);
nand UO_2120 (O_2120,N_24945,N_24859);
nor UO_2121 (O_2121,N_24865,N_24859);
nor UO_2122 (O_2122,N_24926,N_24999);
or UO_2123 (O_2123,N_24820,N_24891);
or UO_2124 (O_2124,N_24814,N_24887);
or UO_2125 (O_2125,N_24954,N_24962);
nand UO_2126 (O_2126,N_24830,N_24972);
nor UO_2127 (O_2127,N_24839,N_24818);
xnor UO_2128 (O_2128,N_24802,N_24892);
nand UO_2129 (O_2129,N_24845,N_24820);
and UO_2130 (O_2130,N_24835,N_24826);
nand UO_2131 (O_2131,N_24854,N_24953);
nand UO_2132 (O_2132,N_24876,N_24802);
nand UO_2133 (O_2133,N_24894,N_24833);
or UO_2134 (O_2134,N_24935,N_24950);
nor UO_2135 (O_2135,N_24984,N_24942);
or UO_2136 (O_2136,N_24940,N_24895);
and UO_2137 (O_2137,N_24995,N_24895);
and UO_2138 (O_2138,N_24940,N_24800);
or UO_2139 (O_2139,N_24963,N_24818);
nand UO_2140 (O_2140,N_24877,N_24980);
nor UO_2141 (O_2141,N_24819,N_24840);
nor UO_2142 (O_2142,N_24967,N_24835);
and UO_2143 (O_2143,N_24891,N_24845);
nand UO_2144 (O_2144,N_24961,N_24819);
nand UO_2145 (O_2145,N_24988,N_24947);
nor UO_2146 (O_2146,N_24835,N_24890);
nor UO_2147 (O_2147,N_24877,N_24911);
and UO_2148 (O_2148,N_24853,N_24922);
nand UO_2149 (O_2149,N_24825,N_24802);
or UO_2150 (O_2150,N_24912,N_24860);
nand UO_2151 (O_2151,N_24951,N_24861);
or UO_2152 (O_2152,N_24881,N_24859);
or UO_2153 (O_2153,N_24871,N_24866);
nand UO_2154 (O_2154,N_24990,N_24875);
and UO_2155 (O_2155,N_24972,N_24930);
nand UO_2156 (O_2156,N_24805,N_24820);
nor UO_2157 (O_2157,N_24880,N_24944);
nor UO_2158 (O_2158,N_24815,N_24949);
and UO_2159 (O_2159,N_24805,N_24881);
or UO_2160 (O_2160,N_24857,N_24933);
nand UO_2161 (O_2161,N_24995,N_24829);
nand UO_2162 (O_2162,N_24968,N_24843);
and UO_2163 (O_2163,N_24956,N_24894);
or UO_2164 (O_2164,N_24843,N_24800);
and UO_2165 (O_2165,N_24930,N_24942);
or UO_2166 (O_2166,N_24994,N_24839);
or UO_2167 (O_2167,N_24931,N_24976);
nand UO_2168 (O_2168,N_24868,N_24863);
nor UO_2169 (O_2169,N_24877,N_24847);
and UO_2170 (O_2170,N_24851,N_24860);
nand UO_2171 (O_2171,N_24948,N_24803);
nor UO_2172 (O_2172,N_24919,N_24856);
nor UO_2173 (O_2173,N_24852,N_24837);
or UO_2174 (O_2174,N_24883,N_24807);
or UO_2175 (O_2175,N_24889,N_24888);
nor UO_2176 (O_2176,N_24910,N_24852);
or UO_2177 (O_2177,N_24841,N_24925);
nand UO_2178 (O_2178,N_24849,N_24822);
nand UO_2179 (O_2179,N_24959,N_24968);
and UO_2180 (O_2180,N_24801,N_24889);
nand UO_2181 (O_2181,N_24865,N_24901);
and UO_2182 (O_2182,N_24910,N_24947);
and UO_2183 (O_2183,N_24942,N_24996);
or UO_2184 (O_2184,N_24873,N_24867);
and UO_2185 (O_2185,N_24834,N_24959);
or UO_2186 (O_2186,N_24943,N_24888);
and UO_2187 (O_2187,N_24812,N_24951);
nor UO_2188 (O_2188,N_24996,N_24832);
and UO_2189 (O_2189,N_24860,N_24822);
nor UO_2190 (O_2190,N_24933,N_24843);
and UO_2191 (O_2191,N_24891,N_24893);
or UO_2192 (O_2192,N_24954,N_24949);
nand UO_2193 (O_2193,N_24828,N_24839);
nand UO_2194 (O_2194,N_24982,N_24995);
nand UO_2195 (O_2195,N_24966,N_24914);
and UO_2196 (O_2196,N_24835,N_24961);
nand UO_2197 (O_2197,N_24962,N_24844);
or UO_2198 (O_2198,N_24867,N_24875);
and UO_2199 (O_2199,N_24969,N_24813);
nand UO_2200 (O_2200,N_24975,N_24887);
nor UO_2201 (O_2201,N_24936,N_24900);
and UO_2202 (O_2202,N_24995,N_24861);
nand UO_2203 (O_2203,N_24823,N_24845);
and UO_2204 (O_2204,N_24878,N_24934);
nor UO_2205 (O_2205,N_24909,N_24997);
nand UO_2206 (O_2206,N_24960,N_24991);
nor UO_2207 (O_2207,N_24802,N_24871);
or UO_2208 (O_2208,N_24959,N_24852);
and UO_2209 (O_2209,N_24802,N_24872);
and UO_2210 (O_2210,N_24836,N_24815);
or UO_2211 (O_2211,N_24897,N_24914);
nand UO_2212 (O_2212,N_24853,N_24870);
and UO_2213 (O_2213,N_24853,N_24944);
nand UO_2214 (O_2214,N_24862,N_24846);
nor UO_2215 (O_2215,N_24991,N_24937);
or UO_2216 (O_2216,N_24863,N_24840);
nand UO_2217 (O_2217,N_24833,N_24851);
or UO_2218 (O_2218,N_24838,N_24974);
or UO_2219 (O_2219,N_24876,N_24983);
nor UO_2220 (O_2220,N_24842,N_24955);
or UO_2221 (O_2221,N_24915,N_24974);
nor UO_2222 (O_2222,N_24977,N_24874);
or UO_2223 (O_2223,N_24900,N_24895);
nor UO_2224 (O_2224,N_24843,N_24808);
nor UO_2225 (O_2225,N_24984,N_24985);
nor UO_2226 (O_2226,N_24927,N_24979);
or UO_2227 (O_2227,N_24987,N_24902);
nor UO_2228 (O_2228,N_24836,N_24879);
and UO_2229 (O_2229,N_24930,N_24944);
or UO_2230 (O_2230,N_24942,N_24873);
or UO_2231 (O_2231,N_24876,N_24882);
or UO_2232 (O_2232,N_24832,N_24990);
nor UO_2233 (O_2233,N_24943,N_24861);
nand UO_2234 (O_2234,N_24924,N_24949);
nor UO_2235 (O_2235,N_24937,N_24852);
nand UO_2236 (O_2236,N_24984,N_24954);
and UO_2237 (O_2237,N_24933,N_24807);
and UO_2238 (O_2238,N_24887,N_24805);
and UO_2239 (O_2239,N_24817,N_24811);
or UO_2240 (O_2240,N_24978,N_24923);
nand UO_2241 (O_2241,N_24867,N_24814);
nand UO_2242 (O_2242,N_24812,N_24905);
nand UO_2243 (O_2243,N_24995,N_24853);
nand UO_2244 (O_2244,N_24934,N_24861);
and UO_2245 (O_2245,N_24954,N_24917);
nand UO_2246 (O_2246,N_24998,N_24852);
nand UO_2247 (O_2247,N_24863,N_24866);
nand UO_2248 (O_2248,N_24867,N_24979);
nand UO_2249 (O_2249,N_24926,N_24975);
nand UO_2250 (O_2250,N_24858,N_24804);
or UO_2251 (O_2251,N_24857,N_24849);
or UO_2252 (O_2252,N_24851,N_24949);
nand UO_2253 (O_2253,N_24854,N_24936);
nor UO_2254 (O_2254,N_24995,N_24934);
nor UO_2255 (O_2255,N_24973,N_24954);
and UO_2256 (O_2256,N_24908,N_24982);
nor UO_2257 (O_2257,N_24832,N_24971);
nand UO_2258 (O_2258,N_24896,N_24945);
nor UO_2259 (O_2259,N_24985,N_24848);
and UO_2260 (O_2260,N_24932,N_24945);
nand UO_2261 (O_2261,N_24944,N_24888);
nor UO_2262 (O_2262,N_24916,N_24947);
nor UO_2263 (O_2263,N_24959,N_24906);
and UO_2264 (O_2264,N_24942,N_24888);
nand UO_2265 (O_2265,N_24866,N_24807);
or UO_2266 (O_2266,N_24950,N_24863);
nand UO_2267 (O_2267,N_24979,N_24882);
nand UO_2268 (O_2268,N_24868,N_24878);
nand UO_2269 (O_2269,N_24902,N_24909);
and UO_2270 (O_2270,N_24941,N_24847);
or UO_2271 (O_2271,N_24940,N_24907);
nor UO_2272 (O_2272,N_24884,N_24925);
or UO_2273 (O_2273,N_24809,N_24910);
nor UO_2274 (O_2274,N_24810,N_24958);
nor UO_2275 (O_2275,N_24817,N_24989);
and UO_2276 (O_2276,N_24935,N_24807);
and UO_2277 (O_2277,N_24828,N_24810);
nor UO_2278 (O_2278,N_24934,N_24800);
nor UO_2279 (O_2279,N_24985,N_24832);
nand UO_2280 (O_2280,N_24926,N_24810);
and UO_2281 (O_2281,N_24916,N_24833);
nor UO_2282 (O_2282,N_24815,N_24854);
nand UO_2283 (O_2283,N_24826,N_24886);
or UO_2284 (O_2284,N_24910,N_24969);
or UO_2285 (O_2285,N_24836,N_24955);
xnor UO_2286 (O_2286,N_24848,N_24990);
nor UO_2287 (O_2287,N_24992,N_24865);
nand UO_2288 (O_2288,N_24903,N_24875);
nand UO_2289 (O_2289,N_24995,N_24960);
nor UO_2290 (O_2290,N_24966,N_24918);
nor UO_2291 (O_2291,N_24946,N_24824);
nor UO_2292 (O_2292,N_24994,N_24882);
and UO_2293 (O_2293,N_24956,N_24910);
or UO_2294 (O_2294,N_24930,N_24849);
nand UO_2295 (O_2295,N_24921,N_24932);
or UO_2296 (O_2296,N_24988,N_24931);
nor UO_2297 (O_2297,N_24926,N_24900);
and UO_2298 (O_2298,N_24982,N_24973);
nand UO_2299 (O_2299,N_24831,N_24904);
or UO_2300 (O_2300,N_24869,N_24958);
nand UO_2301 (O_2301,N_24988,N_24901);
nor UO_2302 (O_2302,N_24945,N_24977);
or UO_2303 (O_2303,N_24998,N_24940);
or UO_2304 (O_2304,N_24912,N_24897);
nand UO_2305 (O_2305,N_24835,N_24972);
nand UO_2306 (O_2306,N_24989,N_24914);
nand UO_2307 (O_2307,N_24809,N_24871);
nand UO_2308 (O_2308,N_24949,N_24938);
and UO_2309 (O_2309,N_24860,N_24838);
nand UO_2310 (O_2310,N_24928,N_24898);
and UO_2311 (O_2311,N_24919,N_24897);
and UO_2312 (O_2312,N_24849,N_24921);
or UO_2313 (O_2313,N_24866,N_24983);
and UO_2314 (O_2314,N_24823,N_24983);
nor UO_2315 (O_2315,N_24853,N_24876);
nand UO_2316 (O_2316,N_24825,N_24834);
nor UO_2317 (O_2317,N_24978,N_24983);
nand UO_2318 (O_2318,N_24966,N_24976);
nand UO_2319 (O_2319,N_24960,N_24845);
nor UO_2320 (O_2320,N_24955,N_24985);
and UO_2321 (O_2321,N_24817,N_24911);
or UO_2322 (O_2322,N_24928,N_24984);
and UO_2323 (O_2323,N_24827,N_24893);
or UO_2324 (O_2324,N_24879,N_24885);
nand UO_2325 (O_2325,N_24863,N_24974);
nor UO_2326 (O_2326,N_24949,N_24883);
and UO_2327 (O_2327,N_24938,N_24812);
or UO_2328 (O_2328,N_24955,N_24881);
and UO_2329 (O_2329,N_24910,N_24944);
nor UO_2330 (O_2330,N_24945,N_24955);
nand UO_2331 (O_2331,N_24902,N_24946);
nor UO_2332 (O_2332,N_24951,N_24859);
nor UO_2333 (O_2333,N_24904,N_24951);
nand UO_2334 (O_2334,N_24861,N_24914);
nand UO_2335 (O_2335,N_24875,N_24908);
and UO_2336 (O_2336,N_24981,N_24815);
nand UO_2337 (O_2337,N_24864,N_24820);
or UO_2338 (O_2338,N_24961,N_24887);
or UO_2339 (O_2339,N_24971,N_24994);
or UO_2340 (O_2340,N_24897,N_24979);
and UO_2341 (O_2341,N_24907,N_24949);
or UO_2342 (O_2342,N_24831,N_24840);
nand UO_2343 (O_2343,N_24905,N_24966);
and UO_2344 (O_2344,N_24939,N_24904);
and UO_2345 (O_2345,N_24983,N_24881);
or UO_2346 (O_2346,N_24874,N_24942);
nor UO_2347 (O_2347,N_24846,N_24892);
and UO_2348 (O_2348,N_24821,N_24897);
nor UO_2349 (O_2349,N_24825,N_24883);
nor UO_2350 (O_2350,N_24900,N_24815);
nor UO_2351 (O_2351,N_24880,N_24853);
or UO_2352 (O_2352,N_24950,N_24920);
nor UO_2353 (O_2353,N_24945,N_24842);
nor UO_2354 (O_2354,N_24883,N_24841);
nand UO_2355 (O_2355,N_24827,N_24994);
and UO_2356 (O_2356,N_24831,N_24943);
and UO_2357 (O_2357,N_24932,N_24899);
or UO_2358 (O_2358,N_24978,N_24896);
nand UO_2359 (O_2359,N_24811,N_24867);
nor UO_2360 (O_2360,N_24933,N_24941);
and UO_2361 (O_2361,N_24957,N_24825);
and UO_2362 (O_2362,N_24952,N_24983);
and UO_2363 (O_2363,N_24845,N_24881);
xor UO_2364 (O_2364,N_24987,N_24842);
or UO_2365 (O_2365,N_24837,N_24964);
nor UO_2366 (O_2366,N_24958,N_24910);
nor UO_2367 (O_2367,N_24992,N_24913);
or UO_2368 (O_2368,N_24813,N_24819);
or UO_2369 (O_2369,N_24801,N_24947);
nor UO_2370 (O_2370,N_24903,N_24801);
and UO_2371 (O_2371,N_24850,N_24849);
and UO_2372 (O_2372,N_24808,N_24832);
nand UO_2373 (O_2373,N_24887,N_24979);
nor UO_2374 (O_2374,N_24808,N_24851);
and UO_2375 (O_2375,N_24951,N_24923);
or UO_2376 (O_2376,N_24807,N_24850);
nand UO_2377 (O_2377,N_24807,N_24896);
or UO_2378 (O_2378,N_24862,N_24868);
nor UO_2379 (O_2379,N_24872,N_24800);
and UO_2380 (O_2380,N_24947,N_24867);
or UO_2381 (O_2381,N_24922,N_24927);
nor UO_2382 (O_2382,N_24879,N_24875);
nand UO_2383 (O_2383,N_24974,N_24865);
or UO_2384 (O_2384,N_24894,N_24862);
nand UO_2385 (O_2385,N_24867,N_24885);
nor UO_2386 (O_2386,N_24882,N_24830);
nor UO_2387 (O_2387,N_24978,N_24973);
and UO_2388 (O_2388,N_24980,N_24945);
nor UO_2389 (O_2389,N_24876,N_24814);
and UO_2390 (O_2390,N_24908,N_24855);
nand UO_2391 (O_2391,N_24983,N_24998);
nand UO_2392 (O_2392,N_24917,N_24809);
nand UO_2393 (O_2393,N_24948,N_24945);
xor UO_2394 (O_2394,N_24997,N_24947);
or UO_2395 (O_2395,N_24806,N_24999);
or UO_2396 (O_2396,N_24887,N_24819);
nor UO_2397 (O_2397,N_24971,N_24892);
and UO_2398 (O_2398,N_24866,N_24849);
nor UO_2399 (O_2399,N_24979,N_24971);
nor UO_2400 (O_2400,N_24947,N_24830);
or UO_2401 (O_2401,N_24927,N_24805);
nand UO_2402 (O_2402,N_24812,N_24989);
nor UO_2403 (O_2403,N_24814,N_24857);
nand UO_2404 (O_2404,N_24836,N_24865);
nor UO_2405 (O_2405,N_24861,N_24808);
and UO_2406 (O_2406,N_24855,N_24992);
and UO_2407 (O_2407,N_24850,N_24954);
nor UO_2408 (O_2408,N_24985,N_24810);
and UO_2409 (O_2409,N_24802,N_24863);
and UO_2410 (O_2410,N_24979,N_24803);
and UO_2411 (O_2411,N_24856,N_24965);
and UO_2412 (O_2412,N_24978,N_24989);
nor UO_2413 (O_2413,N_24910,N_24912);
nand UO_2414 (O_2414,N_24955,N_24863);
nand UO_2415 (O_2415,N_24813,N_24931);
nor UO_2416 (O_2416,N_24929,N_24894);
and UO_2417 (O_2417,N_24911,N_24934);
nor UO_2418 (O_2418,N_24817,N_24954);
and UO_2419 (O_2419,N_24947,N_24907);
nor UO_2420 (O_2420,N_24909,N_24948);
nand UO_2421 (O_2421,N_24860,N_24898);
nor UO_2422 (O_2422,N_24882,N_24850);
nand UO_2423 (O_2423,N_24908,N_24889);
or UO_2424 (O_2424,N_24976,N_24937);
nand UO_2425 (O_2425,N_24866,N_24943);
or UO_2426 (O_2426,N_24894,N_24858);
nand UO_2427 (O_2427,N_24812,N_24887);
and UO_2428 (O_2428,N_24935,N_24953);
and UO_2429 (O_2429,N_24812,N_24944);
or UO_2430 (O_2430,N_24838,N_24905);
nand UO_2431 (O_2431,N_24892,N_24864);
or UO_2432 (O_2432,N_24906,N_24852);
and UO_2433 (O_2433,N_24839,N_24898);
and UO_2434 (O_2434,N_24848,N_24962);
nor UO_2435 (O_2435,N_24885,N_24930);
nor UO_2436 (O_2436,N_24985,N_24931);
or UO_2437 (O_2437,N_24909,N_24850);
nor UO_2438 (O_2438,N_24990,N_24858);
or UO_2439 (O_2439,N_24978,N_24835);
nand UO_2440 (O_2440,N_24997,N_24940);
nor UO_2441 (O_2441,N_24873,N_24917);
and UO_2442 (O_2442,N_24981,N_24908);
and UO_2443 (O_2443,N_24983,N_24870);
or UO_2444 (O_2444,N_24883,N_24814);
and UO_2445 (O_2445,N_24875,N_24980);
or UO_2446 (O_2446,N_24854,N_24968);
nor UO_2447 (O_2447,N_24951,N_24972);
nand UO_2448 (O_2448,N_24967,N_24801);
and UO_2449 (O_2449,N_24815,N_24800);
nand UO_2450 (O_2450,N_24872,N_24880);
nand UO_2451 (O_2451,N_24976,N_24902);
or UO_2452 (O_2452,N_24994,N_24811);
or UO_2453 (O_2453,N_24925,N_24845);
nand UO_2454 (O_2454,N_24819,N_24934);
nand UO_2455 (O_2455,N_24921,N_24961);
nand UO_2456 (O_2456,N_24927,N_24906);
nor UO_2457 (O_2457,N_24898,N_24874);
or UO_2458 (O_2458,N_24803,N_24918);
and UO_2459 (O_2459,N_24901,N_24816);
and UO_2460 (O_2460,N_24982,N_24876);
nand UO_2461 (O_2461,N_24928,N_24972);
nor UO_2462 (O_2462,N_24935,N_24831);
and UO_2463 (O_2463,N_24846,N_24887);
nand UO_2464 (O_2464,N_24967,N_24800);
and UO_2465 (O_2465,N_24857,N_24881);
nor UO_2466 (O_2466,N_24932,N_24985);
nor UO_2467 (O_2467,N_24971,N_24984);
nor UO_2468 (O_2468,N_24896,N_24962);
nand UO_2469 (O_2469,N_24807,N_24939);
or UO_2470 (O_2470,N_24971,N_24808);
nand UO_2471 (O_2471,N_24879,N_24801);
or UO_2472 (O_2472,N_24925,N_24838);
nand UO_2473 (O_2473,N_24992,N_24945);
or UO_2474 (O_2474,N_24914,N_24916);
and UO_2475 (O_2475,N_24980,N_24932);
or UO_2476 (O_2476,N_24871,N_24933);
nor UO_2477 (O_2477,N_24986,N_24984);
nand UO_2478 (O_2478,N_24968,N_24961);
nand UO_2479 (O_2479,N_24918,N_24910);
and UO_2480 (O_2480,N_24899,N_24832);
and UO_2481 (O_2481,N_24831,N_24882);
nand UO_2482 (O_2482,N_24901,N_24902);
nor UO_2483 (O_2483,N_24833,N_24836);
nor UO_2484 (O_2484,N_24905,N_24908);
or UO_2485 (O_2485,N_24819,N_24965);
or UO_2486 (O_2486,N_24884,N_24837);
nor UO_2487 (O_2487,N_24887,N_24917);
nand UO_2488 (O_2488,N_24994,N_24950);
nand UO_2489 (O_2489,N_24994,N_24887);
nor UO_2490 (O_2490,N_24923,N_24955);
nor UO_2491 (O_2491,N_24802,N_24813);
and UO_2492 (O_2492,N_24975,N_24953);
and UO_2493 (O_2493,N_24913,N_24863);
and UO_2494 (O_2494,N_24877,N_24965);
or UO_2495 (O_2495,N_24853,N_24869);
nand UO_2496 (O_2496,N_24980,N_24952);
or UO_2497 (O_2497,N_24824,N_24847);
or UO_2498 (O_2498,N_24889,N_24998);
nor UO_2499 (O_2499,N_24914,N_24995);
nand UO_2500 (O_2500,N_24803,N_24915);
nor UO_2501 (O_2501,N_24993,N_24964);
and UO_2502 (O_2502,N_24854,N_24988);
nor UO_2503 (O_2503,N_24806,N_24936);
nor UO_2504 (O_2504,N_24938,N_24901);
or UO_2505 (O_2505,N_24809,N_24993);
and UO_2506 (O_2506,N_24906,N_24915);
and UO_2507 (O_2507,N_24820,N_24894);
xnor UO_2508 (O_2508,N_24944,N_24870);
and UO_2509 (O_2509,N_24979,N_24981);
and UO_2510 (O_2510,N_24963,N_24927);
nor UO_2511 (O_2511,N_24893,N_24953);
nor UO_2512 (O_2512,N_24976,N_24806);
and UO_2513 (O_2513,N_24838,N_24989);
or UO_2514 (O_2514,N_24982,N_24942);
and UO_2515 (O_2515,N_24852,N_24981);
and UO_2516 (O_2516,N_24999,N_24885);
and UO_2517 (O_2517,N_24906,N_24817);
nor UO_2518 (O_2518,N_24934,N_24983);
nor UO_2519 (O_2519,N_24922,N_24852);
nor UO_2520 (O_2520,N_24965,N_24838);
and UO_2521 (O_2521,N_24982,N_24854);
or UO_2522 (O_2522,N_24942,N_24906);
nand UO_2523 (O_2523,N_24800,N_24973);
and UO_2524 (O_2524,N_24991,N_24847);
or UO_2525 (O_2525,N_24963,N_24954);
nor UO_2526 (O_2526,N_24843,N_24814);
and UO_2527 (O_2527,N_24826,N_24902);
nor UO_2528 (O_2528,N_24976,N_24867);
and UO_2529 (O_2529,N_24984,N_24936);
nor UO_2530 (O_2530,N_24815,N_24987);
nor UO_2531 (O_2531,N_24860,N_24897);
or UO_2532 (O_2532,N_24850,N_24876);
nand UO_2533 (O_2533,N_24931,N_24928);
nor UO_2534 (O_2534,N_24888,N_24800);
and UO_2535 (O_2535,N_24984,N_24876);
nor UO_2536 (O_2536,N_24837,N_24938);
or UO_2537 (O_2537,N_24890,N_24970);
nand UO_2538 (O_2538,N_24816,N_24833);
nor UO_2539 (O_2539,N_24871,N_24907);
and UO_2540 (O_2540,N_24883,N_24920);
nor UO_2541 (O_2541,N_24933,N_24975);
nand UO_2542 (O_2542,N_24843,N_24960);
nor UO_2543 (O_2543,N_24990,N_24901);
or UO_2544 (O_2544,N_24991,N_24815);
or UO_2545 (O_2545,N_24827,N_24914);
nand UO_2546 (O_2546,N_24958,N_24806);
nand UO_2547 (O_2547,N_24952,N_24806);
nor UO_2548 (O_2548,N_24919,N_24994);
or UO_2549 (O_2549,N_24933,N_24924);
nor UO_2550 (O_2550,N_24925,N_24861);
and UO_2551 (O_2551,N_24856,N_24839);
or UO_2552 (O_2552,N_24893,N_24897);
nand UO_2553 (O_2553,N_24872,N_24822);
nand UO_2554 (O_2554,N_24987,N_24857);
and UO_2555 (O_2555,N_24835,N_24859);
nand UO_2556 (O_2556,N_24825,N_24997);
nor UO_2557 (O_2557,N_24892,N_24806);
or UO_2558 (O_2558,N_24946,N_24823);
nor UO_2559 (O_2559,N_24939,N_24960);
nand UO_2560 (O_2560,N_24982,N_24857);
and UO_2561 (O_2561,N_24931,N_24829);
and UO_2562 (O_2562,N_24909,N_24864);
and UO_2563 (O_2563,N_24865,N_24983);
nand UO_2564 (O_2564,N_24844,N_24917);
or UO_2565 (O_2565,N_24850,N_24886);
and UO_2566 (O_2566,N_24983,N_24817);
or UO_2567 (O_2567,N_24913,N_24985);
nand UO_2568 (O_2568,N_24943,N_24925);
nor UO_2569 (O_2569,N_24883,N_24914);
or UO_2570 (O_2570,N_24974,N_24921);
nand UO_2571 (O_2571,N_24844,N_24929);
or UO_2572 (O_2572,N_24818,N_24802);
nand UO_2573 (O_2573,N_24910,N_24808);
nor UO_2574 (O_2574,N_24882,N_24983);
nor UO_2575 (O_2575,N_24823,N_24850);
and UO_2576 (O_2576,N_24898,N_24864);
nor UO_2577 (O_2577,N_24882,N_24846);
nor UO_2578 (O_2578,N_24944,N_24808);
xnor UO_2579 (O_2579,N_24902,N_24997);
nand UO_2580 (O_2580,N_24838,N_24996);
nand UO_2581 (O_2581,N_24823,N_24838);
nand UO_2582 (O_2582,N_24804,N_24838);
or UO_2583 (O_2583,N_24821,N_24818);
or UO_2584 (O_2584,N_24949,N_24993);
or UO_2585 (O_2585,N_24807,N_24981);
nand UO_2586 (O_2586,N_24926,N_24832);
nand UO_2587 (O_2587,N_24969,N_24820);
and UO_2588 (O_2588,N_24972,N_24908);
nor UO_2589 (O_2589,N_24929,N_24930);
or UO_2590 (O_2590,N_24842,N_24819);
nor UO_2591 (O_2591,N_24851,N_24974);
nand UO_2592 (O_2592,N_24849,N_24823);
nand UO_2593 (O_2593,N_24814,N_24826);
nand UO_2594 (O_2594,N_24826,N_24841);
nor UO_2595 (O_2595,N_24877,N_24852);
nand UO_2596 (O_2596,N_24910,N_24806);
nand UO_2597 (O_2597,N_24921,N_24985);
nor UO_2598 (O_2598,N_24901,N_24995);
and UO_2599 (O_2599,N_24870,N_24883);
nand UO_2600 (O_2600,N_24915,N_24916);
or UO_2601 (O_2601,N_24810,N_24816);
and UO_2602 (O_2602,N_24922,N_24990);
nor UO_2603 (O_2603,N_24986,N_24948);
nand UO_2604 (O_2604,N_24905,N_24918);
or UO_2605 (O_2605,N_24867,N_24985);
nand UO_2606 (O_2606,N_24808,N_24989);
or UO_2607 (O_2607,N_24892,N_24908);
and UO_2608 (O_2608,N_24916,N_24832);
and UO_2609 (O_2609,N_24847,N_24987);
or UO_2610 (O_2610,N_24990,N_24993);
and UO_2611 (O_2611,N_24931,N_24878);
nor UO_2612 (O_2612,N_24822,N_24963);
nand UO_2613 (O_2613,N_24885,N_24913);
nand UO_2614 (O_2614,N_24830,N_24824);
and UO_2615 (O_2615,N_24967,N_24956);
nand UO_2616 (O_2616,N_24837,N_24830);
and UO_2617 (O_2617,N_24928,N_24980);
nor UO_2618 (O_2618,N_24887,N_24850);
and UO_2619 (O_2619,N_24918,N_24826);
or UO_2620 (O_2620,N_24924,N_24982);
and UO_2621 (O_2621,N_24817,N_24859);
nor UO_2622 (O_2622,N_24864,N_24968);
nand UO_2623 (O_2623,N_24906,N_24961);
nand UO_2624 (O_2624,N_24899,N_24924);
or UO_2625 (O_2625,N_24810,N_24809);
or UO_2626 (O_2626,N_24946,N_24918);
nand UO_2627 (O_2627,N_24899,N_24825);
nand UO_2628 (O_2628,N_24997,N_24901);
and UO_2629 (O_2629,N_24877,N_24872);
nand UO_2630 (O_2630,N_24874,N_24831);
nand UO_2631 (O_2631,N_24968,N_24837);
nor UO_2632 (O_2632,N_24815,N_24899);
nand UO_2633 (O_2633,N_24828,N_24833);
nand UO_2634 (O_2634,N_24983,N_24935);
nor UO_2635 (O_2635,N_24918,N_24835);
and UO_2636 (O_2636,N_24977,N_24859);
or UO_2637 (O_2637,N_24840,N_24865);
nor UO_2638 (O_2638,N_24886,N_24992);
and UO_2639 (O_2639,N_24950,N_24813);
or UO_2640 (O_2640,N_24885,N_24898);
nor UO_2641 (O_2641,N_24901,N_24957);
nor UO_2642 (O_2642,N_24859,N_24877);
and UO_2643 (O_2643,N_24935,N_24998);
and UO_2644 (O_2644,N_24802,N_24998);
and UO_2645 (O_2645,N_24811,N_24898);
nand UO_2646 (O_2646,N_24986,N_24870);
or UO_2647 (O_2647,N_24806,N_24849);
nand UO_2648 (O_2648,N_24920,N_24849);
and UO_2649 (O_2649,N_24992,N_24849);
nor UO_2650 (O_2650,N_24854,N_24914);
nand UO_2651 (O_2651,N_24985,N_24837);
or UO_2652 (O_2652,N_24949,N_24856);
nand UO_2653 (O_2653,N_24963,N_24944);
nor UO_2654 (O_2654,N_24888,N_24961);
nand UO_2655 (O_2655,N_24811,N_24931);
nor UO_2656 (O_2656,N_24998,N_24915);
or UO_2657 (O_2657,N_24822,N_24994);
nand UO_2658 (O_2658,N_24960,N_24968);
nand UO_2659 (O_2659,N_24889,N_24845);
and UO_2660 (O_2660,N_24815,N_24929);
nand UO_2661 (O_2661,N_24921,N_24847);
nor UO_2662 (O_2662,N_24937,N_24850);
and UO_2663 (O_2663,N_24887,N_24977);
nor UO_2664 (O_2664,N_24842,N_24882);
or UO_2665 (O_2665,N_24864,N_24967);
or UO_2666 (O_2666,N_24933,N_24952);
nand UO_2667 (O_2667,N_24885,N_24894);
or UO_2668 (O_2668,N_24973,N_24810);
and UO_2669 (O_2669,N_24852,N_24931);
and UO_2670 (O_2670,N_24926,N_24922);
nand UO_2671 (O_2671,N_24873,N_24960);
nor UO_2672 (O_2672,N_24847,N_24925);
nand UO_2673 (O_2673,N_24913,N_24915);
nand UO_2674 (O_2674,N_24937,N_24971);
or UO_2675 (O_2675,N_24816,N_24910);
and UO_2676 (O_2676,N_24838,N_24984);
or UO_2677 (O_2677,N_24965,N_24975);
nand UO_2678 (O_2678,N_24999,N_24976);
nand UO_2679 (O_2679,N_24965,N_24935);
and UO_2680 (O_2680,N_24905,N_24903);
and UO_2681 (O_2681,N_24841,N_24965);
or UO_2682 (O_2682,N_24925,N_24962);
nand UO_2683 (O_2683,N_24979,N_24925);
nor UO_2684 (O_2684,N_24925,N_24912);
or UO_2685 (O_2685,N_24863,N_24948);
nor UO_2686 (O_2686,N_24953,N_24891);
and UO_2687 (O_2687,N_24907,N_24928);
or UO_2688 (O_2688,N_24912,N_24908);
nor UO_2689 (O_2689,N_24814,N_24998);
and UO_2690 (O_2690,N_24845,N_24989);
nor UO_2691 (O_2691,N_24830,N_24984);
xnor UO_2692 (O_2692,N_24931,N_24847);
nand UO_2693 (O_2693,N_24853,N_24974);
and UO_2694 (O_2694,N_24875,N_24809);
nor UO_2695 (O_2695,N_24817,N_24830);
or UO_2696 (O_2696,N_24823,N_24888);
nor UO_2697 (O_2697,N_24841,N_24955);
nor UO_2698 (O_2698,N_24955,N_24932);
nand UO_2699 (O_2699,N_24972,N_24956);
nand UO_2700 (O_2700,N_24916,N_24834);
or UO_2701 (O_2701,N_24924,N_24946);
xor UO_2702 (O_2702,N_24859,N_24862);
and UO_2703 (O_2703,N_24981,N_24890);
or UO_2704 (O_2704,N_24954,N_24884);
nand UO_2705 (O_2705,N_24971,N_24975);
nand UO_2706 (O_2706,N_24979,N_24875);
or UO_2707 (O_2707,N_24901,N_24993);
nor UO_2708 (O_2708,N_24933,N_24894);
or UO_2709 (O_2709,N_24926,N_24940);
nor UO_2710 (O_2710,N_24899,N_24868);
or UO_2711 (O_2711,N_24959,N_24840);
or UO_2712 (O_2712,N_24858,N_24841);
nand UO_2713 (O_2713,N_24947,N_24899);
or UO_2714 (O_2714,N_24888,N_24818);
or UO_2715 (O_2715,N_24876,N_24886);
and UO_2716 (O_2716,N_24935,N_24918);
nor UO_2717 (O_2717,N_24869,N_24808);
or UO_2718 (O_2718,N_24950,N_24810);
nor UO_2719 (O_2719,N_24974,N_24814);
nand UO_2720 (O_2720,N_24993,N_24829);
nor UO_2721 (O_2721,N_24926,N_24826);
nor UO_2722 (O_2722,N_24916,N_24837);
nor UO_2723 (O_2723,N_24990,N_24859);
and UO_2724 (O_2724,N_24814,N_24875);
and UO_2725 (O_2725,N_24884,N_24819);
or UO_2726 (O_2726,N_24888,N_24920);
and UO_2727 (O_2727,N_24826,N_24821);
and UO_2728 (O_2728,N_24860,N_24894);
nor UO_2729 (O_2729,N_24900,N_24871);
nor UO_2730 (O_2730,N_24932,N_24800);
nand UO_2731 (O_2731,N_24958,N_24966);
or UO_2732 (O_2732,N_24911,N_24856);
and UO_2733 (O_2733,N_24992,N_24952);
nand UO_2734 (O_2734,N_24915,N_24836);
or UO_2735 (O_2735,N_24902,N_24897);
nand UO_2736 (O_2736,N_24884,N_24934);
nor UO_2737 (O_2737,N_24986,N_24950);
nor UO_2738 (O_2738,N_24821,N_24997);
nor UO_2739 (O_2739,N_24941,N_24822);
xor UO_2740 (O_2740,N_24932,N_24841);
nand UO_2741 (O_2741,N_24843,N_24934);
nand UO_2742 (O_2742,N_24978,N_24867);
nor UO_2743 (O_2743,N_24957,N_24950);
and UO_2744 (O_2744,N_24959,N_24851);
nand UO_2745 (O_2745,N_24934,N_24900);
nand UO_2746 (O_2746,N_24967,N_24847);
and UO_2747 (O_2747,N_24835,N_24908);
and UO_2748 (O_2748,N_24933,N_24845);
nand UO_2749 (O_2749,N_24866,N_24876);
or UO_2750 (O_2750,N_24984,N_24933);
or UO_2751 (O_2751,N_24842,N_24934);
and UO_2752 (O_2752,N_24873,N_24833);
or UO_2753 (O_2753,N_24951,N_24827);
nor UO_2754 (O_2754,N_24843,N_24836);
and UO_2755 (O_2755,N_24826,N_24965);
nand UO_2756 (O_2756,N_24914,N_24886);
or UO_2757 (O_2757,N_24954,N_24865);
and UO_2758 (O_2758,N_24921,N_24843);
and UO_2759 (O_2759,N_24934,N_24968);
nand UO_2760 (O_2760,N_24980,N_24878);
nor UO_2761 (O_2761,N_24917,N_24836);
or UO_2762 (O_2762,N_24859,N_24901);
or UO_2763 (O_2763,N_24961,N_24981);
and UO_2764 (O_2764,N_24830,N_24805);
and UO_2765 (O_2765,N_24914,N_24879);
and UO_2766 (O_2766,N_24928,N_24813);
nand UO_2767 (O_2767,N_24848,N_24951);
or UO_2768 (O_2768,N_24844,N_24894);
and UO_2769 (O_2769,N_24971,N_24992);
nor UO_2770 (O_2770,N_24896,N_24981);
nor UO_2771 (O_2771,N_24897,N_24859);
and UO_2772 (O_2772,N_24866,N_24822);
nand UO_2773 (O_2773,N_24828,N_24989);
and UO_2774 (O_2774,N_24848,N_24807);
and UO_2775 (O_2775,N_24874,N_24888);
nor UO_2776 (O_2776,N_24984,N_24950);
or UO_2777 (O_2777,N_24918,N_24932);
and UO_2778 (O_2778,N_24863,N_24900);
nor UO_2779 (O_2779,N_24988,N_24812);
or UO_2780 (O_2780,N_24839,N_24930);
nor UO_2781 (O_2781,N_24986,N_24951);
and UO_2782 (O_2782,N_24952,N_24896);
nand UO_2783 (O_2783,N_24990,N_24839);
nor UO_2784 (O_2784,N_24894,N_24919);
nand UO_2785 (O_2785,N_24994,N_24982);
nand UO_2786 (O_2786,N_24827,N_24824);
and UO_2787 (O_2787,N_24835,N_24943);
nand UO_2788 (O_2788,N_24884,N_24942);
and UO_2789 (O_2789,N_24836,N_24944);
or UO_2790 (O_2790,N_24852,N_24962);
and UO_2791 (O_2791,N_24915,N_24984);
nor UO_2792 (O_2792,N_24859,N_24910);
nand UO_2793 (O_2793,N_24849,N_24887);
or UO_2794 (O_2794,N_24941,N_24844);
and UO_2795 (O_2795,N_24953,N_24992);
nand UO_2796 (O_2796,N_24851,N_24932);
nand UO_2797 (O_2797,N_24876,N_24900);
nor UO_2798 (O_2798,N_24844,N_24911);
or UO_2799 (O_2799,N_24826,N_24972);
nand UO_2800 (O_2800,N_24880,N_24952);
nor UO_2801 (O_2801,N_24901,N_24828);
nor UO_2802 (O_2802,N_24936,N_24891);
and UO_2803 (O_2803,N_24942,N_24961);
or UO_2804 (O_2804,N_24814,N_24825);
or UO_2805 (O_2805,N_24928,N_24989);
nand UO_2806 (O_2806,N_24992,N_24933);
or UO_2807 (O_2807,N_24989,N_24948);
nand UO_2808 (O_2808,N_24893,N_24899);
nand UO_2809 (O_2809,N_24988,N_24924);
nor UO_2810 (O_2810,N_24929,N_24853);
and UO_2811 (O_2811,N_24877,N_24876);
nor UO_2812 (O_2812,N_24952,N_24882);
nand UO_2813 (O_2813,N_24873,N_24909);
and UO_2814 (O_2814,N_24900,N_24913);
nor UO_2815 (O_2815,N_24927,N_24812);
nand UO_2816 (O_2816,N_24968,N_24829);
and UO_2817 (O_2817,N_24943,N_24991);
and UO_2818 (O_2818,N_24867,N_24842);
or UO_2819 (O_2819,N_24982,N_24805);
nand UO_2820 (O_2820,N_24839,N_24976);
nor UO_2821 (O_2821,N_24938,N_24919);
and UO_2822 (O_2822,N_24997,N_24845);
nand UO_2823 (O_2823,N_24966,N_24853);
or UO_2824 (O_2824,N_24968,N_24931);
nand UO_2825 (O_2825,N_24813,N_24847);
or UO_2826 (O_2826,N_24829,N_24916);
nor UO_2827 (O_2827,N_24960,N_24833);
and UO_2828 (O_2828,N_24917,N_24843);
and UO_2829 (O_2829,N_24880,N_24969);
or UO_2830 (O_2830,N_24878,N_24826);
nand UO_2831 (O_2831,N_24881,N_24839);
and UO_2832 (O_2832,N_24961,N_24839);
or UO_2833 (O_2833,N_24913,N_24924);
and UO_2834 (O_2834,N_24801,N_24913);
xnor UO_2835 (O_2835,N_24949,N_24921);
nor UO_2836 (O_2836,N_24801,N_24881);
nand UO_2837 (O_2837,N_24941,N_24952);
nand UO_2838 (O_2838,N_24879,N_24838);
and UO_2839 (O_2839,N_24803,N_24869);
nand UO_2840 (O_2840,N_24861,N_24848);
nor UO_2841 (O_2841,N_24899,N_24931);
nand UO_2842 (O_2842,N_24842,N_24963);
and UO_2843 (O_2843,N_24861,N_24802);
and UO_2844 (O_2844,N_24880,N_24851);
nand UO_2845 (O_2845,N_24945,N_24957);
nor UO_2846 (O_2846,N_24973,N_24872);
and UO_2847 (O_2847,N_24873,N_24990);
or UO_2848 (O_2848,N_24883,N_24909);
and UO_2849 (O_2849,N_24995,N_24866);
or UO_2850 (O_2850,N_24930,N_24980);
and UO_2851 (O_2851,N_24923,N_24911);
or UO_2852 (O_2852,N_24887,N_24841);
nor UO_2853 (O_2853,N_24815,N_24912);
nand UO_2854 (O_2854,N_24814,N_24958);
and UO_2855 (O_2855,N_24817,N_24933);
nand UO_2856 (O_2856,N_24811,N_24844);
and UO_2857 (O_2857,N_24822,N_24830);
or UO_2858 (O_2858,N_24815,N_24887);
nor UO_2859 (O_2859,N_24907,N_24934);
nor UO_2860 (O_2860,N_24879,N_24871);
or UO_2861 (O_2861,N_24968,N_24824);
nand UO_2862 (O_2862,N_24818,N_24994);
nand UO_2863 (O_2863,N_24854,N_24940);
or UO_2864 (O_2864,N_24811,N_24988);
nand UO_2865 (O_2865,N_24871,N_24942);
and UO_2866 (O_2866,N_24860,N_24907);
and UO_2867 (O_2867,N_24806,N_24987);
or UO_2868 (O_2868,N_24853,N_24845);
nand UO_2869 (O_2869,N_24916,N_24946);
and UO_2870 (O_2870,N_24869,N_24987);
nor UO_2871 (O_2871,N_24873,N_24804);
or UO_2872 (O_2872,N_24817,N_24879);
nor UO_2873 (O_2873,N_24935,N_24969);
nor UO_2874 (O_2874,N_24855,N_24804);
or UO_2875 (O_2875,N_24978,N_24865);
or UO_2876 (O_2876,N_24925,N_24917);
or UO_2877 (O_2877,N_24988,N_24963);
or UO_2878 (O_2878,N_24801,N_24823);
nand UO_2879 (O_2879,N_24994,N_24970);
and UO_2880 (O_2880,N_24808,N_24873);
or UO_2881 (O_2881,N_24888,N_24904);
and UO_2882 (O_2882,N_24915,N_24926);
nand UO_2883 (O_2883,N_24810,N_24811);
xnor UO_2884 (O_2884,N_24972,N_24893);
and UO_2885 (O_2885,N_24803,N_24879);
or UO_2886 (O_2886,N_24994,N_24944);
nor UO_2887 (O_2887,N_24949,N_24803);
nand UO_2888 (O_2888,N_24839,N_24942);
and UO_2889 (O_2889,N_24808,N_24901);
or UO_2890 (O_2890,N_24973,N_24855);
and UO_2891 (O_2891,N_24940,N_24888);
and UO_2892 (O_2892,N_24994,N_24864);
nand UO_2893 (O_2893,N_24908,N_24974);
nand UO_2894 (O_2894,N_24864,N_24844);
or UO_2895 (O_2895,N_24977,N_24966);
nor UO_2896 (O_2896,N_24883,N_24806);
nand UO_2897 (O_2897,N_24921,N_24994);
nor UO_2898 (O_2898,N_24892,N_24828);
nor UO_2899 (O_2899,N_24900,N_24976);
nand UO_2900 (O_2900,N_24940,N_24957);
xor UO_2901 (O_2901,N_24887,N_24853);
or UO_2902 (O_2902,N_24809,N_24951);
nand UO_2903 (O_2903,N_24840,N_24914);
and UO_2904 (O_2904,N_24815,N_24942);
or UO_2905 (O_2905,N_24984,N_24932);
nand UO_2906 (O_2906,N_24849,N_24931);
nor UO_2907 (O_2907,N_24937,N_24929);
and UO_2908 (O_2908,N_24942,N_24954);
and UO_2909 (O_2909,N_24998,N_24974);
nand UO_2910 (O_2910,N_24824,N_24938);
and UO_2911 (O_2911,N_24913,N_24811);
or UO_2912 (O_2912,N_24928,N_24866);
nor UO_2913 (O_2913,N_24865,N_24979);
and UO_2914 (O_2914,N_24994,N_24928);
nor UO_2915 (O_2915,N_24905,N_24889);
or UO_2916 (O_2916,N_24891,N_24878);
or UO_2917 (O_2917,N_24891,N_24813);
nand UO_2918 (O_2918,N_24927,N_24816);
and UO_2919 (O_2919,N_24839,N_24804);
and UO_2920 (O_2920,N_24801,N_24962);
and UO_2921 (O_2921,N_24999,N_24900);
or UO_2922 (O_2922,N_24834,N_24831);
or UO_2923 (O_2923,N_24892,N_24854);
or UO_2924 (O_2924,N_24887,N_24960);
and UO_2925 (O_2925,N_24868,N_24900);
nand UO_2926 (O_2926,N_24995,N_24823);
nand UO_2927 (O_2927,N_24815,N_24853);
nand UO_2928 (O_2928,N_24837,N_24820);
and UO_2929 (O_2929,N_24867,N_24938);
nor UO_2930 (O_2930,N_24830,N_24875);
or UO_2931 (O_2931,N_24941,N_24959);
nor UO_2932 (O_2932,N_24879,N_24950);
nand UO_2933 (O_2933,N_24851,N_24942);
nor UO_2934 (O_2934,N_24811,N_24955);
nor UO_2935 (O_2935,N_24894,N_24942);
or UO_2936 (O_2936,N_24952,N_24912);
or UO_2937 (O_2937,N_24886,N_24999);
nor UO_2938 (O_2938,N_24908,N_24923);
or UO_2939 (O_2939,N_24954,N_24846);
nor UO_2940 (O_2940,N_24881,N_24843);
nor UO_2941 (O_2941,N_24921,N_24986);
and UO_2942 (O_2942,N_24824,N_24971);
or UO_2943 (O_2943,N_24948,N_24983);
or UO_2944 (O_2944,N_24958,N_24865);
or UO_2945 (O_2945,N_24989,N_24936);
or UO_2946 (O_2946,N_24864,N_24955);
and UO_2947 (O_2947,N_24915,N_24880);
or UO_2948 (O_2948,N_24865,N_24945);
nand UO_2949 (O_2949,N_24858,N_24979);
and UO_2950 (O_2950,N_24860,N_24981);
xnor UO_2951 (O_2951,N_24854,N_24917);
xnor UO_2952 (O_2952,N_24805,N_24968);
and UO_2953 (O_2953,N_24871,N_24998);
nand UO_2954 (O_2954,N_24868,N_24828);
or UO_2955 (O_2955,N_24876,N_24825);
or UO_2956 (O_2956,N_24914,N_24891);
or UO_2957 (O_2957,N_24873,N_24992);
nor UO_2958 (O_2958,N_24849,N_24908);
or UO_2959 (O_2959,N_24941,N_24966);
nor UO_2960 (O_2960,N_24800,N_24904);
nand UO_2961 (O_2961,N_24897,N_24812);
nor UO_2962 (O_2962,N_24842,N_24865);
or UO_2963 (O_2963,N_24844,N_24907);
nor UO_2964 (O_2964,N_24982,N_24851);
and UO_2965 (O_2965,N_24945,N_24804);
and UO_2966 (O_2966,N_24849,N_24981);
nor UO_2967 (O_2967,N_24829,N_24813);
nor UO_2968 (O_2968,N_24960,N_24821);
and UO_2969 (O_2969,N_24966,N_24933);
or UO_2970 (O_2970,N_24811,N_24915);
and UO_2971 (O_2971,N_24822,N_24961);
nor UO_2972 (O_2972,N_24902,N_24809);
and UO_2973 (O_2973,N_24910,N_24971);
nand UO_2974 (O_2974,N_24826,N_24800);
or UO_2975 (O_2975,N_24930,N_24833);
nor UO_2976 (O_2976,N_24842,N_24913);
or UO_2977 (O_2977,N_24914,N_24924);
or UO_2978 (O_2978,N_24941,N_24823);
or UO_2979 (O_2979,N_24930,N_24846);
and UO_2980 (O_2980,N_24954,N_24971);
nor UO_2981 (O_2981,N_24907,N_24919);
and UO_2982 (O_2982,N_24909,N_24894);
nand UO_2983 (O_2983,N_24807,N_24863);
nand UO_2984 (O_2984,N_24986,N_24954);
nand UO_2985 (O_2985,N_24901,N_24939);
or UO_2986 (O_2986,N_24900,N_24928);
or UO_2987 (O_2987,N_24924,N_24910);
and UO_2988 (O_2988,N_24850,N_24993);
and UO_2989 (O_2989,N_24995,N_24868);
and UO_2990 (O_2990,N_24990,N_24834);
nor UO_2991 (O_2991,N_24845,N_24826);
and UO_2992 (O_2992,N_24858,N_24869);
or UO_2993 (O_2993,N_24873,N_24915);
nor UO_2994 (O_2994,N_24961,N_24875);
and UO_2995 (O_2995,N_24940,N_24971);
nand UO_2996 (O_2996,N_24933,N_24851);
or UO_2997 (O_2997,N_24961,N_24999);
nand UO_2998 (O_2998,N_24882,N_24918);
and UO_2999 (O_2999,N_24808,N_24918);
endmodule