module basic_500_3000_500_6_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_223,In_123);
or U1 (N_1,In_232,In_91);
xnor U2 (N_2,In_310,In_417);
nand U3 (N_3,In_170,In_155);
and U4 (N_4,In_202,In_243);
and U5 (N_5,In_88,In_346);
nand U6 (N_6,In_372,In_378);
or U7 (N_7,In_463,In_423);
or U8 (N_8,In_366,In_422);
nor U9 (N_9,In_278,In_95);
or U10 (N_10,In_191,In_420);
nor U11 (N_11,In_322,In_269);
nor U12 (N_12,In_20,In_312);
xor U13 (N_13,In_4,In_460);
nor U14 (N_14,In_115,In_31);
xor U15 (N_15,In_410,In_194);
nor U16 (N_16,In_206,In_279);
and U17 (N_17,In_8,In_288);
or U18 (N_18,In_424,In_40);
nand U19 (N_19,In_486,In_135);
nand U20 (N_20,In_474,In_455);
or U21 (N_21,In_401,In_85);
nand U22 (N_22,In_488,In_112);
nand U23 (N_23,In_161,In_497);
nand U24 (N_24,In_73,In_162);
nor U25 (N_25,In_197,In_458);
and U26 (N_26,In_5,In_81);
nand U27 (N_27,In_14,In_52);
nor U28 (N_28,In_308,In_53);
and U29 (N_29,In_114,In_106);
and U30 (N_30,In_76,In_82);
and U31 (N_31,In_55,In_323);
or U32 (N_32,In_61,In_381);
or U33 (N_33,In_118,In_362);
nand U34 (N_34,In_208,In_41);
and U35 (N_35,In_129,In_432);
nand U36 (N_36,In_485,In_169);
or U37 (N_37,In_49,In_148);
and U38 (N_38,In_414,In_176);
nand U39 (N_39,In_304,In_297);
nand U40 (N_40,In_359,In_478);
nand U41 (N_41,In_231,In_200);
nand U42 (N_42,In_350,In_219);
and U43 (N_43,In_303,In_18);
nor U44 (N_44,In_395,In_75);
nor U45 (N_45,In_180,In_425);
and U46 (N_46,In_94,In_442);
nor U47 (N_47,In_30,In_2);
or U48 (N_48,In_313,In_47);
nand U49 (N_49,In_140,In_15);
and U50 (N_50,In_367,In_476);
nand U51 (N_51,In_63,In_168);
nand U52 (N_52,In_260,In_29);
or U53 (N_53,In_457,In_183);
and U54 (N_54,In_364,In_363);
or U55 (N_55,In_182,In_96);
and U56 (N_56,In_371,In_499);
and U57 (N_57,In_327,In_70);
and U58 (N_58,In_396,In_229);
nand U59 (N_59,In_392,In_452);
nand U60 (N_60,In_258,In_245);
nand U61 (N_61,In_300,In_498);
nor U62 (N_62,In_104,In_296);
and U63 (N_63,In_110,In_445);
or U64 (N_64,In_431,In_128);
or U65 (N_65,In_102,In_7);
nand U66 (N_66,In_494,In_482);
nand U67 (N_67,In_286,In_351);
and U68 (N_68,In_496,In_37);
and U69 (N_69,In_309,In_149);
or U70 (N_70,In_121,In_385);
nand U71 (N_71,In_105,In_305);
or U72 (N_72,In_240,In_68);
nor U73 (N_73,In_218,In_487);
nand U74 (N_74,In_133,In_58);
nand U75 (N_75,In_124,In_204);
nand U76 (N_76,In_154,In_316);
or U77 (N_77,In_236,In_60);
nor U78 (N_78,In_145,In_132);
nor U79 (N_79,In_172,In_314);
nand U80 (N_80,In_383,In_326);
nor U81 (N_81,In_440,In_416);
or U82 (N_82,In_59,In_108);
or U83 (N_83,In_150,In_376);
or U84 (N_84,In_292,In_160);
and U85 (N_85,In_280,In_263);
nor U86 (N_86,In_244,In_97);
nor U87 (N_87,In_380,In_146);
and U88 (N_88,In_62,In_107);
nand U89 (N_89,In_449,In_436);
nor U90 (N_90,In_181,In_484);
and U91 (N_91,In_329,In_214);
nand U92 (N_92,In_144,In_227);
nand U93 (N_93,In_131,In_470);
nor U94 (N_94,In_283,In_415);
nor U95 (N_95,In_369,In_464);
nor U96 (N_96,In_492,In_45);
nor U97 (N_97,In_36,In_337);
xnor U98 (N_98,In_64,In_357);
nor U99 (N_99,In_382,In_256);
nand U100 (N_100,In_472,In_66);
nand U101 (N_101,In_237,In_84);
or U102 (N_102,In_101,In_103);
or U103 (N_103,In_126,In_315);
or U104 (N_104,In_490,In_165);
and U105 (N_105,In_265,In_319);
or U106 (N_106,In_468,In_287);
nor U107 (N_107,In_198,In_109);
nand U108 (N_108,In_389,In_35);
nor U109 (N_109,In_259,In_50);
nor U110 (N_110,In_282,In_354);
nor U111 (N_111,In_421,In_273);
or U112 (N_112,In_480,In_388);
and U113 (N_113,In_352,In_17);
nand U114 (N_114,In_409,In_454);
nor U115 (N_115,In_276,In_374);
or U116 (N_116,In_311,In_467);
nor U117 (N_117,In_67,In_407);
or U118 (N_118,In_461,In_493);
nand U119 (N_119,In_138,In_368);
nand U120 (N_120,In_307,In_111);
nor U121 (N_121,In_321,In_384);
nor U122 (N_122,In_57,In_268);
or U123 (N_123,In_437,In_471);
nor U124 (N_124,In_80,In_173);
nor U125 (N_125,In_157,In_167);
nor U126 (N_126,In_334,In_298);
nand U127 (N_127,In_419,In_281);
nor U128 (N_128,In_89,In_216);
nand U129 (N_129,In_171,In_345);
and U130 (N_130,In_90,In_349);
nand U131 (N_131,In_195,In_397);
or U132 (N_132,In_390,In_257);
and U133 (N_133,In_113,In_215);
nor U134 (N_134,In_158,In_86);
nor U135 (N_135,In_0,In_402);
and U136 (N_136,In_32,In_491);
nand U137 (N_137,In_358,In_187);
nor U138 (N_138,In_142,In_74);
nand U139 (N_139,In_430,In_174);
and U140 (N_140,In_250,In_356);
or U141 (N_141,In_246,In_394);
and U142 (N_142,In_324,In_83);
nand U143 (N_143,In_21,In_427);
nand U144 (N_144,In_209,In_295);
nand U145 (N_145,In_185,In_164);
nor U146 (N_146,In_239,In_355);
and U147 (N_147,In_275,In_317);
nand U148 (N_148,In_248,In_344);
nand U149 (N_149,In_247,In_27);
nor U150 (N_150,In_348,In_28);
and U151 (N_151,In_153,In_23);
nor U152 (N_152,In_404,In_365);
and U153 (N_153,In_353,In_56);
nand U154 (N_154,In_117,In_360);
or U155 (N_155,In_361,In_233);
nand U156 (N_156,In_48,In_495);
or U157 (N_157,In_179,In_411);
or U158 (N_158,In_433,In_152);
nand U159 (N_159,In_137,In_373);
and U160 (N_160,In_143,In_72);
or U161 (N_161,In_251,In_221);
or U162 (N_162,In_93,In_222);
and U163 (N_163,In_177,In_147);
nor U164 (N_164,In_299,In_207);
xor U165 (N_165,In_253,In_189);
or U166 (N_166,In_405,In_412);
xor U167 (N_167,In_16,In_429);
nor U168 (N_168,In_193,In_98);
nor U169 (N_169,In_139,In_1);
and U170 (N_170,In_291,In_241);
or U171 (N_171,In_386,In_125);
or U172 (N_172,In_343,In_220);
or U173 (N_173,In_406,In_87);
or U174 (N_174,In_267,In_479);
or U175 (N_175,In_199,In_483);
and U176 (N_176,In_42,In_100);
and U177 (N_177,In_272,In_264);
and U178 (N_178,In_130,In_12);
or U179 (N_179,In_441,In_330);
or U180 (N_180,In_332,In_78);
and U181 (N_181,In_266,In_447);
nand U182 (N_182,In_271,In_448);
or U183 (N_183,In_234,In_6);
or U184 (N_184,In_116,In_306);
and U185 (N_185,In_331,In_39);
nand U186 (N_186,In_341,In_134);
and U187 (N_187,In_285,In_418);
nand U188 (N_188,In_156,In_453);
and U189 (N_189,In_99,In_456);
nand U190 (N_190,In_293,In_428);
and U191 (N_191,In_238,In_462);
and U192 (N_192,In_24,In_469);
and U193 (N_193,In_127,In_277);
or U194 (N_194,In_450,In_159);
nand U195 (N_195,In_475,In_203);
or U196 (N_196,In_230,In_434);
or U197 (N_197,In_443,In_33);
and U198 (N_198,In_370,In_184);
nor U199 (N_199,In_188,In_163);
nor U200 (N_200,In_377,In_122);
or U201 (N_201,In_226,In_210);
nor U202 (N_202,In_413,In_190);
and U203 (N_203,In_224,In_399);
nand U204 (N_204,In_235,In_141);
nor U205 (N_205,In_426,In_44);
and U206 (N_206,In_489,In_205);
or U207 (N_207,In_375,In_481);
xor U208 (N_208,In_290,In_26);
or U209 (N_209,In_400,In_136);
nor U210 (N_210,In_284,In_403);
or U211 (N_211,In_217,In_92);
nor U212 (N_212,In_340,In_178);
nor U213 (N_213,In_34,In_274);
or U214 (N_214,In_225,In_339);
or U215 (N_215,In_249,In_196);
or U216 (N_216,In_255,In_254);
nor U217 (N_217,In_228,In_391);
or U218 (N_218,In_379,In_175);
and U219 (N_219,In_387,In_69);
or U220 (N_220,In_301,In_325);
and U221 (N_221,In_212,In_451);
nand U222 (N_222,In_65,In_192);
and U223 (N_223,In_466,In_38);
and U224 (N_224,In_435,In_459);
or U225 (N_225,In_318,In_270);
and U226 (N_226,In_262,In_10);
or U227 (N_227,In_120,In_328);
nand U228 (N_228,In_242,In_46);
or U229 (N_229,In_261,In_335);
nand U230 (N_230,In_79,In_342);
nand U231 (N_231,In_151,In_336);
nor U232 (N_232,In_408,In_465);
or U233 (N_233,In_13,In_398);
and U234 (N_234,In_3,In_186);
and U235 (N_235,In_347,In_119);
or U236 (N_236,In_54,In_302);
nor U237 (N_237,In_11,In_477);
nand U238 (N_238,In_43,In_166);
or U239 (N_239,In_213,In_438);
nand U240 (N_240,In_393,In_252);
and U241 (N_241,In_320,In_444);
or U242 (N_242,In_333,In_439);
nand U243 (N_243,In_71,In_338);
nand U244 (N_244,In_22,In_294);
nor U245 (N_245,In_19,In_201);
or U246 (N_246,In_77,In_289);
nand U247 (N_247,In_446,In_211);
or U248 (N_248,In_51,In_25);
or U249 (N_249,In_9,In_473);
or U250 (N_250,In_9,In_482);
or U251 (N_251,In_245,In_6);
or U252 (N_252,In_246,In_190);
and U253 (N_253,In_194,In_265);
nor U254 (N_254,In_300,In_311);
nor U255 (N_255,In_492,In_449);
and U256 (N_256,In_420,In_38);
or U257 (N_257,In_195,In_61);
nand U258 (N_258,In_415,In_233);
nand U259 (N_259,In_398,In_245);
nand U260 (N_260,In_341,In_478);
nand U261 (N_261,In_78,In_368);
and U262 (N_262,In_25,In_262);
nand U263 (N_263,In_203,In_129);
or U264 (N_264,In_323,In_128);
or U265 (N_265,In_105,In_416);
or U266 (N_266,In_241,In_144);
nor U267 (N_267,In_332,In_368);
nor U268 (N_268,In_370,In_376);
nor U269 (N_269,In_21,In_47);
or U270 (N_270,In_6,In_217);
or U271 (N_271,In_47,In_132);
nor U272 (N_272,In_312,In_130);
nand U273 (N_273,In_111,In_194);
nand U274 (N_274,In_476,In_454);
nand U275 (N_275,In_211,In_134);
and U276 (N_276,In_275,In_482);
or U277 (N_277,In_79,In_294);
nor U278 (N_278,In_432,In_368);
nand U279 (N_279,In_213,In_386);
nand U280 (N_280,In_81,In_223);
and U281 (N_281,In_37,In_466);
or U282 (N_282,In_42,In_208);
nand U283 (N_283,In_462,In_321);
and U284 (N_284,In_336,In_433);
and U285 (N_285,In_375,In_378);
nor U286 (N_286,In_242,In_40);
and U287 (N_287,In_302,In_264);
or U288 (N_288,In_262,In_271);
and U289 (N_289,In_69,In_498);
and U290 (N_290,In_133,In_379);
nand U291 (N_291,In_30,In_329);
nand U292 (N_292,In_482,In_358);
and U293 (N_293,In_255,In_166);
nor U294 (N_294,In_449,In_140);
and U295 (N_295,In_291,In_286);
nor U296 (N_296,In_156,In_492);
and U297 (N_297,In_105,In_179);
nand U298 (N_298,In_429,In_249);
or U299 (N_299,In_29,In_436);
nor U300 (N_300,In_355,In_475);
and U301 (N_301,In_199,In_99);
and U302 (N_302,In_466,In_342);
nand U303 (N_303,In_444,In_136);
or U304 (N_304,In_97,In_397);
and U305 (N_305,In_208,In_349);
nand U306 (N_306,In_232,In_127);
and U307 (N_307,In_133,In_335);
or U308 (N_308,In_242,In_269);
nor U309 (N_309,In_202,In_158);
and U310 (N_310,In_276,In_318);
or U311 (N_311,In_138,In_466);
nor U312 (N_312,In_218,In_214);
nand U313 (N_313,In_307,In_261);
nor U314 (N_314,In_128,In_98);
nand U315 (N_315,In_466,In_87);
or U316 (N_316,In_9,In_383);
nor U317 (N_317,In_364,In_307);
or U318 (N_318,In_99,In_313);
and U319 (N_319,In_76,In_134);
nor U320 (N_320,In_429,In_48);
or U321 (N_321,In_218,In_204);
xor U322 (N_322,In_223,In_249);
and U323 (N_323,In_181,In_50);
nor U324 (N_324,In_148,In_202);
or U325 (N_325,In_490,In_1);
nor U326 (N_326,In_5,In_243);
or U327 (N_327,In_464,In_446);
nor U328 (N_328,In_70,In_478);
xor U329 (N_329,In_316,In_490);
or U330 (N_330,In_300,In_423);
nor U331 (N_331,In_71,In_335);
nand U332 (N_332,In_20,In_324);
or U333 (N_333,In_265,In_51);
nand U334 (N_334,In_340,In_108);
and U335 (N_335,In_97,In_316);
nand U336 (N_336,In_371,In_324);
and U337 (N_337,In_203,In_277);
and U338 (N_338,In_155,In_461);
and U339 (N_339,In_215,In_463);
or U340 (N_340,In_195,In_122);
or U341 (N_341,In_71,In_173);
xor U342 (N_342,In_473,In_407);
xnor U343 (N_343,In_479,In_77);
or U344 (N_344,In_248,In_228);
nor U345 (N_345,In_352,In_19);
and U346 (N_346,In_348,In_328);
nor U347 (N_347,In_192,In_350);
or U348 (N_348,In_489,In_122);
or U349 (N_349,In_395,In_321);
and U350 (N_350,In_447,In_238);
nand U351 (N_351,In_212,In_121);
nand U352 (N_352,In_421,In_252);
and U353 (N_353,In_74,In_263);
nor U354 (N_354,In_92,In_213);
or U355 (N_355,In_385,In_213);
nor U356 (N_356,In_391,In_182);
or U357 (N_357,In_77,In_173);
or U358 (N_358,In_439,In_111);
nand U359 (N_359,In_268,In_270);
nand U360 (N_360,In_377,In_311);
or U361 (N_361,In_461,In_153);
nor U362 (N_362,In_293,In_407);
nor U363 (N_363,In_70,In_16);
nand U364 (N_364,In_309,In_19);
and U365 (N_365,In_490,In_4);
xor U366 (N_366,In_100,In_277);
nand U367 (N_367,In_306,In_246);
or U368 (N_368,In_274,In_465);
or U369 (N_369,In_381,In_69);
or U370 (N_370,In_111,In_271);
nand U371 (N_371,In_158,In_294);
nor U372 (N_372,In_363,In_43);
nor U373 (N_373,In_261,In_6);
or U374 (N_374,In_134,In_109);
nor U375 (N_375,In_140,In_470);
nand U376 (N_376,In_254,In_2);
or U377 (N_377,In_261,In_118);
nor U378 (N_378,In_331,In_213);
nand U379 (N_379,In_151,In_78);
or U380 (N_380,In_45,In_163);
or U381 (N_381,In_3,In_261);
nand U382 (N_382,In_195,In_477);
nor U383 (N_383,In_343,In_36);
nand U384 (N_384,In_499,In_433);
nor U385 (N_385,In_80,In_341);
nand U386 (N_386,In_309,In_48);
nor U387 (N_387,In_482,In_428);
or U388 (N_388,In_460,In_108);
and U389 (N_389,In_51,In_407);
nand U390 (N_390,In_269,In_32);
nor U391 (N_391,In_219,In_380);
and U392 (N_392,In_338,In_248);
nor U393 (N_393,In_181,In_118);
nand U394 (N_394,In_266,In_215);
and U395 (N_395,In_261,In_332);
nand U396 (N_396,In_461,In_364);
xnor U397 (N_397,In_352,In_41);
nand U398 (N_398,In_4,In_467);
nor U399 (N_399,In_180,In_44);
nor U400 (N_400,In_56,In_185);
xnor U401 (N_401,In_144,In_389);
and U402 (N_402,In_266,In_94);
xnor U403 (N_403,In_150,In_307);
nand U404 (N_404,In_389,In_65);
nand U405 (N_405,In_287,In_307);
or U406 (N_406,In_129,In_433);
nand U407 (N_407,In_34,In_60);
nand U408 (N_408,In_88,In_382);
nand U409 (N_409,In_447,In_305);
nand U410 (N_410,In_336,In_67);
and U411 (N_411,In_189,In_117);
xnor U412 (N_412,In_434,In_375);
nand U413 (N_413,In_425,In_51);
nor U414 (N_414,In_155,In_382);
nor U415 (N_415,In_222,In_130);
nor U416 (N_416,In_231,In_26);
nor U417 (N_417,In_447,In_19);
nand U418 (N_418,In_66,In_351);
nand U419 (N_419,In_126,In_307);
nor U420 (N_420,In_335,In_381);
and U421 (N_421,In_200,In_428);
or U422 (N_422,In_123,In_480);
nand U423 (N_423,In_234,In_11);
or U424 (N_424,In_235,In_315);
nor U425 (N_425,In_137,In_491);
nor U426 (N_426,In_396,In_182);
and U427 (N_427,In_296,In_419);
nor U428 (N_428,In_333,In_127);
nor U429 (N_429,In_314,In_329);
or U430 (N_430,In_139,In_57);
and U431 (N_431,In_31,In_266);
nor U432 (N_432,In_309,In_325);
or U433 (N_433,In_307,In_365);
nand U434 (N_434,In_404,In_203);
nor U435 (N_435,In_238,In_32);
nand U436 (N_436,In_249,In_125);
nor U437 (N_437,In_102,In_157);
nand U438 (N_438,In_29,In_90);
or U439 (N_439,In_379,In_183);
nand U440 (N_440,In_347,In_494);
and U441 (N_441,In_180,In_164);
xnor U442 (N_442,In_476,In_112);
nand U443 (N_443,In_145,In_439);
or U444 (N_444,In_282,In_360);
nand U445 (N_445,In_94,In_163);
xnor U446 (N_446,In_279,In_372);
and U447 (N_447,In_337,In_343);
nand U448 (N_448,In_221,In_218);
or U449 (N_449,In_97,In_214);
nand U450 (N_450,In_278,In_443);
nor U451 (N_451,In_406,In_83);
nand U452 (N_452,In_488,In_475);
nor U453 (N_453,In_405,In_187);
and U454 (N_454,In_426,In_247);
nor U455 (N_455,In_408,In_214);
and U456 (N_456,In_207,In_123);
nand U457 (N_457,In_299,In_66);
or U458 (N_458,In_456,In_464);
nor U459 (N_459,In_452,In_364);
nand U460 (N_460,In_50,In_373);
nor U461 (N_461,In_235,In_95);
nand U462 (N_462,In_397,In_5);
or U463 (N_463,In_107,In_384);
or U464 (N_464,In_120,In_304);
nor U465 (N_465,In_28,In_484);
nor U466 (N_466,In_349,In_312);
or U467 (N_467,In_421,In_491);
nor U468 (N_468,In_185,In_122);
and U469 (N_469,In_493,In_443);
or U470 (N_470,In_207,In_424);
nor U471 (N_471,In_394,In_319);
nor U472 (N_472,In_248,In_414);
nor U473 (N_473,In_416,In_452);
or U474 (N_474,In_489,In_31);
nor U475 (N_475,In_137,In_280);
nor U476 (N_476,In_360,In_253);
or U477 (N_477,In_291,In_273);
or U478 (N_478,In_281,In_104);
or U479 (N_479,In_153,In_111);
nor U480 (N_480,In_390,In_160);
nand U481 (N_481,In_430,In_334);
or U482 (N_482,In_296,In_1);
nand U483 (N_483,In_189,In_351);
or U484 (N_484,In_167,In_251);
nor U485 (N_485,In_187,In_116);
nor U486 (N_486,In_185,In_421);
nor U487 (N_487,In_421,In_162);
and U488 (N_488,In_465,In_463);
nor U489 (N_489,In_319,In_356);
nor U490 (N_490,In_362,In_29);
and U491 (N_491,In_367,In_127);
nor U492 (N_492,In_332,In_413);
and U493 (N_493,In_61,In_422);
or U494 (N_494,In_107,In_171);
nand U495 (N_495,In_471,In_188);
or U496 (N_496,In_315,In_27);
nand U497 (N_497,In_181,In_350);
or U498 (N_498,In_124,In_162);
nor U499 (N_499,In_308,In_367);
nand U500 (N_500,N_455,N_454);
nand U501 (N_501,N_113,N_42);
and U502 (N_502,N_157,N_218);
or U503 (N_503,N_291,N_204);
or U504 (N_504,N_417,N_104);
and U505 (N_505,N_100,N_213);
nor U506 (N_506,N_362,N_98);
nand U507 (N_507,N_324,N_363);
nand U508 (N_508,N_331,N_378);
nor U509 (N_509,N_115,N_51);
or U510 (N_510,N_240,N_97);
nor U511 (N_511,N_321,N_158);
nand U512 (N_512,N_253,N_451);
nor U513 (N_513,N_88,N_339);
nor U514 (N_514,N_193,N_462);
nand U515 (N_515,N_265,N_85);
and U516 (N_516,N_242,N_478);
and U517 (N_517,N_261,N_459);
or U518 (N_518,N_60,N_465);
nor U519 (N_519,N_142,N_195);
nand U520 (N_520,N_189,N_241);
xnor U521 (N_521,N_101,N_427);
and U522 (N_522,N_479,N_401);
nand U523 (N_523,N_174,N_364);
and U524 (N_524,N_44,N_263);
nand U525 (N_525,N_367,N_235);
nand U526 (N_526,N_29,N_143);
nor U527 (N_527,N_288,N_50);
nand U528 (N_528,N_395,N_33);
nand U529 (N_529,N_422,N_39);
or U530 (N_530,N_128,N_262);
nor U531 (N_531,N_238,N_110);
or U532 (N_532,N_251,N_63);
nor U533 (N_533,N_248,N_295);
or U534 (N_534,N_147,N_394);
or U535 (N_535,N_46,N_471);
or U536 (N_536,N_130,N_3);
nor U537 (N_537,N_149,N_173);
nand U538 (N_538,N_168,N_16);
or U539 (N_539,N_172,N_388);
nor U540 (N_540,N_268,N_30);
or U541 (N_541,N_296,N_171);
nand U542 (N_542,N_102,N_223);
nand U543 (N_543,N_65,N_317);
nor U544 (N_544,N_418,N_293);
nand U545 (N_545,N_322,N_413);
nor U546 (N_546,N_20,N_109);
or U547 (N_547,N_164,N_220);
and U548 (N_548,N_430,N_267);
nor U549 (N_549,N_284,N_8);
xnor U550 (N_550,N_239,N_398);
or U551 (N_551,N_396,N_419);
or U552 (N_552,N_209,N_308);
and U553 (N_553,N_494,N_194);
and U554 (N_554,N_304,N_286);
xnor U555 (N_555,N_136,N_337);
or U556 (N_556,N_386,N_498);
or U557 (N_557,N_292,N_469);
nand U558 (N_558,N_230,N_86);
or U559 (N_559,N_305,N_408);
and U560 (N_560,N_146,N_71);
or U561 (N_561,N_370,N_464);
xor U562 (N_562,N_461,N_476);
nor U563 (N_563,N_491,N_256);
nand U564 (N_564,N_225,N_426);
and U565 (N_565,N_151,N_217);
or U566 (N_566,N_332,N_45);
nor U567 (N_567,N_379,N_312);
nand U568 (N_568,N_373,N_446);
or U569 (N_569,N_310,N_325);
nand U570 (N_570,N_120,N_392);
and U571 (N_571,N_202,N_87);
nand U572 (N_572,N_107,N_210);
or U573 (N_573,N_384,N_52);
and U574 (N_574,N_22,N_423);
or U575 (N_575,N_196,N_328);
and U576 (N_576,N_458,N_41);
nand U577 (N_577,N_257,N_409);
nand U578 (N_578,N_404,N_393);
nor U579 (N_579,N_273,N_237);
nor U580 (N_580,N_497,N_117);
and U581 (N_581,N_477,N_59);
and U582 (N_582,N_390,N_91);
nor U583 (N_583,N_485,N_191);
nand U584 (N_584,N_244,N_349);
and U585 (N_585,N_445,N_57);
nand U586 (N_586,N_323,N_319);
or U587 (N_587,N_69,N_429);
and U588 (N_588,N_435,N_152);
nor U589 (N_589,N_473,N_212);
nor U590 (N_590,N_340,N_432);
or U591 (N_591,N_133,N_376);
nand U592 (N_592,N_206,N_54);
nand U593 (N_593,N_68,N_275);
or U594 (N_594,N_391,N_226);
or U595 (N_595,N_350,N_31);
and U596 (N_596,N_166,N_233);
nor U597 (N_597,N_399,N_129);
or U598 (N_598,N_397,N_372);
nand U599 (N_599,N_222,N_474);
or U600 (N_600,N_303,N_90);
or U601 (N_601,N_170,N_12);
or U602 (N_602,N_387,N_5);
nor U603 (N_603,N_407,N_205);
and U604 (N_604,N_442,N_94);
and U605 (N_605,N_326,N_276);
and U606 (N_606,N_377,N_283);
or U607 (N_607,N_499,N_277);
or U608 (N_608,N_258,N_438);
nor U609 (N_609,N_285,N_420);
xor U610 (N_610,N_47,N_389);
and U611 (N_611,N_132,N_301);
nand U612 (N_612,N_99,N_165);
and U613 (N_613,N_467,N_338);
nand U614 (N_614,N_247,N_259);
and U615 (N_615,N_334,N_229);
and U616 (N_616,N_139,N_234);
or U617 (N_617,N_400,N_306);
nor U618 (N_618,N_64,N_314);
or U619 (N_619,N_297,N_403);
nand U620 (N_620,N_181,N_19);
nor U621 (N_621,N_184,N_448);
and U622 (N_622,N_320,N_289);
nand U623 (N_623,N_232,N_468);
nand U624 (N_624,N_23,N_187);
nor U625 (N_625,N_188,N_280);
nor U626 (N_626,N_493,N_126);
and U627 (N_627,N_72,N_495);
or U628 (N_628,N_255,N_178);
and U629 (N_629,N_431,N_375);
and U630 (N_630,N_342,N_0);
nand U631 (N_631,N_211,N_347);
and U632 (N_632,N_36,N_439);
and U633 (N_633,N_300,N_140);
or U634 (N_634,N_333,N_406);
nand U635 (N_635,N_412,N_70);
nand U636 (N_636,N_77,N_249);
xnor U637 (N_637,N_313,N_74);
and U638 (N_638,N_79,N_48);
nor U639 (N_639,N_318,N_252);
or U640 (N_640,N_260,N_484);
or U641 (N_641,N_346,N_203);
and U642 (N_642,N_169,N_298);
and U643 (N_643,N_492,N_245);
and U644 (N_644,N_472,N_282);
nand U645 (N_645,N_161,N_290);
nor U646 (N_646,N_18,N_34);
and U647 (N_647,N_215,N_108);
nor U648 (N_648,N_82,N_433);
and U649 (N_649,N_138,N_201);
or U650 (N_650,N_264,N_4);
and U651 (N_651,N_270,N_311);
or U652 (N_652,N_119,N_227);
nor U653 (N_653,N_14,N_357);
xnor U654 (N_654,N_371,N_32);
or U655 (N_655,N_355,N_344);
nor U656 (N_656,N_2,N_354);
nor U657 (N_657,N_353,N_482);
nand U658 (N_658,N_141,N_121);
nand U659 (N_659,N_341,N_112);
nand U660 (N_660,N_453,N_425);
nor U661 (N_661,N_271,N_95);
or U662 (N_662,N_302,N_281);
xor U663 (N_663,N_254,N_137);
and U664 (N_664,N_374,N_444);
nor U665 (N_665,N_266,N_190);
nand U666 (N_666,N_335,N_221);
nor U667 (N_667,N_352,N_192);
nand U668 (N_668,N_414,N_294);
nand U669 (N_669,N_182,N_150);
nand U670 (N_670,N_410,N_330);
nand U671 (N_671,N_463,N_460);
nor U672 (N_672,N_228,N_197);
nor U673 (N_673,N_160,N_307);
and U674 (N_674,N_27,N_424);
nand U675 (N_675,N_489,N_443);
or U676 (N_676,N_58,N_368);
nor U677 (N_677,N_274,N_483);
and U678 (N_678,N_486,N_84);
and U679 (N_679,N_24,N_200);
nand U680 (N_680,N_421,N_162);
nand U681 (N_681,N_148,N_358);
nand U682 (N_682,N_83,N_207);
or U683 (N_683,N_15,N_124);
nand U684 (N_684,N_76,N_279);
or U685 (N_685,N_134,N_125);
nand U686 (N_686,N_66,N_415);
and U687 (N_687,N_488,N_440);
and U688 (N_688,N_316,N_7);
and U689 (N_689,N_456,N_327);
or U690 (N_690,N_55,N_470);
and U691 (N_691,N_49,N_450);
nand U692 (N_692,N_299,N_176);
and U693 (N_693,N_10,N_447);
or U694 (N_694,N_231,N_236);
nor U695 (N_695,N_361,N_1);
or U696 (N_696,N_40,N_216);
nor U697 (N_697,N_214,N_405);
and U698 (N_698,N_382,N_26);
and U699 (N_699,N_67,N_103);
or U700 (N_700,N_180,N_437);
nor U701 (N_701,N_287,N_345);
or U702 (N_702,N_198,N_336);
and U703 (N_703,N_457,N_123);
nor U704 (N_704,N_28,N_428);
nor U705 (N_705,N_9,N_81);
nand U706 (N_706,N_480,N_369);
nor U707 (N_707,N_177,N_145);
and U708 (N_708,N_53,N_154);
or U709 (N_709,N_411,N_61);
and U710 (N_710,N_466,N_380);
nand U711 (N_711,N_436,N_329);
nor U712 (N_712,N_208,N_402);
nand U713 (N_713,N_315,N_360);
and U714 (N_714,N_343,N_35);
nand U715 (N_715,N_144,N_111);
or U716 (N_716,N_106,N_366);
nand U717 (N_717,N_127,N_269);
or U718 (N_718,N_434,N_348);
nor U719 (N_719,N_131,N_481);
nor U720 (N_720,N_175,N_385);
nor U721 (N_721,N_11,N_73);
or U722 (N_722,N_416,N_356);
nor U723 (N_723,N_75,N_62);
nor U724 (N_724,N_118,N_383);
nor U725 (N_725,N_25,N_359);
nand U726 (N_726,N_116,N_17);
nand U727 (N_727,N_105,N_93);
or U728 (N_728,N_243,N_96);
nand U729 (N_729,N_43,N_122);
nor U730 (N_730,N_89,N_309);
nand U731 (N_731,N_351,N_21);
or U732 (N_732,N_199,N_441);
or U733 (N_733,N_159,N_490);
and U734 (N_734,N_92,N_475);
nor U735 (N_735,N_224,N_13);
and U736 (N_736,N_38,N_155);
and U737 (N_737,N_135,N_487);
nor U738 (N_738,N_167,N_78);
and U739 (N_739,N_80,N_114);
nand U740 (N_740,N_153,N_56);
or U741 (N_741,N_219,N_278);
nand U742 (N_742,N_452,N_6);
nand U743 (N_743,N_250,N_183);
and U744 (N_744,N_272,N_156);
or U745 (N_745,N_163,N_381);
nor U746 (N_746,N_246,N_496);
nand U747 (N_747,N_37,N_185);
or U748 (N_748,N_179,N_186);
xnor U749 (N_749,N_365,N_449);
nor U750 (N_750,N_164,N_125);
nor U751 (N_751,N_295,N_468);
nand U752 (N_752,N_313,N_338);
nand U753 (N_753,N_2,N_151);
or U754 (N_754,N_49,N_177);
and U755 (N_755,N_127,N_347);
nor U756 (N_756,N_39,N_289);
and U757 (N_757,N_349,N_310);
nor U758 (N_758,N_87,N_111);
or U759 (N_759,N_64,N_56);
and U760 (N_760,N_319,N_483);
and U761 (N_761,N_335,N_52);
nand U762 (N_762,N_40,N_203);
or U763 (N_763,N_342,N_396);
or U764 (N_764,N_399,N_82);
and U765 (N_765,N_402,N_119);
or U766 (N_766,N_31,N_299);
nand U767 (N_767,N_156,N_60);
or U768 (N_768,N_491,N_233);
nand U769 (N_769,N_56,N_271);
or U770 (N_770,N_57,N_374);
or U771 (N_771,N_196,N_294);
and U772 (N_772,N_54,N_412);
or U773 (N_773,N_159,N_96);
or U774 (N_774,N_110,N_140);
xnor U775 (N_775,N_416,N_190);
nand U776 (N_776,N_438,N_50);
or U777 (N_777,N_311,N_72);
or U778 (N_778,N_103,N_289);
and U779 (N_779,N_73,N_389);
nor U780 (N_780,N_231,N_163);
nor U781 (N_781,N_377,N_96);
or U782 (N_782,N_28,N_401);
nor U783 (N_783,N_156,N_430);
or U784 (N_784,N_148,N_130);
and U785 (N_785,N_111,N_66);
and U786 (N_786,N_280,N_413);
nand U787 (N_787,N_417,N_212);
nor U788 (N_788,N_155,N_365);
nor U789 (N_789,N_406,N_86);
nand U790 (N_790,N_52,N_439);
nor U791 (N_791,N_397,N_204);
or U792 (N_792,N_348,N_462);
nand U793 (N_793,N_308,N_22);
nand U794 (N_794,N_124,N_39);
nor U795 (N_795,N_385,N_431);
or U796 (N_796,N_171,N_226);
or U797 (N_797,N_404,N_262);
and U798 (N_798,N_319,N_286);
nand U799 (N_799,N_224,N_445);
nand U800 (N_800,N_361,N_157);
or U801 (N_801,N_180,N_70);
nor U802 (N_802,N_306,N_186);
and U803 (N_803,N_313,N_104);
or U804 (N_804,N_2,N_395);
and U805 (N_805,N_11,N_350);
and U806 (N_806,N_463,N_219);
nor U807 (N_807,N_372,N_211);
and U808 (N_808,N_245,N_207);
nor U809 (N_809,N_415,N_481);
nand U810 (N_810,N_476,N_90);
nand U811 (N_811,N_302,N_253);
or U812 (N_812,N_386,N_254);
or U813 (N_813,N_215,N_472);
nand U814 (N_814,N_160,N_243);
and U815 (N_815,N_81,N_31);
and U816 (N_816,N_1,N_106);
nand U817 (N_817,N_52,N_117);
or U818 (N_818,N_294,N_340);
nand U819 (N_819,N_32,N_138);
xor U820 (N_820,N_346,N_132);
nor U821 (N_821,N_100,N_179);
nand U822 (N_822,N_146,N_130);
nor U823 (N_823,N_94,N_57);
nor U824 (N_824,N_142,N_91);
or U825 (N_825,N_219,N_350);
nand U826 (N_826,N_22,N_269);
or U827 (N_827,N_146,N_143);
nand U828 (N_828,N_114,N_64);
and U829 (N_829,N_14,N_25);
nand U830 (N_830,N_310,N_188);
or U831 (N_831,N_188,N_388);
nor U832 (N_832,N_170,N_454);
nand U833 (N_833,N_134,N_225);
xor U834 (N_834,N_125,N_388);
and U835 (N_835,N_135,N_317);
and U836 (N_836,N_373,N_6);
and U837 (N_837,N_307,N_181);
or U838 (N_838,N_127,N_139);
nor U839 (N_839,N_251,N_54);
and U840 (N_840,N_454,N_242);
and U841 (N_841,N_299,N_168);
or U842 (N_842,N_372,N_71);
or U843 (N_843,N_185,N_475);
nand U844 (N_844,N_116,N_68);
xor U845 (N_845,N_365,N_212);
nor U846 (N_846,N_153,N_286);
and U847 (N_847,N_368,N_367);
or U848 (N_848,N_238,N_243);
nand U849 (N_849,N_455,N_138);
or U850 (N_850,N_404,N_130);
nor U851 (N_851,N_248,N_457);
nand U852 (N_852,N_345,N_79);
and U853 (N_853,N_360,N_329);
or U854 (N_854,N_361,N_267);
nor U855 (N_855,N_195,N_220);
nand U856 (N_856,N_194,N_358);
nor U857 (N_857,N_425,N_346);
nor U858 (N_858,N_182,N_175);
nor U859 (N_859,N_54,N_451);
nand U860 (N_860,N_97,N_428);
or U861 (N_861,N_157,N_155);
nand U862 (N_862,N_147,N_75);
nor U863 (N_863,N_96,N_363);
and U864 (N_864,N_161,N_448);
nand U865 (N_865,N_257,N_9);
and U866 (N_866,N_436,N_407);
and U867 (N_867,N_84,N_465);
nor U868 (N_868,N_249,N_28);
or U869 (N_869,N_169,N_99);
or U870 (N_870,N_201,N_20);
or U871 (N_871,N_127,N_11);
nand U872 (N_872,N_484,N_393);
and U873 (N_873,N_427,N_121);
nor U874 (N_874,N_209,N_197);
and U875 (N_875,N_272,N_127);
nand U876 (N_876,N_465,N_280);
nand U877 (N_877,N_333,N_194);
or U878 (N_878,N_104,N_71);
nand U879 (N_879,N_299,N_287);
or U880 (N_880,N_477,N_406);
or U881 (N_881,N_169,N_146);
nor U882 (N_882,N_202,N_30);
or U883 (N_883,N_171,N_283);
nand U884 (N_884,N_420,N_67);
and U885 (N_885,N_168,N_17);
and U886 (N_886,N_83,N_251);
or U887 (N_887,N_435,N_207);
nor U888 (N_888,N_278,N_153);
or U889 (N_889,N_18,N_442);
and U890 (N_890,N_172,N_219);
or U891 (N_891,N_221,N_391);
or U892 (N_892,N_459,N_301);
and U893 (N_893,N_361,N_136);
and U894 (N_894,N_184,N_462);
nand U895 (N_895,N_429,N_453);
nand U896 (N_896,N_186,N_9);
or U897 (N_897,N_40,N_339);
and U898 (N_898,N_376,N_79);
nor U899 (N_899,N_487,N_353);
nor U900 (N_900,N_422,N_243);
nand U901 (N_901,N_424,N_34);
nand U902 (N_902,N_417,N_330);
or U903 (N_903,N_339,N_247);
or U904 (N_904,N_161,N_106);
or U905 (N_905,N_161,N_285);
nor U906 (N_906,N_195,N_210);
nand U907 (N_907,N_273,N_337);
or U908 (N_908,N_163,N_115);
and U909 (N_909,N_411,N_106);
nor U910 (N_910,N_451,N_218);
and U911 (N_911,N_419,N_447);
and U912 (N_912,N_491,N_35);
or U913 (N_913,N_397,N_490);
and U914 (N_914,N_225,N_84);
nand U915 (N_915,N_363,N_482);
nand U916 (N_916,N_199,N_180);
or U917 (N_917,N_220,N_308);
or U918 (N_918,N_414,N_451);
or U919 (N_919,N_150,N_336);
and U920 (N_920,N_372,N_357);
and U921 (N_921,N_323,N_316);
and U922 (N_922,N_221,N_134);
and U923 (N_923,N_297,N_183);
xor U924 (N_924,N_196,N_79);
and U925 (N_925,N_67,N_89);
and U926 (N_926,N_66,N_119);
or U927 (N_927,N_313,N_435);
and U928 (N_928,N_236,N_46);
and U929 (N_929,N_318,N_169);
nor U930 (N_930,N_73,N_481);
nand U931 (N_931,N_260,N_467);
nand U932 (N_932,N_337,N_144);
nand U933 (N_933,N_438,N_255);
nand U934 (N_934,N_458,N_412);
nor U935 (N_935,N_142,N_234);
or U936 (N_936,N_291,N_95);
nor U937 (N_937,N_393,N_280);
xnor U938 (N_938,N_214,N_83);
nand U939 (N_939,N_325,N_253);
nor U940 (N_940,N_63,N_23);
and U941 (N_941,N_39,N_397);
nand U942 (N_942,N_311,N_122);
nor U943 (N_943,N_165,N_275);
nor U944 (N_944,N_367,N_392);
xor U945 (N_945,N_104,N_227);
or U946 (N_946,N_165,N_260);
or U947 (N_947,N_200,N_406);
and U948 (N_948,N_235,N_478);
nand U949 (N_949,N_168,N_356);
and U950 (N_950,N_196,N_482);
nand U951 (N_951,N_394,N_40);
or U952 (N_952,N_128,N_442);
and U953 (N_953,N_56,N_30);
nor U954 (N_954,N_56,N_196);
nor U955 (N_955,N_396,N_349);
or U956 (N_956,N_393,N_227);
xor U957 (N_957,N_454,N_10);
or U958 (N_958,N_265,N_240);
nor U959 (N_959,N_182,N_394);
or U960 (N_960,N_130,N_250);
nor U961 (N_961,N_339,N_153);
nand U962 (N_962,N_75,N_144);
and U963 (N_963,N_459,N_485);
or U964 (N_964,N_16,N_11);
or U965 (N_965,N_18,N_294);
or U966 (N_966,N_303,N_296);
or U967 (N_967,N_483,N_222);
nor U968 (N_968,N_390,N_425);
nor U969 (N_969,N_368,N_44);
or U970 (N_970,N_185,N_441);
or U971 (N_971,N_444,N_292);
and U972 (N_972,N_116,N_36);
and U973 (N_973,N_434,N_460);
nand U974 (N_974,N_183,N_458);
xnor U975 (N_975,N_176,N_461);
or U976 (N_976,N_269,N_232);
nand U977 (N_977,N_455,N_271);
and U978 (N_978,N_272,N_286);
nor U979 (N_979,N_3,N_159);
nor U980 (N_980,N_226,N_290);
nor U981 (N_981,N_384,N_10);
and U982 (N_982,N_498,N_111);
nand U983 (N_983,N_391,N_88);
or U984 (N_984,N_360,N_70);
or U985 (N_985,N_236,N_98);
or U986 (N_986,N_447,N_183);
nand U987 (N_987,N_170,N_234);
nand U988 (N_988,N_117,N_44);
nor U989 (N_989,N_297,N_241);
nand U990 (N_990,N_159,N_218);
nor U991 (N_991,N_83,N_65);
nand U992 (N_992,N_334,N_238);
and U993 (N_993,N_261,N_496);
nor U994 (N_994,N_74,N_163);
nand U995 (N_995,N_9,N_254);
nor U996 (N_996,N_98,N_494);
or U997 (N_997,N_335,N_424);
and U998 (N_998,N_182,N_299);
nor U999 (N_999,N_98,N_130);
or U1000 (N_1000,N_984,N_908);
nand U1001 (N_1001,N_577,N_927);
xor U1002 (N_1002,N_748,N_862);
or U1003 (N_1003,N_688,N_824);
nor U1004 (N_1004,N_872,N_949);
nor U1005 (N_1005,N_605,N_656);
or U1006 (N_1006,N_952,N_550);
nor U1007 (N_1007,N_533,N_669);
or U1008 (N_1008,N_621,N_658);
and U1009 (N_1009,N_822,N_902);
or U1010 (N_1010,N_813,N_585);
xor U1011 (N_1011,N_981,N_840);
nor U1012 (N_1012,N_555,N_523);
and U1013 (N_1013,N_630,N_869);
and U1014 (N_1014,N_809,N_799);
and U1015 (N_1015,N_945,N_801);
nand U1016 (N_1016,N_645,N_744);
nand U1017 (N_1017,N_738,N_566);
and U1018 (N_1018,N_768,N_519);
nor U1019 (N_1019,N_922,N_674);
nor U1020 (N_1020,N_563,N_864);
or U1021 (N_1021,N_561,N_570);
or U1022 (N_1022,N_584,N_646);
and U1023 (N_1023,N_719,N_900);
and U1024 (N_1024,N_884,N_733);
and U1025 (N_1025,N_766,N_863);
or U1026 (N_1026,N_851,N_677);
nor U1027 (N_1027,N_591,N_534);
nor U1028 (N_1028,N_761,N_708);
nand U1029 (N_1029,N_704,N_685);
nor U1030 (N_1030,N_640,N_832);
nand U1031 (N_1031,N_507,N_680);
or U1032 (N_1032,N_700,N_713);
nand U1033 (N_1033,N_589,N_804);
or U1034 (N_1034,N_643,N_966);
nand U1035 (N_1035,N_785,N_702);
nor U1036 (N_1036,N_793,N_556);
or U1037 (N_1037,N_746,N_635);
or U1038 (N_1038,N_641,N_790);
nor U1039 (N_1039,N_559,N_987);
nand U1040 (N_1040,N_762,N_920);
nor U1041 (N_1041,N_609,N_991);
xor U1042 (N_1042,N_564,N_539);
xor U1043 (N_1043,N_831,N_756);
nand U1044 (N_1044,N_871,N_974);
nand U1045 (N_1045,N_812,N_825);
and U1046 (N_1046,N_632,N_509);
or U1047 (N_1047,N_948,N_896);
and U1048 (N_1048,N_633,N_932);
and U1049 (N_1049,N_714,N_676);
and U1050 (N_1050,N_930,N_800);
and U1051 (N_1051,N_619,N_829);
nand U1052 (N_1052,N_520,N_530);
or U1053 (N_1053,N_725,N_972);
nand U1054 (N_1054,N_998,N_703);
or U1055 (N_1055,N_729,N_868);
or U1056 (N_1056,N_717,N_690);
nand U1057 (N_1057,N_882,N_707);
and U1058 (N_1058,N_846,N_529);
and U1059 (N_1059,N_568,N_918);
nor U1060 (N_1060,N_992,N_888);
nand U1061 (N_1061,N_931,N_944);
or U1062 (N_1062,N_755,N_541);
or U1063 (N_1063,N_837,N_592);
and U1064 (N_1064,N_671,N_759);
nor U1065 (N_1065,N_834,N_826);
nand U1066 (N_1066,N_560,N_508);
nor U1067 (N_1067,N_805,N_664);
nor U1068 (N_1068,N_919,N_603);
nand U1069 (N_1069,N_692,N_976);
and U1070 (N_1070,N_522,N_739);
nand U1071 (N_1071,N_540,N_731);
nor U1072 (N_1072,N_623,N_587);
or U1073 (N_1073,N_933,N_955);
nor U1074 (N_1074,N_775,N_629);
and U1075 (N_1075,N_528,N_924);
and U1076 (N_1076,N_960,N_773);
nor U1077 (N_1077,N_861,N_878);
nand U1078 (N_1078,N_810,N_689);
nor U1079 (N_1079,N_890,N_894);
xor U1080 (N_1080,N_770,N_604);
nand U1081 (N_1081,N_705,N_965);
or U1082 (N_1082,N_710,N_916);
and U1083 (N_1083,N_784,N_820);
or U1084 (N_1084,N_501,N_934);
nor U1085 (N_1085,N_600,N_659);
and U1086 (N_1086,N_737,N_835);
nand U1087 (N_1087,N_726,N_736);
nand U1088 (N_1088,N_866,N_682);
nor U1089 (N_1089,N_946,N_767);
nor U1090 (N_1090,N_648,N_780);
or U1091 (N_1091,N_982,N_973);
or U1092 (N_1092,N_986,N_597);
nand U1093 (N_1093,N_819,N_652);
nor U1094 (N_1094,N_712,N_830);
nor U1095 (N_1095,N_625,N_915);
or U1096 (N_1096,N_607,N_673);
and U1097 (N_1097,N_750,N_734);
nand U1098 (N_1098,N_937,N_879);
nor U1099 (N_1099,N_569,N_838);
nor U1100 (N_1100,N_683,N_647);
and U1101 (N_1101,N_985,N_961);
or U1102 (N_1102,N_581,N_663);
and U1103 (N_1103,N_582,N_634);
and U1104 (N_1104,N_665,N_580);
and U1105 (N_1105,N_874,N_613);
and U1106 (N_1106,N_857,N_802);
or U1107 (N_1107,N_660,N_836);
or U1108 (N_1108,N_709,N_886);
nor U1109 (N_1109,N_936,N_903);
and U1110 (N_1110,N_892,N_791);
nand U1111 (N_1111,N_887,N_798);
nand U1112 (N_1112,N_551,N_667);
and U1113 (N_1113,N_867,N_828);
nand U1114 (N_1114,N_576,N_670);
nor U1115 (N_1115,N_516,N_899);
nor U1116 (N_1116,N_891,N_925);
and U1117 (N_1117,N_905,N_769);
nand U1118 (N_1118,N_538,N_814);
nand U1119 (N_1119,N_881,N_661);
and U1120 (N_1120,N_722,N_675);
nor U1121 (N_1121,N_720,N_521);
and U1122 (N_1122,N_907,N_854);
nor U1123 (N_1123,N_792,N_962);
or U1124 (N_1124,N_964,N_914);
nand U1125 (N_1125,N_618,N_574);
nor U1126 (N_1126,N_579,N_525);
nor U1127 (N_1127,N_953,N_990);
or U1128 (N_1128,N_994,N_686);
nand U1129 (N_1129,N_557,N_572);
nor U1130 (N_1130,N_777,N_935);
nand U1131 (N_1131,N_856,N_701);
nand U1132 (N_1132,N_653,N_628);
nand U1133 (N_1133,N_757,N_947);
nor U1134 (N_1134,N_723,N_993);
nand U1135 (N_1135,N_626,N_865);
nand U1136 (N_1136,N_906,N_742);
and U1137 (N_1137,N_558,N_627);
and U1138 (N_1138,N_778,N_841);
or U1139 (N_1139,N_687,N_606);
nand U1140 (N_1140,N_763,N_910);
and U1141 (N_1141,N_850,N_803);
and U1142 (N_1142,N_938,N_532);
nand U1143 (N_1143,N_752,N_913);
nand U1144 (N_1144,N_977,N_855);
or U1145 (N_1145,N_601,N_642);
nand U1146 (N_1146,N_622,N_928);
or U1147 (N_1147,N_715,N_728);
or U1148 (N_1148,N_735,N_997);
or U1149 (N_1149,N_873,N_771);
nor U1150 (N_1150,N_758,N_917);
or U1151 (N_1151,N_624,N_536);
or U1152 (N_1152,N_511,N_885);
or U1153 (N_1153,N_537,N_975);
and U1154 (N_1154,N_679,N_573);
or U1155 (N_1155,N_544,N_612);
nand U1156 (N_1156,N_843,N_706);
nor U1157 (N_1157,N_795,N_833);
and U1158 (N_1158,N_594,N_893);
and U1159 (N_1159,N_583,N_847);
or U1160 (N_1160,N_901,N_988);
xnor U1161 (N_1161,N_514,N_554);
nor U1162 (N_1162,N_839,N_747);
and U1163 (N_1163,N_774,N_786);
and U1164 (N_1164,N_852,N_724);
and U1165 (N_1165,N_921,N_808);
nor U1166 (N_1166,N_950,N_615);
nor U1167 (N_1167,N_904,N_858);
or U1168 (N_1168,N_553,N_788);
and U1169 (N_1169,N_787,N_698);
nand U1170 (N_1170,N_848,N_970);
xor U1171 (N_1171,N_958,N_505);
or U1172 (N_1172,N_876,N_883);
nand U1173 (N_1173,N_989,N_517);
nand U1174 (N_1174,N_562,N_548);
or U1175 (N_1175,N_691,N_753);
nand U1176 (N_1176,N_794,N_806);
or U1177 (N_1177,N_796,N_956);
nand U1178 (N_1178,N_877,N_870);
nand U1179 (N_1179,N_513,N_760);
and U1180 (N_1180,N_510,N_711);
or U1181 (N_1181,N_593,N_929);
nand U1182 (N_1182,N_942,N_897);
nand U1183 (N_1183,N_504,N_655);
nor U1184 (N_1184,N_602,N_821);
or U1185 (N_1185,N_666,N_547);
nand U1186 (N_1186,N_754,N_695);
and U1187 (N_1187,N_542,N_911);
or U1188 (N_1188,N_764,N_979);
nand U1189 (N_1189,N_500,N_781);
or U1190 (N_1190,N_811,N_880);
or U1191 (N_1191,N_730,N_608);
and U1192 (N_1192,N_684,N_662);
or U1193 (N_1193,N_818,N_815);
or U1194 (N_1194,N_860,N_595);
and U1195 (N_1195,N_527,N_611);
or U1196 (N_1196,N_515,N_567);
nand U1197 (N_1197,N_827,N_693);
nand U1198 (N_1198,N_649,N_512);
or U1199 (N_1199,N_939,N_853);
and U1200 (N_1200,N_817,N_816);
nor U1201 (N_1201,N_549,N_616);
nor U1202 (N_1202,N_610,N_971);
or U1203 (N_1203,N_503,N_526);
and U1204 (N_1204,N_650,N_782);
or U1205 (N_1205,N_578,N_639);
and U1206 (N_1206,N_740,N_644);
nor U1207 (N_1207,N_776,N_783);
nor U1208 (N_1208,N_963,N_849);
and U1209 (N_1209,N_518,N_954);
nor U1210 (N_1210,N_651,N_875);
nand U1211 (N_1211,N_749,N_524);
or U1212 (N_1212,N_957,N_909);
and U1213 (N_1213,N_959,N_845);
nand U1214 (N_1214,N_940,N_599);
nand U1215 (N_1215,N_575,N_637);
nand U1216 (N_1216,N_678,N_978);
nand U1217 (N_1217,N_620,N_797);
and U1218 (N_1218,N_745,N_614);
and U1219 (N_1219,N_943,N_842);
nor U1220 (N_1220,N_535,N_545);
nand U1221 (N_1221,N_694,N_941);
and U1222 (N_1222,N_654,N_969);
nor U1223 (N_1223,N_983,N_823);
nor U1224 (N_1224,N_772,N_506);
nor U1225 (N_1225,N_765,N_951);
and U1226 (N_1226,N_968,N_727);
nor U1227 (N_1227,N_681,N_743);
and U1228 (N_1228,N_502,N_980);
nand U1229 (N_1229,N_546,N_617);
nor U1230 (N_1230,N_586,N_889);
and U1231 (N_1231,N_699,N_716);
nand U1232 (N_1232,N_844,N_631);
and U1233 (N_1233,N_588,N_590);
nor U1234 (N_1234,N_696,N_697);
or U1235 (N_1235,N_751,N_638);
nor U1236 (N_1236,N_779,N_895);
and U1237 (N_1237,N_732,N_668);
xnor U1238 (N_1238,N_926,N_741);
or U1239 (N_1239,N_657,N_999);
or U1240 (N_1240,N_672,N_598);
or U1241 (N_1241,N_912,N_543);
or U1242 (N_1242,N_571,N_565);
xor U1243 (N_1243,N_531,N_923);
xnor U1244 (N_1244,N_596,N_967);
nor U1245 (N_1245,N_552,N_636);
nor U1246 (N_1246,N_859,N_721);
nor U1247 (N_1247,N_718,N_995);
or U1248 (N_1248,N_996,N_807);
nand U1249 (N_1249,N_789,N_898);
and U1250 (N_1250,N_855,N_686);
nand U1251 (N_1251,N_803,N_961);
nand U1252 (N_1252,N_535,N_637);
or U1253 (N_1253,N_905,N_841);
or U1254 (N_1254,N_861,N_755);
nand U1255 (N_1255,N_964,N_788);
or U1256 (N_1256,N_740,N_590);
or U1257 (N_1257,N_604,N_972);
nand U1258 (N_1258,N_684,N_640);
and U1259 (N_1259,N_678,N_622);
xor U1260 (N_1260,N_558,N_949);
and U1261 (N_1261,N_950,N_976);
and U1262 (N_1262,N_876,N_649);
and U1263 (N_1263,N_831,N_545);
nand U1264 (N_1264,N_961,N_955);
and U1265 (N_1265,N_757,N_540);
nand U1266 (N_1266,N_768,N_836);
nor U1267 (N_1267,N_700,N_828);
or U1268 (N_1268,N_836,N_981);
or U1269 (N_1269,N_955,N_705);
and U1270 (N_1270,N_882,N_885);
nand U1271 (N_1271,N_594,N_568);
nor U1272 (N_1272,N_565,N_617);
xor U1273 (N_1273,N_754,N_666);
nand U1274 (N_1274,N_781,N_697);
or U1275 (N_1275,N_809,N_697);
and U1276 (N_1276,N_720,N_863);
nand U1277 (N_1277,N_501,N_588);
nor U1278 (N_1278,N_823,N_956);
or U1279 (N_1279,N_865,N_805);
xor U1280 (N_1280,N_978,N_587);
xnor U1281 (N_1281,N_748,N_837);
or U1282 (N_1282,N_921,N_785);
and U1283 (N_1283,N_620,N_565);
nor U1284 (N_1284,N_874,N_873);
nor U1285 (N_1285,N_900,N_987);
nand U1286 (N_1286,N_572,N_597);
xor U1287 (N_1287,N_530,N_501);
nand U1288 (N_1288,N_858,N_864);
nor U1289 (N_1289,N_773,N_834);
nand U1290 (N_1290,N_682,N_632);
nand U1291 (N_1291,N_904,N_920);
nor U1292 (N_1292,N_966,N_780);
or U1293 (N_1293,N_891,N_998);
and U1294 (N_1294,N_913,N_893);
nand U1295 (N_1295,N_798,N_719);
or U1296 (N_1296,N_813,N_890);
nand U1297 (N_1297,N_724,N_803);
nand U1298 (N_1298,N_889,N_766);
nand U1299 (N_1299,N_752,N_980);
nor U1300 (N_1300,N_727,N_746);
or U1301 (N_1301,N_824,N_503);
or U1302 (N_1302,N_758,N_575);
and U1303 (N_1303,N_684,N_687);
nand U1304 (N_1304,N_619,N_606);
nand U1305 (N_1305,N_570,N_714);
nor U1306 (N_1306,N_646,N_923);
nor U1307 (N_1307,N_745,N_607);
nor U1308 (N_1308,N_876,N_917);
and U1309 (N_1309,N_691,N_951);
and U1310 (N_1310,N_896,N_825);
and U1311 (N_1311,N_625,N_801);
nor U1312 (N_1312,N_542,N_549);
or U1313 (N_1313,N_878,N_723);
or U1314 (N_1314,N_620,N_719);
and U1315 (N_1315,N_522,N_711);
nand U1316 (N_1316,N_635,N_610);
nand U1317 (N_1317,N_838,N_583);
nor U1318 (N_1318,N_969,N_595);
nor U1319 (N_1319,N_668,N_704);
nor U1320 (N_1320,N_894,N_930);
nand U1321 (N_1321,N_523,N_661);
nand U1322 (N_1322,N_829,N_613);
nor U1323 (N_1323,N_582,N_975);
or U1324 (N_1324,N_634,N_871);
or U1325 (N_1325,N_798,N_959);
or U1326 (N_1326,N_827,N_500);
nor U1327 (N_1327,N_594,N_698);
or U1328 (N_1328,N_630,N_620);
nand U1329 (N_1329,N_548,N_990);
or U1330 (N_1330,N_607,N_857);
nor U1331 (N_1331,N_938,N_875);
nand U1332 (N_1332,N_956,N_783);
nand U1333 (N_1333,N_898,N_582);
and U1334 (N_1334,N_915,N_980);
nand U1335 (N_1335,N_659,N_848);
and U1336 (N_1336,N_978,N_593);
or U1337 (N_1337,N_638,N_774);
or U1338 (N_1338,N_854,N_970);
and U1339 (N_1339,N_695,N_909);
and U1340 (N_1340,N_682,N_563);
nand U1341 (N_1341,N_736,N_974);
or U1342 (N_1342,N_609,N_889);
and U1343 (N_1343,N_549,N_517);
nor U1344 (N_1344,N_670,N_665);
or U1345 (N_1345,N_938,N_960);
nand U1346 (N_1346,N_970,N_968);
nand U1347 (N_1347,N_621,N_965);
nor U1348 (N_1348,N_506,N_918);
and U1349 (N_1349,N_735,N_557);
or U1350 (N_1350,N_534,N_553);
or U1351 (N_1351,N_685,N_903);
nand U1352 (N_1352,N_848,N_732);
or U1353 (N_1353,N_685,N_849);
and U1354 (N_1354,N_526,N_779);
nand U1355 (N_1355,N_650,N_771);
nor U1356 (N_1356,N_984,N_947);
or U1357 (N_1357,N_967,N_709);
nor U1358 (N_1358,N_783,N_860);
nand U1359 (N_1359,N_982,N_512);
nand U1360 (N_1360,N_519,N_762);
nand U1361 (N_1361,N_824,N_888);
or U1362 (N_1362,N_807,N_524);
nand U1363 (N_1363,N_834,N_530);
and U1364 (N_1364,N_806,N_792);
and U1365 (N_1365,N_680,N_572);
nor U1366 (N_1366,N_925,N_745);
nand U1367 (N_1367,N_576,N_628);
or U1368 (N_1368,N_829,N_989);
nand U1369 (N_1369,N_705,N_937);
nand U1370 (N_1370,N_636,N_880);
and U1371 (N_1371,N_823,N_901);
and U1372 (N_1372,N_823,N_671);
and U1373 (N_1373,N_866,N_699);
or U1374 (N_1374,N_802,N_921);
nand U1375 (N_1375,N_654,N_760);
and U1376 (N_1376,N_745,N_887);
and U1377 (N_1377,N_714,N_715);
and U1378 (N_1378,N_580,N_673);
and U1379 (N_1379,N_939,N_745);
and U1380 (N_1380,N_769,N_977);
or U1381 (N_1381,N_846,N_771);
and U1382 (N_1382,N_915,N_810);
nand U1383 (N_1383,N_704,N_694);
nor U1384 (N_1384,N_550,N_739);
and U1385 (N_1385,N_830,N_528);
nand U1386 (N_1386,N_724,N_938);
nor U1387 (N_1387,N_662,N_813);
and U1388 (N_1388,N_720,N_694);
nor U1389 (N_1389,N_795,N_895);
and U1390 (N_1390,N_808,N_721);
or U1391 (N_1391,N_939,N_814);
nand U1392 (N_1392,N_729,N_999);
or U1393 (N_1393,N_995,N_544);
nand U1394 (N_1394,N_532,N_564);
or U1395 (N_1395,N_739,N_676);
nor U1396 (N_1396,N_796,N_674);
xor U1397 (N_1397,N_741,N_759);
nor U1398 (N_1398,N_786,N_994);
nor U1399 (N_1399,N_535,N_698);
nor U1400 (N_1400,N_574,N_965);
nor U1401 (N_1401,N_977,N_863);
or U1402 (N_1402,N_834,N_774);
nand U1403 (N_1403,N_726,N_802);
nand U1404 (N_1404,N_936,N_520);
nor U1405 (N_1405,N_674,N_914);
nor U1406 (N_1406,N_940,N_749);
or U1407 (N_1407,N_723,N_615);
nor U1408 (N_1408,N_990,N_885);
nor U1409 (N_1409,N_676,N_810);
and U1410 (N_1410,N_741,N_771);
and U1411 (N_1411,N_841,N_663);
and U1412 (N_1412,N_675,N_824);
and U1413 (N_1413,N_814,N_561);
nor U1414 (N_1414,N_759,N_846);
or U1415 (N_1415,N_725,N_556);
or U1416 (N_1416,N_614,N_701);
nand U1417 (N_1417,N_994,N_987);
nand U1418 (N_1418,N_589,N_732);
nor U1419 (N_1419,N_994,N_812);
or U1420 (N_1420,N_786,N_703);
and U1421 (N_1421,N_666,N_723);
and U1422 (N_1422,N_793,N_564);
or U1423 (N_1423,N_808,N_520);
or U1424 (N_1424,N_856,N_637);
nand U1425 (N_1425,N_984,N_963);
nand U1426 (N_1426,N_993,N_659);
or U1427 (N_1427,N_879,N_741);
and U1428 (N_1428,N_826,N_692);
nand U1429 (N_1429,N_995,N_976);
nand U1430 (N_1430,N_719,N_594);
and U1431 (N_1431,N_844,N_948);
or U1432 (N_1432,N_524,N_766);
and U1433 (N_1433,N_793,N_526);
xor U1434 (N_1434,N_787,N_780);
nand U1435 (N_1435,N_737,N_821);
and U1436 (N_1436,N_930,N_607);
or U1437 (N_1437,N_943,N_683);
or U1438 (N_1438,N_529,N_902);
and U1439 (N_1439,N_898,N_902);
and U1440 (N_1440,N_938,N_713);
nor U1441 (N_1441,N_798,N_954);
and U1442 (N_1442,N_857,N_601);
nand U1443 (N_1443,N_782,N_822);
and U1444 (N_1444,N_619,N_978);
nand U1445 (N_1445,N_934,N_536);
or U1446 (N_1446,N_992,N_558);
and U1447 (N_1447,N_968,N_814);
nand U1448 (N_1448,N_588,N_777);
nor U1449 (N_1449,N_738,N_799);
nor U1450 (N_1450,N_547,N_907);
nand U1451 (N_1451,N_762,N_692);
and U1452 (N_1452,N_569,N_654);
nor U1453 (N_1453,N_638,N_954);
nor U1454 (N_1454,N_857,N_536);
nand U1455 (N_1455,N_784,N_637);
and U1456 (N_1456,N_889,N_939);
and U1457 (N_1457,N_722,N_755);
and U1458 (N_1458,N_785,N_803);
nor U1459 (N_1459,N_769,N_767);
nand U1460 (N_1460,N_605,N_788);
nor U1461 (N_1461,N_877,N_773);
nand U1462 (N_1462,N_990,N_790);
or U1463 (N_1463,N_957,N_812);
or U1464 (N_1464,N_867,N_810);
nor U1465 (N_1465,N_734,N_666);
and U1466 (N_1466,N_945,N_960);
and U1467 (N_1467,N_978,N_937);
nand U1468 (N_1468,N_614,N_849);
nand U1469 (N_1469,N_925,N_594);
nand U1470 (N_1470,N_617,N_860);
and U1471 (N_1471,N_692,N_717);
and U1472 (N_1472,N_900,N_818);
nand U1473 (N_1473,N_739,N_797);
and U1474 (N_1474,N_509,N_810);
or U1475 (N_1475,N_711,N_838);
nor U1476 (N_1476,N_711,N_979);
or U1477 (N_1477,N_634,N_934);
or U1478 (N_1478,N_596,N_911);
nand U1479 (N_1479,N_590,N_923);
nand U1480 (N_1480,N_645,N_626);
and U1481 (N_1481,N_767,N_626);
nor U1482 (N_1482,N_788,N_980);
nor U1483 (N_1483,N_823,N_860);
nor U1484 (N_1484,N_742,N_861);
nor U1485 (N_1485,N_797,N_577);
or U1486 (N_1486,N_635,N_796);
and U1487 (N_1487,N_650,N_664);
nand U1488 (N_1488,N_835,N_785);
or U1489 (N_1489,N_865,N_674);
nor U1490 (N_1490,N_516,N_542);
nor U1491 (N_1491,N_961,N_651);
nor U1492 (N_1492,N_877,N_631);
nand U1493 (N_1493,N_970,N_528);
nand U1494 (N_1494,N_905,N_542);
nand U1495 (N_1495,N_689,N_586);
and U1496 (N_1496,N_545,N_839);
nor U1497 (N_1497,N_949,N_786);
nand U1498 (N_1498,N_819,N_944);
nand U1499 (N_1499,N_684,N_663);
nand U1500 (N_1500,N_1218,N_1329);
and U1501 (N_1501,N_1306,N_1336);
or U1502 (N_1502,N_1090,N_1432);
nand U1503 (N_1503,N_1350,N_1077);
and U1504 (N_1504,N_1443,N_1304);
nand U1505 (N_1505,N_1370,N_1495);
or U1506 (N_1506,N_1316,N_1011);
nand U1507 (N_1507,N_1382,N_1444);
nand U1508 (N_1508,N_1481,N_1157);
and U1509 (N_1509,N_1395,N_1486);
nand U1510 (N_1510,N_1437,N_1371);
and U1511 (N_1511,N_1222,N_1409);
or U1512 (N_1512,N_1080,N_1039);
nor U1513 (N_1513,N_1297,N_1285);
or U1514 (N_1514,N_1431,N_1394);
nand U1515 (N_1515,N_1254,N_1472);
nand U1516 (N_1516,N_1128,N_1348);
nand U1517 (N_1517,N_1386,N_1459);
nor U1518 (N_1518,N_1347,N_1092);
nor U1519 (N_1519,N_1230,N_1019);
or U1520 (N_1520,N_1428,N_1118);
nand U1521 (N_1521,N_1260,N_1105);
nor U1522 (N_1522,N_1047,N_1462);
nand U1523 (N_1523,N_1295,N_1342);
nand U1524 (N_1524,N_1068,N_1126);
and U1525 (N_1525,N_1467,N_1102);
nand U1526 (N_1526,N_1429,N_1263);
or U1527 (N_1527,N_1399,N_1108);
or U1528 (N_1528,N_1272,N_1470);
or U1529 (N_1529,N_1076,N_1176);
or U1530 (N_1530,N_1416,N_1216);
nand U1531 (N_1531,N_1026,N_1138);
and U1532 (N_1532,N_1168,N_1145);
and U1533 (N_1533,N_1283,N_1156);
or U1534 (N_1534,N_1065,N_1403);
nand U1535 (N_1535,N_1383,N_1369);
nor U1536 (N_1536,N_1447,N_1318);
nor U1537 (N_1537,N_1086,N_1322);
xnor U1538 (N_1538,N_1130,N_1478);
and U1539 (N_1539,N_1171,N_1335);
nor U1540 (N_1540,N_1441,N_1129);
or U1541 (N_1541,N_1485,N_1004);
or U1542 (N_1542,N_1420,N_1220);
and U1543 (N_1543,N_1286,N_1031);
and U1544 (N_1544,N_1417,N_1192);
or U1545 (N_1545,N_1046,N_1379);
nand U1546 (N_1546,N_1007,N_1387);
nor U1547 (N_1547,N_1201,N_1185);
nand U1548 (N_1548,N_1411,N_1357);
and U1549 (N_1549,N_1334,N_1498);
and U1550 (N_1550,N_1235,N_1361);
and U1551 (N_1551,N_1036,N_1359);
or U1552 (N_1552,N_1255,N_1404);
nand U1553 (N_1553,N_1410,N_1212);
or U1554 (N_1554,N_1231,N_1292);
or U1555 (N_1555,N_1057,N_1389);
and U1556 (N_1556,N_1089,N_1005);
and U1557 (N_1557,N_1349,N_1035);
nand U1558 (N_1558,N_1023,N_1490);
nand U1559 (N_1559,N_1025,N_1343);
nand U1560 (N_1560,N_1071,N_1198);
nand U1561 (N_1561,N_1209,N_1173);
nand U1562 (N_1562,N_1480,N_1450);
xor U1563 (N_1563,N_1058,N_1225);
nand U1564 (N_1564,N_1406,N_1043);
nor U1565 (N_1565,N_1033,N_1149);
nand U1566 (N_1566,N_1448,N_1160);
nand U1567 (N_1567,N_1120,N_1471);
nor U1568 (N_1568,N_1390,N_1119);
and U1569 (N_1569,N_1139,N_1328);
nor U1570 (N_1570,N_1414,N_1484);
nor U1571 (N_1571,N_1352,N_1083);
nor U1572 (N_1572,N_1113,N_1017);
nand U1573 (N_1573,N_1158,N_1264);
nand U1574 (N_1574,N_1008,N_1003);
or U1575 (N_1575,N_1240,N_1466);
nor U1576 (N_1576,N_1131,N_1476);
nand U1577 (N_1577,N_1075,N_1331);
nand U1578 (N_1578,N_1360,N_1069);
and U1579 (N_1579,N_1020,N_1166);
and U1580 (N_1580,N_1274,N_1141);
and U1581 (N_1581,N_1084,N_1238);
and U1582 (N_1582,N_1186,N_1296);
nand U1583 (N_1583,N_1356,N_1364);
and U1584 (N_1584,N_1473,N_1294);
and U1585 (N_1585,N_1167,N_1125);
or U1586 (N_1586,N_1082,N_1140);
nand U1587 (N_1587,N_1422,N_1375);
or U1588 (N_1588,N_1207,N_1165);
or U1589 (N_1589,N_1271,N_1345);
nand U1590 (N_1590,N_1363,N_1170);
or U1591 (N_1591,N_1204,N_1062);
nor U1592 (N_1592,N_1232,N_1457);
nor U1593 (N_1593,N_1028,N_1049);
or U1594 (N_1594,N_1266,N_1172);
and U1595 (N_1595,N_1147,N_1016);
xnor U1596 (N_1596,N_1305,N_1340);
or U1597 (N_1597,N_1099,N_1491);
and U1598 (N_1598,N_1440,N_1096);
nor U1599 (N_1599,N_1194,N_1373);
nand U1600 (N_1600,N_1353,N_1407);
nand U1601 (N_1601,N_1034,N_1116);
nor U1602 (N_1602,N_1135,N_1152);
xor U1603 (N_1603,N_1132,N_1018);
nor U1604 (N_1604,N_1405,N_1001);
or U1605 (N_1605,N_1110,N_1236);
or U1606 (N_1606,N_1246,N_1270);
and U1607 (N_1607,N_1163,N_1122);
nand U1608 (N_1608,N_1079,N_1427);
nor U1609 (N_1609,N_1307,N_1268);
and U1610 (N_1610,N_1205,N_1433);
and U1611 (N_1611,N_1104,N_1257);
or U1612 (N_1612,N_1070,N_1402);
nor U1613 (N_1613,N_1048,N_1449);
nand U1614 (N_1614,N_1468,N_1134);
nand U1615 (N_1615,N_1400,N_1469);
nand U1616 (N_1616,N_1107,N_1208);
xnor U1617 (N_1617,N_1464,N_1434);
nor U1618 (N_1618,N_1234,N_1446);
and U1619 (N_1619,N_1436,N_1398);
and U1620 (N_1620,N_1299,N_1127);
and U1621 (N_1621,N_1064,N_1275);
nand U1622 (N_1622,N_1267,N_1453);
and U1623 (N_1623,N_1325,N_1174);
nor U1624 (N_1624,N_1248,N_1324);
or U1625 (N_1625,N_1239,N_1426);
nand U1626 (N_1626,N_1136,N_1044);
or U1627 (N_1627,N_1150,N_1009);
xnor U1628 (N_1628,N_1094,N_1237);
or U1629 (N_1629,N_1475,N_1042);
nand U1630 (N_1630,N_1377,N_1376);
nand U1631 (N_1631,N_1032,N_1121);
and U1632 (N_1632,N_1424,N_1269);
and U1633 (N_1633,N_1000,N_1095);
and U1634 (N_1634,N_1451,N_1124);
nor U1635 (N_1635,N_1227,N_1323);
nand U1636 (N_1636,N_1053,N_1060);
nand U1637 (N_1637,N_1279,N_1455);
nand U1638 (N_1638,N_1488,N_1418);
or U1639 (N_1639,N_1067,N_1245);
or U1640 (N_1640,N_1252,N_1249);
and U1641 (N_1641,N_1159,N_1351);
and U1642 (N_1642,N_1372,N_1063);
and U1643 (N_1643,N_1114,N_1430);
nor U1644 (N_1644,N_1061,N_1259);
and U1645 (N_1645,N_1337,N_1193);
and U1646 (N_1646,N_1423,N_1038);
and U1647 (N_1647,N_1261,N_1045);
nor U1648 (N_1648,N_1210,N_1052);
or U1649 (N_1649,N_1393,N_1213);
nor U1650 (N_1650,N_1056,N_1041);
nand U1651 (N_1651,N_1384,N_1396);
xor U1652 (N_1652,N_1233,N_1288);
and U1653 (N_1653,N_1435,N_1326);
nand U1654 (N_1654,N_1146,N_1106);
or U1655 (N_1655,N_1487,N_1445);
and U1656 (N_1656,N_1197,N_1415);
or U1657 (N_1657,N_1091,N_1298);
nand U1658 (N_1658,N_1226,N_1101);
nand U1659 (N_1659,N_1289,N_1002);
or U1660 (N_1660,N_1211,N_1228);
and U1661 (N_1661,N_1262,N_1380);
nand U1662 (N_1662,N_1184,N_1365);
and U1663 (N_1663,N_1494,N_1425);
nand U1664 (N_1664,N_1169,N_1314);
nor U1665 (N_1665,N_1300,N_1273);
and U1666 (N_1666,N_1179,N_1217);
nand U1667 (N_1667,N_1155,N_1059);
nand U1668 (N_1668,N_1477,N_1315);
nor U1669 (N_1669,N_1022,N_1175);
nand U1670 (N_1670,N_1392,N_1109);
and U1671 (N_1671,N_1482,N_1489);
or U1672 (N_1672,N_1085,N_1200);
or U1673 (N_1673,N_1180,N_1281);
and U1674 (N_1674,N_1479,N_1241);
nor U1675 (N_1675,N_1247,N_1242);
nand U1676 (N_1676,N_1111,N_1293);
or U1677 (N_1677,N_1278,N_1301);
nand U1678 (N_1678,N_1178,N_1374);
nand U1679 (N_1679,N_1311,N_1013);
nand U1680 (N_1680,N_1339,N_1188);
or U1681 (N_1681,N_1073,N_1143);
nor U1682 (N_1682,N_1421,N_1381);
or U1683 (N_1683,N_1051,N_1330);
or U1684 (N_1684,N_1302,N_1066);
or U1685 (N_1685,N_1358,N_1460);
nand U1686 (N_1686,N_1313,N_1312);
and U1687 (N_1687,N_1215,N_1253);
or U1688 (N_1688,N_1177,N_1303);
nor U1689 (N_1689,N_1072,N_1088);
nor U1690 (N_1690,N_1319,N_1203);
and U1691 (N_1691,N_1093,N_1137);
xor U1692 (N_1692,N_1277,N_1492);
and U1693 (N_1693,N_1117,N_1148);
nand U1694 (N_1694,N_1251,N_1265);
nand U1695 (N_1695,N_1181,N_1401);
and U1696 (N_1696,N_1219,N_1142);
nor U1697 (N_1697,N_1256,N_1112);
nand U1698 (N_1698,N_1103,N_1320);
nor U1699 (N_1699,N_1327,N_1452);
nand U1700 (N_1700,N_1244,N_1413);
nor U1701 (N_1701,N_1442,N_1123);
and U1702 (N_1702,N_1321,N_1182);
or U1703 (N_1703,N_1202,N_1412);
or U1704 (N_1704,N_1287,N_1054);
or U1705 (N_1705,N_1087,N_1497);
and U1706 (N_1706,N_1317,N_1378);
and U1707 (N_1707,N_1229,N_1190);
nand U1708 (N_1708,N_1100,N_1458);
and U1709 (N_1709,N_1367,N_1037);
and U1710 (N_1710,N_1354,N_1474);
nand U1711 (N_1711,N_1223,N_1362);
or U1712 (N_1712,N_1346,N_1098);
and U1713 (N_1713,N_1456,N_1133);
nor U1714 (N_1714,N_1397,N_1154);
nor U1715 (N_1715,N_1014,N_1221);
and U1716 (N_1716,N_1162,N_1015);
and U1717 (N_1717,N_1164,N_1214);
nor U1718 (N_1718,N_1027,N_1191);
or U1719 (N_1719,N_1408,N_1183);
nand U1720 (N_1720,N_1290,N_1368);
and U1721 (N_1721,N_1010,N_1385);
nor U1722 (N_1722,N_1199,N_1040);
nand U1723 (N_1723,N_1366,N_1308);
or U1724 (N_1724,N_1461,N_1338);
nand U1725 (N_1725,N_1024,N_1499);
nor U1726 (N_1726,N_1074,N_1006);
or U1727 (N_1727,N_1050,N_1030);
nand U1728 (N_1728,N_1332,N_1224);
nor U1729 (N_1729,N_1097,N_1151);
and U1730 (N_1730,N_1196,N_1284);
and U1731 (N_1731,N_1078,N_1189);
and U1732 (N_1732,N_1153,N_1454);
or U1733 (N_1733,N_1465,N_1206);
nand U1734 (N_1734,N_1438,N_1344);
or U1735 (N_1735,N_1493,N_1310);
nand U1736 (N_1736,N_1161,N_1280);
nand U1737 (N_1737,N_1243,N_1081);
nand U1738 (N_1738,N_1463,N_1439);
nor U1739 (N_1739,N_1483,N_1021);
nor U1740 (N_1740,N_1258,N_1388);
or U1741 (N_1741,N_1144,N_1419);
nand U1742 (N_1742,N_1276,N_1341);
or U1743 (N_1743,N_1012,N_1391);
and U1744 (N_1744,N_1029,N_1115);
nor U1745 (N_1745,N_1055,N_1496);
or U1746 (N_1746,N_1333,N_1291);
and U1747 (N_1747,N_1195,N_1355);
nor U1748 (N_1748,N_1250,N_1282);
nand U1749 (N_1749,N_1309,N_1187);
nand U1750 (N_1750,N_1434,N_1008);
and U1751 (N_1751,N_1474,N_1212);
or U1752 (N_1752,N_1086,N_1149);
nand U1753 (N_1753,N_1053,N_1384);
and U1754 (N_1754,N_1105,N_1094);
nand U1755 (N_1755,N_1009,N_1083);
nand U1756 (N_1756,N_1288,N_1243);
and U1757 (N_1757,N_1020,N_1051);
nand U1758 (N_1758,N_1475,N_1367);
and U1759 (N_1759,N_1073,N_1065);
nand U1760 (N_1760,N_1461,N_1103);
nand U1761 (N_1761,N_1261,N_1018);
nor U1762 (N_1762,N_1466,N_1238);
and U1763 (N_1763,N_1024,N_1395);
or U1764 (N_1764,N_1174,N_1052);
nor U1765 (N_1765,N_1360,N_1029);
nor U1766 (N_1766,N_1285,N_1050);
and U1767 (N_1767,N_1384,N_1171);
nand U1768 (N_1768,N_1348,N_1407);
or U1769 (N_1769,N_1303,N_1051);
or U1770 (N_1770,N_1190,N_1478);
and U1771 (N_1771,N_1067,N_1447);
and U1772 (N_1772,N_1320,N_1307);
and U1773 (N_1773,N_1308,N_1275);
nor U1774 (N_1774,N_1104,N_1484);
and U1775 (N_1775,N_1441,N_1284);
or U1776 (N_1776,N_1233,N_1133);
or U1777 (N_1777,N_1213,N_1416);
and U1778 (N_1778,N_1257,N_1010);
nand U1779 (N_1779,N_1114,N_1199);
and U1780 (N_1780,N_1124,N_1144);
nand U1781 (N_1781,N_1439,N_1489);
and U1782 (N_1782,N_1422,N_1136);
or U1783 (N_1783,N_1152,N_1336);
or U1784 (N_1784,N_1264,N_1326);
nand U1785 (N_1785,N_1327,N_1208);
xor U1786 (N_1786,N_1178,N_1260);
nor U1787 (N_1787,N_1323,N_1223);
nand U1788 (N_1788,N_1238,N_1010);
and U1789 (N_1789,N_1016,N_1256);
nand U1790 (N_1790,N_1310,N_1448);
or U1791 (N_1791,N_1303,N_1265);
or U1792 (N_1792,N_1002,N_1058);
nand U1793 (N_1793,N_1459,N_1325);
and U1794 (N_1794,N_1128,N_1277);
and U1795 (N_1795,N_1023,N_1398);
or U1796 (N_1796,N_1417,N_1013);
and U1797 (N_1797,N_1155,N_1188);
and U1798 (N_1798,N_1167,N_1473);
xnor U1799 (N_1799,N_1023,N_1325);
and U1800 (N_1800,N_1203,N_1412);
nand U1801 (N_1801,N_1271,N_1132);
nand U1802 (N_1802,N_1028,N_1432);
nand U1803 (N_1803,N_1028,N_1333);
and U1804 (N_1804,N_1200,N_1030);
or U1805 (N_1805,N_1020,N_1304);
nor U1806 (N_1806,N_1428,N_1145);
or U1807 (N_1807,N_1378,N_1245);
and U1808 (N_1808,N_1181,N_1459);
or U1809 (N_1809,N_1134,N_1256);
xnor U1810 (N_1810,N_1080,N_1178);
or U1811 (N_1811,N_1321,N_1193);
nand U1812 (N_1812,N_1483,N_1283);
or U1813 (N_1813,N_1074,N_1004);
or U1814 (N_1814,N_1191,N_1302);
and U1815 (N_1815,N_1087,N_1435);
nand U1816 (N_1816,N_1422,N_1059);
and U1817 (N_1817,N_1321,N_1212);
or U1818 (N_1818,N_1116,N_1327);
nor U1819 (N_1819,N_1176,N_1077);
and U1820 (N_1820,N_1150,N_1360);
and U1821 (N_1821,N_1151,N_1407);
nand U1822 (N_1822,N_1056,N_1072);
and U1823 (N_1823,N_1469,N_1160);
and U1824 (N_1824,N_1122,N_1012);
nand U1825 (N_1825,N_1248,N_1412);
or U1826 (N_1826,N_1304,N_1302);
or U1827 (N_1827,N_1477,N_1485);
or U1828 (N_1828,N_1026,N_1195);
nand U1829 (N_1829,N_1123,N_1467);
nor U1830 (N_1830,N_1272,N_1096);
or U1831 (N_1831,N_1357,N_1257);
and U1832 (N_1832,N_1378,N_1279);
xor U1833 (N_1833,N_1318,N_1274);
nor U1834 (N_1834,N_1080,N_1029);
nand U1835 (N_1835,N_1027,N_1329);
or U1836 (N_1836,N_1151,N_1176);
or U1837 (N_1837,N_1482,N_1438);
nand U1838 (N_1838,N_1210,N_1042);
or U1839 (N_1839,N_1217,N_1119);
or U1840 (N_1840,N_1478,N_1420);
nand U1841 (N_1841,N_1178,N_1134);
nor U1842 (N_1842,N_1467,N_1448);
and U1843 (N_1843,N_1146,N_1090);
nor U1844 (N_1844,N_1242,N_1040);
nand U1845 (N_1845,N_1463,N_1297);
and U1846 (N_1846,N_1111,N_1475);
nor U1847 (N_1847,N_1352,N_1265);
xnor U1848 (N_1848,N_1088,N_1390);
nor U1849 (N_1849,N_1336,N_1338);
or U1850 (N_1850,N_1043,N_1220);
or U1851 (N_1851,N_1205,N_1423);
nor U1852 (N_1852,N_1290,N_1114);
and U1853 (N_1853,N_1236,N_1282);
and U1854 (N_1854,N_1126,N_1031);
nor U1855 (N_1855,N_1284,N_1382);
nor U1856 (N_1856,N_1376,N_1023);
nor U1857 (N_1857,N_1205,N_1007);
and U1858 (N_1858,N_1098,N_1316);
nor U1859 (N_1859,N_1191,N_1121);
or U1860 (N_1860,N_1381,N_1451);
nor U1861 (N_1861,N_1497,N_1219);
or U1862 (N_1862,N_1434,N_1045);
nand U1863 (N_1863,N_1101,N_1256);
and U1864 (N_1864,N_1314,N_1399);
or U1865 (N_1865,N_1326,N_1062);
and U1866 (N_1866,N_1326,N_1068);
and U1867 (N_1867,N_1116,N_1455);
nor U1868 (N_1868,N_1135,N_1394);
and U1869 (N_1869,N_1462,N_1005);
nor U1870 (N_1870,N_1223,N_1241);
nor U1871 (N_1871,N_1313,N_1438);
nor U1872 (N_1872,N_1391,N_1229);
or U1873 (N_1873,N_1234,N_1295);
nor U1874 (N_1874,N_1332,N_1453);
nand U1875 (N_1875,N_1247,N_1209);
and U1876 (N_1876,N_1417,N_1015);
and U1877 (N_1877,N_1218,N_1105);
nor U1878 (N_1878,N_1199,N_1180);
nand U1879 (N_1879,N_1034,N_1374);
and U1880 (N_1880,N_1395,N_1412);
or U1881 (N_1881,N_1353,N_1343);
nand U1882 (N_1882,N_1220,N_1279);
or U1883 (N_1883,N_1158,N_1428);
or U1884 (N_1884,N_1112,N_1290);
and U1885 (N_1885,N_1048,N_1143);
nand U1886 (N_1886,N_1036,N_1301);
and U1887 (N_1887,N_1156,N_1417);
nand U1888 (N_1888,N_1487,N_1462);
nand U1889 (N_1889,N_1337,N_1082);
nand U1890 (N_1890,N_1218,N_1323);
or U1891 (N_1891,N_1180,N_1090);
nand U1892 (N_1892,N_1492,N_1054);
or U1893 (N_1893,N_1164,N_1454);
nor U1894 (N_1894,N_1052,N_1166);
and U1895 (N_1895,N_1002,N_1004);
and U1896 (N_1896,N_1192,N_1057);
nand U1897 (N_1897,N_1033,N_1335);
and U1898 (N_1898,N_1064,N_1268);
nand U1899 (N_1899,N_1022,N_1359);
nor U1900 (N_1900,N_1101,N_1339);
and U1901 (N_1901,N_1125,N_1242);
nor U1902 (N_1902,N_1030,N_1251);
nand U1903 (N_1903,N_1478,N_1314);
nor U1904 (N_1904,N_1216,N_1260);
nor U1905 (N_1905,N_1110,N_1368);
nor U1906 (N_1906,N_1018,N_1113);
and U1907 (N_1907,N_1372,N_1489);
nand U1908 (N_1908,N_1160,N_1074);
or U1909 (N_1909,N_1085,N_1060);
nand U1910 (N_1910,N_1232,N_1253);
and U1911 (N_1911,N_1376,N_1474);
and U1912 (N_1912,N_1460,N_1381);
nand U1913 (N_1913,N_1417,N_1171);
or U1914 (N_1914,N_1153,N_1387);
and U1915 (N_1915,N_1210,N_1306);
and U1916 (N_1916,N_1070,N_1157);
and U1917 (N_1917,N_1277,N_1452);
nor U1918 (N_1918,N_1474,N_1158);
nor U1919 (N_1919,N_1455,N_1260);
or U1920 (N_1920,N_1299,N_1407);
nor U1921 (N_1921,N_1421,N_1490);
and U1922 (N_1922,N_1383,N_1429);
or U1923 (N_1923,N_1047,N_1346);
nor U1924 (N_1924,N_1097,N_1406);
nor U1925 (N_1925,N_1140,N_1055);
nand U1926 (N_1926,N_1424,N_1430);
nand U1927 (N_1927,N_1196,N_1180);
and U1928 (N_1928,N_1381,N_1423);
or U1929 (N_1929,N_1318,N_1371);
or U1930 (N_1930,N_1208,N_1478);
or U1931 (N_1931,N_1069,N_1015);
nor U1932 (N_1932,N_1013,N_1211);
xor U1933 (N_1933,N_1172,N_1141);
nor U1934 (N_1934,N_1450,N_1291);
or U1935 (N_1935,N_1109,N_1396);
nor U1936 (N_1936,N_1047,N_1159);
and U1937 (N_1937,N_1148,N_1459);
and U1938 (N_1938,N_1155,N_1157);
or U1939 (N_1939,N_1146,N_1484);
nor U1940 (N_1940,N_1216,N_1062);
or U1941 (N_1941,N_1132,N_1149);
nand U1942 (N_1942,N_1300,N_1473);
or U1943 (N_1943,N_1181,N_1477);
and U1944 (N_1944,N_1003,N_1141);
nor U1945 (N_1945,N_1081,N_1046);
and U1946 (N_1946,N_1438,N_1226);
nor U1947 (N_1947,N_1326,N_1338);
or U1948 (N_1948,N_1299,N_1000);
nand U1949 (N_1949,N_1135,N_1058);
nor U1950 (N_1950,N_1022,N_1322);
nor U1951 (N_1951,N_1429,N_1066);
nand U1952 (N_1952,N_1172,N_1046);
nor U1953 (N_1953,N_1104,N_1111);
and U1954 (N_1954,N_1272,N_1319);
nand U1955 (N_1955,N_1426,N_1256);
xnor U1956 (N_1956,N_1330,N_1298);
xnor U1957 (N_1957,N_1153,N_1207);
or U1958 (N_1958,N_1417,N_1321);
or U1959 (N_1959,N_1267,N_1257);
or U1960 (N_1960,N_1265,N_1342);
nor U1961 (N_1961,N_1344,N_1231);
or U1962 (N_1962,N_1450,N_1078);
or U1963 (N_1963,N_1156,N_1346);
or U1964 (N_1964,N_1162,N_1335);
or U1965 (N_1965,N_1124,N_1046);
and U1966 (N_1966,N_1332,N_1223);
or U1967 (N_1967,N_1432,N_1403);
nor U1968 (N_1968,N_1319,N_1346);
nand U1969 (N_1969,N_1492,N_1274);
nand U1970 (N_1970,N_1490,N_1111);
nor U1971 (N_1971,N_1106,N_1305);
and U1972 (N_1972,N_1495,N_1196);
or U1973 (N_1973,N_1061,N_1047);
or U1974 (N_1974,N_1458,N_1070);
and U1975 (N_1975,N_1001,N_1185);
xor U1976 (N_1976,N_1282,N_1324);
nor U1977 (N_1977,N_1280,N_1426);
nor U1978 (N_1978,N_1115,N_1444);
or U1979 (N_1979,N_1241,N_1348);
or U1980 (N_1980,N_1229,N_1431);
or U1981 (N_1981,N_1323,N_1040);
and U1982 (N_1982,N_1358,N_1451);
and U1983 (N_1983,N_1277,N_1159);
nand U1984 (N_1984,N_1250,N_1154);
nor U1985 (N_1985,N_1321,N_1396);
or U1986 (N_1986,N_1433,N_1209);
or U1987 (N_1987,N_1423,N_1474);
nand U1988 (N_1988,N_1219,N_1292);
and U1989 (N_1989,N_1125,N_1323);
nand U1990 (N_1990,N_1094,N_1252);
and U1991 (N_1991,N_1486,N_1379);
nor U1992 (N_1992,N_1432,N_1334);
and U1993 (N_1993,N_1278,N_1443);
nor U1994 (N_1994,N_1178,N_1201);
or U1995 (N_1995,N_1357,N_1319);
or U1996 (N_1996,N_1259,N_1367);
and U1997 (N_1997,N_1204,N_1205);
or U1998 (N_1998,N_1068,N_1014);
nand U1999 (N_1999,N_1086,N_1276);
or U2000 (N_2000,N_1698,N_1719);
nand U2001 (N_2001,N_1588,N_1567);
and U2002 (N_2002,N_1653,N_1909);
nor U2003 (N_2003,N_1918,N_1949);
or U2004 (N_2004,N_1657,N_1895);
nor U2005 (N_2005,N_1649,N_1961);
and U2006 (N_2006,N_1855,N_1634);
nor U2007 (N_2007,N_1627,N_1973);
and U2008 (N_2008,N_1507,N_1888);
nand U2009 (N_2009,N_1839,N_1752);
or U2010 (N_2010,N_1705,N_1534);
and U2011 (N_2011,N_1584,N_1622);
nor U2012 (N_2012,N_1645,N_1632);
nand U2013 (N_2013,N_1546,N_1820);
or U2014 (N_2014,N_1970,N_1896);
nand U2015 (N_2015,N_1658,N_1654);
or U2016 (N_2016,N_1718,N_1757);
or U2017 (N_2017,N_1984,N_1730);
nor U2018 (N_2018,N_1945,N_1514);
nor U2019 (N_2019,N_1942,N_1762);
nor U2020 (N_2020,N_1799,N_1966);
or U2021 (N_2021,N_1607,N_1613);
nor U2022 (N_2022,N_1569,N_1579);
or U2023 (N_2023,N_1749,N_1593);
nand U2024 (N_2024,N_1781,N_1891);
and U2025 (N_2025,N_1813,N_1732);
nand U2026 (N_2026,N_1796,N_1672);
nor U2027 (N_2027,N_1722,N_1667);
nand U2028 (N_2028,N_1916,N_1520);
or U2029 (N_2029,N_1755,N_1625);
or U2030 (N_2030,N_1518,N_1544);
nand U2031 (N_2031,N_1501,N_1955);
and U2032 (N_2032,N_1990,N_1929);
or U2033 (N_2033,N_1884,N_1596);
and U2034 (N_2034,N_1852,N_1858);
or U2035 (N_2035,N_1801,N_1582);
nor U2036 (N_2036,N_1992,N_1874);
or U2037 (N_2037,N_1951,N_1890);
or U2038 (N_2038,N_1617,N_1822);
nand U2039 (N_2039,N_1577,N_1527);
or U2040 (N_2040,N_1859,N_1807);
or U2041 (N_2041,N_1530,N_1702);
nor U2042 (N_2042,N_1686,N_1805);
nor U2043 (N_2043,N_1797,N_1887);
nand U2044 (N_2044,N_1503,N_1690);
nand U2045 (N_2045,N_1581,N_1892);
nand U2046 (N_2046,N_1950,N_1713);
or U2047 (N_2047,N_1597,N_1798);
nand U2048 (N_2048,N_1944,N_1599);
nand U2049 (N_2049,N_1900,N_1865);
nor U2050 (N_2050,N_1985,N_1862);
nor U2051 (N_2051,N_1656,N_1703);
nor U2052 (N_2052,N_1628,N_1671);
nor U2053 (N_2053,N_1793,N_1898);
nor U2054 (N_2054,N_1812,N_1742);
nor U2055 (N_2055,N_1693,N_1754);
and U2056 (N_2056,N_1772,N_1743);
nand U2057 (N_2057,N_1689,N_1572);
and U2058 (N_2058,N_1739,N_1775);
and U2059 (N_2059,N_1996,N_1914);
nor U2060 (N_2060,N_1924,N_1678);
and U2061 (N_2061,N_1894,N_1647);
nor U2062 (N_2062,N_1897,N_1525);
nor U2063 (N_2063,N_1776,N_1523);
and U2064 (N_2064,N_1592,N_1779);
or U2065 (N_2065,N_1965,N_1631);
nor U2066 (N_2066,N_1790,N_1680);
and U2067 (N_2067,N_1674,N_1731);
or U2068 (N_2068,N_1921,N_1922);
and U2069 (N_2069,N_1866,N_1991);
nor U2070 (N_2070,N_1619,N_1972);
or U2071 (N_2071,N_1928,N_1711);
nand U2072 (N_2072,N_1681,N_1975);
nand U2073 (N_2073,N_1727,N_1747);
nor U2074 (N_2074,N_1877,N_1623);
or U2075 (N_2075,N_1948,N_1587);
nand U2076 (N_2076,N_1880,N_1676);
nor U2077 (N_2077,N_1978,N_1517);
or U2078 (N_2078,N_1552,N_1618);
or U2079 (N_2079,N_1737,N_1833);
or U2080 (N_2080,N_1923,N_1953);
nand U2081 (N_2081,N_1506,N_1856);
xnor U2082 (N_2082,N_1765,N_1920);
nand U2083 (N_2083,N_1560,N_1557);
nor U2084 (N_2084,N_1620,N_1559);
and U2085 (N_2085,N_1659,N_1626);
and U2086 (N_2086,N_1729,N_1815);
or U2087 (N_2087,N_1967,N_1751);
or U2088 (N_2088,N_1769,N_1802);
and U2089 (N_2089,N_1995,N_1652);
or U2090 (N_2090,N_1930,N_1870);
and U2091 (N_2091,N_1899,N_1778);
or U2092 (N_2092,N_1960,N_1511);
or U2093 (N_2093,N_1881,N_1907);
nor U2094 (N_2094,N_1787,N_1646);
nor U2095 (N_2095,N_1882,N_1906);
nor U2096 (N_2096,N_1533,N_1806);
xnor U2097 (N_2097,N_1639,N_1688);
and U2098 (N_2098,N_1509,N_1675);
nor U2099 (N_2099,N_1771,N_1564);
nand U2100 (N_2100,N_1963,N_1694);
nor U2101 (N_2101,N_1933,N_1700);
nor U2102 (N_2102,N_1935,N_1981);
nand U2103 (N_2103,N_1666,N_1554);
and U2104 (N_2104,N_1635,N_1829);
nand U2105 (N_2105,N_1699,N_1784);
nor U2106 (N_2106,N_1911,N_1828);
nand U2107 (N_2107,N_1570,N_1768);
and U2108 (N_2108,N_1863,N_1538);
nor U2109 (N_2109,N_1957,N_1818);
nand U2110 (N_2110,N_1665,N_1521);
or U2111 (N_2111,N_1746,N_1998);
nand U2112 (N_2112,N_1540,N_1541);
nor U2113 (N_2113,N_1707,N_1603);
nor U2114 (N_2114,N_1549,N_1529);
nand U2115 (N_2115,N_1904,N_1849);
nand U2116 (N_2116,N_1926,N_1615);
nand U2117 (N_2117,N_1941,N_1701);
nor U2118 (N_2118,N_1548,N_1937);
and U2119 (N_2119,N_1841,N_1825);
and U2120 (N_2120,N_1706,N_1591);
or U2121 (N_2121,N_1788,N_1583);
nand U2122 (N_2122,N_1695,N_1962);
xor U2123 (N_2123,N_1766,N_1735);
nand U2124 (N_2124,N_1712,N_1636);
and U2125 (N_2125,N_1565,N_1873);
nor U2126 (N_2126,N_1586,N_1934);
or U2127 (N_2127,N_1679,N_1682);
or U2128 (N_2128,N_1946,N_1893);
nor U2129 (N_2129,N_1931,N_1621);
nor U2130 (N_2130,N_1835,N_1974);
or U2131 (N_2131,N_1600,N_1764);
nor U2132 (N_2132,N_1504,N_1879);
nand U2133 (N_2133,N_1571,N_1744);
nand U2134 (N_2134,N_1854,N_1606);
and U2135 (N_2135,N_1643,N_1651);
nor U2136 (N_2136,N_1748,N_1660);
nand U2137 (N_2137,N_1720,N_1840);
nor U2138 (N_2138,N_1604,N_1902);
or U2139 (N_2139,N_1905,N_1500);
or U2140 (N_2140,N_1589,N_1683);
nor U2141 (N_2141,N_1767,N_1576);
and U2142 (N_2142,N_1616,N_1561);
nor U2143 (N_2143,N_1736,N_1558);
and U2144 (N_2144,N_1968,N_1810);
or U2145 (N_2145,N_1536,N_1629);
or U2146 (N_2146,N_1519,N_1650);
or U2147 (N_2147,N_1709,N_1692);
and U2148 (N_2148,N_1791,N_1508);
and U2149 (N_2149,N_1976,N_1876);
or U2150 (N_2150,N_1537,N_1526);
or U2151 (N_2151,N_1773,N_1585);
and U2152 (N_2152,N_1602,N_1842);
nor U2153 (N_2153,N_1938,N_1919);
or U2154 (N_2154,N_1542,N_1515);
nor U2155 (N_2155,N_1851,N_1824);
nand U2156 (N_2156,N_1803,N_1556);
nor U2157 (N_2157,N_1664,N_1644);
or U2158 (N_2158,N_1915,N_1716);
and U2159 (N_2159,N_1505,N_1573);
or U2160 (N_2160,N_1983,N_1759);
or U2161 (N_2161,N_1939,N_1594);
nand U2162 (N_2162,N_1783,N_1750);
and U2163 (N_2163,N_1816,N_1510);
nand U2164 (N_2164,N_1819,N_1917);
nand U2165 (N_2165,N_1761,N_1687);
nor U2166 (N_2166,N_1925,N_1717);
or U2167 (N_2167,N_1999,N_1648);
nand U2168 (N_2168,N_1550,N_1857);
xor U2169 (N_2169,N_1977,N_1846);
or U2170 (N_2170,N_1831,N_1814);
and U2171 (N_2171,N_1531,N_1792);
nor U2172 (N_2172,N_1563,N_1871);
and U2173 (N_2173,N_1733,N_1610);
and U2174 (N_2174,N_1832,N_1612);
and U2175 (N_2175,N_1710,N_1971);
or U2176 (N_2176,N_1821,N_1913);
and U2177 (N_2177,N_1725,N_1691);
nor U2178 (N_2178,N_1782,N_1997);
or U2179 (N_2179,N_1655,N_1993);
or U2180 (N_2180,N_1969,N_1673);
or U2181 (N_2181,N_1724,N_1844);
or U2182 (N_2182,N_1696,N_1663);
nand U2183 (N_2183,N_1763,N_1875);
or U2184 (N_2184,N_1624,N_1817);
and U2185 (N_2185,N_1547,N_1986);
or U2186 (N_2186,N_1661,N_1677);
and U2187 (N_2187,N_1959,N_1826);
and U2188 (N_2188,N_1513,N_1598);
or U2189 (N_2189,N_1545,N_1721);
or U2190 (N_2190,N_1956,N_1566);
and U2191 (N_2191,N_1595,N_1872);
nand U2192 (N_2192,N_1637,N_1704);
or U2193 (N_2193,N_1987,N_1756);
or U2194 (N_2194,N_1838,N_1568);
and U2195 (N_2195,N_1668,N_1823);
nand U2196 (N_2196,N_1726,N_1994);
nand U2197 (N_2197,N_1611,N_1684);
and U2198 (N_2198,N_1979,N_1535);
nand U2199 (N_2199,N_1685,N_1943);
nand U2200 (N_2200,N_1528,N_1512);
nor U2201 (N_2201,N_1885,N_1605);
and U2202 (N_2202,N_1740,N_1954);
nand U2203 (N_2203,N_1638,N_1789);
xor U2204 (N_2204,N_1947,N_1608);
nor U2205 (N_2205,N_1868,N_1811);
and U2206 (N_2206,N_1850,N_1845);
nand U2207 (N_2207,N_1964,N_1878);
or U2208 (N_2208,N_1760,N_1502);
and U2209 (N_2209,N_1864,N_1578);
nor U2210 (N_2210,N_1853,N_1901);
nand U2211 (N_2211,N_1777,N_1910);
nand U2212 (N_2212,N_1670,N_1903);
nor U2213 (N_2213,N_1795,N_1553);
or U2214 (N_2214,N_1575,N_1601);
nand U2215 (N_2215,N_1936,N_1848);
nor U2216 (N_2216,N_1708,N_1927);
nor U2217 (N_2217,N_1809,N_1562);
and U2218 (N_2218,N_1774,N_1867);
and U2219 (N_2219,N_1989,N_1580);
and U2220 (N_2220,N_1662,N_1640);
xnor U2221 (N_2221,N_1869,N_1715);
or U2222 (N_2222,N_1669,N_1524);
and U2223 (N_2223,N_1834,N_1633);
nand U2224 (N_2224,N_1555,N_1770);
nand U2225 (N_2225,N_1741,N_1516);
or U2226 (N_2226,N_1836,N_1827);
nand U2227 (N_2227,N_1780,N_1614);
nand U2228 (N_2228,N_1539,N_1932);
nor U2229 (N_2229,N_1883,N_1843);
or U2230 (N_2230,N_1728,N_1958);
nand U2231 (N_2231,N_1980,N_1551);
or U2232 (N_2232,N_1800,N_1785);
nand U2233 (N_2233,N_1847,N_1590);
and U2234 (N_2234,N_1745,N_1830);
and U2235 (N_2235,N_1753,N_1808);
nor U2236 (N_2236,N_1889,N_1861);
nand U2237 (N_2237,N_1641,N_1630);
nand U2238 (N_2238,N_1738,N_1940);
nand U2239 (N_2239,N_1860,N_1988);
and U2240 (N_2240,N_1786,N_1912);
or U2241 (N_2241,N_1908,N_1734);
nor U2242 (N_2242,N_1758,N_1697);
and U2243 (N_2243,N_1794,N_1609);
and U2244 (N_2244,N_1952,N_1532);
and U2245 (N_2245,N_1723,N_1642);
nand U2246 (N_2246,N_1804,N_1522);
nand U2247 (N_2247,N_1714,N_1574);
and U2248 (N_2248,N_1543,N_1982);
nand U2249 (N_2249,N_1837,N_1886);
and U2250 (N_2250,N_1754,N_1652);
and U2251 (N_2251,N_1653,N_1602);
nor U2252 (N_2252,N_1679,N_1840);
or U2253 (N_2253,N_1939,N_1758);
or U2254 (N_2254,N_1762,N_1974);
nor U2255 (N_2255,N_1520,N_1714);
xnor U2256 (N_2256,N_1856,N_1575);
nand U2257 (N_2257,N_1556,N_1964);
nor U2258 (N_2258,N_1593,N_1625);
nor U2259 (N_2259,N_1819,N_1663);
and U2260 (N_2260,N_1928,N_1743);
nand U2261 (N_2261,N_1516,N_1778);
and U2262 (N_2262,N_1826,N_1505);
nand U2263 (N_2263,N_1863,N_1825);
nor U2264 (N_2264,N_1693,N_1984);
nor U2265 (N_2265,N_1977,N_1720);
xor U2266 (N_2266,N_1954,N_1769);
nor U2267 (N_2267,N_1999,N_1730);
and U2268 (N_2268,N_1846,N_1587);
or U2269 (N_2269,N_1576,N_1746);
or U2270 (N_2270,N_1887,N_1636);
or U2271 (N_2271,N_1980,N_1509);
or U2272 (N_2272,N_1932,N_1627);
and U2273 (N_2273,N_1735,N_1665);
and U2274 (N_2274,N_1832,N_1911);
xor U2275 (N_2275,N_1998,N_1891);
nand U2276 (N_2276,N_1516,N_1521);
and U2277 (N_2277,N_1823,N_1551);
xor U2278 (N_2278,N_1801,N_1680);
nor U2279 (N_2279,N_1581,N_1812);
nand U2280 (N_2280,N_1503,N_1930);
nand U2281 (N_2281,N_1587,N_1836);
nand U2282 (N_2282,N_1927,N_1572);
and U2283 (N_2283,N_1826,N_1766);
and U2284 (N_2284,N_1574,N_1619);
nand U2285 (N_2285,N_1601,N_1547);
xor U2286 (N_2286,N_1926,N_1679);
and U2287 (N_2287,N_1979,N_1980);
and U2288 (N_2288,N_1801,N_1750);
nand U2289 (N_2289,N_1733,N_1543);
nand U2290 (N_2290,N_1825,N_1930);
or U2291 (N_2291,N_1857,N_1599);
nand U2292 (N_2292,N_1559,N_1817);
or U2293 (N_2293,N_1836,N_1535);
and U2294 (N_2294,N_1940,N_1874);
or U2295 (N_2295,N_1831,N_1987);
xnor U2296 (N_2296,N_1972,N_1895);
or U2297 (N_2297,N_1936,N_1811);
or U2298 (N_2298,N_1538,N_1577);
nand U2299 (N_2299,N_1907,N_1649);
or U2300 (N_2300,N_1970,N_1794);
nand U2301 (N_2301,N_1772,N_1895);
nor U2302 (N_2302,N_1684,N_1791);
nor U2303 (N_2303,N_1985,N_1917);
and U2304 (N_2304,N_1780,N_1611);
and U2305 (N_2305,N_1965,N_1611);
or U2306 (N_2306,N_1690,N_1550);
nor U2307 (N_2307,N_1581,N_1872);
and U2308 (N_2308,N_1753,N_1888);
nand U2309 (N_2309,N_1528,N_1930);
or U2310 (N_2310,N_1643,N_1883);
and U2311 (N_2311,N_1823,N_1971);
nor U2312 (N_2312,N_1553,N_1836);
nand U2313 (N_2313,N_1883,N_1546);
and U2314 (N_2314,N_1606,N_1866);
and U2315 (N_2315,N_1791,N_1863);
or U2316 (N_2316,N_1887,N_1501);
nor U2317 (N_2317,N_1938,N_1764);
or U2318 (N_2318,N_1847,N_1961);
and U2319 (N_2319,N_1834,N_1596);
nor U2320 (N_2320,N_1886,N_1835);
nor U2321 (N_2321,N_1727,N_1952);
or U2322 (N_2322,N_1534,N_1522);
or U2323 (N_2323,N_1947,N_1734);
nand U2324 (N_2324,N_1574,N_1697);
or U2325 (N_2325,N_1604,N_1534);
nand U2326 (N_2326,N_1791,N_1502);
and U2327 (N_2327,N_1928,N_1676);
or U2328 (N_2328,N_1583,N_1820);
and U2329 (N_2329,N_1518,N_1917);
or U2330 (N_2330,N_1862,N_1986);
and U2331 (N_2331,N_1892,N_1862);
or U2332 (N_2332,N_1683,N_1848);
nor U2333 (N_2333,N_1919,N_1762);
nor U2334 (N_2334,N_1588,N_1562);
or U2335 (N_2335,N_1803,N_1969);
or U2336 (N_2336,N_1811,N_1524);
and U2337 (N_2337,N_1582,N_1620);
nor U2338 (N_2338,N_1566,N_1729);
nor U2339 (N_2339,N_1799,N_1767);
nand U2340 (N_2340,N_1826,N_1702);
nor U2341 (N_2341,N_1813,N_1870);
and U2342 (N_2342,N_1774,N_1793);
nor U2343 (N_2343,N_1998,N_1541);
nor U2344 (N_2344,N_1831,N_1693);
nand U2345 (N_2345,N_1832,N_1942);
nand U2346 (N_2346,N_1805,N_1602);
and U2347 (N_2347,N_1854,N_1958);
nor U2348 (N_2348,N_1589,N_1823);
and U2349 (N_2349,N_1685,N_1736);
or U2350 (N_2350,N_1971,N_1708);
nor U2351 (N_2351,N_1517,N_1656);
xor U2352 (N_2352,N_1730,N_1942);
and U2353 (N_2353,N_1951,N_1547);
nand U2354 (N_2354,N_1896,N_1666);
nand U2355 (N_2355,N_1896,N_1744);
or U2356 (N_2356,N_1757,N_1750);
and U2357 (N_2357,N_1605,N_1511);
and U2358 (N_2358,N_1582,N_1740);
or U2359 (N_2359,N_1591,N_1522);
nand U2360 (N_2360,N_1510,N_1840);
nand U2361 (N_2361,N_1831,N_1916);
nand U2362 (N_2362,N_1635,N_1759);
nand U2363 (N_2363,N_1592,N_1512);
and U2364 (N_2364,N_1952,N_1814);
nand U2365 (N_2365,N_1698,N_1981);
and U2366 (N_2366,N_1938,N_1559);
xnor U2367 (N_2367,N_1628,N_1555);
or U2368 (N_2368,N_1958,N_1926);
nor U2369 (N_2369,N_1744,N_1722);
and U2370 (N_2370,N_1564,N_1571);
or U2371 (N_2371,N_1572,N_1618);
or U2372 (N_2372,N_1883,N_1687);
or U2373 (N_2373,N_1660,N_1645);
or U2374 (N_2374,N_1679,N_1542);
nor U2375 (N_2375,N_1939,N_1891);
and U2376 (N_2376,N_1551,N_1816);
nand U2377 (N_2377,N_1598,N_1850);
and U2378 (N_2378,N_1662,N_1516);
nor U2379 (N_2379,N_1889,N_1859);
nor U2380 (N_2380,N_1817,N_1979);
nand U2381 (N_2381,N_1878,N_1685);
and U2382 (N_2382,N_1635,N_1516);
nor U2383 (N_2383,N_1561,N_1908);
xor U2384 (N_2384,N_1503,N_1947);
or U2385 (N_2385,N_1621,N_1933);
nand U2386 (N_2386,N_1958,N_1898);
nor U2387 (N_2387,N_1628,N_1895);
or U2388 (N_2388,N_1562,N_1713);
and U2389 (N_2389,N_1651,N_1758);
and U2390 (N_2390,N_1517,N_1872);
nor U2391 (N_2391,N_1833,N_1960);
nor U2392 (N_2392,N_1788,N_1641);
nor U2393 (N_2393,N_1800,N_1877);
nand U2394 (N_2394,N_1777,N_1966);
or U2395 (N_2395,N_1528,N_1729);
nor U2396 (N_2396,N_1840,N_1929);
nor U2397 (N_2397,N_1642,N_1586);
or U2398 (N_2398,N_1607,N_1880);
nand U2399 (N_2399,N_1533,N_1553);
or U2400 (N_2400,N_1846,N_1569);
nor U2401 (N_2401,N_1976,N_1802);
or U2402 (N_2402,N_1764,N_1895);
nor U2403 (N_2403,N_1799,N_1632);
nor U2404 (N_2404,N_1641,N_1947);
nand U2405 (N_2405,N_1526,N_1897);
nor U2406 (N_2406,N_1877,N_1964);
and U2407 (N_2407,N_1969,N_1664);
and U2408 (N_2408,N_1581,N_1965);
nand U2409 (N_2409,N_1750,N_1528);
nand U2410 (N_2410,N_1914,N_1813);
or U2411 (N_2411,N_1872,N_1804);
or U2412 (N_2412,N_1919,N_1694);
nand U2413 (N_2413,N_1726,N_1944);
nand U2414 (N_2414,N_1605,N_1679);
nand U2415 (N_2415,N_1500,N_1545);
or U2416 (N_2416,N_1979,N_1614);
nand U2417 (N_2417,N_1674,N_1956);
nor U2418 (N_2418,N_1968,N_1975);
nor U2419 (N_2419,N_1907,N_1657);
nand U2420 (N_2420,N_1656,N_1583);
or U2421 (N_2421,N_1500,N_1737);
nor U2422 (N_2422,N_1737,N_1656);
or U2423 (N_2423,N_1956,N_1506);
or U2424 (N_2424,N_1732,N_1627);
nand U2425 (N_2425,N_1713,N_1742);
and U2426 (N_2426,N_1591,N_1857);
nor U2427 (N_2427,N_1572,N_1970);
and U2428 (N_2428,N_1942,N_1905);
and U2429 (N_2429,N_1686,N_1927);
and U2430 (N_2430,N_1619,N_1861);
nand U2431 (N_2431,N_1636,N_1607);
nor U2432 (N_2432,N_1860,N_1787);
nor U2433 (N_2433,N_1991,N_1900);
nor U2434 (N_2434,N_1985,N_1990);
or U2435 (N_2435,N_1713,N_1709);
nand U2436 (N_2436,N_1792,N_1575);
or U2437 (N_2437,N_1681,N_1763);
nor U2438 (N_2438,N_1656,N_1537);
nor U2439 (N_2439,N_1825,N_1651);
and U2440 (N_2440,N_1845,N_1669);
or U2441 (N_2441,N_1776,N_1918);
or U2442 (N_2442,N_1873,N_1693);
nor U2443 (N_2443,N_1795,N_1564);
xor U2444 (N_2444,N_1937,N_1524);
or U2445 (N_2445,N_1824,N_1713);
or U2446 (N_2446,N_1812,N_1915);
nor U2447 (N_2447,N_1952,N_1504);
nand U2448 (N_2448,N_1533,N_1704);
or U2449 (N_2449,N_1834,N_1546);
nor U2450 (N_2450,N_1684,N_1950);
nand U2451 (N_2451,N_1916,N_1917);
and U2452 (N_2452,N_1798,N_1958);
and U2453 (N_2453,N_1917,N_1562);
nand U2454 (N_2454,N_1711,N_1941);
nand U2455 (N_2455,N_1689,N_1934);
and U2456 (N_2456,N_1975,N_1999);
and U2457 (N_2457,N_1723,N_1902);
and U2458 (N_2458,N_1923,N_1940);
nor U2459 (N_2459,N_1858,N_1897);
nor U2460 (N_2460,N_1886,N_1860);
nor U2461 (N_2461,N_1813,N_1617);
nor U2462 (N_2462,N_1957,N_1515);
or U2463 (N_2463,N_1538,N_1647);
and U2464 (N_2464,N_1731,N_1912);
nor U2465 (N_2465,N_1588,N_1631);
or U2466 (N_2466,N_1687,N_1902);
nand U2467 (N_2467,N_1626,N_1543);
or U2468 (N_2468,N_1999,N_1601);
or U2469 (N_2469,N_1523,N_1786);
and U2470 (N_2470,N_1632,N_1993);
nand U2471 (N_2471,N_1884,N_1897);
or U2472 (N_2472,N_1989,N_1512);
or U2473 (N_2473,N_1686,N_1514);
nor U2474 (N_2474,N_1532,N_1954);
and U2475 (N_2475,N_1962,N_1679);
or U2476 (N_2476,N_1690,N_1661);
nand U2477 (N_2477,N_1749,N_1551);
nor U2478 (N_2478,N_1866,N_1980);
nand U2479 (N_2479,N_1538,N_1877);
nor U2480 (N_2480,N_1845,N_1897);
and U2481 (N_2481,N_1639,N_1823);
nand U2482 (N_2482,N_1526,N_1920);
and U2483 (N_2483,N_1621,N_1553);
nor U2484 (N_2484,N_1805,N_1936);
and U2485 (N_2485,N_1611,N_1920);
nand U2486 (N_2486,N_1536,N_1873);
nor U2487 (N_2487,N_1503,N_1749);
nand U2488 (N_2488,N_1505,N_1604);
nor U2489 (N_2489,N_1952,N_1588);
and U2490 (N_2490,N_1992,N_1514);
and U2491 (N_2491,N_1749,N_1573);
and U2492 (N_2492,N_1901,N_1757);
nand U2493 (N_2493,N_1932,N_1662);
nor U2494 (N_2494,N_1811,N_1921);
and U2495 (N_2495,N_1975,N_1972);
or U2496 (N_2496,N_1730,N_1719);
and U2497 (N_2497,N_1525,N_1529);
nand U2498 (N_2498,N_1788,N_1738);
and U2499 (N_2499,N_1981,N_1634);
nor U2500 (N_2500,N_2247,N_2434);
nor U2501 (N_2501,N_2143,N_2311);
or U2502 (N_2502,N_2221,N_2409);
xnor U2503 (N_2503,N_2249,N_2288);
nand U2504 (N_2504,N_2283,N_2363);
or U2505 (N_2505,N_2463,N_2100);
nand U2506 (N_2506,N_2203,N_2345);
nand U2507 (N_2507,N_2286,N_2038);
and U2508 (N_2508,N_2406,N_2414);
or U2509 (N_2509,N_2398,N_2494);
or U2510 (N_2510,N_2240,N_2072);
or U2511 (N_2511,N_2265,N_2448);
or U2512 (N_2512,N_2049,N_2482);
nand U2513 (N_2513,N_2098,N_2354);
and U2514 (N_2514,N_2151,N_2317);
or U2515 (N_2515,N_2300,N_2173);
and U2516 (N_2516,N_2115,N_2337);
and U2517 (N_2517,N_2374,N_2381);
nand U2518 (N_2518,N_2281,N_2070);
nand U2519 (N_2519,N_2295,N_2078);
xnor U2520 (N_2520,N_2382,N_2231);
xnor U2521 (N_2521,N_2040,N_2092);
or U2522 (N_2522,N_2274,N_2485);
or U2523 (N_2523,N_2178,N_2176);
nand U2524 (N_2524,N_2028,N_2370);
nand U2525 (N_2525,N_2459,N_2422);
nor U2526 (N_2526,N_2478,N_2280);
nand U2527 (N_2527,N_2105,N_2157);
nand U2528 (N_2528,N_2056,N_2114);
nand U2529 (N_2529,N_2277,N_2208);
nand U2530 (N_2530,N_2073,N_2312);
nor U2531 (N_2531,N_2356,N_2465);
nor U2532 (N_2532,N_2182,N_2322);
and U2533 (N_2533,N_2267,N_2076);
or U2534 (N_2534,N_2131,N_2170);
or U2535 (N_2535,N_2063,N_2079);
nand U2536 (N_2536,N_2423,N_2321);
or U2537 (N_2537,N_2084,N_2136);
nand U2538 (N_2538,N_2189,N_2426);
and U2539 (N_2539,N_2330,N_2493);
and U2540 (N_2540,N_2287,N_2006);
nor U2541 (N_2541,N_2097,N_2048);
or U2542 (N_2542,N_2066,N_2332);
nand U2543 (N_2543,N_2030,N_2424);
or U2544 (N_2544,N_2145,N_2418);
or U2545 (N_2545,N_2126,N_2452);
nand U2546 (N_2546,N_2230,N_2057);
or U2547 (N_2547,N_2026,N_2325);
or U2548 (N_2548,N_2326,N_2400);
nor U2549 (N_2549,N_2019,N_2349);
or U2550 (N_2550,N_2385,N_2160);
nor U2551 (N_2551,N_2331,N_2109);
nor U2552 (N_2552,N_2137,N_2053);
nor U2553 (N_2553,N_2141,N_2065);
nand U2554 (N_2554,N_2353,N_2154);
nor U2555 (N_2555,N_2215,N_2238);
nand U2556 (N_2556,N_2020,N_2236);
nor U2557 (N_2557,N_2188,N_2456);
nand U2558 (N_2558,N_2217,N_2243);
or U2559 (N_2559,N_2390,N_2439);
or U2560 (N_2560,N_2264,N_2237);
and U2561 (N_2561,N_2405,N_2183);
nand U2562 (N_2562,N_2486,N_2211);
and U2563 (N_2563,N_2016,N_2396);
nand U2564 (N_2564,N_2190,N_2491);
nand U2565 (N_2565,N_2259,N_2153);
nor U2566 (N_2566,N_2239,N_2191);
or U2567 (N_2567,N_2347,N_2244);
nand U2568 (N_2568,N_2474,N_2328);
and U2569 (N_2569,N_2383,N_2445);
or U2570 (N_2570,N_2293,N_2165);
nand U2571 (N_2571,N_2284,N_2175);
nand U2572 (N_2572,N_2446,N_2043);
nand U2573 (N_2573,N_2323,N_2166);
nor U2574 (N_2574,N_2488,N_2179);
and U2575 (N_2575,N_2319,N_2304);
and U2576 (N_2576,N_2301,N_2167);
nor U2577 (N_2577,N_2425,N_2025);
nand U2578 (N_2578,N_2181,N_2432);
nand U2579 (N_2579,N_2021,N_2172);
or U2580 (N_2580,N_2159,N_2348);
nand U2581 (N_2581,N_2343,N_2108);
and U2582 (N_2582,N_2089,N_2000);
nand U2583 (N_2583,N_2450,N_2135);
and U2584 (N_2584,N_2294,N_2483);
and U2585 (N_2585,N_2083,N_2462);
or U2586 (N_2586,N_2260,N_2158);
and U2587 (N_2587,N_2204,N_2226);
nand U2588 (N_2588,N_2024,N_2379);
and U2589 (N_2589,N_2013,N_2121);
nor U2590 (N_2590,N_2392,N_2269);
xnor U2591 (N_2591,N_2177,N_2142);
nand U2592 (N_2592,N_2421,N_2407);
and U2593 (N_2593,N_2275,N_2229);
or U2594 (N_2594,N_2014,N_2479);
or U2595 (N_2595,N_2134,N_2232);
nor U2596 (N_2596,N_2042,N_2252);
and U2597 (N_2597,N_2420,N_2324);
and U2598 (N_2598,N_2359,N_2338);
and U2599 (N_2599,N_2444,N_2192);
nand U2600 (N_2600,N_2438,N_2010);
or U2601 (N_2601,N_2431,N_2087);
xor U2602 (N_2602,N_2313,N_2186);
nand U2603 (N_2603,N_2373,N_2484);
nand U2604 (N_2604,N_2429,N_2086);
or U2605 (N_2605,N_2046,N_2194);
or U2606 (N_2606,N_2298,N_2080);
nor U2607 (N_2607,N_2387,N_2292);
nor U2608 (N_2608,N_2017,N_2029);
and U2609 (N_2609,N_2111,N_2256);
nand U2610 (N_2610,N_2402,N_2473);
nand U2611 (N_2611,N_2362,N_2116);
nor U2612 (N_2612,N_2336,N_2480);
nor U2613 (N_2613,N_2449,N_2271);
and U2614 (N_2614,N_2168,N_2454);
nor U2615 (N_2615,N_2442,N_2412);
nand U2616 (N_2616,N_2437,N_2075);
nor U2617 (N_2617,N_2316,N_2162);
nand U2618 (N_2618,N_2199,N_2443);
nand U2619 (N_2619,N_2380,N_2270);
xor U2620 (N_2620,N_2339,N_2144);
and U2621 (N_2621,N_2045,N_2498);
or U2622 (N_2622,N_2297,N_2218);
xnor U2623 (N_2623,N_2140,N_2302);
nor U2624 (N_2624,N_2015,N_2227);
nand U2625 (N_2625,N_2174,N_2403);
nor U2626 (N_2626,N_2050,N_2401);
or U2627 (N_2627,N_2471,N_2164);
nor U2628 (N_2628,N_2139,N_2487);
xnor U2629 (N_2629,N_2307,N_2453);
nand U2630 (N_2630,N_2455,N_2419);
and U2631 (N_2631,N_2253,N_2433);
or U2632 (N_2632,N_2251,N_2007);
nor U2633 (N_2633,N_2241,N_2315);
nand U2634 (N_2634,N_2246,N_2077);
or U2635 (N_2635,N_2150,N_2228);
nand U2636 (N_2636,N_2268,N_2299);
or U2637 (N_2637,N_2224,N_2254);
nor U2638 (N_2638,N_2138,N_2308);
or U2639 (N_2639,N_2093,N_2052);
or U2640 (N_2640,N_2161,N_2296);
or U2641 (N_2641,N_2250,N_2377);
nor U2642 (N_2642,N_2245,N_2205);
nand U2643 (N_2643,N_2171,N_2059);
and U2644 (N_2644,N_2071,N_2047);
or U2645 (N_2645,N_2068,N_2133);
nand U2646 (N_2646,N_2261,N_2395);
nor U2647 (N_2647,N_2002,N_2372);
and U2648 (N_2648,N_2394,N_2334);
nor U2649 (N_2649,N_2360,N_2263);
nor U2650 (N_2650,N_2351,N_2475);
nand U2651 (N_2651,N_2149,N_2120);
and U2652 (N_2652,N_2104,N_2369);
and U2653 (N_2653,N_2357,N_2096);
or U2654 (N_2654,N_2214,N_2318);
nand U2655 (N_2655,N_2102,N_2365);
or U2656 (N_2656,N_2074,N_2033);
nand U2657 (N_2657,N_2417,N_2430);
nor U2658 (N_2658,N_2408,N_2223);
nand U2659 (N_2659,N_2219,N_2124);
xnor U2660 (N_2660,N_2201,N_2200);
nor U2661 (N_2661,N_2082,N_2397);
nor U2662 (N_2662,N_2212,N_2005);
nor U2663 (N_2663,N_2107,N_2127);
nor U2664 (N_2664,N_2496,N_2340);
and U2665 (N_2665,N_2123,N_2054);
nand U2666 (N_2666,N_2185,N_2146);
or U2667 (N_2667,N_2361,N_2470);
or U2668 (N_2668,N_2037,N_2012);
nand U2669 (N_2669,N_2389,N_2064);
nand U2670 (N_2670,N_2272,N_2344);
nand U2671 (N_2671,N_2461,N_2004);
nand U2672 (N_2672,N_2291,N_2413);
nand U2673 (N_2673,N_2234,N_2466);
or U2674 (N_2674,N_2207,N_2011);
nor U2675 (N_2675,N_2163,N_2058);
and U2676 (N_2676,N_2416,N_2477);
or U2677 (N_2677,N_2341,N_2303);
or U2678 (N_2678,N_2187,N_2088);
nor U2679 (N_2679,N_2220,N_2489);
or U2680 (N_2680,N_2310,N_2113);
nand U2681 (N_2681,N_2495,N_2314);
nor U2682 (N_2682,N_2428,N_2282);
nor U2683 (N_2683,N_2335,N_2130);
nor U2684 (N_2684,N_2447,N_2305);
and U2685 (N_2685,N_2069,N_2391);
nor U2686 (N_2686,N_2320,N_2184);
or U2687 (N_2687,N_2032,N_2044);
or U2688 (N_2688,N_2285,N_2155);
nand U2689 (N_2689,N_2193,N_2350);
nor U2690 (N_2690,N_2112,N_2371);
nand U2691 (N_2691,N_2119,N_2036);
nand U2692 (N_2692,N_2148,N_2067);
and U2693 (N_2693,N_2061,N_2202);
nand U2694 (N_2694,N_2411,N_2085);
nor U2695 (N_2695,N_2290,N_2106);
and U2696 (N_2696,N_2327,N_2384);
nor U2697 (N_2697,N_2008,N_2090);
nor U2698 (N_2698,N_2279,N_2022);
and U2699 (N_2699,N_2342,N_2346);
nor U2700 (N_2700,N_2358,N_2376);
nand U2701 (N_2701,N_2352,N_2329);
nor U2702 (N_2702,N_2180,N_2467);
or U2703 (N_2703,N_2333,N_2415);
or U2704 (N_2704,N_2027,N_2242);
and U2705 (N_2705,N_2122,N_2198);
nor U2706 (N_2706,N_2469,N_2132);
or U2707 (N_2707,N_2041,N_2196);
nor U2708 (N_2708,N_2099,N_2197);
and U2709 (N_2709,N_2476,N_2472);
nand U2710 (N_2710,N_2481,N_2492);
and U2711 (N_2711,N_2147,N_2152);
or U2712 (N_2712,N_2094,N_2366);
and U2713 (N_2713,N_2169,N_2209);
or U2714 (N_2714,N_2278,N_2255);
nor U2715 (N_2715,N_2276,N_2435);
and U2716 (N_2716,N_2110,N_2410);
nor U2717 (N_2717,N_2399,N_2233);
or U2718 (N_2718,N_2035,N_2460);
and U2719 (N_2719,N_2095,N_2091);
nor U2720 (N_2720,N_2386,N_2009);
or U2721 (N_2721,N_2436,N_2388);
and U2722 (N_2722,N_2404,N_2195);
nand U2723 (N_2723,N_2129,N_2464);
or U2724 (N_2724,N_2118,N_2490);
nand U2725 (N_2725,N_2499,N_2216);
or U2726 (N_2726,N_2081,N_2213);
nand U2727 (N_2727,N_2128,N_2206);
and U2728 (N_2728,N_2309,N_2125);
or U2729 (N_2729,N_2210,N_2103);
and U2730 (N_2730,N_2451,N_2156);
and U2731 (N_2731,N_2355,N_2497);
nor U2732 (N_2732,N_2458,N_2468);
nand U2733 (N_2733,N_2051,N_2248);
and U2734 (N_2734,N_2235,N_2031);
and U2735 (N_2735,N_2101,N_2367);
and U2736 (N_2736,N_2060,N_2258);
or U2737 (N_2737,N_2001,N_2457);
nand U2738 (N_2738,N_2266,N_2225);
nor U2739 (N_2739,N_2062,N_2117);
xnor U2740 (N_2740,N_2440,N_2427);
and U2741 (N_2741,N_2018,N_2306);
and U2742 (N_2742,N_2222,N_2393);
nand U2743 (N_2743,N_2368,N_2441);
nor U2744 (N_2744,N_2378,N_2364);
and U2745 (N_2745,N_2375,N_2034);
nand U2746 (N_2746,N_2023,N_2055);
and U2747 (N_2747,N_2273,N_2257);
nand U2748 (N_2748,N_2039,N_2289);
or U2749 (N_2749,N_2262,N_2003);
or U2750 (N_2750,N_2225,N_2353);
nand U2751 (N_2751,N_2384,N_2025);
nor U2752 (N_2752,N_2064,N_2468);
nor U2753 (N_2753,N_2006,N_2463);
nor U2754 (N_2754,N_2167,N_2372);
xnor U2755 (N_2755,N_2091,N_2394);
nand U2756 (N_2756,N_2172,N_2241);
nand U2757 (N_2757,N_2069,N_2116);
nor U2758 (N_2758,N_2291,N_2231);
and U2759 (N_2759,N_2455,N_2161);
nand U2760 (N_2760,N_2284,N_2151);
nand U2761 (N_2761,N_2013,N_2032);
nor U2762 (N_2762,N_2420,N_2253);
and U2763 (N_2763,N_2064,N_2091);
or U2764 (N_2764,N_2107,N_2317);
nand U2765 (N_2765,N_2122,N_2311);
nor U2766 (N_2766,N_2006,N_2383);
xnor U2767 (N_2767,N_2193,N_2188);
nor U2768 (N_2768,N_2127,N_2158);
and U2769 (N_2769,N_2018,N_2327);
xnor U2770 (N_2770,N_2401,N_2164);
nand U2771 (N_2771,N_2102,N_2270);
nand U2772 (N_2772,N_2416,N_2128);
and U2773 (N_2773,N_2261,N_2181);
and U2774 (N_2774,N_2318,N_2405);
or U2775 (N_2775,N_2102,N_2362);
or U2776 (N_2776,N_2175,N_2211);
or U2777 (N_2777,N_2047,N_2086);
nor U2778 (N_2778,N_2411,N_2069);
or U2779 (N_2779,N_2383,N_2172);
nor U2780 (N_2780,N_2255,N_2094);
or U2781 (N_2781,N_2308,N_2153);
xnor U2782 (N_2782,N_2230,N_2408);
or U2783 (N_2783,N_2309,N_2040);
nand U2784 (N_2784,N_2074,N_2112);
nand U2785 (N_2785,N_2385,N_2440);
nor U2786 (N_2786,N_2008,N_2119);
nand U2787 (N_2787,N_2387,N_2004);
or U2788 (N_2788,N_2021,N_2216);
or U2789 (N_2789,N_2095,N_2016);
nor U2790 (N_2790,N_2398,N_2173);
and U2791 (N_2791,N_2378,N_2045);
nor U2792 (N_2792,N_2068,N_2106);
and U2793 (N_2793,N_2462,N_2072);
and U2794 (N_2794,N_2174,N_2486);
or U2795 (N_2795,N_2152,N_2216);
nor U2796 (N_2796,N_2246,N_2049);
and U2797 (N_2797,N_2488,N_2168);
or U2798 (N_2798,N_2244,N_2093);
and U2799 (N_2799,N_2351,N_2303);
nand U2800 (N_2800,N_2003,N_2230);
and U2801 (N_2801,N_2321,N_2204);
or U2802 (N_2802,N_2498,N_2359);
or U2803 (N_2803,N_2364,N_2327);
nand U2804 (N_2804,N_2397,N_2335);
nand U2805 (N_2805,N_2228,N_2465);
nor U2806 (N_2806,N_2155,N_2016);
nand U2807 (N_2807,N_2423,N_2204);
nor U2808 (N_2808,N_2379,N_2214);
and U2809 (N_2809,N_2104,N_2215);
nand U2810 (N_2810,N_2258,N_2148);
nor U2811 (N_2811,N_2132,N_2276);
or U2812 (N_2812,N_2252,N_2263);
or U2813 (N_2813,N_2087,N_2277);
and U2814 (N_2814,N_2332,N_2141);
and U2815 (N_2815,N_2300,N_2482);
and U2816 (N_2816,N_2179,N_2372);
nor U2817 (N_2817,N_2055,N_2211);
or U2818 (N_2818,N_2256,N_2457);
nand U2819 (N_2819,N_2243,N_2442);
and U2820 (N_2820,N_2494,N_2475);
or U2821 (N_2821,N_2452,N_2420);
nand U2822 (N_2822,N_2133,N_2130);
or U2823 (N_2823,N_2132,N_2138);
nand U2824 (N_2824,N_2292,N_2248);
and U2825 (N_2825,N_2076,N_2144);
or U2826 (N_2826,N_2330,N_2125);
and U2827 (N_2827,N_2066,N_2353);
and U2828 (N_2828,N_2457,N_2072);
nor U2829 (N_2829,N_2273,N_2066);
nand U2830 (N_2830,N_2199,N_2491);
nor U2831 (N_2831,N_2384,N_2448);
and U2832 (N_2832,N_2499,N_2062);
and U2833 (N_2833,N_2274,N_2061);
nor U2834 (N_2834,N_2073,N_2430);
nand U2835 (N_2835,N_2432,N_2273);
nand U2836 (N_2836,N_2206,N_2127);
nor U2837 (N_2837,N_2412,N_2257);
nand U2838 (N_2838,N_2473,N_2481);
nand U2839 (N_2839,N_2015,N_2039);
and U2840 (N_2840,N_2150,N_2105);
nand U2841 (N_2841,N_2316,N_2301);
and U2842 (N_2842,N_2289,N_2056);
nand U2843 (N_2843,N_2037,N_2050);
or U2844 (N_2844,N_2432,N_2474);
xnor U2845 (N_2845,N_2390,N_2337);
and U2846 (N_2846,N_2459,N_2086);
or U2847 (N_2847,N_2459,N_2278);
nand U2848 (N_2848,N_2101,N_2335);
nand U2849 (N_2849,N_2331,N_2215);
nand U2850 (N_2850,N_2216,N_2250);
nor U2851 (N_2851,N_2377,N_2046);
nand U2852 (N_2852,N_2087,N_2272);
nor U2853 (N_2853,N_2182,N_2269);
and U2854 (N_2854,N_2300,N_2148);
nand U2855 (N_2855,N_2483,N_2176);
or U2856 (N_2856,N_2353,N_2365);
or U2857 (N_2857,N_2306,N_2337);
nor U2858 (N_2858,N_2016,N_2405);
and U2859 (N_2859,N_2480,N_2073);
nand U2860 (N_2860,N_2430,N_2159);
or U2861 (N_2861,N_2156,N_2173);
nor U2862 (N_2862,N_2394,N_2454);
and U2863 (N_2863,N_2330,N_2333);
and U2864 (N_2864,N_2349,N_2475);
nand U2865 (N_2865,N_2140,N_2454);
and U2866 (N_2866,N_2334,N_2321);
nand U2867 (N_2867,N_2100,N_2434);
and U2868 (N_2868,N_2496,N_2326);
nand U2869 (N_2869,N_2071,N_2073);
nand U2870 (N_2870,N_2222,N_2187);
xnor U2871 (N_2871,N_2021,N_2255);
nand U2872 (N_2872,N_2347,N_2318);
nand U2873 (N_2873,N_2278,N_2238);
nor U2874 (N_2874,N_2460,N_2195);
and U2875 (N_2875,N_2463,N_2153);
nor U2876 (N_2876,N_2233,N_2282);
or U2877 (N_2877,N_2052,N_2335);
nor U2878 (N_2878,N_2206,N_2298);
and U2879 (N_2879,N_2057,N_2060);
and U2880 (N_2880,N_2378,N_2125);
nand U2881 (N_2881,N_2066,N_2390);
nor U2882 (N_2882,N_2016,N_2413);
nor U2883 (N_2883,N_2475,N_2355);
nand U2884 (N_2884,N_2324,N_2244);
nand U2885 (N_2885,N_2469,N_2414);
and U2886 (N_2886,N_2250,N_2110);
nor U2887 (N_2887,N_2124,N_2016);
and U2888 (N_2888,N_2095,N_2015);
or U2889 (N_2889,N_2034,N_2109);
or U2890 (N_2890,N_2404,N_2005);
nor U2891 (N_2891,N_2098,N_2464);
or U2892 (N_2892,N_2251,N_2392);
or U2893 (N_2893,N_2487,N_2422);
or U2894 (N_2894,N_2061,N_2480);
nand U2895 (N_2895,N_2226,N_2249);
nor U2896 (N_2896,N_2426,N_2213);
or U2897 (N_2897,N_2082,N_2210);
and U2898 (N_2898,N_2085,N_2432);
nand U2899 (N_2899,N_2380,N_2070);
xor U2900 (N_2900,N_2165,N_2456);
nor U2901 (N_2901,N_2262,N_2408);
and U2902 (N_2902,N_2402,N_2145);
nor U2903 (N_2903,N_2009,N_2229);
xor U2904 (N_2904,N_2196,N_2183);
and U2905 (N_2905,N_2106,N_2496);
nand U2906 (N_2906,N_2253,N_2062);
nor U2907 (N_2907,N_2030,N_2496);
nor U2908 (N_2908,N_2371,N_2437);
and U2909 (N_2909,N_2115,N_2027);
and U2910 (N_2910,N_2350,N_2458);
nand U2911 (N_2911,N_2372,N_2024);
nand U2912 (N_2912,N_2394,N_2376);
nand U2913 (N_2913,N_2379,N_2469);
and U2914 (N_2914,N_2081,N_2017);
or U2915 (N_2915,N_2043,N_2297);
and U2916 (N_2916,N_2330,N_2439);
and U2917 (N_2917,N_2123,N_2301);
and U2918 (N_2918,N_2005,N_2016);
and U2919 (N_2919,N_2280,N_2467);
nand U2920 (N_2920,N_2102,N_2241);
nor U2921 (N_2921,N_2046,N_2188);
nor U2922 (N_2922,N_2465,N_2136);
or U2923 (N_2923,N_2035,N_2448);
nand U2924 (N_2924,N_2075,N_2104);
or U2925 (N_2925,N_2204,N_2465);
and U2926 (N_2926,N_2378,N_2341);
nor U2927 (N_2927,N_2094,N_2463);
or U2928 (N_2928,N_2020,N_2287);
or U2929 (N_2929,N_2410,N_2136);
nand U2930 (N_2930,N_2112,N_2148);
nand U2931 (N_2931,N_2407,N_2338);
nand U2932 (N_2932,N_2246,N_2382);
or U2933 (N_2933,N_2425,N_2470);
and U2934 (N_2934,N_2091,N_2219);
nor U2935 (N_2935,N_2122,N_2321);
nand U2936 (N_2936,N_2198,N_2188);
nand U2937 (N_2937,N_2358,N_2042);
or U2938 (N_2938,N_2139,N_2071);
nand U2939 (N_2939,N_2024,N_2015);
or U2940 (N_2940,N_2311,N_2155);
nor U2941 (N_2941,N_2006,N_2357);
nor U2942 (N_2942,N_2294,N_2097);
or U2943 (N_2943,N_2380,N_2271);
and U2944 (N_2944,N_2225,N_2006);
or U2945 (N_2945,N_2084,N_2017);
nand U2946 (N_2946,N_2300,N_2033);
or U2947 (N_2947,N_2025,N_2475);
or U2948 (N_2948,N_2441,N_2304);
nor U2949 (N_2949,N_2187,N_2387);
nand U2950 (N_2950,N_2312,N_2350);
nand U2951 (N_2951,N_2434,N_2494);
or U2952 (N_2952,N_2481,N_2465);
nand U2953 (N_2953,N_2209,N_2086);
nor U2954 (N_2954,N_2112,N_2230);
or U2955 (N_2955,N_2474,N_2184);
nand U2956 (N_2956,N_2037,N_2194);
and U2957 (N_2957,N_2431,N_2239);
nand U2958 (N_2958,N_2377,N_2197);
or U2959 (N_2959,N_2355,N_2428);
or U2960 (N_2960,N_2456,N_2284);
nor U2961 (N_2961,N_2363,N_2154);
nand U2962 (N_2962,N_2092,N_2407);
nor U2963 (N_2963,N_2491,N_2193);
and U2964 (N_2964,N_2428,N_2017);
nor U2965 (N_2965,N_2106,N_2449);
or U2966 (N_2966,N_2007,N_2250);
nor U2967 (N_2967,N_2014,N_2373);
nand U2968 (N_2968,N_2433,N_2108);
and U2969 (N_2969,N_2153,N_2395);
and U2970 (N_2970,N_2460,N_2186);
xor U2971 (N_2971,N_2360,N_2050);
and U2972 (N_2972,N_2405,N_2419);
or U2973 (N_2973,N_2029,N_2339);
and U2974 (N_2974,N_2340,N_2092);
and U2975 (N_2975,N_2382,N_2308);
nor U2976 (N_2976,N_2077,N_2189);
or U2977 (N_2977,N_2033,N_2150);
and U2978 (N_2978,N_2153,N_2392);
nor U2979 (N_2979,N_2481,N_2360);
nor U2980 (N_2980,N_2246,N_2342);
or U2981 (N_2981,N_2115,N_2192);
and U2982 (N_2982,N_2061,N_2227);
or U2983 (N_2983,N_2179,N_2023);
nor U2984 (N_2984,N_2136,N_2355);
nor U2985 (N_2985,N_2277,N_2267);
nand U2986 (N_2986,N_2348,N_2404);
nor U2987 (N_2987,N_2072,N_2121);
nor U2988 (N_2988,N_2461,N_2256);
or U2989 (N_2989,N_2314,N_2254);
or U2990 (N_2990,N_2179,N_2030);
and U2991 (N_2991,N_2064,N_2283);
and U2992 (N_2992,N_2056,N_2396);
xnor U2993 (N_2993,N_2020,N_2072);
or U2994 (N_2994,N_2476,N_2314);
or U2995 (N_2995,N_2074,N_2030);
nor U2996 (N_2996,N_2199,N_2251);
or U2997 (N_2997,N_2099,N_2323);
nor U2998 (N_2998,N_2338,N_2045);
or U2999 (N_2999,N_2353,N_2044);
and UO_0 (O_0,N_2918,N_2809);
nand UO_1 (O_1,N_2648,N_2552);
and UO_2 (O_2,N_2910,N_2720);
nand UO_3 (O_3,N_2862,N_2959);
nand UO_4 (O_4,N_2734,N_2963);
nor UO_5 (O_5,N_2729,N_2771);
nand UO_6 (O_6,N_2527,N_2711);
nand UO_7 (O_7,N_2577,N_2861);
and UO_8 (O_8,N_2931,N_2977);
nor UO_9 (O_9,N_2642,N_2851);
and UO_10 (O_10,N_2717,N_2830);
xnor UO_11 (O_11,N_2796,N_2713);
and UO_12 (O_12,N_2900,N_2687);
and UO_13 (O_13,N_2906,N_2555);
and UO_14 (O_14,N_2578,N_2927);
or UO_15 (O_15,N_2509,N_2859);
nor UO_16 (O_16,N_2890,N_2650);
or UO_17 (O_17,N_2854,N_2674);
and UO_18 (O_18,N_2882,N_2945);
nand UO_19 (O_19,N_2602,N_2984);
nand UO_20 (O_20,N_2723,N_2722);
nor UO_21 (O_21,N_2614,N_2735);
nand UO_22 (O_22,N_2948,N_2957);
nor UO_23 (O_23,N_2574,N_2630);
nand UO_24 (O_24,N_2542,N_2865);
nor UO_25 (O_25,N_2995,N_2785);
or UO_26 (O_26,N_2903,N_2522);
nor UO_27 (O_27,N_2606,N_2715);
nand UO_28 (O_28,N_2770,N_2651);
nor UO_29 (O_29,N_2874,N_2609);
and UO_30 (O_30,N_2905,N_2673);
or UO_31 (O_31,N_2936,N_2751);
nand UO_32 (O_32,N_2581,N_2850);
nor UO_33 (O_33,N_2632,N_2562);
or UO_34 (O_34,N_2605,N_2848);
or UO_35 (O_35,N_2636,N_2820);
nor UO_36 (O_36,N_2528,N_2914);
or UO_37 (O_37,N_2965,N_2662);
nor UO_38 (O_38,N_2669,N_2691);
or UO_39 (O_39,N_2658,N_2849);
nand UO_40 (O_40,N_2897,N_2730);
nand UO_41 (O_41,N_2898,N_2917);
or UO_42 (O_42,N_2976,N_2604);
nand UO_43 (O_43,N_2797,N_2500);
nand UO_44 (O_44,N_2647,N_2638);
xor UO_45 (O_45,N_2737,N_2908);
nor UO_46 (O_46,N_2919,N_2736);
nand UO_47 (O_47,N_2641,N_2838);
nand UO_48 (O_48,N_2834,N_2664);
or UO_49 (O_49,N_2686,N_2879);
nor UO_50 (O_50,N_2923,N_2946);
nor UO_51 (O_51,N_2829,N_2966);
or UO_52 (O_52,N_2612,N_2894);
nor UO_53 (O_53,N_2951,N_2800);
or UO_54 (O_54,N_2986,N_2937);
and UO_55 (O_55,N_2991,N_2708);
nor UO_56 (O_56,N_2576,N_2526);
nand UO_57 (O_57,N_2666,N_2875);
nand UO_58 (O_58,N_2613,N_2765);
and UO_59 (O_59,N_2911,N_2626);
nand UO_60 (O_60,N_2808,N_2792);
and UO_61 (O_61,N_2907,N_2913);
nand UO_62 (O_62,N_2858,N_2889);
nor UO_63 (O_63,N_2592,N_2749);
nand UO_64 (O_64,N_2588,N_2795);
nand UO_65 (O_65,N_2503,N_2690);
nor UO_66 (O_66,N_2826,N_2880);
and UO_67 (O_67,N_2961,N_2646);
and UO_68 (O_68,N_2721,N_2960);
and UO_69 (O_69,N_2779,N_2783);
nor UO_70 (O_70,N_2998,N_2703);
nor UO_71 (O_71,N_2530,N_2643);
nand UO_72 (O_72,N_2853,N_2816);
or UO_73 (O_73,N_2827,N_2844);
or UO_74 (O_74,N_2752,N_2583);
nor UO_75 (O_75,N_2627,N_2534);
and UO_76 (O_76,N_2872,N_2563);
nand UO_77 (O_77,N_2596,N_2760);
nand UO_78 (O_78,N_2617,N_2618);
or UO_79 (O_79,N_2981,N_2584);
nor UO_80 (O_80,N_2996,N_2988);
nor UO_81 (O_81,N_2585,N_2504);
nor UO_82 (O_82,N_2663,N_2661);
nor UO_83 (O_83,N_2944,N_2971);
and UO_84 (O_84,N_2788,N_2611);
and UO_85 (O_85,N_2693,N_2989);
nand UO_86 (O_86,N_2529,N_2942);
or UO_87 (O_87,N_2835,N_2575);
or UO_88 (O_88,N_2634,N_2649);
nand UO_89 (O_89,N_2515,N_2746);
nor UO_90 (O_90,N_2544,N_2825);
and UO_91 (O_91,N_2782,N_2706);
or UO_92 (O_92,N_2569,N_2828);
or UO_93 (O_93,N_2599,N_2570);
and UO_94 (O_94,N_2993,N_2671);
nor UO_95 (O_95,N_2840,N_2731);
nor UO_96 (O_96,N_2922,N_2573);
nor UO_97 (O_97,N_2631,N_2695);
nor UO_98 (O_98,N_2501,N_2619);
nand UO_99 (O_99,N_2512,N_2582);
or UO_100 (O_100,N_2644,N_2565);
nand UO_101 (O_101,N_2941,N_2842);
or UO_102 (O_102,N_2759,N_2856);
nand UO_103 (O_103,N_2939,N_2766);
nand UO_104 (O_104,N_2860,N_2777);
nor UO_105 (O_105,N_2550,N_2811);
nor UO_106 (O_106,N_2639,N_2933);
nand UO_107 (O_107,N_2714,N_2786);
nand UO_108 (O_108,N_2652,N_2755);
nor UO_109 (O_109,N_2557,N_2928);
xor UO_110 (O_110,N_2883,N_2677);
or UO_111 (O_111,N_2560,N_2566);
or UO_112 (O_112,N_2982,N_2778);
nand UO_113 (O_113,N_2878,N_2776);
or UO_114 (O_114,N_2997,N_2622);
nand UO_115 (O_115,N_2969,N_2852);
or UO_116 (O_116,N_2832,N_2629);
and UO_117 (O_117,N_2887,N_2615);
nor UO_118 (O_118,N_2885,N_2533);
or UO_119 (O_119,N_2517,N_2537);
or UO_120 (O_120,N_2764,N_2794);
nand UO_121 (O_121,N_2726,N_2524);
nor UO_122 (O_122,N_2683,N_2932);
nor UO_123 (O_123,N_2817,N_2571);
nor UO_124 (O_124,N_2962,N_2950);
or UO_125 (O_125,N_2806,N_2655);
nor UO_126 (O_126,N_2593,N_2864);
or UO_127 (O_127,N_2667,N_2915);
nand UO_128 (O_128,N_2938,N_2926);
nand UO_129 (O_129,N_2798,N_2824);
nor UO_130 (O_130,N_2821,N_2724);
or UO_131 (O_131,N_2679,N_2974);
and UO_132 (O_132,N_2620,N_2819);
nor UO_133 (O_133,N_2520,N_2769);
nor UO_134 (O_134,N_2597,N_2934);
nand UO_135 (O_135,N_2698,N_2902);
nand UO_136 (O_136,N_2833,N_2702);
or UO_137 (O_137,N_2710,N_2733);
xor UO_138 (O_138,N_2892,N_2507);
nand UO_139 (O_139,N_2704,N_2884);
nand UO_140 (O_140,N_2712,N_2675);
and UO_141 (O_141,N_2756,N_2940);
nand UO_142 (O_142,N_2672,N_2625);
or UO_143 (O_143,N_2623,N_2633);
and UO_144 (O_144,N_2754,N_2580);
and UO_145 (O_145,N_2904,N_2546);
nor UO_146 (O_146,N_2701,N_2719);
nand UO_147 (O_147,N_2539,N_2958);
or UO_148 (O_148,N_2610,N_2518);
nand UO_149 (O_149,N_2505,N_2689);
nand UO_150 (O_150,N_2822,N_2983);
nor UO_151 (O_151,N_2670,N_2513);
nand UO_152 (O_152,N_2725,N_2804);
or UO_153 (O_153,N_2543,N_2899);
or UO_154 (O_154,N_2579,N_2743);
nor UO_155 (O_155,N_2799,N_2877);
or UO_156 (O_156,N_2678,N_2600);
or UO_157 (O_157,N_2548,N_2637);
xnor UO_158 (O_158,N_2739,N_2716);
and UO_159 (O_159,N_2978,N_2598);
or UO_160 (O_160,N_2616,N_2553);
and UO_161 (O_161,N_2823,N_2556);
and UO_162 (O_162,N_2909,N_2510);
and UO_163 (O_163,N_2980,N_2893);
and UO_164 (O_164,N_2949,N_2668);
and UO_165 (O_165,N_2564,N_2659);
and UO_166 (O_166,N_2881,N_2531);
and UO_167 (O_167,N_2682,N_2709);
nor UO_168 (O_168,N_2810,N_2845);
and UO_169 (O_169,N_2802,N_2793);
and UO_170 (O_170,N_2591,N_2818);
or UO_171 (O_171,N_2586,N_2547);
nand UO_172 (O_172,N_2930,N_2921);
and UO_173 (O_173,N_2740,N_2727);
nand UO_174 (O_174,N_2867,N_2741);
nand UO_175 (O_175,N_2841,N_2645);
nor UO_176 (O_176,N_2511,N_2803);
nand UO_177 (O_177,N_2567,N_2912);
or UO_178 (O_178,N_2773,N_2814);
nand UO_179 (O_179,N_2685,N_2654);
and UO_180 (O_180,N_2775,N_2888);
nor UO_181 (O_181,N_2813,N_2891);
xnor UO_182 (O_182,N_2943,N_2869);
or UO_183 (O_183,N_2707,N_2601);
nor UO_184 (O_184,N_2545,N_2536);
nor UO_185 (O_185,N_2784,N_2870);
or UO_186 (O_186,N_2753,N_2990);
nor UO_187 (O_187,N_2805,N_2595);
and UO_188 (O_188,N_2863,N_2692);
nor UO_189 (O_189,N_2621,N_2705);
nor UO_190 (O_190,N_2718,N_2968);
or UO_191 (O_191,N_2947,N_2508);
nand UO_192 (O_192,N_2970,N_2697);
nor UO_193 (O_193,N_2767,N_2954);
or UO_194 (O_194,N_2680,N_2768);
and UO_195 (O_195,N_2681,N_2763);
nor UO_196 (O_196,N_2525,N_2837);
nand UO_197 (O_197,N_2973,N_2558);
nor UO_198 (O_198,N_2761,N_2608);
and UO_199 (O_199,N_2757,N_2738);
xor UO_200 (O_200,N_2516,N_2895);
and UO_201 (O_201,N_2985,N_2815);
and UO_202 (O_202,N_2807,N_2559);
or UO_203 (O_203,N_2521,N_2523);
or UO_204 (O_204,N_2538,N_2924);
or UO_205 (O_205,N_2975,N_2772);
or UO_206 (O_206,N_2876,N_2532);
or UO_207 (O_207,N_2953,N_2831);
nand UO_208 (O_208,N_2994,N_2628);
nand UO_209 (O_209,N_2790,N_2781);
nand UO_210 (O_210,N_2561,N_2535);
or UO_211 (O_211,N_2607,N_2624);
nor UO_212 (O_212,N_2886,N_2925);
nand UO_213 (O_213,N_2871,N_2846);
or UO_214 (O_214,N_2987,N_2929);
xor UO_215 (O_215,N_2656,N_2748);
nor UO_216 (O_216,N_2541,N_2660);
and UO_217 (O_217,N_2956,N_2873);
and UO_218 (O_218,N_2747,N_2857);
and UO_219 (O_219,N_2688,N_2999);
nor UO_220 (O_220,N_2676,N_2896);
nor UO_221 (O_221,N_2554,N_2801);
nor UO_222 (O_222,N_2916,N_2836);
or UO_223 (O_223,N_2540,N_2868);
nor UO_224 (O_224,N_2972,N_2568);
and UO_225 (O_225,N_2935,N_2750);
and UO_226 (O_226,N_2847,N_2549);
or UO_227 (O_227,N_2514,N_2732);
or UO_228 (O_228,N_2744,N_2594);
nand UO_229 (O_229,N_2762,N_2955);
xnor UO_230 (O_230,N_2728,N_2901);
or UO_231 (O_231,N_2640,N_2787);
nand UO_232 (O_232,N_2696,N_2791);
nor UO_233 (O_233,N_2694,N_2590);
nor UO_234 (O_234,N_2587,N_2812);
nand UO_235 (O_235,N_2855,N_2758);
and UO_236 (O_236,N_2635,N_2789);
and UO_237 (O_237,N_2742,N_2774);
or UO_238 (O_238,N_2992,N_2551);
or UO_239 (O_239,N_2967,N_2657);
or UO_240 (O_240,N_2699,N_2589);
nor UO_241 (O_241,N_2866,N_2780);
or UO_242 (O_242,N_2653,N_2979);
nand UO_243 (O_243,N_2920,N_2964);
nand UO_244 (O_244,N_2839,N_2745);
or UO_245 (O_245,N_2502,N_2519);
and UO_246 (O_246,N_2700,N_2665);
and UO_247 (O_247,N_2506,N_2684);
and UO_248 (O_248,N_2952,N_2572);
or UO_249 (O_249,N_2843,N_2603);
or UO_250 (O_250,N_2540,N_2818);
nand UO_251 (O_251,N_2767,N_2962);
nand UO_252 (O_252,N_2714,N_2879);
nor UO_253 (O_253,N_2652,N_2891);
and UO_254 (O_254,N_2853,N_2963);
nand UO_255 (O_255,N_2948,N_2910);
and UO_256 (O_256,N_2802,N_2507);
or UO_257 (O_257,N_2973,N_2599);
nor UO_258 (O_258,N_2619,N_2595);
or UO_259 (O_259,N_2880,N_2689);
and UO_260 (O_260,N_2845,N_2986);
or UO_261 (O_261,N_2925,N_2721);
nor UO_262 (O_262,N_2577,N_2827);
and UO_263 (O_263,N_2915,N_2938);
nand UO_264 (O_264,N_2700,N_2654);
and UO_265 (O_265,N_2617,N_2980);
nor UO_266 (O_266,N_2547,N_2572);
and UO_267 (O_267,N_2552,N_2851);
or UO_268 (O_268,N_2590,N_2837);
or UO_269 (O_269,N_2545,N_2636);
and UO_270 (O_270,N_2801,N_2948);
or UO_271 (O_271,N_2924,N_2633);
nor UO_272 (O_272,N_2966,N_2587);
nand UO_273 (O_273,N_2824,N_2994);
nand UO_274 (O_274,N_2720,N_2707);
or UO_275 (O_275,N_2768,N_2734);
nand UO_276 (O_276,N_2934,N_2822);
nor UO_277 (O_277,N_2608,N_2751);
or UO_278 (O_278,N_2693,N_2881);
or UO_279 (O_279,N_2879,N_2683);
nand UO_280 (O_280,N_2817,N_2724);
nor UO_281 (O_281,N_2599,N_2500);
xnor UO_282 (O_282,N_2801,N_2518);
xor UO_283 (O_283,N_2581,N_2584);
and UO_284 (O_284,N_2699,N_2636);
nor UO_285 (O_285,N_2584,N_2608);
and UO_286 (O_286,N_2705,N_2779);
xnor UO_287 (O_287,N_2803,N_2967);
or UO_288 (O_288,N_2540,N_2808);
nor UO_289 (O_289,N_2702,N_2540);
or UO_290 (O_290,N_2507,N_2528);
nor UO_291 (O_291,N_2783,N_2607);
nor UO_292 (O_292,N_2555,N_2748);
nor UO_293 (O_293,N_2607,N_2834);
and UO_294 (O_294,N_2533,N_2561);
or UO_295 (O_295,N_2689,N_2621);
and UO_296 (O_296,N_2907,N_2974);
or UO_297 (O_297,N_2704,N_2615);
or UO_298 (O_298,N_2528,N_2923);
or UO_299 (O_299,N_2819,N_2884);
nand UO_300 (O_300,N_2774,N_2898);
nor UO_301 (O_301,N_2634,N_2618);
nor UO_302 (O_302,N_2761,N_2941);
or UO_303 (O_303,N_2667,N_2945);
nor UO_304 (O_304,N_2629,N_2747);
nor UO_305 (O_305,N_2529,N_2855);
or UO_306 (O_306,N_2643,N_2593);
nor UO_307 (O_307,N_2645,N_2759);
nand UO_308 (O_308,N_2894,N_2750);
or UO_309 (O_309,N_2625,N_2810);
nand UO_310 (O_310,N_2507,N_2858);
or UO_311 (O_311,N_2636,N_2646);
nor UO_312 (O_312,N_2813,N_2597);
nand UO_313 (O_313,N_2890,N_2783);
and UO_314 (O_314,N_2706,N_2591);
nand UO_315 (O_315,N_2816,N_2821);
and UO_316 (O_316,N_2739,N_2650);
or UO_317 (O_317,N_2822,N_2538);
or UO_318 (O_318,N_2565,N_2824);
or UO_319 (O_319,N_2542,N_2796);
or UO_320 (O_320,N_2540,N_2699);
nor UO_321 (O_321,N_2592,N_2570);
or UO_322 (O_322,N_2786,N_2885);
or UO_323 (O_323,N_2500,N_2941);
nand UO_324 (O_324,N_2771,N_2613);
nor UO_325 (O_325,N_2828,N_2560);
nor UO_326 (O_326,N_2692,N_2691);
xnor UO_327 (O_327,N_2651,N_2743);
nand UO_328 (O_328,N_2550,N_2936);
and UO_329 (O_329,N_2912,N_2901);
nor UO_330 (O_330,N_2522,N_2705);
nor UO_331 (O_331,N_2952,N_2725);
nand UO_332 (O_332,N_2843,N_2556);
or UO_333 (O_333,N_2755,N_2911);
or UO_334 (O_334,N_2582,N_2605);
or UO_335 (O_335,N_2876,N_2704);
and UO_336 (O_336,N_2616,N_2754);
and UO_337 (O_337,N_2922,N_2923);
or UO_338 (O_338,N_2595,N_2743);
nor UO_339 (O_339,N_2951,N_2719);
nand UO_340 (O_340,N_2907,N_2981);
nand UO_341 (O_341,N_2528,N_2751);
nand UO_342 (O_342,N_2788,N_2776);
nand UO_343 (O_343,N_2803,N_2710);
nand UO_344 (O_344,N_2812,N_2562);
or UO_345 (O_345,N_2755,N_2852);
or UO_346 (O_346,N_2943,N_2974);
or UO_347 (O_347,N_2762,N_2927);
or UO_348 (O_348,N_2767,N_2893);
nor UO_349 (O_349,N_2779,N_2535);
and UO_350 (O_350,N_2894,N_2793);
nor UO_351 (O_351,N_2522,N_2733);
nand UO_352 (O_352,N_2706,N_2561);
nor UO_353 (O_353,N_2740,N_2713);
or UO_354 (O_354,N_2551,N_2747);
nor UO_355 (O_355,N_2833,N_2903);
nor UO_356 (O_356,N_2939,N_2735);
or UO_357 (O_357,N_2741,N_2846);
or UO_358 (O_358,N_2676,N_2894);
nor UO_359 (O_359,N_2588,N_2703);
and UO_360 (O_360,N_2546,N_2601);
or UO_361 (O_361,N_2539,N_2520);
nor UO_362 (O_362,N_2928,N_2610);
nand UO_363 (O_363,N_2793,N_2912);
nand UO_364 (O_364,N_2567,N_2626);
and UO_365 (O_365,N_2556,N_2714);
or UO_366 (O_366,N_2948,N_2900);
nor UO_367 (O_367,N_2522,N_2831);
nor UO_368 (O_368,N_2831,N_2747);
nand UO_369 (O_369,N_2568,N_2867);
nor UO_370 (O_370,N_2945,N_2602);
nand UO_371 (O_371,N_2664,N_2656);
or UO_372 (O_372,N_2568,N_2961);
nand UO_373 (O_373,N_2922,N_2940);
nor UO_374 (O_374,N_2555,N_2873);
xnor UO_375 (O_375,N_2833,N_2723);
and UO_376 (O_376,N_2615,N_2800);
or UO_377 (O_377,N_2641,N_2944);
or UO_378 (O_378,N_2543,N_2981);
nand UO_379 (O_379,N_2557,N_2733);
nand UO_380 (O_380,N_2917,N_2745);
nor UO_381 (O_381,N_2904,N_2846);
and UO_382 (O_382,N_2790,N_2697);
or UO_383 (O_383,N_2684,N_2977);
and UO_384 (O_384,N_2944,N_2748);
or UO_385 (O_385,N_2948,N_2970);
and UO_386 (O_386,N_2602,N_2505);
and UO_387 (O_387,N_2611,N_2521);
or UO_388 (O_388,N_2780,N_2766);
or UO_389 (O_389,N_2616,N_2868);
and UO_390 (O_390,N_2678,N_2806);
or UO_391 (O_391,N_2514,N_2549);
and UO_392 (O_392,N_2868,N_2977);
nor UO_393 (O_393,N_2627,N_2997);
or UO_394 (O_394,N_2811,N_2988);
nand UO_395 (O_395,N_2916,N_2891);
and UO_396 (O_396,N_2818,N_2503);
and UO_397 (O_397,N_2582,N_2744);
xnor UO_398 (O_398,N_2595,N_2676);
and UO_399 (O_399,N_2689,N_2686);
nor UO_400 (O_400,N_2671,N_2759);
nand UO_401 (O_401,N_2729,N_2658);
xnor UO_402 (O_402,N_2777,N_2773);
nor UO_403 (O_403,N_2570,N_2526);
and UO_404 (O_404,N_2531,N_2983);
and UO_405 (O_405,N_2994,N_2878);
nor UO_406 (O_406,N_2798,N_2709);
nor UO_407 (O_407,N_2824,N_2860);
nand UO_408 (O_408,N_2629,N_2544);
nand UO_409 (O_409,N_2955,N_2634);
and UO_410 (O_410,N_2503,N_2820);
and UO_411 (O_411,N_2564,N_2963);
and UO_412 (O_412,N_2703,N_2624);
nand UO_413 (O_413,N_2675,N_2989);
nand UO_414 (O_414,N_2539,N_2998);
or UO_415 (O_415,N_2550,N_2826);
xor UO_416 (O_416,N_2881,N_2809);
and UO_417 (O_417,N_2832,N_2938);
nor UO_418 (O_418,N_2998,N_2509);
and UO_419 (O_419,N_2891,N_2777);
or UO_420 (O_420,N_2883,N_2594);
nor UO_421 (O_421,N_2535,N_2540);
nand UO_422 (O_422,N_2791,N_2987);
nor UO_423 (O_423,N_2514,N_2819);
and UO_424 (O_424,N_2777,N_2747);
nor UO_425 (O_425,N_2937,N_2893);
xor UO_426 (O_426,N_2884,N_2891);
nor UO_427 (O_427,N_2946,N_2607);
and UO_428 (O_428,N_2859,N_2703);
nor UO_429 (O_429,N_2818,N_2819);
or UO_430 (O_430,N_2573,N_2656);
and UO_431 (O_431,N_2908,N_2682);
and UO_432 (O_432,N_2934,N_2655);
or UO_433 (O_433,N_2618,N_2620);
or UO_434 (O_434,N_2562,N_2521);
nor UO_435 (O_435,N_2519,N_2533);
or UO_436 (O_436,N_2680,N_2852);
nor UO_437 (O_437,N_2853,N_2984);
nand UO_438 (O_438,N_2931,N_2572);
or UO_439 (O_439,N_2884,N_2873);
nand UO_440 (O_440,N_2869,N_2940);
nor UO_441 (O_441,N_2788,N_2882);
nand UO_442 (O_442,N_2656,N_2912);
nand UO_443 (O_443,N_2664,N_2847);
nand UO_444 (O_444,N_2780,N_2541);
and UO_445 (O_445,N_2792,N_2998);
and UO_446 (O_446,N_2845,N_2829);
nand UO_447 (O_447,N_2901,N_2672);
nand UO_448 (O_448,N_2762,N_2846);
and UO_449 (O_449,N_2961,N_2591);
and UO_450 (O_450,N_2915,N_2863);
or UO_451 (O_451,N_2885,N_2740);
and UO_452 (O_452,N_2759,N_2591);
nor UO_453 (O_453,N_2858,N_2647);
nor UO_454 (O_454,N_2857,N_2579);
nor UO_455 (O_455,N_2812,N_2561);
xnor UO_456 (O_456,N_2653,N_2930);
or UO_457 (O_457,N_2618,N_2804);
nor UO_458 (O_458,N_2918,N_2799);
nand UO_459 (O_459,N_2516,N_2589);
nand UO_460 (O_460,N_2546,N_2621);
nor UO_461 (O_461,N_2670,N_2700);
nand UO_462 (O_462,N_2805,N_2728);
or UO_463 (O_463,N_2965,N_2763);
nand UO_464 (O_464,N_2692,N_2651);
xor UO_465 (O_465,N_2603,N_2987);
nor UO_466 (O_466,N_2949,N_2955);
or UO_467 (O_467,N_2651,N_2965);
or UO_468 (O_468,N_2539,N_2615);
nor UO_469 (O_469,N_2773,N_2807);
nor UO_470 (O_470,N_2745,N_2638);
nand UO_471 (O_471,N_2791,N_2627);
and UO_472 (O_472,N_2666,N_2658);
and UO_473 (O_473,N_2697,N_2557);
nor UO_474 (O_474,N_2664,N_2619);
nand UO_475 (O_475,N_2929,N_2758);
or UO_476 (O_476,N_2893,N_2707);
nand UO_477 (O_477,N_2858,N_2951);
nand UO_478 (O_478,N_2925,N_2704);
nand UO_479 (O_479,N_2762,N_2982);
nor UO_480 (O_480,N_2840,N_2956);
nand UO_481 (O_481,N_2582,N_2671);
or UO_482 (O_482,N_2647,N_2504);
xnor UO_483 (O_483,N_2575,N_2685);
nor UO_484 (O_484,N_2713,N_2940);
nand UO_485 (O_485,N_2697,N_2975);
nand UO_486 (O_486,N_2789,N_2878);
nand UO_487 (O_487,N_2551,N_2672);
and UO_488 (O_488,N_2959,N_2597);
nand UO_489 (O_489,N_2636,N_2737);
nor UO_490 (O_490,N_2603,N_2685);
or UO_491 (O_491,N_2784,N_2957);
nand UO_492 (O_492,N_2768,N_2832);
and UO_493 (O_493,N_2726,N_2619);
and UO_494 (O_494,N_2529,N_2954);
nor UO_495 (O_495,N_2966,N_2819);
or UO_496 (O_496,N_2635,N_2832);
or UO_497 (O_497,N_2885,N_2950);
or UO_498 (O_498,N_2638,N_2596);
and UO_499 (O_499,N_2536,N_2913);
endmodule